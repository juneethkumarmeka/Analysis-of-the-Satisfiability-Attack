module basic_1000_10000_1500_10_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_149,In_614);
nor U1 (N_1,In_530,In_164);
or U2 (N_2,In_24,In_228);
nor U3 (N_3,In_954,In_305);
nor U4 (N_4,In_907,In_984);
or U5 (N_5,In_584,In_171);
nand U6 (N_6,In_893,In_860);
and U7 (N_7,In_931,In_822);
or U8 (N_8,In_481,In_196);
nand U9 (N_9,In_669,In_901);
nor U10 (N_10,In_63,In_18);
and U11 (N_11,In_102,In_660);
and U12 (N_12,In_896,In_135);
or U13 (N_13,In_129,In_856);
and U14 (N_14,In_628,In_854);
or U15 (N_15,In_491,In_599);
and U16 (N_16,In_172,In_457);
nand U17 (N_17,In_8,In_52);
or U18 (N_18,In_520,In_683);
nor U19 (N_19,In_69,In_769);
nand U20 (N_20,In_649,In_692);
nand U21 (N_21,In_635,In_430);
and U22 (N_22,In_572,In_147);
and U23 (N_23,In_444,In_209);
nand U24 (N_24,In_809,In_106);
nand U25 (N_25,In_466,In_528);
nand U26 (N_26,In_939,In_682);
and U27 (N_27,In_296,In_990);
nand U28 (N_28,In_337,In_39);
and U29 (N_29,In_743,In_885);
and U30 (N_30,In_206,In_598);
nor U31 (N_31,In_441,In_835);
or U32 (N_32,In_301,In_630);
nor U33 (N_33,In_205,In_74);
and U34 (N_34,In_961,In_929);
or U35 (N_35,In_636,In_312);
nor U36 (N_36,In_233,In_597);
or U37 (N_37,In_420,In_492);
or U38 (N_38,In_982,In_715);
and U39 (N_39,In_125,In_637);
nand U40 (N_40,In_703,In_620);
or U41 (N_41,In_463,In_156);
nand U42 (N_42,In_389,In_718);
nand U43 (N_43,In_775,In_105);
or U44 (N_44,In_140,In_421);
nor U45 (N_45,In_184,In_807);
nor U46 (N_46,In_152,In_333);
nand U47 (N_47,In_792,In_516);
and U48 (N_48,In_243,In_714);
nand U49 (N_49,In_543,In_393);
xnor U50 (N_50,In_639,In_493);
nor U51 (N_51,In_611,In_367);
or U52 (N_52,In_864,In_552);
nand U53 (N_53,In_103,In_988);
and U54 (N_54,In_986,In_123);
or U55 (N_55,In_668,In_407);
and U56 (N_56,In_355,In_454);
nand U57 (N_57,In_532,In_522);
nand U58 (N_58,In_713,In_855);
nand U59 (N_59,In_756,In_357);
or U60 (N_60,In_851,In_542);
nand U61 (N_61,In_912,In_671);
nor U62 (N_62,In_16,In_974);
or U63 (N_63,In_585,In_943);
nand U64 (N_64,In_234,In_953);
and U65 (N_65,In_31,In_388);
or U66 (N_66,In_436,In_776);
nand U67 (N_67,In_956,In_109);
or U68 (N_68,In_398,In_307);
and U69 (N_69,In_541,In_608);
nor U70 (N_70,In_958,In_308);
or U71 (N_71,In_502,In_223);
or U72 (N_72,In_261,In_365);
and U73 (N_73,In_571,In_253);
or U74 (N_74,In_648,In_477);
nand U75 (N_75,In_181,In_558);
nor U76 (N_76,In_42,In_458);
nor U77 (N_77,In_453,In_166);
and U78 (N_78,In_664,In_179);
nand U79 (N_79,In_744,In_394);
xor U80 (N_80,In_705,In_203);
or U81 (N_81,In_804,In_903);
nand U82 (N_82,In_795,In_783);
and U83 (N_83,In_390,In_878);
nand U84 (N_84,In_922,In_936);
and U85 (N_85,In_800,In_902);
and U86 (N_86,In_198,In_805);
or U87 (N_87,In_208,In_447);
nor U88 (N_88,In_918,In_275);
nor U89 (N_89,In_136,In_399);
nor U90 (N_90,In_278,In_364);
nand U91 (N_91,In_487,In_49);
nand U92 (N_92,In_497,In_785);
nand U93 (N_93,In_60,In_68);
or U94 (N_94,In_836,In_863);
and U95 (N_95,In_403,In_495);
or U96 (N_96,In_324,In_507);
or U97 (N_97,In_448,In_122);
or U98 (N_98,In_913,In_20);
nor U99 (N_99,In_633,In_973);
xnor U100 (N_100,In_168,In_794);
nor U101 (N_101,In_554,In_494);
nand U102 (N_102,In_162,In_255);
and U103 (N_103,In_853,In_629);
nand U104 (N_104,In_935,In_29);
or U105 (N_105,In_284,In_91);
nor U106 (N_106,In_274,In_684);
nor U107 (N_107,In_595,In_460);
and U108 (N_108,In_600,In_81);
or U109 (N_109,In_753,In_86);
or U110 (N_110,In_568,In_385);
nor U111 (N_111,In_793,In_663);
nand U112 (N_112,In_348,In_590);
and U113 (N_113,In_64,In_332);
and U114 (N_114,In_362,In_229);
nor U115 (N_115,In_80,In_143);
nand U116 (N_116,In_263,In_277);
nand U117 (N_117,In_919,In_787);
and U118 (N_118,In_730,In_167);
nand U119 (N_119,In_101,In_891);
nor U120 (N_120,In_667,In_601);
nand U121 (N_121,In_376,In_881);
or U122 (N_122,In_952,In_192);
and U123 (N_123,In_911,In_915);
and U124 (N_124,In_717,In_508);
nand U125 (N_125,In_207,In_886);
nand U126 (N_126,In_248,In_183);
or U127 (N_127,In_450,In_158);
and U128 (N_128,In_725,In_659);
nand U129 (N_129,In_297,In_750);
nand U130 (N_130,In_963,In_358);
and U131 (N_131,In_720,In_655);
and U132 (N_132,In_236,In_825);
and U133 (N_133,In_574,In_99);
and U134 (N_134,In_437,In_587);
or U135 (N_135,In_578,In_265);
and U136 (N_136,In_605,In_335);
nor U137 (N_137,In_28,In_104);
and U138 (N_138,In_488,In_877);
nor U139 (N_139,In_857,In_256);
nand U140 (N_140,In_527,In_112);
xor U141 (N_141,In_127,In_279);
nand U142 (N_142,In_113,In_180);
or U143 (N_143,In_526,In_319);
nor U144 (N_144,In_338,In_440);
and U145 (N_145,In_777,In_374);
and U146 (N_146,In_216,In_700);
or U147 (N_147,In_422,In_540);
and U148 (N_148,In_439,In_626);
and U149 (N_149,In_533,In_983);
nand U150 (N_150,In_237,In_560);
or U151 (N_151,In_302,In_318);
and U152 (N_152,In_763,In_615);
and U153 (N_153,In_971,In_521);
or U154 (N_154,In_381,In_613);
or U155 (N_155,In_71,In_425);
or U156 (N_156,In_666,In_503);
and U157 (N_157,In_11,In_772);
nand U158 (N_158,In_652,In_383);
nor U159 (N_159,In_641,In_23);
or U160 (N_160,In_995,In_662);
nand U161 (N_161,In_699,In_813);
or U162 (N_162,In_992,In_197);
nor U163 (N_163,In_947,In_619);
nor U164 (N_164,In_213,In_514);
and U165 (N_165,In_645,In_309);
or U166 (N_166,In_114,In_734);
nand U167 (N_167,In_61,In_980);
or U168 (N_168,In_27,In_3);
and U169 (N_169,In_443,In_926);
and U170 (N_170,In_960,In_326);
and U171 (N_171,In_627,In_12);
or U172 (N_172,In_290,In_799);
and U173 (N_173,In_366,In_806);
or U174 (N_174,In_898,In_282);
nand U175 (N_175,In_830,In_583);
or U176 (N_176,In_375,In_691);
nand U177 (N_177,In_563,In_977);
nor U178 (N_178,In_993,In_449);
nand U179 (N_179,In_716,In_838);
xor U180 (N_180,In_250,In_33);
or U181 (N_181,In_359,In_512);
nand U182 (N_182,In_755,In_827);
nor U183 (N_183,In_538,In_757);
nand U184 (N_184,In_802,In_350);
xor U185 (N_185,In_899,In_85);
nand U186 (N_186,In_218,In_771);
and U187 (N_187,In_252,In_727);
nand U188 (N_188,In_434,In_593);
nand U189 (N_189,In_519,In_1);
or U190 (N_190,In_766,In_694);
or U191 (N_191,In_82,In_934);
or U192 (N_192,In_310,In_537);
and U193 (N_193,In_833,In_928);
xnor U194 (N_194,In_289,In_280);
nand U195 (N_195,In_764,In_246);
nand U196 (N_196,In_523,In_505);
nor U197 (N_197,In_695,In_126);
or U198 (N_198,In_410,In_191);
nor U199 (N_199,In_150,In_824);
and U200 (N_200,In_900,In_401);
nor U201 (N_201,In_97,In_557);
or U202 (N_202,In_665,In_19);
nand U203 (N_203,In_193,In_586);
or U204 (N_204,In_845,In_679);
nand U205 (N_205,In_729,In_451);
or U206 (N_206,In_948,In_876);
and U207 (N_207,In_9,In_978);
or U208 (N_208,In_151,In_550);
nand U209 (N_209,In_658,In_222);
and U210 (N_210,In_553,In_932);
or U211 (N_211,In_214,In_347);
or U212 (N_212,In_490,In_815);
nor U213 (N_213,In_698,In_72);
nand U214 (N_214,In_618,In_624);
nor U215 (N_215,In_83,In_200);
nand U216 (N_216,In_789,In_270);
nand U217 (N_217,In_842,In_178);
and U218 (N_218,In_829,In_94);
or U219 (N_219,In_489,In_589);
and U220 (N_220,In_555,In_920);
or U221 (N_221,In_174,In_621);
or U222 (N_222,In_84,In_782);
or U223 (N_223,In_14,In_832);
and U224 (N_224,In_153,In_549);
nor U225 (N_225,In_905,In_539);
nand U226 (N_226,In_124,In_416);
and U227 (N_227,In_472,In_161);
or U228 (N_228,In_821,In_165);
or U229 (N_229,In_242,In_762);
or U230 (N_230,In_404,In_696);
nand U231 (N_231,In_686,In_504);
and U232 (N_232,In_384,In_369);
or U233 (N_233,In_866,In_858);
nor U234 (N_234,In_859,In_672);
nand U235 (N_235,In_509,In_424);
and U236 (N_236,In_966,In_765);
nor U237 (N_237,In_238,In_266);
nand U238 (N_238,In_330,In_382);
or U239 (N_239,In_157,In_872);
nand U240 (N_240,In_510,In_239);
or U241 (N_241,In_921,In_742);
nor U242 (N_242,In_176,In_603);
or U243 (N_243,In_862,In_498);
or U244 (N_244,In_622,In_117);
nor U245 (N_245,In_499,In_796);
or U246 (N_246,In_10,In_336);
nor U247 (N_247,In_26,In_739);
and U248 (N_248,In_774,In_803);
nand U249 (N_249,In_66,In_464);
nor U250 (N_250,In_461,In_368);
nand U251 (N_251,In_610,In_433);
and U252 (N_252,In_144,In_475);
nor U253 (N_253,In_93,In_220);
nor U254 (N_254,In_767,In_428);
or U255 (N_255,In_107,In_303);
nor U256 (N_256,In_873,In_646);
nor U257 (N_257,In_445,In_90);
nor U258 (N_258,In_689,In_941);
and U259 (N_259,In_861,In_708);
nor U260 (N_260,In_96,In_40);
and U261 (N_261,In_733,In_43);
or U262 (N_262,In_25,In_271);
or U263 (N_263,In_260,In_264);
nand U264 (N_264,In_210,In_67);
nor U265 (N_265,In_139,In_146);
and U266 (N_266,In_592,In_987);
and U267 (N_267,In_15,In_311);
and U268 (N_268,In_741,In_397);
nor U269 (N_269,In_868,In_173);
nor U270 (N_270,In_778,In_98);
nor U271 (N_271,In_132,In_917);
nand U272 (N_272,In_710,In_647);
nor U273 (N_273,In_951,In_247);
and U274 (N_274,In_844,In_726);
nand U275 (N_275,In_643,In_75);
nor U276 (N_276,In_945,In_21);
nor U277 (N_277,In_221,In_894);
and U278 (N_278,In_712,In_955);
nand U279 (N_279,In_235,In_746);
nor U280 (N_280,In_638,In_678);
nor U281 (N_281,In_47,In_329);
or U282 (N_282,In_352,In_968);
nand U283 (N_283,In_480,In_534);
or U284 (N_284,In_199,In_906);
nor U285 (N_285,In_291,In_596);
nand U286 (N_286,In_134,In_511);
nand U287 (N_287,In_426,In_267);
and U288 (N_288,In_298,In_834);
or U289 (N_289,In_41,In_219);
and U290 (N_290,In_989,In_414);
nor U291 (N_291,In_916,In_13);
nand U292 (N_292,In_65,In_950);
or U293 (N_293,In_227,In_59);
and U294 (N_294,In_892,In_848);
or U295 (N_295,In_887,In_115);
or U296 (N_296,In_56,In_964);
nand U297 (N_297,In_418,In_354);
and U298 (N_298,In_930,In_969);
or U299 (N_299,In_865,In_690);
nand U300 (N_300,In_616,In_651);
or U301 (N_301,In_379,In_732);
and U302 (N_302,In_650,In_92);
nand U303 (N_303,In_288,In_339);
and U304 (N_304,In_790,In_251);
or U305 (N_305,In_287,In_138);
nand U306 (N_306,In_575,In_343);
or U307 (N_307,In_631,In_500);
or U308 (N_308,In_602,In_957);
or U309 (N_309,In_561,In_53);
or U310 (N_310,In_736,In_702);
nand U311 (N_311,In_100,In_285);
nand U312 (N_312,In_496,In_131);
nor U313 (N_313,In_44,In_882);
or U314 (N_314,In_293,In_925);
or U315 (N_315,In_476,In_531);
nor U316 (N_316,In_826,In_723);
and U317 (N_317,In_812,In_231);
xor U318 (N_318,In_54,In_545);
or U319 (N_319,In_979,In_190);
and U320 (N_320,In_642,In_780);
nor U321 (N_321,In_37,In_32);
or U322 (N_322,In_914,In_116);
or U323 (N_323,In_429,In_45);
or U324 (N_324,In_320,In_76);
nor U325 (N_325,In_640,In_607);
or U326 (N_326,In_95,In_870);
and U327 (N_327,In_985,In_245);
or U328 (N_328,In_897,In_442);
and U329 (N_329,In_852,In_120);
or U330 (N_330,In_536,In_580);
nand U331 (N_331,In_283,In_788);
or U332 (N_332,In_268,In_770);
nand U333 (N_333,In_972,In_761);
and U334 (N_334,In_976,In_991);
nor U335 (N_335,In_300,In_784);
or U336 (N_336,In_850,In_272);
nand U337 (N_337,In_411,In_680);
nand U338 (N_338,In_944,In_387);
nor U339 (N_339,In_908,In_465);
nand U340 (N_340,In_130,In_604);
or U341 (N_341,In_58,In_748);
nand U342 (N_342,In_483,In_749);
nor U343 (N_343,In_36,In_353);
nand U344 (N_344,In_34,In_693);
or U345 (N_345,In_371,In_315);
nor U346 (N_346,In_632,In_577);
or U347 (N_347,In_820,In_341);
and U348 (N_348,In_996,In_340);
nand U349 (N_349,In_840,In_241);
or U350 (N_350,In_17,In_110);
nor U351 (N_351,In_469,In_159);
or U352 (N_352,In_412,In_547);
or U353 (N_353,In_625,In_808);
or U354 (N_354,In_721,In_467);
nand U355 (N_355,In_435,In_73);
or U356 (N_356,In_513,In_525);
nand U357 (N_357,In_321,In_269);
nand U358 (N_358,In_155,In_924);
and U359 (N_359,In_372,In_257);
nor U360 (N_360,In_759,In_569);
or U361 (N_361,In_728,In_189);
nand U362 (N_362,In_344,In_517);
nand U363 (N_363,In_940,In_738);
or U364 (N_364,In_653,In_35);
and U365 (N_365,In_111,In_688);
nand U366 (N_366,In_6,In_760);
and U367 (N_367,In_810,In_51);
or U368 (N_368,In_46,In_349);
and U369 (N_369,In_0,In_259);
or U370 (N_370,In_923,In_431);
and U371 (N_371,In_828,In_323);
nor U372 (N_372,In_841,In_506);
or U373 (N_373,In_927,In_754);
nor U374 (N_374,In_768,In_276);
and U375 (N_375,In_798,In_673);
nand U376 (N_376,In_195,In_997);
nor U377 (N_377,In_758,In_392);
nand U378 (N_378,In_316,In_406);
nand U379 (N_379,In_215,In_304);
nor U380 (N_380,In_551,In_169);
nand U381 (N_381,In_562,In_87);
and U382 (N_382,In_281,In_817);
nor U383 (N_383,In_831,In_185);
nand U384 (N_384,In_262,In_588);
and U385 (N_385,In_459,In_704);
or U386 (N_386,In_378,In_363);
nor U387 (N_387,In_108,In_89);
nor U388 (N_388,In_322,In_62);
nand U389 (N_389,In_370,In_128);
nor U390 (N_390,In_731,In_142);
and U391 (N_391,In_623,In_949);
and U392 (N_392,In_823,In_524);
or U393 (N_393,In_202,In_186);
nand U394 (N_394,In_701,In_942);
and U395 (N_395,In_88,In_994);
and U396 (N_396,In_141,In_470);
or U397 (N_397,In_473,In_160);
and U398 (N_398,In_773,In_573);
nand U399 (N_399,In_871,In_456);
nor U400 (N_400,In_719,In_438);
and U401 (N_401,In_423,In_306);
and U402 (N_402,In_292,In_249);
nor U403 (N_403,In_462,In_880);
and U404 (N_404,In_468,In_360);
and U405 (N_405,In_79,In_582);
and U406 (N_406,In_559,In_327);
nor U407 (N_407,In_965,In_970);
or U408 (N_408,In_819,In_119);
or U409 (N_409,In_634,In_188);
or U410 (N_410,In_417,In_361);
nor U411 (N_411,In_328,In_334);
or U412 (N_412,In_849,In_975);
nand U413 (N_413,In_224,In_38);
nor U414 (N_414,In_471,In_544);
nor U415 (N_415,In_377,In_345);
nand U416 (N_416,In_883,In_546);
nand U417 (N_417,In_240,In_515);
xnor U418 (N_418,In_654,In_879);
xor U419 (N_419,In_194,In_452);
nor U420 (N_420,In_485,In_843);
and U421 (N_421,In_751,In_211);
xor U422 (N_422,In_846,In_967);
and U423 (N_423,In_867,In_484);
and U424 (N_424,In_446,In_875);
and U425 (N_425,In_201,In_837);
nor U426 (N_426,In_391,In_182);
and U427 (N_427,In_687,In_286);
or U428 (N_428,In_386,In_325);
nor U429 (N_429,In_175,In_317);
nand U430 (N_430,In_501,In_874);
nand U431 (N_431,In_30,In_888);
nand U432 (N_432,In_740,In_869);
nand U433 (N_433,In_722,In_230);
or U434 (N_434,In_212,In_591);
nor U435 (N_435,In_644,In_427);
or U436 (N_436,In_22,In_656);
or U437 (N_437,In_709,In_938);
nor U438 (N_438,In_617,In_7);
or U439 (N_439,In_606,In_55);
nor U440 (N_440,In_737,In_711);
nand U441 (N_441,In_413,In_244);
nor U442 (N_442,In_594,In_818);
or U443 (N_443,In_779,In_847);
nor U444 (N_444,In_154,In_295);
nor U445 (N_445,In_797,In_294);
and U446 (N_446,In_373,In_217);
nor U447 (N_447,In_814,In_946);
nor U448 (N_448,In_409,In_258);
nand U449 (N_449,In_890,In_674);
nor U450 (N_450,In_889,In_981);
or U451 (N_451,In_675,In_752);
or U452 (N_452,In_380,In_565);
and U453 (N_453,In_676,In_5);
or U454 (N_454,In_474,In_118);
nor U455 (N_455,In_884,In_609);
or U456 (N_456,In_77,In_170);
or U457 (N_457,In_148,In_657);
and U458 (N_458,In_351,In_791);
and U459 (N_459,In_478,In_356);
or U460 (N_460,In_581,In_518);
and U461 (N_461,In_400,In_342);
nor U462 (N_462,In_402,In_204);
nand U463 (N_463,In_415,In_163);
nand U464 (N_464,In_408,In_910);
nand U465 (N_465,In_811,In_681);
nand U466 (N_466,In_564,In_962);
and U467 (N_467,In_959,In_816);
nor U468 (N_468,In_801,In_677);
and U469 (N_469,In_482,In_697);
or U470 (N_470,In_839,In_4);
nor U471 (N_471,In_225,In_566);
nand U472 (N_472,In_232,In_904);
and U473 (N_473,In_670,In_2);
nor U474 (N_474,In_707,In_937);
and U475 (N_475,In_786,In_48);
nand U476 (N_476,In_535,In_314);
nor U477 (N_477,In_909,In_177);
and U478 (N_478,In_70,In_121);
and U479 (N_479,In_57,In_486);
and U480 (N_480,In_313,In_556);
nor U481 (N_481,In_432,In_548);
and U482 (N_482,In_145,In_998);
nor U483 (N_483,In_529,In_273);
and U484 (N_484,In_395,In_479);
or U485 (N_485,In_781,In_396);
or U486 (N_486,In_579,In_137);
nand U487 (N_487,In_895,In_745);
and U488 (N_488,In_735,In_187);
or U489 (N_489,In_346,In_747);
nand U490 (N_490,In_133,In_661);
and U491 (N_491,In_999,In_50);
or U492 (N_492,In_419,In_567);
nor U493 (N_493,In_254,In_706);
or U494 (N_494,In_685,In_226);
nor U495 (N_495,In_570,In_724);
or U496 (N_496,In_576,In_331);
and U497 (N_497,In_933,In_78);
or U498 (N_498,In_612,In_455);
and U499 (N_499,In_299,In_405);
nand U500 (N_500,In_483,In_611);
nand U501 (N_501,In_743,In_397);
or U502 (N_502,In_239,In_808);
nor U503 (N_503,In_567,In_188);
nand U504 (N_504,In_419,In_267);
nor U505 (N_505,In_122,In_821);
or U506 (N_506,In_137,In_72);
and U507 (N_507,In_598,In_587);
nand U508 (N_508,In_463,In_312);
nand U509 (N_509,In_941,In_976);
nand U510 (N_510,In_301,In_231);
or U511 (N_511,In_743,In_859);
or U512 (N_512,In_956,In_963);
xor U513 (N_513,In_754,In_921);
nand U514 (N_514,In_948,In_22);
nand U515 (N_515,In_132,In_683);
nand U516 (N_516,In_793,In_973);
nand U517 (N_517,In_455,In_465);
or U518 (N_518,In_549,In_534);
or U519 (N_519,In_741,In_325);
nor U520 (N_520,In_630,In_714);
and U521 (N_521,In_375,In_820);
nor U522 (N_522,In_564,In_687);
nand U523 (N_523,In_293,In_146);
or U524 (N_524,In_897,In_242);
or U525 (N_525,In_638,In_109);
and U526 (N_526,In_272,In_569);
and U527 (N_527,In_7,In_864);
or U528 (N_528,In_21,In_518);
nor U529 (N_529,In_277,In_680);
nand U530 (N_530,In_824,In_850);
nand U531 (N_531,In_888,In_81);
and U532 (N_532,In_5,In_959);
xnor U533 (N_533,In_430,In_644);
nand U534 (N_534,In_96,In_424);
nand U535 (N_535,In_917,In_316);
and U536 (N_536,In_346,In_908);
nor U537 (N_537,In_764,In_893);
or U538 (N_538,In_49,In_177);
or U539 (N_539,In_892,In_898);
nor U540 (N_540,In_481,In_441);
or U541 (N_541,In_418,In_83);
nor U542 (N_542,In_898,In_614);
nand U543 (N_543,In_300,In_930);
nor U544 (N_544,In_46,In_928);
nand U545 (N_545,In_888,In_950);
and U546 (N_546,In_191,In_679);
or U547 (N_547,In_575,In_150);
nand U548 (N_548,In_553,In_315);
xnor U549 (N_549,In_131,In_43);
or U550 (N_550,In_518,In_522);
nand U551 (N_551,In_577,In_406);
and U552 (N_552,In_225,In_943);
nand U553 (N_553,In_384,In_461);
and U554 (N_554,In_482,In_65);
and U555 (N_555,In_146,In_575);
nor U556 (N_556,In_352,In_60);
nor U557 (N_557,In_426,In_671);
and U558 (N_558,In_874,In_69);
or U559 (N_559,In_642,In_711);
xor U560 (N_560,In_638,In_428);
nand U561 (N_561,In_445,In_174);
xnor U562 (N_562,In_580,In_50);
nand U563 (N_563,In_287,In_866);
nand U564 (N_564,In_503,In_140);
and U565 (N_565,In_937,In_649);
nor U566 (N_566,In_844,In_207);
or U567 (N_567,In_49,In_913);
nor U568 (N_568,In_451,In_321);
nor U569 (N_569,In_447,In_775);
or U570 (N_570,In_979,In_2);
nor U571 (N_571,In_616,In_113);
nand U572 (N_572,In_995,In_932);
nand U573 (N_573,In_138,In_659);
or U574 (N_574,In_442,In_617);
or U575 (N_575,In_791,In_595);
nor U576 (N_576,In_23,In_784);
or U577 (N_577,In_177,In_445);
or U578 (N_578,In_420,In_630);
and U579 (N_579,In_595,In_752);
or U580 (N_580,In_889,In_843);
nor U581 (N_581,In_79,In_339);
or U582 (N_582,In_177,In_682);
nand U583 (N_583,In_616,In_632);
nor U584 (N_584,In_364,In_195);
or U585 (N_585,In_25,In_761);
and U586 (N_586,In_543,In_528);
xor U587 (N_587,In_48,In_716);
nand U588 (N_588,In_356,In_922);
or U589 (N_589,In_614,In_699);
nor U590 (N_590,In_605,In_982);
and U591 (N_591,In_690,In_768);
nand U592 (N_592,In_338,In_704);
nor U593 (N_593,In_368,In_217);
nand U594 (N_594,In_916,In_2);
and U595 (N_595,In_231,In_347);
and U596 (N_596,In_87,In_176);
nor U597 (N_597,In_973,In_810);
nand U598 (N_598,In_186,In_997);
or U599 (N_599,In_367,In_823);
nand U600 (N_600,In_622,In_244);
nand U601 (N_601,In_650,In_358);
and U602 (N_602,In_186,In_914);
nand U603 (N_603,In_852,In_135);
nand U604 (N_604,In_610,In_683);
nand U605 (N_605,In_667,In_895);
and U606 (N_606,In_202,In_699);
or U607 (N_607,In_367,In_331);
nor U608 (N_608,In_119,In_163);
and U609 (N_609,In_22,In_170);
xor U610 (N_610,In_843,In_719);
nor U611 (N_611,In_457,In_964);
or U612 (N_612,In_499,In_508);
nor U613 (N_613,In_81,In_981);
nor U614 (N_614,In_526,In_828);
nand U615 (N_615,In_677,In_281);
and U616 (N_616,In_533,In_685);
and U617 (N_617,In_716,In_552);
and U618 (N_618,In_160,In_691);
nand U619 (N_619,In_777,In_409);
or U620 (N_620,In_800,In_86);
nand U621 (N_621,In_817,In_192);
nand U622 (N_622,In_42,In_87);
and U623 (N_623,In_479,In_962);
or U624 (N_624,In_797,In_828);
or U625 (N_625,In_355,In_157);
nand U626 (N_626,In_795,In_396);
nand U627 (N_627,In_521,In_816);
nor U628 (N_628,In_486,In_252);
nand U629 (N_629,In_295,In_275);
nor U630 (N_630,In_436,In_549);
nand U631 (N_631,In_800,In_418);
and U632 (N_632,In_904,In_671);
nor U633 (N_633,In_679,In_397);
or U634 (N_634,In_767,In_572);
nor U635 (N_635,In_814,In_398);
and U636 (N_636,In_656,In_916);
and U637 (N_637,In_391,In_295);
nor U638 (N_638,In_51,In_71);
or U639 (N_639,In_573,In_537);
or U640 (N_640,In_153,In_997);
and U641 (N_641,In_475,In_318);
and U642 (N_642,In_414,In_126);
and U643 (N_643,In_704,In_916);
nand U644 (N_644,In_950,In_153);
and U645 (N_645,In_165,In_304);
nor U646 (N_646,In_715,In_264);
and U647 (N_647,In_384,In_290);
and U648 (N_648,In_465,In_806);
nand U649 (N_649,In_747,In_472);
or U650 (N_650,In_680,In_767);
nand U651 (N_651,In_393,In_74);
and U652 (N_652,In_687,In_60);
and U653 (N_653,In_843,In_861);
or U654 (N_654,In_334,In_206);
or U655 (N_655,In_313,In_204);
nor U656 (N_656,In_889,In_709);
or U657 (N_657,In_424,In_196);
nor U658 (N_658,In_503,In_112);
nor U659 (N_659,In_931,In_982);
and U660 (N_660,In_515,In_203);
and U661 (N_661,In_301,In_482);
and U662 (N_662,In_718,In_478);
nand U663 (N_663,In_517,In_661);
or U664 (N_664,In_946,In_987);
and U665 (N_665,In_487,In_517);
and U666 (N_666,In_599,In_38);
nor U667 (N_667,In_475,In_416);
nor U668 (N_668,In_723,In_150);
or U669 (N_669,In_975,In_611);
nand U670 (N_670,In_398,In_402);
and U671 (N_671,In_819,In_167);
nand U672 (N_672,In_512,In_616);
nor U673 (N_673,In_976,In_391);
nand U674 (N_674,In_106,In_602);
nor U675 (N_675,In_731,In_514);
and U676 (N_676,In_318,In_295);
and U677 (N_677,In_632,In_459);
or U678 (N_678,In_60,In_469);
and U679 (N_679,In_159,In_919);
or U680 (N_680,In_764,In_345);
nor U681 (N_681,In_502,In_186);
and U682 (N_682,In_217,In_383);
nor U683 (N_683,In_36,In_240);
nand U684 (N_684,In_143,In_730);
nor U685 (N_685,In_984,In_990);
or U686 (N_686,In_879,In_18);
and U687 (N_687,In_626,In_358);
or U688 (N_688,In_393,In_126);
nand U689 (N_689,In_80,In_586);
nand U690 (N_690,In_262,In_155);
and U691 (N_691,In_78,In_87);
and U692 (N_692,In_413,In_979);
nor U693 (N_693,In_961,In_778);
nand U694 (N_694,In_140,In_602);
and U695 (N_695,In_507,In_95);
or U696 (N_696,In_697,In_526);
nor U697 (N_697,In_423,In_206);
or U698 (N_698,In_771,In_948);
and U699 (N_699,In_755,In_375);
or U700 (N_700,In_832,In_390);
nor U701 (N_701,In_141,In_754);
nand U702 (N_702,In_706,In_172);
and U703 (N_703,In_75,In_996);
nor U704 (N_704,In_778,In_208);
nor U705 (N_705,In_302,In_674);
nor U706 (N_706,In_600,In_816);
or U707 (N_707,In_831,In_923);
and U708 (N_708,In_227,In_127);
or U709 (N_709,In_311,In_116);
nand U710 (N_710,In_677,In_416);
or U711 (N_711,In_599,In_402);
or U712 (N_712,In_207,In_868);
or U713 (N_713,In_644,In_520);
xnor U714 (N_714,In_822,In_433);
and U715 (N_715,In_417,In_621);
or U716 (N_716,In_737,In_508);
or U717 (N_717,In_203,In_308);
and U718 (N_718,In_828,In_270);
or U719 (N_719,In_688,In_667);
nand U720 (N_720,In_652,In_440);
nor U721 (N_721,In_844,In_863);
and U722 (N_722,In_45,In_22);
nand U723 (N_723,In_244,In_158);
nand U724 (N_724,In_147,In_450);
nand U725 (N_725,In_186,In_937);
nor U726 (N_726,In_994,In_597);
nand U727 (N_727,In_75,In_827);
and U728 (N_728,In_2,In_478);
and U729 (N_729,In_579,In_298);
nand U730 (N_730,In_574,In_636);
nand U731 (N_731,In_295,In_942);
or U732 (N_732,In_952,In_719);
or U733 (N_733,In_224,In_440);
and U734 (N_734,In_80,In_961);
or U735 (N_735,In_232,In_774);
or U736 (N_736,In_32,In_127);
or U737 (N_737,In_553,In_35);
nor U738 (N_738,In_135,In_475);
and U739 (N_739,In_283,In_416);
nand U740 (N_740,In_464,In_310);
and U741 (N_741,In_798,In_491);
nor U742 (N_742,In_845,In_810);
and U743 (N_743,In_83,In_478);
and U744 (N_744,In_223,In_468);
and U745 (N_745,In_167,In_869);
or U746 (N_746,In_575,In_394);
or U747 (N_747,In_39,In_52);
nand U748 (N_748,In_991,In_179);
and U749 (N_749,In_723,In_204);
and U750 (N_750,In_750,In_687);
and U751 (N_751,In_796,In_20);
nand U752 (N_752,In_379,In_313);
nand U753 (N_753,In_655,In_641);
and U754 (N_754,In_600,In_648);
and U755 (N_755,In_640,In_611);
and U756 (N_756,In_706,In_435);
nand U757 (N_757,In_603,In_881);
nand U758 (N_758,In_233,In_850);
and U759 (N_759,In_223,In_357);
and U760 (N_760,In_509,In_87);
nand U761 (N_761,In_445,In_561);
nor U762 (N_762,In_881,In_573);
nand U763 (N_763,In_332,In_789);
nor U764 (N_764,In_430,In_207);
or U765 (N_765,In_756,In_269);
nor U766 (N_766,In_888,In_491);
nand U767 (N_767,In_605,In_367);
or U768 (N_768,In_73,In_330);
and U769 (N_769,In_743,In_440);
or U770 (N_770,In_494,In_683);
nor U771 (N_771,In_782,In_961);
nand U772 (N_772,In_652,In_673);
nor U773 (N_773,In_152,In_545);
nand U774 (N_774,In_54,In_847);
nor U775 (N_775,In_489,In_102);
and U776 (N_776,In_149,In_848);
or U777 (N_777,In_99,In_321);
and U778 (N_778,In_316,In_308);
nand U779 (N_779,In_182,In_631);
nand U780 (N_780,In_478,In_954);
and U781 (N_781,In_740,In_108);
nor U782 (N_782,In_536,In_18);
nand U783 (N_783,In_346,In_27);
or U784 (N_784,In_808,In_997);
nor U785 (N_785,In_376,In_340);
nor U786 (N_786,In_203,In_904);
and U787 (N_787,In_611,In_143);
nand U788 (N_788,In_475,In_302);
or U789 (N_789,In_685,In_192);
xnor U790 (N_790,In_453,In_640);
nand U791 (N_791,In_306,In_329);
and U792 (N_792,In_188,In_462);
nor U793 (N_793,In_462,In_534);
nor U794 (N_794,In_728,In_364);
and U795 (N_795,In_392,In_720);
and U796 (N_796,In_794,In_542);
nor U797 (N_797,In_615,In_977);
or U798 (N_798,In_493,In_541);
and U799 (N_799,In_583,In_87);
nand U800 (N_800,In_159,In_96);
or U801 (N_801,In_444,In_464);
or U802 (N_802,In_656,In_409);
and U803 (N_803,In_18,In_574);
and U804 (N_804,In_200,In_0);
or U805 (N_805,In_460,In_449);
nand U806 (N_806,In_134,In_904);
and U807 (N_807,In_306,In_969);
and U808 (N_808,In_521,In_941);
nand U809 (N_809,In_497,In_939);
nor U810 (N_810,In_852,In_409);
xnor U811 (N_811,In_299,In_463);
nor U812 (N_812,In_542,In_979);
or U813 (N_813,In_377,In_620);
nand U814 (N_814,In_725,In_323);
nand U815 (N_815,In_577,In_834);
and U816 (N_816,In_737,In_206);
and U817 (N_817,In_875,In_697);
nor U818 (N_818,In_231,In_248);
and U819 (N_819,In_64,In_835);
nor U820 (N_820,In_64,In_475);
and U821 (N_821,In_273,In_230);
nor U822 (N_822,In_503,In_500);
or U823 (N_823,In_981,In_130);
nand U824 (N_824,In_214,In_983);
and U825 (N_825,In_471,In_896);
and U826 (N_826,In_116,In_114);
nor U827 (N_827,In_101,In_515);
or U828 (N_828,In_116,In_476);
and U829 (N_829,In_141,In_694);
or U830 (N_830,In_473,In_522);
or U831 (N_831,In_396,In_304);
nand U832 (N_832,In_670,In_664);
or U833 (N_833,In_261,In_181);
nor U834 (N_834,In_794,In_380);
nor U835 (N_835,In_977,In_197);
nand U836 (N_836,In_836,In_462);
nand U837 (N_837,In_198,In_715);
or U838 (N_838,In_110,In_858);
nor U839 (N_839,In_256,In_626);
nor U840 (N_840,In_816,In_870);
nand U841 (N_841,In_689,In_676);
or U842 (N_842,In_768,In_221);
or U843 (N_843,In_679,In_142);
and U844 (N_844,In_106,In_194);
and U845 (N_845,In_561,In_774);
or U846 (N_846,In_464,In_546);
nand U847 (N_847,In_711,In_2);
or U848 (N_848,In_468,In_797);
nand U849 (N_849,In_994,In_538);
or U850 (N_850,In_918,In_120);
nand U851 (N_851,In_718,In_331);
nand U852 (N_852,In_496,In_754);
nor U853 (N_853,In_167,In_281);
nor U854 (N_854,In_559,In_677);
nand U855 (N_855,In_68,In_285);
and U856 (N_856,In_247,In_487);
nor U857 (N_857,In_787,In_813);
and U858 (N_858,In_709,In_870);
or U859 (N_859,In_640,In_275);
or U860 (N_860,In_155,In_712);
and U861 (N_861,In_519,In_427);
and U862 (N_862,In_658,In_904);
and U863 (N_863,In_75,In_911);
nand U864 (N_864,In_405,In_513);
or U865 (N_865,In_670,In_46);
and U866 (N_866,In_597,In_345);
nand U867 (N_867,In_209,In_962);
nand U868 (N_868,In_514,In_636);
or U869 (N_869,In_27,In_672);
or U870 (N_870,In_855,In_616);
nor U871 (N_871,In_950,In_159);
nand U872 (N_872,In_179,In_994);
and U873 (N_873,In_355,In_620);
nor U874 (N_874,In_472,In_860);
nor U875 (N_875,In_963,In_46);
and U876 (N_876,In_548,In_519);
nor U877 (N_877,In_24,In_49);
nor U878 (N_878,In_746,In_742);
or U879 (N_879,In_131,In_338);
and U880 (N_880,In_0,In_4);
nand U881 (N_881,In_448,In_858);
nor U882 (N_882,In_82,In_774);
nand U883 (N_883,In_988,In_440);
or U884 (N_884,In_211,In_716);
nor U885 (N_885,In_110,In_670);
or U886 (N_886,In_69,In_936);
and U887 (N_887,In_840,In_919);
nor U888 (N_888,In_705,In_259);
nand U889 (N_889,In_802,In_320);
nor U890 (N_890,In_549,In_127);
or U891 (N_891,In_647,In_670);
nand U892 (N_892,In_679,In_434);
and U893 (N_893,In_317,In_571);
and U894 (N_894,In_152,In_929);
nor U895 (N_895,In_424,In_447);
nor U896 (N_896,In_88,In_872);
and U897 (N_897,In_227,In_947);
and U898 (N_898,In_355,In_349);
and U899 (N_899,In_512,In_821);
or U900 (N_900,In_836,In_801);
and U901 (N_901,In_231,In_792);
or U902 (N_902,In_530,In_464);
and U903 (N_903,In_801,In_714);
and U904 (N_904,In_3,In_182);
nand U905 (N_905,In_308,In_21);
nor U906 (N_906,In_695,In_615);
nand U907 (N_907,In_676,In_356);
nand U908 (N_908,In_494,In_285);
nand U909 (N_909,In_330,In_831);
nand U910 (N_910,In_193,In_452);
nand U911 (N_911,In_670,In_401);
nand U912 (N_912,In_215,In_588);
nor U913 (N_913,In_659,In_621);
nor U914 (N_914,In_792,In_618);
and U915 (N_915,In_533,In_688);
nand U916 (N_916,In_855,In_770);
nand U917 (N_917,In_341,In_666);
nor U918 (N_918,In_285,In_956);
nand U919 (N_919,In_874,In_34);
nor U920 (N_920,In_64,In_772);
and U921 (N_921,In_986,In_106);
and U922 (N_922,In_531,In_872);
or U923 (N_923,In_670,In_507);
or U924 (N_924,In_483,In_571);
and U925 (N_925,In_28,In_425);
nand U926 (N_926,In_222,In_867);
or U927 (N_927,In_172,In_467);
and U928 (N_928,In_263,In_433);
and U929 (N_929,In_446,In_582);
nand U930 (N_930,In_581,In_345);
or U931 (N_931,In_62,In_736);
and U932 (N_932,In_123,In_636);
nor U933 (N_933,In_521,In_298);
nand U934 (N_934,In_735,In_933);
and U935 (N_935,In_904,In_613);
nor U936 (N_936,In_801,In_698);
or U937 (N_937,In_349,In_921);
or U938 (N_938,In_334,In_547);
or U939 (N_939,In_465,In_960);
and U940 (N_940,In_341,In_19);
or U941 (N_941,In_362,In_684);
nand U942 (N_942,In_323,In_986);
nand U943 (N_943,In_244,In_399);
and U944 (N_944,In_923,In_799);
xor U945 (N_945,In_934,In_983);
nand U946 (N_946,In_160,In_289);
and U947 (N_947,In_46,In_84);
and U948 (N_948,In_407,In_893);
and U949 (N_949,In_643,In_107);
nor U950 (N_950,In_757,In_838);
nor U951 (N_951,In_63,In_457);
nand U952 (N_952,In_121,In_815);
or U953 (N_953,In_795,In_921);
nor U954 (N_954,In_672,In_440);
nor U955 (N_955,In_310,In_11);
nor U956 (N_956,In_613,In_814);
or U957 (N_957,In_964,In_154);
and U958 (N_958,In_556,In_912);
and U959 (N_959,In_163,In_95);
or U960 (N_960,In_987,In_943);
and U961 (N_961,In_995,In_905);
and U962 (N_962,In_657,In_244);
nor U963 (N_963,In_758,In_423);
nand U964 (N_964,In_423,In_661);
or U965 (N_965,In_272,In_860);
nor U966 (N_966,In_431,In_114);
nand U967 (N_967,In_464,In_747);
and U968 (N_968,In_149,In_62);
nor U969 (N_969,In_664,In_974);
nand U970 (N_970,In_832,In_227);
nor U971 (N_971,In_59,In_104);
nand U972 (N_972,In_476,In_834);
and U973 (N_973,In_154,In_322);
or U974 (N_974,In_44,In_113);
or U975 (N_975,In_571,In_465);
nor U976 (N_976,In_948,In_476);
nand U977 (N_977,In_809,In_166);
and U978 (N_978,In_934,In_358);
or U979 (N_979,In_784,In_551);
or U980 (N_980,In_419,In_387);
or U981 (N_981,In_628,In_713);
nand U982 (N_982,In_778,In_995);
nand U983 (N_983,In_941,In_361);
or U984 (N_984,In_74,In_660);
and U985 (N_985,In_163,In_344);
nor U986 (N_986,In_919,In_132);
and U987 (N_987,In_652,In_979);
and U988 (N_988,In_657,In_222);
and U989 (N_989,In_309,In_854);
and U990 (N_990,In_194,In_193);
and U991 (N_991,In_853,In_674);
or U992 (N_992,In_866,In_760);
and U993 (N_993,In_445,In_133);
nor U994 (N_994,In_756,In_171);
nand U995 (N_995,In_743,In_1);
nor U996 (N_996,In_480,In_447);
and U997 (N_997,In_554,In_211);
nand U998 (N_998,In_864,In_565);
or U999 (N_999,In_49,In_698);
and U1000 (N_1000,N_246,N_405);
and U1001 (N_1001,N_181,N_262);
nor U1002 (N_1002,N_212,N_614);
and U1003 (N_1003,N_373,N_433);
and U1004 (N_1004,N_970,N_680);
nor U1005 (N_1005,N_389,N_860);
and U1006 (N_1006,N_504,N_741);
nand U1007 (N_1007,N_498,N_626);
and U1008 (N_1008,N_320,N_382);
nand U1009 (N_1009,N_79,N_134);
or U1010 (N_1010,N_146,N_50);
nor U1011 (N_1011,N_829,N_166);
and U1012 (N_1012,N_426,N_378);
or U1013 (N_1013,N_334,N_75);
and U1014 (N_1014,N_862,N_818);
or U1015 (N_1015,N_623,N_419);
xor U1016 (N_1016,N_423,N_745);
or U1017 (N_1017,N_38,N_497);
nor U1018 (N_1018,N_179,N_150);
or U1019 (N_1019,N_210,N_324);
and U1020 (N_1020,N_797,N_70);
and U1021 (N_1021,N_448,N_951);
nand U1022 (N_1022,N_94,N_314);
and U1023 (N_1023,N_335,N_697);
and U1024 (N_1024,N_774,N_330);
and U1025 (N_1025,N_625,N_55);
and U1026 (N_1026,N_294,N_587);
and U1027 (N_1027,N_293,N_435);
or U1028 (N_1028,N_197,N_113);
and U1029 (N_1029,N_71,N_783);
nand U1030 (N_1030,N_615,N_726);
and U1031 (N_1031,N_450,N_515);
nor U1032 (N_1032,N_949,N_296);
and U1033 (N_1033,N_944,N_112);
or U1034 (N_1034,N_861,N_41);
nand U1035 (N_1035,N_182,N_612);
nand U1036 (N_1036,N_718,N_821);
nor U1037 (N_1037,N_369,N_830);
and U1038 (N_1038,N_201,N_183);
nand U1039 (N_1039,N_743,N_310);
or U1040 (N_1040,N_388,N_586);
or U1041 (N_1041,N_319,N_813);
nand U1042 (N_1042,N_239,N_957);
or U1043 (N_1043,N_338,N_863);
nand U1044 (N_1044,N_39,N_82);
nand U1045 (N_1045,N_922,N_493);
and U1046 (N_1046,N_795,N_888);
nor U1047 (N_1047,N_375,N_751);
nand U1048 (N_1048,N_43,N_844);
and U1049 (N_1049,N_540,N_896);
and U1050 (N_1050,N_152,N_171);
nand U1051 (N_1051,N_479,N_880);
and U1052 (N_1052,N_823,N_29);
and U1053 (N_1053,N_557,N_424);
or U1054 (N_1054,N_732,N_403);
and U1055 (N_1055,N_693,N_740);
or U1056 (N_1056,N_617,N_509);
or U1057 (N_1057,N_337,N_907);
nand U1058 (N_1058,N_824,N_354);
and U1059 (N_1059,N_366,N_139);
and U1060 (N_1060,N_675,N_108);
or U1061 (N_1061,N_787,N_281);
nor U1062 (N_1062,N_577,N_782);
nor U1063 (N_1063,N_431,N_123);
nand U1064 (N_1064,N_621,N_464);
or U1065 (N_1065,N_92,N_25);
and U1066 (N_1066,N_505,N_457);
and U1067 (N_1067,N_6,N_611);
nor U1068 (N_1068,N_215,N_799);
and U1069 (N_1069,N_528,N_395);
and U1070 (N_1070,N_807,N_328);
or U1071 (N_1071,N_537,N_287);
nand U1072 (N_1072,N_561,N_659);
nor U1073 (N_1073,N_959,N_875);
and U1074 (N_1074,N_952,N_673);
nor U1075 (N_1075,N_800,N_316);
nand U1076 (N_1076,N_727,N_651);
nor U1077 (N_1077,N_298,N_418);
nand U1078 (N_1078,N_376,N_129);
nand U1079 (N_1079,N_802,N_748);
or U1080 (N_1080,N_760,N_284);
and U1081 (N_1081,N_677,N_962);
and U1082 (N_1082,N_307,N_332);
nand U1083 (N_1083,N_638,N_977);
or U1084 (N_1084,N_219,N_456);
and U1085 (N_1085,N_706,N_409);
and U1086 (N_1086,N_891,N_730);
nor U1087 (N_1087,N_646,N_989);
nor U1088 (N_1088,N_415,N_656);
or U1089 (N_1089,N_755,N_77);
or U1090 (N_1090,N_822,N_21);
nor U1091 (N_1091,N_979,N_434);
and U1092 (N_1092,N_905,N_696);
nor U1093 (N_1093,N_243,N_902);
nand U1094 (N_1094,N_728,N_67);
and U1095 (N_1095,N_652,N_927);
nor U1096 (N_1096,N_278,N_444);
and U1097 (N_1097,N_876,N_360);
or U1098 (N_1098,N_480,N_443);
nand U1099 (N_1099,N_202,N_681);
or U1100 (N_1100,N_381,N_591);
nor U1101 (N_1101,N_211,N_11);
or U1102 (N_1102,N_42,N_806);
or U1103 (N_1103,N_749,N_442);
nor U1104 (N_1104,N_761,N_470);
and U1105 (N_1105,N_58,N_746);
nor U1106 (N_1106,N_174,N_966);
nand U1107 (N_1107,N_897,N_941);
nand U1108 (N_1108,N_453,N_449);
or U1109 (N_1109,N_54,N_855);
nand U1110 (N_1110,N_546,N_489);
nor U1111 (N_1111,N_57,N_141);
or U1112 (N_1112,N_170,N_705);
or U1113 (N_1113,N_639,N_785);
or U1114 (N_1114,N_585,N_130);
nor U1115 (N_1115,N_257,N_793);
xor U1116 (N_1116,N_921,N_766);
or U1117 (N_1117,N_819,N_616);
and U1118 (N_1118,N_44,N_304);
or U1119 (N_1119,N_72,N_474);
or U1120 (N_1120,N_380,N_955);
and U1121 (N_1121,N_613,N_637);
nand U1122 (N_1122,N_144,N_685);
nand U1123 (N_1123,N_884,N_88);
or U1124 (N_1124,N_347,N_187);
or U1125 (N_1125,N_910,N_967);
nand U1126 (N_1126,N_394,N_544);
nand U1127 (N_1127,N_916,N_349);
or U1128 (N_1128,N_837,N_943);
nor U1129 (N_1129,N_752,N_826);
nand U1130 (N_1130,N_814,N_859);
and U1131 (N_1131,N_7,N_221);
nor U1132 (N_1132,N_156,N_632);
nor U1133 (N_1133,N_993,N_898);
nand U1134 (N_1134,N_530,N_960);
and U1135 (N_1135,N_410,N_580);
or U1136 (N_1136,N_687,N_241);
or U1137 (N_1137,N_85,N_868);
or U1138 (N_1138,N_145,N_886);
nand U1139 (N_1139,N_400,N_95);
or U1140 (N_1140,N_532,N_991);
and U1141 (N_1141,N_533,N_622);
nor U1142 (N_1142,N_121,N_280);
and U1143 (N_1143,N_606,N_348);
and U1144 (N_1144,N_683,N_820);
nor U1145 (N_1145,N_45,N_708);
nor U1146 (N_1146,N_213,N_512);
or U1147 (N_1147,N_231,N_176);
or U1148 (N_1148,N_322,N_279);
and U1149 (N_1149,N_5,N_3);
nand U1150 (N_1150,N_191,N_574);
nor U1151 (N_1151,N_40,N_199);
nor U1152 (N_1152,N_570,N_758);
and U1153 (N_1153,N_356,N_147);
nand U1154 (N_1154,N_244,N_481);
and U1155 (N_1155,N_306,N_850);
or U1156 (N_1156,N_282,N_900);
nand U1157 (N_1157,N_392,N_290);
nand U1158 (N_1158,N_37,N_76);
or U1159 (N_1159,N_620,N_119);
nand U1160 (N_1160,N_90,N_274);
nand U1161 (N_1161,N_735,N_817);
nand U1162 (N_1162,N_869,N_260);
nor U1163 (N_1163,N_317,N_522);
and U1164 (N_1164,N_458,N_168);
nor U1165 (N_1165,N_265,N_153);
nand U1166 (N_1166,N_894,N_940);
or U1167 (N_1167,N_224,N_116);
or U1168 (N_1168,N_430,N_240);
nor U1169 (N_1169,N_981,N_329);
and U1170 (N_1170,N_520,N_581);
or U1171 (N_1171,N_105,N_674);
and U1172 (N_1172,N_190,N_678);
nor U1173 (N_1173,N_253,N_593);
and U1174 (N_1174,N_261,N_325);
xor U1175 (N_1175,N_416,N_536);
and U1176 (N_1176,N_102,N_469);
nor U1177 (N_1177,N_556,N_23);
nand U1178 (N_1178,N_487,N_873);
nor U1179 (N_1179,N_247,N_914);
and U1180 (N_1180,N_524,N_689);
and U1181 (N_1181,N_465,N_948);
nor U1182 (N_1182,N_635,N_729);
nand U1183 (N_1183,N_657,N_340);
nand U1184 (N_1184,N_477,N_971);
or U1185 (N_1185,N_200,N_703);
nor U1186 (N_1186,N_441,N_839);
nand U1187 (N_1187,N_890,N_214);
nor U1188 (N_1188,N_964,N_535);
or U1189 (N_1189,N_973,N_374);
nand U1190 (N_1190,N_313,N_399);
and U1191 (N_1191,N_552,N_836);
and U1192 (N_1192,N_180,N_136);
nand U1193 (N_1193,N_929,N_391);
or U1194 (N_1194,N_663,N_589);
xnor U1195 (N_1195,N_628,N_848);
and U1196 (N_1196,N_994,N_676);
nor U1197 (N_1197,N_816,N_909);
nor U1198 (N_1198,N_695,N_852);
or U1199 (N_1199,N_545,N_52);
and U1200 (N_1200,N_650,N_438);
nand U1201 (N_1201,N_935,N_341);
nor U1202 (N_1202,N_359,N_292);
or U1203 (N_1203,N_361,N_779);
nor U1204 (N_1204,N_59,N_547);
and U1205 (N_1205,N_984,N_733);
nand U1206 (N_1206,N_510,N_185);
nand U1207 (N_1207,N_775,N_513);
nor U1208 (N_1208,N_28,N_149);
or U1209 (N_1209,N_812,N_216);
nand U1210 (N_1210,N_120,N_588);
nand U1211 (N_1211,N_326,N_866);
and U1212 (N_1212,N_173,N_60);
nor U1213 (N_1213,N_83,N_331);
nand U1214 (N_1214,N_534,N_872);
nor U1215 (N_1215,N_798,N_710);
or U1216 (N_1216,N_143,N_383);
nor U1217 (N_1217,N_100,N_669);
or U1218 (N_1218,N_122,N_186);
nand U1219 (N_1219,N_756,N_161);
nor U1220 (N_1220,N_849,N_932);
nand U1221 (N_1221,N_351,N_867);
nand U1222 (N_1222,N_63,N_901);
nor U1223 (N_1223,N_237,N_508);
and U1224 (N_1224,N_609,N_472);
nand U1225 (N_1225,N_188,N_767);
nand U1226 (N_1226,N_539,N_634);
and U1227 (N_1227,N_579,N_305);
nor U1228 (N_1228,N_835,N_499);
nand U1229 (N_1229,N_664,N_562);
or U1230 (N_1230,N_169,N_18);
and U1231 (N_1231,N_682,N_759);
nand U1232 (N_1232,N_700,N_365);
and U1233 (N_1233,N_908,N_658);
nor U1234 (N_1234,N_327,N_911);
and U1235 (N_1235,N_89,N_87);
nor U1236 (N_1236,N_20,N_98);
or U1237 (N_1237,N_953,N_297);
and U1238 (N_1238,N_670,N_109);
nand U1239 (N_1239,N_507,N_990);
nand U1240 (N_1240,N_406,N_791);
nand U1241 (N_1241,N_968,N_492);
nor U1242 (N_1242,N_488,N_963);
and U1243 (N_1243,N_289,N_398);
and U1244 (N_1244,N_350,N_584);
or U1245 (N_1245,N_572,N_14);
and U1246 (N_1246,N_466,N_601);
or U1247 (N_1247,N_704,N_242);
and U1248 (N_1248,N_414,N_600);
nand U1249 (N_1249,N_462,N_471);
nand U1250 (N_1250,N_51,N_47);
and U1251 (N_1251,N_969,N_525);
and U1252 (N_1252,N_636,N_716);
nand U1253 (N_1253,N_889,N_714);
nand U1254 (N_1254,N_654,N_346);
nand U1255 (N_1255,N_46,N_934);
nand U1256 (N_1256,N_645,N_235);
nand U1257 (N_1257,N_691,N_140);
nand U1258 (N_1258,N_596,N_15);
nor U1259 (N_1259,N_846,N_753);
xnor U1260 (N_1260,N_773,N_159);
or U1261 (N_1261,N_516,N_148);
nand U1262 (N_1262,N_277,N_938);
nand U1263 (N_1263,N_106,N_750);
nor U1264 (N_1264,N_203,N_1);
nor U1265 (N_1265,N_128,N_649);
nor U1266 (N_1266,N_734,N_97);
and U1267 (N_1267,N_267,N_2);
nand U1268 (N_1268,N_563,N_368);
nand U1269 (N_1269,N_854,N_421);
or U1270 (N_1270,N_565,N_223);
or U1271 (N_1271,N_93,N_878);
or U1272 (N_1272,N_363,N_906);
or U1273 (N_1273,N_286,N_554);
nand U1274 (N_1274,N_222,N_496);
nor U1275 (N_1275,N_160,N_566);
and U1276 (N_1276,N_323,N_895);
nand U1277 (N_1277,N_299,N_269);
nand U1278 (N_1278,N_372,N_437);
or U1279 (N_1279,N_619,N_560);
and U1280 (N_1280,N_127,N_576);
nor U1281 (N_1281,N_825,N_643);
or U1282 (N_1282,N_251,N_762);
xnor U1283 (N_1283,N_460,N_80);
and U1284 (N_1284,N_111,N_803);
nor U1285 (N_1285,N_805,N_234);
nand U1286 (N_1286,N_110,N_523);
xor U1287 (N_1287,N_204,N_847);
and U1288 (N_1288,N_980,N_519);
and U1289 (N_1289,N_856,N_833);
or U1290 (N_1290,N_427,N_899);
and U1291 (N_1291,N_428,N_64);
or U1292 (N_1292,N_412,N_396);
and U1293 (N_1293,N_958,N_841);
nand U1294 (N_1294,N_165,N_62);
nand U1295 (N_1295,N_74,N_49);
nor U1296 (N_1296,N_135,N_312);
and U1297 (N_1297,N_594,N_781);
nor U1298 (N_1298,N_151,N_384);
and U1299 (N_1299,N_404,N_192);
nor U1300 (N_1300,N_553,N_468);
nor U1301 (N_1301,N_425,N_961);
and U1302 (N_1302,N_925,N_81);
nor U1303 (N_1303,N_16,N_238);
nand U1304 (N_1304,N_975,N_486);
or U1305 (N_1305,N_358,N_86);
nand U1306 (N_1306,N_411,N_920);
nor U1307 (N_1307,N_629,N_701);
nor U1308 (N_1308,N_357,N_715);
and U1309 (N_1309,N_692,N_671);
and U1310 (N_1310,N_809,N_476);
and U1311 (N_1311,N_194,N_624);
nor U1312 (N_1312,N_690,N_254);
and U1313 (N_1313,N_995,N_717);
nand U1314 (N_1314,N_724,N_402);
and U1315 (N_1315,N_882,N_569);
nand U1316 (N_1316,N_285,N_114);
nor U1317 (N_1317,N_947,N_722);
or U1318 (N_1318,N_737,N_838);
and U1319 (N_1319,N_436,N_827);
nor U1320 (N_1320,N_229,N_336);
or U1321 (N_1321,N_24,N_686);
or U1322 (N_1322,N_367,N_408);
or U1323 (N_1323,N_273,N_684);
or U1324 (N_1324,N_65,N_840);
and U1325 (N_1325,N_455,N_739);
nand U1326 (N_1326,N_503,N_271);
and U1327 (N_1327,N_521,N_193);
and U1328 (N_1328,N_543,N_440);
or U1329 (N_1329,N_272,N_912);
and U1330 (N_1330,N_871,N_550);
or U1331 (N_1331,N_205,N_256);
or U1332 (N_1332,N_780,N_834);
or U1333 (N_1333,N_778,N_974);
or U1334 (N_1334,N_608,N_452);
and U1335 (N_1335,N_885,N_9);
and U1336 (N_1336,N_987,N_68);
nor U1337 (N_1337,N_506,N_551);
or U1338 (N_1338,N_870,N_397);
xor U1339 (N_1339,N_931,N_502);
or U1340 (N_1340,N_725,N_924);
and U1341 (N_1341,N_195,N_107);
or U1342 (N_1342,N_473,N_432);
nor U1343 (N_1343,N_318,N_484);
nand U1344 (N_1344,N_607,N_747);
nand U1345 (N_1345,N_245,N_104);
or U1346 (N_1346,N_810,N_933);
nor U1347 (N_1347,N_407,N_34);
and U1348 (N_1348,N_0,N_309);
and U1349 (N_1349,N_19,N_660);
nor U1350 (N_1350,N_568,N_655);
nor U1351 (N_1351,N_288,N_291);
nand U1352 (N_1352,N_592,N_447);
nand U1353 (N_1353,N_857,N_178);
nor U1354 (N_1354,N_998,N_258);
nor U1355 (N_1355,N_571,N_459);
nand U1356 (N_1356,N_988,N_61);
nor U1357 (N_1357,N_248,N_757);
and U1358 (N_1358,N_598,N_48);
nand U1359 (N_1359,N_218,N_263);
or U1360 (N_1360,N_232,N_661);
and U1361 (N_1361,N_698,N_723);
or U1362 (N_1362,N_352,N_694);
nand U1363 (N_1363,N_485,N_117);
and U1364 (N_1364,N_483,N_220);
nor U1365 (N_1365,N_514,N_919);
or U1366 (N_1366,N_720,N_500);
nor U1367 (N_1367,N_390,N_230);
or U1368 (N_1368,N_946,N_56);
nor U1369 (N_1369,N_362,N_731);
or U1370 (N_1370,N_930,N_618);
nand U1371 (N_1371,N_567,N_228);
and U1372 (N_1372,N_22,N_903);
and U1373 (N_1373,N_879,N_662);
nor U1374 (N_1374,N_937,N_642);
and U1375 (N_1375,N_84,N_422);
nand U1376 (N_1376,N_776,N_131);
or U1377 (N_1377,N_445,N_99);
nor U1378 (N_1378,N_978,N_982);
or U1379 (N_1379,N_549,N_478);
nand U1380 (N_1380,N_255,N_198);
or U1381 (N_1381,N_463,N_482);
nand U1382 (N_1382,N_252,N_501);
or U1383 (N_1383,N_385,N_184);
and U1384 (N_1384,N_4,N_754);
and U1385 (N_1385,N_167,N_163);
nor U1386 (N_1386,N_804,N_883);
and U1387 (N_1387,N_33,N_233);
nand U1388 (N_1388,N_264,N_393);
nor U1389 (N_1389,N_495,N_124);
or U1390 (N_1390,N_702,N_225);
and U1391 (N_1391,N_155,N_490);
and U1392 (N_1392,N_603,N_339);
and U1393 (N_1393,N_118,N_125);
and U1394 (N_1394,N_542,N_858);
and U1395 (N_1395,N_913,N_648);
or U1396 (N_1396,N_792,N_853);
and U1397 (N_1397,N_172,N_790);
or U1398 (N_1398,N_832,N_712);
nand U1399 (N_1399,N_275,N_688);
and U1400 (N_1400,N_582,N_877);
nand U1401 (N_1401,N_610,N_413);
and U1402 (N_1402,N_672,N_771);
nor U1403 (N_1403,N_864,N_17);
and U1404 (N_1404,N_796,N_531);
nor U1405 (N_1405,N_605,N_132);
or U1406 (N_1406,N_559,N_942);
and U1407 (N_1407,N_301,N_851);
and U1408 (N_1408,N_259,N_377);
and U1409 (N_1409,N_788,N_302);
nand U1410 (N_1410,N_770,N_454);
nor U1411 (N_1411,N_764,N_30);
and U1412 (N_1412,N_207,N_226);
nand U1413 (N_1413,N_177,N_78);
nor U1414 (N_1414,N_811,N_446);
or U1415 (N_1415,N_815,N_420);
nor U1416 (N_1416,N_831,N_986);
nand U1417 (N_1417,N_517,N_548);
nand U1418 (N_1418,N_308,N_53);
or U1419 (N_1419,N_158,N_887);
and U1420 (N_1420,N_196,N_138);
or U1421 (N_1421,N_491,N_26);
and U1422 (N_1422,N_137,N_142);
or U1423 (N_1423,N_8,N_604);
nand U1424 (N_1424,N_157,N_928);
nand U1425 (N_1425,N_379,N_27);
and U1426 (N_1426,N_845,N_794);
and U1427 (N_1427,N_709,N_36);
and U1428 (N_1428,N_526,N_633);
nand U1429 (N_1429,N_699,N_653);
nor U1430 (N_1430,N_333,N_926);
or U1431 (N_1431,N_249,N_765);
or U1432 (N_1432,N_208,N_541);
or U1433 (N_1433,N_511,N_641);
nor U1434 (N_1434,N_939,N_719);
nor U1435 (N_1435,N_268,N_315);
nand U1436 (N_1436,N_915,N_164);
and U1437 (N_1437,N_162,N_768);
nand U1438 (N_1438,N_538,N_401);
nand U1439 (N_1439,N_801,N_965);
nor U1440 (N_1440,N_429,N_564);
nand U1441 (N_1441,N_370,N_999);
and U1442 (N_1442,N_772,N_69);
nor U1443 (N_1443,N_666,N_630);
or U1444 (N_1444,N_721,N_595);
nand U1445 (N_1445,N_386,N_276);
and U1446 (N_1446,N_917,N_992);
and U1447 (N_1447,N_342,N_73);
and U1448 (N_1448,N_985,N_13);
and U1449 (N_1449,N_769,N_972);
and U1450 (N_1450,N_189,N_627);
and U1451 (N_1451,N_527,N_91);
nand U1452 (N_1452,N_679,N_843);
and U1453 (N_1453,N_923,N_573);
nand U1454 (N_1454,N_956,N_439);
or U1455 (N_1455,N_738,N_353);
and U1456 (N_1456,N_784,N_555);
or U1457 (N_1457,N_461,N_343);
and U1458 (N_1458,N_874,N_936);
nand U1459 (N_1459,N_996,N_602);
and U1460 (N_1460,N_35,N_997);
nor U1461 (N_1461,N_154,N_126);
nor U1462 (N_1462,N_945,N_976);
nand U1463 (N_1463,N_206,N_590);
or U1464 (N_1464,N_345,N_364);
and U1465 (N_1465,N_744,N_494);
or U1466 (N_1466,N_417,N_865);
and U1467 (N_1467,N_893,N_133);
or U1468 (N_1468,N_518,N_10);
nor U1469 (N_1469,N_904,N_371);
nor U1470 (N_1470,N_283,N_344);
nand U1471 (N_1471,N_558,N_578);
nor U1472 (N_1472,N_667,N_236);
nand U1473 (N_1473,N_707,N_640);
nor U1474 (N_1474,N_175,N_31);
or U1475 (N_1475,N_115,N_217);
nor U1476 (N_1476,N_266,N_983);
nor U1477 (N_1477,N_475,N_892);
nand U1478 (N_1478,N_842,N_668);
or U1479 (N_1479,N_270,N_950);
and U1480 (N_1480,N_665,N_808);
or U1481 (N_1481,N_713,N_32);
nand U1482 (N_1482,N_631,N_303);
nor U1483 (N_1483,N_529,N_644);
nor U1484 (N_1484,N_599,N_250);
and U1485 (N_1485,N_786,N_12);
nand U1486 (N_1486,N_387,N_227);
nand U1487 (N_1487,N_742,N_300);
nand U1488 (N_1488,N_954,N_828);
nor U1489 (N_1489,N_103,N_355);
nand U1490 (N_1490,N_597,N_101);
and U1491 (N_1491,N_711,N_311);
or U1492 (N_1492,N_918,N_647);
and U1493 (N_1493,N_451,N_467);
or U1494 (N_1494,N_575,N_583);
and U1495 (N_1495,N_295,N_881);
nor U1496 (N_1496,N_763,N_777);
nand U1497 (N_1497,N_789,N_736);
or U1498 (N_1498,N_96,N_321);
or U1499 (N_1499,N_66,N_209);
and U1500 (N_1500,N_404,N_55);
and U1501 (N_1501,N_259,N_805);
and U1502 (N_1502,N_497,N_145);
or U1503 (N_1503,N_816,N_574);
or U1504 (N_1504,N_492,N_168);
nand U1505 (N_1505,N_352,N_662);
nand U1506 (N_1506,N_781,N_23);
and U1507 (N_1507,N_55,N_680);
nor U1508 (N_1508,N_599,N_910);
nand U1509 (N_1509,N_29,N_367);
nor U1510 (N_1510,N_993,N_259);
nor U1511 (N_1511,N_550,N_783);
nand U1512 (N_1512,N_522,N_235);
nand U1513 (N_1513,N_757,N_409);
or U1514 (N_1514,N_236,N_210);
and U1515 (N_1515,N_754,N_242);
nor U1516 (N_1516,N_111,N_248);
xor U1517 (N_1517,N_638,N_518);
nor U1518 (N_1518,N_470,N_540);
or U1519 (N_1519,N_852,N_466);
or U1520 (N_1520,N_281,N_520);
nor U1521 (N_1521,N_534,N_125);
or U1522 (N_1522,N_151,N_792);
nor U1523 (N_1523,N_649,N_10);
and U1524 (N_1524,N_208,N_215);
nor U1525 (N_1525,N_135,N_735);
nand U1526 (N_1526,N_130,N_289);
or U1527 (N_1527,N_222,N_71);
or U1528 (N_1528,N_45,N_179);
and U1529 (N_1529,N_3,N_198);
nand U1530 (N_1530,N_631,N_756);
nand U1531 (N_1531,N_693,N_651);
or U1532 (N_1532,N_798,N_287);
nor U1533 (N_1533,N_581,N_130);
or U1534 (N_1534,N_281,N_937);
or U1535 (N_1535,N_818,N_595);
nand U1536 (N_1536,N_805,N_970);
nand U1537 (N_1537,N_360,N_336);
nor U1538 (N_1538,N_927,N_412);
or U1539 (N_1539,N_345,N_909);
or U1540 (N_1540,N_75,N_867);
nand U1541 (N_1541,N_647,N_699);
and U1542 (N_1542,N_961,N_680);
or U1543 (N_1543,N_452,N_284);
or U1544 (N_1544,N_948,N_414);
or U1545 (N_1545,N_342,N_810);
nand U1546 (N_1546,N_34,N_377);
nand U1547 (N_1547,N_745,N_918);
nand U1548 (N_1548,N_195,N_95);
nand U1549 (N_1549,N_289,N_596);
nor U1550 (N_1550,N_735,N_876);
nor U1551 (N_1551,N_542,N_490);
nand U1552 (N_1552,N_464,N_320);
or U1553 (N_1553,N_511,N_168);
and U1554 (N_1554,N_296,N_957);
nor U1555 (N_1555,N_583,N_360);
nand U1556 (N_1556,N_374,N_558);
nand U1557 (N_1557,N_653,N_949);
nor U1558 (N_1558,N_847,N_384);
nor U1559 (N_1559,N_207,N_16);
nand U1560 (N_1560,N_158,N_844);
and U1561 (N_1561,N_761,N_206);
and U1562 (N_1562,N_560,N_411);
nand U1563 (N_1563,N_615,N_413);
and U1564 (N_1564,N_282,N_526);
or U1565 (N_1565,N_9,N_698);
nor U1566 (N_1566,N_27,N_81);
nor U1567 (N_1567,N_197,N_768);
nand U1568 (N_1568,N_736,N_491);
nor U1569 (N_1569,N_509,N_919);
nor U1570 (N_1570,N_131,N_312);
and U1571 (N_1571,N_25,N_727);
and U1572 (N_1572,N_611,N_974);
nand U1573 (N_1573,N_998,N_806);
or U1574 (N_1574,N_52,N_38);
and U1575 (N_1575,N_787,N_391);
and U1576 (N_1576,N_894,N_151);
nand U1577 (N_1577,N_35,N_884);
nor U1578 (N_1578,N_918,N_869);
nand U1579 (N_1579,N_759,N_974);
nor U1580 (N_1580,N_237,N_396);
or U1581 (N_1581,N_471,N_199);
nor U1582 (N_1582,N_813,N_188);
and U1583 (N_1583,N_459,N_757);
or U1584 (N_1584,N_152,N_935);
or U1585 (N_1585,N_673,N_75);
or U1586 (N_1586,N_403,N_673);
nor U1587 (N_1587,N_672,N_686);
or U1588 (N_1588,N_596,N_819);
nand U1589 (N_1589,N_996,N_20);
and U1590 (N_1590,N_364,N_128);
or U1591 (N_1591,N_348,N_409);
or U1592 (N_1592,N_559,N_524);
nand U1593 (N_1593,N_463,N_457);
nand U1594 (N_1594,N_145,N_978);
nand U1595 (N_1595,N_960,N_188);
or U1596 (N_1596,N_867,N_23);
nand U1597 (N_1597,N_10,N_455);
nand U1598 (N_1598,N_857,N_158);
or U1599 (N_1599,N_979,N_806);
nand U1600 (N_1600,N_61,N_233);
nand U1601 (N_1601,N_549,N_799);
or U1602 (N_1602,N_581,N_984);
and U1603 (N_1603,N_84,N_668);
nor U1604 (N_1604,N_92,N_891);
nand U1605 (N_1605,N_428,N_866);
nand U1606 (N_1606,N_916,N_837);
nand U1607 (N_1607,N_422,N_366);
nor U1608 (N_1608,N_471,N_699);
nor U1609 (N_1609,N_825,N_884);
and U1610 (N_1610,N_586,N_526);
nand U1611 (N_1611,N_520,N_230);
nor U1612 (N_1612,N_667,N_42);
and U1613 (N_1613,N_369,N_177);
or U1614 (N_1614,N_253,N_140);
and U1615 (N_1615,N_443,N_295);
nand U1616 (N_1616,N_366,N_145);
xnor U1617 (N_1617,N_817,N_371);
and U1618 (N_1618,N_244,N_731);
nor U1619 (N_1619,N_962,N_117);
xnor U1620 (N_1620,N_318,N_481);
and U1621 (N_1621,N_168,N_271);
nor U1622 (N_1622,N_284,N_417);
and U1623 (N_1623,N_396,N_91);
nand U1624 (N_1624,N_207,N_416);
nor U1625 (N_1625,N_860,N_755);
nand U1626 (N_1626,N_81,N_511);
nor U1627 (N_1627,N_277,N_609);
or U1628 (N_1628,N_610,N_906);
and U1629 (N_1629,N_325,N_354);
nor U1630 (N_1630,N_395,N_956);
or U1631 (N_1631,N_902,N_24);
and U1632 (N_1632,N_395,N_998);
and U1633 (N_1633,N_634,N_254);
nand U1634 (N_1634,N_219,N_316);
nor U1635 (N_1635,N_29,N_953);
and U1636 (N_1636,N_379,N_885);
nand U1637 (N_1637,N_721,N_860);
or U1638 (N_1638,N_832,N_762);
nand U1639 (N_1639,N_797,N_173);
nor U1640 (N_1640,N_280,N_935);
xnor U1641 (N_1641,N_390,N_689);
nand U1642 (N_1642,N_290,N_856);
and U1643 (N_1643,N_602,N_705);
and U1644 (N_1644,N_920,N_982);
and U1645 (N_1645,N_995,N_616);
nor U1646 (N_1646,N_272,N_743);
nand U1647 (N_1647,N_83,N_71);
xor U1648 (N_1648,N_870,N_269);
nor U1649 (N_1649,N_179,N_471);
nand U1650 (N_1650,N_90,N_945);
and U1651 (N_1651,N_24,N_135);
and U1652 (N_1652,N_619,N_510);
nand U1653 (N_1653,N_399,N_784);
nor U1654 (N_1654,N_447,N_267);
nor U1655 (N_1655,N_269,N_779);
nor U1656 (N_1656,N_644,N_750);
nand U1657 (N_1657,N_375,N_771);
and U1658 (N_1658,N_38,N_549);
nor U1659 (N_1659,N_97,N_646);
or U1660 (N_1660,N_572,N_886);
nor U1661 (N_1661,N_710,N_516);
and U1662 (N_1662,N_865,N_851);
nor U1663 (N_1663,N_99,N_384);
nor U1664 (N_1664,N_433,N_585);
nor U1665 (N_1665,N_372,N_688);
or U1666 (N_1666,N_42,N_113);
nand U1667 (N_1667,N_676,N_356);
nor U1668 (N_1668,N_203,N_168);
nor U1669 (N_1669,N_663,N_548);
nor U1670 (N_1670,N_146,N_609);
or U1671 (N_1671,N_383,N_459);
nor U1672 (N_1672,N_732,N_385);
nand U1673 (N_1673,N_994,N_140);
and U1674 (N_1674,N_441,N_604);
or U1675 (N_1675,N_48,N_436);
and U1676 (N_1676,N_158,N_132);
nor U1677 (N_1677,N_326,N_786);
nand U1678 (N_1678,N_653,N_980);
nand U1679 (N_1679,N_321,N_230);
nor U1680 (N_1680,N_625,N_149);
and U1681 (N_1681,N_945,N_473);
or U1682 (N_1682,N_654,N_220);
and U1683 (N_1683,N_790,N_672);
and U1684 (N_1684,N_341,N_548);
and U1685 (N_1685,N_749,N_50);
nand U1686 (N_1686,N_208,N_406);
nor U1687 (N_1687,N_96,N_232);
nand U1688 (N_1688,N_891,N_716);
nand U1689 (N_1689,N_555,N_565);
nor U1690 (N_1690,N_127,N_67);
or U1691 (N_1691,N_125,N_766);
and U1692 (N_1692,N_563,N_46);
or U1693 (N_1693,N_414,N_221);
nor U1694 (N_1694,N_845,N_523);
nor U1695 (N_1695,N_409,N_890);
or U1696 (N_1696,N_958,N_272);
nand U1697 (N_1697,N_877,N_298);
or U1698 (N_1698,N_731,N_432);
or U1699 (N_1699,N_865,N_24);
nor U1700 (N_1700,N_991,N_968);
and U1701 (N_1701,N_370,N_337);
nand U1702 (N_1702,N_251,N_467);
and U1703 (N_1703,N_861,N_469);
and U1704 (N_1704,N_241,N_487);
or U1705 (N_1705,N_337,N_360);
nor U1706 (N_1706,N_679,N_371);
nand U1707 (N_1707,N_548,N_842);
and U1708 (N_1708,N_586,N_313);
nand U1709 (N_1709,N_619,N_424);
and U1710 (N_1710,N_68,N_298);
nand U1711 (N_1711,N_937,N_259);
or U1712 (N_1712,N_692,N_414);
or U1713 (N_1713,N_544,N_427);
nor U1714 (N_1714,N_347,N_941);
nand U1715 (N_1715,N_651,N_659);
nor U1716 (N_1716,N_759,N_288);
and U1717 (N_1717,N_263,N_327);
nand U1718 (N_1718,N_638,N_827);
or U1719 (N_1719,N_712,N_726);
or U1720 (N_1720,N_382,N_62);
or U1721 (N_1721,N_457,N_846);
or U1722 (N_1722,N_158,N_708);
nor U1723 (N_1723,N_585,N_818);
or U1724 (N_1724,N_184,N_427);
nand U1725 (N_1725,N_542,N_191);
nor U1726 (N_1726,N_59,N_922);
or U1727 (N_1727,N_850,N_646);
nand U1728 (N_1728,N_52,N_362);
and U1729 (N_1729,N_71,N_210);
xnor U1730 (N_1730,N_655,N_598);
and U1731 (N_1731,N_769,N_475);
or U1732 (N_1732,N_36,N_152);
nor U1733 (N_1733,N_51,N_995);
or U1734 (N_1734,N_907,N_162);
nand U1735 (N_1735,N_883,N_179);
nor U1736 (N_1736,N_741,N_213);
and U1737 (N_1737,N_849,N_12);
nand U1738 (N_1738,N_288,N_276);
or U1739 (N_1739,N_36,N_113);
or U1740 (N_1740,N_366,N_539);
nand U1741 (N_1741,N_453,N_891);
nor U1742 (N_1742,N_122,N_150);
nand U1743 (N_1743,N_529,N_43);
nor U1744 (N_1744,N_165,N_664);
nand U1745 (N_1745,N_776,N_530);
nand U1746 (N_1746,N_2,N_51);
and U1747 (N_1747,N_16,N_657);
nor U1748 (N_1748,N_866,N_148);
nor U1749 (N_1749,N_772,N_898);
nand U1750 (N_1750,N_404,N_308);
or U1751 (N_1751,N_694,N_474);
nor U1752 (N_1752,N_720,N_386);
or U1753 (N_1753,N_0,N_55);
nand U1754 (N_1754,N_927,N_74);
and U1755 (N_1755,N_690,N_544);
nor U1756 (N_1756,N_518,N_687);
nor U1757 (N_1757,N_897,N_29);
and U1758 (N_1758,N_207,N_560);
or U1759 (N_1759,N_943,N_879);
and U1760 (N_1760,N_834,N_53);
and U1761 (N_1761,N_872,N_12);
nand U1762 (N_1762,N_27,N_767);
nand U1763 (N_1763,N_758,N_81);
nand U1764 (N_1764,N_513,N_630);
and U1765 (N_1765,N_472,N_736);
nand U1766 (N_1766,N_328,N_300);
and U1767 (N_1767,N_13,N_556);
nand U1768 (N_1768,N_791,N_545);
or U1769 (N_1769,N_462,N_295);
or U1770 (N_1770,N_326,N_682);
and U1771 (N_1771,N_521,N_683);
nor U1772 (N_1772,N_70,N_213);
and U1773 (N_1773,N_132,N_624);
and U1774 (N_1774,N_170,N_120);
nand U1775 (N_1775,N_837,N_138);
nand U1776 (N_1776,N_730,N_296);
and U1777 (N_1777,N_946,N_557);
xor U1778 (N_1778,N_986,N_339);
or U1779 (N_1779,N_762,N_300);
nand U1780 (N_1780,N_21,N_113);
nand U1781 (N_1781,N_404,N_509);
and U1782 (N_1782,N_705,N_780);
xnor U1783 (N_1783,N_104,N_729);
nand U1784 (N_1784,N_576,N_842);
xor U1785 (N_1785,N_775,N_562);
nand U1786 (N_1786,N_142,N_339);
nor U1787 (N_1787,N_9,N_36);
and U1788 (N_1788,N_806,N_204);
and U1789 (N_1789,N_454,N_886);
nand U1790 (N_1790,N_130,N_91);
and U1791 (N_1791,N_140,N_268);
nor U1792 (N_1792,N_458,N_839);
nand U1793 (N_1793,N_615,N_969);
and U1794 (N_1794,N_18,N_724);
and U1795 (N_1795,N_589,N_274);
and U1796 (N_1796,N_531,N_342);
and U1797 (N_1797,N_913,N_218);
and U1798 (N_1798,N_353,N_680);
nand U1799 (N_1799,N_532,N_298);
or U1800 (N_1800,N_19,N_20);
and U1801 (N_1801,N_118,N_923);
nor U1802 (N_1802,N_304,N_288);
nand U1803 (N_1803,N_204,N_285);
or U1804 (N_1804,N_260,N_351);
nand U1805 (N_1805,N_105,N_318);
nand U1806 (N_1806,N_133,N_648);
nor U1807 (N_1807,N_717,N_888);
or U1808 (N_1808,N_843,N_406);
nand U1809 (N_1809,N_910,N_566);
and U1810 (N_1810,N_383,N_176);
nand U1811 (N_1811,N_648,N_549);
nor U1812 (N_1812,N_829,N_155);
and U1813 (N_1813,N_253,N_866);
nor U1814 (N_1814,N_430,N_933);
nand U1815 (N_1815,N_855,N_167);
or U1816 (N_1816,N_526,N_765);
nand U1817 (N_1817,N_739,N_547);
or U1818 (N_1818,N_194,N_440);
and U1819 (N_1819,N_183,N_323);
nor U1820 (N_1820,N_876,N_470);
nand U1821 (N_1821,N_483,N_190);
nor U1822 (N_1822,N_739,N_242);
and U1823 (N_1823,N_247,N_649);
or U1824 (N_1824,N_686,N_94);
and U1825 (N_1825,N_219,N_669);
nand U1826 (N_1826,N_472,N_674);
nor U1827 (N_1827,N_186,N_577);
nor U1828 (N_1828,N_663,N_83);
and U1829 (N_1829,N_257,N_169);
nor U1830 (N_1830,N_975,N_732);
or U1831 (N_1831,N_901,N_332);
or U1832 (N_1832,N_205,N_924);
and U1833 (N_1833,N_718,N_960);
and U1834 (N_1834,N_506,N_441);
or U1835 (N_1835,N_341,N_995);
and U1836 (N_1836,N_350,N_945);
nor U1837 (N_1837,N_150,N_641);
xor U1838 (N_1838,N_473,N_612);
nor U1839 (N_1839,N_988,N_985);
nand U1840 (N_1840,N_812,N_41);
nor U1841 (N_1841,N_42,N_402);
nor U1842 (N_1842,N_10,N_924);
and U1843 (N_1843,N_70,N_174);
and U1844 (N_1844,N_769,N_893);
nand U1845 (N_1845,N_49,N_581);
nand U1846 (N_1846,N_188,N_247);
nor U1847 (N_1847,N_545,N_891);
nor U1848 (N_1848,N_431,N_255);
nor U1849 (N_1849,N_85,N_447);
and U1850 (N_1850,N_6,N_549);
nand U1851 (N_1851,N_80,N_269);
or U1852 (N_1852,N_780,N_379);
or U1853 (N_1853,N_877,N_823);
or U1854 (N_1854,N_777,N_764);
xnor U1855 (N_1855,N_447,N_301);
nor U1856 (N_1856,N_912,N_909);
nand U1857 (N_1857,N_350,N_136);
or U1858 (N_1858,N_131,N_181);
nor U1859 (N_1859,N_356,N_607);
nand U1860 (N_1860,N_845,N_244);
or U1861 (N_1861,N_482,N_202);
or U1862 (N_1862,N_786,N_139);
or U1863 (N_1863,N_650,N_918);
nand U1864 (N_1864,N_806,N_418);
nor U1865 (N_1865,N_200,N_448);
nand U1866 (N_1866,N_159,N_385);
and U1867 (N_1867,N_669,N_195);
nor U1868 (N_1868,N_878,N_853);
and U1869 (N_1869,N_181,N_41);
nand U1870 (N_1870,N_746,N_321);
or U1871 (N_1871,N_571,N_19);
or U1872 (N_1872,N_518,N_996);
nor U1873 (N_1873,N_802,N_909);
and U1874 (N_1874,N_934,N_363);
or U1875 (N_1875,N_443,N_555);
and U1876 (N_1876,N_607,N_149);
and U1877 (N_1877,N_704,N_208);
and U1878 (N_1878,N_646,N_903);
nand U1879 (N_1879,N_339,N_87);
nor U1880 (N_1880,N_631,N_9);
xor U1881 (N_1881,N_581,N_735);
nor U1882 (N_1882,N_343,N_599);
nand U1883 (N_1883,N_114,N_295);
nor U1884 (N_1884,N_991,N_161);
or U1885 (N_1885,N_815,N_37);
or U1886 (N_1886,N_755,N_361);
and U1887 (N_1887,N_346,N_889);
or U1888 (N_1888,N_344,N_230);
nor U1889 (N_1889,N_563,N_875);
nor U1890 (N_1890,N_875,N_76);
and U1891 (N_1891,N_517,N_306);
or U1892 (N_1892,N_589,N_620);
or U1893 (N_1893,N_72,N_167);
nor U1894 (N_1894,N_205,N_461);
and U1895 (N_1895,N_23,N_465);
or U1896 (N_1896,N_212,N_914);
nand U1897 (N_1897,N_515,N_749);
nand U1898 (N_1898,N_238,N_496);
nand U1899 (N_1899,N_984,N_213);
or U1900 (N_1900,N_533,N_844);
nor U1901 (N_1901,N_934,N_525);
nor U1902 (N_1902,N_176,N_940);
and U1903 (N_1903,N_909,N_44);
or U1904 (N_1904,N_625,N_388);
nand U1905 (N_1905,N_582,N_408);
or U1906 (N_1906,N_260,N_838);
nor U1907 (N_1907,N_968,N_162);
nand U1908 (N_1908,N_226,N_300);
and U1909 (N_1909,N_643,N_47);
nand U1910 (N_1910,N_468,N_222);
nor U1911 (N_1911,N_408,N_890);
or U1912 (N_1912,N_501,N_992);
or U1913 (N_1913,N_871,N_924);
nand U1914 (N_1914,N_859,N_615);
nor U1915 (N_1915,N_270,N_37);
nand U1916 (N_1916,N_435,N_975);
and U1917 (N_1917,N_287,N_395);
or U1918 (N_1918,N_971,N_703);
or U1919 (N_1919,N_699,N_50);
and U1920 (N_1920,N_635,N_129);
nor U1921 (N_1921,N_529,N_846);
or U1922 (N_1922,N_979,N_25);
or U1923 (N_1923,N_575,N_492);
and U1924 (N_1924,N_18,N_749);
nor U1925 (N_1925,N_72,N_789);
and U1926 (N_1926,N_275,N_550);
or U1927 (N_1927,N_23,N_779);
nor U1928 (N_1928,N_533,N_397);
and U1929 (N_1929,N_859,N_596);
or U1930 (N_1930,N_762,N_726);
nand U1931 (N_1931,N_573,N_830);
or U1932 (N_1932,N_253,N_586);
nand U1933 (N_1933,N_180,N_738);
and U1934 (N_1934,N_321,N_583);
nand U1935 (N_1935,N_974,N_534);
nand U1936 (N_1936,N_644,N_386);
and U1937 (N_1937,N_950,N_475);
nand U1938 (N_1938,N_581,N_757);
and U1939 (N_1939,N_340,N_29);
nor U1940 (N_1940,N_697,N_488);
nor U1941 (N_1941,N_551,N_186);
nor U1942 (N_1942,N_116,N_311);
or U1943 (N_1943,N_120,N_559);
nand U1944 (N_1944,N_663,N_81);
nor U1945 (N_1945,N_655,N_794);
nand U1946 (N_1946,N_567,N_857);
nor U1947 (N_1947,N_367,N_277);
nor U1948 (N_1948,N_254,N_499);
nand U1949 (N_1949,N_752,N_54);
or U1950 (N_1950,N_866,N_811);
and U1951 (N_1951,N_131,N_91);
nand U1952 (N_1952,N_660,N_975);
nor U1953 (N_1953,N_560,N_70);
nor U1954 (N_1954,N_540,N_939);
nor U1955 (N_1955,N_222,N_630);
and U1956 (N_1956,N_738,N_668);
or U1957 (N_1957,N_858,N_797);
or U1958 (N_1958,N_145,N_15);
or U1959 (N_1959,N_282,N_348);
nor U1960 (N_1960,N_660,N_456);
nand U1961 (N_1961,N_9,N_959);
nand U1962 (N_1962,N_141,N_132);
and U1963 (N_1963,N_871,N_617);
and U1964 (N_1964,N_760,N_684);
nor U1965 (N_1965,N_795,N_457);
nand U1966 (N_1966,N_984,N_775);
nor U1967 (N_1967,N_211,N_335);
nor U1968 (N_1968,N_32,N_957);
nor U1969 (N_1969,N_961,N_457);
or U1970 (N_1970,N_901,N_157);
and U1971 (N_1971,N_239,N_105);
nor U1972 (N_1972,N_268,N_826);
nor U1973 (N_1973,N_562,N_710);
and U1974 (N_1974,N_897,N_365);
and U1975 (N_1975,N_874,N_847);
and U1976 (N_1976,N_390,N_560);
and U1977 (N_1977,N_961,N_326);
or U1978 (N_1978,N_501,N_668);
nand U1979 (N_1979,N_377,N_456);
nor U1980 (N_1980,N_340,N_225);
nor U1981 (N_1981,N_732,N_368);
nand U1982 (N_1982,N_374,N_353);
and U1983 (N_1983,N_887,N_684);
nand U1984 (N_1984,N_389,N_661);
or U1985 (N_1985,N_318,N_4);
and U1986 (N_1986,N_880,N_313);
or U1987 (N_1987,N_49,N_522);
nor U1988 (N_1988,N_596,N_849);
and U1989 (N_1989,N_891,N_13);
nor U1990 (N_1990,N_384,N_140);
nand U1991 (N_1991,N_418,N_109);
nand U1992 (N_1992,N_881,N_208);
or U1993 (N_1993,N_522,N_342);
nand U1994 (N_1994,N_718,N_161);
and U1995 (N_1995,N_234,N_946);
and U1996 (N_1996,N_647,N_531);
nor U1997 (N_1997,N_142,N_184);
nor U1998 (N_1998,N_753,N_67);
or U1999 (N_1999,N_672,N_249);
and U2000 (N_2000,N_1111,N_1003);
nor U2001 (N_2001,N_1127,N_1477);
and U2002 (N_2002,N_1972,N_1348);
and U2003 (N_2003,N_1522,N_1746);
and U2004 (N_2004,N_1354,N_1406);
nand U2005 (N_2005,N_1027,N_1496);
nand U2006 (N_2006,N_1474,N_1543);
and U2007 (N_2007,N_1575,N_1766);
nor U2008 (N_2008,N_1687,N_1779);
nor U2009 (N_2009,N_1770,N_1559);
or U2010 (N_2010,N_1061,N_1536);
or U2011 (N_2011,N_1789,N_1236);
or U2012 (N_2012,N_1119,N_1084);
and U2013 (N_2013,N_1197,N_1023);
nor U2014 (N_2014,N_1892,N_1918);
or U2015 (N_2015,N_1498,N_1100);
and U2016 (N_2016,N_1605,N_1514);
or U2017 (N_2017,N_1372,N_1211);
and U2018 (N_2018,N_1167,N_1499);
nor U2019 (N_2019,N_1884,N_1855);
or U2020 (N_2020,N_1070,N_1396);
or U2021 (N_2021,N_1753,N_1161);
nand U2022 (N_2022,N_1307,N_1908);
and U2023 (N_2023,N_1278,N_1482);
and U2024 (N_2024,N_1337,N_1114);
or U2025 (N_2025,N_1057,N_1568);
nand U2026 (N_2026,N_1875,N_1738);
nand U2027 (N_2027,N_1077,N_1137);
nor U2028 (N_2028,N_1535,N_1518);
or U2029 (N_2029,N_1022,N_1800);
nand U2030 (N_2030,N_1887,N_1312);
or U2031 (N_2031,N_1610,N_1511);
xor U2032 (N_2032,N_1683,N_1204);
xnor U2033 (N_2033,N_1504,N_1828);
and U2034 (N_2034,N_1836,N_1181);
xnor U2035 (N_2035,N_1270,N_1253);
nor U2036 (N_2036,N_1302,N_1798);
nand U2037 (N_2037,N_1890,N_1520);
or U2038 (N_2038,N_1633,N_1059);
or U2039 (N_2039,N_1885,N_1924);
nor U2040 (N_2040,N_1370,N_1635);
xnor U2041 (N_2041,N_1627,N_1615);
and U2042 (N_2042,N_1229,N_1716);
or U2043 (N_2043,N_1184,N_1437);
nand U2044 (N_2044,N_1851,N_1072);
and U2045 (N_2045,N_1400,N_1411);
nor U2046 (N_2046,N_1018,N_1228);
nor U2047 (N_2047,N_1539,N_1684);
nand U2048 (N_2048,N_1203,N_1345);
or U2049 (N_2049,N_1927,N_1313);
nor U2050 (N_2050,N_1825,N_1826);
or U2051 (N_2051,N_1930,N_1093);
nor U2052 (N_2052,N_1943,N_1816);
nand U2053 (N_2053,N_1830,N_1021);
and U2054 (N_2054,N_1419,N_1958);
and U2055 (N_2055,N_1448,N_1799);
and U2056 (N_2056,N_1421,N_1802);
or U2057 (N_2057,N_1858,N_1447);
or U2058 (N_2058,N_1174,N_1439);
and U2059 (N_2059,N_1443,N_1068);
and U2060 (N_2060,N_1284,N_1979);
nor U2061 (N_2061,N_1842,N_1945);
nor U2062 (N_2062,N_1444,N_1168);
nor U2063 (N_2063,N_1326,N_1860);
nor U2064 (N_2064,N_1827,N_1234);
or U2065 (N_2065,N_1462,N_1237);
nor U2066 (N_2066,N_1516,N_1880);
nor U2067 (N_2067,N_1777,N_1637);
nor U2068 (N_2068,N_1628,N_1612);
and U2069 (N_2069,N_1654,N_1846);
nor U2070 (N_2070,N_1220,N_1316);
nor U2071 (N_2071,N_1048,N_1865);
nand U2072 (N_2072,N_1926,N_1973);
nand U2073 (N_2073,N_1910,N_1105);
and U2074 (N_2074,N_1831,N_1937);
nand U2075 (N_2075,N_1676,N_1224);
nor U2076 (N_2076,N_1721,N_1032);
nor U2077 (N_2077,N_1269,N_1931);
nor U2078 (N_2078,N_1863,N_1704);
nand U2079 (N_2079,N_1121,N_1506);
and U2080 (N_2080,N_1634,N_1352);
or U2081 (N_2081,N_1581,N_1573);
or U2082 (N_2082,N_1192,N_1639);
and U2083 (N_2083,N_1445,N_1467);
or U2084 (N_2084,N_1727,N_1432);
and U2085 (N_2085,N_1953,N_1709);
and U2086 (N_2086,N_1784,N_1452);
and U2087 (N_2087,N_1383,N_1690);
and U2088 (N_2088,N_1940,N_1173);
nor U2089 (N_2089,N_1135,N_1378);
nand U2090 (N_2090,N_1668,N_1285);
nor U2091 (N_2091,N_1614,N_1702);
nand U2092 (N_2092,N_1899,N_1917);
nor U2093 (N_2093,N_1963,N_1685);
nor U2094 (N_2094,N_1975,N_1981);
and U2095 (N_2095,N_1146,N_1646);
or U2096 (N_2096,N_1889,N_1929);
nor U2097 (N_2097,N_1056,N_1182);
nor U2098 (N_2098,N_1758,N_1076);
nor U2099 (N_2099,N_1814,N_1970);
nor U2100 (N_2100,N_1571,N_1366);
nor U2101 (N_2101,N_1371,N_1155);
and U2102 (N_2102,N_1956,N_1706);
nand U2103 (N_2103,N_1948,N_1576);
nand U2104 (N_2104,N_1742,N_1916);
nand U2105 (N_2105,N_1081,N_1896);
and U2106 (N_2106,N_1636,N_1153);
nand U2107 (N_2107,N_1856,N_1459);
and U2108 (N_2108,N_1780,N_1233);
nand U2109 (N_2109,N_1425,N_1381);
nand U2110 (N_2110,N_1235,N_1095);
or U2111 (N_2111,N_1598,N_1824);
nor U2112 (N_2112,N_1544,N_1115);
or U2113 (N_2113,N_1607,N_1431);
nor U2114 (N_2114,N_1098,N_1672);
nor U2115 (N_2115,N_1271,N_1942);
nand U2116 (N_2116,N_1148,N_1810);
and U2117 (N_2117,N_1418,N_1531);
or U2118 (N_2118,N_1509,N_1004);
nand U2119 (N_2119,N_1440,N_1208);
or U2120 (N_2120,N_1349,N_1643);
and U2121 (N_2121,N_1151,N_1407);
and U2122 (N_2122,N_1232,N_1388);
and U2123 (N_2123,N_1176,N_1853);
and U2124 (N_2124,N_1397,N_1546);
nor U2125 (N_2125,N_1398,N_1703);
nor U2126 (N_2126,N_1997,N_1261);
nor U2127 (N_2127,N_1662,N_1919);
and U2128 (N_2128,N_1014,N_1707);
nand U2129 (N_2129,N_1750,N_1239);
and U2130 (N_2130,N_1124,N_1964);
nor U2131 (N_2131,N_1650,N_1868);
or U2132 (N_2132,N_1590,N_1794);
nand U2133 (N_2133,N_1013,N_1163);
nand U2134 (N_2134,N_1774,N_1202);
nand U2135 (N_2135,N_1620,N_1286);
or U2136 (N_2136,N_1688,N_1120);
nand U2137 (N_2137,N_1955,N_1218);
or U2138 (N_2138,N_1624,N_1879);
nand U2139 (N_2139,N_1251,N_1075);
nand U2140 (N_2140,N_1257,N_1751);
nand U2141 (N_2141,N_1821,N_1722);
or U2142 (N_2142,N_1734,N_1730);
and U2143 (N_2143,N_1062,N_1745);
nor U2144 (N_2144,N_1936,N_1213);
nor U2145 (N_2145,N_1438,N_1954);
or U2146 (N_2146,N_1888,N_1999);
and U2147 (N_2147,N_1570,N_1334);
nor U2148 (N_2148,N_1992,N_1723);
nor U2149 (N_2149,N_1085,N_1142);
and U2150 (N_2150,N_1260,N_1043);
nor U2151 (N_2151,N_1033,N_1519);
and U2152 (N_2152,N_1413,N_1330);
nor U2153 (N_2153,N_1243,N_1392);
and U2154 (N_2154,N_1912,N_1698);
and U2155 (N_2155,N_1225,N_1869);
and U2156 (N_2156,N_1262,N_1123);
or U2157 (N_2157,N_1030,N_1808);
nor U2158 (N_2158,N_1078,N_1409);
and U2159 (N_2159,N_1939,N_1580);
and U2160 (N_2160,N_1292,N_1510);
nand U2161 (N_2161,N_1719,N_1281);
or U2162 (N_2162,N_1053,N_1140);
nand U2163 (N_2163,N_1876,N_1364);
nand U2164 (N_2164,N_1558,N_1631);
or U2165 (N_2165,N_1343,N_1223);
or U2166 (N_2166,N_1304,N_1569);
nand U2167 (N_2167,N_1982,N_1424);
or U2168 (N_2168,N_1433,N_1741);
nor U2169 (N_2169,N_1350,N_1288);
or U2170 (N_2170,N_1870,N_1214);
nor U2171 (N_2171,N_1695,N_1338);
nand U2172 (N_2172,N_1139,N_1670);
or U2173 (N_2173,N_1403,N_1667);
nand U2174 (N_2174,N_1007,N_1221);
and U2175 (N_2175,N_1086,N_1198);
or U2176 (N_2176,N_1380,N_1162);
and U2177 (N_2177,N_1542,N_1834);
and U2178 (N_2178,N_1386,N_1454);
or U2179 (N_2179,N_1408,N_1359);
nand U2180 (N_2180,N_1932,N_1323);
or U2181 (N_2181,N_1944,N_1259);
nor U2182 (N_2182,N_1857,N_1893);
or U2183 (N_2183,N_1562,N_1980);
and U2184 (N_2184,N_1274,N_1622);
nand U2185 (N_2185,N_1394,N_1527);
or U2186 (N_2186,N_1282,N_1661);
nor U2187 (N_2187,N_1042,N_1490);
xnor U2188 (N_2188,N_1156,N_1178);
nor U2189 (N_2189,N_1475,N_1845);
nand U2190 (N_2190,N_1160,N_1039);
nand U2191 (N_2191,N_1949,N_1756);
and U2192 (N_2192,N_1675,N_1905);
and U2193 (N_2193,N_1792,N_1012);
nand U2194 (N_2194,N_1547,N_1500);
nand U2195 (N_2195,N_1376,N_1995);
nand U2196 (N_2196,N_1523,N_1130);
nor U2197 (N_2197,N_1548,N_1107);
and U2198 (N_2198,N_1689,N_1739);
and U2199 (N_2199,N_1616,N_1382);
nor U2200 (N_2200,N_1147,N_1387);
or U2201 (N_2201,N_1487,N_1708);
and U2202 (N_2202,N_1938,N_1881);
or U2203 (N_2203,N_1602,N_1657);
and U2204 (N_2204,N_1180,N_1066);
nand U2205 (N_2205,N_1143,N_1529);
nand U2206 (N_2206,N_1906,N_1480);
and U2207 (N_2207,N_1333,N_1347);
or U2208 (N_2208,N_1484,N_1928);
or U2209 (N_2209,N_1854,N_1618);
or U2210 (N_2210,N_1754,N_1097);
nand U2211 (N_2211,N_1671,N_1242);
nor U2212 (N_2212,N_1638,N_1728);
nand U2213 (N_2213,N_1862,N_1577);
and U2214 (N_2214,N_1256,N_1501);
or U2215 (N_2215,N_1951,N_1469);
or U2216 (N_2216,N_1472,N_1453);
and U2217 (N_2217,N_1346,N_1886);
nand U2218 (N_2218,N_1199,N_1325);
nor U2219 (N_2219,N_1217,N_1720);
nand U2220 (N_2220,N_1045,N_1904);
xnor U2221 (N_2221,N_1265,N_1781);
and U2222 (N_2222,N_1898,N_1976);
or U2223 (N_2223,N_1089,N_1250);
or U2224 (N_2224,N_1363,N_1154);
nand U2225 (N_2225,N_1761,N_1989);
nor U2226 (N_2226,N_1852,N_1092);
or U2227 (N_2227,N_1950,N_1299);
nand U2228 (N_2228,N_1254,N_1849);
nand U2229 (N_2229,N_1110,N_1512);
and U2230 (N_2230,N_1327,N_1169);
nor U2231 (N_2231,N_1505,N_1310);
or U2232 (N_2232,N_1065,N_1818);
nand U2233 (N_2233,N_1621,N_1172);
nor U2234 (N_2234,N_1405,N_1212);
and U2235 (N_2235,N_1769,N_1451);
nand U2236 (N_2236,N_1112,N_1150);
nand U2237 (N_2237,N_1787,N_1268);
and U2238 (N_2238,N_1416,N_1665);
nand U2239 (N_2239,N_1080,N_1049);
nand U2240 (N_2240,N_1537,N_1219);
nand U2241 (N_2241,N_1578,N_1663);
nand U2242 (N_2242,N_1272,N_1900);
and U2243 (N_2243,N_1915,N_1566);
nand U2244 (N_2244,N_1247,N_1907);
nand U2245 (N_2245,N_1055,N_1832);
or U2246 (N_2246,N_1656,N_1128);
or U2247 (N_2247,N_1489,N_1373);
or U2248 (N_2248,N_1426,N_1494);
and U2249 (N_2249,N_1790,N_1587);
xnor U2250 (N_2250,N_1414,N_1692);
nor U2251 (N_2251,N_1417,N_1693);
nor U2252 (N_2252,N_1320,N_1118);
xor U2253 (N_2253,N_1660,N_1882);
or U2254 (N_2254,N_1877,N_1641);
nand U2255 (N_2255,N_1149,N_1395);
and U2256 (N_2256,N_1492,N_1812);
or U2257 (N_2257,N_1017,N_1589);
nor U2258 (N_2258,N_1666,N_1244);
nand U2259 (N_2259,N_1835,N_1549);
nand U2260 (N_2260,N_1507,N_1399);
nor U2261 (N_2261,N_1113,N_1129);
and U2262 (N_2262,N_1867,N_1036);
and U2263 (N_2263,N_1277,N_1691);
nor U2264 (N_2264,N_1914,N_1674);
and U2265 (N_2265,N_1743,N_1874);
or U2266 (N_2266,N_1962,N_1597);
nor U2267 (N_2267,N_1289,N_1988);
and U2268 (N_2268,N_1360,N_1460);
xor U2269 (N_2269,N_1328,N_1177);
or U2270 (N_2270,N_1673,N_1553);
or U2271 (N_2271,N_1434,N_1933);
nand U2272 (N_2272,N_1028,N_1594);
or U2273 (N_2273,N_1786,N_1138);
or U2274 (N_2274,N_1369,N_1596);
nor U2275 (N_2275,N_1749,N_1785);
and U2276 (N_2276,N_1358,N_1171);
and U2277 (N_2277,N_1306,N_1194);
and U2278 (N_2278,N_1592,N_1427);
and U2279 (N_2279,N_1700,N_1508);
and U2280 (N_2280,N_1541,N_1336);
or U2281 (N_2281,N_1170,N_1034);
or U2282 (N_2282,N_1415,N_1340);
nand U2283 (N_2283,N_1755,N_1206);
or U2284 (N_2284,N_1807,N_1471);
nor U2285 (N_2285,N_1822,N_1210);
nand U2286 (N_2286,N_1771,N_1805);
nor U2287 (N_2287,N_1934,N_1079);
and U2288 (N_2288,N_1355,N_1966);
nor U2289 (N_2289,N_1744,N_1450);
nand U2290 (N_2290,N_1240,N_1010);
and U2291 (N_2291,N_1911,N_1186);
and U2292 (N_2292,N_1967,N_1318);
and U2293 (N_2293,N_1303,N_1132);
and U2294 (N_2294,N_1248,N_1651);
and U2295 (N_2295,N_1195,N_1677);
nor U2296 (N_2296,N_1478,N_1455);
or U2297 (N_2297,N_1891,N_1909);
or U2298 (N_2298,N_1300,N_1102);
nand U2299 (N_2299,N_1724,N_1503);
and U2300 (N_2300,N_1809,N_1696);
nor U2301 (N_2301,N_1998,N_1046);
or U2302 (N_2302,N_1763,N_1583);
nand U2303 (N_2303,N_1008,N_1901);
xnor U2304 (N_2304,N_1362,N_1002);
or U2305 (N_2305,N_1157,N_1071);
and U2306 (N_2306,N_1861,N_1588);
nand U2307 (N_2307,N_1599,N_1356);
nor U2308 (N_2308,N_1488,N_1629);
or U2309 (N_2309,N_1361,N_1099);
xnor U2310 (N_2310,N_1465,N_1913);
or U2311 (N_2311,N_1773,N_1778);
or U2312 (N_2312,N_1483,N_1747);
nand U2313 (N_2313,N_1903,N_1732);
or U2314 (N_2314,N_1804,N_1601);
or U2315 (N_2315,N_1301,N_1844);
or U2316 (N_2316,N_1871,N_1040);
and U2317 (N_2317,N_1461,N_1957);
nor U2318 (N_2318,N_1843,N_1344);
and U2319 (N_2319,N_1803,N_1185);
nor U2320 (N_2320,N_1054,N_1920);
nor U2321 (N_2321,N_1019,N_1319);
nand U2322 (N_2322,N_1561,N_1025);
nor U2323 (N_2323,N_1829,N_1391);
nor U2324 (N_2324,N_1682,N_1109);
xor U2325 (N_2325,N_1735,N_1820);
nor U2326 (N_2326,N_1215,N_1922);
and U2327 (N_2327,N_1859,N_1189);
or U2328 (N_2328,N_1626,N_1517);
or U2329 (N_2329,N_1158,N_1617);
and U2330 (N_2330,N_1379,N_1694);
or U2331 (N_2331,N_1538,N_1593);
and U2332 (N_2332,N_1969,N_1442);
nor U2333 (N_2333,N_1193,N_1144);
nor U2334 (N_2334,N_1481,N_1767);
nor U2335 (N_2335,N_1996,N_1864);
and U2336 (N_2336,N_1757,N_1353);
nand U2337 (N_2337,N_1556,N_1994);
nor U2338 (N_2338,N_1159,N_1041);
nor U2339 (N_2339,N_1902,N_1974);
nand U2340 (N_2340,N_1491,N_1315);
nor U2341 (N_2341,N_1686,N_1275);
nor U2342 (N_2342,N_1623,N_1765);
nand U2343 (N_2343,N_1729,N_1819);
nor U2344 (N_2344,N_1096,N_1793);
nor U2345 (N_2345,N_1005,N_1552);
nor U2346 (N_2346,N_1551,N_1020);
nor U2347 (N_2347,N_1290,N_1390);
nand U2348 (N_2348,N_1298,N_1280);
nor U2349 (N_2349,N_1293,N_1365);
nand U2350 (N_2350,N_1287,N_1585);
or U2351 (N_2351,N_1026,N_1579);
nor U2352 (N_2352,N_1231,N_1001);
or U2353 (N_2353,N_1873,N_1725);
nand U2354 (N_2354,N_1644,N_1679);
or U2355 (N_2355,N_1710,N_1058);
and U2356 (N_2356,N_1841,N_1713);
and U2357 (N_2357,N_1630,N_1227);
or U2358 (N_2358,N_1101,N_1850);
and U2359 (N_2359,N_1374,N_1625);
xor U2360 (N_2360,N_1083,N_1322);
or U2361 (N_2361,N_1420,N_1717);
nand U2362 (N_2362,N_1782,N_1968);
or U2363 (N_2363,N_1015,N_1464);
and U2364 (N_2364,N_1731,N_1305);
or U2365 (N_2365,N_1466,N_1458);
nand U2366 (N_2366,N_1377,N_1190);
and U2367 (N_2367,N_1681,N_1252);
xnor U2368 (N_2368,N_1091,N_1035);
nand U2369 (N_2369,N_1647,N_1152);
and U2370 (N_2370,N_1051,N_1833);
xnor U2371 (N_2371,N_1457,N_1495);
nand U2372 (N_2372,N_1776,N_1332);
nor U2373 (N_2373,N_1883,N_1640);
and U2374 (N_2374,N_1000,N_1216);
nor U2375 (N_2375,N_1817,N_1166);
and U2376 (N_2376,N_1715,N_1752);
or U2377 (N_2377,N_1430,N_1246);
nand U2378 (N_2378,N_1619,N_1106);
nor U2379 (N_2379,N_1357,N_1797);
nand U2380 (N_2380,N_1540,N_1295);
and U2381 (N_2381,N_1991,N_1011);
or U2382 (N_2382,N_1473,N_1878);
nor U2383 (N_2383,N_1582,N_1047);
or U2384 (N_2384,N_1133,N_1165);
nor U2385 (N_2385,N_1436,N_1669);
nand U2386 (N_2386,N_1664,N_1606);
or U2387 (N_2387,N_1515,N_1116);
nand U2388 (N_2388,N_1565,N_1314);
or U2389 (N_2389,N_1191,N_1342);
and U2390 (N_2390,N_1476,N_1368);
or U2391 (N_2391,N_1200,N_1952);
and U2392 (N_2392,N_1435,N_1645);
or U2393 (N_2393,N_1648,N_1052);
nand U2394 (N_2394,N_1308,N_1678);
nor U2395 (N_2395,N_1317,N_1329);
nand U2396 (N_2396,N_1737,N_1241);
or U2397 (N_2397,N_1103,N_1983);
nand U2398 (N_2398,N_1608,N_1872);
nor U2399 (N_2399,N_1067,N_1230);
or U2400 (N_2400,N_1574,N_1470);
nand U2401 (N_2401,N_1179,N_1971);
nor U2402 (N_2402,N_1530,N_1532);
and U2403 (N_2403,N_1572,N_1733);
or U2404 (N_2404,N_1063,N_1273);
nand U2405 (N_2405,N_1712,N_1393);
nand U2406 (N_2406,N_1526,N_1987);
nand U2407 (N_2407,N_1209,N_1009);
nand U2408 (N_2408,N_1764,N_1117);
nor U2409 (N_2409,N_1533,N_1074);
and U2410 (N_2410,N_1897,N_1961);
and U2411 (N_2411,N_1485,N_1563);
nand U2412 (N_2412,N_1550,N_1164);
nand U2413 (N_2413,N_1921,N_1813);
and U2414 (N_2414,N_1655,N_1136);
nand U2415 (N_2415,N_1263,N_1090);
nand U2416 (N_2416,N_1423,N_1772);
or U2417 (N_2417,N_1613,N_1131);
nor U2418 (N_2418,N_1094,N_1060);
nand U2419 (N_2419,N_1959,N_1309);
nand U2420 (N_2420,N_1375,N_1925);
and U2421 (N_2421,N_1701,N_1449);
or U2422 (N_2422,N_1788,N_1497);
or U2423 (N_2423,N_1984,N_1296);
nand U2424 (N_2424,N_1486,N_1525);
nand U2425 (N_2425,N_1126,N_1990);
nor U2426 (N_2426,N_1632,N_1711);
nand U2427 (N_2427,N_1207,N_1294);
or U2428 (N_2428,N_1965,N_1276);
nor U2429 (N_2429,N_1145,N_1652);
nor U2430 (N_2430,N_1479,N_1029);
nor U2431 (N_2431,N_1141,N_1064);
or U2432 (N_2432,N_1429,N_1187);
nand U2433 (N_2433,N_1188,N_1087);
or U2434 (N_2434,N_1923,N_1604);
nand U2435 (N_2435,N_1866,N_1557);
nor U2436 (N_2436,N_1653,N_1775);
nor U2437 (N_2437,N_1238,N_1649);
nand U2438 (N_2438,N_1502,N_1796);
or U2439 (N_2439,N_1806,N_1446);
nand U2440 (N_2440,N_1038,N_1266);
or U2441 (N_2441,N_1456,N_1759);
nor U2442 (N_2442,N_1255,N_1811);
or U2443 (N_2443,N_1801,N_1993);
and U2444 (N_2444,N_1960,N_1245);
or U2445 (N_2445,N_1339,N_1082);
nand U2446 (N_2446,N_1385,N_1279);
nand U2447 (N_2447,N_1341,N_1545);
nand U2448 (N_2448,N_1249,N_1324);
or U2449 (N_2449,N_1412,N_1222);
nor U2450 (N_2450,N_1384,N_1680);
nor U2451 (N_2451,N_1521,N_1718);
or U2452 (N_2452,N_1226,N_1947);
and U2453 (N_2453,N_1699,N_1321);
nor U2454 (N_2454,N_1659,N_1528);
nand U2455 (N_2455,N_1410,N_1205);
and U2456 (N_2456,N_1762,N_1714);
nand U2457 (N_2457,N_1264,N_1611);
and U2458 (N_2458,N_1609,N_1795);
and U2459 (N_2459,N_1351,N_1748);
nand U2460 (N_2460,N_1283,N_1267);
and U2461 (N_2461,N_1402,N_1555);
and U2462 (N_2462,N_1175,N_1258);
nand U2463 (N_2463,N_1468,N_1838);
and U2464 (N_2464,N_1428,N_1847);
nand U2465 (N_2465,N_1331,N_1122);
xnor U2466 (N_2466,N_1840,N_1367);
nor U2467 (N_2467,N_1335,N_1567);
or U2468 (N_2468,N_1404,N_1125);
nor U2469 (N_2469,N_1524,N_1815);
or U2470 (N_2470,N_1894,N_1044);
nand U2471 (N_2471,N_1554,N_1493);
nor U2472 (N_2472,N_1031,N_1291);
nand U2473 (N_2473,N_1513,N_1560);
or U2474 (N_2474,N_1740,N_1985);
and U2475 (N_2475,N_1760,N_1705);
nor U2476 (N_2476,N_1422,N_1848);
nor U2477 (N_2477,N_1658,N_1389);
and U2478 (N_2478,N_1642,N_1016);
or U2479 (N_2479,N_1595,N_1823);
and U2480 (N_2480,N_1463,N_1791);
or U2481 (N_2481,N_1297,N_1006);
nand U2482 (N_2482,N_1134,N_1073);
nor U2483 (N_2483,N_1088,N_1050);
nand U2484 (N_2484,N_1586,N_1977);
and U2485 (N_2485,N_1534,N_1564);
and U2486 (N_2486,N_1600,N_1591);
or U2487 (N_2487,N_1069,N_1726);
or U2488 (N_2488,N_1837,N_1941);
nand U2489 (N_2489,N_1104,N_1736);
and U2490 (N_2490,N_1441,N_1108);
nand U2491 (N_2491,N_1311,N_1196);
or U2492 (N_2492,N_1978,N_1201);
nor U2493 (N_2493,N_1986,N_1603);
and U2494 (N_2494,N_1401,N_1935);
nand U2495 (N_2495,N_1895,N_1037);
nand U2496 (N_2496,N_1768,N_1584);
and U2497 (N_2497,N_1697,N_1024);
nor U2498 (N_2498,N_1783,N_1839);
or U2499 (N_2499,N_1946,N_1183);
nor U2500 (N_2500,N_1168,N_1933);
or U2501 (N_2501,N_1035,N_1422);
and U2502 (N_2502,N_1973,N_1268);
and U2503 (N_2503,N_1319,N_1876);
nor U2504 (N_2504,N_1858,N_1778);
and U2505 (N_2505,N_1505,N_1271);
nor U2506 (N_2506,N_1396,N_1895);
nor U2507 (N_2507,N_1789,N_1240);
nor U2508 (N_2508,N_1352,N_1895);
or U2509 (N_2509,N_1989,N_1496);
or U2510 (N_2510,N_1742,N_1064);
and U2511 (N_2511,N_1503,N_1087);
xor U2512 (N_2512,N_1162,N_1579);
xnor U2513 (N_2513,N_1384,N_1606);
nor U2514 (N_2514,N_1739,N_1191);
or U2515 (N_2515,N_1380,N_1044);
or U2516 (N_2516,N_1497,N_1968);
nor U2517 (N_2517,N_1354,N_1793);
nand U2518 (N_2518,N_1826,N_1979);
nand U2519 (N_2519,N_1002,N_1942);
or U2520 (N_2520,N_1939,N_1744);
or U2521 (N_2521,N_1916,N_1817);
or U2522 (N_2522,N_1391,N_1471);
nor U2523 (N_2523,N_1108,N_1493);
and U2524 (N_2524,N_1252,N_1910);
nand U2525 (N_2525,N_1846,N_1806);
nand U2526 (N_2526,N_1027,N_1260);
nand U2527 (N_2527,N_1166,N_1326);
nor U2528 (N_2528,N_1956,N_1183);
nor U2529 (N_2529,N_1492,N_1817);
nand U2530 (N_2530,N_1138,N_1529);
or U2531 (N_2531,N_1031,N_1203);
nor U2532 (N_2532,N_1976,N_1628);
nor U2533 (N_2533,N_1139,N_1574);
nor U2534 (N_2534,N_1493,N_1497);
or U2535 (N_2535,N_1309,N_1839);
or U2536 (N_2536,N_1995,N_1374);
and U2537 (N_2537,N_1047,N_1964);
or U2538 (N_2538,N_1707,N_1716);
nand U2539 (N_2539,N_1288,N_1398);
and U2540 (N_2540,N_1189,N_1375);
and U2541 (N_2541,N_1680,N_1959);
xor U2542 (N_2542,N_1359,N_1124);
or U2543 (N_2543,N_1513,N_1854);
or U2544 (N_2544,N_1235,N_1646);
and U2545 (N_2545,N_1533,N_1660);
or U2546 (N_2546,N_1009,N_1730);
xnor U2547 (N_2547,N_1142,N_1497);
or U2548 (N_2548,N_1080,N_1191);
nor U2549 (N_2549,N_1539,N_1422);
nor U2550 (N_2550,N_1204,N_1582);
and U2551 (N_2551,N_1715,N_1735);
nand U2552 (N_2552,N_1154,N_1573);
or U2553 (N_2553,N_1080,N_1285);
nand U2554 (N_2554,N_1974,N_1768);
or U2555 (N_2555,N_1963,N_1572);
and U2556 (N_2556,N_1468,N_1701);
nand U2557 (N_2557,N_1250,N_1186);
or U2558 (N_2558,N_1558,N_1432);
and U2559 (N_2559,N_1246,N_1900);
and U2560 (N_2560,N_1368,N_1574);
xor U2561 (N_2561,N_1678,N_1374);
and U2562 (N_2562,N_1695,N_1597);
or U2563 (N_2563,N_1794,N_1458);
nor U2564 (N_2564,N_1490,N_1469);
or U2565 (N_2565,N_1568,N_1780);
and U2566 (N_2566,N_1191,N_1089);
nor U2567 (N_2567,N_1961,N_1199);
and U2568 (N_2568,N_1850,N_1788);
or U2569 (N_2569,N_1318,N_1006);
or U2570 (N_2570,N_1957,N_1043);
or U2571 (N_2571,N_1510,N_1291);
nand U2572 (N_2572,N_1379,N_1458);
or U2573 (N_2573,N_1534,N_1294);
nor U2574 (N_2574,N_1900,N_1781);
nand U2575 (N_2575,N_1613,N_1300);
nor U2576 (N_2576,N_1744,N_1105);
nand U2577 (N_2577,N_1781,N_1277);
and U2578 (N_2578,N_1946,N_1372);
nor U2579 (N_2579,N_1239,N_1459);
or U2580 (N_2580,N_1217,N_1133);
and U2581 (N_2581,N_1136,N_1373);
and U2582 (N_2582,N_1327,N_1777);
nor U2583 (N_2583,N_1531,N_1583);
nand U2584 (N_2584,N_1632,N_1802);
and U2585 (N_2585,N_1593,N_1433);
or U2586 (N_2586,N_1876,N_1229);
nand U2587 (N_2587,N_1954,N_1621);
and U2588 (N_2588,N_1242,N_1980);
or U2589 (N_2589,N_1436,N_1594);
and U2590 (N_2590,N_1909,N_1212);
and U2591 (N_2591,N_1352,N_1693);
and U2592 (N_2592,N_1521,N_1017);
nor U2593 (N_2593,N_1423,N_1884);
and U2594 (N_2594,N_1138,N_1059);
or U2595 (N_2595,N_1038,N_1148);
and U2596 (N_2596,N_1682,N_1240);
or U2597 (N_2597,N_1131,N_1908);
and U2598 (N_2598,N_1742,N_1305);
nor U2599 (N_2599,N_1337,N_1142);
nor U2600 (N_2600,N_1738,N_1987);
nor U2601 (N_2601,N_1786,N_1231);
and U2602 (N_2602,N_1278,N_1775);
nor U2603 (N_2603,N_1956,N_1808);
and U2604 (N_2604,N_1959,N_1585);
or U2605 (N_2605,N_1056,N_1138);
or U2606 (N_2606,N_1299,N_1574);
nand U2607 (N_2607,N_1314,N_1596);
xor U2608 (N_2608,N_1866,N_1556);
or U2609 (N_2609,N_1413,N_1040);
and U2610 (N_2610,N_1304,N_1348);
nor U2611 (N_2611,N_1354,N_1084);
nor U2612 (N_2612,N_1750,N_1811);
or U2613 (N_2613,N_1271,N_1802);
nand U2614 (N_2614,N_1697,N_1657);
and U2615 (N_2615,N_1287,N_1534);
nand U2616 (N_2616,N_1832,N_1186);
nor U2617 (N_2617,N_1038,N_1302);
nor U2618 (N_2618,N_1762,N_1520);
and U2619 (N_2619,N_1067,N_1072);
nor U2620 (N_2620,N_1200,N_1161);
and U2621 (N_2621,N_1773,N_1012);
nor U2622 (N_2622,N_1477,N_1645);
nor U2623 (N_2623,N_1825,N_1024);
and U2624 (N_2624,N_1420,N_1377);
nand U2625 (N_2625,N_1317,N_1507);
nor U2626 (N_2626,N_1581,N_1276);
or U2627 (N_2627,N_1297,N_1158);
nand U2628 (N_2628,N_1432,N_1794);
nand U2629 (N_2629,N_1430,N_1497);
nor U2630 (N_2630,N_1269,N_1769);
nand U2631 (N_2631,N_1132,N_1148);
or U2632 (N_2632,N_1070,N_1215);
nor U2633 (N_2633,N_1921,N_1238);
nor U2634 (N_2634,N_1185,N_1462);
and U2635 (N_2635,N_1805,N_1872);
or U2636 (N_2636,N_1026,N_1274);
or U2637 (N_2637,N_1548,N_1991);
and U2638 (N_2638,N_1629,N_1789);
nor U2639 (N_2639,N_1599,N_1605);
or U2640 (N_2640,N_1828,N_1235);
and U2641 (N_2641,N_1453,N_1229);
nor U2642 (N_2642,N_1829,N_1680);
nor U2643 (N_2643,N_1339,N_1050);
or U2644 (N_2644,N_1874,N_1349);
nand U2645 (N_2645,N_1524,N_1237);
nand U2646 (N_2646,N_1320,N_1691);
nor U2647 (N_2647,N_1750,N_1116);
nand U2648 (N_2648,N_1519,N_1938);
nand U2649 (N_2649,N_1794,N_1020);
or U2650 (N_2650,N_1565,N_1119);
nand U2651 (N_2651,N_1417,N_1501);
nor U2652 (N_2652,N_1239,N_1935);
nor U2653 (N_2653,N_1426,N_1944);
or U2654 (N_2654,N_1813,N_1435);
or U2655 (N_2655,N_1467,N_1621);
and U2656 (N_2656,N_1596,N_1562);
and U2657 (N_2657,N_1403,N_1694);
nand U2658 (N_2658,N_1879,N_1483);
nand U2659 (N_2659,N_1503,N_1770);
and U2660 (N_2660,N_1328,N_1312);
and U2661 (N_2661,N_1137,N_1175);
or U2662 (N_2662,N_1964,N_1300);
nor U2663 (N_2663,N_1772,N_1660);
and U2664 (N_2664,N_1826,N_1517);
nor U2665 (N_2665,N_1970,N_1251);
or U2666 (N_2666,N_1051,N_1351);
or U2667 (N_2667,N_1651,N_1791);
nand U2668 (N_2668,N_1010,N_1769);
or U2669 (N_2669,N_1374,N_1271);
nand U2670 (N_2670,N_1239,N_1088);
nand U2671 (N_2671,N_1297,N_1451);
nand U2672 (N_2672,N_1177,N_1226);
and U2673 (N_2673,N_1399,N_1652);
and U2674 (N_2674,N_1521,N_1839);
nand U2675 (N_2675,N_1864,N_1224);
and U2676 (N_2676,N_1085,N_1988);
and U2677 (N_2677,N_1567,N_1845);
nand U2678 (N_2678,N_1819,N_1539);
nor U2679 (N_2679,N_1321,N_1260);
nand U2680 (N_2680,N_1757,N_1700);
or U2681 (N_2681,N_1576,N_1540);
nor U2682 (N_2682,N_1276,N_1060);
and U2683 (N_2683,N_1605,N_1838);
nand U2684 (N_2684,N_1638,N_1136);
nand U2685 (N_2685,N_1710,N_1875);
nand U2686 (N_2686,N_1847,N_1247);
and U2687 (N_2687,N_1854,N_1215);
nor U2688 (N_2688,N_1678,N_1375);
nor U2689 (N_2689,N_1966,N_1351);
nand U2690 (N_2690,N_1163,N_1495);
or U2691 (N_2691,N_1532,N_1144);
nor U2692 (N_2692,N_1552,N_1490);
nor U2693 (N_2693,N_1472,N_1723);
or U2694 (N_2694,N_1703,N_1512);
and U2695 (N_2695,N_1374,N_1838);
nor U2696 (N_2696,N_1301,N_1231);
or U2697 (N_2697,N_1839,N_1194);
nor U2698 (N_2698,N_1462,N_1374);
nand U2699 (N_2699,N_1189,N_1709);
and U2700 (N_2700,N_1840,N_1006);
nand U2701 (N_2701,N_1837,N_1058);
nor U2702 (N_2702,N_1767,N_1338);
nor U2703 (N_2703,N_1472,N_1846);
nand U2704 (N_2704,N_1774,N_1239);
nand U2705 (N_2705,N_1454,N_1489);
or U2706 (N_2706,N_1721,N_1416);
nand U2707 (N_2707,N_1671,N_1933);
and U2708 (N_2708,N_1214,N_1733);
or U2709 (N_2709,N_1978,N_1821);
nor U2710 (N_2710,N_1789,N_1252);
and U2711 (N_2711,N_1191,N_1408);
and U2712 (N_2712,N_1872,N_1003);
nand U2713 (N_2713,N_1348,N_1758);
nor U2714 (N_2714,N_1202,N_1557);
and U2715 (N_2715,N_1879,N_1923);
nand U2716 (N_2716,N_1598,N_1149);
or U2717 (N_2717,N_1775,N_1527);
nand U2718 (N_2718,N_1133,N_1623);
nand U2719 (N_2719,N_1970,N_1085);
and U2720 (N_2720,N_1565,N_1777);
and U2721 (N_2721,N_1627,N_1417);
nand U2722 (N_2722,N_1965,N_1186);
nor U2723 (N_2723,N_1830,N_1338);
and U2724 (N_2724,N_1159,N_1648);
nand U2725 (N_2725,N_1332,N_1077);
nand U2726 (N_2726,N_1117,N_1158);
nor U2727 (N_2727,N_1970,N_1402);
and U2728 (N_2728,N_1877,N_1872);
nand U2729 (N_2729,N_1333,N_1169);
nand U2730 (N_2730,N_1880,N_1125);
or U2731 (N_2731,N_1885,N_1769);
or U2732 (N_2732,N_1119,N_1991);
or U2733 (N_2733,N_1005,N_1365);
and U2734 (N_2734,N_1555,N_1515);
nand U2735 (N_2735,N_1211,N_1225);
or U2736 (N_2736,N_1546,N_1071);
nor U2737 (N_2737,N_1661,N_1391);
nor U2738 (N_2738,N_1924,N_1109);
nand U2739 (N_2739,N_1234,N_1997);
nor U2740 (N_2740,N_1657,N_1622);
or U2741 (N_2741,N_1285,N_1179);
nand U2742 (N_2742,N_1457,N_1397);
nand U2743 (N_2743,N_1414,N_1160);
or U2744 (N_2744,N_1868,N_1358);
and U2745 (N_2745,N_1392,N_1414);
or U2746 (N_2746,N_1028,N_1121);
xor U2747 (N_2747,N_1242,N_1099);
nand U2748 (N_2748,N_1683,N_1701);
or U2749 (N_2749,N_1516,N_1223);
nor U2750 (N_2750,N_1262,N_1448);
or U2751 (N_2751,N_1800,N_1634);
nand U2752 (N_2752,N_1371,N_1260);
nor U2753 (N_2753,N_1388,N_1988);
nor U2754 (N_2754,N_1791,N_1894);
and U2755 (N_2755,N_1117,N_1182);
and U2756 (N_2756,N_1119,N_1841);
nor U2757 (N_2757,N_1048,N_1890);
nand U2758 (N_2758,N_1053,N_1768);
or U2759 (N_2759,N_1280,N_1227);
or U2760 (N_2760,N_1070,N_1082);
and U2761 (N_2761,N_1633,N_1391);
and U2762 (N_2762,N_1121,N_1463);
nand U2763 (N_2763,N_1222,N_1328);
or U2764 (N_2764,N_1048,N_1655);
nor U2765 (N_2765,N_1236,N_1817);
nand U2766 (N_2766,N_1878,N_1147);
nand U2767 (N_2767,N_1219,N_1231);
or U2768 (N_2768,N_1542,N_1974);
or U2769 (N_2769,N_1143,N_1240);
or U2770 (N_2770,N_1304,N_1960);
nor U2771 (N_2771,N_1519,N_1811);
nor U2772 (N_2772,N_1348,N_1830);
and U2773 (N_2773,N_1294,N_1195);
nand U2774 (N_2774,N_1778,N_1877);
and U2775 (N_2775,N_1637,N_1799);
nand U2776 (N_2776,N_1910,N_1715);
and U2777 (N_2777,N_1974,N_1588);
nor U2778 (N_2778,N_1927,N_1845);
and U2779 (N_2779,N_1481,N_1247);
or U2780 (N_2780,N_1094,N_1249);
and U2781 (N_2781,N_1981,N_1726);
or U2782 (N_2782,N_1696,N_1646);
nor U2783 (N_2783,N_1091,N_1376);
nor U2784 (N_2784,N_1285,N_1605);
or U2785 (N_2785,N_1982,N_1137);
or U2786 (N_2786,N_1416,N_1913);
and U2787 (N_2787,N_1960,N_1555);
nor U2788 (N_2788,N_1697,N_1366);
nor U2789 (N_2789,N_1288,N_1942);
nand U2790 (N_2790,N_1043,N_1965);
or U2791 (N_2791,N_1733,N_1941);
nor U2792 (N_2792,N_1699,N_1515);
or U2793 (N_2793,N_1681,N_1709);
nand U2794 (N_2794,N_1528,N_1523);
nand U2795 (N_2795,N_1539,N_1970);
nor U2796 (N_2796,N_1079,N_1376);
nor U2797 (N_2797,N_1097,N_1709);
and U2798 (N_2798,N_1747,N_1320);
xnor U2799 (N_2799,N_1496,N_1702);
or U2800 (N_2800,N_1300,N_1301);
or U2801 (N_2801,N_1599,N_1256);
nand U2802 (N_2802,N_1727,N_1950);
or U2803 (N_2803,N_1588,N_1303);
or U2804 (N_2804,N_1591,N_1706);
nor U2805 (N_2805,N_1766,N_1036);
nand U2806 (N_2806,N_1345,N_1579);
and U2807 (N_2807,N_1576,N_1887);
nor U2808 (N_2808,N_1407,N_1614);
and U2809 (N_2809,N_1711,N_1158);
nand U2810 (N_2810,N_1738,N_1549);
and U2811 (N_2811,N_1176,N_1973);
nand U2812 (N_2812,N_1758,N_1360);
and U2813 (N_2813,N_1772,N_1947);
xnor U2814 (N_2814,N_1714,N_1133);
nor U2815 (N_2815,N_1128,N_1060);
and U2816 (N_2816,N_1753,N_1170);
nand U2817 (N_2817,N_1981,N_1336);
nor U2818 (N_2818,N_1622,N_1370);
nor U2819 (N_2819,N_1802,N_1931);
or U2820 (N_2820,N_1740,N_1114);
or U2821 (N_2821,N_1651,N_1851);
nand U2822 (N_2822,N_1904,N_1573);
and U2823 (N_2823,N_1544,N_1948);
nand U2824 (N_2824,N_1147,N_1635);
nor U2825 (N_2825,N_1227,N_1387);
nor U2826 (N_2826,N_1714,N_1864);
or U2827 (N_2827,N_1185,N_1562);
or U2828 (N_2828,N_1896,N_1922);
and U2829 (N_2829,N_1337,N_1624);
nor U2830 (N_2830,N_1863,N_1367);
or U2831 (N_2831,N_1556,N_1729);
and U2832 (N_2832,N_1464,N_1236);
nor U2833 (N_2833,N_1230,N_1451);
nand U2834 (N_2834,N_1576,N_1321);
nand U2835 (N_2835,N_1790,N_1489);
nand U2836 (N_2836,N_1624,N_1889);
nand U2837 (N_2837,N_1214,N_1820);
or U2838 (N_2838,N_1520,N_1935);
and U2839 (N_2839,N_1794,N_1909);
and U2840 (N_2840,N_1017,N_1028);
or U2841 (N_2841,N_1056,N_1743);
and U2842 (N_2842,N_1389,N_1628);
and U2843 (N_2843,N_1628,N_1112);
and U2844 (N_2844,N_1600,N_1955);
nand U2845 (N_2845,N_1871,N_1544);
or U2846 (N_2846,N_1176,N_1633);
nand U2847 (N_2847,N_1384,N_1357);
or U2848 (N_2848,N_1873,N_1563);
nor U2849 (N_2849,N_1023,N_1067);
nor U2850 (N_2850,N_1872,N_1108);
or U2851 (N_2851,N_1033,N_1316);
nor U2852 (N_2852,N_1810,N_1953);
or U2853 (N_2853,N_1418,N_1570);
or U2854 (N_2854,N_1790,N_1448);
nor U2855 (N_2855,N_1667,N_1197);
nor U2856 (N_2856,N_1404,N_1959);
nand U2857 (N_2857,N_1143,N_1455);
or U2858 (N_2858,N_1234,N_1999);
or U2859 (N_2859,N_1009,N_1671);
nor U2860 (N_2860,N_1687,N_1206);
nor U2861 (N_2861,N_1094,N_1563);
nand U2862 (N_2862,N_1281,N_1036);
nand U2863 (N_2863,N_1338,N_1192);
or U2864 (N_2864,N_1873,N_1024);
and U2865 (N_2865,N_1740,N_1770);
nor U2866 (N_2866,N_1027,N_1734);
nor U2867 (N_2867,N_1437,N_1526);
nand U2868 (N_2868,N_1177,N_1641);
nand U2869 (N_2869,N_1832,N_1291);
or U2870 (N_2870,N_1653,N_1445);
or U2871 (N_2871,N_1582,N_1631);
nand U2872 (N_2872,N_1723,N_1106);
or U2873 (N_2873,N_1188,N_1162);
and U2874 (N_2874,N_1957,N_1151);
nand U2875 (N_2875,N_1961,N_1894);
nor U2876 (N_2876,N_1422,N_1677);
or U2877 (N_2877,N_1259,N_1424);
nand U2878 (N_2878,N_1422,N_1849);
nor U2879 (N_2879,N_1584,N_1767);
nand U2880 (N_2880,N_1895,N_1269);
and U2881 (N_2881,N_1773,N_1982);
xor U2882 (N_2882,N_1645,N_1763);
and U2883 (N_2883,N_1708,N_1739);
nor U2884 (N_2884,N_1451,N_1360);
nand U2885 (N_2885,N_1834,N_1821);
and U2886 (N_2886,N_1473,N_1955);
nand U2887 (N_2887,N_1833,N_1928);
and U2888 (N_2888,N_1022,N_1670);
and U2889 (N_2889,N_1017,N_1261);
or U2890 (N_2890,N_1089,N_1736);
nor U2891 (N_2891,N_1582,N_1104);
nor U2892 (N_2892,N_1941,N_1312);
nor U2893 (N_2893,N_1754,N_1465);
nor U2894 (N_2894,N_1304,N_1036);
or U2895 (N_2895,N_1749,N_1392);
or U2896 (N_2896,N_1094,N_1100);
nor U2897 (N_2897,N_1819,N_1756);
and U2898 (N_2898,N_1045,N_1192);
and U2899 (N_2899,N_1435,N_1905);
nor U2900 (N_2900,N_1603,N_1555);
nor U2901 (N_2901,N_1812,N_1664);
and U2902 (N_2902,N_1869,N_1743);
nand U2903 (N_2903,N_1854,N_1107);
xnor U2904 (N_2904,N_1796,N_1413);
and U2905 (N_2905,N_1237,N_1651);
nor U2906 (N_2906,N_1247,N_1267);
nor U2907 (N_2907,N_1481,N_1795);
nand U2908 (N_2908,N_1497,N_1501);
or U2909 (N_2909,N_1921,N_1026);
and U2910 (N_2910,N_1947,N_1619);
nand U2911 (N_2911,N_1485,N_1204);
or U2912 (N_2912,N_1789,N_1835);
nor U2913 (N_2913,N_1660,N_1731);
nor U2914 (N_2914,N_1190,N_1143);
or U2915 (N_2915,N_1407,N_1989);
or U2916 (N_2916,N_1329,N_1138);
nand U2917 (N_2917,N_1985,N_1957);
nor U2918 (N_2918,N_1922,N_1455);
nor U2919 (N_2919,N_1781,N_1414);
nor U2920 (N_2920,N_1961,N_1855);
nand U2921 (N_2921,N_1966,N_1056);
nor U2922 (N_2922,N_1524,N_1888);
xnor U2923 (N_2923,N_1880,N_1686);
or U2924 (N_2924,N_1940,N_1943);
nand U2925 (N_2925,N_1930,N_1089);
nor U2926 (N_2926,N_1738,N_1868);
and U2927 (N_2927,N_1943,N_1369);
or U2928 (N_2928,N_1677,N_1275);
nand U2929 (N_2929,N_1186,N_1675);
and U2930 (N_2930,N_1338,N_1293);
nor U2931 (N_2931,N_1723,N_1852);
or U2932 (N_2932,N_1577,N_1637);
nand U2933 (N_2933,N_1227,N_1318);
nand U2934 (N_2934,N_1161,N_1243);
nand U2935 (N_2935,N_1609,N_1553);
and U2936 (N_2936,N_1306,N_1007);
or U2937 (N_2937,N_1330,N_1779);
nand U2938 (N_2938,N_1681,N_1360);
and U2939 (N_2939,N_1832,N_1851);
or U2940 (N_2940,N_1150,N_1794);
nand U2941 (N_2941,N_1663,N_1401);
nand U2942 (N_2942,N_1520,N_1180);
nor U2943 (N_2943,N_1295,N_1444);
and U2944 (N_2944,N_1889,N_1211);
nor U2945 (N_2945,N_1817,N_1255);
or U2946 (N_2946,N_1475,N_1818);
nor U2947 (N_2947,N_1980,N_1785);
nor U2948 (N_2948,N_1835,N_1871);
nand U2949 (N_2949,N_1743,N_1841);
nor U2950 (N_2950,N_1760,N_1751);
or U2951 (N_2951,N_1899,N_1694);
and U2952 (N_2952,N_1165,N_1783);
and U2953 (N_2953,N_1315,N_1454);
or U2954 (N_2954,N_1116,N_1947);
nand U2955 (N_2955,N_1170,N_1721);
nor U2956 (N_2956,N_1001,N_1007);
nor U2957 (N_2957,N_1508,N_1855);
or U2958 (N_2958,N_1609,N_1542);
or U2959 (N_2959,N_1948,N_1269);
or U2960 (N_2960,N_1822,N_1296);
nand U2961 (N_2961,N_1148,N_1243);
nor U2962 (N_2962,N_1130,N_1448);
nor U2963 (N_2963,N_1953,N_1635);
and U2964 (N_2964,N_1146,N_1636);
and U2965 (N_2965,N_1903,N_1801);
nor U2966 (N_2966,N_1394,N_1720);
and U2967 (N_2967,N_1979,N_1729);
nor U2968 (N_2968,N_1954,N_1254);
nor U2969 (N_2969,N_1017,N_1400);
and U2970 (N_2970,N_1341,N_1655);
nor U2971 (N_2971,N_1161,N_1366);
or U2972 (N_2972,N_1123,N_1310);
or U2973 (N_2973,N_1150,N_1429);
or U2974 (N_2974,N_1731,N_1686);
nor U2975 (N_2975,N_1366,N_1354);
nor U2976 (N_2976,N_1409,N_1423);
and U2977 (N_2977,N_1970,N_1404);
nand U2978 (N_2978,N_1019,N_1720);
and U2979 (N_2979,N_1000,N_1485);
or U2980 (N_2980,N_1937,N_1226);
nand U2981 (N_2981,N_1523,N_1730);
or U2982 (N_2982,N_1981,N_1229);
or U2983 (N_2983,N_1759,N_1460);
or U2984 (N_2984,N_1189,N_1422);
and U2985 (N_2985,N_1626,N_1955);
nand U2986 (N_2986,N_1234,N_1628);
and U2987 (N_2987,N_1634,N_1226);
xor U2988 (N_2988,N_1968,N_1989);
nor U2989 (N_2989,N_1973,N_1732);
or U2990 (N_2990,N_1569,N_1603);
and U2991 (N_2991,N_1873,N_1871);
or U2992 (N_2992,N_1740,N_1694);
and U2993 (N_2993,N_1694,N_1236);
and U2994 (N_2994,N_1655,N_1424);
or U2995 (N_2995,N_1464,N_1769);
and U2996 (N_2996,N_1551,N_1574);
nor U2997 (N_2997,N_1808,N_1508);
nand U2998 (N_2998,N_1851,N_1335);
or U2999 (N_2999,N_1019,N_1847);
nor U3000 (N_3000,N_2151,N_2610);
or U3001 (N_3001,N_2917,N_2464);
nand U3002 (N_3002,N_2758,N_2815);
nand U3003 (N_3003,N_2527,N_2003);
or U3004 (N_3004,N_2104,N_2285);
nand U3005 (N_3005,N_2178,N_2352);
nand U3006 (N_3006,N_2692,N_2969);
or U3007 (N_3007,N_2417,N_2712);
and U3008 (N_3008,N_2592,N_2273);
nand U3009 (N_3009,N_2808,N_2000);
nand U3010 (N_3010,N_2287,N_2376);
nor U3011 (N_3011,N_2588,N_2092);
or U3012 (N_3012,N_2233,N_2560);
nor U3013 (N_3013,N_2910,N_2659);
xnor U3014 (N_3014,N_2813,N_2223);
nor U3015 (N_3015,N_2451,N_2792);
nor U3016 (N_3016,N_2953,N_2165);
or U3017 (N_3017,N_2374,N_2900);
or U3018 (N_3018,N_2097,N_2932);
or U3019 (N_3019,N_2617,N_2749);
nand U3020 (N_3020,N_2055,N_2909);
nor U3021 (N_3021,N_2234,N_2961);
and U3022 (N_3022,N_2257,N_2978);
nor U3023 (N_3023,N_2553,N_2936);
nor U3024 (N_3024,N_2486,N_2912);
nand U3025 (N_3025,N_2558,N_2297);
nor U3026 (N_3026,N_2227,N_2767);
or U3027 (N_3027,N_2479,N_2773);
and U3028 (N_3028,N_2298,N_2720);
nor U3029 (N_3029,N_2728,N_2838);
nand U3030 (N_3030,N_2741,N_2312);
nand U3031 (N_3031,N_2836,N_2807);
nand U3032 (N_3032,N_2511,N_2576);
and U3033 (N_3033,N_2131,N_2389);
and U3034 (N_3034,N_2076,N_2409);
or U3035 (N_3035,N_2256,N_2655);
nand U3036 (N_3036,N_2858,N_2426);
nand U3037 (N_3037,N_2416,N_2149);
nor U3038 (N_3038,N_2864,N_2848);
or U3039 (N_3039,N_2860,N_2137);
or U3040 (N_3040,N_2489,N_2595);
nor U3041 (N_3041,N_2903,N_2011);
or U3042 (N_3042,N_2517,N_2455);
nand U3043 (N_3043,N_2252,N_2843);
nor U3044 (N_3044,N_2032,N_2648);
nor U3045 (N_3045,N_2759,N_2056);
nor U3046 (N_3046,N_2791,N_2533);
or U3047 (N_3047,N_2545,N_2833);
and U3048 (N_3048,N_2886,N_2070);
and U3049 (N_3049,N_2316,N_2265);
nor U3050 (N_3050,N_2962,N_2362);
xnor U3051 (N_3051,N_2038,N_2259);
and U3052 (N_3052,N_2211,N_2125);
and U3053 (N_3053,N_2872,N_2048);
nand U3054 (N_3054,N_2831,N_2175);
and U3055 (N_3055,N_2616,N_2529);
nand U3056 (N_3056,N_2340,N_2508);
nand U3057 (N_3057,N_2505,N_2307);
and U3058 (N_3058,N_2667,N_2779);
or U3059 (N_3059,N_2201,N_2447);
nor U3060 (N_3060,N_2103,N_2670);
and U3061 (N_3061,N_2295,N_2793);
and U3062 (N_3062,N_2320,N_2706);
nand U3063 (N_3063,N_2929,N_2817);
nand U3064 (N_3064,N_2777,N_2168);
and U3065 (N_3065,N_2005,N_2493);
nand U3066 (N_3066,N_2857,N_2315);
or U3067 (N_3067,N_2629,N_2523);
or U3068 (N_3068,N_2457,N_2448);
nor U3069 (N_3069,N_2786,N_2124);
nor U3070 (N_3070,N_2608,N_2439);
nor U3071 (N_3071,N_2438,N_2141);
nor U3072 (N_3072,N_2769,N_2713);
and U3073 (N_3073,N_2431,N_2377);
or U3074 (N_3074,N_2441,N_2206);
nand U3075 (N_3075,N_2427,N_2332);
and U3076 (N_3076,N_2901,N_2108);
nor U3077 (N_3077,N_2618,N_2981);
or U3078 (N_3078,N_2293,N_2499);
or U3079 (N_3079,N_2844,N_2009);
or U3080 (N_3080,N_2171,N_2771);
nand U3081 (N_3081,N_2437,N_2622);
and U3082 (N_3082,N_2044,N_2176);
or U3083 (N_3083,N_2361,N_2931);
and U3084 (N_3084,N_2536,N_2509);
or U3085 (N_3085,N_2550,N_2222);
nor U3086 (N_3086,N_2760,N_2270);
nand U3087 (N_3087,N_2572,N_2944);
nand U3088 (N_3088,N_2326,N_2183);
nor U3089 (N_3089,N_2675,N_2887);
nor U3090 (N_3090,N_2145,N_2753);
or U3091 (N_3091,N_2244,N_2894);
and U3092 (N_3092,N_2300,N_2415);
or U3093 (N_3093,N_2065,N_2952);
and U3094 (N_3094,N_2161,N_2650);
nand U3095 (N_3095,N_2896,N_2224);
nand U3096 (N_3096,N_2094,N_2294);
or U3097 (N_3097,N_2052,N_2991);
and U3098 (N_3098,N_2232,N_2513);
nand U3099 (N_3099,N_2177,N_2845);
and U3100 (N_3100,N_2724,N_2875);
or U3101 (N_3101,N_2794,N_2620);
and U3102 (N_3102,N_2174,N_2189);
nand U3103 (N_3103,N_2840,N_2449);
nor U3104 (N_3104,N_2306,N_2481);
nand U3105 (N_3105,N_2026,N_2333);
or U3106 (N_3106,N_2263,N_2514);
or U3107 (N_3107,N_2642,N_2601);
nand U3108 (N_3108,N_2852,N_2080);
or U3109 (N_3109,N_2585,N_2869);
and U3110 (N_3110,N_2460,N_2207);
nand U3111 (N_3111,N_2353,N_2812);
or U3112 (N_3112,N_2990,N_2391);
nand U3113 (N_3113,N_2384,N_2686);
and U3114 (N_3114,N_2017,N_2607);
nor U3115 (N_3115,N_2275,N_2614);
or U3116 (N_3116,N_2379,N_2682);
and U3117 (N_3117,N_2129,N_2619);
nand U3118 (N_3118,N_2700,N_2693);
or U3119 (N_3119,N_2491,N_2940);
and U3120 (N_3120,N_2243,N_2945);
nor U3121 (N_3121,N_2877,N_2281);
xor U3122 (N_3122,N_2407,N_2898);
nor U3123 (N_3123,N_2213,N_2110);
and U3124 (N_3124,N_2630,N_2640);
nor U3125 (N_3125,N_2762,N_2819);
nand U3126 (N_3126,N_2816,N_2106);
and U3127 (N_3127,N_2229,N_2412);
nor U3128 (N_3128,N_2078,N_2107);
nand U3129 (N_3129,N_2747,N_2600);
or U3130 (N_3130,N_2182,N_2972);
nand U3131 (N_3131,N_2347,N_2564);
nand U3132 (N_3132,N_2188,N_2432);
or U3133 (N_3133,N_2568,N_2378);
nand U3134 (N_3134,N_2166,N_2837);
nor U3135 (N_3135,N_2299,N_2488);
nand U3136 (N_3136,N_2268,N_2049);
or U3137 (N_3137,N_2956,N_2975);
or U3138 (N_3138,N_2995,N_2450);
nand U3139 (N_3139,N_2043,N_2500);
nand U3140 (N_3140,N_2050,N_2388);
or U3141 (N_3141,N_2718,N_2756);
and U3142 (N_3142,N_2475,N_2521);
nand U3143 (N_3143,N_2633,N_2160);
or U3144 (N_3144,N_2212,N_2696);
nor U3145 (N_3145,N_2238,N_2789);
or U3146 (N_3146,N_2284,N_2606);
or U3147 (N_3147,N_2582,N_2249);
and U3148 (N_3148,N_2661,N_2303);
or U3149 (N_3149,N_2856,N_2590);
nor U3150 (N_3150,N_2704,N_2539);
and U3151 (N_3151,N_2541,N_2918);
or U3152 (N_3152,N_2459,N_2750);
and U3153 (N_3153,N_2001,N_2863);
nor U3154 (N_3154,N_2302,N_2531);
and U3155 (N_3155,N_2904,N_2507);
nand U3156 (N_3156,N_2878,N_2943);
nor U3157 (N_3157,N_2116,N_2102);
or U3158 (N_3158,N_2370,N_2308);
and U3159 (N_3159,N_2986,N_2751);
and U3160 (N_3160,N_2069,N_2034);
nor U3161 (N_3161,N_2784,N_2429);
nand U3162 (N_3162,N_2136,N_2854);
nand U3163 (N_3163,N_2061,N_2716);
nand U3164 (N_3164,N_2732,N_2057);
and U3165 (N_3165,N_2935,N_2355);
or U3166 (N_3166,N_2323,N_2472);
or U3167 (N_3167,N_2520,N_2674);
nor U3168 (N_3168,N_2556,N_2804);
or U3169 (N_3169,N_2310,N_2077);
nor U3170 (N_3170,N_2827,N_2025);
nand U3171 (N_3171,N_2707,N_2516);
nor U3172 (N_3172,N_2525,N_2660);
nor U3173 (N_3173,N_2778,N_2487);
or U3174 (N_3174,N_2510,N_2698);
nand U3175 (N_3175,N_2369,N_2825);
nand U3176 (N_3176,N_2730,N_2989);
or U3177 (N_3177,N_2597,N_2113);
or U3178 (N_3178,N_2859,N_2906);
or U3179 (N_3179,N_2433,N_2949);
or U3180 (N_3180,N_2652,N_2383);
nor U3181 (N_3181,N_2645,N_2835);
nand U3182 (N_3182,N_2334,N_2911);
nor U3183 (N_3183,N_2428,N_2461);
or U3184 (N_3184,N_2723,N_2882);
or U3185 (N_3185,N_2470,N_2013);
nand U3186 (N_3186,N_2423,N_2084);
nor U3187 (N_3187,N_2360,N_2914);
or U3188 (N_3188,N_2088,N_2186);
or U3189 (N_3189,N_2130,N_2871);
xnor U3190 (N_3190,N_2466,N_2811);
or U3191 (N_3191,N_2566,N_2734);
or U3192 (N_3192,N_2480,N_2555);
nand U3193 (N_3193,N_2714,N_2276);
and U3194 (N_3194,N_2185,N_2037);
nand U3195 (N_3195,N_2963,N_2471);
or U3196 (N_3196,N_2853,N_2846);
or U3197 (N_3197,N_2537,N_2715);
nor U3198 (N_3198,N_2795,N_2063);
nor U3199 (N_3199,N_2436,N_2473);
nand U3200 (N_3200,N_2452,N_2635);
or U3201 (N_3201,N_2549,N_2913);
or U3202 (N_3202,N_2062,N_2885);
nand U3203 (N_3203,N_2271,N_2279);
or U3204 (N_3204,N_2970,N_2678);
nor U3205 (N_3205,N_2538,N_2602);
or U3206 (N_3206,N_2283,N_2033);
and U3207 (N_3207,N_2515,N_2198);
and U3208 (N_3208,N_2982,N_2385);
and U3209 (N_3209,N_2120,N_2221);
and U3210 (N_3210,N_2163,N_2478);
nor U3211 (N_3211,N_2651,N_2408);
nand U3212 (N_3212,N_2623,N_2023);
or U3213 (N_3213,N_2357,N_2624);
nor U3214 (N_3214,N_2689,N_2386);
nor U3215 (N_3215,N_2775,N_2117);
nor U3216 (N_3216,N_2880,N_2096);
and U3217 (N_3217,N_2596,N_2787);
nor U3218 (N_3218,N_2567,N_2147);
nor U3219 (N_3219,N_2274,N_2327);
nor U3220 (N_3220,N_2121,N_2519);
or U3221 (N_3221,N_2208,N_2925);
nand U3222 (N_3222,N_2868,N_2960);
or U3223 (N_3223,N_2167,N_2483);
nand U3224 (N_3224,N_2095,N_2824);
and U3225 (N_3225,N_2637,N_2994);
nand U3226 (N_3226,N_2364,N_2041);
nand U3227 (N_3227,N_2143,N_2035);
or U3228 (N_3228,N_2855,N_2593);
or U3229 (N_3229,N_2122,N_2810);
and U3230 (N_3230,N_2641,N_2251);
or U3231 (N_3231,N_2939,N_2395);
nand U3232 (N_3232,N_2926,N_2586);
nor U3233 (N_3233,N_2318,N_2047);
nand U3234 (N_3234,N_2397,N_2228);
nand U3235 (N_3235,N_2598,N_2218);
and U3236 (N_3236,N_2403,N_2892);
nand U3237 (N_3237,N_2456,N_2351);
and U3238 (N_3238,N_2705,N_2322);
or U3239 (N_3239,N_2862,N_2764);
and U3240 (N_3240,N_2286,N_2304);
and U3241 (N_3241,N_2742,N_2317);
nor U3242 (N_3242,N_2551,N_2059);
or U3243 (N_3243,N_2691,N_2087);
or U3244 (N_3244,N_2446,N_2090);
nor U3245 (N_3245,N_2669,N_2031);
or U3246 (N_3246,N_2973,N_2468);
nor U3247 (N_3247,N_2123,N_2162);
nor U3248 (N_3248,N_2611,N_2266);
nand U3249 (N_3249,N_2703,N_2899);
nor U3250 (N_3250,N_2802,N_2766);
and U3251 (N_3251,N_2225,N_2851);
or U3252 (N_3252,N_2923,N_2280);
or U3253 (N_3253,N_2893,N_2927);
nor U3254 (N_3254,N_2993,N_2202);
nor U3255 (N_3255,N_2905,N_2425);
nand U3256 (N_3256,N_2947,N_2343);
or U3257 (N_3257,N_2921,N_2561);
nor U3258 (N_3258,N_2115,N_2976);
and U3259 (N_3259,N_2242,N_2656);
or U3260 (N_3260,N_2609,N_2027);
and U3261 (N_3261,N_2150,N_2337);
or U3262 (N_3262,N_2967,N_2241);
and U3263 (N_3263,N_2979,N_2396);
nand U3264 (N_3264,N_2170,N_2677);
or U3265 (N_3265,N_2405,N_2870);
nand U3266 (N_3266,N_2540,N_2876);
nor U3267 (N_3267,N_2554,N_2688);
and U3268 (N_3268,N_2255,N_2021);
nor U3269 (N_3269,N_2068,N_2890);
nor U3270 (N_3270,N_2442,N_2731);
or U3271 (N_3271,N_2022,N_2010);
nor U3272 (N_3272,N_2098,N_2954);
nand U3273 (N_3273,N_2269,N_2443);
nor U3274 (N_3274,N_2319,N_2546);
or U3275 (N_3275,N_2687,N_2371);
nor U3276 (N_3276,N_2400,N_2955);
or U3277 (N_3277,N_2019,N_2799);
and U3278 (N_3278,N_2654,N_2072);
and U3279 (N_3279,N_2339,N_2708);
nor U3280 (N_3280,N_2613,N_2236);
nand U3281 (N_3281,N_2577,N_2559);
nor U3282 (N_3282,N_2435,N_2359);
xnor U3283 (N_3283,N_2148,N_2235);
or U3284 (N_3284,N_2100,N_2354);
and U3285 (N_3285,N_2702,N_2336);
nand U3286 (N_3286,N_2153,N_2644);
nor U3287 (N_3287,N_2544,N_2373);
or U3288 (N_3288,N_2342,N_2458);
nor U3289 (N_3289,N_2946,N_2562);
and U3290 (N_3290,N_2467,N_2746);
nor U3291 (N_3291,N_2528,N_2016);
and U3292 (N_3292,N_2058,N_2152);
nor U3293 (N_3293,N_2997,N_2192);
or U3294 (N_3294,N_2366,N_2727);
or U3295 (N_3295,N_2980,N_2745);
nor U3296 (N_3296,N_2169,N_2101);
or U3297 (N_3297,N_2245,N_2144);
or U3298 (N_3298,N_2282,N_2114);
or U3299 (N_3299,N_2462,N_2127);
and U3300 (N_3300,N_2907,N_2335);
nor U3301 (N_3301,N_2411,N_2007);
and U3302 (N_3302,N_2823,N_2413);
nand U3303 (N_3303,N_2030,N_2599);
nand U3304 (N_3304,N_2889,N_2998);
or U3305 (N_3305,N_2552,N_2226);
nand U3306 (N_3306,N_2649,N_2180);
or U3307 (N_3307,N_2119,N_2179);
and U3308 (N_3308,N_2289,N_2676);
and U3309 (N_3309,N_2134,N_2673);
or U3310 (N_3310,N_2584,N_2111);
nand U3311 (N_3311,N_2250,N_2805);
or U3312 (N_3312,N_2053,N_2841);
or U3313 (N_3313,N_2064,N_2757);
and U3314 (N_3314,N_2082,N_2679);
or U3315 (N_3315,N_2338,N_2341);
nand U3316 (N_3316,N_2490,N_2164);
or U3317 (N_3317,N_2197,N_2205);
or U3318 (N_3318,N_2512,N_2574);
nor U3319 (N_3319,N_2463,N_2783);
nand U3320 (N_3320,N_2496,N_2083);
nand U3321 (N_3321,N_2847,N_2958);
nor U3322 (N_3322,N_2381,N_2085);
nor U3323 (N_3323,N_2663,N_2133);
or U3324 (N_3324,N_2522,N_2262);
or U3325 (N_3325,N_2135,N_2938);
and U3326 (N_3326,N_2036,N_2701);
nor U3327 (N_3327,N_2631,N_2220);
nor U3328 (N_3328,N_2191,N_2173);
nand U3329 (N_3329,N_2798,N_2996);
nand U3330 (N_3330,N_2748,N_2331);
nand U3331 (N_3331,N_2004,N_2722);
and U3332 (N_3332,N_2638,N_2419);
or U3333 (N_3333,N_2612,N_2046);
nor U3334 (N_3334,N_2401,N_2542);
and U3335 (N_3335,N_2012,N_2888);
nand U3336 (N_3336,N_2203,N_2781);
and U3337 (N_3337,N_2261,N_2184);
and U3338 (N_3338,N_2985,N_2711);
nor U3339 (N_3339,N_2328,N_2363);
nor U3340 (N_3340,N_2915,N_2726);
nand U3341 (N_3341,N_2344,N_2492);
nand U3342 (N_3342,N_2765,N_2482);
or U3343 (N_3343,N_2345,N_2404);
and U3344 (N_3344,N_2603,N_2028);
nor U3345 (N_3345,N_2934,N_2636);
nand U3346 (N_3346,N_2504,N_2140);
or U3347 (N_3347,N_2666,N_2814);
or U3348 (N_3348,N_2821,N_2356);
and U3349 (N_3349,N_2776,N_2964);
nand U3350 (N_3350,N_2524,N_2440);
nor U3351 (N_3351,N_2729,N_2215);
nor U3352 (N_3352,N_2420,N_2358);
nand U3353 (N_3353,N_2685,N_2755);
nor U3354 (N_3354,N_2752,N_2658);
or U3355 (N_3355,N_2216,N_2118);
nand U3356 (N_3356,N_2563,N_2879);
or U3357 (N_3357,N_2253,N_2465);
nand U3358 (N_3358,N_2625,N_2365);
and U3359 (N_3359,N_2190,N_2829);
or U3360 (N_3360,N_2089,N_2763);
or U3361 (N_3361,N_2782,N_2959);
and U3362 (N_3362,N_2581,N_2690);
or U3363 (N_3363,N_2329,N_2210);
nand U3364 (N_3364,N_2534,N_2067);
or U3365 (N_3365,N_2424,N_2453);
or U3366 (N_3366,N_2497,N_2834);
nand U3367 (N_3367,N_2393,N_2040);
or U3368 (N_3368,N_2296,N_2494);
nand U3369 (N_3369,N_2873,N_2313);
nor U3370 (N_3370,N_2474,N_2039);
and U3371 (N_3371,N_2739,N_2951);
or U3372 (N_3372,N_2091,N_2809);
nor U3373 (N_3373,N_2941,N_2006);
and U3374 (N_3374,N_2414,N_2800);
nor U3375 (N_3375,N_2883,N_2719);
nand U3376 (N_3376,N_2818,N_2024);
and U3377 (N_3377,N_2867,N_2231);
xnor U3378 (N_3378,N_2736,N_2430);
nor U3379 (N_3379,N_2093,N_2790);
and U3380 (N_3380,N_2849,N_2671);
and U3381 (N_3381,N_2485,N_2785);
nor U3382 (N_3382,N_2382,N_2881);
and U3383 (N_3383,N_2874,N_2984);
or U3384 (N_3384,N_2589,N_2288);
or U3385 (N_3385,N_2272,N_2948);
nand U3386 (N_3386,N_2128,N_2254);
and U3387 (N_3387,N_2583,N_2683);
and U3388 (N_3388,N_2394,N_2621);
nor U3389 (N_3389,N_2662,N_2350);
nor U3390 (N_3390,N_2291,N_2780);
or U3391 (N_3391,N_2657,N_2375);
or U3392 (N_3392,N_2842,N_2977);
nand U3393 (N_3393,N_2806,N_2647);
and U3394 (N_3394,N_2737,N_2526);
nand U3395 (N_3395,N_2664,N_2247);
or U3396 (N_3396,N_2548,N_2725);
nand U3397 (N_3397,N_2797,N_2126);
or U3398 (N_3398,N_2684,N_2421);
nand U3399 (N_3399,N_2015,N_2074);
nor U3400 (N_3400,N_2680,N_2081);
nor U3401 (N_3401,N_2916,N_2733);
or U3402 (N_3402,N_2754,N_2073);
and U3403 (N_3403,N_2695,N_2158);
or U3404 (N_3404,N_2897,N_2278);
nor U3405 (N_3405,N_2042,N_2957);
and U3406 (N_3406,N_2109,N_2861);
nand U3407 (N_3407,N_2258,N_2761);
or U3408 (N_3408,N_2579,N_2214);
and U3409 (N_3409,N_2099,N_2665);
and U3410 (N_3410,N_2950,N_2305);
nor U3411 (N_3411,N_2721,N_2498);
xnor U3412 (N_3412,N_2418,N_2587);
nand U3413 (N_3413,N_2681,N_2992);
or U3414 (N_3414,N_2591,N_2142);
and U3415 (N_3415,N_2830,N_2292);
nor U3416 (N_3416,N_2477,N_2246);
nor U3417 (N_3417,N_2054,N_2155);
nand U3418 (N_3418,N_2902,N_2971);
nor U3419 (N_3419,N_2699,N_2828);
nor U3420 (N_3420,N_2768,N_2387);
or U3421 (N_3421,N_2146,N_2930);
and U3422 (N_3422,N_2196,N_2735);
nand U3423 (N_3423,N_2646,N_2919);
nand U3424 (N_3424,N_2820,N_2965);
or U3425 (N_3425,N_2002,N_2324);
and U3426 (N_3426,N_2105,N_2573);
nor U3427 (N_3427,N_2788,N_2518);
nand U3428 (N_3428,N_2264,N_2398);
nor U3429 (N_3429,N_2924,N_2014);
nand U3430 (N_3430,N_2571,N_2071);
and U3431 (N_3431,N_2346,N_2066);
or U3432 (N_3432,N_2372,N_2639);
or U3433 (N_3433,N_2248,N_2632);
or U3434 (N_3434,N_2045,N_2410);
and U3435 (N_3435,N_2260,N_2501);
nor U3436 (N_3436,N_2209,N_2772);
nor U3437 (N_3437,N_2740,N_2839);
or U3438 (N_3438,N_2826,N_2301);
and U3439 (N_3439,N_2634,N_2454);
and U3440 (N_3440,N_2895,N_2569);
nand U3441 (N_3441,N_2543,N_2928);
or U3442 (N_3442,N_2204,N_2311);
nand U3443 (N_3443,N_2503,N_2132);
or U3444 (N_3444,N_2668,N_2187);
nor U3445 (N_3445,N_2694,N_2193);
and U3446 (N_3446,N_2277,N_2942);
nor U3447 (N_3447,N_2392,N_2506);
or U3448 (N_3448,N_2349,N_2709);
or U3449 (N_3449,N_2051,N_2230);
and U3450 (N_3450,N_2615,N_2822);
and U3451 (N_3451,N_2217,N_2968);
nor U3452 (N_3452,N_2974,N_2884);
xnor U3453 (N_3453,N_2139,N_2181);
and U3454 (N_3454,N_2570,N_2200);
nor U3455 (N_3455,N_2626,N_2801);
or U3456 (N_3456,N_2348,N_2380);
nand U3457 (N_3457,N_2159,N_2653);
nand U3458 (N_3458,N_2445,N_2484);
and U3459 (N_3459,N_2469,N_2770);
nor U3460 (N_3460,N_2075,N_2239);
nand U3461 (N_3461,N_2643,N_2154);
and U3462 (N_3462,N_2565,N_2434);
or U3463 (N_3463,N_2743,N_2983);
and U3464 (N_3464,N_2717,N_2156);
nand U3465 (N_3465,N_2219,N_2672);
and U3466 (N_3466,N_2240,N_2138);
nor U3467 (N_3467,N_2476,N_2086);
and U3468 (N_3468,N_2891,N_2920);
and U3469 (N_3469,N_2325,N_2194);
nand U3470 (N_3470,N_2422,N_2988);
nor U3471 (N_3471,N_2697,N_2399);
or U3472 (N_3472,N_2390,N_2195);
or U3473 (N_3473,N_2367,N_2502);
and U3474 (N_3474,N_2605,N_2157);
or U3475 (N_3475,N_2237,N_2079);
and U3476 (N_3476,N_2020,N_2199);
nand U3477 (N_3477,N_2832,N_2744);
or U3478 (N_3478,N_2966,N_2803);
nand U3479 (N_3479,N_2060,N_2267);
nand U3480 (N_3480,N_2495,N_2578);
nand U3481 (N_3481,N_2368,N_2532);
nor U3482 (N_3482,N_2406,N_2999);
and U3483 (N_3483,N_2850,N_2172);
or U3484 (N_3484,N_2547,N_2444);
and U3485 (N_3485,N_2937,N_2627);
nand U3486 (N_3486,N_2738,N_2933);
nor U3487 (N_3487,N_2330,N_2290);
and U3488 (N_3488,N_2535,N_2557);
nor U3489 (N_3489,N_2580,N_2628);
nor U3490 (N_3490,N_2865,N_2309);
and U3491 (N_3491,N_2029,N_2604);
nor U3492 (N_3492,N_2530,N_2008);
and U3493 (N_3493,N_2710,N_2321);
nor U3494 (N_3494,N_2908,N_2987);
or U3495 (N_3495,N_2774,N_2112);
and U3496 (N_3496,N_2575,N_2922);
or U3497 (N_3497,N_2796,N_2018);
nor U3498 (N_3498,N_2402,N_2866);
or U3499 (N_3499,N_2314,N_2594);
and U3500 (N_3500,N_2193,N_2555);
nand U3501 (N_3501,N_2064,N_2009);
and U3502 (N_3502,N_2246,N_2975);
and U3503 (N_3503,N_2593,N_2651);
nand U3504 (N_3504,N_2918,N_2617);
and U3505 (N_3505,N_2491,N_2786);
or U3506 (N_3506,N_2864,N_2884);
nor U3507 (N_3507,N_2380,N_2948);
nand U3508 (N_3508,N_2741,N_2136);
or U3509 (N_3509,N_2134,N_2537);
and U3510 (N_3510,N_2656,N_2720);
nand U3511 (N_3511,N_2969,N_2835);
nor U3512 (N_3512,N_2276,N_2026);
nand U3513 (N_3513,N_2911,N_2317);
nor U3514 (N_3514,N_2000,N_2884);
nor U3515 (N_3515,N_2265,N_2679);
nand U3516 (N_3516,N_2782,N_2071);
and U3517 (N_3517,N_2456,N_2681);
and U3518 (N_3518,N_2568,N_2067);
or U3519 (N_3519,N_2714,N_2304);
or U3520 (N_3520,N_2716,N_2738);
or U3521 (N_3521,N_2254,N_2370);
nand U3522 (N_3522,N_2596,N_2850);
or U3523 (N_3523,N_2341,N_2407);
nand U3524 (N_3524,N_2335,N_2022);
or U3525 (N_3525,N_2149,N_2492);
nand U3526 (N_3526,N_2789,N_2523);
nand U3527 (N_3527,N_2461,N_2851);
nand U3528 (N_3528,N_2362,N_2696);
nand U3529 (N_3529,N_2491,N_2658);
and U3530 (N_3530,N_2295,N_2205);
nand U3531 (N_3531,N_2085,N_2061);
nand U3532 (N_3532,N_2315,N_2833);
or U3533 (N_3533,N_2153,N_2167);
nand U3534 (N_3534,N_2275,N_2813);
nor U3535 (N_3535,N_2555,N_2016);
nor U3536 (N_3536,N_2184,N_2808);
nand U3537 (N_3537,N_2441,N_2638);
nor U3538 (N_3538,N_2203,N_2239);
or U3539 (N_3539,N_2561,N_2911);
and U3540 (N_3540,N_2589,N_2203);
nand U3541 (N_3541,N_2485,N_2804);
nand U3542 (N_3542,N_2775,N_2498);
or U3543 (N_3543,N_2495,N_2029);
or U3544 (N_3544,N_2694,N_2162);
nand U3545 (N_3545,N_2726,N_2098);
and U3546 (N_3546,N_2280,N_2721);
nand U3547 (N_3547,N_2332,N_2011);
nand U3548 (N_3548,N_2186,N_2061);
nor U3549 (N_3549,N_2409,N_2223);
and U3550 (N_3550,N_2034,N_2796);
nand U3551 (N_3551,N_2303,N_2077);
and U3552 (N_3552,N_2925,N_2068);
and U3553 (N_3553,N_2234,N_2221);
or U3554 (N_3554,N_2207,N_2124);
nand U3555 (N_3555,N_2283,N_2431);
or U3556 (N_3556,N_2046,N_2567);
nor U3557 (N_3557,N_2576,N_2287);
and U3558 (N_3558,N_2286,N_2912);
nand U3559 (N_3559,N_2136,N_2592);
and U3560 (N_3560,N_2813,N_2508);
nand U3561 (N_3561,N_2168,N_2051);
or U3562 (N_3562,N_2833,N_2736);
nand U3563 (N_3563,N_2304,N_2770);
and U3564 (N_3564,N_2725,N_2124);
nor U3565 (N_3565,N_2542,N_2715);
or U3566 (N_3566,N_2525,N_2481);
and U3567 (N_3567,N_2960,N_2273);
nand U3568 (N_3568,N_2299,N_2860);
and U3569 (N_3569,N_2336,N_2968);
and U3570 (N_3570,N_2506,N_2097);
nand U3571 (N_3571,N_2623,N_2776);
or U3572 (N_3572,N_2736,N_2485);
nand U3573 (N_3573,N_2703,N_2555);
nor U3574 (N_3574,N_2097,N_2836);
nor U3575 (N_3575,N_2101,N_2258);
or U3576 (N_3576,N_2872,N_2812);
or U3577 (N_3577,N_2267,N_2256);
nor U3578 (N_3578,N_2396,N_2847);
nand U3579 (N_3579,N_2167,N_2178);
nor U3580 (N_3580,N_2015,N_2525);
and U3581 (N_3581,N_2365,N_2703);
nand U3582 (N_3582,N_2772,N_2724);
nor U3583 (N_3583,N_2836,N_2104);
or U3584 (N_3584,N_2382,N_2373);
nor U3585 (N_3585,N_2303,N_2446);
and U3586 (N_3586,N_2434,N_2429);
nand U3587 (N_3587,N_2174,N_2431);
and U3588 (N_3588,N_2774,N_2927);
or U3589 (N_3589,N_2744,N_2226);
nand U3590 (N_3590,N_2202,N_2209);
and U3591 (N_3591,N_2935,N_2838);
nor U3592 (N_3592,N_2292,N_2544);
or U3593 (N_3593,N_2281,N_2693);
nor U3594 (N_3594,N_2741,N_2355);
nor U3595 (N_3595,N_2359,N_2242);
or U3596 (N_3596,N_2220,N_2145);
and U3597 (N_3597,N_2170,N_2630);
or U3598 (N_3598,N_2429,N_2121);
or U3599 (N_3599,N_2030,N_2340);
nor U3600 (N_3600,N_2791,N_2434);
nor U3601 (N_3601,N_2045,N_2253);
nand U3602 (N_3602,N_2432,N_2452);
nand U3603 (N_3603,N_2022,N_2259);
and U3604 (N_3604,N_2248,N_2570);
and U3605 (N_3605,N_2034,N_2423);
or U3606 (N_3606,N_2042,N_2456);
nand U3607 (N_3607,N_2540,N_2662);
nand U3608 (N_3608,N_2163,N_2678);
nand U3609 (N_3609,N_2705,N_2718);
nor U3610 (N_3610,N_2854,N_2761);
nor U3611 (N_3611,N_2370,N_2447);
nand U3612 (N_3612,N_2892,N_2291);
nor U3613 (N_3613,N_2944,N_2098);
and U3614 (N_3614,N_2737,N_2732);
and U3615 (N_3615,N_2605,N_2460);
nand U3616 (N_3616,N_2641,N_2957);
and U3617 (N_3617,N_2444,N_2910);
and U3618 (N_3618,N_2425,N_2244);
xor U3619 (N_3619,N_2590,N_2331);
or U3620 (N_3620,N_2772,N_2272);
nand U3621 (N_3621,N_2310,N_2530);
and U3622 (N_3622,N_2839,N_2075);
nand U3623 (N_3623,N_2272,N_2664);
nand U3624 (N_3624,N_2985,N_2293);
nor U3625 (N_3625,N_2796,N_2478);
nand U3626 (N_3626,N_2790,N_2261);
or U3627 (N_3627,N_2128,N_2900);
nand U3628 (N_3628,N_2854,N_2973);
nor U3629 (N_3629,N_2659,N_2726);
and U3630 (N_3630,N_2322,N_2885);
nor U3631 (N_3631,N_2307,N_2285);
nand U3632 (N_3632,N_2445,N_2468);
nand U3633 (N_3633,N_2354,N_2030);
nand U3634 (N_3634,N_2117,N_2552);
nand U3635 (N_3635,N_2220,N_2639);
and U3636 (N_3636,N_2058,N_2484);
or U3637 (N_3637,N_2818,N_2348);
and U3638 (N_3638,N_2262,N_2392);
nand U3639 (N_3639,N_2745,N_2995);
and U3640 (N_3640,N_2022,N_2905);
nor U3641 (N_3641,N_2829,N_2118);
and U3642 (N_3642,N_2796,N_2167);
nor U3643 (N_3643,N_2683,N_2054);
nand U3644 (N_3644,N_2741,N_2501);
or U3645 (N_3645,N_2909,N_2364);
nand U3646 (N_3646,N_2772,N_2827);
and U3647 (N_3647,N_2423,N_2644);
and U3648 (N_3648,N_2384,N_2685);
and U3649 (N_3649,N_2548,N_2862);
or U3650 (N_3650,N_2355,N_2930);
or U3651 (N_3651,N_2141,N_2944);
and U3652 (N_3652,N_2139,N_2017);
nand U3653 (N_3653,N_2670,N_2488);
nand U3654 (N_3654,N_2128,N_2104);
or U3655 (N_3655,N_2346,N_2114);
nor U3656 (N_3656,N_2255,N_2514);
and U3657 (N_3657,N_2713,N_2111);
and U3658 (N_3658,N_2157,N_2893);
nand U3659 (N_3659,N_2814,N_2599);
and U3660 (N_3660,N_2581,N_2932);
or U3661 (N_3661,N_2759,N_2185);
nand U3662 (N_3662,N_2381,N_2149);
nor U3663 (N_3663,N_2944,N_2303);
and U3664 (N_3664,N_2526,N_2750);
nor U3665 (N_3665,N_2513,N_2682);
or U3666 (N_3666,N_2586,N_2616);
nand U3667 (N_3667,N_2272,N_2086);
or U3668 (N_3668,N_2634,N_2258);
nand U3669 (N_3669,N_2605,N_2441);
nand U3670 (N_3670,N_2739,N_2026);
nand U3671 (N_3671,N_2588,N_2807);
nor U3672 (N_3672,N_2249,N_2012);
nand U3673 (N_3673,N_2296,N_2776);
and U3674 (N_3674,N_2800,N_2958);
nor U3675 (N_3675,N_2514,N_2623);
nand U3676 (N_3676,N_2854,N_2965);
or U3677 (N_3677,N_2351,N_2992);
and U3678 (N_3678,N_2382,N_2677);
or U3679 (N_3679,N_2737,N_2864);
nor U3680 (N_3680,N_2499,N_2988);
or U3681 (N_3681,N_2047,N_2601);
nand U3682 (N_3682,N_2117,N_2847);
nand U3683 (N_3683,N_2901,N_2486);
or U3684 (N_3684,N_2868,N_2752);
nor U3685 (N_3685,N_2759,N_2188);
nand U3686 (N_3686,N_2822,N_2251);
nor U3687 (N_3687,N_2229,N_2791);
nor U3688 (N_3688,N_2010,N_2327);
and U3689 (N_3689,N_2716,N_2938);
nor U3690 (N_3690,N_2599,N_2649);
nor U3691 (N_3691,N_2704,N_2958);
nor U3692 (N_3692,N_2605,N_2380);
and U3693 (N_3693,N_2146,N_2883);
or U3694 (N_3694,N_2178,N_2142);
and U3695 (N_3695,N_2562,N_2960);
and U3696 (N_3696,N_2947,N_2640);
or U3697 (N_3697,N_2084,N_2280);
or U3698 (N_3698,N_2362,N_2442);
nor U3699 (N_3699,N_2129,N_2245);
nand U3700 (N_3700,N_2669,N_2612);
and U3701 (N_3701,N_2418,N_2495);
nor U3702 (N_3702,N_2774,N_2641);
nand U3703 (N_3703,N_2573,N_2829);
nand U3704 (N_3704,N_2174,N_2049);
nor U3705 (N_3705,N_2376,N_2824);
nand U3706 (N_3706,N_2612,N_2210);
nand U3707 (N_3707,N_2756,N_2537);
nand U3708 (N_3708,N_2228,N_2426);
and U3709 (N_3709,N_2520,N_2335);
nor U3710 (N_3710,N_2550,N_2547);
or U3711 (N_3711,N_2903,N_2213);
and U3712 (N_3712,N_2082,N_2946);
or U3713 (N_3713,N_2516,N_2072);
xor U3714 (N_3714,N_2438,N_2068);
and U3715 (N_3715,N_2032,N_2586);
nand U3716 (N_3716,N_2350,N_2819);
nand U3717 (N_3717,N_2015,N_2001);
or U3718 (N_3718,N_2704,N_2018);
or U3719 (N_3719,N_2148,N_2927);
nand U3720 (N_3720,N_2180,N_2615);
nand U3721 (N_3721,N_2453,N_2308);
or U3722 (N_3722,N_2551,N_2407);
nor U3723 (N_3723,N_2803,N_2870);
and U3724 (N_3724,N_2990,N_2462);
nor U3725 (N_3725,N_2316,N_2731);
nand U3726 (N_3726,N_2604,N_2833);
and U3727 (N_3727,N_2277,N_2524);
nand U3728 (N_3728,N_2746,N_2708);
nor U3729 (N_3729,N_2512,N_2571);
xnor U3730 (N_3730,N_2661,N_2480);
and U3731 (N_3731,N_2051,N_2303);
and U3732 (N_3732,N_2685,N_2260);
nand U3733 (N_3733,N_2973,N_2828);
or U3734 (N_3734,N_2932,N_2858);
or U3735 (N_3735,N_2272,N_2173);
and U3736 (N_3736,N_2121,N_2143);
nand U3737 (N_3737,N_2045,N_2867);
nand U3738 (N_3738,N_2081,N_2069);
or U3739 (N_3739,N_2770,N_2608);
nor U3740 (N_3740,N_2184,N_2420);
nand U3741 (N_3741,N_2928,N_2456);
or U3742 (N_3742,N_2014,N_2144);
nand U3743 (N_3743,N_2823,N_2086);
nor U3744 (N_3744,N_2581,N_2595);
and U3745 (N_3745,N_2149,N_2389);
nand U3746 (N_3746,N_2742,N_2415);
nor U3747 (N_3747,N_2007,N_2774);
nand U3748 (N_3748,N_2358,N_2697);
and U3749 (N_3749,N_2555,N_2834);
or U3750 (N_3750,N_2032,N_2033);
and U3751 (N_3751,N_2482,N_2632);
or U3752 (N_3752,N_2998,N_2037);
or U3753 (N_3753,N_2458,N_2376);
or U3754 (N_3754,N_2449,N_2635);
nand U3755 (N_3755,N_2559,N_2426);
nand U3756 (N_3756,N_2264,N_2490);
nor U3757 (N_3757,N_2107,N_2840);
nor U3758 (N_3758,N_2772,N_2395);
nor U3759 (N_3759,N_2958,N_2643);
and U3760 (N_3760,N_2108,N_2387);
or U3761 (N_3761,N_2079,N_2788);
nor U3762 (N_3762,N_2199,N_2187);
and U3763 (N_3763,N_2423,N_2047);
nor U3764 (N_3764,N_2207,N_2843);
or U3765 (N_3765,N_2365,N_2244);
or U3766 (N_3766,N_2362,N_2789);
and U3767 (N_3767,N_2679,N_2517);
or U3768 (N_3768,N_2170,N_2738);
nand U3769 (N_3769,N_2409,N_2160);
and U3770 (N_3770,N_2328,N_2894);
and U3771 (N_3771,N_2355,N_2268);
nand U3772 (N_3772,N_2634,N_2330);
or U3773 (N_3773,N_2148,N_2030);
xnor U3774 (N_3774,N_2518,N_2294);
nand U3775 (N_3775,N_2070,N_2416);
nand U3776 (N_3776,N_2386,N_2129);
and U3777 (N_3777,N_2798,N_2506);
and U3778 (N_3778,N_2388,N_2617);
or U3779 (N_3779,N_2566,N_2696);
or U3780 (N_3780,N_2864,N_2722);
and U3781 (N_3781,N_2471,N_2165);
nor U3782 (N_3782,N_2686,N_2912);
nor U3783 (N_3783,N_2168,N_2016);
nor U3784 (N_3784,N_2686,N_2909);
or U3785 (N_3785,N_2385,N_2773);
nand U3786 (N_3786,N_2912,N_2565);
nor U3787 (N_3787,N_2045,N_2802);
nand U3788 (N_3788,N_2103,N_2567);
nor U3789 (N_3789,N_2828,N_2340);
and U3790 (N_3790,N_2129,N_2830);
nor U3791 (N_3791,N_2540,N_2584);
xor U3792 (N_3792,N_2017,N_2325);
and U3793 (N_3793,N_2573,N_2831);
nor U3794 (N_3794,N_2906,N_2282);
and U3795 (N_3795,N_2337,N_2833);
nand U3796 (N_3796,N_2122,N_2601);
or U3797 (N_3797,N_2799,N_2430);
nand U3798 (N_3798,N_2945,N_2734);
or U3799 (N_3799,N_2212,N_2751);
nor U3800 (N_3800,N_2274,N_2375);
or U3801 (N_3801,N_2628,N_2214);
or U3802 (N_3802,N_2738,N_2753);
and U3803 (N_3803,N_2385,N_2406);
nand U3804 (N_3804,N_2296,N_2589);
and U3805 (N_3805,N_2371,N_2622);
or U3806 (N_3806,N_2215,N_2643);
nand U3807 (N_3807,N_2468,N_2541);
and U3808 (N_3808,N_2014,N_2226);
nand U3809 (N_3809,N_2302,N_2944);
nor U3810 (N_3810,N_2156,N_2017);
and U3811 (N_3811,N_2698,N_2690);
nand U3812 (N_3812,N_2046,N_2683);
and U3813 (N_3813,N_2757,N_2745);
nand U3814 (N_3814,N_2066,N_2547);
or U3815 (N_3815,N_2333,N_2727);
nor U3816 (N_3816,N_2999,N_2983);
nor U3817 (N_3817,N_2162,N_2921);
nand U3818 (N_3818,N_2671,N_2962);
and U3819 (N_3819,N_2023,N_2862);
nor U3820 (N_3820,N_2541,N_2122);
nor U3821 (N_3821,N_2836,N_2791);
nor U3822 (N_3822,N_2089,N_2245);
and U3823 (N_3823,N_2243,N_2931);
and U3824 (N_3824,N_2640,N_2296);
nand U3825 (N_3825,N_2635,N_2216);
nor U3826 (N_3826,N_2483,N_2773);
nand U3827 (N_3827,N_2602,N_2283);
nand U3828 (N_3828,N_2512,N_2412);
and U3829 (N_3829,N_2412,N_2679);
nor U3830 (N_3830,N_2462,N_2439);
nand U3831 (N_3831,N_2723,N_2867);
xor U3832 (N_3832,N_2418,N_2658);
and U3833 (N_3833,N_2797,N_2320);
nor U3834 (N_3834,N_2519,N_2675);
nand U3835 (N_3835,N_2615,N_2590);
and U3836 (N_3836,N_2785,N_2574);
nor U3837 (N_3837,N_2523,N_2070);
nand U3838 (N_3838,N_2541,N_2720);
and U3839 (N_3839,N_2361,N_2500);
or U3840 (N_3840,N_2568,N_2056);
or U3841 (N_3841,N_2973,N_2392);
and U3842 (N_3842,N_2979,N_2950);
nand U3843 (N_3843,N_2231,N_2307);
nor U3844 (N_3844,N_2540,N_2929);
nor U3845 (N_3845,N_2480,N_2921);
nand U3846 (N_3846,N_2075,N_2504);
or U3847 (N_3847,N_2379,N_2214);
and U3848 (N_3848,N_2214,N_2206);
and U3849 (N_3849,N_2871,N_2352);
and U3850 (N_3850,N_2640,N_2492);
or U3851 (N_3851,N_2825,N_2906);
nor U3852 (N_3852,N_2818,N_2702);
nand U3853 (N_3853,N_2160,N_2423);
or U3854 (N_3854,N_2422,N_2748);
or U3855 (N_3855,N_2761,N_2568);
nor U3856 (N_3856,N_2584,N_2115);
and U3857 (N_3857,N_2600,N_2061);
or U3858 (N_3858,N_2898,N_2367);
or U3859 (N_3859,N_2258,N_2046);
and U3860 (N_3860,N_2040,N_2260);
nor U3861 (N_3861,N_2565,N_2849);
xor U3862 (N_3862,N_2520,N_2891);
nand U3863 (N_3863,N_2978,N_2461);
nand U3864 (N_3864,N_2877,N_2935);
nand U3865 (N_3865,N_2586,N_2937);
and U3866 (N_3866,N_2702,N_2489);
and U3867 (N_3867,N_2679,N_2472);
or U3868 (N_3868,N_2700,N_2544);
nand U3869 (N_3869,N_2021,N_2228);
or U3870 (N_3870,N_2188,N_2060);
or U3871 (N_3871,N_2914,N_2594);
nand U3872 (N_3872,N_2010,N_2231);
nand U3873 (N_3873,N_2848,N_2539);
and U3874 (N_3874,N_2231,N_2079);
nand U3875 (N_3875,N_2221,N_2718);
nand U3876 (N_3876,N_2443,N_2649);
nand U3877 (N_3877,N_2162,N_2996);
and U3878 (N_3878,N_2060,N_2627);
or U3879 (N_3879,N_2493,N_2762);
nand U3880 (N_3880,N_2325,N_2232);
and U3881 (N_3881,N_2560,N_2684);
or U3882 (N_3882,N_2037,N_2472);
or U3883 (N_3883,N_2388,N_2819);
and U3884 (N_3884,N_2719,N_2698);
and U3885 (N_3885,N_2682,N_2621);
nand U3886 (N_3886,N_2282,N_2985);
nor U3887 (N_3887,N_2335,N_2222);
or U3888 (N_3888,N_2313,N_2868);
and U3889 (N_3889,N_2278,N_2450);
and U3890 (N_3890,N_2697,N_2040);
nor U3891 (N_3891,N_2123,N_2895);
or U3892 (N_3892,N_2248,N_2834);
and U3893 (N_3893,N_2820,N_2635);
nand U3894 (N_3894,N_2483,N_2910);
or U3895 (N_3895,N_2895,N_2793);
nor U3896 (N_3896,N_2732,N_2538);
or U3897 (N_3897,N_2804,N_2801);
nor U3898 (N_3898,N_2983,N_2576);
or U3899 (N_3899,N_2383,N_2648);
nand U3900 (N_3900,N_2808,N_2210);
nor U3901 (N_3901,N_2997,N_2819);
nand U3902 (N_3902,N_2490,N_2858);
xnor U3903 (N_3903,N_2401,N_2697);
nand U3904 (N_3904,N_2517,N_2257);
nor U3905 (N_3905,N_2540,N_2243);
and U3906 (N_3906,N_2725,N_2601);
nor U3907 (N_3907,N_2234,N_2471);
nor U3908 (N_3908,N_2134,N_2269);
nand U3909 (N_3909,N_2290,N_2790);
nor U3910 (N_3910,N_2329,N_2536);
and U3911 (N_3911,N_2335,N_2803);
nor U3912 (N_3912,N_2474,N_2465);
and U3913 (N_3913,N_2932,N_2077);
nor U3914 (N_3914,N_2175,N_2661);
nand U3915 (N_3915,N_2360,N_2980);
nand U3916 (N_3916,N_2730,N_2456);
or U3917 (N_3917,N_2748,N_2278);
or U3918 (N_3918,N_2132,N_2260);
and U3919 (N_3919,N_2989,N_2802);
or U3920 (N_3920,N_2436,N_2891);
and U3921 (N_3921,N_2807,N_2328);
or U3922 (N_3922,N_2227,N_2191);
or U3923 (N_3923,N_2964,N_2391);
nand U3924 (N_3924,N_2997,N_2535);
or U3925 (N_3925,N_2443,N_2109);
nor U3926 (N_3926,N_2477,N_2451);
nor U3927 (N_3927,N_2454,N_2305);
nor U3928 (N_3928,N_2564,N_2416);
nand U3929 (N_3929,N_2138,N_2996);
nand U3930 (N_3930,N_2044,N_2608);
and U3931 (N_3931,N_2687,N_2072);
or U3932 (N_3932,N_2454,N_2229);
or U3933 (N_3933,N_2374,N_2039);
and U3934 (N_3934,N_2951,N_2062);
and U3935 (N_3935,N_2765,N_2546);
or U3936 (N_3936,N_2443,N_2856);
nand U3937 (N_3937,N_2297,N_2837);
nor U3938 (N_3938,N_2058,N_2500);
and U3939 (N_3939,N_2341,N_2173);
or U3940 (N_3940,N_2401,N_2320);
or U3941 (N_3941,N_2217,N_2303);
or U3942 (N_3942,N_2905,N_2635);
or U3943 (N_3943,N_2354,N_2678);
and U3944 (N_3944,N_2710,N_2580);
or U3945 (N_3945,N_2306,N_2182);
xor U3946 (N_3946,N_2894,N_2259);
nor U3947 (N_3947,N_2273,N_2596);
and U3948 (N_3948,N_2141,N_2602);
and U3949 (N_3949,N_2391,N_2348);
and U3950 (N_3950,N_2983,N_2628);
nor U3951 (N_3951,N_2443,N_2943);
nand U3952 (N_3952,N_2896,N_2559);
nand U3953 (N_3953,N_2140,N_2916);
and U3954 (N_3954,N_2942,N_2882);
nor U3955 (N_3955,N_2132,N_2339);
nor U3956 (N_3956,N_2547,N_2875);
or U3957 (N_3957,N_2783,N_2622);
or U3958 (N_3958,N_2466,N_2000);
and U3959 (N_3959,N_2606,N_2976);
nand U3960 (N_3960,N_2339,N_2332);
nor U3961 (N_3961,N_2812,N_2021);
nor U3962 (N_3962,N_2568,N_2336);
or U3963 (N_3963,N_2760,N_2287);
or U3964 (N_3964,N_2995,N_2015);
xor U3965 (N_3965,N_2608,N_2397);
and U3966 (N_3966,N_2651,N_2266);
nor U3967 (N_3967,N_2502,N_2001);
or U3968 (N_3968,N_2850,N_2474);
nand U3969 (N_3969,N_2005,N_2074);
nor U3970 (N_3970,N_2915,N_2350);
nand U3971 (N_3971,N_2486,N_2462);
and U3972 (N_3972,N_2603,N_2509);
nand U3973 (N_3973,N_2030,N_2304);
nor U3974 (N_3974,N_2786,N_2835);
nand U3975 (N_3975,N_2090,N_2599);
nor U3976 (N_3976,N_2661,N_2963);
or U3977 (N_3977,N_2634,N_2837);
and U3978 (N_3978,N_2823,N_2214);
nor U3979 (N_3979,N_2345,N_2152);
or U3980 (N_3980,N_2189,N_2551);
and U3981 (N_3981,N_2582,N_2862);
nand U3982 (N_3982,N_2289,N_2116);
or U3983 (N_3983,N_2577,N_2686);
and U3984 (N_3984,N_2256,N_2974);
nand U3985 (N_3985,N_2893,N_2510);
and U3986 (N_3986,N_2874,N_2273);
nand U3987 (N_3987,N_2232,N_2869);
or U3988 (N_3988,N_2979,N_2074);
nor U3989 (N_3989,N_2756,N_2430);
nor U3990 (N_3990,N_2808,N_2049);
or U3991 (N_3991,N_2365,N_2228);
or U3992 (N_3992,N_2669,N_2005);
nor U3993 (N_3993,N_2255,N_2165);
nand U3994 (N_3994,N_2893,N_2365);
nor U3995 (N_3995,N_2827,N_2843);
or U3996 (N_3996,N_2280,N_2668);
nor U3997 (N_3997,N_2827,N_2894);
and U3998 (N_3998,N_2288,N_2981);
or U3999 (N_3999,N_2451,N_2755);
or U4000 (N_4000,N_3418,N_3100);
nand U4001 (N_4001,N_3490,N_3306);
or U4002 (N_4002,N_3785,N_3009);
nor U4003 (N_4003,N_3104,N_3386);
nor U4004 (N_4004,N_3141,N_3071);
nand U4005 (N_4005,N_3112,N_3154);
nand U4006 (N_4006,N_3321,N_3970);
or U4007 (N_4007,N_3671,N_3819);
nand U4008 (N_4008,N_3413,N_3797);
nor U4009 (N_4009,N_3642,N_3768);
nor U4010 (N_4010,N_3981,N_3274);
or U4011 (N_4011,N_3007,N_3194);
or U4012 (N_4012,N_3215,N_3103);
or U4013 (N_4013,N_3001,N_3500);
or U4014 (N_4014,N_3199,N_3551);
nor U4015 (N_4015,N_3209,N_3412);
or U4016 (N_4016,N_3822,N_3808);
nor U4017 (N_4017,N_3210,N_3099);
nor U4018 (N_4018,N_3085,N_3213);
and U4019 (N_4019,N_3143,N_3656);
nand U4020 (N_4020,N_3515,N_3392);
and U4021 (N_4021,N_3157,N_3381);
and U4022 (N_4022,N_3982,N_3180);
or U4023 (N_4023,N_3409,N_3844);
and U4024 (N_4024,N_3593,N_3816);
nor U4025 (N_4025,N_3063,N_3929);
nor U4026 (N_4026,N_3297,N_3932);
nor U4027 (N_4027,N_3953,N_3246);
nor U4028 (N_4028,N_3097,N_3153);
nor U4029 (N_4029,N_3528,N_3996);
or U4030 (N_4030,N_3400,N_3331);
or U4031 (N_4031,N_3193,N_3526);
nor U4032 (N_4032,N_3948,N_3156);
or U4033 (N_4033,N_3757,N_3689);
nor U4034 (N_4034,N_3842,N_3573);
and U4035 (N_4035,N_3545,N_3602);
nand U4036 (N_4036,N_3655,N_3339);
nand U4037 (N_4037,N_3232,N_3544);
nand U4038 (N_4038,N_3423,N_3444);
nor U4039 (N_4039,N_3295,N_3968);
nor U4040 (N_4040,N_3479,N_3938);
and U4041 (N_4041,N_3991,N_3442);
nor U4042 (N_4042,N_3150,N_3491);
nand U4043 (N_4043,N_3342,N_3627);
nand U4044 (N_4044,N_3315,N_3145);
nand U4045 (N_4045,N_3108,N_3709);
or U4046 (N_4046,N_3497,N_3975);
and U4047 (N_4047,N_3841,N_3292);
or U4048 (N_4048,N_3588,N_3184);
or U4049 (N_4049,N_3231,N_3512);
nand U4050 (N_4050,N_3595,N_3269);
nand U4051 (N_4051,N_3467,N_3674);
nor U4052 (N_4052,N_3114,N_3237);
nand U4053 (N_4053,N_3893,N_3020);
and U4054 (N_4054,N_3823,N_3238);
or U4055 (N_4055,N_3169,N_3926);
and U4056 (N_4056,N_3662,N_3185);
or U4057 (N_4057,N_3802,N_3972);
or U4058 (N_4058,N_3736,N_3234);
xor U4059 (N_4059,N_3459,N_3728);
nor U4060 (N_4060,N_3755,N_3658);
nand U4061 (N_4061,N_3590,N_3850);
or U4062 (N_4062,N_3620,N_3189);
nor U4063 (N_4063,N_3918,N_3920);
nor U4064 (N_4064,N_3033,N_3688);
and U4065 (N_4065,N_3142,N_3317);
and U4066 (N_4066,N_3079,N_3705);
nand U4067 (N_4067,N_3075,N_3503);
nor U4068 (N_4068,N_3446,N_3690);
and U4069 (N_4069,N_3307,N_3628);
nand U4070 (N_4070,N_3597,N_3319);
nor U4071 (N_4071,N_3687,N_3083);
nand U4072 (N_4072,N_3577,N_3041);
nand U4073 (N_4073,N_3566,N_3228);
nor U4074 (N_4074,N_3300,N_3366);
nor U4075 (N_4075,N_3496,N_3152);
nor U4076 (N_4076,N_3048,N_3149);
nor U4077 (N_4077,N_3259,N_3026);
nor U4078 (N_4078,N_3477,N_3725);
nor U4079 (N_4079,N_3264,N_3860);
and U4080 (N_4080,N_3128,N_3188);
nor U4081 (N_4081,N_3879,N_3046);
nand U4082 (N_4082,N_3651,N_3166);
or U4083 (N_4083,N_3583,N_3520);
nand U4084 (N_4084,N_3610,N_3028);
nor U4085 (N_4085,N_3135,N_3223);
and U4086 (N_4086,N_3378,N_3691);
or U4087 (N_4087,N_3022,N_3700);
nand U4088 (N_4088,N_3469,N_3622);
nor U4089 (N_4089,N_3021,N_3482);
or U4090 (N_4090,N_3277,N_3778);
nor U4091 (N_4091,N_3758,N_3186);
or U4092 (N_4092,N_3943,N_3115);
nand U4093 (N_4093,N_3456,N_3582);
and U4094 (N_4094,N_3127,N_3834);
and U4095 (N_4095,N_3208,N_3639);
or U4096 (N_4096,N_3624,N_3694);
or U4097 (N_4097,N_3084,N_3043);
nor U4098 (N_4098,N_3276,N_3570);
nor U4099 (N_4099,N_3887,N_3296);
nand U4100 (N_4100,N_3502,N_3096);
and U4101 (N_4101,N_3164,N_3343);
nor U4102 (N_4102,N_3712,N_3181);
and U4103 (N_4103,N_3645,N_3334);
or U4104 (N_4104,N_3915,N_3191);
or U4105 (N_4105,N_3762,N_3042);
and U4106 (N_4106,N_3977,N_3513);
and U4107 (N_4107,N_3522,N_3717);
or U4108 (N_4108,N_3966,N_3944);
and U4109 (N_4109,N_3441,N_3810);
nand U4110 (N_4110,N_3495,N_3748);
nand U4111 (N_4111,N_3037,N_3643);
nor U4112 (N_4112,N_3449,N_3554);
and U4113 (N_4113,N_3813,N_3427);
nand U4114 (N_4114,N_3793,N_3359);
or U4115 (N_4115,N_3062,N_3950);
nand U4116 (N_4116,N_3747,N_3068);
and U4117 (N_4117,N_3571,N_3167);
nor U4118 (N_4118,N_3455,N_3616);
nand U4119 (N_4119,N_3776,N_3775);
and U4120 (N_4120,N_3010,N_3777);
and U4121 (N_4121,N_3330,N_3473);
nor U4122 (N_4122,N_3971,N_3326);
nor U4123 (N_4123,N_3867,N_3067);
nor U4124 (N_4124,N_3931,N_3242);
nand U4125 (N_4125,N_3124,N_3325);
nand U4126 (N_4126,N_3634,N_3052);
nor U4127 (N_4127,N_3155,N_3871);
and U4128 (N_4128,N_3407,N_3572);
nor U4129 (N_4129,N_3290,N_3849);
nand U4130 (N_4130,N_3447,N_3175);
nand U4131 (N_4131,N_3692,N_3621);
and U4132 (N_4132,N_3241,N_3388);
nor U4133 (N_4133,N_3091,N_3752);
or U4134 (N_4134,N_3458,N_3675);
or U4135 (N_4135,N_3555,N_3744);
or U4136 (N_4136,N_3187,N_3465);
and U4137 (N_4137,N_3222,N_3078);
or U4138 (N_4138,N_3393,N_3680);
or U4139 (N_4139,N_3925,N_3422);
nor U4140 (N_4140,N_3303,N_3288);
and U4141 (N_4141,N_3013,N_3499);
or U4142 (N_4142,N_3909,N_3106);
nand U4143 (N_4143,N_3924,N_3698);
nand U4144 (N_4144,N_3756,N_3023);
or U4145 (N_4145,N_3450,N_3608);
and U4146 (N_4146,N_3333,N_3677);
nand U4147 (N_4147,N_3148,N_3707);
or U4148 (N_4148,N_3815,N_3769);
nor U4149 (N_4149,N_3786,N_3270);
and U4150 (N_4150,N_3864,N_3137);
nor U4151 (N_4151,N_3875,N_3019);
nand U4152 (N_4152,N_3481,N_3484);
or U4153 (N_4153,N_3192,N_3764);
nand U4154 (N_4154,N_3840,N_3685);
nand U4155 (N_4155,N_3733,N_3064);
or U4156 (N_4156,N_3601,N_3575);
nor U4157 (N_4157,N_3569,N_3561);
nand U4158 (N_4158,N_3701,N_3695);
or U4159 (N_4159,N_3094,N_3890);
nor U4160 (N_4160,N_3506,N_3082);
nor U4161 (N_4161,N_3789,N_3548);
nor U4162 (N_4162,N_3603,N_3576);
and U4163 (N_4163,N_3804,N_3941);
nand U4164 (N_4164,N_3719,N_3611);
nand U4165 (N_4165,N_3088,N_3221);
nor U4166 (N_4166,N_3913,N_3792);
or U4167 (N_4167,N_3781,N_3766);
nand U4168 (N_4168,N_3293,N_3371);
nand U4169 (N_4169,N_3002,N_3947);
or U4170 (N_4170,N_3439,N_3424);
nand U4171 (N_4171,N_3735,N_3868);
and U4172 (N_4172,N_3126,N_3814);
nand U4173 (N_4173,N_3908,N_3396);
nor U4174 (N_4174,N_3825,N_3251);
nand U4175 (N_4175,N_3087,N_3606);
nand U4176 (N_4176,N_3648,N_3183);
nor U4177 (N_4177,N_3335,N_3179);
nor U4178 (N_4178,N_3653,N_3962);
nor U4179 (N_4179,N_3217,N_3759);
or U4180 (N_4180,N_3765,N_3865);
nor U4181 (N_4181,N_3877,N_3345);
nand U4182 (N_4182,N_3811,N_3668);
nand U4183 (N_4183,N_3410,N_3726);
nor U4184 (N_4184,N_3745,N_3873);
nand U4185 (N_4185,N_3605,N_3767);
or U4186 (N_4186,N_3980,N_3483);
nor U4187 (N_4187,N_3951,N_3451);
or U4188 (N_4188,N_3942,N_3952);
or U4189 (N_4189,N_3957,N_3667);
and U4190 (N_4190,N_3669,N_3015);
and U4191 (N_4191,N_3612,N_3861);
nor U4192 (N_4192,N_3074,N_3433);
nor U4193 (N_4193,N_3809,N_3937);
or U4194 (N_4194,N_3579,N_3132);
or U4195 (N_4195,N_3696,N_3494);
nor U4196 (N_4196,N_3284,N_3742);
nor U4197 (N_4197,N_3090,N_3430);
or U4198 (N_4198,N_3262,N_3539);
nor U4199 (N_4199,N_3031,N_3111);
nor U4200 (N_4200,N_3580,N_3492);
nand U4201 (N_4201,N_3462,N_3406);
and U4202 (N_4202,N_3955,N_3660);
nand U4203 (N_4203,N_3626,N_3302);
nand U4204 (N_4204,N_3640,N_3732);
nor U4205 (N_4205,N_3344,N_3403);
or U4206 (N_4206,N_3714,N_3693);
nor U4207 (N_4207,N_3305,N_3738);
nor U4208 (N_4208,N_3934,N_3054);
nand U4209 (N_4209,N_3702,N_3049);
and U4210 (N_4210,N_3391,N_3699);
and U4211 (N_4211,N_3994,N_3939);
and U4212 (N_4212,N_3346,N_3516);
or U4213 (N_4213,N_3587,N_3471);
nand U4214 (N_4214,N_3637,N_3349);
or U4215 (N_4215,N_3165,N_3965);
nor U4216 (N_4216,N_3904,N_3383);
or U4217 (N_4217,N_3058,N_3435);
nor U4218 (N_4218,N_3652,N_3846);
or U4219 (N_4219,N_3843,N_3011);
and U4220 (N_4220,N_3585,N_3003);
nand U4221 (N_4221,N_3990,N_3235);
or U4222 (N_4222,N_3831,N_3623);
nor U4223 (N_4223,N_3927,N_3830);
and U4224 (N_4224,N_3255,N_3060);
nand U4225 (N_4225,N_3151,N_3959);
nand U4226 (N_4226,N_3059,N_3045);
nor U4227 (N_4227,N_3686,N_3273);
or U4228 (N_4228,N_3105,N_3564);
nand U4229 (N_4229,N_3379,N_3654);
nor U4230 (N_4230,N_3676,N_3487);
nor U4231 (N_4231,N_3529,N_3987);
nor U4232 (N_4232,N_3466,N_3380);
nor U4233 (N_4233,N_3604,N_3531);
nor U4234 (N_4234,N_3214,N_3443);
and U4235 (N_4235,N_3684,N_3140);
nor U4236 (N_4236,N_3558,N_3250);
nand U4237 (N_4237,N_3886,N_3282);
or U4238 (N_4238,N_3212,N_3835);
and U4239 (N_4239,N_3207,N_3314);
and U4240 (N_4240,N_3275,N_3417);
and U4241 (N_4241,N_3807,N_3229);
nor U4242 (N_4242,N_3710,N_3508);
nor U4243 (N_4243,N_3289,N_3369);
or U4244 (N_4244,N_3404,N_3069);
nor U4245 (N_4245,N_3395,N_3619);
nor U4246 (N_4246,N_3129,N_3357);
or U4247 (N_4247,N_3988,N_3517);
nand U4248 (N_4248,N_3800,N_3788);
or U4249 (N_4249,N_3532,N_3614);
xor U4250 (N_4250,N_3445,N_3928);
nor U4251 (N_4251,N_3704,N_3697);
nand U4252 (N_4252,N_3287,N_3113);
nand U4253 (N_4253,N_3859,N_3974);
nand U4254 (N_4254,N_3883,N_3631);
nand U4255 (N_4255,N_3102,N_3452);
nor U4256 (N_4256,N_3472,N_3552);
xor U4257 (N_4257,N_3741,N_3266);
and U4258 (N_4258,N_3826,N_3964);
nand U4259 (N_4259,N_3598,N_3795);
nand U4260 (N_4260,N_3901,N_3415);
or U4261 (N_4261,N_3363,N_3408);
nor U4262 (N_4262,N_3116,N_3190);
and U4263 (N_4263,N_3252,N_3592);
nand U4264 (N_4264,N_3428,N_3018);
or U4265 (N_4265,N_3464,N_3897);
nand U4266 (N_4266,N_3556,N_3527);
nand U4267 (N_4267,N_3382,N_3236);
nor U4268 (N_4268,N_3336,N_3182);
and U4269 (N_4269,N_3838,N_3540);
or U4270 (N_4270,N_3485,N_3905);
or U4271 (N_4271,N_3414,N_3322);
nor U4272 (N_4272,N_3387,N_3787);
and U4273 (N_4273,N_3425,N_3411);
and U4274 (N_4274,N_3420,N_3377);
and U4275 (N_4275,N_3254,N_3353);
and U4276 (N_4276,N_3374,N_3737);
nor U4277 (N_4277,N_3659,N_3978);
nor U4278 (N_4278,N_3881,N_3159);
nor U4279 (N_4279,N_3872,N_3541);
and U4280 (N_4280,N_3956,N_3286);
or U4281 (N_4281,N_3761,N_3912);
and U4282 (N_4282,N_3036,N_3311);
and U4283 (N_4283,N_3098,N_3607);
nor U4284 (N_4284,N_3711,N_3316);
or U4285 (N_4285,N_3895,N_3120);
nor U4286 (N_4286,N_3783,N_3770);
nor U4287 (N_4287,N_3914,N_3780);
or U4288 (N_4288,N_3081,N_3833);
xnor U4289 (N_4289,N_3727,N_3440);
or U4290 (N_4290,N_3664,N_3240);
and U4291 (N_4291,N_3313,N_3304);
or U4292 (N_4292,N_3954,N_3935);
or U4293 (N_4293,N_3878,N_3550);
or U4294 (N_4294,N_3205,N_3799);
and U4295 (N_4295,N_3900,N_3560);
nor U4296 (N_4296,N_3754,N_3853);
nor U4297 (N_4297,N_3239,N_3683);
nor U4298 (N_4298,N_3753,N_3794);
nor U4299 (N_4299,N_3751,N_3072);
nor U4300 (N_4300,N_3201,N_3646);
nor U4301 (N_4301,N_3076,N_3862);
or U4302 (N_4302,N_3848,N_3524);
nor U4303 (N_4303,N_3923,N_3244);
and U4304 (N_4304,N_3206,N_3347);
and U4305 (N_4305,N_3249,N_3874);
or U4306 (N_4306,N_3828,N_3945);
or U4307 (N_4307,N_3567,N_3749);
nand U4308 (N_4308,N_3613,N_3168);
and U4309 (N_4309,N_3734,N_3260);
nor U4310 (N_4310,N_3549,N_3352);
nand U4311 (N_4311,N_3869,N_3448);
and U4312 (N_4312,N_3958,N_3372);
nor U4313 (N_4313,N_3933,N_3461);
or U4314 (N_4314,N_3504,N_3257);
xor U4315 (N_4315,N_3723,N_3638);
xnor U4316 (N_4316,N_3801,N_3518);
nor U4317 (N_4317,N_3921,N_3044);
nor U4318 (N_4318,N_3636,N_3029);
or U4319 (N_4319,N_3258,N_3219);
and U4320 (N_4320,N_3581,N_3324);
nor U4321 (N_4321,N_3419,N_3092);
nor U4322 (N_4322,N_3973,N_3534);
nand U4323 (N_4323,N_3650,N_3498);
nand U4324 (N_4324,N_3227,N_3530);
nand U4325 (N_4325,N_3586,N_3715);
nor U4326 (N_4326,N_3855,N_3030);
or U4327 (N_4327,N_3509,N_3332);
nor U4328 (N_4328,N_3401,N_3438);
and U4329 (N_4329,N_3327,N_3599);
nor U4330 (N_4330,N_3421,N_3892);
or U4331 (N_4331,N_3117,N_3230);
and U4332 (N_4332,N_3278,N_3323);
xnor U4333 (N_4333,N_3782,N_3385);
and U4334 (N_4334,N_3040,N_3678);
nand U4335 (N_4335,N_3203,N_3746);
and U4336 (N_4336,N_3839,N_3673);
or U4337 (N_4337,N_3930,N_3337);
nor U4338 (N_4338,N_3301,N_3474);
nor U4339 (N_4339,N_3122,N_3995);
nor U4340 (N_4340,N_3008,N_3247);
or U4341 (N_4341,N_3220,N_3969);
or U4342 (N_4342,N_3774,N_3125);
or U4343 (N_4343,N_3121,N_3470);
nor U4344 (N_4344,N_3546,N_3589);
nand U4345 (N_4345,N_3004,N_3429);
or U4346 (N_4346,N_3310,N_3837);
nand U4347 (N_4347,N_3389,N_3489);
and U4348 (N_4348,N_3773,N_3635);
and U4349 (N_4349,N_3817,N_3594);
or U4350 (N_4350,N_3053,N_3625);
nand U4351 (N_4351,N_3703,N_3390);
nor U4352 (N_4352,N_3880,N_3158);
nand U4353 (N_4353,N_3478,N_3600);
nand U4354 (N_4354,N_3178,N_3827);
and U4355 (N_4355,N_3731,N_3641);
or U4356 (N_4356,N_3894,N_3961);
or U4357 (N_4357,N_3218,N_3967);
nor U4358 (N_4358,N_3110,N_3328);
and U4359 (N_4359,N_3261,N_3468);
nor U4360 (N_4360,N_3056,N_3364);
nand U4361 (N_4361,N_3146,N_3176);
or U4362 (N_4362,N_3398,N_3279);
nor U4363 (N_4363,N_3061,N_3657);
nor U4364 (N_4364,N_3716,N_3362);
nor U4365 (N_4365,N_3535,N_3501);
nand U4366 (N_4366,N_3463,N_3505);
nor U4367 (N_4367,N_3351,N_3888);
nand U4368 (N_4368,N_3682,N_3784);
nor U4369 (N_4369,N_3162,N_3596);
nand U4370 (N_4370,N_3163,N_3866);
and U4371 (N_4371,N_3457,N_3584);
or U4372 (N_4372,N_3373,N_3134);
nor U4373 (N_4373,N_3005,N_3565);
nor U4374 (N_4374,N_3976,N_3946);
or U4375 (N_4375,N_3453,N_3899);
nor U4376 (N_4376,N_3722,N_3298);
and U4377 (N_4377,N_3665,N_3666);
or U4378 (N_4378,N_3730,N_3476);
nor U4379 (N_4379,N_3245,N_3173);
or U4380 (N_4380,N_3820,N_3211);
nor U4381 (N_4381,N_3089,N_3216);
nand U4382 (N_4382,N_3025,N_3718);
nand U4383 (N_4383,N_3910,N_3233);
nor U4384 (N_4384,N_3488,N_3035);
or U4385 (N_4385,N_3320,N_3521);
nand U4386 (N_4386,N_3519,N_3174);
nand U4387 (N_4387,N_3633,N_3574);
nand U4388 (N_4388,N_3000,N_3243);
nand U4389 (N_4389,N_3055,N_3202);
or U4390 (N_4390,N_3559,N_3437);
nand U4391 (N_4391,N_3902,N_3032);
or U4392 (N_4392,N_3720,N_3291);
nand U4393 (N_4393,N_3992,N_3647);
or U4394 (N_4394,N_3891,N_3983);
and U4395 (N_4395,N_3708,N_3138);
nand U4396 (N_4396,N_3989,N_3204);
or U4397 (N_4397,N_3397,N_3779);
nor U4398 (N_4398,N_3960,N_3402);
nor U4399 (N_4399,N_3256,N_3514);
or U4400 (N_4400,N_3538,N_3365);
or U4401 (N_4401,N_3077,N_3012);
or U4402 (N_4402,N_3267,N_3917);
or U4403 (N_4403,N_3024,N_3014);
nor U4404 (N_4404,N_3940,N_3171);
and U4405 (N_4405,N_3985,N_3368);
nand U4406 (N_4406,N_3006,N_3361);
or U4407 (N_4407,N_3729,N_3663);
nor U4408 (N_4408,N_3681,N_3405);
and U4409 (N_4409,N_3805,N_3394);
and U4410 (N_4410,N_3760,N_3740);
nor U4411 (N_4411,N_3147,N_3568);
nand U4412 (N_4412,N_3537,N_3283);
nand U4413 (N_4413,N_3460,N_3309);
nor U4414 (N_4414,N_3889,N_3856);
or U4415 (N_4415,N_3318,N_3161);
and U4416 (N_4416,N_3824,N_3426);
and U4417 (N_4417,N_3454,N_3578);
nor U4418 (N_4418,N_3047,N_3341);
and U4419 (N_4419,N_3027,N_3851);
nor U4420 (N_4420,N_3272,N_3039);
and U4421 (N_4421,N_3118,N_3195);
nor U4422 (N_4422,N_3329,N_3870);
and U4423 (N_4423,N_3706,N_3818);
nand U4424 (N_4424,N_3858,N_3863);
and U4425 (N_4425,N_3493,N_3130);
nor U4426 (N_4426,N_3907,N_3644);
and U4427 (N_4427,N_3355,N_3070);
nand U4428 (N_4428,N_3997,N_3743);
nand U4429 (N_4429,N_3107,N_3198);
nor U4430 (N_4430,N_3119,N_3095);
or U4431 (N_4431,N_3172,N_3226);
and U4432 (N_4432,N_3821,N_3615);
and U4433 (N_4433,N_3144,N_3370);
and U4434 (N_4434,N_3949,N_3523);
nor U4435 (N_4435,N_3017,N_3525);
nor U4436 (N_4436,N_3016,N_3066);
nor U4437 (N_4437,N_3536,N_3050);
or U4438 (N_4438,N_3798,N_3312);
nand U4439 (N_4439,N_3280,N_3486);
nand U4440 (N_4440,N_3253,N_3763);
nor U4441 (N_4441,N_3547,N_3375);
and U4442 (N_4442,N_3771,N_3791);
nor U4443 (N_4443,N_3649,N_3903);
nand U4444 (N_4444,N_3562,N_3101);
or U4445 (N_4445,N_3739,N_3884);
nand U4446 (N_4446,N_3563,N_3533);
or U4447 (N_4447,N_3542,N_3832);
and U4448 (N_4448,N_3436,N_3922);
nor U4449 (N_4449,N_3271,N_3224);
and U4450 (N_4450,N_3896,N_3916);
and U4451 (N_4451,N_3845,N_3854);
and U4452 (N_4452,N_3750,N_3384);
or U4453 (N_4453,N_3200,N_3416);
or U4454 (N_4454,N_3553,N_3225);
and U4455 (N_4455,N_3609,N_3360);
nand U4456 (N_4456,N_3836,N_3963);
and U4457 (N_4457,N_3661,N_3618);
and U4458 (N_4458,N_3507,N_3340);
or U4459 (N_4459,N_3557,N_3591);
or U4460 (N_4460,N_3434,N_3984);
or U4461 (N_4461,N_3721,N_3812);
nor U4462 (N_4462,N_3263,N_3109);
or U4463 (N_4463,N_3057,N_3131);
nand U4464 (N_4464,N_3630,N_3265);
nor U4465 (N_4465,N_3160,N_3170);
and U4466 (N_4466,N_3086,N_3399);
nand U4467 (N_4467,N_3480,N_3617);
and U4468 (N_4468,N_3772,N_3358);
or U4469 (N_4469,N_3432,N_3898);
or U4470 (N_4470,N_3724,N_3294);
or U4471 (N_4471,N_3713,N_3367);
or U4472 (N_4472,N_3629,N_3034);
or U4473 (N_4473,N_3998,N_3281);
nand U4474 (N_4474,N_3073,N_3123);
or U4475 (N_4475,N_3876,N_3093);
nand U4476 (N_4476,N_3911,N_3510);
or U4477 (N_4477,N_3803,N_3356);
nor U4478 (N_4478,N_3196,N_3354);
nor U4479 (N_4479,N_3065,N_3350);
and U4480 (N_4480,N_3268,N_3885);
or U4481 (N_4481,N_3806,N_3919);
nor U4482 (N_4482,N_3882,N_3080);
or U4483 (N_4483,N_3986,N_3348);
or U4484 (N_4484,N_3285,N_3829);
and U4485 (N_4485,N_3847,N_3670);
nand U4486 (N_4486,N_3857,N_3248);
nor U4487 (N_4487,N_3177,N_3511);
nor U4488 (N_4488,N_3790,N_3999);
and U4489 (N_4489,N_3299,N_3308);
nand U4490 (N_4490,N_3936,N_3475);
and U4491 (N_4491,N_3672,N_3796);
or U4492 (N_4492,N_3543,N_3136);
nand U4493 (N_4493,N_3051,N_3979);
or U4494 (N_4494,N_3038,N_3852);
nand U4495 (N_4495,N_3338,N_3679);
and U4496 (N_4496,N_3133,N_3376);
nand U4497 (N_4497,N_3139,N_3632);
or U4498 (N_4498,N_3993,N_3431);
nand U4499 (N_4499,N_3197,N_3906);
or U4500 (N_4500,N_3614,N_3439);
nor U4501 (N_4501,N_3938,N_3567);
or U4502 (N_4502,N_3242,N_3158);
and U4503 (N_4503,N_3809,N_3612);
nand U4504 (N_4504,N_3619,N_3856);
nor U4505 (N_4505,N_3616,N_3990);
nand U4506 (N_4506,N_3272,N_3831);
nor U4507 (N_4507,N_3825,N_3142);
and U4508 (N_4508,N_3843,N_3495);
and U4509 (N_4509,N_3152,N_3131);
or U4510 (N_4510,N_3538,N_3179);
nand U4511 (N_4511,N_3688,N_3514);
and U4512 (N_4512,N_3980,N_3213);
nand U4513 (N_4513,N_3220,N_3398);
nor U4514 (N_4514,N_3173,N_3181);
nand U4515 (N_4515,N_3513,N_3354);
nor U4516 (N_4516,N_3261,N_3864);
or U4517 (N_4517,N_3739,N_3867);
nand U4518 (N_4518,N_3231,N_3800);
or U4519 (N_4519,N_3244,N_3720);
or U4520 (N_4520,N_3306,N_3514);
nand U4521 (N_4521,N_3456,N_3390);
and U4522 (N_4522,N_3477,N_3802);
nor U4523 (N_4523,N_3854,N_3597);
nand U4524 (N_4524,N_3560,N_3806);
nand U4525 (N_4525,N_3740,N_3037);
xnor U4526 (N_4526,N_3378,N_3043);
and U4527 (N_4527,N_3077,N_3104);
nand U4528 (N_4528,N_3340,N_3040);
nor U4529 (N_4529,N_3253,N_3681);
or U4530 (N_4530,N_3170,N_3381);
nor U4531 (N_4531,N_3661,N_3411);
or U4532 (N_4532,N_3508,N_3307);
nor U4533 (N_4533,N_3112,N_3805);
or U4534 (N_4534,N_3500,N_3247);
and U4535 (N_4535,N_3452,N_3449);
or U4536 (N_4536,N_3617,N_3767);
or U4537 (N_4537,N_3930,N_3743);
and U4538 (N_4538,N_3438,N_3293);
or U4539 (N_4539,N_3831,N_3652);
or U4540 (N_4540,N_3660,N_3374);
nand U4541 (N_4541,N_3219,N_3505);
nand U4542 (N_4542,N_3581,N_3462);
and U4543 (N_4543,N_3318,N_3064);
and U4544 (N_4544,N_3743,N_3966);
and U4545 (N_4545,N_3705,N_3757);
nand U4546 (N_4546,N_3435,N_3127);
nand U4547 (N_4547,N_3504,N_3842);
or U4548 (N_4548,N_3514,N_3196);
or U4549 (N_4549,N_3925,N_3111);
and U4550 (N_4550,N_3210,N_3474);
nand U4551 (N_4551,N_3260,N_3751);
nor U4552 (N_4552,N_3143,N_3432);
and U4553 (N_4553,N_3047,N_3869);
and U4554 (N_4554,N_3196,N_3023);
or U4555 (N_4555,N_3240,N_3223);
nand U4556 (N_4556,N_3213,N_3831);
or U4557 (N_4557,N_3912,N_3836);
nand U4558 (N_4558,N_3638,N_3242);
and U4559 (N_4559,N_3589,N_3600);
and U4560 (N_4560,N_3632,N_3934);
or U4561 (N_4561,N_3067,N_3298);
or U4562 (N_4562,N_3291,N_3064);
or U4563 (N_4563,N_3112,N_3670);
or U4564 (N_4564,N_3389,N_3719);
nand U4565 (N_4565,N_3071,N_3091);
nor U4566 (N_4566,N_3038,N_3160);
or U4567 (N_4567,N_3154,N_3105);
xor U4568 (N_4568,N_3041,N_3789);
or U4569 (N_4569,N_3419,N_3026);
and U4570 (N_4570,N_3134,N_3678);
and U4571 (N_4571,N_3282,N_3145);
nand U4572 (N_4572,N_3528,N_3828);
and U4573 (N_4573,N_3171,N_3924);
nor U4574 (N_4574,N_3367,N_3574);
and U4575 (N_4575,N_3247,N_3603);
or U4576 (N_4576,N_3789,N_3609);
or U4577 (N_4577,N_3921,N_3006);
and U4578 (N_4578,N_3999,N_3004);
and U4579 (N_4579,N_3317,N_3975);
nor U4580 (N_4580,N_3196,N_3225);
nand U4581 (N_4581,N_3590,N_3532);
and U4582 (N_4582,N_3500,N_3654);
nor U4583 (N_4583,N_3256,N_3392);
nor U4584 (N_4584,N_3734,N_3335);
nor U4585 (N_4585,N_3871,N_3702);
nor U4586 (N_4586,N_3739,N_3209);
nor U4587 (N_4587,N_3375,N_3857);
nor U4588 (N_4588,N_3934,N_3940);
nand U4589 (N_4589,N_3738,N_3722);
and U4590 (N_4590,N_3813,N_3569);
nand U4591 (N_4591,N_3355,N_3311);
nor U4592 (N_4592,N_3421,N_3407);
or U4593 (N_4593,N_3382,N_3402);
or U4594 (N_4594,N_3890,N_3460);
nand U4595 (N_4595,N_3905,N_3910);
nor U4596 (N_4596,N_3142,N_3542);
nand U4597 (N_4597,N_3653,N_3259);
nor U4598 (N_4598,N_3464,N_3443);
nor U4599 (N_4599,N_3657,N_3753);
or U4600 (N_4600,N_3489,N_3813);
nand U4601 (N_4601,N_3806,N_3684);
nand U4602 (N_4602,N_3685,N_3944);
nand U4603 (N_4603,N_3171,N_3464);
or U4604 (N_4604,N_3011,N_3535);
or U4605 (N_4605,N_3546,N_3633);
nand U4606 (N_4606,N_3999,N_3268);
or U4607 (N_4607,N_3020,N_3883);
nor U4608 (N_4608,N_3784,N_3024);
nor U4609 (N_4609,N_3608,N_3026);
or U4610 (N_4610,N_3530,N_3931);
or U4611 (N_4611,N_3776,N_3735);
or U4612 (N_4612,N_3232,N_3358);
or U4613 (N_4613,N_3523,N_3746);
nor U4614 (N_4614,N_3756,N_3016);
and U4615 (N_4615,N_3829,N_3895);
and U4616 (N_4616,N_3007,N_3390);
and U4617 (N_4617,N_3766,N_3398);
or U4618 (N_4618,N_3619,N_3687);
nand U4619 (N_4619,N_3656,N_3441);
or U4620 (N_4620,N_3110,N_3806);
nand U4621 (N_4621,N_3964,N_3095);
or U4622 (N_4622,N_3450,N_3074);
nor U4623 (N_4623,N_3883,N_3740);
nand U4624 (N_4624,N_3781,N_3723);
nor U4625 (N_4625,N_3467,N_3020);
xor U4626 (N_4626,N_3885,N_3509);
and U4627 (N_4627,N_3413,N_3641);
nand U4628 (N_4628,N_3644,N_3049);
and U4629 (N_4629,N_3702,N_3777);
or U4630 (N_4630,N_3580,N_3565);
nand U4631 (N_4631,N_3826,N_3915);
and U4632 (N_4632,N_3648,N_3805);
nor U4633 (N_4633,N_3332,N_3050);
nand U4634 (N_4634,N_3946,N_3484);
or U4635 (N_4635,N_3662,N_3348);
and U4636 (N_4636,N_3068,N_3882);
and U4637 (N_4637,N_3274,N_3246);
nand U4638 (N_4638,N_3199,N_3964);
nor U4639 (N_4639,N_3103,N_3574);
nor U4640 (N_4640,N_3139,N_3837);
and U4641 (N_4641,N_3624,N_3884);
and U4642 (N_4642,N_3594,N_3575);
nor U4643 (N_4643,N_3438,N_3485);
nor U4644 (N_4644,N_3944,N_3505);
nand U4645 (N_4645,N_3661,N_3570);
and U4646 (N_4646,N_3259,N_3817);
or U4647 (N_4647,N_3356,N_3864);
and U4648 (N_4648,N_3606,N_3351);
nand U4649 (N_4649,N_3193,N_3306);
nor U4650 (N_4650,N_3385,N_3070);
or U4651 (N_4651,N_3659,N_3752);
and U4652 (N_4652,N_3832,N_3889);
nor U4653 (N_4653,N_3915,N_3889);
or U4654 (N_4654,N_3975,N_3584);
or U4655 (N_4655,N_3074,N_3381);
nand U4656 (N_4656,N_3217,N_3351);
or U4657 (N_4657,N_3344,N_3876);
and U4658 (N_4658,N_3380,N_3065);
and U4659 (N_4659,N_3581,N_3814);
nand U4660 (N_4660,N_3288,N_3230);
and U4661 (N_4661,N_3103,N_3121);
or U4662 (N_4662,N_3614,N_3590);
and U4663 (N_4663,N_3545,N_3351);
and U4664 (N_4664,N_3220,N_3446);
or U4665 (N_4665,N_3890,N_3965);
or U4666 (N_4666,N_3431,N_3016);
nand U4667 (N_4667,N_3831,N_3442);
nand U4668 (N_4668,N_3355,N_3465);
or U4669 (N_4669,N_3309,N_3458);
nor U4670 (N_4670,N_3137,N_3712);
nand U4671 (N_4671,N_3424,N_3325);
nor U4672 (N_4672,N_3545,N_3232);
and U4673 (N_4673,N_3108,N_3705);
and U4674 (N_4674,N_3526,N_3413);
and U4675 (N_4675,N_3508,N_3716);
nand U4676 (N_4676,N_3820,N_3074);
or U4677 (N_4677,N_3536,N_3201);
nor U4678 (N_4678,N_3550,N_3755);
nor U4679 (N_4679,N_3194,N_3865);
or U4680 (N_4680,N_3763,N_3742);
nand U4681 (N_4681,N_3626,N_3519);
nand U4682 (N_4682,N_3805,N_3882);
nor U4683 (N_4683,N_3062,N_3503);
nor U4684 (N_4684,N_3183,N_3657);
or U4685 (N_4685,N_3830,N_3538);
nor U4686 (N_4686,N_3485,N_3901);
nand U4687 (N_4687,N_3835,N_3208);
nand U4688 (N_4688,N_3552,N_3861);
xor U4689 (N_4689,N_3617,N_3277);
nor U4690 (N_4690,N_3024,N_3006);
and U4691 (N_4691,N_3184,N_3311);
nor U4692 (N_4692,N_3188,N_3069);
nor U4693 (N_4693,N_3958,N_3507);
nand U4694 (N_4694,N_3486,N_3913);
and U4695 (N_4695,N_3382,N_3580);
or U4696 (N_4696,N_3281,N_3997);
nor U4697 (N_4697,N_3956,N_3572);
or U4698 (N_4698,N_3607,N_3606);
nor U4699 (N_4699,N_3726,N_3336);
nor U4700 (N_4700,N_3005,N_3321);
xnor U4701 (N_4701,N_3390,N_3793);
nand U4702 (N_4702,N_3103,N_3287);
nand U4703 (N_4703,N_3471,N_3589);
or U4704 (N_4704,N_3777,N_3567);
nand U4705 (N_4705,N_3079,N_3906);
and U4706 (N_4706,N_3541,N_3550);
or U4707 (N_4707,N_3341,N_3270);
or U4708 (N_4708,N_3267,N_3648);
or U4709 (N_4709,N_3498,N_3970);
and U4710 (N_4710,N_3205,N_3507);
nor U4711 (N_4711,N_3792,N_3093);
or U4712 (N_4712,N_3362,N_3058);
xor U4713 (N_4713,N_3388,N_3705);
nor U4714 (N_4714,N_3778,N_3397);
and U4715 (N_4715,N_3628,N_3166);
or U4716 (N_4716,N_3887,N_3120);
nand U4717 (N_4717,N_3196,N_3922);
nor U4718 (N_4718,N_3940,N_3615);
or U4719 (N_4719,N_3486,N_3201);
and U4720 (N_4720,N_3208,N_3812);
nand U4721 (N_4721,N_3553,N_3490);
nor U4722 (N_4722,N_3489,N_3630);
nor U4723 (N_4723,N_3211,N_3394);
and U4724 (N_4724,N_3987,N_3628);
nand U4725 (N_4725,N_3958,N_3851);
or U4726 (N_4726,N_3890,N_3631);
or U4727 (N_4727,N_3320,N_3048);
or U4728 (N_4728,N_3504,N_3060);
nor U4729 (N_4729,N_3442,N_3776);
nand U4730 (N_4730,N_3723,N_3257);
or U4731 (N_4731,N_3378,N_3524);
nand U4732 (N_4732,N_3512,N_3756);
nand U4733 (N_4733,N_3452,N_3475);
nor U4734 (N_4734,N_3954,N_3923);
xor U4735 (N_4735,N_3524,N_3227);
nor U4736 (N_4736,N_3328,N_3235);
or U4737 (N_4737,N_3309,N_3440);
nor U4738 (N_4738,N_3857,N_3475);
and U4739 (N_4739,N_3720,N_3812);
or U4740 (N_4740,N_3854,N_3510);
nor U4741 (N_4741,N_3503,N_3845);
or U4742 (N_4742,N_3518,N_3123);
and U4743 (N_4743,N_3172,N_3489);
nor U4744 (N_4744,N_3318,N_3776);
nor U4745 (N_4745,N_3822,N_3100);
and U4746 (N_4746,N_3127,N_3628);
and U4747 (N_4747,N_3274,N_3598);
nor U4748 (N_4748,N_3047,N_3943);
nor U4749 (N_4749,N_3920,N_3893);
nand U4750 (N_4750,N_3655,N_3780);
nor U4751 (N_4751,N_3775,N_3671);
nand U4752 (N_4752,N_3972,N_3797);
or U4753 (N_4753,N_3442,N_3694);
or U4754 (N_4754,N_3658,N_3580);
or U4755 (N_4755,N_3008,N_3429);
and U4756 (N_4756,N_3301,N_3611);
and U4757 (N_4757,N_3184,N_3587);
nor U4758 (N_4758,N_3350,N_3888);
nor U4759 (N_4759,N_3345,N_3357);
nor U4760 (N_4760,N_3403,N_3521);
and U4761 (N_4761,N_3542,N_3818);
nand U4762 (N_4762,N_3583,N_3374);
or U4763 (N_4763,N_3278,N_3907);
and U4764 (N_4764,N_3536,N_3684);
or U4765 (N_4765,N_3569,N_3760);
nor U4766 (N_4766,N_3797,N_3290);
nand U4767 (N_4767,N_3830,N_3900);
nor U4768 (N_4768,N_3273,N_3063);
nand U4769 (N_4769,N_3003,N_3198);
or U4770 (N_4770,N_3827,N_3153);
nand U4771 (N_4771,N_3607,N_3252);
and U4772 (N_4772,N_3455,N_3260);
nand U4773 (N_4773,N_3135,N_3910);
nand U4774 (N_4774,N_3830,N_3576);
nor U4775 (N_4775,N_3891,N_3314);
and U4776 (N_4776,N_3736,N_3342);
or U4777 (N_4777,N_3876,N_3788);
and U4778 (N_4778,N_3629,N_3263);
nand U4779 (N_4779,N_3897,N_3581);
nand U4780 (N_4780,N_3340,N_3257);
and U4781 (N_4781,N_3674,N_3967);
xor U4782 (N_4782,N_3342,N_3314);
and U4783 (N_4783,N_3328,N_3446);
nand U4784 (N_4784,N_3673,N_3465);
and U4785 (N_4785,N_3855,N_3094);
nand U4786 (N_4786,N_3477,N_3099);
and U4787 (N_4787,N_3335,N_3457);
or U4788 (N_4788,N_3257,N_3133);
nand U4789 (N_4789,N_3751,N_3631);
and U4790 (N_4790,N_3649,N_3043);
or U4791 (N_4791,N_3454,N_3749);
or U4792 (N_4792,N_3055,N_3097);
nor U4793 (N_4793,N_3981,N_3213);
nand U4794 (N_4794,N_3407,N_3743);
and U4795 (N_4795,N_3739,N_3814);
and U4796 (N_4796,N_3939,N_3594);
nand U4797 (N_4797,N_3632,N_3367);
nand U4798 (N_4798,N_3319,N_3557);
nor U4799 (N_4799,N_3336,N_3683);
and U4800 (N_4800,N_3303,N_3308);
nand U4801 (N_4801,N_3331,N_3560);
nand U4802 (N_4802,N_3238,N_3895);
and U4803 (N_4803,N_3824,N_3764);
or U4804 (N_4804,N_3681,N_3908);
nand U4805 (N_4805,N_3050,N_3308);
or U4806 (N_4806,N_3892,N_3781);
nand U4807 (N_4807,N_3021,N_3864);
and U4808 (N_4808,N_3687,N_3094);
nor U4809 (N_4809,N_3876,N_3831);
xnor U4810 (N_4810,N_3092,N_3498);
and U4811 (N_4811,N_3815,N_3894);
or U4812 (N_4812,N_3805,N_3854);
nor U4813 (N_4813,N_3875,N_3089);
and U4814 (N_4814,N_3159,N_3279);
nor U4815 (N_4815,N_3404,N_3162);
or U4816 (N_4816,N_3212,N_3397);
nor U4817 (N_4817,N_3582,N_3197);
and U4818 (N_4818,N_3081,N_3656);
and U4819 (N_4819,N_3668,N_3840);
and U4820 (N_4820,N_3675,N_3454);
and U4821 (N_4821,N_3910,N_3995);
and U4822 (N_4822,N_3980,N_3163);
nand U4823 (N_4823,N_3572,N_3057);
nand U4824 (N_4824,N_3672,N_3731);
nand U4825 (N_4825,N_3990,N_3891);
nand U4826 (N_4826,N_3854,N_3002);
or U4827 (N_4827,N_3770,N_3724);
nor U4828 (N_4828,N_3191,N_3260);
nor U4829 (N_4829,N_3610,N_3586);
or U4830 (N_4830,N_3408,N_3959);
nand U4831 (N_4831,N_3472,N_3960);
nand U4832 (N_4832,N_3638,N_3794);
nand U4833 (N_4833,N_3785,N_3545);
nor U4834 (N_4834,N_3035,N_3158);
xor U4835 (N_4835,N_3810,N_3360);
nand U4836 (N_4836,N_3702,N_3037);
nor U4837 (N_4837,N_3842,N_3986);
nor U4838 (N_4838,N_3548,N_3896);
or U4839 (N_4839,N_3136,N_3805);
nand U4840 (N_4840,N_3922,N_3231);
nor U4841 (N_4841,N_3718,N_3626);
nand U4842 (N_4842,N_3154,N_3056);
nand U4843 (N_4843,N_3326,N_3531);
and U4844 (N_4844,N_3236,N_3635);
nor U4845 (N_4845,N_3072,N_3506);
nand U4846 (N_4846,N_3478,N_3833);
and U4847 (N_4847,N_3127,N_3926);
nand U4848 (N_4848,N_3158,N_3433);
or U4849 (N_4849,N_3639,N_3876);
nor U4850 (N_4850,N_3578,N_3168);
nand U4851 (N_4851,N_3257,N_3175);
or U4852 (N_4852,N_3384,N_3093);
or U4853 (N_4853,N_3341,N_3324);
nor U4854 (N_4854,N_3187,N_3121);
nor U4855 (N_4855,N_3164,N_3553);
or U4856 (N_4856,N_3085,N_3248);
nor U4857 (N_4857,N_3651,N_3596);
nand U4858 (N_4858,N_3202,N_3338);
or U4859 (N_4859,N_3911,N_3595);
nand U4860 (N_4860,N_3315,N_3881);
or U4861 (N_4861,N_3779,N_3325);
or U4862 (N_4862,N_3547,N_3615);
and U4863 (N_4863,N_3451,N_3226);
nor U4864 (N_4864,N_3184,N_3633);
nand U4865 (N_4865,N_3956,N_3746);
or U4866 (N_4866,N_3683,N_3606);
nor U4867 (N_4867,N_3857,N_3357);
nor U4868 (N_4868,N_3380,N_3960);
and U4869 (N_4869,N_3330,N_3879);
nand U4870 (N_4870,N_3713,N_3784);
nor U4871 (N_4871,N_3711,N_3976);
nand U4872 (N_4872,N_3676,N_3558);
nand U4873 (N_4873,N_3456,N_3651);
nand U4874 (N_4874,N_3840,N_3342);
nor U4875 (N_4875,N_3371,N_3305);
nand U4876 (N_4876,N_3294,N_3458);
and U4877 (N_4877,N_3361,N_3180);
or U4878 (N_4878,N_3458,N_3941);
and U4879 (N_4879,N_3417,N_3057);
and U4880 (N_4880,N_3859,N_3635);
or U4881 (N_4881,N_3467,N_3575);
nand U4882 (N_4882,N_3340,N_3450);
xnor U4883 (N_4883,N_3618,N_3498);
nand U4884 (N_4884,N_3200,N_3869);
and U4885 (N_4885,N_3241,N_3379);
nor U4886 (N_4886,N_3451,N_3821);
and U4887 (N_4887,N_3545,N_3040);
and U4888 (N_4888,N_3566,N_3572);
nor U4889 (N_4889,N_3354,N_3653);
nand U4890 (N_4890,N_3977,N_3091);
nor U4891 (N_4891,N_3737,N_3714);
and U4892 (N_4892,N_3420,N_3740);
or U4893 (N_4893,N_3571,N_3896);
nor U4894 (N_4894,N_3767,N_3676);
nand U4895 (N_4895,N_3702,N_3051);
and U4896 (N_4896,N_3091,N_3228);
nor U4897 (N_4897,N_3409,N_3896);
nand U4898 (N_4898,N_3482,N_3700);
or U4899 (N_4899,N_3211,N_3589);
or U4900 (N_4900,N_3423,N_3490);
and U4901 (N_4901,N_3813,N_3354);
or U4902 (N_4902,N_3705,N_3399);
and U4903 (N_4903,N_3616,N_3543);
nand U4904 (N_4904,N_3065,N_3936);
or U4905 (N_4905,N_3468,N_3909);
or U4906 (N_4906,N_3810,N_3249);
or U4907 (N_4907,N_3166,N_3853);
and U4908 (N_4908,N_3926,N_3092);
and U4909 (N_4909,N_3964,N_3396);
and U4910 (N_4910,N_3653,N_3547);
nand U4911 (N_4911,N_3873,N_3142);
nor U4912 (N_4912,N_3923,N_3163);
and U4913 (N_4913,N_3771,N_3941);
or U4914 (N_4914,N_3374,N_3216);
nor U4915 (N_4915,N_3847,N_3090);
and U4916 (N_4916,N_3576,N_3632);
nor U4917 (N_4917,N_3859,N_3619);
or U4918 (N_4918,N_3516,N_3552);
or U4919 (N_4919,N_3553,N_3572);
or U4920 (N_4920,N_3297,N_3094);
nand U4921 (N_4921,N_3096,N_3441);
and U4922 (N_4922,N_3143,N_3073);
nor U4923 (N_4923,N_3586,N_3941);
or U4924 (N_4924,N_3313,N_3125);
and U4925 (N_4925,N_3883,N_3785);
nand U4926 (N_4926,N_3904,N_3361);
and U4927 (N_4927,N_3051,N_3408);
and U4928 (N_4928,N_3555,N_3069);
or U4929 (N_4929,N_3919,N_3611);
or U4930 (N_4930,N_3004,N_3731);
nand U4931 (N_4931,N_3836,N_3003);
or U4932 (N_4932,N_3415,N_3030);
nor U4933 (N_4933,N_3741,N_3356);
and U4934 (N_4934,N_3726,N_3851);
xnor U4935 (N_4935,N_3465,N_3239);
or U4936 (N_4936,N_3897,N_3534);
and U4937 (N_4937,N_3858,N_3545);
or U4938 (N_4938,N_3596,N_3816);
nand U4939 (N_4939,N_3651,N_3971);
and U4940 (N_4940,N_3253,N_3454);
nand U4941 (N_4941,N_3727,N_3297);
or U4942 (N_4942,N_3301,N_3288);
nand U4943 (N_4943,N_3396,N_3926);
nor U4944 (N_4944,N_3864,N_3482);
nand U4945 (N_4945,N_3465,N_3800);
nor U4946 (N_4946,N_3183,N_3561);
and U4947 (N_4947,N_3804,N_3126);
and U4948 (N_4948,N_3552,N_3934);
or U4949 (N_4949,N_3362,N_3443);
and U4950 (N_4950,N_3839,N_3476);
nand U4951 (N_4951,N_3574,N_3645);
nor U4952 (N_4952,N_3106,N_3112);
or U4953 (N_4953,N_3322,N_3808);
nor U4954 (N_4954,N_3244,N_3159);
nand U4955 (N_4955,N_3267,N_3498);
or U4956 (N_4956,N_3273,N_3897);
nor U4957 (N_4957,N_3279,N_3117);
nand U4958 (N_4958,N_3273,N_3582);
nor U4959 (N_4959,N_3780,N_3576);
or U4960 (N_4960,N_3741,N_3297);
or U4961 (N_4961,N_3709,N_3004);
nand U4962 (N_4962,N_3263,N_3752);
or U4963 (N_4963,N_3447,N_3102);
nor U4964 (N_4964,N_3168,N_3355);
nor U4965 (N_4965,N_3614,N_3509);
and U4966 (N_4966,N_3078,N_3755);
nand U4967 (N_4967,N_3995,N_3008);
or U4968 (N_4968,N_3165,N_3796);
nand U4969 (N_4969,N_3871,N_3572);
nor U4970 (N_4970,N_3324,N_3398);
or U4971 (N_4971,N_3286,N_3788);
and U4972 (N_4972,N_3995,N_3587);
nor U4973 (N_4973,N_3852,N_3436);
nand U4974 (N_4974,N_3564,N_3680);
nor U4975 (N_4975,N_3773,N_3660);
and U4976 (N_4976,N_3467,N_3262);
and U4977 (N_4977,N_3425,N_3029);
nor U4978 (N_4978,N_3928,N_3295);
nand U4979 (N_4979,N_3788,N_3562);
nor U4980 (N_4980,N_3323,N_3472);
nor U4981 (N_4981,N_3970,N_3240);
or U4982 (N_4982,N_3927,N_3078);
or U4983 (N_4983,N_3088,N_3071);
and U4984 (N_4984,N_3090,N_3207);
or U4985 (N_4985,N_3388,N_3332);
nand U4986 (N_4986,N_3483,N_3781);
nand U4987 (N_4987,N_3554,N_3096);
nor U4988 (N_4988,N_3754,N_3189);
nand U4989 (N_4989,N_3748,N_3733);
or U4990 (N_4990,N_3390,N_3389);
nand U4991 (N_4991,N_3465,N_3144);
nand U4992 (N_4992,N_3659,N_3317);
and U4993 (N_4993,N_3708,N_3576);
and U4994 (N_4994,N_3761,N_3375);
nand U4995 (N_4995,N_3416,N_3921);
and U4996 (N_4996,N_3745,N_3300);
or U4997 (N_4997,N_3770,N_3290);
nor U4998 (N_4998,N_3649,N_3321);
nor U4999 (N_4999,N_3773,N_3158);
nor U5000 (N_5000,N_4152,N_4160);
nand U5001 (N_5001,N_4514,N_4953);
nor U5002 (N_5002,N_4841,N_4333);
nand U5003 (N_5003,N_4158,N_4422);
or U5004 (N_5004,N_4682,N_4190);
or U5005 (N_5005,N_4178,N_4449);
nor U5006 (N_5006,N_4957,N_4390);
nor U5007 (N_5007,N_4576,N_4181);
and U5008 (N_5008,N_4891,N_4496);
nor U5009 (N_5009,N_4579,N_4804);
nor U5010 (N_5010,N_4939,N_4300);
nor U5011 (N_5011,N_4136,N_4216);
or U5012 (N_5012,N_4272,N_4527);
nor U5013 (N_5013,N_4958,N_4137);
and U5014 (N_5014,N_4836,N_4033);
nand U5015 (N_5015,N_4481,N_4297);
and U5016 (N_5016,N_4569,N_4290);
or U5017 (N_5017,N_4826,N_4821);
nand U5018 (N_5018,N_4961,N_4519);
and U5019 (N_5019,N_4327,N_4684);
and U5020 (N_5020,N_4208,N_4285);
nand U5021 (N_5021,N_4001,N_4938);
or U5022 (N_5022,N_4313,N_4164);
nor U5023 (N_5023,N_4697,N_4323);
nor U5024 (N_5024,N_4125,N_4774);
and U5025 (N_5025,N_4265,N_4976);
xnor U5026 (N_5026,N_4256,N_4713);
xnor U5027 (N_5027,N_4411,N_4171);
and U5028 (N_5028,N_4986,N_4515);
nand U5029 (N_5029,N_4444,N_4104);
or U5030 (N_5030,N_4611,N_4161);
nor U5031 (N_5031,N_4577,N_4420);
and U5032 (N_5032,N_4544,N_4074);
nor U5033 (N_5033,N_4346,N_4644);
nand U5034 (N_5034,N_4029,N_4893);
nor U5035 (N_5035,N_4546,N_4773);
nor U5036 (N_5036,N_4215,N_4824);
nor U5037 (N_5037,N_4360,N_4944);
and U5038 (N_5038,N_4874,N_4548);
or U5039 (N_5039,N_4570,N_4461);
nor U5040 (N_5040,N_4562,N_4812);
and U5041 (N_5041,N_4348,N_4406);
nand U5042 (N_5042,N_4009,N_4431);
and U5043 (N_5043,N_4022,N_4670);
nand U5044 (N_5044,N_4652,N_4226);
nand U5045 (N_5045,N_4879,N_4207);
nand U5046 (N_5046,N_4643,N_4105);
or U5047 (N_5047,N_4989,N_4084);
nor U5048 (N_5048,N_4842,N_4219);
nand U5049 (N_5049,N_4249,N_4720);
nor U5050 (N_5050,N_4479,N_4717);
nand U5051 (N_5051,N_4484,N_4759);
and U5052 (N_5052,N_4992,N_4377);
or U5053 (N_5053,N_4004,N_4385);
nor U5054 (N_5054,N_4988,N_4371);
or U5055 (N_5055,N_4531,N_4292);
or U5056 (N_5056,N_4977,N_4097);
nor U5057 (N_5057,N_4808,N_4474);
nand U5058 (N_5058,N_4967,N_4554);
nor U5059 (N_5059,N_4102,N_4810);
and U5060 (N_5060,N_4610,N_4495);
nor U5061 (N_5061,N_4250,N_4182);
or U5062 (N_5062,N_4294,N_4044);
nand U5063 (N_5063,N_4419,N_4445);
and U5064 (N_5064,N_4511,N_4082);
and U5065 (N_5065,N_4231,N_4845);
nor U5066 (N_5066,N_4195,N_4590);
xnor U5067 (N_5067,N_4241,N_4919);
nor U5068 (N_5068,N_4426,N_4379);
or U5069 (N_5069,N_4786,N_4897);
or U5070 (N_5070,N_4480,N_4264);
or U5071 (N_5071,N_4424,N_4396);
nor U5072 (N_5072,N_4601,N_4395);
nor U5073 (N_5073,N_4526,N_4017);
or U5074 (N_5074,N_4080,N_4817);
nor U5075 (N_5075,N_4439,N_4947);
nor U5076 (N_5076,N_4870,N_4334);
and U5077 (N_5077,N_4413,N_4352);
nor U5078 (N_5078,N_4530,N_4251);
or U5079 (N_5079,N_4330,N_4726);
nand U5080 (N_5080,N_4112,N_4437);
and U5081 (N_5081,N_4894,N_4863);
nor U5082 (N_5082,N_4067,N_4521);
nor U5083 (N_5083,N_4245,N_4796);
or U5084 (N_5084,N_4884,N_4301);
and U5085 (N_5085,N_4397,N_4864);
nor U5086 (N_5086,N_4750,N_4010);
and U5087 (N_5087,N_4254,N_4775);
and U5088 (N_5088,N_4013,N_4532);
and U5089 (N_5089,N_4131,N_4647);
or U5090 (N_5090,N_4429,N_4200);
nor U5091 (N_5091,N_4491,N_4428);
nand U5092 (N_5092,N_4686,N_4452);
and U5093 (N_5093,N_4937,N_4176);
and U5094 (N_5094,N_4941,N_4831);
nor U5095 (N_5095,N_4175,N_4315);
nor U5096 (N_5096,N_4908,N_4517);
and U5097 (N_5097,N_4163,N_4571);
nor U5098 (N_5098,N_4132,N_4659);
or U5099 (N_5099,N_4578,N_4706);
nor U5100 (N_5100,N_4099,N_4676);
and U5101 (N_5101,N_4673,N_4153);
or U5102 (N_5102,N_4165,N_4685);
xor U5103 (N_5103,N_4996,N_4769);
nor U5104 (N_5104,N_4277,N_4118);
or U5105 (N_5105,N_4928,N_4971);
or U5106 (N_5106,N_4573,N_4316);
or U5107 (N_5107,N_4954,N_4613);
and U5108 (N_5108,N_4935,N_4784);
nor U5109 (N_5109,N_4409,N_4000);
and U5110 (N_5110,N_4625,N_4197);
nand U5111 (N_5111,N_4753,N_4851);
nand U5112 (N_5112,N_4933,N_4718);
nand U5113 (N_5113,N_4350,N_4075);
nand U5114 (N_5114,N_4233,N_4036);
nand U5115 (N_5115,N_4756,N_4145);
or U5116 (N_5116,N_4667,N_4557);
nor U5117 (N_5117,N_4225,N_4122);
and U5118 (N_5118,N_4843,N_4146);
and U5119 (N_5119,N_4932,N_4096);
and U5120 (N_5120,N_4525,N_4690);
and U5121 (N_5121,N_4014,N_4621);
nand U5122 (N_5122,N_4787,N_4120);
nor U5123 (N_5123,N_4997,N_4159);
and U5124 (N_5124,N_4539,N_4493);
or U5125 (N_5125,N_4142,N_4952);
or U5126 (N_5126,N_4353,N_4465);
nor U5127 (N_5127,N_4622,N_4595);
or U5128 (N_5128,N_4069,N_4835);
nor U5129 (N_5129,N_4993,N_4030);
and U5130 (N_5130,N_4415,N_4980);
or U5131 (N_5131,N_4202,N_4361);
and U5132 (N_5132,N_4561,N_4306);
or U5133 (N_5133,N_4357,N_4711);
xor U5134 (N_5134,N_4708,N_4403);
nand U5135 (N_5135,N_4740,N_4741);
nor U5136 (N_5136,N_4612,N_4898);
or U5137 (N_5137,N_4778,N_4979);
and U5138 (N_5138,N_4995,N_4653);
nor U5139 (N_5139,N_4901,N_4110);
nor U5140 (N_5140,N_4721,N_4473);
nor U5141 (N_5141,N_4349,N_4263);
nand U5142 (N_5142,N_4949,N_4078);
and U5143 (N_5143,N_4459,N_4365);
and U5144 (N_5144,N_4128,N_4991);
and U5145 (N_5145,N_4776,N_4288);
or U5146 (N_5146,N_4257,N_4701);
and U5147 (N_5147,N_4599,N_4443);
and U5148 (N_5148,N_4543,N_4564);
nand U5149 (N_5149,N_4224,N_4303);
and U5150 (N_5150,N_4133,N_4869);
nand U5151 (N_5151,N_4111,N_4608);
nand U5152 (N_5152,N_4923,N_4978);
and U5153 (N_5153,N_4326,N_4085);
or U5154 (N_5154,N_4885,N_4281);
and U5155 (N_5155,N_4631,N_4130);
and U5156 (N_5156,N_4402,N_4803);
nand U5157 (N_5157,N_4948,N_4304);
or U5158 (N_5158,N_4559,N_4744);
nand U5159 (N_5159,N_4144,N_4309);
nor U5160 (N_5160,N_4286,N_4049);
and U5161 (N_5161,N_4743,N_4704);
nand U5162 (N_5162,N_4909,N_4668);
nor U5163 (N_5163,N_4512,N_4018);
or U5164 (N_5164,N_4849,N_4438);
and U5165 (N_5165,N_4283,N_4699);
nand U5166 (N_5166,N_4765,N_4951);
or U5167 (N_5167,N_4794,N_4296);
or U5168 (N_5168,N_4139,N_4770);
or U5169 (N_5169,N_4834,N_4098);
and U5170 (N_5170,N_4848,N_4974);
or U5171 (N_5171,N_4584,N_4478);
or U5172 (N_5172,N_4271,N_4269);
nor U5173 (N_5173,N_4023,N_4827);
nor U5174 (N_5174,N_4077,N_4401);
and U5175 (N_5175,N_4041,N_4464);
nand U5176 (N_5176,N_4983,N_4068);
or U5177 (N_5177,N_4063,N_4883);
nor U5178 (N_5178,N_4083,N_4691);
nand U5179 (N_5179,N_4031,N_4696);
nand U5180 (N_5180,N_4114,N_4907);
nand U5181 (N_5181,N_4628,N_4038);
xor U5182 (N_5182,N_4679,N_4966);
nor U5183 (N_5183,N_4861,N_4729);
or U5184 (N_5184,N_4867,N_4963);
and U5185 (N_5185,N_4700,N_4275);
nand U5186 (N_5186,N_4337,N_4423);
nor U5187 (N_5187,N_4039,N_4934);
nand U5188 (N_5188,N_4592,N_4232);
and U5189 (N_5189,N_4282,N_4730);
and U5190 (N_5190,N_4727,N_4430);
xnor U5191 (N_5191,N_4661,N_4026);
nor U5192 (N_5192,N_4284,N_4506);
or U5193 (N_5193,N_4565,N_4258);
or U5194 (N_5194,N_4732,N_4688);
and U5195 (N_5195,N_4633,N_4735);
and U5196 (N_5196,N_4280,N_4196);
nor U5197 (N_5197,N_4143,N_4545);
nor U5198 (N_5198,N_4243,N_4179);
nand U5199 (N_5199,N_4081,N_4866);
or U5200 (N_5200,N_4193,N_4150);
or U5201 (N_5201,N_4307,N_4220);
nor U5202 (N_5202,N_4797,N_4582);
or U5203 (N_5203,N_4781,N_4008);
and U5204 (N_5204,N_4844,N_4779);
or U5205 (N_5205,N_4270,N_4343);
nand U5206 (N_5206,N_4830,N_4542);
or U5207 (N_5207,N_4820,N_4722);
nand U5208 (N_5208,N_4368,N_4126);
or U5209 (N_5209,N_4965,N_4508);
nand U5210 (N_5210,N_4680,N_4322);
and U5211 (N_5211,N_4448,N_4335);
or U5212 (N_5212,N_4016,N_4522);
or U5213 (N_5213,N_4692,N_4556);
nor U5214 (N_5214,N_4677,N_4191);
or U5215 (N_5215,N_4453,N_4738);
nand U5216 (N_5216,N_4823,N_4341);
nand U5217 (N_5217,N_4734,N_4210);
or U5218 (N_5218,N_4550,N_4320);
and U5219 (N_5219,N_4091,N_4651);
and U5220 (N_5220,N_4975,N_4815);
nor U5221 (N_5221,N_4043,N_4833);
nor U5222 (N_5222,N_4054,N_4498);
and U5223 (N_5223,N_4760,N_4355);
xor U5224 (N_5224,N_4956,N_4062);
or U5225 (N_5225,N_4064,N_4056);
and U5226 (N_5226,N_4623,N_4308);
and U5227 (N_5227,N_4212,N_4683);
and U5228 (N_5228,N_4324,N_4529);
and U5229 (N_5229,N_4764,N_4180);
nor U5230 (N_5230,N_4393,N_4962);
nor U5231 (N_5231,N_4540,N_4969);
or U5232 (N_5232,N_4558,N_4689);
xor U5233 (N_5233,N_4758,N_4751);
and U5234 (N_5234,N_4593,N_4372);
xor U5235 (N_5235,N_4945,N_4418);
and U5236 (N_5236,N_4340,N_4339);
nand U5237 (N_5237,N_4373,N_4655);
nand U5238 (N_5238,N_4253,N_4881);
and U5239 (N_5239,N_4436,N_4076);
nor U5240 (N_5240,N_4342,N_4211);
and U5241 (N_5241,N_4828,N_4414);
or U5242 (N_5242,N_4509,N_4305);
nor U5243 (N_5243,N_4050,N_4871);
or U5244 (N_5244,N_4467,N_4138);
and U5245 (N_5245,N_4186,N_4501);
nand U5246 (N_5246,N_4737,N_4020);
and U5247 (N_5247,N_4586,N_4234);
nor U5248 (N_5248,N_4172,N_4376);
or U5249 (N_5249,N_4603,N_4053);
nor U5250 (N_5250,N_4793,N_4746);
and U5251 (N_5251,N_4581,N_4490);
nor U5252 (N_5252,N_4606,N_4747);
and U5253 (N_5253,N_4410,N_4433);
nor U5254 (N_5254,N_4624,N_4061);
and U5255 (N_5255,N_4950,N_4547);
and U5256 (N_5256,N_4669,N_4329);
nor U5257 (N_5257,N_4273,N_4440);
nand U5258 (N_5258,N_4011,N_4538);
and U5259 (N_5259,N_4888,N_4640);
nor U5260 (N_5260,N_4940,N_4147);
and U5261 (N_5261,N_4100,N_4405);
nand U5262 (N_5262,N_4638,N_4347);
nand U5263 (N_5263,N_4895,N_4239);
nand U5264 (N_5264,N_4914,N_4777);
or U5265 (N_5265,N_4968,N_4850);
and U5266 (N_5266,N_4451,N_4757);
nand U5267 (N_5267,N_4795,N_4752);
nand U5268 (N_5268,N_4497,N_4154);
nor U5269 (N_5269,N_4374,N_4537);
or U5270 (N_5270,N_4536,N_4905);
or U5271 (N_5271,N_4607,N_4763);
and U5272 (N_5272,N_4214,N_4380);
and U5273 (N_5273,N_4121,N_4598);
nor U5274 (N_5274,N_4148,N_4442);
or U5275 (N_5275,N_4802,N_4472);
nor U5276 (N_5276,N_4338,N_4040);
nand U5277 (N_5277,N_4681,N_4170);
nand U5278 (N_5278,N_4089,N_4911);
nand U5279 (N_5279,N_4441,N_4252);
or U5280 (N_5280,N_4614,N_4173);
nor U5281 (N_5281,N_4635,N_4748);
or U5282 (N_5282,N_4242,N_4505);
nand U5283 (N_5283,N_4920,N_4177);
nor U5284 (N_5284,N_4310,N_4388);
and U5285 (N_5285,N_4336,N_4768);
and U5286 (N_5286,N_4025,N_4609);
nand U5287 (N_5287,N_4930,N_4293);
and U5288 (N_5288,N_4789,N_4520);
nand U5289 (N_5289,N_4492,N_4618);
nand U5290 (N_5290,N_4123,N_4344);
nand U5291 (N_5291,N_4970,N_4500);
nor U5292 (N_5292,N_4858,N_4446);
nand U5293 (N_5293,N_4312,N_4615);
and U5294 (N_5294,N_4065,N_4616);
or U5295 (N_5295,N_4872,N_4518);
nor U5296 (N_5296,N_4714,N_4356);
or U5297 (N_5297,N_4189,N_4859);
nand U5298 (N_5298,N_4917,N_4626);
nor U5299 (N_5299,N_4860,N_4057);
and U5300 (N_5300,N_4523,N_4407);
and U5301 (N_5301,N_4602,N_4002);
or U5302 (N_5302,N_4227,N_4915);
and U5303 (N_5303,N_4151,N_4351);
or U5304 (N_5304,N_4364,N_4596);
nand U5305 (N_5305,N_4024,N_4149);
nor U5306 (N_5306,N_4311,N_4092);
nor U5307 (N_5307,N_4432,N_4882);
and U5308 (N_5308,N_4597,N_4516);
and U5309 (N_5309,N_4731,N_4903);
or U5310 (N_5310,N_4274,N_4627);
and U5311 (N_5311,N_4006,N_4761);
nor U5312 (N_5312,N_4421,N_4246);
or U5313 (N_5313,N_4955,N_4382);
nand U5314 (N_5314,N_4665,N_4055);
nor U5315 (N_5315,N_4630,N_4213);
and U5316 (N_5316,N_4739,N_4391);
and U5317 (N_5317,N_4916,N_4456);
nand U5318 (N_5318,N_4460,N_4476);
nor U5319 (N_5319,N_4814,N_4332);
and U5320 (N_5320,N_4591,N_4719);
nor U5321 (N_5321,N_4093,N_4325);
nand U5322 (N_5322,N_4389,N_4267);
nand U5323 (N_5323,N_4218,N_4399);
nand U5324 (N_5324,N_4555,N_4892);
nor U5325 (N_5325,N_4887,N_4837);
nand U5326 (N_5326,N_4244,N_4455);
nand U5327 (N_5327,N_4910,N_4946);
or U5328 (N_5328,N_4103,N_4780);
nand U5329 (N_5329,N_4847,N_4184);
nor U5330 (N_5330,N_4675,N_4839);
nor U5331 (N_5331,N_4922,N_4936);
nor U5332 (N_5332,N_4217,N_4192);
nor U5333 (N_5333,N_4733,N_4878);
nand U5334 (N_5334,N_4299,N_4646);
and U5335 (N_5335,N_4657,N_4563);
or U5336 (N_5336,N_4899,N_4771);
and U5337 (N_5337,N_4567,N_4378);
nor U5338 (N_5338,N_4749,N_4902);
nor U5339 (N_5339,N_4412,N_4641);
and U5340 (N_5340,N_4999,N_4801);
and U5341 (N_5341,N_4155,N_4829);
nor U5342 (N_5342,N_4375,N_4106);
and U5343 (N_5343,N_4483,N_4058);
and U5344 (N_5344,N_4594,N_4021);
nor U5345 (N_5345,N_4742,N_4047);
nand U5346 (N_5346,N_4560,N_4007);
or U5347 (N_5347,N_4513,N_4856);
and U5348 (N_5348,N_4664,N_4620);
nor U5349 (N_5349,N_4925,N_4987);
or U5350 (N_5350,N_4381,N_4066);
or U5351 (N_5351,N_4012,N_4059);
nor U5352 (N_5352,N_4115,N_4416);
nand U5353 (N_5353,N_4921,N_4931);
nor U5354 (N_5354,N_4822,N_4398);
and U5355 (N_5355,N_4317,N_4629);
nand U5356 (N_5356,N_4551,N_4832);
nor U5357 (N_5357,N_4427,N_4129);
or U5358 (N_5358,N_4658,N_4087);
or U5359 (N_5359,N_4754,N_4188);
or U5360 (N_5360,N_4857,N_4205);
xor U5361 (N_5361,N_4201,N_4240);
nand U5362 (N_5362,N_4725,N_4799);
and U5363 (N_5363,N_4702,N_4943);
nor U5364 (N_5364,N_4485,N_4783);
nor U5365 (N_5365,N_4666,N_4482);
nor U5366 (N_5366,N_4468,N_4052);
nand U5367 (N_5367,N_4141,N_4463);
xnor U5368 (N_5368,N_4383,N_4086);
nor U5369 (N_5369,N_4117,N_4238);
and U5370 (N_5370,N_4868,N_4805);
and U5371 (N_5371,N_4846,N_4574);
nor U5372 (N_5372,N_4865,N_4094);
or U5373 (N_5373,N_4877,N_4709);
and U5374 (N_5374,N_4107,N_4672);
and U5375 (N_5375,N_4502,N_4425);
and U5376 (N_5376,N_4223,N_4457);
or U5377 (N_5377,N_4674,N_4876);
and U5378 (N_5378,N_4712,N_4964);
nand U5379 (N_5379,N_4985,N_4228);
nand U5380 (N_5380,N_4694,N_4134);
nor U5381 (N_5381,N_4650,N_4209);
nand U5382 (N_5382,N_4462,N_4255);
nor U5383 (N_5383,N_4345,N_4116);
or U5384 (N_5384,N_4203,N_4693);
nand U5385 (N_5385,N_4278,N_4302);
nor U5386 (N_5386,N_4806,N_4073);
nor U5387 (N_5387,N_4417,N_4745);
nor U5388 (N_5388,N_4528,N_4855);
nand U5389 (N_5389,N_4541,N_4477);
nor U5390 (N_5390,N_4321,N_4095);
and U5391 (N_5391,N_4504,N_4807);
nor U5392 (N_5392,N_4268,N_4162);
nand U5393 (N_5393,N_4716,N_4929);
nor U5394 (N_5394,N_4235,N_4762);
nand U5395 (N_5395,N_4384,N_4392);
nor U5396 (N_5396,N_4572,N_4568);
or U5397 (N_5397,N_4494,N_4071);
nand U5398 (N_5398,N_4705,N_4101);
or U5399 (N_5399,N_4072,N_4328);
or U5400 (N_5400,N_4318,N_4369);
nor U5401 (N_5401,N_4724,N_4221);
or U5402 (N_5402,N_4656,N_4470);
nor U5403 (N_5403,N_4488,N_4587);
or U5404 (N_5404,N_4359,N_4792);
nand U5405 (N_5405,N_4486,N_4019);
or U5406 (N_5406,N_4875,N_4354);
or U5407 (N_5407,N_4135,N_4982);
nand U5408 (N_5408,N_4404,N_4552);
and U5409 (N_5409,N_4510,N_4589);
nand U5410 (N_5410,N_4051,N_4818);
and U5411 (N_5411,N_4088,N_4533);
and U5412 (N_5412,N_4194,N_4167);
nand U5413 (N_5413,N_4654,N_4998);
nand U5414 (N_5414,N_4157,N_4639);
or U5415 (N_5415,N_4015,N_4813);
nor U5416 (N_5416,N_4634,N_4649);
nor U5417 (N_5417,N_4926,N_4434);
and U5418 (N_5418,N_4553,N_4108);
nor U5419 (N_5419,N_4791,N_4788);
or U5420 (N_5420,N_4687,N_4906);
or U5421 (N_5421,N_4663,N_4032);
nand U5422 (N_5422,N_4972,N_4840);
or U5423 (N_5423,N_4912,N_4862);
or U5424 (N_5424,N_4660,N_4723);
and U5425 (N_5425,N_4266,N_4904);
nand U5426 (N_5426,N_4852,N_4604);
or U5427 (N_5427,N_4109,N_4048);
and U5428 (N_5428,N_4045,N_4466);
nor U5429 (N_5429,N_4005,N_4187);
and U5430 (N_5430,N_4295,N_4489);
and U5431 (N_5431,N_4767,N_4671);
nand U5432 (N_5432,N_4291,N_4535);
and U5433 (N_5433,N_4447,N_4174);
or U5434 (N_5434,N_4703,N_4471);
or U5435 (N_5435,N_4960,N_4499);
nand U5436 (N_5436,N_4942,N_4798);
nand U5437 (N_5437,N_4825,N_4695);
or U5438 (N_5438,N_4637,N_4782);
nor U5439 (N_5439,N_4838,N_4236);
nand U5440 (N_5440,N_4617,N_4168);
nor U5441 (N_5441,N_4169,N_4619);
nand U5442 (N_5442,N_4636,N_4319);
or U5443 (N_5443,N_4698,N_4222);
nand U5444 (N_5444,N_4262,N_4800);
or U5445 (N_5445,N_4583,N_4259);
or U5446 (N_5446,N_4816,N_4707);
or U5447 (N_5447,N_4276,N_4090);
nor U5448 (N_5448,N_4183,N_4819);
and U5449 (N_5449,N_4853,N_4386);
nor U5450 (N_5450,N_4715,N_4454);
and U5451 (N_5451,N_4549,N_4766);
or U5452 (N_5452,N_4632,N_4642);
nand U5453 (N_5453,N_4896,N_4140);
nor U5454 (N_5454,N_4575,N_4206);
or U5455 (N_5455,N_4450,N_4503);
nand U5456 (N_5456,N_4229,N_4678);
nor U5457 (N_5457,N_4811,N_4873);
and U5458 (N_5458,N_4886,N_4469);
nand U5459 (N_5459,N_4534,N_4900);
and U5460 (N_5460,N_4854,N_4287);
and U5461 (N_5461,N_4918,N_4124);
nand U5462 (N_5462,N_4366,N_4247);
and U5463 (N_5463,N_4362,N_4566);
or U5464 (N_5464,N_4199,N_4728);
and U5465 (N_5465,N_4990,N_4710);
or U5466 (N_5466,N_4890,N_4166);
or U5467 (N_5467,N_4261,N_4984);
nor U5468 (N_5468,N_4435,N_4959);
nor U5469 (N_5469,N_4973,N_4248);
and U5470 (N_5470,N_4198,N_4331);
xnor U5471 (N_5471,N_4037,N_4237);
and U5472 (N_5472,N_4367,N_4034);
and U5473 (N_5473,N_4585,N_4028);
and U5474 (N_5474,N_4475,N_4279);
and U5475 (N_5475,N_4662,N_4314);
xor U5476 (N_5476,N_4070,N_4408);
nand U5477 (N_5477,N_4927,N_4772);
nor U5478 (N_5478,N_4079,N_4046);
or U5479 (N_5479,N_4648,N_4042);
nor U5480 (N_5480,N_4524,N_4394);
nor U5481 (N_5481,N_4880,N_4458);
nor U5482 (N_5482,N_4790,N_4260);
nor U5483 (N_5483,N_4913,N_4370);
and U5484 (N_5484,N_4600,N_4185);
nand U5485 (N_5485,N_4924,N_4113);
and U5486 (N_5486,N_4035,N_4127);
and U5487 (N_5487,N_4230,N_4487);
nand U5488 (N_5488,N_4507,N_4289);
or U5489 (N_5489,N_4889,N_4060);
nand U5490 (N_5490,N_4605,N_4204);
nand U5491 (N_5491,N_4994,N_4027);
or U5492 (N_5492,N_4736,N_4981);
nand U5493 (N_5493,N_4645,N_4298);
or U5494 (N_5494,N_4387,N_4785);
and U5495 (N_5495,N_4580,N_4156);
and U5496 (N_5496,N_4119,N_4363);
nand U5497 (N_5497,N_4588,N_4755);
nor U5498 (N_5498,N_4003,N_4358);
nand U5499 (N_5499,N_4400,N_4809);
nor U5500 (N_5500,N_4052,N_4251);
nand U5501 (N_5501,N_4913,N_4274);
nor U5502 (N_5502,N_4606,N_4265);
nor U5503 (N_5503,N_4425,N_4458);
and U5504 (N_5504,N_4889,N_4499);
or U5505 (N_5505,N_4502,N_4683);
nand U5506 (N_5506,N_4461,N_4359);
or U5507 (N_5507,N_4827,N_4917);
nor U5508 (N_5508,N_4854,N_4828);
or U5509 (N_5509,N_4426,N_4903);
nand U5510 (N_5510,N_4634,N_4812);
and U5511 (N_5511,N_4526,N_4750);
and U5512 (N_5512,N_4130,N_4594);
or U5513 (N_5513,N_4567,N_4815);
nand U5514 (N_5514,N_4939,N_4948);
and U5515 (N_5515,N_4730,N_4523);
nor U5516 (N_5516,N_4645,N_4127);
nand U5517 (N_5517,N_4032,N_4880);
nor U5518 (N_5518,N_4455,N_4437);
and U5519 (N_5519,N_4150,N_4206);
or U5520 (N_5520,N_4251,N_4867);
nand U5521 (N_5521,N_4783,N_4158);
nor U5522 (N_5522,N_4324,N_4917);
nand U5523 (N_5523,N_4379,N_4347);
nor U5524 (N_5524,N_4722,N_4006);
or U5525 (N_5525,N_4702,N_4014);
and U5526 (N_5526,N_4224,N_4778);
or U5527 (N_5527,N_4201,N_4067);
nand U5528 (N_5528,N_4548,N_4138);
nand U5529 (N_5529,N_4498,N_4877);
nor U5530 (N_5530,N_4110,N_4523);
and U5531 (N_5531,N_4296,N_4864);
nor U5532 (N_5532,N_4004,N_4837);
nor U5533 (N_5533,N_4314,N_4501);
nor U5534 (N_5534,N_4633,N_4828);
nor U5535 (N_5535,N_4030,N_4909);
and U5536 (N_5536,N_4950,N_4122);
and U5537 (N_5537,N_4636,N_4262);
or U5538 (N_5538,N_4175,N_4431);
nor U5539 (N_5539,N_4709,N_4941);
nor U5540 (N_5540,N_4720,N_4834);
and U5541 (N_5541,N_4978,N_4166);
or U5542 (N_5542,N_4985,N_4853);
or U5543 (N_5543,N_4968,N_4797);
nor U5544 (N_5544,N_4447,N_4644);
and U5545 (N_5545,N_4210,N_4406);
nand U5546 (N_5546,N_4026,N_4944);
nand U5547 (N_5547,N_4440,N_4024);
nor U5548 (N_5548,N_4830,N_4905);
nor U5549 (N_5549,N_4548,N_4715);
and U5550 (N_5550,N_4721,N_4983);
nand U5551 (N_5551,N_4508,N_4171);
and U5552 (N_5552,N_4077,N_4886);
or U5553 (N_5553,N_4337,N_4538);
and U5554 (N_5554,N_4012,N_4995);
nand U5555 (N_5555,N_4553,N_4386);
and U5556 (N_5556,N_4235,N_4267);
nand U5557 (N_5557,N_4699,N_4910);
or U5558 (N_5558,N_4262,N_4961);
nand U5559 (N_5559,N_4775,N_4048);
nor U5560 (N_5560,N_4003,N_4507);
or U5561 (N_5561,N_4076,N_4570);
nor U5562 (N_5562,N_4839,N_4214);
nor U5563 (N_5563,N_4640,N_4683);
and U5564 (N_5564,N_4817,N_4569);
or U5565 (N_5565,N_4519,N_4482);
or U5566 (N_5566,N_4974,N_4710);
or U5567 (N_5567,N_4548,N_4566);
nand U5568 (N_5568,N_4828,N_4852);
nor U5569 (N_5569,N_4469,N_4440);
and U5570 (N_5570,N_4254,N_4330);
or U5571 (N_5571,N_4940,N_4800);
or U5572 (N_5572,N_4707,N_4314);
nand U5573 (N_5573,N_4926,N_4228);
and U5574 (N_5574,N_4933,N_4400);
or U5575 (N_5575,N_4228,N_4690);
and U5576 (N_5576,N_4171,N_4825);
and U5577 (N_5577,N_4906,N_4692);
nor U5578 (N_5578,N_4508,N_4122);
or U5579 (N_5579,N_4892,N_4576);
nor U5580 (N_5580,N_4256,N_4775);
and U5581 (N_5581,N_4400,N_4492);
and U5582 (N_5582,N_4365,N_4809);
nor U5583 (N_5583,N_4838,N_4374);
nor U5584 (N_5584,N_4777,N_4436);
nand U5585 (N_5585,N_4356,N_4997);
nand U5586 (N_5586,N_4906,N_4664);
nor U5587 (N_5587,N_4752,N_4321);
nor U5588 (N_5588,N_4319,N_4793);
nand U5589 (N_5589,N_4420,N_4581);
nor U5590 (N_5590,N_4350,N_4008);
and U5591 (N_5591,N_4130,N_4042);
and U5592 (N_5592,N_4999,N_4051);
or U5593 (N_5593,N_4399,N_4159);
and U5594 (N_5594,N_4254,N_4312);
nor U5595 (N_5595,N_4190,N_4035);
nor U5596 (N_5596,N_4091,N_4128);
and U5597 (N_5597,N_4475,N_4220);
and U5598 (N_5598,N_4393,N_4445);
nand U5599 (N_5599,N_4440,N_4729);
and U5600 (N_5600,N_4314,N_4045);
nand U5601 (N_5601,N_4065,N_4090);
nor U5602 (N_5602,N_4968,N_4204);
or U5603 (N_5603,N_4026,N_4236);
and U5604 (N_5604,N_4010,N_4728);
and U5605 (N_5605,N_4926,N_4241);
and U5606 (N_5606,N_4403,N_4658);
nor U5607 (N_5607,N_4134,N_4035);
and U5608 (N_5608,N_4790,N_4646);
nor U5609 (N_5609,N_4735,N_4205);
and U5610 (N_5610,N_4073,N_4708);
or U5611 (N_5611,N_4483,N_4937);
nor U5612 (N_5612,N_4577,N_4630);
and U5613 (N_5613,N_4759,N_4860);
nand U5614 (N_5614,N_4768,N_4050);
or U5615 (N_5615,N_4485,N_4243);
nand U5616 (N_5616,N_4881,N_4841);
and U5617 (N_5617,N_4779,N_4543);
and U5618 (N_5618,N_4894,N_4289);
or U5619 (N_5619,N_4225,N_4330);
and U5620 (N_5620,N_4096,N_4650);
or U5621 (N_5621,N_4333,N_4814);
nand U5622 (N_5622,N_4341,N_4131);
and U5623 (N_5623,N_4154,N_4099);
nand U5624 (N_5624,N_4942,N_4247);
xor U5625 (N_5625,N_4148,N_4342);
or U5626 (N_5626,N_4185,N_4637);
and U5627 (N_5627,N_4085,N_4549);
xnor U5628 (N_5628,N_4417,N_4034);
nor U5629 (N_5629,N_4814,N_4084);
nand U5630 (N_5630,N_4783,N_4731);
and U5631 (N_5631,N_4598,N_4297);
nor U5632 (N_5632,N_4055,N_4972);
and U5633 (N_5633,N_4545,N_4500);
and U5634 (N_5634,N_4805,N_4079);
or U5635 (N_5635,N_4364,N_4554);
nand U5636 (N_5636,N_4033,N_4158);
nand U5637 (N_5637,N_4790,N_4807);
and U5638 (N_5638,N_4596,N_4447);
nor U5639 (N_5639,N_4764,N_4137);
nand U5640 (N_5640,N_4142,N_4571);
nand U5641 (N_5641,N_4114,N_4203);
nor U5642 (N_5642,N_4342,N_4763);
nand U5643 (N_5643,N_4532,N_4616);
nor U5644 (N_5644,N_4673,N_4605);
and U5645 (N_5645,N_4224,N_4937);
nand U5646 (N_5646,N_4143,N_4551);
nor U5647 (N_5647,N_4131,N_4543);
or U5648 (N_5648,N_4576,N_4014);
nor U5649 (N_5649,N_4063,N_4678);
or U5650 (N_5650,N_4444,N_4474);
nand U5651 (N_5651,N_4986,N_4291);
or U5652 (N_5652,N_4630,N_4642);
nor U5653 (N_5653,N_4014,N_4267);
nor U5654 (N_5654,N_4379,N_4969);
nand U5655 (N_5655,N_4192,N_4125);
nand U5656 (N_5656,N_4459,N_4008);
nor U5657 (N_5657,N_4486,N_4306);
nor U5658 (N_5658,N_4993,N_4897);
nand U5659 (N_5659,N_4435,N_4085);
or U5660 (N_5660,N_4551,N_4747);
and U5661 (N_5661,N_4940,N_4283);
or U5662 (N_5662,N_4380,N_4042);
or U5663 (N_5663,N_4160,N_4493);
nand U5664 (N_5664,N_4475,N_4068);
and U5665 (N_5665,N_4164,N_4924);
and U5666 (N_5666,N_4410,N_4108);
nor U5667 (N_5667,N_4756,N_4207);
nor U5668 (N_5668,N_4448,N_4735);
nor U5669 (N_5669,N_4284,N_4068);
xnor U5670 (N_5670,N_4459,N_4930);
nand U5671 (N_5671,N_4343,N_4205);
and U5672 (N_5672,N_4675,N_4824);
nor U5673 (N_5673,N_4921,N_4478);
and U5674 (N_5674,N_4909,N_4360);
and U5675 (N_5675,N_4655,N_4138);
nor U5676 (N_5676,N_4362,N_4878);
or U5677 (N_5677,N_4405,N_4942);
xor U5678 (N_5678,N_4453,N_4636);
nor U5679 (N_5679,N_4239,N_4875);
and U5680 (N_5680,N_4000,N_4987);
and U5681 (N_5681,N_4393,N_4020);
nand U5682 (N_5682,N_4754,N_4376);
and U5683 (N_5683,N_4977,N_4477);
nand U5684 (N_5684,N_4500,N_4774);
or U5685 (N_5685,N_4279,N_4855);
nand U5686 (N_5686,N_4256,N_4463);
nor U5687 (N_5687,N_4385,N_4665);
and U5688 (N_5688,N_4006,N_4099);
nor U5689 (N_5689,N_4108,N_4293);
nor U5690 (N_5690,N_4612,N_4305);
and U5691 (N_5691,N_4480,N_4467);
nor U5692 (N_5692,N_4311,N_4071);
and U5693 (N_5693,N_4220,N_4680);
nand U5694 (N_5694,N_4172,N_4807);
nor U5695 (N_5695,N_4408,N_4166);
nand U5696 (N_5696,N_4504,N_4770);
nand U5697 (N_5697,N_4308,N_4976);
and U5698 (N_5698,N_4441,N_4593);
and U5699 (N_5699,N_4091,N_4662);
or U5700 (N_5700,N_4442,N_4408);
nand U5701 (N_5701,N_4829,N_4749);
nor U5702 (N_5702,N_4131,N_4468);
and U5703 (N_5703,N_4396,N_4846);
or U5704 (N_5704,N_4065,N_4159);
or U5705 (N_5705,N_4924,N_4822);
and U5706 (N_5706,N_4651,N_4081);
or U5707 (N_5707,N_4166,N_4781);
or U5708 (N_5708,N_4076,N_4243);
and U5709 (N_5709,N_4116,N_4681);
nor U5710 (N_5710,N_4955,N_4457);
or U5711 (N_5711,N_4956,N_4409);
nand U5712 (N_5712,N_4835,N_4002);
nand U5713 (N_5713,N_4823,N_4959);
and U5714 (N_5714,N_4452,N_4897);
nand U5715 (N_5715,N_4519,N_4776);
nor U5716 (N_5716,N_4573,N_4193);
nor U5717 (N_5717,N_4124,N_4967);
nor U5718 (N_5718,N_4867,N_4320);
nor U5719 (N_5719,N_4192,N_4808);
nand U5720 (N_5720,N_4086,N_4540);
or U5721 (N_5721,N_4212,N_4123);
nor U5722 (N_5722,N_4221,N_4710);
xnor U5723 (N_5723,N_4837,N_4646);
nand U5724 (N_5724,N_4293,N_4093);
and U5725 (N_5725,N_4316,N_4729);
nor U5726 (N_5726,N_4881,N_4619);
or U5727 (N_5727,N_4847,N_4853);
and U5728 (N_5728,N_4104,N_4002);
and U5729 (N_5729,N_4627,N_4688);
and U5730 (N_5730,N_4747,N_4764);
or U5731 (N_5731,N_4692,N_4618);
nand U5732 (N_5732,N_4847,N_4277);
nand U5733 (N_5733,N_4140,N_4764);
nor U5734 (N_5734,N_4136,N_4389);
or U5735 (N_5735,N_4118,N_4490);
or U5736 (N_5736,N_4318,N_4565);
and U5737 (N_5737,N_4439,N_4969);
or U5738 (N_5738,N_4364,N_4570);
nand U5739 (N_5739,N_4028,N_4730);
or U5740 (N_5740,N_4669,N_4849);
or U5741 (N_5741,N_4411,N_4339);
or U5742 (N_5742,N_4298,N_4847);
nand U5743 (N_5743,N_4843,N_4083);
or U5744 (N_5744,N_4890,N_4406);
or U5745 (N_5745,N_4376,N_4149);
or U5746 (N_5746,N_4722,N_4591);
nor U5747 (N_5747,N_4839,N_4602);
nor U5748 (N_5748,N_4806,N_4898);
nor U5749 (N_5749,N_4338,N_4524);
xor U5750 (N_5750,N_4889,N_4075);
or U5751 (N_5751,N_4180,N_4706);
nand U5752 (N_5752,N_4382,N_4590);
and U5753 (N_5753,N_4925,N_4153);
and U5754 (N_5754,N_4274,N_4012);
nor U5755 (N_5755,N_4010,N_4357);
or U5756 (N_5756,N_4721,N_4580);
nand U5757 (N_5757,N_4890,N_4515);
nor U5758 (N_5758,N_4727,N_4389);
nor U5759 (N_5759,N_4051,N_4217);
and U5760 (N_5760,N_4227,N_4057);
or U5761 (N_5761,N_4164,N_4236);
or U5762 (N_5762,N_4419,N_4646);
nor U5763 (N_5763,N_4177,N_4214);
nor U5764 (N_5764,N_4968,N_4852);
and U5765 (N_5765,N_4406,N_4097);
xor U5766 (N_5766,N_4587,N_4248);
and U5767 (N_5767,N_4302,N_4245);
nand U5768 (N_5768,N_4240,N_4708);
and U5769 (N_5769,N_4967,N_4677);
nor U5770 (N_5770,N_4835,N_4191);
nand U5771 (N_5771,N_4714,N_4880);
or U5772 (N_5772,N_4281,N_4719);
or U5773 (N_5773,N_4824,N_4365);
or U5774 (N_5774,N_4892,N_4197);
and U5775 (N_5775,N_4448,N_4087);
or U5776 (N_5776,N_4100,N_4905);
nor U5777 (N_5777,N_4186,N_4887);
nor U5778 (N_5778,N_4651,N_4203);
or U5779 (N_5779,N_4489,N_4257);
or U5780 (N_5780,N_4847,N_4944);
nand U5781 (N_5781,N_4780,N_4207);
nor U5782 (N_5782,N_4275,N_4962);
and U5783 (N_5783,N_4201,N_4379);
or U5784 (N_5784,N_4774,N_4115);
and U5785 (N_5785,N_4421,N_4977);
nand U5786 (N_5786,N_4931,N_4540);
nand U5787 (N_5787,N_4344,N_4691);
and U5788 (N_5788,N_4069,N_4930);
nor U5789 (N_5789,N_4207,N_4502);
or U5790 (N_5790,N_4050,N_4667);
and U5791 (N_5791,N_4277,N_4807);
nand U5792 (N_5792,N_4603,N_4958);
xor U5793 (N_5793,N_4618,N_4012);
and U5794 (N_5794,N_4191,N_4351);
and U5795 (N_5795,N_4489,N_4919);
or U5796 (N_5796,N_4815,N_4580);
nand U5797 (N_5797,N_4475,N_4714);
or U5798 (N_5798,N_4547,N_4778);
and U5799 (N_5799,N_4475,N_4804);
or U5800 (N_5800,N_4492,N_4577);
nand U5801 (N_5801,N_4992,N_4054);
or U5802 (N_5802,N_4204,N_4109);
or U5803 (N_5803,N_4796,N_4480);
nor U5804 (N_5804,N_4166,N_4357);
or U5805 (N_5805,N_4119,N_4082);
and U5806 (N_5806,N_4959,N_4354);
and U5807 (N_5807,N_4535,N_4197);
or U5808 (N_5808,N_4809,N_4441);
nand U5809 (N_5809,N_4014,N_4603);
nor U5810 (N_5810,N_4497,N_4257);
or U5811 (N_5811,N_4410,N_4298);
or U5812 (N_5812,N_4744,N_4164);
nand U5813 (N_5813,N_4598,N_4795);
nor U5814 (N_5814,N_4781,N_4078);
or U5815 (N_5815,N_4687,N_4135);
nor U5816 (N_5816,N_4194,N_4664);
nor U5817 (N_5817,N_4851,N_4442);
and U5818 (N_5818,N_4600,N_4576);
nand U5819 (N_5819,N_4374,N_4448);
or U5820 (N_5820,N_4826,N_4961);
or U5821 (N_5821,N_4341,N_4477);
and U5822 (N_5822,N_4308,N_4376);
nor U5823 (N_5823,N_4710,N_4107);
and U5824 (N_5824,N_4356,N_4368);
nand U5825 (N_5825,N_4137,N_4464);
nand U5826 (N_5826,N_4474,N_4460);
nand U5827 (N_5827,N_4534,N_4178);
and U5828 (N_5828,N_4451,N_4950);
nor U5829 (N_5829,N_4057,N_4848);
nor U5830 (N_5830,N_4244,N_4531);
nand U5831 (N_5831,N_4769,N_4036);
and U5832 (N_5832,N_4478,N_4370);
and U5833 (N_5833,N_4967,N_4931);
nor U5834 (N_5834,N_4091,N_4594);
nand U5835 (N_5835,N_4467,N_4071);
or U5836 (N_5836,N_4330,N_4272);
or U5837 (N_5837,N_4505,N_4677);
xor U5838 (N_5838,N_4681,N_4837);
nand U5839 (N_5839,N_4010,N_4560);
or U5840 (N_5840,N_4617,N_4243);
nor U5841 (N_5841,N_4960,N_4351);
and U5842 (N_5842,N_4858,N_4365);
nor U5843 (N_5843,N_4064,N_4283);
or U5844 (N_5844,N_4487,N_4133);
or U5845 (N_5845,N_4723,N_4663);
and U5846 (N_5846,N_4217,N_4305);
nor U5847 (N_5847,N_4973,N_4942);
nand U5848 (N_5848,N_4262,N_4980);
nand U5849 (N_5849,N_4842,N_4864);
and U5850 (N_5850,N_4145,N_4973);
or U5851 (N_5851,N_4139,N_4061);
or U5852 (N_5852,N_4203,N_4770);
and U5853 (N_5853,N_4704,N_4668);
nor U5854 (N_5854,N_4304,N_4496);
or U5855 (N_5855,N_4638,N_4743);
and U5856 (N_5856,N_4743,N_4300);
or U5857 (N_5857,N_4554,N_4424);
nor U5858 (N_5858,N_4303,N_4610);
nor U5859 (N_5859,N_4225,N_4985);
and U5860 (N_5860,N_4227,N_4112);
nand U5861 (N_5861,N_4955,N_4694);
nand U5862 (N_5862,N_4641,N_4681);
nor U5863 (N_5863,N_4918,N_4697);
nor U5864 (N_5864,N_4667,N_4264);
nor U5865 (N_5865,N_4664,N_4492);
or U5866 (N_5866,N_4626,N_4971);
nor U5867 (N_5867,N_4053,N_4311);
nor U5868 (N_5868,N_4501,N_4518);
or U5869 (N_5869,N_4534,N_4474);
nor U5870 (N_5870,N_4926,N_4110);
or U5871 (N_5871,N_4993,N_4838);
xnor U5872 (N_5872,N_4978,N_4046);
nand U5873 (N_5873,N_4533,N_4539);
nand U5874 (N_5874,N_4747,N_4984);
nor U5875 (N_5875,N_4646,N_4061);
or U5876 (N_5876,N_4087,N_4300);
nand U5877 (N_5877,N_4836,N_4173);
nand U5878 (N_5878,N_4981,N_4829);
or U5879 (N_5879,N_4583,N_4362);
or U5880 (N_5880,N_4095,N_4492);
and U5881 (N_5881,N_4795,N_4182);
or U5882 (N_5882,N_4187,N_4692);
nor U5883 (N_5883,N_4567,N_4532);
or U5884 (N_5884,N_4870,N_4335);
nand U5885 (N_5885,N_4812,N_4431);
and U5886 (N_5886,N_4131,N_4937);
xor U5887 (N_5887,N_4037,N_4958);
and U5888 (N_5888,N_4451,N_4084);
nor U5889 (N_5889,N_4756,N_4808);
nor U5890 (N_5890,N_4683,N_4671);
or U5891 (N_5891,N_4798,N_4058);
or U5892 (N_5892,N_4069,N_4285);
or U5893 (N_5893,N_4711,N_4814);
or U5894 (N_5894,N_4604,N_4034);
or U5895 (N_5895,N_4019,N_4433);
or U5896 (N_5896,N_4497,N_4139);
nor U5897 (N_5897,N_4098,N_4875);
or U5898 (N_5898,N_4911,N_4292);
and U5899 (N_5899,N_4364,N_4564);
nor U5900 (N_5900,N_4544,N_4515);
nand U5901 (N_5901,N_4676,N_4812);
or U5902 (N_5902,N_4071,N_4049);
nand U5903 (N_5903,N_4956,N_4123);
nor U5904 (N_5904,N_4940,N_4996);
xor U5905 (N_5905,N_4023,N_4051);
nand U5906 (N_5906,N_4305,N_4838);
nand U5907 (N_5907,N_4443,N_4154);
nand U5908 (N_5908,N_4813,N_4560);
nand U5909 (N_5909,N_4044,N_4096);
nor U5910 (N_5910,N_4495,N_4527);
nor U5911 (N_5911,N_4810,N_4151);
or U5912 (N_5912,N_4033,N_4679);
nor U5913 (N_5913,N_4089,N_4889);
or U5914 (N_5914,N_4609,N_4556);
nand U5915 (N_5915,N_4960,N_4879);
and U5916 (N_5916,N_4641,N_4217);
or U5917 (N_5917,N_4212,N_4094);
nand U5918 (N_5918,N_4654,N_4013);
or U5919 (N_5919,N_4770,N_4516);
nor U5920 (N_5920,N_4386,N_4987);
nor U5921 (N_5921,N_4784,N_4942);
nand U5922 (N_5922,N_4253,N_4476);
nand U5923 (N_5923,N_4563,N_4643);
or U5924 (N_5924,N_4012,N_4201);
nand U5925 (N_5925,N_4501,N_4276);
nor U5926 (N_5926,N_4088,N_4601);
or U5927 (N_5927,N_4203,N_4789);
and U5928 (N_5928,N_4617,N_4335);
and U5929 (N_5929,N_4603,N_4474);
nor U5930 (N_5930,N_4847,N_4275);
or U5931 (N_5931,N_4002,N_4937);
and U5932 (N_5932,N_4762,N_4738);
nor U5933 (N_5933,N_4967,N_4137);
and U5934 (N_5934,N_4241,N_4216);
nand U5935 (N_5935,N_4796,N_4560);
nor U5936 (N_5936,N_4348,N_4893);
and U5937 (N_5937,N_4449,N_4943);
nand U5938 (N_5938,N_4974,N_4499);
and U5939 (N_5939,N_4650,N_4300);
or U5940 (N_5940,N_4920,N_4104);
nand U5941 (N_5941,N_4951,N_4888);
nand U5942 (N_5942,N_4008,N_4799);
and U5943 (N_5943,N_4408,N_4848);
nor U5944 (N_5944,N_4679,N_4260);
nor U5945 (N_5945,N_4024,N_4556);
or U5946 (N_5946,N_4424,N_4950);
or U5947 (N_5947,N_4659,N_4663);
nor U5948 (N_5948,N_4999,N_4854);
nand U5949 (N_5949,N_4823,N_4976);
nor U5950 (N_5950,N_4290,N_4376);
nand U5951 (N_5951,N_4332,N_4344);
or U5952 (N_5952,N_4740,N_4147);
or U5953 (N_5953,N_4091,N_4210);
xnor U5954 (N_5954,N_4476,N_4478);
nor U5955 (N_5955,N_4997,N_4399);
nor U5956 (N_5956,N_4720,N_4008);
nand U5957 (N_5957,N_4525,N_4863);
or U5958 (N_5958,N_4186,N_4346);
and U5959 (N_5959,N_4720,N_4007);
nand U5960 (N_5960,N_4095,N_4909);
or U5961 (N_5961,N_4080,N_4202);
nor U5962 (N_5962,N_4073,N_4535);
nor U5963 (N_5963,N_4484,N_4875);
and U5964 (N_5964,N_4137,N_4419);
and U5965 (N_5965,N_4140,N_4731);
nor U5966 (N_5966,N_4275,N_4631);
or U5967 (N_5967,N_4171,N_4120);
nor U5968 (N_5968,N_4297,N_4410);
nand U5969 (N_5969,N_4504,N_4902);
and U5970 (N_5970,N_4299,N_4166);
nor U5971 (N_5971,N_4195,N_4632);
and U5972 (N_5972,N_4473,N_4278);
nand U5973 (N_5973,N_4174,N_4326);
or U5974 (N_5974,N_4337,N_4777);
nand U5975 (N_5975,N_4679,N_4693);
nand U5976 (N_5976,N_4595,N_4415);
or U5977 (N_5977,N_4750,N_4539);
or U5978 (N_5978,N_4276,N_4825);
nor U5979 (N_5979,N_4847,N_4522);
nor U5980 (N_5980,N_4380,N_4890);
nand U5981 (N_5981,N_4304,N_4266);
nand U5982 (N_5982,N_4665,N_4939);
and U5983 (N_5983,N_4357,N_4275);
and U5984 (N_5984,N_4299,N_4205);
or U5985 (N_5985,N_4969,N_4437);
nand U5986 (N_5986,N_4585,N_4180);
nor U5987 (N_5987,N_4645,N_4895);
nand U5988 (N_5988,N_4753,N_4550);
or U5989 (N_5989,N_4985,N_4003);
and U5990 (N_5990,N_4121,N_4462);
nand U5991 (N_5991,N_4046,N_4210);
nand U5992 (N_5992,N_4199,N_4960);
nand U5993 (N_5993,N_4834,N_4605);
or U5994 (N_5994,N_4308,N_4853);
or U5995 (N_5995,N_4554,N_4482);
nor U5996 (N_5996,N_4063,N_4446);
or U5997 (N_5997,N_4383,N_4627);
and U5998 (N_5998,N_4609,N_4608);
or U5999 (N_5999,N_4351,N_4345);
nor U6000 (N_6000,N_5756,N_5541);
or U6001 (N_6001,N_5392,N_5795);
nand U6002 (N_6002,N_5087,N_5474);
and U6003 (N_6003,N_5202,N_5394);
or U6004 (N_6004,N_5857,N_5010);
nand U6005 (N_6005,N_5567,N_5179);
nor U6006 (N_6006,N_5557,N_5686);
and U6007 (N_6007,N_5965,N_5054);
nand U6008 (N_6008,N_5661,N_5806);
nor U6009 (N_6009,N_5414,N_5442);
and U6010 (N_6010,N_5568,N_5552);
nor U6011 (N_6011,N_5006,N_5055);
nor U6012 (N_6012,N_5307,N_5116);
nor U6013 (N_6013,N_5781,N_5282);
and U6014 (N_6014,N_5449,N_5141);
or U6015 (N_6015,N_5764,N_5165);
and U6016 (N_6016,N_5953,N_5652);
nand U6017 (N_6017,N_5802,N_5124);
and U6018 (N_6018,N_5289,N_5025);
and U6019 (N_6019,N_5709,N_5695);
and U6020 (N_6020,N_5560,N_5934);
nand U6021 (N_6021,N_5177,N_5245);
and U6022 (N_6022,N_5901,N_5873);
nand U6023 (N_6023,N_5765,N_5311);
nand U6024 (N_6024,N_5822,N_5098);
nor U6025 (N_6025,N_5396,N_5489);
and U6026 (N_6026,N_5349,N_5636);
nand U6027 (N_6027,N_5607,N_5785);
nor U6028 (N_6028,N_5689,N_5227);
nand U6029 (N_6029,N_5915,N_5947);
and U6030 (N_6030,N_5342,N_5451);
nand U6031 (N_6031,N_5883,N_5382);
and U6032 (N_6032,N_5432,N_5330);
or U6033 (N_6033,N_5621,N_5559);
or U6034 (N_6034,N_5160,N_5036);
and U6035 (N_6035,N_5800,N_5155);
nand U6036 (N_6036,N_5164,N_5103);
nor U6037 (N_6037,N_5867,N_5536);
or U6038 (N_6038,N_5108,N_5153);
nor U6039 (N_6039,N_5618,N_5970);
nand U6040 (N_6040,N_5790,N_5954);
and U6041 (N_6041,N_5705,N_5121);
and U6042 (N_6042,N_5602,N_5412);
nor U6043 (N_6043,N_5902,N_5539);
nand U6044 (N_6044,N_5452,N_5679);
and U6045 (N_6045,N_5182,N_5273);
or U6046 (N_6046,N_5700,N_5562);
and U6047 (N_6047,N_5018,N_5550);
or U6048 (N_6048,N_5105,N_5584);
nand U6049 (N_6049,N_5738,N_5810);
nand U6050 (N_6050,N_5749,N_5453);
or U6051 (N_6051,N_5657,N_5356);
and U6052 (N_6052,N_5587,N_5376);
nor U6053 (N_6053,N_5250,N_5920);
nand U6054 (N_6054,N_5511,N_5032);
and U6055 (N_6055,N_5737,N_5157);
or U6056 (N_6056,N_5077,N_5713);
or U6057 (N_6057,N_5670,N_5029);
nand U6058 (N_6058,N_5281,N_5234);
and U6059 (N_6059,N_5870,N_5385);
nand U6060 (N_6060,N_5880,N_5325);
or U6061 (N_6061,N_5174,N_5007);
nand U6062 (N_6062,N_5861,N_5564);
and U6063 (N_6063,N_5850,N_5506);
nand U6064 (N_6064,N_5491,N_5251);
nor U6065 (N_6065,N_5329,N_5669);
nor U6066 (N_6066,N_5122,N_5910);
nor U6067 (N_6067,N_5386,N_5338);
nand U6068 (N_6068,N_5823,N_5192);
nand U6069 (N_6069,N_5914,N_5668);
and U6070 (N_6070,N_5359,N_5379);
or U6071 (N_6071,N_5095,N_5928);
and U6072 (N_6072,N_5983,N_5466);
nand U6073 (N_6073,N_5093,N_5891);
nand U6074 (N_6074,N_5257,N_5839);
nor U6075 (N_6075,N_5316,N_5014);
nand U6076 (N_6076,N_5882,N_5404);
nor U6077 (N_6077,N_5242,N_5369);
nand U6078 (N_6078,N_5752,N_5318);
or U6079 (N_6079,N_5285,N_5012);
nor U6080 (N_6080,N_5183,N_5892);
nand U6081 (N_6081,N_5859,N_5588);
or U6082 (N_6082,N_5648,N_5403);
nand U6083 (N_6083,N_5254,N_5677);
nand U6084 (N_6084,N_5745,N_5156);
nor U6085 (N_6085,N_5894,N_5678);
and U6086 (N_6086,N_5258,N_5389);
or U6087 (N_6087,N_5381,N_5181);
nand U6088 (N_6088,N_5016,N_5310);
or U6089 (N_6089,N_5935,N_5692);
xnor U6090 (N_6090,N_5555,N_5889);
nand U6091 (N_6091,N_5653,N_5704);
or U6092 (N_6092,N_5465,N_5331);
or U6093 (N_6093,N_5175,N_5685);
nand U6094 (N_6094,N_5081,N_5730);
or U6095 (N_6095,N_5924,N_5593);
and U6096 (N_6096,N_5523,N_5145);
or U6097 (N_6097,N_5461,N_5266);
and U6098 (N_6098,N_5305,N_5723);
or U6099 (N_6099,N_5803,N_5278);
or U6100 (N_6100,N_5957,N_5626);
nand U6101 (N_6101,N_5586,N_5643);
and U6102 (N_6102,N_5230,N_5645);
nor U6103 (N_6103,N_5968,N_5913);
or U6104 (N_6104,N_5650,N_5042);
and U6105 (N_6105,N_5972,N_5372);
nor U6106 (N_6106,N_5346,N_5774);
nor U6107 (N_6107,N_5527,N_5193);
nand U6108 (N_6108,N_5480,N_5200);
and U6109 (N_6109,N_5946,N_5110);
or U6110 (N_6110,N_5345,N_5878);
or U6111 (N_6111,N_5438,N_5231);
and U6112 (N_6112,N_5868,N_5874);
nand U6113 (N_6113,N_5654,N_5428);
and U6114 (N_6114,N_5931,N_5722);
or U6115 (N_6115,N_5485,N_5547);
nand U6116 (N_6116,N_5464,N_5732);
nand U6117 (N_6117,N_5092,N_5350);
or U6118 (N_6118,N_5300,N_5472);
or U6119 (N_6119,N_5005,N_5641);
or U6120 (N_6120,N_5760,N_5622);
nand U6121 (N_6121,N_5731,N_5630);
nor U6122 (N_6122,N_5952,N_5696);
and U6123 (N_6123,N_5225,N_5979);
nor U6124 (N_6124,N_5963,N_5221);
or U6125 (N_6125,N_5191,N_5013);
or U6126 (N_6126,N_5462,N_5406);
or U6127 (N_6127,N_5071,N_5573);
nor U6128 (N_6128,N_5027,N_5797);
or U6129 (N_6129,N_5097,N_5792);
nor U6130 (N_6130,N_5773,N_5306);
nand U6131 (N_6131,N_5493,N_5619);
and U6132 (N_6132,N_5603,N_5646);
nor U6133 (N_6133,N_5017,N_5690);
nor U6134 (N_6134,N_5180,N_5053);
or U6135 (N_6135,N_5409,N_5158);
or U6136 (N_6136,N_5875,N_5624);
nand U6137 (N_6137,N_5344,N_5682);
nand U6138 (N_6138,N_5966,N_5906);
nand U6139 (N_6139,N_5353,N_5606);
nand U6140 (N_6140,N_5767,N_5707);
or U6141 (N_6141,N_5577,N_5959);
nor U6142 (N_6142,N_5333,N_5829);
or U6143 (N_6143,N_5268,N_5496);
and U6144 (N_6144,N_5267,N_5127);
nor U6145 (N_6145,N_5783,N_5111);
nand U6146 (N_6146,N_5131,N_5213);
nand U6147 (N_6147,N_5253,N_5069);
nor U6148 (N_6148,N_5549,N_5526);
and U6149 (N_6149,N_5241,N_5943);
nand U6150 (N_6150,N_5799,N_5150);
and U6151 (N_6151,N_5067,N_5048);
or U6152 (N_6152,N_5877,N_5498);
nand U6153 (N_6153,N_5178,N_5524);
and U6154 (N_6154,N_5317,N_5287);
nand U6155 (N_6155,N_5494,N_5635);
nand U6156 (N_6156,N_5687,N_5410);
nand U6157 (N_6157,N_5303,N_5084);
or U6158 (N_6158,N_5236,N_5594);
or U6159 (N_6159,N_5352,N_5746);
nand U6160 (N_6160,N_5063,N_5964);
and U6161 (N_6161,N_5365,N_5189);
nor U6162 (N_6162,N_5589,N_5431);
nand U6163 (N_6163,N_5008,N_5985);
xor U6164 (N_6164,N_5206,N_5529);
nand U6165 (N_6165,N_5222,N_5497);
or U6166 (N_6166,N_5437,N_5060);
nand U6167 (N_6167,N_5426,N_5154);
nand U6168 (N_6168,N_5582,N_5681);
nor U6169 (N_6169,N_5517,N_5443);
nand U6170 (N_6170,N_5988,N_5520);
nor U6171 (N_6171,N_5816,N_5120);
nor U6172 (N_6172,N_5632,N_5417);
nand U6173 (N_6173,N_5446,N_5610);
nand U6174 (N_6174,N_5512,N_5041);
nor U6175 (N_6175,N_5718,N_5265);
nor U6176 (N_6176,N_5051,N_5728);
nand U6177 (N_6177,N_5215,N_5644);
nand U6178 (N_6178,N_5291,N_5845);
and U6179 (N_6179,N_5929,N_5400);
and U6180 (N_6180,N_5831,N_5667);
and U6181 (N_6181,N_5421,N_5444);
nor U6182 (N_6182,N_5134,N_5038);
xor U6183 (N_6183,N_5383,N_5739);
and U6184 (N_6184,N_5384,N_5298);
and U6185 (N_6185,N_5827,N_5735);
or U6186 (N_6186,N_5411,N_5272);
nand U6187 (N_6187,N_5605,N_5777);
nand U6188 (N_6188,N_5515,N_5940);
and U6189 (N_6189,N_5944,N_5364);
or U6190 (N_6190,N_5469,N_5509);
nor U6191 (N_6191,N_5960,N_5532);
nand U6192 (N_6192,N_5712,N_5118);
and U6193 (N_6193,N_5601,N_5371);
or U6194 (N_6194,N_5537,N_5917);
and U6195 (N_6195,N_5322,N_5842);
and U6196 (N_6196,N_5275,N_5862);
nor U6197 (N_6197,N_5355,N_5470);
and U6198 (N_6198,N_5212,N_5837);
nand U6199 (N_6199,N_5424,N_5378);
or U6200 (N_6200,N_5495,N_5533);
nor U6201 (N_6201,N_5980,N_5327);
or U6202 (N_6202,N_5675,N_5613);
or U6203 (N_6203,N_5763,N_5834);
or U6204 (N_6204,N_5255,N_5633);
and U6205 (N_6205,N_5339,N_5659);
and U6206 (N_6206,N_5720,N_5858);
and U6207 (N_6207,N_5534,N_5982);
or U6208 (N_6208,N_5741,N_5194);
and U6209 (N_6209,N_5321,N_5228);
or U6210 (N_6210,N_5721,N_5436);
nand U6211 (N_6211,N_5904,N_5569);
nor U6212 (N_6212,N_5173,N_5820);
and U6213 (N_6213,N_5548,N_5370);
nor U6214 (N_6214,N_5059,N_5297);
and U6215 (N_6215,N_5185,N_5091);
nand U6216 (N_6216,N_5912,N_5725);
nand U6217 (N_6217,N_5544,N_5079);
and U6218 (N_6218,N_5240,N_5142);
and U6219 (N_6219,N_5471,N_5864);
and U6220 (N_6220,N_5684,N_5841);
nand U6221 (N_6221,N_5948,N_5719);
and U6222 (N_6222,N_5479,N_5631);
nor U6223 (N_6223,N_5490,N_5237);
and U6224 (N_6224,N_5101,N_5791);
nand U6225 (N_6225,N_5759,N_5172);
nor U6226 (N_6226,N_5843,N_5138);
or U6227 (N_6227,N_5224,N_5301);
and U6228 (N_6228,N_5701,N_5057);
and U6229 (N_6229,N_5852,N_5244);
nand U6230 (N_6230,N_5280,N_5269);
nand U6231 (N_6231,N_5402,N_5768);
and U6232 (N_6232,N_5430,N_5152);
or U6233 (N_6233,N_5276,N_5796);
nand U6234 (N_6234,N_5037,N_5778);
nor U6235 (N_6235,N_5500,N_5604);
or U6236 (N_6236,N_5736,N_5000);
or U6237 (N_6237,N_5047,N_5503);
nand U6238 (N_6238,N_5727,N_5513);
and U6239 (N_6239,N_5293,N_5617);
or U6240 (N_6240,N_5933,N_5439);
nor U6241 (N_6241,N_5981,N_5542);
or U6242 (N_6242,N_5387,N_5058);
or U6243 (N_6243,N_5805,N_5238);
and U6244 (N_6244,N_5832,N_5075);
nor U6245 (N_6245,N_5450,N_5425);
or U6246 (N_6246,N_5994,N_5961);
nand U6247 (N_6247,N_5885,N_5769);
nand U6248 (N_6248,N_5459,N_5990);
or U6249 (N_6249,N_5754,N_5572);
and U6250 (N_6250,N_5854,N_5726);
nand U6251 (N_6251,N_5220,N_5969);
nand U6252 (N_6252,N_5197,N_5232);
and U6253 (N_6253,N_5551,N_5112);
nand U6254 (N_6254,N_5585,N_5226);
and U6255 (N_6255,N_5697,N_5698);
and U6256 (N_6256,N_5922,N_5186);
nand U6257 (N_6257,N_5518,N_5104);
or U6258 (N_6258,N_5936,N_5395);
or U6259 (N_6259,N_5419,N_5418);
nor U6260 (N_6260,N_5066,N_5997);
and U6261 (N_6261,N_5872,N_5591);
nor U6262 (N_6262,N_5137,N_5256);
and U6263 (N_6263,N_5210,N_5085);
and U6264 (N_6264,N_5729,N_5611);
or U6265 (N_6265,N_5218,N_5088);
nor U6266 (N_6266,N_5407,N_5072);
nor U6267 (N_6267,N_5897,N_5993);
and U6268 (N_6268,N_5538,N_5065);
and U6269 (N_6269,N_5888,N_5162);
or U6270 (N_6270,N_5710,N_5184);
and U6271 (N_6271,N_5949,N_5628);
nor U6272 (N_6272,N_5853,N_5900);
and U6273 (N_6273,N_5627,N_5592);
nand U6274 (N_6274,N_5740,N_5814);
nor U6275 (N_6275,N_5879,N_5235);
nand U6276 (N_6276,N_5286,N_5660);
or U6277 (N_6277,N_5296,N_5742);
nor U6278 (N_6278,N_5958,N_5304);
and U6279 (N_6279,N_5457,N_5898);
nand U6280 (N_6280,N_5579,N_5114);
nand U6281 (N_6281,N_5094,N_5565);
nand U6282 (N_6282,N_5324,N_5638);
nor U6283 (N_6283,N_5161,N_5784);
and U6284 (N_6284,N_5043,N_5671);
nand U6285 (N_6285,N_5895,N_5986);
nor U6286 (N_6286,N_5999,N_5107);
nand U6287 (N_6287,N_5168,N_5283);
and U6288 (N_6288,N_5855,N_5445);
nor U6289 (N_6289,N_5460,N_5334);
or U6290 (N_6290,N_5119,N_5320);
or U6291 (N_6291,N_5477,N_5502);
nor U6292 (N_6292,N_5649,N_5919);
or U6293 (N_6293,N_5019,N_5945);
nor U6294 (N_6294,N_5195,N_5708);
and U6295 (N_6295,N_5312,N_5824);
or U6296 (N_6296,N_5420,N_5612);
or U6297 (N_6297,N_5393,N_5751);
nor U6298 (N_6298,N_5347,N_5575);
nor U6299 (N_6299,N_5308,N_5505);
and U6300 (N_6300,N_5003,N_5563);
nor U6301 (N_6301,N_5198,N_5614);
nor U6302 (N_6302,N_5416,N_5380);
nand U6303 (N_6303,N_5249,N_5423);
nor U6304 (N_6304,N_5399,N_5580);
nor U6305 (N_6305,N_5033,N_5779);
or U6306 (N_6306,N_5989,N_5620);
nand U6307 (N_6307,N_5836,N_5776);
and U6308 (N_6308,N_5361,N_5911);
nor U6309 (N_6309,N_5336,N_5061);
or U6310 (N_6310,N_5656,N_5804);
and U6311 (N_6311,N_5714,N_5642);
and U6312 (N_6312,N_5941,N_5292);
nand U6313 (N_6313,N_5117,N_5052);
nand U6314 (N_6314,N_5833,N_5204);
nand U6315 (N_6315,N_5757,N_5531);
nand U6316 (N_6316,N_5899,N_5408);
nand U6317 (N_6317,N_5514,N_5651);
nand U6318 (N_6318,N_5772,N_5045);
nand U6319 (N_6319,N_5973,N_5358);
and U6320 (N_6320,N_5570,N_5821);
or U6321 (N_6321,N_5488,N_5566);
and U6322 (N_6322,N_5089,N_5926);
and U6323 (N_6323,N_5733,N_5113);
or U6324 (N_6324,N_5024,N_5170);
and U6325 (N_6325,N_5148,N_5397);
nand U6326 (N_6326,N_5844,N_5561);
or U6327 (N_6327,N_5373,N_5484);
or U6328 (N_6328,N_5354,N_5476);
nand U6329 (N_6329,N_5664,N_5553);
or U6330 (N_6330,N_5299,N_5367);
nand U6331 (N_6331,N_5332,N_5277);
or U6332 (N_6332,N_5998,N_5263);
or U6333 (N_6333,N_5674,N_5683);
or U6334 (N_6334,N_5893,N_5467);
nand U6335 (N_6335,N_5747,N_5374);
nor U6336 (N_6336,N_5753,N_5615);
and U6337 (N_6337,N_5481,N_5597);
nor U6338 (N_6338,N_5096,N_5448);
and U6339 (N_6339,N_5216,N_5422);
or U6340 (N_6340,N_5835,N_5942);
and U6341 (N_6341,N_5992,N_5319);
nor U6342 (N_6342,N_5521,N_5454);
or U6343 (N_6343,N_5413,N_5229);
nor U6344 (N_6344,N_5673,N_5483);
and U6345 (N_6345,N_5039,N_5716);
and U6346 (N_6346,N_5554,N_5083);
or U6347 (N_6347,N_5159,N_5596);
nand U6348 (N_6348,N_5128,N_5004);
nand U6349 (N_6349,N_5270,N_5530);
and U6350 (N_6350,N_5717,N_5264);
or U6351 (N_6351,N_5151,N_5830);
and U6352 (N_6352,N_5658,N_5815);
or U6353 (N_6353,N_5343,N_5188);
or U6354 (N_6354,N_5932,N_5074);
nor U6355 (N_6355,N_5907,N_5026);
and U6356 (N_6356,N_5288,N_5456);
nor U6357 (N_6357,N_5595,N_5434);
and U6358 (N_6358,N_5743,N_5702);
and U6359 (N_6359,N_5558,N_5508);
nor U6360 (N_6360,N_5223,N_5528);
nand U6361 (N_6361,N_5629,N_5616);
or U6362 (N_6362,N_5851,N_5543);
or U6363 (N_6363,N_5556,N_5099);
and U6364 (N_6364,N_5724,N_5261);
and U6365 (N_6365,N_5140,N_5368);
and U6366 (N_6366,N_5762,N_5205);
nand U6367 (N_6367,N_5391,N_5540);
nand U6368 (N_6368,N_5046,N_5987);
nor U6369 (N_6369,N_5028,N_5187);
and U6370 (N_6370,N_5598,N_5035);
nor U6371 (N_6371,N_5313,N_5734);
nor U6372 (N_6372,N_5259,N_5499);
or U6373 (N_6373,N_5123,N_5758);
nor U6374 (N_6374,N_5786,N_5706);
nand U6375 (N_6375,N_5865,N_5590);
nand U6376 (N_6376,N_5828,N_5576);
and U6377 (N_6377,N_5441,N_5921);
and U6378 (N_6378,N_5447,N_5233);
or U6379 (N_6379,N_5908,N_5519);
and U6380 (N_6380,N_5640,N_5787);
nand U6381 (N_6381,N_5903,N_5748);
nor U6382 (N_6382,N_5860,N_5144);
or U6383 (N_6383,N_5243,N_5167);
or U6384 (N_6384,N_5199,N_5715);
or U6385 (N_6385,N_5294,N_5314);
nor U6386 (N_6386,N_5637,N_5106);
and U6387 (N_6387,N_5871,N_5847);
nor U6388 (N_6388,N_5070,N_5335);
or U6389 (N_6389,N_5711,N_5390);
and U6390 (N_6390,N_5176,N_5415);
nand U6391 (N_6391,N_5248,N_5482);
or U6392 (N_6392,N_5309,N_5817);
nor U6393 (N_6393,N_5050,N_5647);
and U6394 (N_6394,N_5744,N_5939);
and U6395 (N_6395,N_5545,N_5672);
and U6396 (N_6396,N_5009,N_5574);
nand U6397 (N_6397,N_5351,N_5022);
nand U6398 (N_6398,N_5031,N_5798);
nor U6399 (N_6399,N_5073,N_5608);
xnor U6400 (N_6400,N_5262,N_5086);
nand U6401 (N_6401,N_5040,N_5271);
or U6402 (N_6402,N_5360,N_5789);
or U6403 (N_6403,N_5501,N_5956);
or U6404 (N_6404,N_5473,N_5896);
and U6405 (N_6405,N_5771,N_5950);
or U6406 (N_6406,N_5295,N_5955);
nand U6407 (N_6407,N_5869,N_5363);
nor U6408 (N_6408,N_5260,N_5977);
or U6409 (N_6409,N_5463,N_5146);
nor U6410 (N_6410,N_5062,N_5109);
nand U6411 (N_6411,N_5995,N_5147);
nor U6412 (N_6412,N_5405,N_5535);
nor U6413 (N_6413,N_5818,N_5886);
nor U6414 (N_6414,N_5819,N_5290);
or U6415 (N_6415,N_5583,N_5775);
nand U6416 (N_6416,N_5132,N_5348);
or U6417 (N_6417,N_5435,N_5337);
nand U6418 (N_6418,N_5196,N_5468);
nand U6419 (N_6419,N_5207,N_5209);
nand U6420 (N_6420,N_5962,N_5665);
or U6421 (N_6421,N_5688,N_5925);
nand U6422 (N_6422,N_5487,N_5486);
nor U6423 (N_6423,N_5049,N_5881);
nand U6424 (N_6424,N_5429,N_5849);
and U6425 (N_6425,N_5581,N_5315);
and U6426 (N_6426,N_5102,N_5478);
and U6427 (N_6427,N_5100,N_5133);
and U6428 (N_6428,N_5694,N_5876);
and U6429 (N_6429,N_5504,N_5082);
nor U6430 (N_6430,N_5578,N_5976);
nor U6431 (N_6431,N_5021,N_5809);
and U6432 (N_6432,N_5978,N_5149);
nor U6433 (N_6433,N_5130,N_5918);
nand U6434 (N_6434,N_5884,N_5770);
or U6435 (N_6435,N_5056,N_5625);
nand U6436 (N_6436,N_5699,N_5680);
and U6437 (N_6437,N_5846,N_5011);
and U6438 (N_6438,N_5923,N_5020);
nand U6439 (N_6439,N_5801,N_5996);
and U6440 (N_6440,N_5510,N_5274);
and U6441 (N_6441,N_5115,N_5974);
nor U6442 (N_6442,N_5201,N_5938);
or U6443 (N_6443,N_5826,N_5930);
nor U6444 (N_6444,N_5794,N_5916);
and U6445 (N_6445,N_5433,N_5323);
or U6446 (N_6446,N_5252,N_5927);
and U6447 (N_6447,N_5340,N_5971);
nand U6448 (N_6448,N_5326,N_5546);
and U6449 (N_6449,N_5341,N_5139);
nand U6450 (N_6450,N_5492,N_5357);
nand U6451 (N_6451,N_5171,N_5427);
nand U6452 (N_6452,N_5691,N_5525);
nand U6453 (N_6453,N_5984,N_5693);
and U6454 (N_6454,N_5401,N_5666);
nand U6455 (N_6455,N_5793,N_5440);
or U6456 (N_6456,N_5388,N_5676);
or U6457 (N_6457,N_5366,N_5090);
xnor U6458 (N_6458,N_5655,N_5848);
nand U6459 (N_6459,N_5609,N_5217);
nor U6460 (N_6460,N_5838,N_5135);
nand U6461 (N_6461,N_5143,N_5890);
nor U6462 (N_6462,N_5455,N_5516);
or U6463 (N_6463,N_5937,N_5522);
and U6464 (N_6464,N_5166,N_5782);
or U6465 (N_6465,N_5002,N_5788);
or U6466 (N_6466,N_5211,N_5755);
nand U6467 (N_6467,N_5163,N_5203);
and U6468 (N_6468,N_5169,N_5811);
and U6469 (N_6469,N_5662,N_5125);
nand U6470 (N_6470,N_5507,N_5840);
or U6471 (N_6471,N_5362,N_5905);
or U6472 (N_6472,N_5856,N_5034);
nor U6473 (N_6473,N_5812,N_5623);
and U6474 (N_6474,N_5375,N_5023);
nor U6475 (N_6475,N_5571,N_5600);
nor U6476 (N_6476,N_5766,N_5813);
nor U6477 (N_6477,N_5909,N_5780);
nor U6478 (N_6478,N_5078,N_5068);
nand U6479 (N_6479,N_5064,N_5750);
and U6480 (N_6480,N_5136,N_5219);
nand U6481 (N_6481,N_5458,N_5076);
or U6482 (N_6482,N_5080,N_5284);
or U6483 (N_6483,N_5246,N_5807);
and U6484 (N_6484,N_5044,N_5634);
and U6485 (N_6485,N_5214,N_5967);
nor U6486 (N_6486,N_5126,N_5703);
or U6487 (N_6487,N_5887,N_5015);
nor U6488 (N_6488,N_5808,N_5991);
nand U6489 (N_6489,N_5247,N_5761);
and U6490 (N_6490,N_5475,N_5825);
or U6491 (N_6491,N_5863,N_5377);
nor U6492 (N_6492,N_5208,N_5129);
nand U6493 (N_6493,N_5398,N_5951);
xnor U6494 (N_6494,N_5190,N_5866);
or U6495 (N_6495,N_5279,N_5328);
and U6496 (N_6496,N_5030,N_5239);
and U6497 (N_6497,N_5639,N_5302);
and U6498 (N_6498,N_5599,N_5975);
and U6499 (N_6499,N_5663,N_5001);
nor U6500 (N_6500,N_5572,N_5346);
and U6501 (N_6501,N_5485,N_5003);
and U6502 (N_6502,N_5195,N_5218);
and U6503 (N_6503,N_5463,N_5324);
nand U6504 (N_6504,N_5605,N_5166);
or U6505 (N_6505,N_5370,N_5513);
and U6506 (N_6506,N_5744,N_5451);
or U6507 (N_6507,N_5226,N_5640);
nor U6508 (N_6508,N_5042,N_5267);
and U6509 (N_6509,N_5430,N_5310);
and U6510 (N_6510,N_5208,N_5432);
and U6511 (N_6511,N_5116,N_5345);
nand U6512 (N_6512,N_5024,N_5109);
and U6513 (N_6513,N_5497,N_5345);
nor U6514 (N_6514,N_5376,N_5157);
and U6515 (N_6515,N_5105,N_5519);
and U6516 (N_6516,N_5118,N_5398);
nor U6517 (N_6517,N_5613,N_5345);
nor U6518 (N_6518,N_5482,N_5714);
nand U6519 (N_6519,N_5250,N_5901);
nor U6520 (N_6520,N_5092,N_5483);
nand U6521 (N_6521,N_5328,N_5632);
and U6522 (N_6522,N_5654,N_5691);
nand U6523 (N_6523,N_5973,N_5961);
nand U6524 (N_6524,N_5369,N_5402);
and U6525 (N_6525,N_5256,N_5194);
and U6526 (N_6526,N_5488,N_5389);
or U6527 (N_6527,N_5294,N_5712);
nor U6528 (N_6528,N_5725,N_5447);
and U6529 (N_6529,N_5179,N_5437);
or U6530 (N_6530,N_5551,N_5386);
nand U6531 (N_6531,N_5510,N_5944);
nor U6532 (N_6532,N_5873,N_5082);
nand U6533 (N_6533,N_5414,N_5367);
nand U6534 (N_6534,N_5939,N_5422);
nor U6535 (N_6535,N_5291,N_5270);
or U6536 (N_6536,N_5870,N_5320);
or U6537 (N_6537,N_5057,N_5299);
nor U6538 (N_6538,N_5641,N_5213);
or U6539 (N_6539,N_5207,N_5378);
or U6540 (N_6540,N_5547,N_5197);
nand U6541 (N_6541,N_5126,N_5851);
or U6542 (N_6542,N_5863,N_5355);
nor U6543 (N_6543,N_5092,N_5976);
or U6544 (N_6544,N_5798,N_5414);
nor U6545 (N_6545,N_5105,N_5577);
and U6546 (N_6546,N_5591,N_5587);
nor U6547 (N_6547,N_5148,N_5154);
and U6548 (N_6548,N_5949,N_5576);
or U6549 (N_6549,N_5116,N_5456);
or U6550 (N_6550,N_5598,N_5191);
and U6551 (N_6551,N_5905,N_5974);
nand U6552 (N_6552,N_5290,N_5292);
and U6553 (N_6553,N_5917,N_5614);
nand U6554 (N_6554,N_5217,N_5871);
and U6555 (N_6555,N_5547,N_5267);
or U6556 (N_6556,N_5969,N_5831);
nor U6557 (N_6557,N_5383,N_5714);
or U6558 (N_6558,N_5831,N_5730);
nor U6559 (N_6559,N_5772,N_5397);
or U6560 (N_6560,N_5852,N_5256);
nor U6561 (N_6561,N_5718,N_5842);
nor U6562 (N_6562,N_5312,N_5131);
or U6563 (N_6563,N_5566,N_5062);
and U6564 (N_6564,N_5534,N_5193);
nor U6565 (N_6565,N_5976,N_5570);
and U6566 (N_6566,N_5396,N_5636);
or U6567 (N_6567,N_5692,N_5147);
nor U6568 (N_6568,N_5984,N_5355);
or U6569 (N_6569,N_5465,N_5527);
nand U6570 (N_6570,N_5320,N_5389);
nand U6571 (N_6571,N_5735,N_5641);
nor U6572 (N_6572,N_5159,N_5494);
nand U6573 (N_6573,N_5572,N_5528);
and U6574 (N_6574,N_5680,N_5104);
and U6575 (N_6575,N_5027,N_5213);
nor U6576 (N_6576,N_5110,N_5653);
nand U6577 (N_6577,N_5525,N_5289);
and U6578 (N_6578,N_5688,N_5634);
and U6579 (N_6579,N_5933,N_5321);
nor U6580 (N_6580,N_5349,N_5859);
nand U6581 (N_6581,N_5788,N_5854);
or U6582 (N_6582,N_5301,N_5264);
and U6583 (N_6583,N_5658,N_5486);
or U6584 (N_6584,N_5782,N_5084);
nor U6585 (N_6585,N_5865,N_5578);
nand U6586 (N_6586,N_5679,N_5008);
or U6587 (N_6587,N_5039,N_5073);
nor U6588 (N_6588,N_5272,N_5863);
nor U6589 (N_6589,N_5179,N_5960);
nor U6590 (N_6590,N_5702,N_5451);
nand U6591 (N_6591,N_5679,N_5605);
nand U6592 (N_6592,N_5675,N_5261);
nor U6593 (N_6593,N_5215,N_5531);
or U6594 (N_6594,N_5205,N_5420);
and U6595 (N_6595,N_5798,N_5135);
and U6596 (N_6596,N_5919,N_5697);
nor U6597 (N_6597,N_5521,N_5601);
nor U6598 (N_6598,N_5410,N_5394);
and U6599 (N_6599,N_5063,N_5615);
xor U6600 (N_6600,N_5829,N_5149);
or U6601 (N_6601,N_5947,N_5561);
nand U6602 (N_6602,N_5013,N_5880);
nand U6603 (N_6603,N_5774,N_5475);
and U6604 (N_6604,N_5739,N_5717);
or U6605 (N_6605,N_5809,N_5721);
and U6606 (N_6606,N_5381,N_5302);
or U6607 (N_6607,N_5451,N_5591);
and U6608 (N_6608,N_5501,N_5138);
nand U6609 (N_6609,N_5555,N_5121);
nand U6610 (N_6610,N_5642,N_5904);
xor U6611 (N_6611,N_5378,N_5629);
or U6612 (N_6612,N_5926,N_5884);
or U6613 (N_6613,N_5138,N_5810);
and U6614 (N_6614,N_5205,N_5098);
or U6615 (N_6615,N_5169,N_5015);
or U6616 (N_6616,N_5484,N_5217);
nor U6617 (N_6617,N_5969,N_5189);
and U6618 (N_6618,N_5962,N_5718);
or U6619 (N_6619,N_5394,N_5209);
nor U6620 (N_6620,N_5222,N_5849);
and U6621 (N_6621,N_5701,N_5197);
nand U6622 (N_6622,N_5329,N_5339);
nor U6623 (N_6623,N_5622,N_5307);
nor U6624 (N_6624,N_5866,N_5843);
and U6625 (N_6625,N_5664,N_5500);
and U6626 (N_6626,N_5573,N_5892);
nand U6627 (N_6627,N_5501,N_5949);
nor U6628 (N_6628,N_5448,N_5609);
nand U6629 (N_6629,N_5164,N_5136);
nand U6630 (N_6630,N_5122,N_5939);
nand U6631 (N_6631,N_5897,N_5819);
and U6632 (N_6632,N_5185,N_5794);
and U6633 (N_6633,N_5632,N_5653);
nand U6634 (N_6634,N_5824,N_5788);
nor U6635 (N_6635,N_5375,N_5208);
and U6636 (N_6636,N_5401,N_5775);
or U6637 (N_6637,N_5761,N_5498);
or U6638 (N_6638,N_5106,N_5928);
or U6639 (N_6639,N_5995,N_5575);
or U6640 (N_6640,N_5796,N_5638);
and U6641 (N_6641,N_5958,N_5442);
and U6642 (N_6642,N_5939,N_5859);
or U6643 (N_6643,N_5800,N_5260);
nand U6644 (N_6644,N_5026,N_5796);
or U6645 (N_6645,N_5252,N_5295);
nor U6646 (N_6646,N_5676,N_5412);
nand U6647 (N_6647,N_5327,N_5516);
or U6648 (N_6648,N_5664,N_5841);
nand U6649 (N_6649,N_5843,N_5363);
nand U6650 (N_6650,N_5161,N_5475);
or U6651 (N_6651,N_5018,N_5688);
nor U6652 (N_6652,N_5911,N_5611);
nand U6653 (N_6653,N_5221,N_5106);
nand U6654 (N_6654,N_5818,N_5131);
nor U6655 (N_6655,N_5261,N_5876);
nand U6656 (N_6656,N_5924,N_5528);
and U6657 (N_6657,N_5185,N_5073);
and U6658 (N_6658,N_5631,N_5028);
and U6659 (N_6659,N_5424,N_5975);
and U6660 (N_6660,N_5460,N_5365);
nor U6661 (N_6661,N_5955,N_5668);
and U6662 (N_6662,N_5903,N_5637);
nand U6663 (N_6663,N_5041,N_5625);
nor U6664 (N_6664,N_5339,N_5356);
nor U6665 (N_6665,N_5027,N_5138);
or U6666 (N_6666,N_5797,N_5176);
nor U6667 (N_6667,N_5258,N_5588);
nand U6668 (N_6668,N_5341,N_5672);
or U6669 (N_6669,N_5127,N_5718);
and U6670 (N_6670,N_5028,N_5499);
nand U6671 (N_6671,N_5793,N_5770);
or U6672 (N_6672,N_5238,N_5791);
and U6673 (N_6673,N_5010,N_5725);
or U6674 (N_6674,N_5824,N_5405);
xor U6675 (N_6675,N_5024,N_5265);
nor U6676 (N_6676,N_5187,N_5695);
and U6677 (N_6677,N_5465,N_5247);
nand U6678 (N_6678,N_5159,N_5987);
nor U6679 (N_6679,N_5014,N_5496);
nand U6680 (N_6680,N_5241,N_5400);
or U6681 (N_6681,N_5754,N_5002);
or U6682 (N_6682,N_5934,N_5548);
and U6683 (N_6683,N_5809,N_5466);
nor U6684 (N_6684,N_5017,N_5425);
or U6685 (N_6685,N_5805,N_5204);
nor U6686 (N_6686,N_5465,N_5773);
or U6687 (N_6687,N_5806,N_5306);
nand U6688 (N_6688,N_5809,N_5276);
nand U6689 (N_6689,N_5043,N_5720);
nand U6690 (N_6690,N_5658,N_5273);
or U6691 (N_6691,N_5138,N_5734);
nand U6692 (N_6692,N_5204,N_5711);
nor U6693 (N_6693,N_5164,N_5524);
and U6694 (N_6694,N_5547,N_5404);
and U6695 (N_6695,N_5418,N_5458);
nor U6696 (N_6696,N_5456,N_5213);
and U6697 (N_6697,N_5550,N_5177);
and U6698 (N_6698,N_5238,N_5889);
and U6699 (N_6699,N_5335,N_5468);
and U6700 (N_6700,N_5430,N_5112);
nor U6701 (N_6701,N_5424,N_5715);
nand U6702 (N_6702,N_5564,N_5820);
and U6703 (N_6703,N_5195,N_5727);
nor U6704 (N_6704,N_5228,N_5884);
xor U6705 (N_6705,N_5665,N_5966);
or U6706 (N_6706,N_5785,N_5363);
or U6707 (N_6707,N_5648,N_5248);
and U6708 (N_6708,N_5100,N_5364);
and U6709 (N_6709,N_5717,N_5332);
nor U6710 (N_6710,N_5447,N_5074);
and U6711 (N_6711,N_5736,N_5122);
and U6712 (N_6712,N_5785,N_5897);
and U6713 (N_6713,N_5646,N_5062);
or U6714 (N_6714,N_5533,N_5284);
nand U6715 (N_6715,N_5505,N_5333);
and U6716 (N_6716,N_5272,N_5102);
or U6717 (N_6717,N_5133,N_5305);
nand U6718 (N_6718,N_5996,N_5599);
nand U6719 (N_6719,N_5687,N_5367);
or U6720 (N_6720,N_5670,N_5812);
or U6721 (N_6721,N_5205,N_5182);
and U6722 (N_6722,N_5549,N_5072);
nor U6723 (N_6723,N_5905,N_5958);
nand U6724 (N_6724,N_5234,N_5222);
or U6725 (N_6725,N_5240,N_5007);
or U6726 (N_6726,N_5817,N_5242);
and U6727 (N_6727,N_5644,N_5517);
or U6728 (N_6728,N_5245,N_5413);
nor U6729 (N_6729,N_5144,N_5361);
nand U6730 (N_6730,N_5251,N_5518);
or U6731 (N_6731,N_5828,N_5982);
nand U6732 (N_6732,N_5512,N_5982);
or U6733 (N_6733,N_5815,N_5259);
nand U6734 (N_6734,N_5557,N_5608);
and U6735 (N_6735,N_5104,N_5614);
nor U6736 (N_6736,N_5829,N_5423);
nand U6737 (N_6737,N_5227,N_5839);
nand U6738 (N_6738,N_5674,N_5162);
nand U6739 (N_6739,N_5523,N_5322);
or U6740 (N_6740,N_5865,N_5494);
and U6741 (N_6741,N_5514,N_5836);
nand U6742 (N_6742,N_5023,N_5287);
nand U6743 (N_6743,N_5405,N_5205);
or U6744 (N_6744,N_5008,N_5460);
or U6745 (N_6745,N_5456,N_5169);
or U6746 (N_6746,N_5160,N_5737);
nor U6747 (N_6747,N_5605,N_5505);
nand U6748 (N_6748,N_5209,N_5700);
xnor U6749 (N_6749,N_5381,N_5983);
and U6750 (N_6750,N_5924,N_5905);
nand U6751 (N_6751,N_5576,N_5586);
nor U6752 (N_6752,N_5260,N_5991);
nand U6753 (N_6753,N_5601,N_5643);
or U6754 (N_6754,N_5891,N_5261);
nand U6755 (N_6755,N_5046,N_5946);
or U6756 (N_6756,N_5552,N_5069);
and U6757 (N_6757,N_5098,N_5635);
nand U6758 (N_6758,N_5900,N_5264);
nand U6759 (N_6759,N_5943,N_5671);
and U6760 (N_6760,N_5288,N_5744);
nor U6761 (N_6761,N_5319,N_5031);
nor U6762 (N_6762,N_5351,N_5165);
or U6763 (N_6763,N_5954,N_5784);
nand U6764 (N_6764,N_5461,N_5321);
and U6765 (N_6765,N_5207,N_5902);
or U6766 (N_6766,N_5680,N_5300);
nor U6767 (N_6767,N_5027,N_5849);
nor U6768 (N_6768,N_5602,N_5095);
or U6769 (N_6769,N_5059,N_5496);
nor U6770 (N_6770,N_5479,N_5820);
nor U6771 (N_6771,N_5229,N_5638);
and U6772 (N_6772,N_5412,N_5082);
and U6773 (N_6773,N_5178,N_5588);
nor U6774 (N_6774,N_5767,N_5213);
nor U6775 (N_6775,N_5808,N_5685);
nor U6776 (N_6776,N_5043,N_5960);
and U6777 (N_6777,N_5567,N_5185);
or U6778 (N_6778,N_5598,N_5286);
and U6779 (N_6779,N_5576,N_5859);
nor U6780 (N_6780,N_5716,N_5060);
nor U6781 (N_6781,N_5679,N_5007);
nor U6782 (N_6782,N_5085,N_5856);
and U6783 (N_6783,N_5133,N_5977);
and U6784 (N_6784,N_5516,N_5225);
nor U6785 (N_6785,N_5854,N_5034);
nor U6786 (N_6786,N_5264,N_5835);
nor U6787 (N_6787,N_5697,N_5529);
or U6788 (N_6788,N_5133,N_5033);
nor U6789 (N_6789,N_5191,N_5945);
or U6790 (N_6790,N_5664,N_5786);
nor U6791 (N_6791,N_5142,N_5541);
nor U6792 (N_6792,N_5786,N_5779);
nor U6793 (N_6793,N_5627,N_5588);
and U6794 (N_6794,N_5538,N_5219);
nor U6795 (N_6795,N_5414,N_5621);
or U6796 (N_6796,N_5937,N_5301);
nand U6797 (N_6797,N_5952,N_5082);
and U6798 (N_6798,N_5993,N_5803);
nor U6799 (N_6799,N_5637,N_5438);
nor U6800 (N_6800,N_5940,N_5389);
nand U6801 (N_6801,N_5002,N_5432);
nor U6802 (N_6802,N_5529,N_5588);
nand U6803 (N_6803,N_5718,N_5629);
or U6804 (N_6804,N_5516,N_5205);
nand U6805 (N_6805,N_5946,N_5706);
nor U6806 (N_6806,N_5248,N_5753);
nor U6807 (N_6807,N_5271,N_5319);
and U6808 (N_6808,N_5187,N_5601);
nor U6809 (N_6809,N_5862,N_5041);
and U6810 (N_6810,N_5364,N_5586);
nor U6811 (N_6811,N_5816,N_5012);
nand U6812 (N_6812,N_5023,N_5918);
or U6813 (N_6813,N_5367,N_5811);
nor U6814 (N_6814,N_5631,N_5652);
or U6815 (N_6815,N_5910,N_5195);
and U6816 (N_6816,N_5136,N_5224);
nor U6817 (N_6817,N_5009,N_5804);
and U6818 (N_6818,N_5339,N_5393);
nor U6819 (N_6819,N_5049,N_5458);
nor U6820 (N_6820,N_5958,N_5455);
nand U6821 (N_6821,N_5643,N_5187);
nand U6822 (N_6822,N_5877,N_5597);
nand U6823 (N_6823,N_5982,N_5095);
nand U6824 (N_6824,N_5891,N_5574);
nor U6825 (N_6825,N_5700,N_5454);
nand U6826 (N_6826,N_5264,N_5420);
and U6827 (N_6827,N_5883,N_5362);
nand U6828 (N_6828,N_5003,N_5278);
or U6829 (N_6829,N_5499,N_5502);
nand U6830 (N_6830,N_5675,N_5203);
nand U6831 (N_6831,N_5727,N_5815);
or U6832 (N_6832,N_5311,N_5671);
and U6833 (N_6833,N_5626,N_5879);
or U6834 (N_6834,N_5569,N_5581);
nand U6835 (N_6835,N_5574,N_5716);
and U6836 (N_6836,N_5189,N_5014);
nor U6837 (N_6837,N_5132,N_5145);
or U6838 (N_6838,N_5482,N_5369);
or U6839 (N_6839,N_5397,N_5423);
and U6840 (N_6840,N_5038,N_5811);
and U6841 (N_6841,N_5053,N_5564);
or U6842 (N_6842,N_5242,N_5935);
nor U6843 (N_6843,N_5425,N_5187);
nor U6844 (N_6844,N_5911,N_5476);
or U6845 (N_6845,N_5512,N_5689);
or U6846 (N_6846,N_5996,N_5335);
nand U6847 (N_6847,N_5805,N_5693);
and U6848 (N_6848,N_5873,N_5987);
nor U6849 (N_6849,N_5274,N_5470);
and U6850 (N_6850,N_5646,N_5844);
and U6851 (N_6851,N_5961,N_5597);
and U6852 (N_6852,N_5652,N_5801);
nand U6853 (N_6853,N_5493,N_5301);
and U6854 (N_6854,N_5135,N_5189);
or U6855 (N_6855,N_5181,N_5686);
nor U6856 (N_6856,N_5314,N_5470);
or U6857 (N_6857,N_5900,N_5145);
nor U6858 (N_6858,N_5748,N_5620);
nor U6859 (N_6859,N_5206,N_5002);
or U6860 (N_6860,N_5845,N_5010);
nand U6861 (N_6861,N_5821,N_5043);
nand U6862 (N_6862,N_5743,N_5419);
or U6863 (N_6863,N_5720,N_5592);
or U6864 (N_6864,N_5537,N_5724);
nor U6865 (N_6865,N_5926,N_5292);
or U6866 (N_6866,N_5730,N_5599);
nand U6867 (N_6867,N_5541,N_5070);
nand U6868 (N_6868,N_5156,N_5006);
and U6869 (N_6869,N_5389,N_5693);
or U6870 (N_6870,N_5919,N_5132);
and U6871 (N_6871,N_5419,N_5333);
nor U6872 (N_6872,N_5418,N_5563);
or U6873 (N_6873,N_5090,N_5837);
and U6874 (N_6874,N_5652,N_5176);
and U6875 (N_6875,N_5919,N_5592);
or U6876 (N_6876,N_5676,N_5613);
and U6877 (N_6877,N_5147,N_5658);
nor U6878 (N_6878,N_5236,N_5596);
or U6879 (N_6879,N_5885,N_5584);
nor U6880 (N_6880,N_5318,N_5721);
or U6881 (N_6881,N_5696,N_5660);
nand U6882 (N_6882,N_5856,N_5539);
nand U6883 (N_6883,N_5764,N_5453);
or U6884 (N_6884,N_5833,N_5047);
and U6885 (N_6885,N_5210,N_5473);
nor U6886 (N_6886,N_5132,N_5818);
or U6887 (N_6887,N_5539,N_5780);
and U6888 (N_6888,N_5678,N_5765);
and U6889 (N_6889,N_5386,N_5467);
and U6890 (N_6890,N_5423,N_5533);
and U6891 (N_6891,N_5267,N_5370);
nand U6892 (N_6892,N_5400,N_5837);
nand U6893 (N_6893,N_5235,N_5967);
or U6894 (N_6894,N_5620,N_5759);
nor U6895 (N_6895,N_5769,N_5081);
nand U6896 (N_6896,N_5992,N_5957);
nand U6897 (N_6897,N_5983,N_5771);
or U6898 (N_6898,N_5896,N_5293);
nor U6899 (N_6899,N_5952,N_5127);
or U6900 (N_6900,N_5313,N_5591);
nand U6901 (N_6901,N_5260,N_5325);
nor U6902 (N_6902,N_5538,N_5718);
nand U6903 (N_6903,N_5328,N_5246);
or U6904 (N_6904,N_5873,N_5637);
and U6905 (N_6905,N_5100,N_5502);
nor U6906 (N_6906,N_5909,N_5124);
nor U6907 (N_6907,N_5371,N_5899);
and U6908 (N_6908,N_5818,N_5418);
and U6909 (N_6909,N_5007,N_5126);
and U6910 (N_6910,N_5289,N_5597);
nor U6911 (N_6911,N_5270,N_5504);
nor U6912 (N_6912,N_5276,N_5856);
or U6913 (N_6913,N_5790,N_5451);
or U6914 (N_6914,N_5782,N_5069);
nor U6915 (N_6915,N_5083,N_5185);
or U6916 (N_6916,N_5730,N_5013);
and U6917 (N_6917,N_5065,N_5235);
nor U6918 (N_6918,N_5191,N_5161);
or U6919 (N_6919,N_5478,N_5745);
and U6920 (N_6920,N_5918,N_5693);
and U6921 (N_6921,N_5635,N_5941);
nand U6922 (N_6922,N_5330,N_5194);
and U6923 (N_6923,N_5042,N_5615);
or U6924 (N_6924,N_5259,N_5736);
or U6925 (N_6925,N_5300,N_5178);
nor U6926 (N_6926,N_5948,N_5722);
nand U6927 (N_6927,N_5017,N_5592);
or U6928 (N_6928,N_5524,N_5785);
nand U6929 (N_6929,N_5424,N_5120);
and U6930 (N_6930,N_5818,N_5773);
or U6931 (N_6931,N_5687,N_5733);
nand U6932 (N_6932,N_5569,N_5834);
or U6933 (N_6933,N_5448,N_5225);
nand U6934 (N_6934,N_5697,N_5390);
and U6935 (N_6935,N_5493,N_5582);
or U6936 (N_6936,N_5043,N_5922);
nand U6937 (N_6937,N_5571,N_5115);
or U6938 (N_6938,N_5723,N_5467);
nor U6939 (N_6939,N_5402,N_5638);
nand U6940 (N_6940,N_5496,N_5943);
and U6941 (N_6941,N_5817,N_5048);
nor U6942 (N_6942,N_5320,N_5359);
and U6943 (N_6943,N_5536,N_5145);
nor U6944 (N_6944,N_5528,N_5502);
and U6945 (N_6945,N_5829,N_5607);
or U6946 (N_6946,N_5967,N_5203);
xor U6947 (N_6947,N_5405,N_5032);
and U6948 (N_6948,N_5140,N_5164);
and U6949 (N_6949,N_5487,N_5080);
and U6950 (N_6950,N_5578,N_5034);
or U6951 (N_6951,N_5339,N_5951);
nand U6952 (N_6952,N_5789,N_5865);
or U6953 (N_6953,N_5153,N_5761);
and U6954 (N_6954,N_5134,N_5688);
nor U6955 (N_6955,N_5992,N_5221);
and U6956 (N_6956,N_5911,N_5986);
or U6957 (N_6957,N_5828,N_5146);
nor U6958 (N_6958,N_5244,N_5126);
or U6959 (N_6959,N_5908,N_5919);
or U6960 (N_6960,N_5747,N_5523);
and U6961 (N_6961,N_5431,N_5889);
nor U6962 (N_6962,N_5446,N_5838);
nand U6963 (N_6963,N_5834,N_5253);
nand U6964 (N_6964,N_5274,N_5319);
and U6965 (N_6965,N_5734,N_5846);
and U6966 (N_6966,N_5702,N_5687);
or U6967 (N_6967,N_5253,N_5615);
nand U6968 (N_6968,N_5997,N_5742);
nor U6969 (N_6969,N_5035,N_5523);
or U6970 (N_6970,N_5303,N_5203);
nor U6971 (N_6971,N_5692,N_5482);
or U6972 (N_6972,N_5423,N_5017);
or U6973 (N_6973,N_5775,N_5223);
xor U6974 (N_6974,N_5166,N_5802);
nor U6975 (N_6975,N_5702,N_5222);
or U6976 (N_6976,N_5773,N_5864);
and U6977 (N_6977,N_5858,N_5939);
nand U6978 (N_6978,N_5620,N_5248);
nand U6979 (N_6979,N_5108,N_5746);
and U6980 (N_6980,N_5962,N_5480);
nand U6981 (N_6981,N_5391,N_5842);
nand U6982 (N_6982,N_5115,N_5283);
and U6983 (N_6983,N_5794,N_5813);
nor U6984 (N_6984,N_5279,N_5134);
nor U6985 (N_6985,N_5363,N_5327);
and U6986 (N_6986,N_5841,N_5960);
and U6987 (N_6987,N_5232,N_5431);
or U6988 (N_6988,N_5155,N_5468);
or U6989 (N_6989,N_5731,N_5236);
nand U6990 (N_6990,N_5954,N_5036);
nand U6991 (N_6991,N_5330,N_5223);
or U6992 (N_6992,N_5564,N_5265);
and U6993 (N_6993,N_5704,N_5110);
and U6994 (N_6994,N_5977,N_5054);
nand U6995 (N_6995,N_5422,N_5187);
nand U6996 (N_6996,N_5524,N_5244);
nor U6997 (N_6997,N_5979,N_5643);
nand U6998 (N_6998,N_5435,N_5441);
nand U6999 (N_6999,N_5362,N_5870);
or U7000 (N_7000,N_6673,N_6837);
and U7001 (N_7001,N_6128,N_6008);
and U7002 (N_7002,N_6378,N_6505);
and U7003 (N_7003,N_6232,N_6050);
nand U7004 (N_7004,N_6330,N_6353);
nor U7005 (N_7005,N_6731,N_6918);
nand U7006 (N_7006,N_6937,N_6254);
nor U7007 (N_7007,N_6829,N_6181);
and U7008 (N_7008,N_6500,N_6688);
nand U7009 (N_7009,N_6896,N_6068);
and U7010 (N_7010,N_6938,N_6146);
nand U7011 (N_7011,N_6780,N_6917);
nand U7012 (N_7012,N_6321,N_6377);
nor U7013 (N_7013,N_6222,N_6549);
nor U7014 (N_7014,N_6558,N_6887);
or U7015 (N_7015,N_6230,N_6596);
nand U7016 (N_7016,N_6809,N_6812);
nand U7017 (N_7017,N_6901,N_6478);
nand U7018 (N_7018,N_6432,N_6934);
or U7019 (N_7019,N_6618,N_6269);
and U7020 (N_7020,N_6376,N_6773);
or U7021 (N_7021,N_6899,N_6644);
or U7022 (N_7022,N_6648,N_6808);
and U7023 (N_7023,N_6294,N_6924);
nand U7024 (N_7024,N_6411,N_6295);
nand U7025 (N_7025,N_6891,N_6234);
and U7026 (N_7026,N_6779,N_6586);
nand U7027 (N_7027,N_6886,N_6667);
nand U7028 (N_7028,N_6297,N_6540);
nand U7029 (N_7029,N_6952,N_6959);
nor U7030 (N_7030,N_6863,N_6341);
and U7031 (N_7031,N_6038,N_6753);
or U7032 (N_7032,N_6656,N_6594);
and U7033 (N_7033,N_6970,N_6554);
nand U7034 (N_7034,N_6125,N_6249);
nand U7035 (N_7035,N_6717,N_6971);
nand U7036 (N_7036,N_6360,N_6787);
and U7037 (N_7037,N_6289,N_6607);
nand U7038 (N_7038,N_6977,N_6592);
and U7039 (N_7039,N_6501,N_6526);
nand U7040 (N_7040,N_6851,N_6010);
or U7041 (N_7041,N_6778,N_6075);
and U7042 (N_7042,N_6845,N_6444);
or U7043 (N_7043,N_6794,N_6331);
nor U7044 (N_7044,N_6923,N_6898);
or U7045 (N_7045,N_6528,N_6218);
and U7046 (N_7046,N_6916,N_6797);
or U7047 (N_7047,N_6091,N_6314);
or U7048 (N_7048,N_6132,N_6534);
nor U7049 (N_7049,N_6102,N_6951);
and U7050 (N_7050,N_6270,N_6827);
nor U7051 (N_7051,N_6978,N_6196);
and U7052 (N_7052,N_6097,N_6548);
and U7053 (N_7053,N_6749,N_6859);
nand U7054 (N_7054,N_6383,N_6697);
nand U7055 (N_7055,N_6271,N_6490);
nor U7056 (N_7056,N_6210,N_6318);
nor U7057 (N_7057,N_6202,N_6035);
nor U7058 (N_7058,N_6395,N_6171);
and U7059 (N_7059,N_6718,N_6198);
xor U7060 (N_7060,N_6735,N_6416);
nand U7061 (N_7061,N_6519,N_6909);
or U7062 (N_7062,N_6724,N_6908);
and U7063 (N_7063,N_6776,N_6538);
nand U7064 (N_7064,N_6518,N_6872);
nand U7065 (N_7065,N_6085,N_6728);
nor U7066 (N_7066,N_6083,N_6458);
nand U7067 (N_7067,N_6374,N_6742);
or U7068 (N_7068,N_6087,N_6180);
or U7069 (N_7069,N_6743,N_6134);
nor U7070 (N_7070,N_6893,N_6373);
and U7071 (N_7071,N_6720,N_6939);
and U7072 (N_7072,N_6203,N_6228);
nor U7073 (N_7073,N_6092,N_6459);
or U7074 (N_7074,N_6604,N_6616);
or U7075 (N_7075,N_6640,N_6026);
nand U7076 (N_7076,N_6841,N_6105);
nor U7077 (N_7077,N_6094,N_6461);
nand U7078 (N_7078,N_6400,N_6600);
nand U7079 (N_7079,N_6802,N_6036);
and U7080 (N_7080,N_6191,N_6159);
nand U7081 (N_7081,N_6873,N_6860);
nor U7082 (N_7082,N_6523,N_6991);
or U7083 (N_7083,N_6089,N_6283);
nor U7084 (N_7084,N_6771,N_6848);
or U7085 (N_7085,N_6398,N_6646);
nor U7086 (N_7086,N_6713,N_6452);
nand U7087 (N_7087,N_6960,N_6947);
and U7088 (N_7088,N_6357,N_6264);
and U7089 (N_7089,N_6814,N_6804);
or U7090 (N_7090,N_6754,N_6462);
nand U7091 (N_7091,N_6765,N_6372);
nand U7092 (N_7092,N_6054,N_6682);
nor U7093 (N_7093,N_6073,N_6474);
or U7094 (N_7094,N_6403,N_6961);
nand U7095 (N_7095,N_6763,N_6935);
and U7096 (N_7096,N_6063,N_6869);
nor U7097 (N_7097,N_6621,N_6429);
nand U7098 (N_7098,N_6129,N_6530);
or U7099 (N_7099,N_6431,N_6581);
nor U7100 (N_7100,N_6066,N_6868);
and U7101 (N_7101,N_6172,N_6926);
and U7102 (N_7102,N_6605,N_6883);
xnor U7103 (N_7103,N_6986,N_6030);
nor U7104 (N_7104,N_6488,N_6155);
and U7105 (N_7105,N_6948,N_6525);
and U7106 (N_7106,N_6854,N_6984);
nand U7107 (N_7107,N_6906,N_6447);
nor U7108 (N_7108,N_6571,N_6866);
or U7109 (N_7109,N_6856,N_6072);
or U7110 (N_7110,N_6520,N_6288);
or U7111 (N_7111,N_6703,N_6052);
and U7112 (N_7112,N_6685,N_6897);
and U7113 (N_7113,N_6792,N_6274);
or U7114 (N_7114,N_6093,N_6996);
and U7115 (N_7115,N_6839,N_6903);
or U7116 (N_7116,N_6811,N_6699);
nor U7117 (N_7117,N_6700,N_6055);
nor U7118 (N_7118,N_6857,N_6838);
and U7119 (N_7119,N_6821,N_6136);
nor U7120 (N_7120,N_6497,N_6413);
nor U7121 (N_7121,N_6291,N_6529);
and U7122 (N_7122,N_6608,N_6610);
nand U7123 (N_7123,N_6723,N_6788);
or U7124 (N_7124,N_6775,N_6828);
and U7125 (N_7125,N_6211,N_6850);
and U7126 (N_7126,N_6243,N_6455);
or U7127 (N_7127,N_6624,N_6290);
or U7128 (N_7128,N_6645,N_6527);
or U7129 (N_7129,N_6840,N_6875);
nor U7130 (N_7130,N_6456,N_6510);
nor U7131 (N_7131,N_6823,N_6483);
or U7132 (N_7132,N_6547,N_6692);
nand U7133 (N_7133,N_6207,N_6106);
nor U7134 (N_7134,N_6985,N_6589);
nor U7135 (N_7135,N_6339,N_6852);
nand U7136 (N_7136,N_6932,N_6709);
and U7137 (N_7137,N_6074,N_6200);
nor U7138 (N_7138,N_6630,N_6084);
nor U7139 (N_7139,N_6966,N_6433);
nor U7140 (N_7140,N_6298,N_6414);
and U7141 (N_7141,N_6406,N_6698);
nand U7142 (N_7142,N_6936,N_6079);
nand U7143 (N_7143,N_6407,N_6800);
nor U7144 (N_7144,N_6475,N_6541);
nand U7145 (N_7145,N_6322,N_6681);
nand U7146 (N_7146,N_6384,N_6757);
nand U7147 (N_7147,N_6120,N_6810);
or U7148 (N_7148,N_6332,N_6964);
nand U7149 (N_7149,N_6992,N_6994);
or U7150 (N_7150,N_6195,N_6954);
or U7151 (N_7151,N_6774,N_6049);
nor U7152 (N_7152,N_6065,N_6516);
nor U7153 (N_7153,N_6722,N_6399);
and U7154 (N_7154,N_6577,N_6791);
or U7155 (N_7155,N_6409,N_6843);
and U7156 (N_7156,N_6153,N_6597);
and U7157 (N_7157,N_6205,N_6347);
and U7158 (N_7158,N_6263,N_6144);
and U7159 (N_7159,N_6613,N_6284);
or U7160 (N_7160,N_6212,N_6423);
and U7161 (N_7161,N_6362,N_6649);
and U7162 (N_7162,N_6498,N_6311);
nor U7163 (N_7163,N_6062,N_6436);
or U7164 (N_7164,N_6729,N_6216);
or U7165 (N_7165,N_6691,N_6336);
or U7166 (N_7166,N_6865,N_6018);
or U7167 (N_7167,N_6912,N_6585);
nand U7168 (N_7168,N_6273,N_6486);
nand U7169 (N_7169,N_6424,N_6714);
or U7170 (N_7170,N_6004,N_6037);
nand U7171 (N_7171,N_6428,N_6150);
nor U7172 (N_7172,N_6027,N_6515);
nand U7173 (N_7173,N_6612,N_6641);
nand U7174 (N_7174,N_6046,N_6024);
or U7175 (N_7175,N_6477,N_6513);
and U7176 (N_7176,N_6669,N_6081);
nand U7177 (N_7177,N_6250,N_6042);
or U7178 (N_7178,N_6166,N_6408);
nand U7179 (N_7179,N_6485,N_6217);
or U7180 (N_7180,N_6326,N_6175);
or U7181 (N_7181,N_6450,N_6048);
nor U7182 (N_7182,N_6178,N_6426);
xor U7183 (N_7183,N_6256,N_6257);
nand U7184 (N_7184,N_6664,N_6759);
or U7185 (N_7185,N_6696,N_6920);
and U7186 (N_7186,N_6242,N_6338);
and U7187 (N_7187,N_6005,N_6067);
nor U7188 (N_7188,N_6337,N_6580);
nor U7189 (N_7189,N_6739,N_6041);
nand U7190 (N_7190,N_6504,N_6014);
nor U7191 (N_7191,N_6650,N_6110);
and U7192 (N_7192,N_6118,N_6878);
nand U7193 (N_7193,N_6793,N_6312);
or U7194 (N_7194,N_6660,N_6358);
and U7195 (N_7195,N_6517,N_6296);
or U7196 (N_7196,N_6546,N_6417);
nand U7197 (N_7197,N_6394,N_6405);
nor U7198 (N_7198,N_6315,N_6238);
and U7199 (N_7199,N_6231,N_6975);
nor U7200 (N_7200,N_6340,N_6382);
or U7201 (N_7201,N_6979,N_6001);
nand U7202 (N_7202,N_6492,N_6747);
nand U7203 (N_7203,N_6642,N_6388);
nand U7204 (N_7204,N_6354,N_6100);
nor U7205 (N_7205,N_6012,N_6738);
or U7206 (N_7206,N_6675,N_6441);
nand U7207 (N_7207,N_6595,N_6190);
nand U7208 (N_7208,N_6545,N_6633);
or U7209 (N_7209,N_6109,N_6434);
nand U7210 (N_7210,N_6777,N_6715);
or U7211 (N_7211,N_6189,N_6997);
nand U7212 (N_7212,N_6152,N_6929);
and U7213 (N_7213,N_6907,N_6647);
nand U7214 (N_7214,N_6583,N_6987);
nand U7215 (N_7215,N_6278,N_6532);
nand U7216 (N_7216,N_6016,N_6188);
nand U7217 (N_7217,N_6366,N_6522);
and U7218 (N_7218,N_6367,N_6080);
nand U7219 (N_7219,N_6389,N_6834);
and U7220 (N_7220,N_6884,N_6862);
or U7221 (N_7221,N_6861,N_6849);
nor U7222 (N_7222,N_6168,N_6327);
nand U7223 (N_7223,N_6151,N_6575);
nand U7224 (N_7224,N_6652,N_6602);
or U7225 (N_7225,N_6858,N_6401);
nand U7226 (N_7226,N_6043,N_6380);
and U7227 (N_7227,N_6846,N_6201);
nand U7228 (N_7228,N_6396,N_6512);
nand U7229 (N_7229,N_6437,N_6040);
nor U7230 (N_7230,N_6686,N_6412);
or U7231 (N_7231,N_6603,N_6625);
nand U7232 (N_7232,N_6045,N_6184);
and U7233 (N_7233,N_6162,N_6782);
or U7234 (N_7234,N_6798,N_6535);
and U7235 (N_7235,N_6343,N_6847);
nor U7236 (N_7236,N_6945,N_6069);
or U7237 (N_7237,N_6364,N_6941);
nor U7238 (N_7238,N_6033,N_6761);
nand U7239 (N_7239,N_6557,N_6344);
or U7240 (N_7240,N_6114,N_6721);
nand U7241 (N_7241,N_6221,N_6113);
and U7242 (N_7242,N_6116,N_6174);
and U7243 (N_7243,N_6126,N_6748);
and U7244 (N_7244,N_6160,N_6556);
or U7245 (N_7245,N_6371,N_6694);
nand U7246 (N_7246,N_6768,N_6261);
nand U7247 (N_7247,N_6300,N_6259);
or U7248 (N_7248,N_6363,N_6825);
nand U7249 (N_7249,N_6468,N_6689);
nand U7250 (N_7250,N_6308,N_6995);
nand U7251 (N_7251,N_6781,N_6919);
nand U7252 (N_7252,N_6208,N_6017);
nand U7253 (N_7253,N_6659,N_6764);
and U7254 (N_7254,N_6310,N_6668);
or U7255 (N_7255,N_6506,N_6487);
or U7256 (N_7256,N_6157,N_6870);
and U7257 (N_7257,N_6021,N_6766);
or U7258 (N_7258,N_6143,N_6223);
or U7259 (N_7259,N_6895,N_6598);
nor U7260 (N_7260,N_6836,N_6573);
and U7261 (N_7261,N_6135,N_6149);
and U7262 (N_7262,N_6957,N_6197);
or U7263 (N_7263,N_6785,N_6022);
and U7264 (N_7264,N_6281,N_6922);
nor U7265 (N_7265,N_6484,N_6756);
nand U7266 (N_7266,N_6246,N_6544);
nor U7267 (N_7267,N_6307,N_6940);
nand U7268 (N_7268,N_6427,N_6955);
nand U7269 (N_7269,N_6440,N_6702);
nand U7270 (N_7270,N_6819,N_6816);
or U7271 (N_7271,N_6684,N_6931);
nor U7272 (N_7272,N_6031,N_6569);
nor U7273 (N_7273,N_6572,N_6333);
nor U7274 (N_7274,N_6983,N_6561);
nor U7275 (N_7275,N_6795,N_6750);
or U7276 (N_7276,N_6565,N_6039);
and U7277 (N_7277,N_6348,N_6265);
and U7278 (N_7278,N_6889,N_6508);
nand U7279 (N_7279,N_6524,N_6240);
or U7280 (N_7280,N_6141,N_6982);
nor U7281 (N_7281,N_6730,N_6734);
or U7282 (N_7282,N_6442,N_6831);
nand U7283 (N_7283,N_6391,N_6824);
nor U7284 (N_7284,N_6783,N_6044);
and U7285 (N_7285,N_6051,N_6993);
and U7286 (N_7286,N_6905,N_6509);
nor U7287 (N_7287,N_6064,N_6453);
nand U7288 (N_7288,N_6158,N_6639);
nor U7289 (N_7289,N_6751,N_6272);
or U7290 (N_7290,N_6111,N_6193);
nor U7291 (N_7291,N_6933,N_6784);
or U7292 (N_7292,N_6334,N_6627);
and U7293 (N_7293,N_6591,N_6306);
nor U7294 (N_7294,N_6489,N_6454);
or U7295 (N_7295,N_6710,N_6539);
or U7296 (N_7296,N_6855,N_6117);
nand U7297 (N_7297,N_6293,N_6266);
nor U7298 (N_7298,N_6705,N_6536);
nand U7299 (N_7299,N_6302,N_6204);
or U7300 (N_7300,N_6762,N_6107);
nor U7301 (N_7301,N_6495,N_6361);
or U7302 (N_7302,N_6457,N_6615);
nor U7303 (N_7303,N_6614,N_6167);
nand U7304 (N_7304,N_6566,N_6365);
and U7305 (N_7305,N_6385,N_6451);
or U7306 (N_7306,N_6187,N_6507);
nor U7307 (N_7307,N_6179,N_6275);
or U7308 (N_7308,N_6199,N_6672);
and U7309 (N_7309,N_6606,N_6422);
or U7310 (N_7310,N_6770,N_6185);
nor U7311 (N_7311,N_6386,N_6767);
nor U7312 (N_7312,N_6220,N_6588);
nor U7313 (N_7313,N_6568,N_6786);
nand U7314 (N_7314,N_6680,N_6472);
nand U7315 (N_7315,N_6328,N_6567);
or U7316 (N_7316,N_6636,N_6769);
and U7317 (N_7317,N_6976,N_6148);
nor U7318 (N_7318,N_6192,N_6131);
nor U7319 (N_7319,N_6349,N_6009);
and U7320 (N_7320,N_6708,N_6020);
and U7321 (N_7321,N_6099,N_6127);
or U7322 (N_7322,N_6369,N_6746);
or U7323 (N_7323,N_6570,N_6463);
nand U7324 (N_7324,N_6842,N_6313);
and U7325 (N_7325,N_6981,N_6942);
nand U7326 (N_7326,N_6262,N_6023);
or U7327 (N_7327,N_6582,N_6058);
and U7328 (N_7328,N_6236,N_6438);
and U7329 (N_7329,N_6635,N_6758);
or U7330 (N_7330,N_6552,N_6835);
and U7331 (N_7331,N_6972,N_6059);
and U7332 (N_7332,N_6415,N_6402);
nor U7333 (N_7333,N_6690,N_6285);
nor U7334 (N_7334,N_6355,N_6820);
and U7335 (N_7335,N_6213,N_6177);
or U7336 (N_7336,N_6287,N_6006);
and U7337 (N_7337,N_6946,N_6305);
or U7338 (N_7338,N_6695,N_6988);
or U7339 (N_7339,N_6317,N_6279);
nand U7340 (N_7340,N_6643,N_6482);
nor U7341 (N_7341,N_6480,N_6445);
and U7342 (N_7342,N_6460,N_6973);
and U7343 (N_7343,N_6393,N_6090);
and U7344 (N_7344,N_6502,N_6956);
nand U7345 (N_7345,N_6927,N_6258);
nor U7346 (N_7346,N_6493,N_6551);
nor U7347 (N_7347,N_6430,N_6011);
or U7348 (N_7348,N_6224,N_6410);
nor U7349 (N_7349,N_6880,N_6282);
nor U7350 (N_7350,N_6252,N_6712);
nor U7351 (N_7351,N_6601,N_6247);
or U7352 (N_7352,N_6304,N_6163);
nand U7353 (N_7353,N_6219,N_6733);
and U7354 (N_7354,N_6170,N_6741);
nor U7355 (N_7355,N_6392,N_6803);
nand U7356 (N_7356,N_6950,N_6425);
nor U7357 (N_7357,N_6632,N_6805);
xnor U7358 (N_7358,N_6292,N_6514);
nand U7359 (N_7359,N_6013,N_6704);
nor U7360 (N_7360,N_6491,N_6679);
nand U7361 (N_7361,N_6822,N_6418);
and U7362 (N_7362,N_6584,N_6299);
or U7363 (N_7363,N_6745,N_6876);
or U7364 (N_7364,N_6755,N_6826);
nor U7365 (N_7365,N_6235,N_6958);
or U7366 (N_7366,N_6060,N_6998);
nor U7367 (N_7367,N_6662,N_6818);
and U7368 (N_7368,N_6631,N_6142);
and U7369 (N_7369,N_6320,N_6732);
or U7370 (N_7370,N_6470,N_6587);
and U7371 (N_7371,N_6944,N_6359);
nand U7372 (N_7372,N_6503,N_6481);
and U7373 (N_7373,N_6325,N_6626);
nor U7374 (N_7374,N_6760,N_6095);
nor U7375 (N_7375,N_6071,N_6629);
nor U7376 (N_7376,N_6368,N_6471);
and U7377 (N_7377,N_6356,N_6864);
or U7378 (N_7378,N_6871,N_6687);
nand U7379 (N_7379,N_6375,N_6658);
nor U7380 (N_7380,N_6115,N_6342);
and U7381 (N_7381,N_6056,N_6108);
and U7382 (N_7382,N_6233,N_6053);
and U7383 (N_7383,N_6555,N_6226);
nor U7384 (N_7384,N_6676,N_6677);
nand U7385 (N_7385,N_6173,N_6161);
nand U7386 (N_7386,N_6622,N_6737);
and U7387 (N_7387,N_6209,N_6000);
or U7388 (N_7388,N_6140,N_6882);
nand U7389 (N_7389,N_6542,N_6186);
nor U7390 (N_7390,N_6449,N_6752);
and U7391 (N_7391,N_6902,N_6494);
or U7392 (N_7392,N_6531,N_6194);
or U7393 (N_7393,N_6323,N_6473);
nand U7394 (N_7394,N_6915,N_6370);
or U7395 (N_7395,N_6911,N_6711);
nor U7396 (N_7396,N_6707,N_6082);
and U7397 (N_7397,N_6421,N_6351);
and U7398 (N_7398,N_6674,N_6693);
nand U7399 (N_7399,N_6553,N_6799);
or U7400 (N_7400,N_6467,N_6772);
or U7401 (N_7401,N_6466,N_6335);
and U7402 (N_7402,N_6446,N_6346);
nand U7403 (N_7403,N_6088,N_6599);
nor U7404 (N_7404,N_6047,N_6678);
or U7405 (N_7405,N_6706,N_6229);
and U7406 (N_7406,N_6007,N_6874);
nand U7407 (N_7407,N_6448,N_6593);
and U7408 (N_7408,N_6404,N_6815);
nor U7409 (N_7409,N_6379,N_6154);
and U7410 (N_7410,N_6904,N_6309);
nor U7411 (N_7411,N_6465,N_6499);
or U7412 (N_7412,N_6653,N_6953);
or U7413 (N_7413,N_6806,N_6086);
or U7414 (N_7414,N_6137,N_6464);
and U7415 (N_7415,N_6119,N_6807);
nor U7416 (N_7416,N_6655,N_6890);
or U7417 (N_7417,N_6239,N_6104);
xnor U7418 (N_7418,N_6138,N_6830);
nand U7419 (N_7419,N_6268,N_6182);
and U7420 (N_7420,N_6352,N_6533);
nor U7421 (N_7421,N_6562,N_6439);
nor U7422 (N_7422,N_6537,N_6654);
nor U7423 (N_7423,N_6183,N_6435);
nand U7424 (N_7424,N_6885,N_6900);
nor U7425 (N_7425,N_6139,N_6101);
nand U7426 (N_7426,N_6867,N_6241);
nand U7427 (N_7427,N_6476,N_6003);
or U7428 (N_7428,N_6133,N_6002);
nor U7429 (N_7429,N_6248,N_6949);
nand U7430 (N_7430,N_6663,N_6560);
and U7431 (N_7431,N_6253,N_6657);
nand U7432 (N_7432,N_6479,N_6965);
and U7433 (N_7433,N_6564,N_6251);
nor U7434 (N_7434,N_6034,N_6319);
and U7435 (N_7435,N_6559,N_6877);
and U7436 (N_7436,N_6928,N_6719);
nor U7437 (N_7437,N_6276,N_6930);
and U7438 (N_7438,N_6670,N_6521);
nand U7439 (N_7439,N_6623,N_6130);
and U7440 (N_7440,N_6833,N_6963);
nand U7441 (N_7441,N_6980,N_6796);
nor U7442 (N_7442,N_6215,N_6578);
nor U7443 (N_7443,N_6543,N_6716);
nor U7444 (N_7444,N_6881,N_6124);
and U7445 (N_7445,N_6025,N_6967);
nor U7446 (N_7446,N_6892,N_6853);
or U7447 (N_7447,N_6078,N_6666);
or U7448 (N_7448,N_6390,N_6244);
nand U7449 (N_7449,N_6619,N_6329);
and U7450 (N_7450,N_6879,N_6943);
nor U7451 (N_7451,N_6028,N_6303);
or U7452 (N_7452,N_6122,N_6661);
nand U7453 (N_7453,N_6727,N_6070);
nor U7454 (N_7454,N_6611,N_6096);
or U7455 (N_7455,N_6225,N_6345);
or U7456 (N_7456,N_6894,N_6962);
or U7457 (N_7457,N_6350,N_6634);
and U7458 (N_7458,N_6701,N_6077);
nand U7459 (N_7459,N_6832,N_6651);
nor U7460 (N_7460,N_6736,N_6112);
nor U7461 (N_7461,N_6397,N_6638);
and U7462 (N_7462,N_6913,N_6620);
and U7463 (N_7463,N_6164,N_6277);
or U7464 (N_7464,N_6324,N_6563);
and U7465 (N_7465,N_6790,N_6260);
and U7466 (N_7466,N_6801,N_6176);
and U7467 (N_7467,N_6156,N_6999);
or U7468 (N_7468,N_6029,N_6057);
nor U7469 (N_7469,N_6637,N_6590);
and U7470 (N_7470,N_6910,N_6381);
and U7471 (N_7471,N_6267,N_6789);
and U7472 (N_7472,N_6061,N_6726);
nand U7473 (N_7473,N_6286,N_6725);
and U7474 (N_7474,N_6969,N_6227);
nand U7475 (N_7475,N_6813,N_6316);
nor U7476 (N_7476,N_6744,N_6550);
nor U7477 (N_7477,N_6169,N_6103);
nor U7478 (N_7478,N_6511,N_6496);
or U7479 (N_7479,N_6990,N_6989);
or U7480 (N_7480,N_6579,N_6032);
or U7481 (N_7481,N_6671,N_6443);
nor U7482 (N_7482,N_6237,N_6740);
nor U7483 (N_7483,N_6145,N_6123);
and U7484 (N_7484,N_6255,N_6214);
and U7485 (N_7485,N_6098,N_6974);
and U7486 (N_7486,N_6844,N_6420);
xnor U7487 (N_7487,N_6469,N_6121);
nor U7488 (N_7488,N_6576,N_6076);
nor U7489 (N_7489,N_6147,N_6925);
nor U7490 (N_7490,N_6206,N_6387);
and U7491 (N_7491,N_6015,N_6888);
or U7492 (N_7492,N_6245,N_6914);
or U7493 (N_7493,N_6921,N_6665);
nand U7494 (N_7494,N_6817,N_6574);
nor U7495 (N_7495,N_6628,N_6609);
nand U7496 (N_7496,N_6683,N_6617);
xnor U7497 (N_7497,N_6165,N_6301);
nand U7498 (N_7498,N_6019,N_6968);
nand U7499 (N_7499,N_6419,N_6280);
or U7500 (N_7500,N_6662,N_6848);
and U7501 (N_7501,N_6371,N_6894);
nand U7502 (N_7502,N_6480,N_6113);
nand U7503 (N_7503,N_6902,N_6137);
nand U7504 (N_7504,N_6139,N_6687);
nand U7505 (N_7505,N_6667,N_6488);
nand U7506 (N_7506,N_6247,N_6220);
and U7507 (N_7507,N_6201,N_6704);
and U7508 (N_7508,N_6764,N_6278);
and U7509 (N_7509,N_6231,N_6879);
nand U7510 (N_7510,N_6499,N_6741);
nand U7511 (N_7511,N_6321,N_6918);
nand U7512 (N_7512,N_6773,N_6959);
and U7513 (N_7513,N_6069,N_6350);
or U7514 (N_7514,N_6554,N_6199);
nor U7515 (N_7515,N_6960,N_6279);
and U7516 (N_7516,N_6585,N_6395);
nor U7517 (N_7517,N_6549,N_6987);
or U7518 (N_7518,N_6198,N_6803);
and U7519 (N_7519,N_6329,N_6916);
or U7520 (N_7520,N_6131,N_6716);
and U7521 (N_7521,N_6498,N_6090);
nand U7522 (N_7522,N_6984,N_6326);
or U7523 (N_7523,N_6893,N_6295);
nand U7524 (N_7524,N_6157,N_6381);
and U7525 (N_7525,N_6836,N_6718);
and U7526 (N_7526,N_6532,N_6594);
nor U7527 (N_7527,N_6740,N_6250);
or U7528 (N_7528,N_6935,N_6074);
and U7529 (N_7529,N_6769,N_6152);
nor U7530 (N_7530,N_6460,N_6539);
or U7531 (N_7531,N_6594,N_6916);
or U7532 (N_7532,N_6798,N_6928);
nor U7533 (N_7533,N_6841,N_6743);
nor U7534 (N_7534,N_6376,N_6587);
nand U7535 (N_7535,N_6554,N_6010);
nand U7536 (N_7536,N_6508,N_6059);
and U7537 (N_7537,N_6578,N_6366);
or U7538 (N_7538,N_6767,N_6666);
or U7539 (N_7539,N_6202,N_6514);
or U7540 (N_7540,N_6265,N_6409);
xnor U7541 (N_7541,N_6703,N_6023);
nand U7542 (N_7542,N_6581,N_6304);
nor U7543 (N_7543,N_6309,N_6467);
and U7544 (N_7544,N_6988,N_6555);
and U7545 (N_7545,N_6590,N_6596);
and U7546 (N_7546,N_6971,N_6818);
nand U7547 (N_7547,N_6800,N_6199);
nand U7548 (N_7548,N_6826,N_6041);
nand U7549 (N_7549,N_6347,N_6001);
and U7550 (N_7550,N_6067,N_6631);
nor U7551 (N_7551,N_6695,N_6002);
or U7552 (N_7552,N_6148,N_6274);
nor U7553 (N_7553,N_6571,N_6121);
nor U7554 (N_7554,N_6246,N_6418);
or U7555 (N_7555,N_6043,N_6913);
nand U7556 (N_7556,N_6606,N_6152);
and U7557 (N_7557,N_6968,N_6198);
and U7558 (N_7558,N_6909,N_6102);
nor U7559 (N_7559,N_6241,N_6638);
nor U7560 (N_7560,N_6503,N_6914);
nor U7561 (N_7561,N_6734,N_6545);
and U7562 (N_7562,N_6927,N_6902);
and U7563 (N_7563,N_6761,N_6766);
or U7564 (N_7564,N_6131,N_6017);
or U7565 (N_7565,N_6108,N_6595);
nor U7566 (N_7566,N_6155,N_6777);
and U7567 (N_7567,N_6010,N_6342);
nor U7568 (N_7568,N_6726,N_6293);
or U7569 (N_7569,N_6937,N_6468);
nor U7570 (N_7570,N_6780,N_6642);
nand U7571 (N_7571,N_6660,N_6263);
or U7572 (N_7572,N_6848,N_6576);
and U7573 (N_7573,N_6427,N_6931);
and U7574 (N_7574,N_6792,N_6396);
nand U7575 (N_7575,N_6541,N_6005);
nand U7576 (N_7576,N_6077,N_6856);
nand U7577 (N_7577,N_6276,N_6620);
and U7578 (N_7578,N_6663,N_6581);
nand U7579 (N_7579,N_6541,N_6247);
and U7580 (N_7580,N_6068,N_6079);
nor U7581 (N_7581,N_6243,N_6931);
nor U7582 (N_7582,N_6874,N_6981);
or U7583 (N_7583,N_6016,N_6989);
and U7584 (N_7584,N_6612,N_6984);
or U7585 (N_7585,N_6938,N_6498);
nand U7586 (N_7586,N_6575,N_6769);
and U7587 (N_7587,N_6641,N_6381);
and U7588 (N_7588,N_6032,N_6360);
nor U7589 (N_7589,N_6678,N_6241);
or U7590 (N_7590,N_6419,N_6126);
and U7591 (N_7591,N_6528,N_6130);
and U7592 (N_7592,N_6053,N_6770);
nand U7593 (N_7593,N_6977,N_6685);
or U7594 (N_7594,N_6646,N_6345);
or U7595 (N_7595,N_6813,N_6843);
or U7596 (N_7596,N_6064,N_6528);
nor U7597 (N_7597,N_6039,N_6122);
nor U7598 (N_7598,N_6140,N_6117);
or U7599 (N_7599,N_6063,N_6941);
nor U7600 (N_7600,N_6066,N_6403);
or U7601 (N_7601,N_6987,N_6211);
nand U7602 (N_7602,N_6747,N_6606);
nor U7603 (N_7603,N_6197,N_6368);
and U7604 (N_7604,N_6262,N_6265);
or U7605 (N_7605,N_6103,N_6959);
and U7606 (N_7606,N_6277,N_6244);
and U7607 (N_7607,N_6591,N_6940);
nor U7608 (N_7608,N_6316,N_6847);
nand U7609 (N_7609,N_6748,N_6362);
and U7610 (N_7610,N_6975,N_6295);
or U7611 (N_7611,N_6518,N_6530);
and U7612 (N_7612,N_6979,N_6099);
nand U7613 (N_7613,N_6358,N_6846);
or U7614 (N_7614,N_6059,N_6725);
and U7615 (N_7615,N_6963,N_6703);
nor U7616 (N_7616,N_6255,N_6817);
nand U7617 (N_7617,N_6003,N_6619);
and U7618 (N_7618,N_6566,N_6643);
and U7619 (N_7619,N_6965,N_6998);
and U7620 (N_7620,N_6240,N_6377);
nor U7621 (N_7621,N_6053,N_6541);
nand U7622 (N_7622,N_6294,N_6522);
nor U7623 (N_7623,N_6665,N_6866);
and U7624 (N_7624,N_6086,N_6350);
or U7625 (N_7625,N_6371,N_6477);
nor U7626 (N_7626,N_6809,N_6024);
and U7627 (N_7627,N_6692,N_6613);
nor U7628 (N_7628,N_6012,N_6023);
and U7629 (N_7629,N_6556,N_6625);
nand U7630 (N_7630,N_6752,N_6689);
nor U7631 (N_7631,N_6002,N_6209);
and U7632 (N_7632,N_6726,N_6535);
and U7633 (N_7633,N_6823,N_6039);
nor U7634 (N_7634,N_6111,N_6002);
nand U7635 (N_7635,N_6338,N_6434);
nor U7636 (N_7636,N_6778,N_6993);
and U7637 (N_7637,N_6842,N_6962);
nand U7638 (N_7638,N_6113,N_6145);
and U7639 (N_7639,N_6593,N_6602);
and U7640 (N_7640,N_6856,N_6582);
and U7641 (N_7641,N_6231,N_6178);
nor U7642 (N_7642,N_6603,N_6834);
and U7643 (N_7643,N_6205,N_6102);
nand U7644 (N_7644,N_6818,N_6428);
or U7645 (N_7645,N_6564,N_6856);
nand U7646 (N_7646,N_6296,N_6006);
and U7647 (N_7647,N_6240,N_6009);
nor U7648 (N_7648,N_6096,N_6702);
nor U7649 (N_7649,N_6300,N_6145);
and U7650 (N_7650,N_6786,N_6053);
or U7651 (N_7651,N_6618,N_6247);
nand U7652 (N_7652,N_6383,N_6248);
nor U7653 (N_7653,N_6507,N_6351);
nand U7654 (N_7654,N_6086,N_6437);
and U7655 (N_7655,N_6109,N_6254);
or U7656 (N_7656,N_6825,N_6198);
or U7657 (N_7657,N_6586,N_6557);
nor U7658 (N_7658,N_6776,N_6329);
nor U7659 (N_7659,N_6710,N_6735);
and U7660 (N_7660,N_6391,N_6389);
or U7661 (N_7661,N_6880,N_6990);
nand U7662 (N_7662,N_6290,N_6960);
nor U7663 (N_7663,N_6626,N_6989);
and U7664 (N_7664,N_6238,N_6518);
nor U7665 (N_7665,N_6297,N_6733);
nor U7666 (N_7666,N_6457,N_6001);
or U7667 (N_7667,N_6636,N_6491);
nand U7668 (N_7668,N_6950,N_6244);
nor U7669 (N_7669,N_6668,N_6798);
nand U7670 (N_7670,N_6865,N_6786);
nand U7671 (N_7671,N_6175,N_6411);
or U7672 (N_7672,N_6187,N_6362);
nor U7673 (N_7673,N_6093,N_6526);
or U7674 (N_7674,N_6779,N_6006);
and U7675 (N_7675,N_6810,N_6491);
nand U7676 (N_7676,N_6223,N_6259);
or U7677 (N_7677,N_6130,N_6173);
nor U7678 (N_7678,N_6803,N_6094);
or U7679 (N_7679,N_6124,N_6700);
nor U7680 (N_7680,N_6615,N_6927);
nor U7681 (N_7681,N_6065,N_6980);
or U7682 (N_7682,N_6745,N_6113);
or U7683 (N_7683,N_6931,N_6766);
or U7684 (N_7684,N_6502,N_6242);
or U7685 (N_7685,N_6046,N_6610);
or U7686 (N_7686,N_6697,N_6971);
nand U7687 (N_7687,N_6466,N_6947);
and U7688 (N_7688,N_6662,N_6672);
nor U7689 (N_7689,N_6839,N_6880);
and U7690 (N_7690,N_6654,N_6897);
nor U7691 (N_7691,N_6053,N_6969);
or U7692 (N_7692,N_6549,N_6648);
and U7693 (N_7693,N_6726,N_6193);
nor U7694 (N_7694,N_6233,N_6019);
nand U7695 (N_7695,N_6802,N_6450);
nand U7696 (N_7696,N_6985,N_6791);
and U7697 (N_7697,N_6618,N_6791);
and U7698 (N_7698,N_6058,N_6362);
or U7699 (N_7699,N_6570,N_6853);
and U7700 (N_7700,N_6603,N_6496);
nand U7701 (N_7701,N_6208,N_6784);
nor U7702 (N_7702,N_6113,N_6378);
or U7703 (N_7703,N_6365,N_6831);
and U7704 (N_7704,N_6690,N_6833);
nand U7705 (N_7705,N_6934,N_6183);
or U7706 (N_7706,N_6881,N_6370);
and U7707 (N_7707,N_6461,N_6944);
and U7708 (N_7708,N_6089,N_6392);
nor U7709 (N_7709,N_6703,N_6126);
nor U7710 (N_7710,N_6496,N_6219);
or U7711 (N_7711,N_6722,N_6937);
nor U7712 (N_7712,N_6040,N_6693);
and U7713 (N_7713,N_6605,N_6865);
and U7714 (N_7714,N_6358,N_6753);
xor U7715 (N_7715,N_6226,N_6307);
nor U7716 (N_7716,N_6736,N_6320);
nor U7717 (N_7717,N_6071,N_6245);
and U7718 (N_7718,N_6567,N_6231);
nand U7719 (N_7719,N_6546,N_6019);
and U7720 (N_7720,N_6835,N_6719);
nor U7721 (N_7721,N_6278,N_6794);
or U7722 (N_7722,N_6949,N_6084);
or U7723 (N_7723,N_6468,N_6775);
or U7724 (N_7724,N_6110,N_6932);
nor U7725 (N_7725,N_6394,N_6859);
nor U7726 (N_7726,N_6687,N_6974);
nand U7727 (N_7727,N_6849,N_6026);
or U7728 (N_7728,N_6700,N_6189);
or U7729 (N_7729,N_6696,N_6290);
nand U7730 (N_7730,N_6005,N_6360);
or U7731 (N_7731,N_6616,N_6542);
and U7732 (N_7732,N_6424,N_6292);
or U7733 (N_7733,N_6545,N_6614);
and U7734 (N_7734,N_6089,N_6577);
or U7735 (N_7735,N_6724,N_6468);
and U7736 (N_7736,N_6968,N_6500);
and U7737 (N_7737,N_6295,N_6796);
nor U7738 (N_7738,N_6135,N_6100);
nor U7739 (N_7739,N_6623,N_6444);
nor U7740 (N_7740,N_6449,N_6118);
or U7741 (N_7741,N_6975,N_6806);
and U7742 (N_7742,N_6997,N_6601);
nand U7743 (N_7743,N_6488,N_6780);
nor U7744 (N_7744,N_6649,N_6288);
or U7745 (N_7745,N_6296,N_6500);
and U7746 (N_7746,N_6556,N_6125);
nand U7747 (N_7747,N_6309,N_6169);
or U7748 (N_7748,N_6712,N_6590);
and U7749 (N_7749,N_6139,N_6185);
and U7750 (N_7750,N_6659,N_6870);
nor U7751 (N_7751,N_6348,N_6295);
nor U7752 (N_7752,N_6595,N_6069);
nand U7753 (N_7753,N_6158,N_6894);
and U7754 (N_7754,N_6052,N_6327);
nor U7755 (N_7755,N_6187,N_6729);
and U7756 (N_7756,N_6033,N_6869);
nor U7757 (N_7757,N_6662,N_6751);
and U7758 (N_7758,N_6407,N_6527);
and U7759 (N_7759,N_6086,N_6828);
nor U7760 (N_7760,N_6442,N_6179);
nor U7761 (N_7761,N_6165,N_6769);
and U7762 (N_7762,N_6100,N_6431);
nor U7763 (N_7763,N_6974,N_6864);
nand U7764 (N_7764,N_6218,N_6702);
nand U7765 (N_7765,N_6452,N_6634);
nor U7766 (N_7766,N_6631,N_6508);
and U7767 (N_7767,N_6682,N_6225);
nor U7768 (N_7768,N_6002,N_6722);
or U7769 (N_7769,N_6274,N_6301);
and U7770 (N_7770,N_6850,N_6951);
nand U7771 (N_7771,N_6793,N_6306);
nor U7772 (N_7772,N_6418,N_6804);
nor U7773 (N_7773,N_6440,N_6550);
or U7774 (N_7774,N_6361,N_6210);
nor U7775 (N_7775,N_6675,N_6222);
or U7776 (N_7776,N_6251,N_6048);
and U7777 (N_7777,N_6543,N_6225);
nand U7778 (N_7778,N_6290,N_6468);
or U7779 (N_7779,N_6202,N_6387);
and U7780 (N_7780,N_6237,N_6735);
nor U7781 (N_7781,N_6649,N_6507);
nand U7782 (N_7782,N_6361,N_6998);
or U7783 (N_7783,N_6777,N_6419);
nor U7784 (N_7784,N_6857,N_6978);
and U7785 (N_7785,N_6871,N_6050);
nand U7786 (N_7786,N_6161,N_6736);
nand U7787 (N_7787,N_6016,N_6025);
nand U7788 (N_7788,N_6541,N_6088);
nor U7789 (N_7789,N_6780,N_6312);
nand U7790 (N_7790,N_6660,N_6487);
and U7791 (N_7791,N_6210,N_6673);
nor U7792 (N_7792,N_6427,N_6204);
nor U7793 (N_7793,N_6828,N_6461);
nor U7794 (N_7794,N_6156,N_6023);
xnor U7795 (N_7795,N_6744,N_6075);
and U7796 (N_7796,N_6177,N_6576);
nor U7797 (N_7797,N_6024,N_6071);
and U7798 (N_7798,N_6202,N_6025);
nor U7799 (N_7799,N_6830,N_6534);
nand U7800 (N_7800,N_6171,N_6316);
and U7801 (N_7801,N_6932,N_6774);
or U7802 (N_7802,N_6900,N_6874);
nand U7803 (N_7803,N_6324,N_6421);
and U7804 (N_7804,N_6265,N_6453);
nor U7805 (N_7805,N_6386,N_6576);
or U7806 (N_7806,N_6243,N_6271);
nor U7807 (N_7807,N_6393,N_6917);
and U7808 (N_7808,N_6299,N_6761);
nand U7809 (N_7809,N_6349,N_6698);
nor U7810 (N_7810,N_6102,N_6311);
or U7811 (N_7811,N_6601,N_6740);
and U7812 (N_7812,N_6768,N_6322);
and U7813 (N_7813,N_6282,N_6031);
nand U7814 (N_7814,N_6098,N_6308);
or U7815 (N_7815,N_6774,N_6702);
nand U7816 (N_7816,N_6175,N_6513);
nor U7817 (N_7817,N_6069,N_6707);
or U7818 (N_7818,N_6413,N_6950);
xnor U7819 (N_7819,N_6421,N_6970);
and U7820 (N_7820,N_6944,N_6706);
and U7821 (N_7821,N_6387,N_6885);
and U7822 (N_7822,N_6931,N_6018);
nor U7823 (N_7823,N_6744,N_6886);
nand U7824 (N_7824,N_6238,N_6393);
nor U7825 (N_7825,N_6734,N_6616);
and U7826 (N_7826,N_6022,N_6003);
or U7827 (N_7827,N_6372,N_6146);
and U7828 (N_7828,N_6146,N_6377);
nand U7829 (N_7829,N_6989,N_6665);
nor U7830 (N_7830,N_6445,N_6515);
nor U7831 (N_7831,N_6031,N_6168);
nor U7832 (N_7832,N_6372,N_6855);
or U7833 (N_7833,N_6808,N_6537);
or U7834 (N_7834,N_6714,N_6116);
and U7835 (N_7835,N_6265,N_6443);
nand U7836 (N_7836,N_6034,N_6721);
nand U7837 (N_7837,N_6514,N_6618);
nand U7838 (N_7838,N_6135,N_6101);
and U7839 (N_7839,N_6874,N_6442);
or U7840 (N_7840,N_6954,N_6899);
nor U7841 (N_7841,N_6304,N_6840);
and U7842 (N_7842,N_6043,N_6669);
nor U7843 (N_7843,N_6421,N_6924);
or U7844 (N_7844,N_6110,N_6869);
nand U7845 (N_7845,N_6698,N_6718);
and U7846 (N_7846,N_6226,N_6105);
and U7847 (N_7847,N_6395,N_6207);
and U7848 (N_7848,N_6462,N_6667);
nand U7849 (N_7849,N_6022,N_6302);
and U7850 (N_7850,N_6707,N_6416);
nand U7851 (N_7851,N_6078,N_6773);
or U7852 (N_7852,N_6506,N_6341);
nand U7853 (N_7853,N_6941,N_6253);
nor U7854 (N_7854,N_6478,N_6372);
nand U7855 (N_7855,N_6517,N_6975);
and U7856 (N_7856,N_6582,N_6629);
and U7857 (N_7857,N_6292,N_6360);
nor U7858 (N_7858,N_6574,N_6617);
nand U7859 (N_7859,N_6005,N_6789);
or U7860 (N_7860,N_6524,N_6023);
and U7861 (N_7861,N_6460,N_6597);
or U7862 (N_7862,N_6648,N_6100);
nor U7863 (N_7863,N_6945,N_6708);
or U7864 (N_7864,N_6218,N_6732);
or U7865 (N_7865,N_6879,N_6706);
nor U7866 (N_7866,N_6676,N_6600);
or U7867 (N_7867,N_6070,N_6311);
nand U7868 (N_7868,N_6230,N_6246);
nor U7869 (N_7869,N_6478,N_6407);
or U7870 (N_7870,N_6186,N_6784);
nor U7871 (N_7871,N_6545,N_6728);
or U7872 (N_7872,N_6918,N_6605);
and U7873 (N_7873,N_6315,N_6939);
and U7874 (N_7874,N_6254,N_6608);
nand U7875 (N_7875,N_6423,N_6858);
nand U7876 (N_7876,N_6114,N_6848);
or U7877 (N_7877,N_6077,N_6086);
or U7878 (N_7878,N_6862,N_6005);
nor U7879 (N_7879,N_6446,N_6486);
nor U7880 (N_7880,N_6912,N_6584);
and U7881 (N_7881,N_6907,N_6804);
nand U7882 (N_7882,N_6225,N_6609);
nor U7883 (N_7883,N_6288,N_6602);
nor U7884 (N_7884,N_6131,N_6363);
nor U7885 (N_7885,N_6829,N_6430);
nand U7886 (N_7886,N_6938,N_6317);
or U7887 (N_7887,N_6101,N_6417);
nand U7888 (N_7888,N_6575,N_6700);
nor U7889 (N_7889,N_6465,N_6119);
nand U7890 (N_7890,N_6532,N_6266);
and U7891 (N_7891,N_6805,N_6039);
nand U7892 (N_7892,N_6343,N_6631);
nand U7893 (N_7893,N_6286,N_6990);
or U7894 (N_7894,N_6949,N_6538);
nor U7895 (N_7895,N_6105,N_6633);
nor U7896 (N_7896,N_6482,N_6944);
and U7897 (N_7897,N_6207,N_6675);
and U7898 (N_7898,N_6894,N_6147);
and U7899 (N_7899,N_6731,N_6732);
nor U7900 (N_7900,N_6487,N_6122);
nor U7901 (N_7901,N_6765,N_6892);
nor U7902 (N_7902,N_6975,N_6629);
and U7903 (N_7903,N_6253,N_6437);
nor U7904 (N_7904,N_6532,N_6780);
nor U7905 (N_7905,N_6812,N_6553);
and U7906 (N_7906,N_6558,N_6321);
nor U7907 (N_7907,N_6519,N_6430);
or U7908 (N_7908,N_6713,N_6136);
nor U7909 (N_7909,N_6141,N_6753);
or U7910 (N_7910,N_6695,N_6537);
and U7911 (N_7911,N_6247,N_6827);
and U7912 (N_7912,N_6055,N_6889);
nand U7913 (N_7913,N_6876,N_6049);
nor U7914 (N_7914,N_6894,N_6941);
or U7915 (N_7915,N_6431,N_6148);
or U7916 (N_7916,N_6579,N_6515);
nor U7917 (N_7917,N_6584,N_6159);
nand U7918 (N_7918,N_6826,N_6633);
or U7919 (N_7919,N_6072,N_6543);
and U7920 (N_7920,N_6526,N_6217);
nand U7921 (N_7921,N_6703,N_6850);
nand U7922 (N_7922,N_6552,N_6339);
nand U7923 (N_7923,N_6560,N_6847);
and U7924 (N_7924,N_6274,N_6074);
nand U7925 (N_7925,N_6121,N_6879);
nor U7926 (N_7926,N_6047,N_6823);
nor U7927 (N_7927,N_6624,N_6680);
nand U7928 (N_7928,N_6421,N_6636);
or U7929 (N_7929,N_6403,N_6234);
nor U7930 (N_7930,N_6234,N_6585);
nor U7931 (N_7931,N_6733,N_6187);
or U7932 (N_7932,N_6099,N_6255);
nor U7933 (N_7933,N_6694,N_6173);
and U7934 (N_7934,N_6828,N_6854);
or U7935 (N_7935,N_6561,N_6109);
nand U7936 (N_7936,N_6296,N_6075);
nor U7937 (N_7937,N_6613,N_6836);
nand U7938 (N_7938,N_6321,N_6488);
nor U7939 (N_7939,N_6729,N_6160);
or U7940 (N_7940,N_6311,N_6732);
and U7941 (N_7941,N_6368,N_6921);
or U7942 (N_7942,N_6430,N_6873);
or U7943 (N_7943,N_6715,N_6746);
nor U7944 (N_7944,N_6958,N_6628);
or U7945 (N_7945,N_6414,N_6670);
and U7946 (N_7946,N_6281,N_6522);
or U7947 (N_7947,N_6515,N_6325);
nand U7948 (N_7948,N_6715,N_6981);
and U7949 (N_7949,N_6464,N_6479);
nand U7950 (N_7950,N_6276,N_6343);
nor U7951 (N_7951,N_6712,N_6427);
nor U7952 (N_7952,N_6577,N_6142);
nand U7953 (N_7953,N_6356,N_6225);
nor U7954 (N_7954,N_6319,N_6465);
and U7955 (N_7955,N_6186,N_6797);
nor U7956 (N_7956,N_6295,N_6223);
nor U7957 (N_7957,N_6644,N_6937);
nor U7958 (N_7958,N_6387,N_6987);
nor U7959 (N_7959,N_6413,N_6925);
or U7960 (N_7960,N_6732,N_6299);
nor U7961 (N_7961,N_6880,N_6757);
and U7962 (N_7962,N_6247,N_6740);
nor U7963 (N_7963,N_6427,N_6710);
and U7964 (N_7964,N_6657,N_6370);
and U7965 (N_7965,N_6344,N_6562);
and U7966 (N_7966,N_6422,N_6121);
nor U7967 (N_7967,N_6780,N_6049);
nor U7968 (N_7968,N_6339,N_6026);
nand U7969 (N_7969,N_6125,N_6582);
nor U7970 (N_7970,N_6220,N_6317);
nor U7971 (N_7971,N_6710,N_6915);
and U7972 (N_7972,N_6551,N_6246);
nand U7973 (N_7973,N_6617,N_6687);
nand U7974 (N_7974,N_6428,N_6295);
nand U7975 (N_7975,N_6078,N_6256);
nor U7976 (N_7976,N_6340,N_6791);
and U7977 (N_7977,N_6425,N_6850);
nand U7978 (N_7978,N_6193,N_6435);
nand U7979 (N_7979,N_6278,N_6038);
nor U7980 (N_7980,N_6524,N_6125);
or U7981 (N_7981,N_6857,N_6832);
nand U7982 (N_7982,N_6471,N_6323);
nand U7983 (N_7983,N_6241,N_6665);
and U7984 (N_7984,N_6385,N_6924);
or U7985 (N_7985,N_6071,N_6981);
or U7986 (N_7986,N_6919,N_6249);
nor U7987 (N_7987,N_6493,N_6625);
or U7988 (N_7988,N_6645,N_6681);
and U7989 (N_7989,N_6777,N_6200);
nand U7990 (N_7990,N_6821,N_6725);
xor U7991 (N_7991,N_6120,N_6738);
or U7992 (N_7992,N_6939,N_6274);
or U7993 (N_7993,N_6247,N_6061);
nand U7994 (N_7994,N_6559,N_6564);
or U7995 (N_7995,N_6424,N_6825);
nor U7996 (N_7996,N_6843,N_6419);
or U7997 (N_7997,N_6038,N_6560);
nand U7998 (N_7998,N_6753,N_6647);
or U7999 (N_7999,N_6077,N_6019);
nor U8000 (N_8000,N_7107,N_7056);
or U8001 (N_8001,N_7766,N_7287);
nand U8002 (N_8002,N_7232,N_7020);
and U8003 (N_8003,N_7743,N_7532);
and U8004 (N_8004,N_7045,N_7952);
and U8005 (N_8005,N_7876,N_7350);
nor U8006 (N_8006,N_7471,N_7327);
nor U8007 (N_8007,N_7799,N_7758);
nand U8008 (N_8008,N_7230,N_7291);
nor U8009 (N_8009,N_7523,N_7186);
nand U8010 (N_8010,N_7535,N_7326);
nor U8011 (N_8011,N_7409,N_7256);
or U8012 (N_8012,N_7832,N_7813);
and U8013 (N_8013,N_7285,N_7501);
or U8014 (N_8014,N_7640,N_7600);
nand U8015 (N_8015,N_7863,N_7564);
xor U8016 (N_8016,N_7652,N_7148);
or U8017 (N_8017,N_7774,N_7831);
and U8018 (N_8018,N_7916,N_7092);
or U8019 (N_8019,N_7996,N_7764);
or U8020 (N_8020,N_7777,N_7142);
nor U8021 (N_8021,N_7354,N_7245);
and U8022 (N_8022,N_7982,N_7980);
and U8023 (N_8023,N_7599,N_7117);
nand U8024 (N_8024,N_7431,N_7448);
and U8025 (N_8025,N_7626,N_7132);
and U8026 (N_8026,N_7641,N_7836);
nand U8027 (N_8027,N_7006,N_7397);
and U8028 (N_8028,N_7096,N_7457);
and U8029 (N_8029,N_7213,N_7218);
or U8030 (N_8030,N_7054,N_7234);
or U8031 (N_8031,N_7243,N_7637);
nand U8032 (N_8032,N_7377,N_7533);
and U8033 (N_8033,N_7417,N_7169);
nand U8034 (N_8034,N_7461,N_7469);
or U8035 (N_8035,N_7322,N_7144);
and U8036 (N_8036,N_7864,N_7769);
or U8037 (N_8037,N_7792,N_7375);
nor U8038 (N_8038,N_7435,N_7429);
and U8039 (N_8039,N_7536,N_7210);
and U8040 (N_8040,N_7882,N_7833);
and U8041 (N_8041,N_7085,N_7805);
and U8042 (N_8042,N_7602,N_7166);
nand U8043 (N_8043,N_7353,N_7058);
nor U8044 (N_8044,N_7632,N_7046);
nor U8045 (N_8045,N_7221,N_7981);
or U8046 (N_8046,N_7992,N_7312);
or U8047 (N_8047,N_7951,N_7464);
or U8048 (N_8048,N_7752,N_7164);
nand U8049 (N_8049,N_7156,N_7502);
nor U8050 (N_8050,N_7986,N_7133);
nand U8051 (N_8051,N_7562,N_7699);
nand U8052 (N_8052,N_7781,N_7822);
nor U8053 (N_8053,N_7030,N_7360);
and U8054 (N_8054,N_7888,N_7177);
or U8055 (N_8055,N_7624,N_7499);
nand U8056 (N_8056,N_7715,N_7840);
nor U8057 (N_8057,N_7567,N_7378);
nand U8058 (N_8058,N_7609,N_7995);
nor U8059 (N_8059,N_7317,N_7630);
and U8060 (N_8060,N_7668,N_7627);
or U8061 (N_8061,N_7829,N_7505);
nand U8062 (N_8062,N_7519,N_7147);
nor U8063 (N_8063,N_7052,N_7563);
nor U8064 (N_8064,N_7154,N_7441);
or U8065 (N_8065,N_7479,N_7314);
nor U8066 (N_8066,N_7530,N_7733);
and U8067 (N_8067,N_7549,N_7239);
nand U8068 (N_8068,N_7347,N_7406);
nor U8069 (N_8069,N_7901,N_7428);
or U8070 (N_8070,N_7047,N_7800);
nor U8071 (N_8071,N_7442,N_7507);
or U8072 (N_8072,N_7659,N_7565);
nor U8073 (N_8073,N_7911,N_7797);
or U8074 (N_8074,N_7604,N_7925);
and U8075 (N_8075,N_7313,N_7427);
nor U8076 (N_8076,N_7012,N_7595);
nand U8077 (N_8077,N_7447,N_7947);
nand U8078 (N_8078,N_7454,N_7053);
and U8079 (N_8079,N_7828,N_7003);
and U8080 (N_8080,N_7987,N_7233);
and U8081 (N_8081,N_7124,N_7349);
nand U8082 (N_8082,N_7290,N_7954);
nand U8083 (N_8083,N_7773,N_7994);
and U8084 (N_8084,N_7513,N_7373);
nand U8085 (N_8085,N_7226,N_7212);
and U8086 (N_8086,N_7906,N_7979);
nand U8087 (N_8087,N_7491,N_7307);
and U8088 (N_8088,N_7810,N_7948);
nor U8089 (N_8089,N_7883,N_7645);
or U8090 (N_8090,N_7946,N_7500);
or U8091 (N_8091,N_7439,N_7618);
nor U8092 (N_8092,N_7008,N_7275);
xnor U8093 (N_8093,N_7255,N_7267);
and U8094 (N_8094,N_7517,N_7845);
or U8095 (N_8095,N_7975,N_7231);
nor U8096 (N_8096,N_7109,N_7685);
nand U8097 (N_8097,N_7286,N_7506);
nor U8098 (N_8098,N_7497,N_7136);
or U8099 (N_8099,N_7574,N_7735);
or U8100 (N_8100,N_7180,N_7190);
or U8101 (N_8101,N_7035,N_7859);
nor U8102 (N_8102,N_7049,N_7515);
and U8103 (N_8103,N_7712,N_7258);
or U8104 (N_8104,N_7744,N_7265);
nor U8105 (N_8105,N_7971,N_7250);
nand U8106 (N_8106,N_7896,N_7670);
or U8107 (N_8107,N_7129,N_7474);
and U8108 (N_8108,N_7485,N_7451);
or U8109 (N_8109,N_7698,N_7036);
nor U8110 (N_8110,N_7582,N_7550);
and U8111 (N_8111,N_7671,N_7208);
nor U8112 (N_8112,N_7912,N_7727);
or U8113 (N_8113,N_7319,N_7104);
or U8114 (N_8114,N_7650,N_7466);
nor U8115 (N_8115,N_7651,N_7097);
nor U8116 (N_8116,N_7108,N_7419);
or U8117 (N_8117,N_7592,N_7135);
or U8118 (N_8118,N_7498,N_7470);
nand U8119 (N_8119,N_7486,N_7615);
and U8120 (N_8120,N_7157,N_7811);
and U8121 (N_8121,N_7661,N_7426);
or U8122 (N_8122,N_7335,N_7696);
and U8123 (N_8123,N_7140,N_7934);
nor U8124 (N_8124,N_7207,N_7776);
nand U8125 (N_8125,N_7956,N_7689);
or U8126 (N_8126,N_7521,N_7666);
nor U8127 (N_8127,N_7063,N_7960);
or U8128 (N_8128,N_7083,N_7838);
or U8129 (N_8129,N_7669,N_7033);
or U8130 (N_8130,N_7029,N_7418);
and U8131 (N_8131,N_7588,N_7529);
and U8132 (N_8132,N_7543,N_7573);
nor U8133 (N_8133,N_7162,N_7939);
nor U8134 (N_8134,N_7134,N_7309);
nor U8135 (N_8135,N_7837,N_7824);
nand U8136 (N_8136,N_7711,N_7382);
nand U8137 (N_8137,N_7393,N_7988);
nor U8138 (N_8138,N_7344,N_7421);
nand U8139 (N_8139,N_7415,N_7205);
or U8140 (N_8140,N_7680,N_7511);
nand U8141 (N_8141,N_7779,N_7112);
nor U8142 (N_8142,N_7809,N_7569);
or U8143 (N_8143,N_7355,N_7293);
nor U8144 (N_8144,N_7961,N_7141);
nor U8145 (N_8145,N_7926,N_7551);
nor U8146 (N_8146,N_7333,N_7933);
nand U8147 (N_8147,N_7158,N_7178);
nand U8148 (N_8148,N_7062,N_7422);
nand U8149 (N_8149,N_7751,N_7620);
nand U8150 (N_8150,N_7363,N_7885);
and U8151 (N_8151,N_7560,N_7276);
nor U8152 (N_8152,N_7137,N_7197);
nor U8153 (N_8153,N_7189,N_7271);
nor U8154 (N_8154,N_7119,N_7289);
and U8155 (N_8155,N_7617,N_7789);
nor U8156 (N_8156,N_7238,N_7953);
or U8157 (N_8157,N_7855,N_7761);
nand U8158 (N_8158,N_7403,N_7907);
or U8159 (N_8159,N_7007,N_7115);
nor U8160 (N_8160,N_7930,N_7253);
and U8161 (N_8161,N_7940,N_7816);
nand U8162 (N_8162,N_7437,N_7379);
or U8163 (N_8163,N_7026,N_7941);
or U8164 (N_8164,N_7184,N_7942);
and U8165 (N_8165,N_7897,N_7522);
nand U8166 (N_8166,N_7042,N_7125);
nand U8167 (N_8167,N_7440,N_7893);
nand U8168 (N_8168,N_7346,N_7153);
nor U8169 (N_8169,N_7721,N_7913);
and U8170 (N_8170,N_7308,N_7202);
or U8171 (N_8171,N_7163,N_7796);
or U8172 (N_8172,N_7384,N_7443);
and U8173 (N_8173,N_7570,N_7316);
nand U8174 (N_8174,N_7358,N_7702);
nand U8175 (N_8175,N_7635,N_7890);
and U8176 (N_8176,N_7749,N_7420);
nand U8177 (N_8177,N_7552,N_7928);
and U8178 (N_8178,N_7264,N_7009);
and U8179 (N_8179,N_7955,N_7219);
nand U8180 (N_8180,N_7462,N_7572);
nor U8181 (N_8181,N_7667,N_7296);
and U8182 (N_8182,N_7100,N_7775);
or U8183 (N_8183,N_7581,N_7392);
nor U8184 (N_8184,N_7340,N_7705);
nand U8185 (N_8185,N_7639,N_7073);
and U8186 (N_8186,N_7410,N_7160);
nor U8187 (N_8187,N_7182,N_7084);
nand U8188 (N_8188,N_7895,N_7820);
nand U8189 (N_8189,N_7904,N_7405);
nand U8190 (N_8190,N_7222,N_7585);
or U8191 (N_8191,N_7694,N_7784);
nor U8192 (N_8192,N_7528,N_7539);
and U8193 (N_8193,N_7780,N_7606);
nor U8194 (N_8194,N_7116,N_7086);
or U8195 (N_8195,N_7962,N_7456);
and U8196 (N_8196,N_7731,N_7717);
nor U8197 (N_8197,N_7851,N_7217);
nor U8198 (N_8198,N_7983,N_7272);
nand U8199 (N_8199,N_7559,N_7648);
nor U8200 (N_8200,N_7959,N_7179);
nor U8201 (N_8201,N_7725,N_7806);
nand U8202 (N_8202,N_7692,N_7772);
and U8203 (N_8203,N_7311,N_7400);
or U8204 (N_8204,N_7587,N_7002);
and U8205 (N_8205,N_7050,N_7807);
or U8206 (N_8206,N_7057,N_7943);
and U8207 (N_8207,N_7937,N_7005);
nor U8208 (N_8208,N_7783,N_7646);
nor U8209 (N_8209,N_7077,N_7999);
nor U8210 (N_8210,N_7300,N_7873);
nand U8211 (N_8211,N_7282,N_7737);
nor U8212 (N_8212,N_7199,N_7345);
nand U8213 (N_8213,N_7281,N_7488);
or U8214 (N_8214,N_7191,N_7424);
and U8215 (N_8215,N_7338,N_7452);
nor U8216 (N_8216,N_7093,N_7066);
or U8217 (N_8217,N_7894,N_7388);
and U8218 (N_8218,N_7371,N_7544);
nand U8219 (N_8219,N_7608,N_7817);
nor U8220 (N_8220,N_7558,N_7802);
nor U8221 (N_8221,N_7173,N_7295);
xnor U8222 (N_8222,N_7803,N_7301);
nand U8223 (N_8223,N_7854,N_7143);
nor U8224 (N_8224,N_7459,N_7801);
and U8225 (N_8225,N_7328,N_7741);
and U8226 (N_8226,N_7525,N_7259);
or U8227 (N_8227,N_7788,N_7524);
nand U8228 (N_8228,N_7674,N_7174);
or U8229 (N_8229,N_7976,N_7188);
or U8230 (N_8230,N_7575,N_7763);
nand U8231 (N_8231,N_7554,N_7172);
nor U8232 (N_8232,N_7480,N_7181);
and U8233 (N_8233,N_7413,N_7938);
and U8234 (N_8234,N_7747,N_7019);
nand U8235 (N_8235,N_7915,N_7681);
nand U8236 (N_8236,N_7381,N_7654);
and U8237 (N_8237,N_7745,N_7075);
nand U8238 (N_8238,N_7481,N_7280);
nand U8239 (N_8239,N_7545,N_7923);
xnor U8240 (N_8240,N_7339,N_7254);
or U8241 (N_8241,N_7825,N_7849);
or U8242 (N_8242,N_7399,N_7483);
or U8243 (N_8243,N_7579,N_7204);
or U8244 (N_8244,N_7453,N_7734);
and U8245 (N_8245,N_7105,N_7446);
or U8246 (N_8246,N_7716,N_7819);
nand U8247 (N_8247,N_7682,N_7871);
nor U8248 (N_8248,N_7812,N_7623);
and U8249 (N_8249,N_7414,N_7677);
and U8250 (N_8250,N_7875,N_7138);
nand U8251 (N_8251,N_7880,N_7458);
nand U8252 (N_8252,N_7038,N_7298);
or U8253 (N_8253,N_7061,N_7161);
nand U8254 (N_8254,N_7324,N_7991);
nand U8255 (N_8255,N_7279,N_7631);
xnor U8256 (N_8256,N_7542,N_7114);
nor U8257 (N_8257,N_7611,N_7069);
nand U8258 (N_8258,N_7701,N_7847);
or U8259 (N_8259,N_7127,N_7103);
or U8260 (N_8260,N_7315,N_7430);
nand U8261 (N_8261,N_7843,N_7850);
or U8262 (N_8262,N_7887,N_7278);
and U8263 (N_8263,N_7768,N_7736);
nand U8264 (N_8264,N_7242,N_7868);
nor U8265 (N_8265,N_7059,N_7228);
nand U8266 (N_8266,N_7739,N_7357);
or U8267 (N_8267,N_7193,N_7998);
and U8268 (N_8268,N_7889,N_7706);
or U8269 (N_8269,N_7914,N_7957);
or U8270 (N_8270,N_7740,N_7770);
or U8271 (N_8271,N_7856,N_7438);
and U8272 (N_8272,N_7794,N_7589);
and U8273 (N_8273,N_7899,N_7978);
or U8274 (N_8274,N_7229,N_7593);
nand U8275 (N_8275,N_7274,N_7821);
or U8276 (N_8276,N_7455,N_7647);
or U8277 (N_8277,N_7936,N_7762);
nor U8278 (N_8278,N_7149,N_7472);
nand U8279 (N_8279,N_7935,N_7898);
nor U8280 (N_8280,N_7244,N_7055);
nor U8281 (N_8281,N_7755,N_7014);
or U8282 (N_8282,N_7621,N_7676);
or U8283 (N_8283,N_7321,N_7330);
and U8284 (N_8284,N_7703,N_7917);
or U8285 (N_8285,N_7015,N_7372);
and U8286 (N_8286,N_7607,N_7118);
and U8287 (N_8287,N_7016,N_7804);
xnor U8288 (N_8288,N_7918,N_7760);
nor U8289 (N_8289,N_7394,N_7071);
nand U8290 (N_8290,N_7336,N_7984);
or U8291 (N_8291,N_7476,N_7827);
nand U8292 (N_8292,N_7512,N_7842);
nor U8293 (N_8293,N_7288,N_7225);
nor U8294 (N_8294,N_7223,N_7432);
xor U8295 (N_8295,N_7067,N_7248);
or U8296 (N_8296,N_7629,N_7151);
nor U8297 (N_8297,N_7094,N_7150);
nor U8298 (N_8298,N_7700,N_7434);
or U8299 (N_8299,N_7969,N_7678);
and U8300 (N_8300,N_7765,N_7714);
nand U8301 (N_8301,N_7292,N_7080);
nor U8302 (N_8302,N_7929,N_7835);
and U8303 (N_8303,N_7060,N_7520);
nand U8304 (N_8304,N_7516,N_7538);
nor U8305 (N_8305,N_7892,N_7862);
nand U8306 (N_8306,N_7642,N_7089);
nor U8307 (N_8307,N_7237,N_7449);
or U8308 (N_8308,N_7852,N_7619);
or U8309 (N_8309,N_7380,N_7878);
nor U8310 (N_8310,N_7396,N_7398);
and U8311 (N_8311,N_7269,N_7070);
or U8312 (N_8312,N_7601,N_7710);
nand U8313 (N_8313,N_7302,N_7120);
and U8314 (N_8314,N_7341,N_7495);
nor U8315 (N_8315,N_7106,N_7920);
nor U8316 (N_8316,N_7910,N_7068);
nand U8317 (N_8317,N_7131,N_7509);
and U8318 (N_8318,N_7728,N_7860);
and U8319 (N_8319,N_7571,N_7908);
nor U8320 (N_8320,N_7098,N_7241);
nand U8321 (N_8321,N_7478,N_7660);
nor U8322 (N_8322,N_7556,N_7808);
nand U8323 (N_8323,N_7235,N_7924);
nand U8324 (N_8324,N_7465,N_7385);
or U8325 (N_8325,N_7277,N_7304);
nand U8326 (N_8326,N_7944,N_7407);
and U8327 (N_8327,N_7695,N_7081);
nor U8328 (N_8328,N_7622,N_7778);
or U8329 (N_8329,N_7257,N_7203);
nand U8330 (N_8330,N_7704,N_7331);
nand U8331 (N_8331,N_7099,N_7738);
nand U8332 (N_8332,N_7541,N_7260);
or U8333 (N_8333,N_7170,N_7320);
nand U8334 (N_8334,N_7266,N_7425);
nor U8335 (N_8335,N_7122,N_7433);
nand U8336 (N_8336,N_7369,N_7128);
nand U8337 (N_8337,N_7625,N_7356);
nor U8338 (N_8338,N_7795,N_7989);
nand U8339 (N_8339,N_7508,N_7310);
or U8340 (N_8340,N_7332,N_7548);
nand U8341 (N_8341,N_7171,N_7527);
nor U8342 (N_8342,N_7395,N_7101);
nand U8343 (N_8343,N_7598,N_7844);
and U8344 (N_8344,N_7964,N_7351);
nand U8345 (N_8345,N_7283,N_7482);
and U8346 (N_8346,N_7262,N_7473);
and U8347 (N_8347,N_7644,N_7510);
or U8348 (N_8348,N_7662,N_7201);
nand U8349 (N_8349,N_7401,N_7367);
nand U8350 (N_8350,N_7445,N_7436);
and U8351 (N_8351,N_7065,N_7963);
and U8352 (N_8352,N_7649,N_7683);
nor U8353 (N_8353,N_7475,N_7076);
or U8354 (N_8354,N_7412,N_7352);
or U8355 (N_8355,N_7633,N_7968);
and U8356 (N_8356,N_7823,N_7636);
or U8357 (N_8357,N_7787,N_7023);
nand U8358 (N_8358,N_7111,N_7224);
xnor U8359 (N_8359,N_7753,N_7130);
nor U8360 (N_8360,N_7663,N_7577);
or U8361 (N_8361,N_7489,N_7022);
nor U8362 (N_8362,N_7909,N_7493);
nand U8363 (N_8363,N_7997,N_7209);
or U8364 (N_8364,N_7043,N_7504);
nand U8365 (N_8365,N_7390,N_7653);
and U8366 (N_8366,N_7730,N_7616);
nor U8367 (N_8367,N_7553,N_7869);
nor U8368 (N_8368,N_7329,N_7113);
and U8369 (N_8369,N_7198,N_7757);
nor U8370 (N_8370,N_7168,N_7011);
nor U8371 (N_8371,N_7830,N_7672);
and U8372 (N_8372,N_7318,N_7546);
nor U8373 (N_8373,N_7323,N_7467);
or U8374 (N_8374,N_7534,N_7665);
nand U8375 (N_8375,N_7251,N_7759);
and U8376 (N_8376,N_7273,N_7826);
nand U8377 (N_8377,N_7927,N_7900);
nand U8378 (N_8378,N_7145,N_7690);
and U8379 (N_8379,N_7713,N_7246);
or U8380 (N_8380,N_7072,N_7684);
nor U8381 (N_8381,N_7000,N_7970);
and U8382 (N_8382,N_7922,N_7594);
nor U8383 (N_8383,N_7767,N_7343);
and U8384 (N_8384,N_7404,N_7634);
xor U8385 (N_8385,N_7958,N_7921);
and U8386 (N_8386,N_7884,N_7596);
or U8387 (N_8387,N_7110,N_7102);
nor U8388 (N_8388,N_7165,N_7366);
nand U8389 (N_8389,N_7965,N_7815);
and U8390 (N_8390,N_7643,N_7841);
xnor U8391 (N_8391,N_7487,N_7628);
and U8392 (N_8392,N_7919,N_7568);
nor U8393 (N_8393,N_7391,N_7610);
nor U8394 (N_8394,N_7790,N_7192);
nor U8395 (N_8395,N_7613,N_7603);
or U8396 (N_8396,N_7723,N_7656);
nor U8397 (N_8397,N_7268,N_7638);
nand U8398 (N_8398,N_7655,N_7614);
and U8399 (N_8399,N_7786,N_7748);
and U8400 (N_8400,N_7719,N_7051);
nor U8401 (N_8401,N_7902,N_7079);
nor U8402 (N_8402,N_7537,N_7612);
or U8403 (N_8403,N_7031,N_7708);
and U8404 (N_8404,N_7408,N_7041);
nand U8405 (N_8405,N_7756,N_7215);
nand U8406 (N_8406,N_7402,N_7793);
nand U8407 (N_8407,N_7870,N_7973);
and U8408 (N_8408,N_7249,N_7305);
nand U8409 (N_8409,N_7194,N_7966);
nand U8410 (N_8410,N_7196,N_7657);
nand U8411 (N_8411,N_7389,N_7879);
nand U8412 (N_8412,N_7095,N_7039);
nor U8413 (N_8413,N_7152,N_7306);
or U8414 (N_8414,N_7074,N_7949);
nand U8415 (N_8415,N_7746,N_7082);
or U8416 (N_8416,N_7200,N_7503);
or U8417 (N_8417,N_7123,N_7531);
nor U8418 (N_8418,N_7139,N_7416);
nor U8419 (N_8419,N_7028,N_7025);
and U8420 (N_8420,N_7021,N_7010);
nand U8421 (N_8421,N_7693,N_7270);
and U8422 (N_8422,N_7444,N_7048);
nand U8423 (N_8423,N_7557,N_7368);
nor U8424 (N_8424,N_7032,N_7468);
nor U8425 (N_8425,N_7342,N_7974);
nor U8426 (N_8426,N_7578,N_7175);
nor U8427 (N_8427,N_7865,N_7294);
nand U8428 (N_8428,N_7707,N_7364);
nor U8429 (N_8429,N_7018,N_7017);
nor U8430 (N_8430,N_7782,N_7566);
and U8431 (N_8431,N_7853,N_7176);
nor U8432 (N_8432,N_7463,N_7263);
nor U8433 (N_8433,N_7159,N_7686);
and U8434 (N_8434,N_7679,N_7903);
nand U8435 (N_8435,N_7460,N_7742);
nand U8436 (N_8436,N_7490,N_7881);
nand U8437 (N_8437,N_7167,N_7325);
nor U8438 (N_8438,N_7724,N_7675);
and U8439 (N_8439,N_7697,N_7586);
nor U8440 (N_8440,N_7362,N_7024);
and U8441 (N_8441,N_7387,N_7227);
nor U8442 (N_8442,N_7518,N_7261);
and U8443 (N_8443,N_7126,N_7590);
or U8444 (N_8444,N_7771,N_7359);
or U8445 (N_8445,N_7195,N_7605);
or U8446 (N_8446,N_7858,N_7374);
nand U8447 (N_8447,N_7183,N_7886);
nand U8448 (N_8448,N_7726,N_7297);
or U8449 (N_8449,N_7334,N_7088);
nand U8450 (N_8450,N_7874,N_7121);
nor U8451 (N_8451,N_7846,N_7754);
nand U8452 (N_8452,N_7064,N_7972);
nor U8453 (N_8453,N_7484,N_7004);
and U8454 (N_8454,N_7798,N_7785);
nor U8455 (N_8455,N_7729,N_7576);
and U8456 (N_8456,N_7688,N_7411);
or U8457 (N_8457,N_7044,N_7839);
nand U8458 (N_8458,N_7877,N_7185);
and U8459 (N_8459,N_7977,N_7361);
and U8460 (N_8460,N_7848,N_7386);
and U8461 (N_8461,N_7146,N_7040);
nor U8462 (N_8462,N_7732,N_7492);
nand U8463 (N_8463,N_7861,N_7664);
nor U8464 (N_8464,N_7597,N_7155);
nand U8465 (N_8465,N_7365,N_7220);
nor U8466 (N_8466,N_7087,N_7950);
nand U8467 (N_8467,N_7376,N_7580);
or U8468 (N_8468,N_7791,N_7872);
or U8469 (N_8469,N_7691,N_7658);
or U8470 (N_8470,N_7370,N_7001);
nand U8471 (N_8471,N_7967,N_7078);
nor U8472 (N_8472,N_7547,N_7091);
nor U8473 (N_8473,N_7555,N_7514);
or U8474 (N_8474,N_7945,N_7037);
or U8475 (N_8475,N_7583,N_7383);
or U8476 (N_8476,N_7687,N_7673);
nand U8477 (N_8477,N_7990,N_7299);
nand U8478 (N_8478,N_7931,N_7561);
nand U8479 (N_8479,N_7187,N_7709);
or U8480 (N_8480,N_7526,N_7993);
and U8481 (N_8481,N_7034,N_7013);
or U8482 (N_8482,N_7477,N_7985);
nor U8483 (N_8483,N_7866,N_7932);
and U8484 (N_8484,N_7216,N_7090);
nand U8485 (N_8485,N_7337,N_7303);
and U8486 (N_8486,N_7867,N_7720);
nor U8487 (N_8487,N_7348,N_7750);
nand U8488 (N_8488,N_7584,N_7247);
nor U8489 (N_8489,N_7905,N_7818);
and U8490 (N_8490,N_7450,N_7027);
and U8491 (N_8491,N_7591,N_7252);
nor U8492 (N_8492,N_7284,N_7540);
or U8493 (N_8493,N_7814,N_7240);
nand U8494 (N_8494,N_7857,N_7494);
nand U8495 (N_8495,N_7722,N_7834);
nor U8496 (N_8496,N_7211,N_7496);
or U8497 (N_8497,N_7423,N_7206);
nand U8498 (N_8498,N_7891,N_7718);
nor U8499 (N_8499,N_7236,N_7214);
nor U8500 (N_8500,N_7776,N_7501);
nand U8501 (N_8501,N_7635,N_7683);
or U8502 (N_8502,N_7060,N_7873);
nor U8503 (N_8503,N_7714,N_7911);
nand U8504 (N_8504,N_7660,N_7902);
or U8505 (N_8505,N_7262,N_7729);
nand U8506 (N_8506,N_7475,N_7250);
nand U8507 (N_8507,N_7453,N_7563);
and U8508 (N_8508,N_7176,N_7886);
nand U8509 (N_8509,N_7201,N_7541);
nand U8510 (N_8510,N_7146,N_7920);
or U8511 (N_8511,N_7505,N_7490);
and U8512 (N_8512,N_7039,N_7832);
nor U8513 (N_8513,N_7446,N_7932);
nand U8514 (N_8514,N_7035,N_7227);
and U8515 (N_8515,N_7874,N_7631);
nand U8516 (N_8516,N_7054,N_7374);
nor U8517 (N_8517,N_7896,N_7693);
and U8518 (N_8518,N_7606,N_7449);
and U8519 (N_8519,N_7378,N_7829);
nand U8520 (N_8520,N_7579,N_7354);
nand U8521 (N_8521,N_7074,N_7283);
nor U8522 (N_8522,N_7252,N_7135);
nand U8523 (N_8523,N_7365,N_7377);
nand U8524 (N_8524,N_7135,N_7416);
xnor U8525 (N_8525,N_7040,N_7578);
nand U8526 (N_8526,N_7665,N_7149);
or U8527 (N_8527,N_7298,N_7102);
nor U8528 (N_8528,N_7069,N_7122);
and U8529 (N_8529,N_7597,N_7377);
nand U8530 (N_8530,N_7303,N_7018);
nor U8531 (N_8531,N_7599,N_7469);
and U8532 (N_8532,N_7425,N_7320);
nand U8533 (N_8533,N_7757,N_7586);
and U8534 (N_8534,N_7079,N_7274);
or U8535 (N_8535,N_7325,N_7813);
or U8536 (N_8536,N_7195,N_7870);
and U8537 (N_8537,N_7964,N_7352);
nand U8538 (N_8538,N_7116,N_7589);
and U8539 (N_8539,N_7263,N_7647);
and U8540 (N_8540,N_7833,N_7637);
or U8541 (N_8541,N_7911,N_7970);
nand U8542 (N_8542,N_7273,N_7296);
nor U8543 (N_8543,N_7926,N_7241);
or U8544 (N_8544,N_7999,N_7270);
nor U8545 (N_8545,N_7926,N_7865);
and U8546 (N_8546,N_7522,N_7423);
or U8547 (N_8547,N_7396,N_7436);
nor U8548 (N_8548,N_7843,N_7634);
or U8549 (N_8549,N_7355,N_7816);
and U8550 (N_8550,N_7208,N_7275);
nor U8551 (N_8551,N_7668,N_7693);
or U8552 (N_8552,N_7354,N_7348);
nand U8553 (N_8553,N_7057,N_7985);
nand U8554 (N_8554,N_7037,N_7723);
or U8555 (N_8555,N_7294,N_7662);
nand U8556 (N_8556,N_7670,N_7789);
xnor U8557 (N_8557,N_7796,N_7683);
and U8558 (N_8558,N_7115,N_7898);
nor U8559 (N_8559,N_7595,N_7751);
nand U8560 (N_8560,N_7297,N_7764);
nand U8561 (N_8561,N_7202,N_7326);
nor U8562 (N_8562,N_7076,N_7327);
nor U8563 (N_8563,N_7854,N_7743);
nor U8564 (N_8564,N_7966,N_7893);
nor U8565 (N_8565,N_7307,N_7953);
and U8566 (N_8566,N_7951,N_7014);
and U8567 (N_8567,N_7836,N_7680);
nand U8568 (N_8568,N_7526,N_7919);
nand U8569 (N_8569,N_7934,N_7044);
or U8570 (N_8570,N_7406,N_7643);
nand U8571 (N_8571,N_7149,N_7368);
or U8572 (N_8572,N_7123,N_7126);
nor U8573 (N_8573,N_7419,N_7530);
nor U8574 (N_8574,N_7254,N_7206);
or U8575 (N_8575,N_7086,N_7007);
nor U8576 (N_8576,N_7411,N_7737);
nand U8577 (N_8577,N_7459,N_7418);
or U8578 (N_8578,N_7176,N_7090);
and U8579 (N_8579,N_7694,N_7301);
and U8580 (N_8580,N_7843,N_7232);
and U8581 (N_8581,N_7354,N_7100);
or U8582 (N_8582,N_7846,N_7319);
nand U8583 (N_8583,N_7704,N_7191);
nand U8584 (N_8584,N_7462,N_7801);
nor U8585 (N_8585,N_7435,N_7711);
nor U8586 (N_8586,N_7890,N_7786);
nor U8587 (N_8587,N_7524,N_7981);
and U8588 (N_8588,N_7421,N_7048);
and U8589 (N_8589,N_7787,N_7771);
nor U8590 (N_8590,N_7619,N_7884);
nand U8591 (N_8591,N_7622,N_7559);
and U8592 (N_8592,N_7613,N_7460);
nor U8593 (N_8593,N_7804,N_7115);
or U8594 (N_8594,N_7269,N_7442);
nand U8595 (N_8595,N_7445,N_7544);
nand U8596 (N_8596,N_7191,N_7892);
or U8597 (N_8597,N_7121,N_7137);
or U8598 (N_8598,N_7084,N_7870);
nand U8599 (N_8599,N_7052,N_7776);
nand U8600 (N_8600,N_7309,N_7071);
or U8601 (N_8601,N_7088,N_7722);
and U8602 (N_8602,N_7690,N_7893);
and U8603 (N_8603,N_7282,N_7243);
and U8604 (N_8604,N_7027,N_7288);
nand U8605 (N_8605,N_7742,N_7200);
and U8606 (N_8606,N_7572,N_7502);
nand U8607 (N_8607,N_7827,N_7266);
nand U8608 (N_8608,N_7256,N_7682);
nand U8609 (N_8609,N_7978,N_7979);
nor U8610 (N_8610,N_7586,N_7420);
nand U8611 (N_8611,N_7972,N_7739);
nor U8612 (N_8612,N_7269,N_7760);
or U8613 (N_8613,N_7272,N_7838);
nand U8614 (N_8614,N_7421,N_7195);
nand U8615 (N_8615,N_7048,N_7785);
and U8616 (N_8616,N_7112,N_7362);
and U8617 (N_8617,N_7417,N_7866);
nor U8618 (N_8618,N_7687,N_7128);
and U8619 (N_8619,N_7666,N_7464);
and U8620 (N_8620,N_7754,N_7920);
or U8621 (N_8621,N_7549,N_7561);
and U8622 (N_8622,N_7641,N_7686);
or U8623 (N_8623,N_7675,N_7054);
nor U8624 (N_8624,N_7032,N_7875);
or U8625 (N_8625,N_7632,N_7038);
and U8626 (N_8626,N_7265,N_7731);
or U8627 (N_8627,N_7481,N_7120);
nand U8628 (N_8628,N_7706,N_7679);
and U8629 (N_8629,N_7414,N_7128);
or U8630 (N_8630,N_7076,N_7586);
or U8631 (N_8631,N_7096,N_7190);
nand U8632 (N_8632,N_7843,N_7294);
nand U8633 (N_8633,N_7015,N_7318);
nand U8634 (N_8634,N_7426,N_7113);
nand U8635 (N_8635,N_7576,N_7166);
or U8636 (N_8636,N_7190,N_7274);
nand U8637 (N_8637,N_7411,N_7003);
nand U8638 (N_8638,N_7706,N_7350);
and U8639 (N_8639,N_7604,N_7420);
nor U8640 (N_8640,N_7477,N_7839);
nand U8641 (N_8641,N_7967,N_7863);
or U8642 (N_8642,N_7481,N_7704);
or U8643 (N_8643,N_7094,N_7552);
and U8644 (N_8644,N_7734,N_7496);
nor U8645 (N_8645,N_7407,N_7391);
or U8646 (N_8646,N_7035,N_7098);
nand U8647 (N_8647,N_7195,N_7380);
nand U8648 (N_8648,N_7423,N_7146);
nor U8649 (N_8649,N_7411,N_7435);
and U8650 (N_8650,N_7096,N_7407);
and U8651 (N_8651,N_7212,N_7444);
and U8652 (N_8652,N_7543,N_7312);
and U8653 (N_8653,N_7682,N_7167);
and U8654 (N_8654,N_7222,N_7357);
nand U8655 (N_8655,N_7925,N_7333);
nor U8656 (N_8656,N_7043,N_7062);
or U8657 (N_8657,N_7494,N_7870);
nand U8658 (N_8658,N_7290,N_7560);
nand U8659 (N_8659,N_7700,N_7037);
or U8660 (N_8660,N_7475,N_7207);
nand U8661 (N_8661,N_7496,N_7052);
nand U8662 (N_8662,N_7630,N_7615);
nand U8663 (N_8663,N_7975,N_7891);
nor U8664 (N_8664,N_7086,N_7394);
and U8665 (N_8665,N_7864,N_7535);
and U8666 (N_8666,N_7287,N_7240);
nand U8667 (N_8667,N_7758,N_7967);
nor U8668 (N_8668,N_7742,N_7774);
nand U8669 (N_8669,N_7639,N_7202);
nor U8670 (N_8670,N_7269,N_7863);
nor U8671 (N_8671,N_7436,N_7318);
and U8672 (N_8672,N_7055,N_7338);
and U8673 (N_8673,N_7961,N_7488);
nor U8674 (N_8674,N_7884,N_7472);
nor U8675 (N_8675,N_7514,N_7928);
nand U8676 (N_8676,N_7795,N_7964);
nor U8677 (N_8677,N_7208,N_7044);
nand U8678 (N_8678,N_7764,N_7401);
nor U8679 (N_8679,N_7826,N_7530);
nor U8680 (N_8680,N_7621,N_7195);
nand U8681 (N_8681,N_7578,N_7690);
and U8682 (N_8682,N_7748,N_7274);
nor U8683 (N_8683,N_7802,N_7521);
or U8684 (N_8684,N_7068,N_7541);
and U8685 (N_8685,N_7888,N_7638);
or U8686 (N_8686,N_7006,N_7172);
and U8687 (N_8687,N_7707,N_7793);
nand U8688 (N_8688,N_7704,N_7917);
nor U8689 (N_8689,N_7343,N_7103);
or U8690 (N_8690,N_7714,N_7944);
nor U8691 (N_8691,N_7700,N_7109);
or U8692 (N_8692,N_7461,N_7618);
nand U8693 (N_8693,N_7230,N_7200);
nor U8694 (N_8694,N_7696,N_7969);
nand U8695 (N_8695,N_7959,N_7115);
and U8696 (N_8696,N_7755,N_7017);
or U8697 (N_8697,N_7003,N_7151);
nand U8698 (N_8698,N_7366,N_7592);
nor U8699 (N_8699,N_7542,N_7318);
or U8700 (N_8700,N_7683,N_7003);
or U8701 (N_8701,N_7885,N_7963);
or U8702 (N_8702,N_7010,N_7866);
nor U8703 (N_8703,N_7375,N_7870);
nand U8704 (N_8704,N_7861,N_7976);
nand U8705 (N_8705,N_7738,N_7575);
or U8706 (N_8706,N_7347,N_7616);
nand U8707 (N_8707,N_7488,N_7946);
nand U8708 (N_8708,N_7236,N_7213);
or U8709 (N_8709,N_7471,N_7020);
nand U8710 (N_8710,N_7072,N_7914);
nand U8711 (N_8711,N_7427,N_7135);
nor U8712 (N_8712,N_7901,N_7198);
or U8713 (N_8713,N_7955,N_7791);
and U8714 (N_8714,N_7402,N_7845);
nand U8715 (N_8715,N_7183,N_7213);
nand U8716 (N_8716,N_7812,N_7143);
nand U8717 (N_8717,N_7491,N_7187);
or U8718 (N_8718,N_7300,N_7790);
and U8719 (N_8719,N_7014,N_7824);
or U8720 (N_8720,N_7527,N_7560);
nand U8721 (N_8721,N_7750,N_7679);
nand U8722 (N_8722,N_7234,N_7466);
nand U8723 (N_8723,N_7540,N_7651);
nor U8724 (N_8724,N_7654,N_7863);
nand U8725 (N_8725,N_7060,N_7001);
and U8726 (N_8726,N_7094,N_7378);
and U8727 (N_8727,N_7527,N_7952);
nand U8728 (N_8728,N_7720,N_7208);
and U8729 (N_8729,N_7174,N_7350);
and U8730 (N_8730,N_7965,N_7564);
and U8731 (N_8731,N_7067,N_7048);
nand U8732 (N_8732,N_7797,N_7873);
nor U8733 (N_8733,N_7005,N_7079);
or U8734 (N_8734,N_7356,N_7089);
or U8735 (N_8735,N_7427,N_7512);
and U8736 (N_8736,N_7699,N_7933);
nand U8737 (N_8737,N_7388,N_7167);
or U8738 (N_8738,N_7028,N_7033);
and U8739 (N_8739,N_7019,N_7439);
and U8740 (N_8740,N_7203,N_7983);
or U8741 (N_8741,N_7901,N_7541);
or U8742 (N_8742,N_7620,N_7662);
nand U8743 (N_8743,N_7096,N_7101);
and U8744 (N_8744,N_7414,N_7702);
or U8745 (N_8745,N_7528,N_7781);
or U8746 (N_8746,N_7392,N_7531);
nor U8747 (N_8747,N_7741,N_7226);
and U8748 (N_8748,N_7356,N_7211);
nor U8749 (N_8749,N_7151,N_7034);
or U8750 (N_8750,N_7461,N_7281);
and U8751 (N_8751,N_7959,N_7867);
and U8752 (N_8752,N_7285,N_7245);
nor U8753 (N_8753,N_7759,N_7649);
nor U8754 (N_8754,N_7480,N_7930);
or U8755 (N_8755,N_7123,N_7188);
and U8756 (N_8756,N_7282,N_7679);
or U8757 (N_8757,N_7340,N_7898);
and U8758 (N_8758,N_7073,N_7438);
or U8759 (N_8759,N_7255,N_7838);
or U8760 (N_8760,N_7683,N_7803);
and U8761 (N_8761,N_7957,N_7777);
or U8762 (N_8762,N_7998,N_7903);
nand U8763 (N_8763,N_7745,N_7364);
or U8764 (N_8764,N_7136,N_7111);
and U8765 (N_8765,N_7227,N_7922);
nand U8766 (N_8766,N_7845,N_7733);
and U8767 (N_8767,N_7015,N_7139);
and U8768 (N_8768,N_7061,N_7518);
nor U8769 (N_8769,N_7260,N_7887);
or U8770 (N_8770,N_7687,N_7968);
and U8771 (N_8771,N_7747,N_7690);
nand U8772 (N_8772,N_7698,N_7446);
or U8773 (N_8773,N_7081,N_7641);
and U8774 (N_8774,N_7806,N_7314);
nor U8775 (N_8775,N_7917,N_7898);
and U8776 (N_8776,N_7552,N_7000);
and U8777 (N_8777,N_7508,N_7368);
nor U8778 (N_8778,N_7273,N_7220);
or U8779 (N_8779,N_7494,N_7288);
and U8780 (N_8780,N_7642,N_7777);
and U8781 (N_8781,N_7972,N_7230);
and U8782 (N_8782,N_7658,N_7532);
nand U8783 (N_8783,N_7356,N_7014);
nand U8784 (N_8784,N_7134,N_7914);
nand U8785 (N_8785,N_7193,N_7970);
or U8786 (N_8786,N_7203,N_7138);
nor U8787 (N_8787,N_7061,N_7568);
nor U8788 (N_8788,N_7254,N_7721);
and U8789 (N_8789,N_7731,N_7019);
or U8790 (N_8790,N_7073,N_7921);
or U8791 (N_8791,N_7696,N_7528);
and U8792 (N_8792,N_7558,N_7131);
or U8793 (N_8793,N_7704,N_7122);
nand U8794 (N_8794,N_7414,N_7913);
nand U8795 (N_8795,N_7929,N_7806);
or U8796 (N_8796,N_7063,N_7380);
or U8797 (N_8797,N_7451,N_7295);
nand U8798 (N_8798,N_7809,N_7953);
and U8799 (N_8799,N_7727,N_7983);
or U8800 (N_8800,N_7084,N_7959);
or U8801 (N_8801,N_7827,N_7293);
or U8802 (N_8802,N_7817,N_7241);
and U8803 (N_8803,N_7742,N_7338);
and U8804 (N_8804,N_7894,N_7437);
or U8805 (N_8805,N_7122,N_7261);
or U8806 (N_8806,N_7902,N_7110);
nor U8807 (N_8807,N_7306,N_7070);
and U8808 (N_8808,N_7966,N_7904);
and U8809 (N_8809,N_7473,N_7991);
nand U8810 (N_8810,N_7438,N_7786);
or U8811 (N_8811,N_7293,N_7150);
and U8812 (N_8812,N_7275,N_7023);
nand U8813 (N_8813,N_7805,N_7169);
nand U8814 (N_8814,N_7509,N_7088);
nor U8815 (N_8815,N_7968,N_7084);
nand U8816 (N_8816,N_7475,N_7002);
nor U8817 (N_8817,N_7153,N_7393);
nand U8818 (N_8818,N_7346,N_7140);
nand U8819 (N_8819,N_7131,N_7362);
nor U8820 (N_8820,N_7334,N_7007);
nand U8821 (N_8821,N_7515,N_7870);
nand U8822 (N_8822,N_7850,N_7136);
and U8823 (N_8823,N_7947,N_7793);
nor U8824 (N_8824,N_7647,N_7990);
or U8825 (N_8825,N_7873,N_7309);
xnor U8826 (N_8826,N_7781,N_7324);
or U8827 (N_8827,N_7478,N_7514);
or U8828 (N_8828,N_7409,N_7046);
or U8829 (N_8829,N_7663,N_7956);
nor U8830 (N_8830,N_7978,N_7783);
nand U8831 (N_8831,N_7230,N_7117);
xnor U8832 (N_8832,N_7362,N_7906);
or U8833 (N_8833,N_7913,N_7953);
or U8834 (N_8834,N_7928,N_7084);
and U8835 (N_8835,N_7364,N_7948);
and U8836 (N_8836,N_7743,N_7424);
or U8837 (N_8837,N_7497,N_7769);
or U8838 (N_8838,N_7390,N_7021);
and U8839 (N_8839,N_7164,N_7125);
nor U8840 (N_8840,N_7019,N_7093);
and U8841 (N_8841,N_7652,N_7664);
or U8842 (N_8842,N_7971,N_7616);
nand U8843 (N_8843,N_7184,N_7566);
nand U8844 (N_8844,N_7565,N_7208);
nor U8845 (N_8845,N_7541,N_7082);
nor U8846 (N_8846,N_7528,N_7304);
and U8847 (N_8847,N_7369,N_7298);
and U8848 (N_8848,N_7689,N_7954);
or U8849 (N_8849,N_7385,N_7368);
nor U8850 (N_8850,N_7948,N_7807);
nand U8851 (N_8851,N_7941,N_7634);
and U8852 (N_8852,N_7905,N_7440);
nand U8853 (N_8853,N_7251,N_7982);
and U8854 (N_8854,N_7750,N_7534);
or U8855 (N_8855,N_7330,N_7974);
nand U8856 (N_8856,N_7228,N_7929);
nor U8857 (N_8857,N_7030,N_7406);
or U8858 (N_8858,N_7483,N_7216);
nor U8859 (N_8859,N_7130,N_7434);
or U8860 (N_8860,N_7460,N_7046);
nor U8861 (N_8861,N_7312,N_7846);
xnor U8862 (N_8862,N_7800,N_7070);
and U8863 (N_8863,N_7217,N_7670);
nand U8864 (N_8864,N_7026,N_7738);
or U8865 (N_8865,N_7982,N_7476);
nand U8866 (N_8866,N_7815,N_7200);
nand U8867 (N_8867,N_7583,N_7762);
and U8868 (N_8868,N_7534,N_7782);
or U8869 (N_8869,N_7902,N_7571);
and U8870 (N_8870,N_7518,N_7760);
nand U8871 (N_8871,N_7619,N_7935);
nand U8872 (N_8872,N_7958,N_7675);
nand U8873 (N_8873,N_7505,N_7519);
nand U8874 (N_8874,N_7260,N_7484);
nand U8875 (N_8875,N_7366,N_7164);
nand U8876 (N_8876,N_7519,N_7899);
nor U8877 (N_8877,N_7999,N_7098);
or U8878 (N_8878,N_7413,N_7316);
or U8879 (N_8879,N_7696,N_7027);
nand U8880 (N_8880,N_7331,N_7488);
and U8881 (N_8881,N_7453,N_7068);
and U8882 (N_8882,N_7094,N_7333);
nand U8883 (N_8883,N_7457,N_7661);
or U8884 (N_8884,N_7084,N_7657);
or U8885 (N_8885,N_7796,N_7311);
or U8886 (N_8886,N_7638,N_7301);
or U8887 (N_8887,N_7460,N_7903);
and U8888 (N_8888,N_7010,N_7960);
xnor U8889 (N_8889,N_7135,N_7883);
or U8890 (N_8890,N_7668,N_7450);
nand U8891 (N_8891,N_7776,N_7071);
nand U8892 (N_8892,N_7005,N_7896);
or U8893 (N_8893,N_7035,N_7016);
or U8894 (N_8894,N_7679,N_7953);
nor U8895 (N_8895,N_7432,N_7624);
and U8896 (N_8896,N_7911,N_7921);
and U8897 (N_8897,N_7568,N_7845);
or U8898 (N_8898,N_7822,N_7541);
or U8899 (N_8899,N_7797,N_7452);
or U8900 (N_8900,N_7254,N_7798);
and U8901 (N_8901,N_7370,N_7353);
and U8902 (N_8902,N_7163,N_7277);
or U8903 (N_8903,N_7958,N_7213);
nand U8904 (N_8904,N_7752,N_7344);
or U8905 (N_8905,N_7541,N_7542);
and U8906 (N_8906,N_7244,N_7713);
nand U8907 (N_8907,N_7786,N_7833);
or U8908 (N_8908,N_7299,N_7367);
nand U8909 (N_8909,N_7809,N_7950);
or U8910 (N_8910,N_7824,N_7551);
nor U8911 (N_8911,N_7659,N_7468);
nand U8912 (N_8912,N_7506,N_7193);
nor U8913 (N_8913,N_7729,N_7065);
or U8914 (N_8914,N_7553,N_7032);
nor U8915 (N_8915,N_7595,N_7815);
and U8916 (N_8916,N_7759,N_7417);
and U8917 (N_8917,N_7446,N_7253);
or U8918 (N_8918,N_7506,N_7966);
nand U8919 (N_8919,N_7712,N_7720);
and U8920 (N_8920,N_7178,N_7634);
nand U8921 (N_8921,N_7030,N_7118);
nand U8922 (N_8922,N_7928,N_7183);
and U8923 (N_8923,N_7563,N_7008);
nor U8924 (N_8924,N_7581,N_7607);
nand U8925 (N_8925,N_7833,N_7701);
or U8926 (N_8926,N_7651,N_7647);
nor U8927 (N_8927,N_7459,N_7410);
or U8928 (N_8928,N_7648,N_7908);
and U8929 (N_8929,N_7309,N_7695);
and U8930 (N_8930,N_7921,N_7859);
or U8931 (N_8931,N_7623,N_7213);
nor U8932 (N_8932,N_7106,N_7234);
and U8933 (N_8933,N_7628,N_7444);
and U8934 (N_8934,N_7774,N_7570);
or U8935 (N_8935,N_7983,N_7441);
and U8936 (N_8936,N_7007,N_7987);
and U8937 (N_8937,N_7772,N_7881);
or U8938 (N_8938,N_7897,N_7482);
and U8939 (N_8939,N_7738,N_7038);
or U8940 (N_8940,N_7794,N_7767);
nor U8941 (N_8941,N_7818,N_7822);
or U8942 (N_8942,N_7557,N_7162);
nand U8943 (N_8943,N_7320,N_7148);
nor U8944 (N_8944,N_7997,N_7013);
nor U8945 (N_8945,N_7125,N_7466);
or U8946 (N_8946,N_7429,N_7972);
nor U8947 (N_8947,N_7263,N_7340);
nand U8948 (N_8948,N_7657,N_7373);
and U8949 (N_8949,N_7762,N_7120);
nand U8950 (N_8950,N_7682,N_7986);
nor U8951 (N_8951,N_7633,N_7536);
and U8952 (N_8952,N_7483,N_7555);
nand U8953 (N_8953,N_7190,N_7501);
or U8954 (N_8954,N_7287,N_7311);
nor U8955 (N_8955,N_7914,N_7055);
nand U8956 (N_8956,N_7472,N_7895);
nand U8957 (N_8957,N_7945,N_7922);
nor U8958 (N_8958,N_7532,N_7197);
and U8959 (N_8959,N_7582,N_7058);
and U8960 (N_8960,N_7429,N_7703);
or U8961 (N_8961,N_7827,N_7759);
nor U8962 (N_8962,N_7539,N_7561);
nand U8963 (N_8963,N_7601,N_7548);
nor U8964 (N_8964,N_7161,N_7408);
or U8965 (N_8965,N_7305,N_7182);
and U8966 (N_8966,N_7811,N_7756);
nand U8967 (N_8967,N_7398,N_7721);
xor U8968 (N_8968,N_7802,N_7577);
nand U8969 (N_8969,N_7699,N_7305);
or U8970 (N_8970,N_7770,N_7478);
nand U8971 (N_8971,N_7140,N_7772);
or U8972 (N_8972,N_7578,N_7699);
and U8973 (N_8973,N_7349,N_7455);
or U8974 (N_8974,N_7330,N_7003);
nand U8975 (N_8975,N_7217,N_7891);
nor U8976 (N_8976,N_7432,N_7054);
or U8977 (N_8977,N_7187,N_7710);
nand U8978 (N_8978,N_7891,N_7978);
or U8979 (N_8979,N_7239,N_7813);
nor U8980 (N_8980,N_7188,N_7262);
nor U8981 (N_8981,N_7034,N_7414);
and U8982 (N_8982,N_7785,N_7828);
nor U8983 (N_8983,N_7488,N_7969);
nor U8984 (N_8984,N_7722,N_7987);
nand U8985 (N_8985,N_7277,N_7564);
and U8986 (N_8986,N_7571,N_7081);
nand U8987 (N_8987,N_7477,N_7090);
nand U8988 (N_8988,N_7101,N_7462);
nand U8989 (N_8989,N_7256,N_7224);
or U8990 (N_8990,N_7406,N_7424);
nand U8991 (N_8991,N_7223,N_7975);
nor U8992 (N_8992,N_7621,N_7538);
nand U8993 (N_8993,N_7679,N_7393);
and U8994 (N_8994,N_7467,N_7892);
nand U8995 (N_8995,N_7365,N_7284);
and U8996 (N_8996,N_7678,N_7874);
nand U8997 (N_8997,N_7186,N_7748);
nor U8998 (N_8998,N_7827,N_7532);
or U8999 (N_8999,N_7313,N_7730);
nand U9000 (N_9000,N_8760,N_8851);
or U9001 (N_9001,N_8818,N_8267);
and U9002 (N_9002,N_8703,N_8946);
nor U9003 (N_9003,N_8385,N_8016);
and U9004 (N_9004,N_8673,N_8455);
nand U9005 (N_9005,N_8330,N_8697);
nor U9006 (N_9006,N_8966,N_8753);
nor U9007 (N_9007,N_8684,N_8291);
or U9008 (N_9008,N_8632,N_8453);
nand U9009 (N_9009,N_8489,N_8250);
or U9010 (N_9010,N_8492,N_8417);
or U9011 (N_9011,N_8032,N_8985);
and U9012 (N_9012,N_8925,N_8205);
or U9013 (N_9013,N_8853,N_8070);
nor U9014 (N_9014,N_8692,N_8962);
and U9015 (N_9015,N_8174,N_8980);
nor U9016 (N_9016,N_8161,N_8126);
and U9017 (N_9017,N_8058,N_8483);
and U9018 (N_9018,N_8369,N_8309);
nand U9019 (N_9019,N_8781,N_8638);
nor U9020 (N_9020,N_8912,N_8235);
nand U9021 (N_9021,N_8829,N_8444);
or U9022 (N_9022,N_8939,N_8326);
nor U9023 (N_9023,N_8854,N_8850);
and U9024 (N_9024,N_8571,N_8775);
nor U9025 (N_9025,N_8322,N_8486);
or U9026 (N_9026,N_8176,N_8334);
and U9027 (N_9027,N_8628,N_8215);
nand U9028 (N_9028,N_8091,N_8252);
nand U9029 (N_9029,N_8332,N_8393);
and U9030 (N_9030,N_8436,N_8941);
nand U9031 (N_9031,N_8248,N_8389);
or U9032 (N_9032,N_8631,N_8314);
or U9033 (N_9033,N_8724,N_8635);
and U9034 (N_9034,N_8062,N_8924);
nand U9035 (N_9035,N_8297,N_8415);
nand U9036 (N_9036,N_8147,N_8481);
and U9037 (N_9037,N_8814,N_8173);
nor U9038 (N_9038,N_8101,N_8034);
nor U9039 (N_9039,N_8838,N_8596);
nand U9040 (N_9040,N_8266,N_8410);
and U9041 (N_9041,N_8038,N_8433);
or U9042 (N_9042,N_8458,N_8637);
and U9043 (N_9043,N_8157,N_8808);
nand U9044 (N_9044,N_8262,N_8527);
nor U9045 (N_9045,N_8194,N_8499);
and U9046 (N_9046,N_8895,N_8054);
nand U9047 (N_9047,N_8493,N_8669);
and U9048 (N_9048,N_8747,N_8471);
nand U9049 (N_9049,N_8689,N_8022);
or U9050 (N_9050,N_8856,N_8013);
or U9051 (N_9051,N_8019,N_8357);
nand U9052 (N_9052,N_8382,N_8464);
nand U9053 (N_9053,N_8447,N_8963);
nor U9054 (N_9054,N_8365,N_8052);
or U9055 (N_9055,N_8594,N_8435);
or U9056 (N_9056,N_8193,N_8535);
nor U9057 (N_9057,N_8813,N_8111);
or U9058 (N_9058,N_8236,N_8220);
nor U9059 (N_9059,N_8354,N_8894);
and U9060 (N_9060,N_8618,N_8118);
nand U9061 (N_9061,N_8706,N_8796);
nor U9062 (N_9062,N_8621,N_8336);
nand U9063 (N_9063,N_8822,N_8816);
nor U9064 (N_9064,N_8782,N_8619);
and U9065 (N_9065,N_8408,N_8356);
nand U9066 (N_9066,N_8974,N_8636);
or U9067 (N_9067,N_8209,N_8454);
and U9068 (N_9068,N_8456,N_8682);
nand U9069 (N_9069,N_8112,N_8418);
nand U9070 (N_9070,N_8053,N_8146);
nand U9071 (N_9071,N_8092,N_8694);
nor U9072 (N_9072,N_8578,N_8559);
nor U9073 (N_9073,N_8475,N_8949);
and U9074 (N_9074,N_8374,N_8687);
nand U9075 (N_9075,N_8473,N_8109);
or U9076 (N_9076,N_8608,N_8798);
nand U9077 (N_9077,N_8242,N_8707);
and U9078 (N_9078,N_8617,N_8983);
and U9079 (N_9079,N_8756,N_8353);
nand U9080 (N_9080,N_8595,N_8024);
and U9081 (N_9081,N_8730,N_8523);
nor U9082 (N_9082,N_8922,N_8461);
or U9083 (N_9083,N_8411,N_8386);
nor U9084 (N_9084,N_8565,N_8218);
nor U9085 (N_9085,N_8546,N_8195);
and U9086 (N_9086,N_8751,N_8178);
and U9087 (N_9087,N_8343,N_8529);
xnor U9088 (N_9088,N_8133,N_8391);
nor U9089 (N_9089,N_8642,N_8355);
nor U9090 (N_9090,N_8167,N_8819);
nor U9091 (N_9091,N_8001,N_8691);
or U9092 (N_9092,N_8197,N_8733);
nand U9093 (N_9093,N_8875,N_8153);
nand U9094 (N_9094,N_8539,N_8044);
nand U9095 (N_9095,N_8807,N_8294);
nand U9096 (N_9096,N_8046,N_8863);
nand U9097 (N_9097,N_8422,N_8287);
or U9098 (N_9098,N_8237,N_8679);
xor U9099 (N_9099,N_8379,N_8975);
nor U9100 (N_9100,N_8114,N_8906);
or U9101 (N_9101,N_8340,N_8260);
nor U9102 (N_9102,N_8584,N_8081);
and U9103 (N_9103,N_8779,N_8186);
or U9104 (N_9104,N_8509,N_8900);
or U9105 (N_9105,N_8738,N_8725);
and U9106 (N_9106,N_8893,N_8289);
nand U9107 (N_9107,N_8520,N_8352);
nor U9108 (N_9108,N_8071,N_8590);
nand U9109 (N_9109,N_8095,N_8791);
and U9110 (N_9110,N_8213,N_8858);
nor U9111 (N_9111,N_8898,N_8362);
or U9112 (N_9112,N_8478,N_8373);
nor U9113 (N_9113,N_8469,N_8166);
nor U9114 (N_9114,N_8093,N_8364);
nand U9115 (N_9115,N_8904,N_8006);
xnor U9116 (N_9116,N_8639,N_8686);
and U9117 (N_9117,N_8712,N_8304);
nor U9118 (N_9118,N_8238,N_8168);
nor U9119 (N_9119,N_8564,N_8954);
nor U9120 (N_9120,N_8171,N_8026);
or U9121 (N_9121,N_8901,N_8459);
and U9122 (N_9122,N_8698,N_8870);
nor U9123 (N_9123,N_8605,N_8263);
or U9124 (N_9124,N_8667,N_8398);
or U9125 (N_9125,N_8347,N_8744);
and U9126 (N_9126,N_8778,N_8871);
nand U9127 (N_9127,N_8059,N_8315);
and U9128 (N_9128,N_8131,N_8116);
and U9129 (N_9129,N_8843,N_8548);
nand U9130 (N_9130,N_8042,N_8606);
nor U9131 (N_9131,N_8028,N_8562);
nand U9132 (N_9132,N_8494,N_8510);
nor U9133 (N_9133,N_8857,N_8011);
nor U9134 (N_9134,N_8407,N_8221);
or U9135 (N_9135,N_8283,N_8089);
nand U9136 (N_9136,N_8570,N_8083);
or U9137 (N_9137,N_8976,N_8107);
xnor U9138 (N_9138,N_8414,N_8795);
nand U9139 (N_9139,N_8793,N_8251);
or U9140 (N_9140,N_8395,N_8349);
nor U9141 (N_9141,N_8233,N_8652);
nand U9142 (N_9142,N_8105,N_8031);
or U9143 (N_9143,N_8285,N_8224);
and U9144 (N_9144,N_8427,N_8501);
or U9145 (N_9145,N_8067,N_8214);
nand U9146 (N_9146,N_8310,N_8345);
and U9147 (N_9147,N_8537,N_8358);
or U9148 (N_9148,N_8479,N_8230);
and U9149 (N_9149,N_8384,N_8592);
nor U9150 (N_9150,N_8948,N_8074);
and U9151 (N_9151,N_8869,N_8246);
and U9152 (N_9152,N_8512,N_8463);
and U9153 (N_9153,N_8879,N_8005);
or U9154 (N_9154,N_8069,N_8002);
nor U9155 (N_9155,N_8327,N_8833);
or U9156 (N_9156,N_8401,N_8615);
and U9157 (N_9157,N_8583,N_8518);
nor U9158 (N_9158,N_8862,N_8634);
nand U9159 (N_9159,N_8579,N_8553);
and U9160 (N_9160,N_8700,N_8317);
and U9161 (N_9161,N_8280,N_8312);
nand U9162 (N_9162,N_8409,N_8487);
nand U9163 (N_9163,N_8203,N_8713);
nand U9164 (N_9164,N_8018,N_8702);
nor U9165 (N_9165,N_8423,N_8204);
nor U9166 (N_9166,N_8367,N_8908);
nor U9167 (N_9167,N_8574,N_8556);
or U9168 (N_9168,N_8826,N_8566);
nor U9169 (N_9169,N_8094,N_8909);
nand U9170 (N_9170,N_8223,N_8557);
nor U9171 (N_9171,N_8338,N_8625);
nor U9172 (N_9172,N_8086,N_8387);
nand U9173 (N_9173,N_8140,N_8545);
nor U9174 (N_9174,N_8268,N_8511);
and U9175 (N_9175,N_8844,N_8947);
or U9176 (N_9176,N_8035,N_8586);
or U9177 (N_9177,N_8658,N_8959);
nor U9178 (N_9178,N_8416,N_8245);
nor U9179 (N_9179,N_8569,N_8211);
nor U9180 (N_9180,N_8405,N_8255);
nor U9181 (N_9181,N_8175,N_8467);
and U9182 (N_9182,N_8797,N_8764);
and U9183 (N_9183,N_8158,N_8425);
nor U9184 (N_9184,N_8803,N_8728);
or U9185 (N_9185,N_8572,N_8426);
or U9186 (N_9186,N_8599,N_8977);
nor U9187 (N_9187,N_8430,N_8699);
and U9188 (N_9188,N_8505,N_8735);
nor U9189 (N_9189,N_8122,N_8716);
nor U9190 (N_9190,N_8288,N_8602);
xor U9191 (N_9191,N_8688,N_8377);
nor U9192 (N_9192,N_8614,N_8182);
and U9193 (N_9193,N_8806,N_8729);
or U9194 (N_9194,N_8012,N_8141);
and U9195 (N_9195,N_8627,N_8325);
or U9196 (N_9196,N_8229,N_8080);
or U9197 (N_9197,N_8644,N_8732);
nor U9198 (N_9198,N_8295,N_8342);
and U9199 (N_9199,N_8143,N_8008);
xnor U9200 (N_9200,N_8810,N_8664);
or U9201 (N_9201,N_8978,N_8240);
nor U9202 (N_9202,N_8884,N_8531);
and U9203 (N_9203,N_8905,N_8249);
nor U9204 (N_9204,N_8897,N_8500);
or U9205 (N_9205,N_8923,N_8498);
nor U9206 (N_9206,N_8270,N_8676);
nand U9207 (N_9207,N_8544,N_8568);
and U9208 (N_9208,N_8787,N_8555);
and U9209 (N_9209,N_8282,N_8281);
nand U9210 (N_9210,N_8257,N_8050);
or U9211 (N_9211,N_8683,N_8671);
or U9212 (N_9212,N_8451,N_8861);
nor U9213 (N_9213,N_8480,N_8219);
or U9214 (N_9214,N_8956,N_8232);
and U9215 (N_9215,N_8726,N_8284);
nand U9216 (N_9216,N_8241,N_8891);
and U9217 (N_9217,N_8137,N_8462);
or U9218 (N_9218,N_8573,N_8341);
nand U9219 (N_9219,N_8953,N_8630);
nor U9220 (N_9220,N_8404,N_8704);
and U9221 (N_9221,N_8457,N_8936);
nand U9222 (N_9222,N_8296,N_8899);
nand U9223 (N_9223,N_8651,N_8622);
or U9224 (N_9224,N_8275,N_8402);
nor U9225 (N_9225,N_8534,N_8460);
nand U9226 (N_9226,N_8199,N_8030);
and U9227 (N_9227,N_8477,N_8420);
nor U9228 (N_9228,N_8227,N_8129);
nand U9229 (N_9229,N_8029,N_8656);
nor U9230 (N_9230,N_8017,N_8885);
and U9231 (N_9231,N_8938,N_8629);
and U9232 (N_9232,N_8811,N_8931);
and U9233 (N_9233,N_8892,N_8311);
nand U9234 (N_9234,N_8485,N_8072);
and U9235 (N_9235,N_8540,N_8828);
or U9236 (N_9236,N_8560,N_8169);
nand U9237 (N_9237,N_8145,N_8913);
nand U9238 (N_9238,N_8766,N_8279);
and U9239 (N_9239,N_8339,N_8945);
nand U9240 (N_9240,N_8705,N_8261);
or U9241 (N_9241,N_8533,N_8039);
nor U9242 (N_9242,N_8701,N_8023);
or U9243 (N_9243,N_8591,N_8999);
or U9244 (N_9244,N_8748,N_8769);
nor U9245 (N_9245,N_8099,N_8835);
nand U9246 (N_9246,N_8274,N_8247);
or U9247 (N_9247,N_8889,N_8033);
or U9248 (N_9248,N_8867,N_8876);
or U9249 (N_9249,N_8660,N_8832);
nand U9250 (N_9250,N_8646,N_8964);
and U9251 (N_9251,N_8256,N_8051);
and U9252 (N_9252,N_8333,N_8363);
and U9253 (N_9253,N_8823,N_8258);
and U9254 (N_9254,N_8502,N_8916);
nand U9255 (N_9255,N_8097,N_8967);
nand U9256 (N_9256,N_8329,N_8055);
nor U9257 (N_9257,N_8004,N_8727);
or U9258 (N_9258,N_8239,N_8654);
or U9259 (N_9259,N_8715,N_8066);
nor U9260 (N_9260,N_8525,N_8929);
nand U9261 (N_9261,N_8695,N_8987);
nor U9262 (N_9262,N_8484,N_8626);
and U9263 (N_9263,N_8522,N_8670);
or U9264 (N_9264,N_8761,N_8910);
nand U9265 (N_9265,N_8077,N_8376);
and U9266 (N_9266,N_8809,N_8973);
and U9267 (N_9267,N_8049,N_8014);
and U9268 (N_9268,N_8666,N_8997);
or U9269 (N_9269,N_8440,N_8866);
nand U9270 (N_9270,N_8736,N_8743);
nor U9271 (N_9271,N_8647,N_8346);
and U9272 (N_9272,N_8466,N_8788);
and U9273 (N_9273,N_8604,N_8078);
and U9274 (N_9274,N_8717,N_8757);
nand U9275 (N_9275,N_8613,N_8935);
nand U9276 (N_9276,N_8162,N_8763);
or U9277 (N_9277,N_8108,N_8234);
nor U9278 (N_9278,N_8771,N_8576);
and U9279 (N_9279,N_8624,N_8655);
and U9280 (N_9280,N_8061,N_8138);
nor U9281 (N_9281,N_8872,N_8971);
nor U9282 (N_9282,N_8841,N_8740);
and U9283 (N_9283,N_8010,N_8693);
nor U9284 (N_9284,N_8836,N_8780);
nand U9285 (N_9285,N_8914,N_8037);
nand U9286 (N_9286,N_8490,N_8388);
nor U9287 (N_9287,N_8643,N_8981);
nand U9288 (N_9288,N_8496,N_8383);
or U9289 (N_9289,N_8952,N_8177);
nor U9290 (N_9290,N_8007,N_8272);
nor U9291 (N_9291,N_8961,N_8096);
and U9292 (N_9292,N_8128,N_8720);
nand U9293 (N_9293,N_8768,N_8503);
and U9294 (N_9294,N_8657,N_8351);
nand U9295 (N_9295,N_8675,N_8513);
nand U9296 (N_9296,N_8542,N_8216);
or U9297 (N_9297,N_8888,N_8864);
nand U9298 (N_9298,N_8350,N_8665);
nor U9299 (N_9299,N_8855,N_8119);
nor U9300 (N_9300,N_8917,N_8585);
nor U9301 (N_9301,N_8316,N_8731);
nor U9302 (N_9302,N_8449,N_8714);
or U9303 (N_9303,N_8125,N_8882);
nor U9304 (N_9304,N_8378,N_8392);
nor U9305 (N_9305,N_8372,N_8597);
and U9306 (N_9306,N_8612,N_8025);
and U9307 (N_9307,N_8820,N_8276);
nor U9308 (N_9308,N_8244,N_8984);
and U9309 (N_9309,N_8770,N_8068);
or U9310 (N_9310,N_8805,N_8318);
nor U9311 (N_9311,N_8514,N_8886);
or U9312 (N_9312,N_8121,N_8040);
or U9313 (N_9313,N_8491,N_8543);
and U9314 (N_9314,N_8045,N_8206);
or U9315 (N_9315,N_8434,N_8359);
and U9316 (N_9316,N_8043,N_8874);
nor U9317 (N_9317,N_8225,N_8000);
nor U9318 (N_9318,N_8827,N_8450);
and U9319 (N_9319,N_8321,N_8439);
nand U9320 (N_9320,N_8696,N_8603);
nor U9321 (N_9321,N_8972,N_8982);
nor U9322 (N_9322,N_8222,N_8142);
or U9323 (N_9323,N_8253,N_8746);
nor U9324 (N_9324,N_8880,N_8907);
or U9325 (N_9325,N_8428,N_8942);
or U9326 (N_9326,N_8915,N_8200);
nor U9327 (N_9327,N_8127,N_8027);
nor U9328 (N_9328,N_8663,N_8381);
or U9329 (N_9329,N_8846,N_8741);
and U9330 (N_9330,N_8593,N_8303);
nor U9331 (N_9331,N_8117,N_8881);
and U9332 (N_9332,N_8100,N_8149);
nor U9333 (N_9333,N_8998,N_8765);
and U9334 (N_9334,N_8824,N_8192);
nor U9335 (N_9335,N_8516,N_8718);
and U9336 (N_9336,N_8259,N_8950);
and U9337 (N_9337,N_8802,N_8064);
nor U9338 (N_9338,N_8293,N_8812);
or U9339 (N_9339,N_8887,N_8210);
nand U9340 (N_9340,N_8759,N_8290);
nor U9341 (N_9341,N_8208,N_8659);
nor U9342 (N_9342,N_8988,N_8709);
nand U9343 (N_9343,N_8611,N_8930);
nor U9344 (N_9344,N_8390,N_8723);
and U9345 (N_9345,N_8600,N_8506);
and U9346 (N_9346,N_8551,N_8650);
nand U9347 (N_9347,N_8773,N_8226);
nor U9348 (N_9348,N_8890,N_8419);
nand U9349 (N_9349,N_8344,N_8549);
or U9350 (N_9350,N_8470,N_8476);
or U9351 (N_9351,N_8181,N_8184);
nor U9352 (N_9352,N_8313,N_8845);
and U9353 (N_9353,N_8020,N_8970);
nor U9354 (N_9354,N_8421,N_8380);
or U9355 (N_9355,N_8801,N_8519);
nand U9356 (N_9356,N_8598,N_8524);
nand U9357 (N_9357,N_8842,N_8530);
nand U9358 (N_9358,N_8995,N_8685);
nand U9359 (N_9359,N_8106,N_8927);
or U9360 (N_9360,N_8429,N_8431);
nor U9361 (N_9361,N_8207,N_8164);
or U9362 (N_9362,N_8468,N_8424);
nor U9363 (N_9363,N_8933,N_8155);
and U9364 (N_9364,N_8928,N_8300);
nor U9365 (N_9365,N_8085,N_8335);
nor U9366 (N_9366,N_8582,N_8446);
nand U9367 (N_9367,N_8366,N_8151);
or U9368 (N_9368,N_8159,N_8076);
or U9369 (N_9369,N_8170,N_8079);
nor U9370 (N_9370,N_8674,N_8552);
and U9371 (N_9371,N_8120,N_8737);
and U9372 (N_9372,N_8774,N_8443);
or U9373 (N_9373,N_8690,N_8903);
and U9374 (N_9374,N_8968,N_8075);
and U9375 (N_9375,N_8989,N_8063);
nand U9376 (N_9376,N_8508,N_8817);
and U9377 (N_9377,N_8292,N_8231);
nor U9378 (N_9378,N_8677,N_8859);
nor U9379 (N_9379,N_8198,N_8641);
or U9380 (N_9380,N_8849,N_8616);
nand U9381 (N_9381,N_8815,N_8406);
or U9382 (N_9382,N_8442,N_8441);
nand U9383 (N_9383,N_8990,N_8228);
and U9384 (N_9384,N_8577,N_8957);
or U9385 (N_9385,N_8088,N_8951);
nand U9386 (N_9386,N_8507,N_8394);
and U9387 (N_9387,N_8134,N_8784);
nand U9388 (N_9388,N_8515,N_8589);
nand U9389 (N_9389,N_8777,N_8087);
nor U9390 (N_9390,N_8790,N_8269);
and U9391 (N_9391,N_8587,N_8320);
nand U9392 (N_9392,N_8821,N_8965);
or U9393 (N_9393,N_8575,N_8722);
or U9394 (N_9394,N_8645,N_8474);
nand U9395 (N_9395,N_8403,N_8607);
nand U9396 (N_9396,N_8561,N_8848);
and U9397 (N_9397,N_8920,N_8009);
nor U9398 (N_9398,N_8581,N_8368);
or U9399 (N_9399,N_8986,N_8452);
nor U9400 (N_9400,N_8799,N_8448);
and U9401 (N_9401,N_8115,N_8755);
nand U9402 (N_9402,N_8286,N_8662);
nand U9403 (N_9403,N_8413,N_8073);
and U9404 (N_9404,N_8776,N_8943);
nand U9405 (N_9405,N_8152,N_8550);
or U9406 (N_9406,N_8563,N_8337);
and U9407 (N_9407,N_8136,N_8994);
nor U9408 (N_9408,N_8264,N_8580);
nand U9409 (N_9409,N_8517,N_8609);
or U9410 (N_9410,N_8640,N_8745);
or U9411 (N_9411,N_8179,N_8919);
nor U9412 (N_9412,N_8794,N_8567);
or U9413 (N_9413,N_8180,N_8749);
or U9414 (N_9414,N_8056,N_8786);
nor U9415 (N_9415,N_8102,N_8150);
nand U9416 (N_9416,N_8324,N_8649);
nand U9417 (N_9417,N_8960,N_8783);
or U9418 (N_9418,N_8710,N_8437);
nand U9419 (N_9419,N_8538,N_8762);
nand U9420 (N_9420,N_8847,N_8993);
nor U9421 (N_9421,N_8370,N_8212);
nor U9422 (N_9422,N_8397,N_8772);
or U9423 (N_9423,N_8877,N_8189);
and U9424 (N_9424,N_8830,N_8328);
and U9425 (N_9425,N_8661,N_8969);
and U9426 (N_9426,N_8302,N_8495);
nor U9427 (N_9427,N_8254,N_8139);
nand U9428 (N_9428,N_8708,N_8432);
nor U9429 (N_9429,N_8465,N_8041);
and U9430 (N_9430,N_8648,N_8825);
nor U9431 (N_9431,N_8932,N_8057);
and U9432 (N_9432,N_8541,N_8721);
and U9433 (N_9433,N_8532,N_8852);
nor U9434 (N_9434,N_8165,N_8399);
and U9435 (N_9435,N_8265,N_8060);
or U9436 (N_9436,N_8065,N_8319);
nand U9437 (N_9437,N_8445,N_8837);
nor U9438 (N_9438,N_8156,N_8678);
and U9439 (N_9439,N_8504,N_8883);
or U9440 (N_9440,N_8348,N_8191);
nand U9441 (N_9441,N_8488,N_8396);
or U9442 (N_9442,N_8183,N_8921);
nand U9443 (N_9443,N_8187,N_8048);
nor U9444 (N_9444,N_8185,N_8148);
or U9445 (N_9445,N_8201,N_8132);
nand U9446 (N_9446,N_8588,N_8497);
or U9447 (N_9447,N_8082,N_8878);
nor U9448 (N_9448,N_8371,N_8800);
or U9449 (N_9449,N_8934,N_8902);
or U9450 (N_9450,N_8036,N_8789);
and U9451 (N_9451,N_8601,N_8668);
nor U9452 (N_9452,N_8271,N_8301);
and U9453 (N_9453,N_8438,N_8172);
nand U9454 (N_9454,N_8739,N_8163);
nor U9455 (N_9455,N_8554,N_8767);
and U9456 (N_9456,N_8785,N_8911);
or U9457 (N_9457,N_8308,N_8991);
and U9458 (N_9458,N_8110,N_8190);
and U9459 (N_9459,N_8196,N_8672);
and U9460 (N_9460,N_8681,N_8273);
nand U9461 (N_9461,N_8375,N_8719);
nand U9462 (N_9462,N_8124,N_8558);
nand U9463 (N_9463,N_8217,N_8623);
nor U9464 (N_9464,N_8160,N_8918);
and U9465 (N_9465,N_8526,N_8955);
nand U9466 (N_9466,N_8750,N_8752);
nor U9467 (N_9467,N_8792,N_8015);
or U9468 (N_9468,N_8979,N_8680);
and U9469 (N_9469,N_8521,N_8400);
or U9470 (N_9470,N_8144,N_8742);
nand U9471 (N_9471,N_8873,N_8243);
nand U9472 (N_9472,N_8135,N_8361);
or U9473 (N_9473,N_8992,N_8130);
nor U9474 (N_9474,N_8323,N_8047);
nor U9475 (N_9475,N_8758,N_8754);
and U9476 (N_9476,N_8307,N_8896);
or U9477 (N_9477,N_8021,N_8278);
or U9478 (N_9478,N_8834,N_8472);
or U9479 (N_9479,N_8653,N_8958);
and U9480 (N_9480,N_8547,N_8734);
and U9481 (N_9481,N_8865,N_8084);
nor U9482 (N_9482,N_8360,N_8412);
nand U9483 (N_9483,N_8831,N_8482);
nand U9484 (N_9484,N_8711,N_8003);
nand U9485 (N_9485,N_8940,N_8944);
nand U9486 (N_9486,N_8937,N_8202);
nor U9487 (N_9487,N_8620,N_8633);
or U9488 (N_9488,N_8926,N_8306);
nand U9489 (N_9489,N_8113,N_8331);
or U9490 (N_9490,N_8277,N_8839);
or U9491 (N_9491,N_8090,N_8528);
or U9492 (N_9492,N_8840,N_8536);
and U9493 (N_9493,N_8860,N_8104);
nand U9494 (N_9494,N_8868,N_8610);
or U9495 (N_9495,N_8305,N_8154);
and U9496 (N_9496,N_8123,N_8996);
and U9497 (N_9497,N_8188,N_8299);
nand U9498 (N_9498,N_8804,N_8098);
or U9499 (N_9499,N_8298,N_8103);
and U9500 (N_9500,N_8945,N_8653);
nor U9501 (N_9501,N_8319,N_8280);
nor U9502 (N_9502,N_8300,N_8548);
or U9503 (N_9503,N_8219,N_8760);
nand U9504 (N_9504,N_8241,N_8470);
nand U9505 (N_9505,N_8923,N_8039);
and U9506 (N_9506,N_8183,N_8047);
nand U9507 (N_9507,N_8036,N_8430);
nor U9508 (N_9508,N_8177,N_8040);
and U9509 (N_9509,N_8655,N_8045);
or U9510 (N_9510,N_8976,N_8148);
and U9511 (N_9511,N_8396,N_8248);
nand U9512 (N_9512,N_8708,N_8379);
nand U9513 (N_9513,N_8171,N_8081);
nand U9514 (N_9514,N_8193,N_8987);
nand U9515 (N_9515,N_8238,N_8862);
and U9516 (N_9516,N_8488,N_8567);
nor U9517 (N_9517,N_8479,N_8637);
nand U9518 (N_9518,N_8820,N_8322);
nand U9519 (N_9519,N_8289,N_8881);
or U9520 (N_9520,N_8997,N_8152);
or U9521 (N_9521,N_8506,N_8444);
nand U9522 (N_9522,N_8699,N_8443);
nor U9523 (N_9523,N_8357,N_8343);
and U9524 (N_9524,N_8861,N_8977);
or U9525 (N_9525,N_8889,N_8140);
or U9526 (N_9526,N_8488,N_8981);
nor U9527 (N_9527,N_8202,N_8913);
nor U9528 (N_9528,N_8851,N_8826);
nor U9529 (N_9529,N_8261,N_8486);
nand U9530 (N_9530,N_8758,N_8187);
and U9531 (N_9531,N_8879,N_8985);
nor U9532 (N_9532,N_8495,N_8574);
and U9533 (N_9533,N_8051,N_8465);
nor U9534 (N_9534,N_8213,N_8115);
nor U9535 (N_9535,N_8825,N_8704);
or U9536 (N_9536,N_8170,N_8136);
and U9537 (N_9537,N_8765,N_8987);
nand U9538 (N_9538,N_8431,N_8074);
nand U9539 (N_9539,N_8300,N_8900);
or U9540 (N_9540,N_8399,N_8996);
nand U9541 (N_9541,N_8260,N_8208);
nor U9542 (N_9542,N_8269,N_8064);
or U9543 (N_9543,N_8971,N_8781);
and U9544 (N_9544,N_8800,N_8770);
nor U9545 (N_9545,N_8135,N_8302);
nand U9546 (N_9546,N_8321,N_8746);
and U9547 (N_9547,N_8121,N_8216);
and U9548 (N_9548,N_8152,N_8208);
and U9549 (N_9549,N_8077,N_8640);
nand U9550 (N_9550,N_8472,N_8333);
or U9551 (N_9551,N_8591,N_8057);
or U9552 (N_9552,N_8515,N_8828);
nor U9553 (N_9553,N_8841,N_8671);
nand U9554 (N_9554,N_8855,N_8384);
nand U9555 (N_9555,N_8707,N_8675);
or U9556 (N_9556,N_8942,N_8494);
and U9557 (N_9557,N_8528,N_8428);
nand U9558 (N_9558,N_8642,N_8824);
nand U9559 (N_9559,N_8544,N_8444);
nand U9560 (N_9560,N_8160,N_8466);
or U9561 (N_9561,N_8360,N_8278);
nor U9562 (N_9562,N_8412,N_8532);
and U9563 (N_9563,N_8993,N_8829);
or U9564 (N_9564,N_8157,N_8290);
nor U9565 (N_9565,N_8626,N_8508);
or U9566 (N_9566,N_8168,N_8776);
nor U9567 (N_9567,N_8513,N_8118);
nand U9568 (N_9568,N_8389,N_8896);
nor U9569 (N_9569,N_8932,N_8807);
and U9570 (N_9570,N_8484,N_8420);
and U9571 (N_9571,N_8777,N_8486);
nand U9572 (N_9572,N_8672,N_8743);
and U9573 (N_9573,N_8794,N_8695);
nand U9574 (N_9574,N_8796,N_8360);
nor U9575 (N_9575,N_8526,N_8444);
and U9576 (N_9576,N_8575,N_8037);
nor U9577 (N_9577,N_8712,N_8512);
or U9578 (N_9578,N_8268,N_8805);
and U9579 (N_9579,N_8805,N_8391);
or U9580 (N_9580,N_8823,N_8443);
nand U9581 (N_9581,N_8235,N_8208);
xor U9582 (N_9582,N_8514,N_8075);
or U9583 (N_9583,N_8899,N_8228);
nand U9584 (N_9584,N_8292,N_8814);
nand U9585 (N_9585,N_8049,N_8294);
and U9586 (N_9586,N_8899,N_8194);
and U9587 (N_9587,N_8305,N_8269);
or U9588 (N_9588,N_8586,N_8118);
and U9589 (N_9589,N_8224,N_8534);
and U9590 (N_9590,N_8383,N_8097);
or U9591 (N_9591,N_8798,N_8956);
nand U9592 (N_9592,N_8614,N_8063);
nor U9593 (N_9593,N_8292,N_8034);
nor U9594 (N_9594,N_8618,N_8979);
nand U9595 (N_9595,N_8258,N_8982);
or U9596 (N_9596,N_8756,N_8137);
nand U9597 (N_9597,N_8502,N_8579);
nand U9598 (N_9598,N_8402,N_8114);
and U9599 (N_9599,N_8566,N_8380);
nand U9600 (N_9600,N_8409,N_8259);
nand U9601 (N_9601,N_8701,N_8539);
and U9602 (N_9602,N_8525,N_8061);
nor U9603 (N_9603,N_8472,N_8611);
and U9604 (N_9604,N_8175,N_8662);
and U9605 (N_9605,N_8294,N_8522);
or U9606 (N_9606,N_8507,N_8562);
and U9607 (N_9607,N_8474,N_8340);
or U9608 (N_9608,N_8143,N_8071);
and U9609 (N_9609,N_8938,N_8032);
or U9610 (N_9610,N_8635,N_8610);
and U9611 (N_9611,N_8788,N_8682);
nor U9612 (N_9612,N_8595,N_8369);
nand U9613 (N_9613,N_8283,N_8551);
and U9614 (N_9614,N_8028,N_8525);
nor U9615 (N_9615,N_8362,N_8558);
and U9616 (N_9616,N_8065,N_8715);
nor U9617 (N_9617,N_8899,N_8746);
nor U9618 (N_9618,N_8634,N_8286);
or U9619 (N_9619,N_8604,N_8274);
or U9620 (N_9620,N_8521,N_8265);
nand U9621 (N_9621,N_8384,N_8481);
and U9622 (N_9622,N_8076,N_8604);
or U9623 (N_9623,N_8171,N_8595);
nand U9624 (N_9624,N_8812,N_8628);
nor U9625 (N_9625,N_8430,N_8775);
nand U9626 (N_9626,N_8470,N_8872);
and U9627 (N_9627,N_8091,N_8840);
or U9628 (N_9628,N_8799,N_8411);
or U9629 (N_9629,N_8456,N_8291);
xnor U9630 (N_9630,N_8120,N_8972);
nand U9631 (N_9631,N_8282,N_8852);
nand U9632 (N_9632,N_8116,N_8779);
and U9633 (N_9633,N_8707,N_8601);
nor U9634 (N_9634,N_8599,N_8011);
and U9635 (N_9635,N_8677,N_8954);
and U9636 (N_9636,N_8771,N_8613);
or U9637 (N_9637,N_8983,N_8905);
nor U9638 (N_9638,N_8037,N_8230);
nor U9639 (N_9639,N_8510,N_8527);
or U9640 (N_9640,N_8015,N_8436);
nor U9641 (N_9641,N_8209,N_8435);
and U9642 (N_9642,N_8331,N_8925);
and U9643 (N_9643,N_8531,N_8876);
or U9644 (N_9644,N_8492,N_8471);
nand U9645 (N_9645,N_8224,N_8060);
and U9646 (N_9646,N_8329,N_8278);
or U9647 (N_9647,N_8804,N_8935);
nand U9648 (N_9648,N_8504,N_8148);
nand U9649 (N_9649,N_8090,N_8702);
nor U9650 (N_9650,N_8682,N_8018);
and U9651 (N_9651,N_8287,N_8892);
or U9652 (N_9652,N_8233,N_8840);
nor U9653 (N_9653,N_8034,N_8878);
nor U9654 (N_9654,N_8627,N_8451);
nor U9655 (N_9655,N_8841,N_8484);
nor U9656 (N_9656,N_8235,N_8245);
nor U9657 (N_9657,N_8553,N_8599);
or U9658 (N_9658,N_8654,N_8052);
nor U9659 (N_9659,N_8960,N_8655);
nand U9660 (N_9660,N_8548,N_8485);
or U9661 (N_9661,N_8939,N_8009);
nand U9662 (N_9662,N_8157,N_8837);
nand U9663 (N_9663,N_8810,N_8782);
or U9664 (N_9664,N_8480,N_8843);
nor U9665 (N_9665,N_8622,N_8992);
nand U9666 (N_9666,N_8339,N_8583);
and U9667 (N_9667,N_8600,N_8284);
or U9668 (N_9668,N_8146,N_8885);
or U9669 (N_9669,N_8524,N_8621);
nand U9670 (N_9670,N_8850,N_8616);
nor U9671 (N_9671,N_8200,N_8513);
and U9672 (N_9672,N_8123,N_8780);
and U9673 (N_9673,N_8419,N_8169);
and U9674 (N_9674,N_8952,N_8152);
nand U9675 (N_9675,N_8840,N_8360);
or U9676 (N_9676,N_8668,N_8485);
and U9677 (N_9677,N_8033,N_8857);
nand U9678 (N_9678,N_8791,N_8277);
and U9679 (N_9679,N_8854,N_8975);
and U9680 (N_9680,N_8729,N_8548);
or U9681 (N_9681,N_8546,N_8114);
or U9682 (N_9682,N_8509,N_8708);
and U9683 (N_9683,N_8531,N_8762);
nand U9684 (N_9684,N_8143,N_8631);
nand U9685 (N_9685,N_8123,N_8345);
nor U9686 (N_9686,N_8172,N_8942);
nand U9687 (N_9687,N_8893,N_8585);
and U9688 (N_9688,N_8676,N_8689);
nand U9689 (N_9689,N_8368,N_8119);
nand U9690 (N_9690,N_8523,N_8558);
nand U9691 (N_9691,N_8747,N_8484);
or U9692 (N_9692,N_8596,N_8166);
nor U9693 (N_9693,N_8479,N_8239);
and U9694 (N_9694,N_8323,N_8756);
and U9695 (N_9695,N_8240,N_8783);
nand U9696 (N_9696,N_8513,N_8734);
nor U9697 (N_9697,N_8421,N_8995);
or U9698 (N_9698,N_8330,N_8278);
nor U9699 (N_9699,N_8649,N_8552);
or U9700 (N_9700,N_8762,N_8950);
or U9701 (N_9701,N_8379,N_8660);
or U9702 (N_9702,N_8819,N_8976);
nand U9703 (N_9703,N_8468,N_8033);
and U9704 (N_9704,N_8944,N_8051);
or U9705 (N_9705,N_8785,N_8643);
nor U9706 (N_9706,N_8031,N_8184);
nor U9707 (N_9707,N_8165,N_8865);
and U9708 (N_9708,N_8254,N_8479);
nor U9709 (N_9709,N_8900,N_8925);
nor U9710 (N_9710,N_8198,N_8228);
nor U9711 (N_9711,N_8660,N_8651);
and U9712 (N_9712,N_8687,N_8320);
or U9713 (N_9713,N_8850,N_8040);
nand U9714 (N_9714,N_8840,N_8372);
or U9715 (N_9715,N_8765,N_8616);
nand U9716 (N_9716,N_8838,N_8451);
and U9717 (N_9717,N_8944,N_8933);
and U9718 (N_9718,N_8541,N_8620);
and U9719 (N_9719,N_8662,N_8281);
nand U9720 (N_9720,N_8155,N_8298);
or U9721 (N_9721,N_8443,N_8469);
nor U9722 (N_9722,N_8931,N_8822);
nor U9723 (N_9723,N_8572,N_8731);
or U9724 (N_9724,N_8974,N_8078);
nor U9725 (N_9725,N_8847,N_8469);
nor U9726 (N_9726,N_8283,N_8829);
or U9727 (N_9727,N_8735,N_8785);
or U9728 (N_9728,N_8090,N_8311);
and U9729 (N_9729,N_8230,N_8023);
nand U9730 (N_9730,N_8056,N_8527);
or U9731 (N_9731,N_8137,N_8504);
and U9732 (N_9732,N_8594,N_8542);
and U9733 (N_9733,N_8327,N_8424);
nand U9734 (N_9734,N_8645,N_8103);
or U9735 (N_9735,N_8697,N_8903);
or U9736 (N_9736,N_8089,N_8493);
xor U9737 (N_9737,N_8665,N_8238);
nand U9738 (N_9738,N_8758,N_8039);
nor U9739 (N_9739,N_8294,N_8513);
nor U9740 (N_9740,N_8481,N_8169);
nor U9741 (N_9741,N_8707,N_8595);
or U9742 (N_9742,N_8706,N_8633);
nor U9743 (N_9743,N_8510,N_8818);
or U9744 (N_9744,N_8416,N_8827);
nand U9745 (N_9745,N_8073,N_8935);
nor U9746 (N_9746,N_8745,N_8065);
and U9747 (N_9747,N_8709,N_8350);
nor U9748 (N_9748,N_8448,N_8373);
or U9749 (N_9749,N_8720,N_8135);
and U9750 (N_9750,N_8072,N_8699);
nand U9751 (N_9751,N_8706,N_8969);
or U9752 (N_9752,N_8654,N_8694);
nor U9753 (N_9753,N_8567,N_8589);
or U9754 (N_9754,N_8280,N_8817);
nor U9755 (N_9755,N_8559,N_8655);
and U9756 (N_9756,N_8395,N_8913);
nor U9757 (N_9757,N_8103,N_8834);
nand U9758 (N_9758,N_8687,N_8022);
nand U9759 (N_9759,N_8137,N_8097);
and U9760 (N_9760,N_8669,N_8028);
nand U9761 (N_9761,N_8582,N_8639);
nand U9762 (N_9762,N_8336,N_8744);
or U9763 (N_9763,N_8499,N_8557);
nor U9764 (N_9764,N_8241,N_8444);
and U9765 (N_9765,N_8374,N_8247);
nand U9766 (N_9766,N_8855,N_8142);
nor U9767 (N_9767,N_8734,N_8058);
nor U9768 (N_9768,N_8981,N_8771);
nand U9769 (N_9769,N_8343,N_8727);
and U9770 (N_9770,N_8532,N_8297);
or U9771 (N_9771,N_8822,N_8252);
or U9772 (N_9772,N_8445,N_8874);
and U9773 (N_9773,N_8298,N_8816);
and U9774 (N_9774,N_8500,N_8763);
nand U9775 (N_9775,N_8876,N_8643);
or U9776 (N_9776,N_8313,N_8171);
and U9777 (N_9777,N_8951,N_8182);
nand U9778 (N_9778,N_8444,N_8745);
nor U9779 (N_9779,N_8680,N_8244);
or U9780 (N_9780,N_8260,N_8697);
and U9781 (N_9781,N_8081,N_8927);
nand U9782 (N_9782,N_8440,N_8683);
nor U9783 (N_9783,N_8470,N_8633);
nor U9784 (N_9784,N_8365,N_8920);
nor U9785 (N_9785,N_8621,N_8778);
nand U9786 (N_9786,N_8484,N_8849);
and U9787 (N_9787,N_8109,N_8860);
nand U9788 (N_9788,N_8071,N_8628);
nor U9789 (N_9789,N_8204,N_8262);
and U9790 (N_9790,N_8377,N_8293);
or U9791 (N_9791,N_8786,N_8790);
or U9792 (N_9792,N_8539,N_8500);
nand U9793 (N_9793,N_8430,N_8689);
and U9794 (N_9794,N_8921,N_8086);
nor U9795 (N_9795,N_8439,N_8798);
nand U9796 (N_9796,N_8641,N_8949);
and U9797 (N_9797,N_8548,N_8133);
and U9798 (N_9798,N_8352,N_8178);
or U9799 (N_9799,N_8701,N_8641);
and U9800 (N_9800,N_8454,N_8817);
nand U9801 (N_9801,N_8469,N_8751);
and U9802 (N_9802,N_8530,N_8498);
nand U9803 (N_9803,N_8852,N_8183);
nand U9804 (N_9804,N_8799,N_8148);
nand U9805 (N_9805,N_8154,N_8952);
nor U9806 (N_9806,N_8168,N_8381);
and U9807 (N_9807,N_8946,N_8771);
and U9808 (N_9808,N_8503,N_8017);
or U9809 (N_9809,N_8934,N_8615);
nor U9810 (N_9810,N_8256,N_8787);
and U9811 (N_9811,N_8989,N_8056);
nor U9812 (N_9812,N_8915,N_8380);
and U9813 (N_9813,N_8072,N_8866);
nor U9814 (N_9814,N_8589,N_8548);
xnor U9815 (N_9815,N_8125,N_8388);
nand U9816 (N_9816,N_8480,N_8994);
nand U9817 (N_9817,N_8946,N_8504);
nand U9818 (N_9818,N_8610,N_8520);
nand U9819 (N_9819,N_8504,N_8758);
nand U9820 (N_9820,N_8082,N_8487);
or U9821 (N_9821,N_8106,N_8293);
and U9822 (N_9822,N_8951,N_8552);
xor U9823 (N_9823,N_8820,N_8924);
nand U9824 (N_9824,N_8917,N_8998);
nor U9825 (N_9825,N_8703,N_8197);
nor U9826 (N_9826,N_8708,N_8503);
nor U9827 (N_9827,N_8890,N_8444);
or U9828 (N_9828,N_8806,N_8679);
or U9829 (N_9829,N_8390,N_8439);
nor U9830 (N_9830,N_8195,N_8508);
or U9831 (N_9831,N_8813,N_8107);
nand U9832 (N_9832,N_8132,N_8348);
nor U9833 (N_9833,N_8415,N_8242);
nor U9834 (N_9834,N_8004,N_8165);
and U9835 (N_9835,N_8506,N_8745);
nand U9836 (N_9836,N_8152,N_8583);
nand U9837 (N_9837,N_8200,N_8036);
or U9838 (N_9838,N_8720,N_8799);
nand U9839 (N_9839,N_8421,N_8239);
or U9840 (N_9840,N_8484,N_8055);
nor U9841 (N_9841,N_8588,N_8743);
nor U9842 (N_9842,N_8154,N_8474);
or U9843 (N_9843,N_8615,N_8323);
nand U9844 (N_9844,N_8855,N_8652);
nand U9845 (N_9845,N_8609,N_8115);
and U9846 (N_9846,N_8485,N_8371);
nand U9847 (N_9847,N_8573,N_8997);
nand U9848 (N_9848,N_8353,N_8256);
nand U9849 (N_9849,N_8373,N_8691);
nand U9850 (N_9850,N_8656,N_8464);
or U9851 (N_9851,N_8987,N_8154);
nor U9852 (N_9852,N_8720,N_8204);
nand U9853 (N_9853,N_8599,N_8942);
nand U9854 (N_9854,N_8802,N_8271);
or U9855 (N_9855,N_8202,N_8218);
nand U9856 (N_9856,N_8019,N_8026);
and U9857 (N_9857,N_8877,N_8779);
nand U9858 (N_9858,N_8637,N_8070);
xnor U9859 (N_9859,N_8806,N_8912);
or U9860 (N_9860,N_8412,N_8361);
or U9861 (N_9861,N_8188,N_8876);
nand U9862 (N_9862,N_8946,N_8548);
or U9863 (N_9863,N_8954,N_8973);
nor U9864 (N_9864,N_8277,N_8835);
or U9865 (N_9865,N_8624,N_8539);
or U9866 (N_9866,N_8187,N_8222);
nand U9867 (N_9867,N_8189,N_8597);
nand U9868 (N_9868,N_8051,N_8839);
and U9869 (N_9869,N_8199,N_8460);
nor U9870 (N_9870,N_8586,N_8538);
nor U9871 (N_9871,N_8317,N_8073);
or U9872 (N_9872,N_8982,N_8708);
nor U9873 (N_9873,N_8576,N_8262);
or U9874 (N_9874,N_8411,N_8754);
and U9875 (N_9875,N_8055,N_8201);
nor U9876 (N_9876,N_8663,N_8252);
xnor U9877 (N_9877,N_8302,N_8711);
and U9878 (N_9878,N_8099,N_8075);
and U9879 (N_9879,N_8833,N_8421);
nand U9880 (N_9880,N_8497,N_8712);
nor U9881 (N_9881,N_8365,N_8637);
and U9882 (N_9882,N_8767,N_8330);
nand U9883 (N_9883,N_8064,N_8867);
and U9884 (N_9884,N_8404,N_8964);
nand U9885 (N_9885,N_8583,N_8076);
nor U9886 (N_9886,N_8066,N_8270);
or U9887 (N_9887,N_8156,N_8524);
or U9888 (N_9888,N_8601,N_8796);
and U9889 (N_9889,N_8501,N_8139);
nand U9890 (N_9890,N_8004,N_8109);
nand U9891 (N_9891,N_8509,N_8581);
nand U9892 (N_9892,N_8387,N_8831);
nor U9893 (N_9893,N_8133,N_8223);
nand U9894 (N_9894,N_8140,N_8984);
nand U9895 (N_9895,N_8937,N_8366);
nor U9896 (N_9896,N_8817,N_8863);
nor U9897 (N_9897,N_8991,N_8412);
nand U9898 (N_9898,N_8742,N_8307);
nor U9899 (N_9899,N_8091,N_8632);
nand U9900 (N_9900,N_8036,N_8691);
or U9901 (N_9901,N_8662,N_8646);
nor U9902 (N_9902,N_8694,N_8089);
nor U9903 (N_9903,N_8250,N_8691);
nor U9904 (N_9904,N_8828,N_8984);
and U9905 (N_9905,N_8675,N_8854);
or U9906 (N_9906,N_8031,N_8408);
or U9907 (N_9907,N_8092,N_8612);
and U9908 (N_9908,N_8909,N_8965);
and U9909 (N_9909,N_8834,N_8045);
or U9910 (N_9910,N_8662,N_8490);
nor U9911 (N_9911,N_8507,N_8382);
nor U9912 (N_9912,N_8409,N_8844);
or U9913 (N_9913,N_8336,N_8942);
and U9914 (N_9914,N_8423,N_8709);
nor U9915 (N_9915,N_8609,N_8788);
nor U9916 (N_9916,N_8251,N_8742);
and U9917 (N_9917,N_8538,N_8255);
nand U9918 (N_9918,N_8968,N_8594);
or U9919 (N_9919,N_8712,N_8358);
or U9920 (N_9920,N_8766,N_8555);
and U9921 (N_9921,N_8662,N_8978);
nor U9922 (N_9922,N_8234,N_8979);
and U9923 (N_9923,N_8538,N_8870);
or U9924 (N_9924,N_8029,N_8434);
nand U9925 (N_9925,N_8157,N_8679);
and U9926 (N_9926,N_8725,N_8592);
nor U9927 (N_9927,N_8910,N_8305);
and U9928 (N_9928,N_8738,N_8210);
nor U9929 (N_9929,N_8955,N_8164);
nor U9930 (N_9930,N_8715,N_8986);
and U9931 (N_9931,N_8675,N_8443);
nor U9932 (N_9932,N_8759,N_8058);
and U9933 (N_9933,N_8939,N_8330);
and U9934 (N_9934,N_8021,N_8246);
nor U9935 (N_9935,N_8959,N_8727);
and U9936 (N_9936,N_8620,N_8845);
nor U9937 (N_9937,N_8654,N_8969);
and U9938 (N_9938,N_8407,N_8699);
and U9939 (N_9939,N_8128,N_8605);
nor U9940 (N_9940,N_8364,N_8049);
or U9941 (N_9941,N_8833,N_8321);
and U9942 (N_9942,N_8518,N_8888);
nor U9943 (N_9943,N_8809,N_8615);
nor U9944 (N_9944,N_8419,N_8103);
or U9945 (N_9945,N_8363,N_8916);
nor U9946 (N_9946,N_8826,N_8247);
and U9947 (N_9947,N_8909,N_8428);
nand U9948 (N_9948,N_8281,N_8710);
or U9949 (N_9949,N_8051,N_8163);
and U9950 (N_9950,N_8354,N_8381);
and U9951 (N_9951,N_8548,N_8936);
nand U9952 (N_9952,N_8832,N_8105);
nand U9953 (N_9953,N_8414,N_8663);
nand U9954 (N_9954,N_8325,N_8942);
or U9955 (N_9955,N_8118,N_8001);
or U9956 (N_9956,N_8188,N_8432);
or U9957 (N_9957,N_8385,N_8219);
or U9958 (N_9958,N_8368,N_8257);
nor U9959 (N_9959,N_8900,N_8454);
nor U9960 (N_9960,N_8755,N_8047);
or U9961 (N_9961,N_8587,N_8548);
and U9962 (N_9962,N_8712,N_8331);
nand U9963 (N_9963,N_8295,N_8538);
nor U9964 (N_9964,N_8624,N_8087);
nor U9965 (N_9965,N_8057,N_8158);
and U9966 (N_9966,N_8089,N_8079);
or U9967 (N_9967,N_8656,N_8929);
or U9968 (N_9968,N_8212,N_8351);
nand U9969 (N_9969,N_8767,N_8275);
nor U9970 (N_9970,N_8265,N_8284);
nand U9971 (N_9971,N_8239,N_8474);
nand U9972 (N_9972,N_8058,N_8815);
and U9973 (N_9973,N_8985,N_8698);
nor U9974 (N_9974,N_8355,N_8381);
or U9975 (N_9975,N_8219,N_8842);
nor U9976 (N_9976,N_8218,N_8027);
and U9977 (N_9977,N_8143,N_8740);
and U9978 (N_9978,N_8637,N_8501);
nor U9979 (N_9979,N_8187,N_8415);
and U9980 (N_9980,N_8885,N_8596);
nand U9981 (N_9981,N_8448,N_8769);
nand U9982 (N_9982,N_8560,N_8721);
or U9983 (N_9983,N_8073,N_8872);
nand U9984 (N_9984,N_8141,N_8256);
nor U9985 (N_9985,N_8017,N_8888);
nor U9986 (N_9986,N_8170,N_8244);
or U9987 (N_9987,N_8634,N_8261);
and U9988 (N_9988,N_8594,N_8129);
or U9989 (N_9989,N_8627,N_8826);
nand U9990 (N_9990,N_8021,N_8086);
nand U9991 (N_9991,N_8645,N_8162);
nand U9992 (N_9992,N_8751,N_8010);
nor U9993 (N_9993,N_8431,N_8311);
nor U9994 (N_9994,N_8068,N_8402);
and U9995 (N_9995,N_8558,N_8288);
nor U9996 (N_9996,N_8786,N_8129);
nor U9997 (N_9997,N_8044,N_8198);
nor U9998 (N_9998,N_8935,N_8701);
nor U9999 (N_9999,N_8383,N_8762);
nand UO_0 (O_0,N_9812,N_9354);
nand UO_1 (O_1,N_9362,N_9509);
or UO_2 (O_2,N_9564,N_9542);
xnor UO_3 (O_3,N_9648,N_9809);
and UO_4 (O_4,N_9656,N_9810);
nand UO_5 (O_5,N_9008,N_9644);
and UO_6 (O_6,N_9862,N_9954);
nor UO_7 (O_7,N_9983,N_9702);
nor UO_8 (O_8,N_9156,N_9449);
and UO_9 (O_9,N_9691,N_9858);
and UO_10 (O_10,N_9334,N_9508);
nor UO_11 (O_11,N_9474,N_9063);
or UO_12 (O_12,N_9692,N_9381);
nand UO_13 (O_13,N_9207,N_9328);
nor UO_14 (O_14,N_9489,N_9382);
and UO_15 (O_15,N_9415,N_9473);
or UO_16 (O_16,N_9628,N_9853);
nand UO_17 (O_17,N_9397,N_9022);
nor UO_18 (O_18,N_9857,N_9337);
or UO_19 (O_19,N_9766,N_9392);
nand UO_20 (O_20,N_9657,N_9726);
nor UO_21 (O_21,N_9505,N_9827);
nand UO_22 (O_22,N_9268,N_9002);
nand UO_23 (O_23,N_9230,N_9499);
nor UO_24 (O_24,N_9945,N_9781);
and UO_25 (O_25,N_9330,N_9209);
nor UO_26 (O_26,N_9735,N_9188);
or UO_27 (O_27,N_9922,N_9347);
or UO_28 (O_28,N_9071,N_9897);
nand UO_29 (O_29,N_9256,N_9470);
and UO_30 (O_30,N_9590,N_9106);
nand UO_31 (O_31,N_9562,N_9970);
xor UO_32 (O_32,N_9369,N_9316);
nand UO_33 (O_33,N_9249,N_9741);
nor UO_34 (O_34,N_9361,N_9183);
and UO_35 (O_35,N_9376,N_9246);
and UO_36 (O_36,N_9166,N_9677);
xnor UO_37 (O_37,N_9228,N_9890);
and UO_38 (O_38,N_9313,N_9588);
and UO_39 (O_39,N_9651,N_9295);
nand UO_40 (O_40,N_9434,N_9211);
or UO_41 (O_41,N_9331,N_9048);
and UO_42 (O_42,N_9736,N_9550);
nand UO_43 (O_43,N_9130,N_9513);
and UO_44 (O_44,N_9877,N_9296);
or UO_45 (O_45,N_9447,N_9275);
nand UO_46 (O_46,N_9969,N_9335);
nor UO_47 (O_47,N_9639,N_9602);
or UO_48 (O_48,N_9097,N_9044);
xor UO_49 (O_49,N_9751,N_9925);
or UO_50 (O_50,N_9072,N_9503);
nor UO_51 (O_51,N_9611,N_9524);
and UO_52 (O_52,N_9795,N_9554);
and UO_53 (O_53,N_9600,N_9757);
and UO_54 (O_54,N_9032,N_9703);
and UO_55 (O_55,N_9446,N_9116);
or UO_56 (O_56,N_9258,N_9941);
and UO_57 (O_57,N_9973,N_9310);
nand UO_58 (O_58,N_9494,N_9760);
and UO_59 (O_59,N_9966,N_9225);
and UO_60 (O_60,N_9041,N_9900);
nor UO_61 (O_61,N_9278,N_9823);
nand UO_62 (O_62,N_9064,N_9529);
or UO_63 (O_63,N_9687,N_9901);
nand UO_64 (O_64,N_9341,N_9774);
nor UO_65 (O_65,N_9806,N_9797);
or UO_66 (O_66,N_9199,N_9972);
and UO_67 (O_67,N_9034,N_9592);
or UO_68 (O_68,N_9998,N_9536);
and UO_69 (O_69,N_9979,N_9108);
nand UO_70 (O_70,N_9383,N_9396);
and UO_71 (O_71,N_9530,N_9915);
or UO_72 (O_72,N_9248,N_9899);
nand UO_73 (O_73,N_9923,N_9788);
nor UO_74 (O_74,N_9582,N_9525);
or UO_75 (O_75,N_9663,N_9716);
and UO_76 (O_76,N_9488,N_9872);
nor UO_77 (O_77,N_9682,N_9984);
nand UO_78 (O_78,N_9802,N_9187);
xor UO_79 (O_79,N_9668,N_9838);
nor UO_80 (O_80,N_9908,N_9830);
nand UO_81 (O_81,N_9237,N_9649);
and UO_82 (O_82,N_9832,N_9960);
nor UO_83 (O_83,N_9010,N_9539);
or UO_84 (O_84,N_9798,N_9579);
nor UO_85 (O_85,N_9410,N_9526);
nor UO_86 (O_86,N_9195,N_9424);
nand UO_87 (O_87,N_9443,N_9861);
or UO_88 (O_88,N_9866,N_9532);
and UO_89 (O_89,N_9087,N_9917);
nor UO_90 (O_90,N_9995,N_9303);
nand UO_91 (O_91,N_9342,N_9953);
or UO_92 (O_92,N_9412,N_9120);
nor UO_93 (O_93,N_9033,N_9796);
nand UO_94 (O_94,N_9365,N_9986);
or UO_95 (O_95,N_9546,N_9787);
and UO_96 (O_96,N_9596,N_9783);
and UO_97 (O_97,N_9150,N_9623);
and UO_98 (O_98,N_9180,N_9472);
or UO_99 (O_99,N_9836,N_9348);
or UO_100 (O_100,N_9684,N_9585);
nand UO_101 (O_101,N_9152,N_9723);
nor UO_102 (O_102,N_9438,N_9164);
nand UO_103 (O_103,N_9799,N_9119);
or UO_104 (O_104,N_9645,N_9770);
or UO_105 (O_105,N_9436,N_9360);
or UO_106 (O_106,N_9052,N_9732);
or UO_107 (O_107,N_9133,N_9765);
and UO_108 (O_108,N_9358,N_9626);
nand UO_109 (O_109,N_9398,N_9194);
nand UO_110 (O_110,N_9015,N_9715);
nor UO_111 (O_111,N_9767,N_9074);
or UO_112 (O_112,N_9614,N_9794);
nand UO_113 (O_113,N_9521,N_9320);
or UO_114 (O_114,N_9367,N_9101);
or UO_115 (O_115,N_9740,N_9580);
and UO_116 (O_116,N_9759,N_9835);
or UO_117 (O_117,N_9882,N_9117);
nand UO_118 (O_118,N_9886,N_9949);
nor UO_119 (O_119,N_9870,N_9563);
or UO_120 (O_120,N_9151,N_9982);
nand UO_121 (O_121,N_9111,N_9988);
nor UO_122 (O_122,N_9411,N_9846);
or UO_123 (O_123,N_9170,N_9233);
nor UO_124 (O_124,N_9753,N_9423);
xor UO_125 (O_125,N_9629,N_9744);
or UO_126 (O_126,N_9025,N_9699);
nand UO_127 (O_127,N_9676,N_9340);
and UO_128 (O_128,N_9871,N_9286);
and UO_129 (O_129,N_9589,N_9786);
or UO_130 (O_130,N_9161,N_9828);
nand UO_131 (O_131,N_9652,N_9069);
and UO_132 (O_132,N_9764,N_9189);
nor UO_133 (O_133,N_9378,N_9975);
xor UO_134 (O_134,N_9387,N_9062);
nand UO_135 (O_135,N_9670,N_9840);
nand UO_136 (O_136,N_9807,N_9815);
nor UO_137 (O_137,N_9245,N_9038);
or UO_138 (O_138,N_9281,N_9216);
and UO_139 (O_139,N_9952,N_9076);
and UO_140 (O_140,N_9421,N_9476);
and UO_141 (O_141,N_9292,N_9658);
nor UO_142 (O_142,N_9926,N_9191);
nand UO_143 (O_143,N_9479,N_9356);
and UO_144 (O_144,N_9154,N_9617);
nand UO_145 (O_145,N_9567,N_9635);
nand UO_146 (O_146,N_9553,N_9566);
nand UO_147 (O_147,N_9834,N_9747);
nand UO_148 (O_148,N_9305,N_9962);
and UO_149 (O_149,N_9214,N_9904);
and UO_150 (O_150,N_9463,N_9920);
or UO_151 (O_151,N_9441,N_9731);
or UO_152 (O_152,N_9583,N_9577);
and UO_153 (O_153,N_9790,N_9420);
nor UO_154 (O_154,N_9223,N_9094);
and UO_155 (O_155,N_9433,N_9024);
or UO_156 (O_156,N_9455,N_9819);
and UO_157 (O_157,N_9704,N_9486);
nor UO_158 (O_158,N_9028,N_9671);
or UO_159 (O_159,N_9375,N_9641);
nand UO_160 (O_160,N_9586,N_9750);
nand UO_161 (O_161,N_9132,N_9679);
or UO_162 (O_162,N_9919,N_9528);
nand UO_163 (O_163,N_9234,N_9714);
nand UO_164 (O_164,N_9318,N_9126);
nand UO_165 (O_165,N_9200,N_9182);
and UO_166 (O_166,N_9856,N_9535);
or UO_167 (O_167,N_9414,N_9067);
nor UO_168 (O_168,N_9801,N_9338);
nor UO_169 (O_169,N_9018,N_9314);
nor UO_170 (O_170,N_9707,N_9005);
nand UO_171 (O_171,N_9036,N_9311);
and UO_172 (O_172,N_9329,N_9843);
nand UO_173 (O_173,N_9053,N_9058);
or UO_174 (O_174,N_9950,N_9102);
and UO_175 (O_175,N_9162,N_9239);
and UO_176 (O_176,N_9581,N_9938);
or UO_177 (O_177,N_9839,N_9673);
xor UO_178 (O_178,N_9190,N_9604);
or UO_179 (O_179,N_9255,N_9854);
or UO_180 (O_180,N_9752,N_9619);
or UO_181 (O_181,N_9066,N_9302);
nor UO_182 (O_182,N_9357,N_9096);
nand UO_183 (O_183,N_9711,N_9388);
nand UO_184 (O_184,N_9855,N_9298);
or UO_185 (O_185,N_9304,N_9098);
nand UO_186 (O_186,N_9393,N_9265);
nand UO_187 (O_187,N_9867,N_9930);
nand UO_188 (O_188,N_9625,N_9203);
nand UO_189 (O_189,N_9370,N_9612);
and UO_190 (O_190,N_9215,N_9000);
nand UO_191 (O_191,N_9934,N_9533);
or UO_192 (O_192,N_9468,N_9879);
nand UO_193 (O_193,N_9779,N_9371);
or UO_194 (O_194,N_9510,N_9517);
nor UO_195 (O_195,N_9667,N_9889);
nand UO_196 (O_196,N_9805,N_9647);
nand UO_197 (O_197,N_9439,N_9850);
nor UO_198 (O_198,N_9409,N_9017);
nor UO_199 (O_199,N_9864,N_9413);
nand UO_200 (O_200,N_9056,N_9083);
nand UO_201 (O_201,N_9813,N_9353);
or UO_202 (O_202,N_9883,N_9457);
nor UO_203 (O_203,N_9822,N_9964);
or UO_204 (O_204,N_9777,N_9955);
and UO_205 (O_205,N_9860,N_9669);
nor UO_206 (O_206,N_9696,N_9896);
nand UO_207 (O_207,N_9148,N_9837);
or UO_208 (O_208,N_9933,N_9548);
and UO_209 (O_209,N_9432,N_9921);
nand UO_210 (O_210,N_9709,N_9205);
xor UO_211 (O_211,N_9755,N_9380);
or UO_212 (O_212,N_9491,N_9250);
or UO_213 (O_213,N_9299,N_9878);
and UO_214 (O_214,N_9327,N_9636);
nand UO_215 (O_215,N_9322,N_9713);
and UO_216 (O_216,N_9729,N_9487);
or UO_217 (O_217,N_9451,N_9814);
nand UO_218 (O_218,N_9880,N_9681);
nand UO_219 (O_219,N_9029,N_9541);
nand UO_220 (O_220,N_9492,N_9547);
and UO_221 (O_221,N_9165,N_9021);
and UO_222 (O_222,N_9294,N_9257);
or UO_223 (O_223,N_9936,N_9321);
or UO_224 (O_224,N_9570,N_9104);
nor UO_225 (O_225,N_9477,N_9538);
xnor UO_226 (O_226,N_9003,N_9168);
nor UO_227 (O_227,N_9721,N_9958);
nor UO_228 (O_228,N_9218,N_9907);
nand UO_229 (O_229,N_9031,N_9927);
and UO_230 (O_230,N_9394,N_9020);
or UO_231 (O_231,N_9448,N_9425);
nand UO_232 (O_232,N_9113,N_9282);
and UO_233 (O_233,N_9893,N_9089);
nor UO_234 (O_234,N_9050,N_9947);
or UO_235 (O_235,N_9607,N_9993);
or UO_236 (O_236,N_9201,N_9210);
nand UO_237 (O_237,N_9622,N_9105);
or UO_238 (O_238,N_9224,N_9591);
or UO_239 (O_239,N_9458,N_9504);
or UO_240 (O_240,N_9638,N_9829);
nand UO_241 (O_241,N_9288,N_9306);
and UO_242 (O_242,N_9100,N_9276);
nor UO_243 (O_243,N_9660,N_9266);
nand UO_244 (O_244,N_9372,N_9418);
and UO_245 (O_245,N_9742,N_9519);
and UO_246 (O_246,N_9171,N_9987);
and UO_247 (O_247,N_9875,N_9627);
nand UO_248 (O_248,N_9019,N_9963);
nand UO_249 (O_249,N_9202,N_9027);
nand UO_250 (O_250,N_9466,N_9279);
nor UO_251 (O_251,N_9138,N_9693);
nor UO_252 (O_252,N_9518,N_9666);
nor UO_253 (O_253,N_9431,N_9198);
and UO_254 (O_254,N_9219,N_9841);
nand UO_255 (O_255,N_9599,N_9459);
nand UO_256 (O_256,N_9131,N_9937);
nand UO_257 (O_257,N_9820,N_9842);
or UO_258 (O_258,N_9724,N_9047);
nor UO_259 (O_259,N_9733,N_9999);
nand UO_260 (O_260,N_9618,N_9939);
and UO_261 (O_261,N_9943,N_9483);
nand UO_262 (O_262,N_9037,N_9235);
or UO_263 (O_263,N_9985,N_9039);
or UO_264 (O_264,N_9107,N_9654);
nand UO_265 (O_265,N_9789,N_9243);
nor UO_266 (O_266,N_9968,N_9484);
and UO_267 (O_267,N_9873,N_9776);
nor UO_268 (O_268,N_9309,N_9368);
and UO_269 (O_269,N_9971,N_9754);
or UO_270 (O_270,N_9727,N_9804);
and UO_271 (O_271,N_9139,N_9332);
nor UO_272 (O_272,N_9502,N_9730);
or UO_273 (O_273,N_9137,N_9259);
or UO_274 (O_274,N_9469,N_9226);
and UO_275 (O_275,N_9159,N_9391);
nand UO_276 (O_276,N_9763,N_9859);
nand UO_277 (O_277,N_9605,N_9389);
nor UO_278 (O_278,N_9977,N_9826);
nand UO_279 (O_279,N_9642,N_9948);
nand UO_280 (O_280,N_9465,N_9012);
nand UO_281 (O_281,N_9323,N_9140);
nand UO_282 (O_282,N_9419,N_9613);
nor UO_283 (O_283,N_9646,N_9848);
and UO_284 (O_284,N_9086,N_9997);
and UO_285 (O_285,N_9147,N_9527);
nor UO_286 (O_286,N_9307,N_9743);
and UO_287 (O_287,N_9336,N_9127);
or UO_288 (O_288,N_9902,N_9242);
and UO_289 (O_289,N_9430,N_9109);
and UO_290 (O_290,N_9204,N_9339);
nor UO_291 (O_291,N_9768,N_9718);
nand UO_292 (O_292,N_9345,N_9495);
nor UO_293 (O_293,N_9792,N_9643);
and UO_294 (O_294,N_9762,N_9006);
and UO_295 (O_295,N_9260,N_9800);
or UO_296 (O_296,N_9088,N_9630);
or UO_297 (O_297,N_9672,N_9452);
or UO_298 (O_298,N_9270,N_9175);
nand UO_299 (O_299,N_9906,N_9009);
nand UO_300 (O_300,N_9051,N_9573);
or UO_301 (O_301,N_9057,N_9831);
or UO_302 (O_302,N_9445,N_9549);
nand UO_303 (O_303,N_9112,N_9269);
or UO_304 (O_304,N_9514,N_9888);
nand UO_305 (O_305,N_9910,N_9070);
or UO_306 (O_306,N_9640,N_9981);
nand UO_307 (O_307,N_9167,N_9594);
or UO_308 (O_308,N_9515,N_9179);
nand UO_309 (O_309,N_9475,N_9885);
and UO_310 (O_310,N_9373,N_9688);
and UO_311 (O_311,N_9808,N_9406);
nand UO_312 (O_312,N_9569,N_9771);
nand UO_313 (O_313,N_9887,N_9782);
nand UO_314 (O_314,N_9507,N_9157);
nor UO_315 (O_315,N_9697,N_9055);
nand UO_316 (O_316,N_9324,N_9467);
xor UO_317 (O_317,N_9217,N_9701);
nor UO_318 (O_318,N_9163,N_9891);
or UO_319 (O_319,N_9385,N_9444);
or UO_320 (O_320,N_9293,N_9632);
or UO_321 (O_321,N_9758,N_9746);
nor UO_322 (O_322,N_9608,N_9516);
or UO_323 (O_323,N_9174,N_9931);
or UO_324 (O_324,N_9912,N_9422);
nor UO_325 (O_325,N_9143,N_9653);
nand UO_326 (O_326,N_9450,N_9996);
and UO_327 (O_327,N_9262,N_9780);
nand UO_328 (O_328,N_9146,N_9990);
or UO_329 (O_329,N_9485,N_9994);
and UO_330 (O_330,N_9080,N_9075);
nor UO_331 (O_331,N_9099,N_9991);
nand UO_332 (O_332,N_9685,N_9942);
or UO_333 (O_333,N_9534,N_9719);
and UO_334 (O_334,N_9405,N_9091);
or UO_335 (O_335,N_9749,N_9903);
or UO_336 (O_336,N_9122,N_9349);
nand UO_337 (O_337,N_9916,N_9158);
and UO_338 (O_338,N_9196,N_9892);
nand UO_339 (O_339,N_9737,N_9197);
and UO_340 (O_340,N_9609,N_9905);
or UO_341 (O_341,N_9869,N_9557);
and UO_342 (O_342,N_9374,N_9844);
or UO_343 (O_343,N_9956,N_9054);
nor UO_344 (O_344,N_9169,N_9634);
nand UO_345 (O_345,N_9407,N_9913);
or UO_346 (O_346,N_9574,N_9090);
nand UO_347 (O_347,N_9390,N_9352);
and UO_348 (O_348,N_9176,N_9784);
nand UO_349 (O_349,N_9325,N_9650);
nand UO_350 (O_350,N_9959,N_9791);
and UO_351 (O_351,N_9144,N_9222);
nand UO_352 (O_352,N_9576,N_9428);
nor UO_353 (O_353,N_9346,N_9114);
or UO_354 (O_354,N_9403,N_9178);
nand UO_355 (O_355,N_9621,N_9016);
nand UO_356 (O_356,N_9384,N_9427);
or UO_357 (O_357,N_9496,N_9500);
or UO_358 (O_358,N_9290,N_9399);
nor UO_359 (O_359,N_9655,N_9285);
and UO_360 (O_360,N_9825,N_9935);
xnor UO_361 (O_361,N_9456,N_9748);
nor UO_362 (O_362,N_9659,N_9584);
nor UO_363 (O_363,N_9572,N_9772);
or UO_364 (O_364,N_9461,N_9142);
or UO_365 (O_365,N_9552,N_9277);
nor UO_366 (O_366,N_9350,N_9435);
nand UO_367 (O_367,N_9123,N_9155);
and UO_368 (O_368,N_9606,N_9847);
nor UO_369 (O_369,N_9283,N_9043);
and UO_370 (O_370,N_9725,N_9700);
nor UO_371 (O_371,N_9976,N_9961);
or UO_372 (O_372,N_9664,N_9620);
nor UO_373 (O_373,N_9355,N_9965);
nand UO_374 (O_374,N_9482,N_9408);
nor UO_375 (O_375,N_9710,N_9555);
nand UO_376 (O_376,N_9271,N_9134);
nand UO_377 (O_377,N_9631,N_9705);
and UO_378 (O_378,N_9125,N_9236);
or UO_379 (O_379,N_9252,N_9537);
nor UO_380 (O_380,N_9932,N_9675);
nor UO_381 (O_381,N_9739,N_9253);
nand UO_382 (O_382,N_9816,N_9284);
nor UO_383 (O_383,N_9480,N_9833);
or UO_384 (O_384,N_9035,N_9221);
and UO_385 (O_385,N_9181,N_9501);
and UO_386 (O_386,N_9312,N_9478);
nand UO_387 (O_387,N_9079,N_9454);
nand UO_388 (O_388,N_9545,N_9453);
nand UO_389 (O_389,N_9193,N_9065);
nor UO_390 (O_390,N_9229,N_9115);
nand UO_391 (O_391,N_9129,N_9192);
and UO_392 (O_392,N_9734,N_9402);
nand UO_393 (O_393,N_9437,N_9013);
and UO_394 (O_394,N_9212,N_9177);
nand UO_395 (O_395,N_9894,N_9030);
or UO_396 (O_396,N_9287,N_9238);
nor UO_397 (O_397,N_9722,N_9811);
nor UO_398 (O_398,N_9587,N_9980);
nand UO_399 (O_399,N_9674,N_9560);
and UO_400 (O_400,N_9881,N_9308);
and UO_401 (O_401,N_9462,N_9363);
or UO_402 (O_402,N_9863,N_9662);
or UO_403 (O_403,N_9706,N_9989);
or UO_404 (O_404,N_9978,N_9267);
nor UO_405 (O_405,N_9046,N_9232);
nand UO_406 (O_406,N_9231,N_9884);
nor UO_407 (O_407,N_9565,N_9173);
and UO_408 (O_408,N_9426,N_9481);
and UO_409 (O_409,N_9558,N_9084);
and UO_410 (O_410,N_9615,N_9624);
or UO_411 (O_411,N_9551,N_9610);
nor UO_412 (O_412,N_9992,N_9001);
and UO_413 (O_413,N_9556,N_9957);
and UO_414 (O_414,N_9400,N_9110);
and UO_415 (O_415,N_9121,N_9343);
and UO_416 (O_416,N_9206,N_9918);
and UO_417 (O_417,N_9379,N_9092);
or UO_418 (O_418,N_9506,N_9460);
and UO_419 (O_419,N_9124,N_9490);
or UO_420 (O_420,N_9665,N_9540);
nor UO_421 (O_421,N_9720,N_9289);
nor UO_422 (O_422,N_9061,N_9523);
nor UO_423 (O_423,N_9471,N_9601);
and UO_424 (O_424,N_9068,N_9683);
nor UO_425 (O_425,N_9698,N_9366);
nor UO_426 (O_426,N_9404,N_9082);
or UO_427 (O_427,N_9728,N_9049);
nor UO_428 (O_428,N_9011,N_9603);
or UO_429 (O_429,N_9186,N_9301);
nand UO_430 (O_430,N_9865,N_9690);
nand UO_431 (O_431,N_9007,N_9637);
nand UO_432 (O_432,N_9023,N_9543);
and UO_433 (O_433,N_9045,N_9440);
nand UO_434 (O_434,N_9273,N_9571);
nand UO_435 (O_435,N_9694,N_9326);
nor UO_436 (O_436,N_9172,N_9251);
nand UO_437 (O_437,N_9544,N_9849);
and UO_438 (O_438,N_9145,N_9185);
and UO_439 (O_439,N_9845,N_9773);
or UO_440 (O_440,N_9785,N_9712);
and UO_441 (O_441,N_9769,N_9416);
or UO_442 (O_442,N_9333,N_9775);
nor UO_443 (O_443,N_9464,N_9598);
nand UO_444 (O_444,N_9940,N_9876);
and UO_445 (O_445,N_9678,N_9395);
or UO_446 (O_446,N_9272,N_9240);
and UO_447 (O_447,N_9661,N_9059);
nand UO_448 (O_448,N_9756,N_9895);
or UO_449 (O_449,N_9909,N_9263);
nand UO_450 (O_450,N_9208,N_9081);
nand UO_451 (O_451,N_9512,N_9442);
or UO_452 (O_452,N_9085,N_9103);
or UO_453 (O_453,N_9531,N_9929);
and UO_454 (O_454,N_9578,N_9351);
nand UO_455 (O_455,N_9274,N_9633);
nand UO_456 (O_456,N_9559,N_9136);
nor UO_457 (O_457,N_9004,N_9498);
nand UO_458 (O_458,N_9924,N_9874);
nand UO_459 (O_459,N_9315,N_9297);
and UO_460 (O_460,N_9014,N_9280);
nand UO_461 (O_461,N_9317,N_9497);
nand UO_462 (O_462,N_9708,N_9686);
or UO_463 (O_463,N_9689,N_9818);
and UO_464 (O_464,N_9247,N_9745);
and UO_465 (O_465,N_9928,N_9149);
nand UO_466 (O_466,N_9738,N_9153);
and UO_467 (O_467,N_9244,N_9561);
xnor UO_468 (O_468,N_9220,N_9821);
nor UO_469 (O_469,N_9344,N_9616);
nor UO_470 (O_470,N_9695,N_9595);
nand UO_471 (O_471,N_9429,N_9946);
nor UO_472 (O_472,N_9401,N_9493);
nand UO_473 (O_473,N_9803,N_9520);
or UO_474 (O_474,N_9319,N_9898);
or UO_475 (O_475,N_9241,N_9261);
nand UO_476 (O_476,N_9568,N_9254);
nor UO_477 (O_477,N_9073,N_9974);
and UO_478 (O_478,N_9093,N_9135);
and UO_479 (O_479,N_9077,N_9377);
or UO_480 (O_480,N_9141,N_9868);
nand UO_481 (O_481,N_9817,N_9040);
and UO_482 (O_482,N_9522,N_9160);
and UO_483 (O_483,N_9951,N_9793);
nor UO_484 (O_484,N_9386,N_9944);
nor UO_485 (O_485,N_9078,N_9851);
nor UO_486 (O_486,N_9227,N_9359);
or UO_487 (O_487,N_9095,N_9911);
nand UO_488 (O_488,N_9778,N_9026);
nor UO_489 (O_489,N_9060,N_9128);
nand UO_490 (O_490,N_9761,N_9852);
nand UO_491 (O_491,N_9593,N_9300);
nor UO_492 (O_492,N_9417,N_9291);
nor UO_493 (O_493,N_9597,N_9967);
and UO_494 (O_494,N_9184,N_9717);
nand UO_495 (O_495,N_9575,N_9264);
xor UO_496 (O_496,N_9511,N_9914);
nor UO_497 (O_497,N_9680,N_9824);
and UO_498 (O_498,N_9042,N_9118);
nand UO_499 (O_499,N_9364,N_9213);
and UO_500 (O_500,N_9403,N_9231);
or UO_501 (O_501,N_9587,N_9554);
and UO_502 (O_502,N_9985,N_9566);
or UO_503 (O_503,N_9274,N_9472);
nor UO_504 (O_504,N_9201,N_9608);
nor UO_505 (O_505,N_9630,N_9412);
nor UO_506 (O_506,N_9294,N_9593);
nand UO_507 (O_507,N_9146,N_9594);
nand UO_508 (O_508,N_9567,N_9017);
or UO_509 (O_509,N_9718,N_9947);
or UO_510 (O_510,N_9844,N_9636);
nand UO_511 (O_511,N_9154,N_9608);
or UO_512 (O_512,N_9838,N_9624);
nor UO_513 (O_513,N_9412,N_9638);
or UO_514 (O_514,N_9830,N_9094);
nor UO_515 (O_515,N_9553,N_9238);
and UO_516 (O_516,N_9876,N_9974);
nor UO_517 (O_517,N_9192,N_9711);
nor UO_518 (O_518,N_9458,N_9926);
nor UO_519 (O_519,N_9234,N_9273);
nand UO_520 (O_520,N_9114,N_9359);
nand UO_521 (O_521,N_9302,N_9166);
nand UO_522 (O_522,N_9612,N_9253);
nand UO_523 (O_523,N_9337,N_9029);
nor UO_524 (O_524,N_9459,N_9048);
or UO_525 (O_525,N_9962,N_9469);
nor UO_526 (O_526,N_9398,N_9464);
or UO_527 (O_527,N_9316,N_9144);
or UO_528 (O_528,N_9275,N_9515);
or UO_529 (O_529,N_9362,N_9154);
and UO_530 (O_530,N_9571,N_9880);
and UO_531 (O_531,N_9837,N_9063);
and UO_532 (O_532,N_9685,N_9668);
nor UO_533 (O_533,N_9363,N_9004);
and UO_534 (O_534,N_9452,N_9020);
nand UO_535 (O_535,N_9471,N_9492);
and UO_536 (O_536,N_9589,N_9046);
and UO_537 (O_537,N_9295,N_9301);
or UO_538 (O_538,N_9412,N_9040);
and UO_539 (O_539,N_9398,N_9158);
nand UO_540 (O_540,N_9313,N_9532);
or UO_541 (O_541,N_9299,N_9410);
nand UO_542 (O_542,N_9168,N_9490);
nor UO_543 (O_543,N_9329,N_9704);
and UO_544 (O_544,N_9281,N_9547);
or UO_545 (O_545,N_9400,N_9237);
or UO_546 (O_546,N_9208,N_9335);
and UO_547 (O_547,N_9783,N_9806);
and UO_548 (O_548,N_9891,N_9741);
and UO_549 (O_549,N_9615,N_9942);
nor UO_550 (O_550,N_9069,N_9159);
and UO_551 (O_551,N_9903,N_9376);
nand UO_552 (O_552,N_9365,N_9294);
nor UO_553 (O_553,N_9935,N_9735);
or UO_554 (O_554,N_9330,N_9178);
nand UO_555 (O_555,N_9507,N_9009);
nor UO_556 (O_556,N_9733,N_9960);
and UO_557 (O_557,N_9114,N_9072);
and UO_558 (O_558,N_9767,N_9190);
nor UO_559 (O_559,N_9675,N_9293);
nor UO_560 (O_560,N_9994,N_9047);
and UO_561 (O_561,N_9097,N_9493);
or UO_562 (O_562,N_9706,N_9713);
and UO_563 (O_563,N_9317,N_9650);
nand UO_564 (O_564,N_9017,N_9822);
nand UO_565 (O_565,N_9016,N_9428);
and UO_566 (O_566,N_9413,N_9565);
and UO_567 (O_567,N_9846,N_9960);
nand UO_568 (O_568,N_9583,N_9326);
nor UO_569 (O_569,N_9565,N_9593);
or UO_570 (O_570,N_9433,N_9079);
or UO_571 (O_571,N_9759,N_9853);
nor UO_572 (O_572,N_9133,N_9684);
or UO_573 (O_573,N_9233,N_9020);
nor UO_574 (O_574,N_9347,N_9675);
nand UO_575 (O_575,N_9018,N_9507);
nand UO_576 (O_576,N_9410,N_9252);
nor UO_577 (O_577,N_9838,N_9260);
or UO_578 (O_578,N_9275,N_9880);
nand UO_579 (O_579,N_9194,N_9084);
nor UO_580 (O_580,N_9668,N_9625);
and UO_581 (O_581,N_9881,N_9494);
nor UO_582 (O_582,N_9512,N_9168);
nand UO_583 (O_583,N_9375,N_9670);
nor UO_584 (O_584,N_9539,N_9933);
nor UO_585 (O_585,N_9434,N_9619);
nor UO_586 (O_586,N_9767,N_9598);
nand UO_587 (O_587,N_9863,N_9693);
and UO_588 (O_588,N_9128,N_9515);
or UO_589 (O_589,N_9828,N_9368);
nor UO_590 (O_590,N_9293,N_9394);
and UO_591 (O_591,N_9532,N_9729);
nand UO_592 (O_592,N_9518,N_9221);
nor UO_593 (O_593,N_9763,N_9657);
and UO_594 (O_594,N_9980,N_9765);
or UO_595 (O_595,N_9512,N_9982);
or UO_596 (O_596,N_9445,N_9588);
or UO_597 (O_597,N_9954,N_9285);
and UO_598 (O_598,N_9337,N_9213);
and UO_599 (O_599,N_9539,N_9908);
and UO_600 (O_600,N_9915,N_9025);
nor UO_601 (O_601,N_9530,N_9242);
nor UO_602 (O_602,N_9635,N_9100);
nor UO_603 (O_603,N_9217,N_9136);
and UO_604 (O_604,N_9977,N_9757);
nand UO_605 (O_605,N_9471,N_9530);
nor UO_606 (O_606,N_9226,N_9434);
nand UO_607 (O_607,N_9915,N_9004);
or UO_608 (O_608,N_9424,N_9372);
nand UO_609 (O_609,N_9943,N_9477);
or UO_610 (O_610,N_9531,N_9941);
nand UO_611 (O_611,N_9067,N_9535);
nand UO_612 (O_612,N_9042,N_9753);
nand UO_613 (O_613,N_9859,N_9878);
and UO_614 (O_614,N_9111,N_9937);
nand UO_615 (O_615,N_9816,N_9203);
and UO_616 (O_616,N_9789,N_9930);
and UO_617 (O_617,N_9364,N_9882);
or UO_618 (O_618,N_9313,N_9884);
and UO_619 (O_619,N_9562,N_9327);
or UO_620 (O_620,N_9243,N_9549);
nand UO_621 (O_621,N_9069,N_9125);
or UO_622 (O_622,N_9572,N_9827);
nor UO_623 (O_623,N_9515,N_9493);
nor UO_624 (O_624,N_9973,N_9052);
nor UO_625 (O_625,N_9337,N_9730);
and UO_626 (O_626,N_9502,N_9330);
nand UO_627 (O_627,N_9130,N_9073);
nand UO_628 (O_628,N_9254,N_9984);
nand UO_629 (O_629,N_9970,N_9855);
or UO_630 (O_630,N_9524,N_9811);
nor UO_631 (O_631,N_9283,N_9892);
nand UO_632 (O_632,N_9722,N_9417);
nor UO_633 (O_633,N_9126,N_9561);
or UO_634 (O_634,N_9750,N_9319);
nor UO_635 (O_635,N_9504,N_9723);
nand UO_636 (O_636,N_9665,N_9800);
nand UO_637 (O_637,N_9559,N_9519);
and UO_638 (O_638,N_9713,N_9746);
and UO_639 (O_639,N_9455,N_9744);
nor UO_640 (O_640,N_9148,N_9325);
or UO_641 (O_641,N_9690,N_9095);
nand UO_642 (O_642,N_9163,N_9068);
and UO_643 (O_643,N_9009,N_9054);
or UO_644 (O_644,N_9201,N_9699);
or UO_645 (O_645,N_9928,N_9355);
nand UO_646 (O_646,N_9305,N_9640);
nor UO_647 (O_647,N_9538,N_9539);
nand UO_648 (O_648,N_9530,N_9628);
nor UO_649 (O_649,N_9212,N_9716);
nor UO_650 (O_650,N_9867,N_9430);
or UO_651 (O_651,N_9210,N_9556);
nor UO_652 (O_652,N_9843,N_9250);
or UO_653 (O_653,N_9656,N_9968);
and UO_654 (O_654,N_9738,N_9604);
nor UO_655 (O_655,N_9831,N_9061);
nor UO_656 (O_656,N_9935,N_9062);
nand UO_657 (O_657,N_9570,N_9074);
nand UO_658 (O_658,N_9668,N_9472);
nor UO_659 (O_659,N_9457,N_9509);
nor UO_660 (O_660,N_9023,N_9050);
nor UO_661 (O_661,N_9044,N_9972);
nor UO_662 (O_662,N_9915,N_9408);
or UO_663 (O_663,N_9085,N_9087);
nor UO_664 (O_664,N_9075,N_9628);
nor UO_665 (O_665,N_9197,N_9037);
and UO_666 (O_666,N_9821,N_9829);
and UO_667 (O_667,N_9664,N_9769);
nand UO_668 (O_668,N_9801,N_9888);
and UO_669 (O_669,N_9412,N_9440);
and UO_670 (O_670,N_9695,N_9057);
and UO_671 (O_671,N_9164,N_9524);
nand UO_672 (O_672,N_9184,N_9468);
or UO_673 (O_673,N_9082,N_9217);
nand UO_674 (O_674,N_9418,N_9545);
or UO_675 (O_675,N_9070,N_9022);
nand UO_676 (O_676,N_9090,N_9668);
nand UO_677 (O_677,N_9150,N_9461);
or UO_678 (O_678,N_9760,N_9519);
nand UO_679 (O_679,N_9020,N_9848);
nand UO_680 (O_680,N_9798,N_9611);
nand UO_681 (O_681,N_9067,N_9703);
nand UO_682 (O_682,N_9353,N_9836);
or UO_683 (O_683,N_9292,N_9581);
or UO_684 (O_684,N_9489,N_9790);
or UO_685 (O_685,N_9077,N_9149);
or UO_686 (O_686,N_9958,N_9513);
nor UO_687 (O_687,N_9403,N_9673);
or UO_688 (O_688,N_9820,N_9831);
nand UO_689 (O_689,N_9741,N_9819);
nand UO_690 (O_690,N_9852,N_9876);
and UO_691 (O_691,N_9190,N_9173);
nor UO_692 (O_692,N_9884,N_9304);
nor UO_693 (O_693,N_9300,N_9068);
nand UO_694 (O_694,N_9576,N_9619);
and UO_695 (O_695,N_9159,N_9584);
and UO_696 (O_696,N_9896,N_9500);
nor UO_697 (O_697,N_9533,N_9161);
nand UO_698 (O_698,N_9695,N_9860);
and UO_699 (O_699,N_9367,N_9018);
nor UO_700 (O_700,N_9879,N_9202);
nor UO_701 (O_701,N_9709,N_9264);
and UO_702 (O_702,N_9534,N_9112);
nor UO_703 (O_703,N_9273,N_9514);
nand UO_704 (O_704,N_9397,N_9641);
nor UO_705 (O_705,N_9008,N_9105);
and UO_706 (O_706,N_9009,N_9393);
nand UO_707 (O_707,N_9890,N_9896);
and UO_708 (O_708,N_9392,N_9966);
and UO_709 (O_709,N_9307,N_9480);
nand UO_710 (O_710,N_9705,N_9696);
nand UO_711 (O_711,N_9246,N_9596);
nor UO_712 (O_712,N_9705,N_9737);
nand UO_713 (O_713,N_9580,N_9896);
nand UO_714 (O_714,N_9320,N_9646);
and UO_715 (O_715,N_9717,N_9779);
or UO_716 (O_716,N_9569,N_9380);
nand UO_717 (O_717,N_9488,N_9657);
or UO_718 (O_718,N_9744,N_9223);
and UO_719 (O_719,N_9105,N_9563);
nor UO_720 (O_720,N_9492,N_9909);
and UO_721 (O_721,N_9929,N_9818);
or UO_722 (O_722,N_9843,N_9454);
and UO_723 (O_723,N_9283,N_9538);
and UO_724 (O_724,N_9562,N_9382);
nand UO_725 (O_725,N_9519,N_9228);
nand UO_726 (O_726,N_9456,N_9481);
nand UO_727 (O_727,N_9423,N_9928);
or UO_728 (O_728,N_9138,N_9739);
nor UO_729 (O_729,N_9405,N_9675);
nor UO_730 (O_730,N_9562,N_9683);
nand UO_731 (O_731,N_9279,N_9594);
nand UO_732 (O_732,N_9926,N_9899);
or UO_733 (O_733,N_9503,N_9767);
nor UO_734 (O_734,N_9984,N_9802);
and UO_735 (O_735,N_9711,N_9112);
or UO_736 (O_736,N_9876,N_9127);
nand UO_737 (O_737,N_9039,N_9160);
and UO_738 (O_738,N_9003,N_9432);
or UO_739 (O_739,N_9724,N_9556);
nand UO_740 (O_740,N_9791,N_9018);
or UO_741 (O_741,N_9908,N_9017);
nor UO_742 (O_742,N_9003,N_9597);
or UO_743 (O_743,N_9611,N_9769);
nand UO_744 (O_744,N_9495,N_9202);
or UO_745 (O_745,N_9362,N_9634);
or UO_746 (O_746,N_9565,N_9427);
nand UO_747 (O_747,N_9718,N_9262);
or UO_748 (O_748,N_9506,N_9992);
nor UO_749 (O_749,N_9996,N_9623);
nand UO_750 (O_750,N_9552,N_9618);
nand UO_751 (O_751,N_9352,N_9406);
and UO_752 (O_752,N_9737,N_9527);
nand UO_753 (O_753,N_9142,N_9044);
and UO_754 (O_754,N_9693,N_9244);
nor UO_755 (O_755,N_9715,N_9373);
and UO_756 (O_756,N_9968,N_9606);
or UO_757 (O_757,N_9064,N_9649);
and UO_758 (O_758,N_9763,N_9921);
nor UO_759 (O_759,N_9637,N_9591);
and UO_760 (O_760,N_9949,N_9285);
or UO_761 (O_761,N_9003,N_9408);
and UO_762 (O_762,N_9464,N_9533);
xor UO_763 (O_763,N_9126,N_9798);
nor UO_764 (O_764,N_9044,N_9754);
nor UO_765 (O_765,N_9679,N_9448);
and UO_766 (O_766,N_9586,N_9889);
or UO_767 (O_767,N_9858,N_9095);
or UO_768 (O_768,N_9133,N_9720);
nor UO_769 (O_769,N_9160,N_9218);
nor UO_770 (O_770,N_9528,N_9757);
or UO_771 (O_771,N_9233,N_9534);
nand UO_772 (O_772,N_9741,N_9386);
or UO_773 (O_773,N_9025,N_9981);
nand UO_774 (O_774,N_9893,N_9990);
nand UO_775 (O_775,N_9730,N_9614);
or UO_776 (O_776,N_9158,N_9081);
or UO_777 (O_777,N_9450,N_9580);
nor UO_778 (O_778,N_9277,N_9666);
or UO_779 (O_779,N_9126,N_9034);
nor UO_780 (O_780,N_9855,N_9463);
nor UO_781 (O_781,N_9328,N_9566);
nand UO_782 (O_782,N_9177,N_9454);
and UO_783 (O_783,N_9569,N_9219);
or UO_784 (O_784,N_9219,N_9344);
or UO_785 (O_785,N_9781,N_9668);
and UO_786 (O_786,N_9824,N_9416);
xnor UO_787 (O_787,N_9296,N_9817);
nor UO_788 (O_788,N_9424,N_9203);
or UO_789 (O_789,N_9254,N_9630);
and UO_790 (O_790,N_9036,N_9456);
and UO_791 (O_791,N_9111,N_9942);
or UO_792 (O_792,N_9287,N_9672);
and UO_793 (O_793,N_9153,N_9286);
and UO_794 (O_794,N_9450,N_9164);
nor UO_795 (O_795,N_9923,N_9189);
and UO_796 (O_796,N_9768,N_9205);
nand UO_797 (O_797,N_9107,N_9628);
and UO_798 (O_798,N_9043,N_9629);
and UO_799 (O_799,N_9237,N_9808);
and UO_800 (O_800,N_9633,N_9970);
nor UO_801 (O_801,N_9654,N_9866);
or UO_802 (O_802,N_9612,N_9044);
or UO_803 (O_803,N_9311,N_9187);
nor UO_804 (O_804,N_9225,N_9929);
nor UO_805 (O_805,N_9475,N_9650);
nand UO_806 (O_806,N_9027,N_9174);
or UO_807 (O_807,N_9478,N_9573);
or UO_808 (O_808,N_9743,N_9111);
and UO_809 (O_809,N_9308,N_9653);
or UO_810 (O_810,N_9817,N_9796);
nand UO_811 (O_811,N_9484,N_9545);
or UO_812 (O_812,N_9774,N_9984);
and UO_813 (O_813,N_9680,N_9973);
and UO_814 (O_814,N_9297,N_9681);
and UO_815 (O_815,N_9303,N_9759);
nor UO_816 (O_816,N_9371,N_9873);
and UO_817 (O_817,N_9392,N_9329);
or UO_818 (O_818,N_9812,N_9595);
and UO_819 (O_819,N_9672,N_9792);
or UO_820 (O_820,N_9512,N_9908);
nand UO_821 (O_821,N_9067,N_9784);
or UO_822 (O_822,N_9007,N_9253);
and UO_823 (O_823,N_9060,N_9172);
or UO_824 (O_824,N_9934,N_9948);
nand UO_825 (O_825,N_9646,N_9737);
nor UO_826 (O_826,N_9909,N_9800);
or UO_827 (O_827,N_9527,N_9655);
or UO_828 (O_828,N_9922,N_9652);
or UO_829 (O_829,N_9304,N_9391);
nand UO_830 (O_830,N_9155,N_9620);
nor UO_831 (O_831,N_9221,N_9781);
nand UO_832 (O_832,N_9969,N_9984);
nand UO_833 (O_833,N_9192,N_9911);
nor UO_834 (O_834,N_9428,N_9045);
and UO_835 (O_835,N_9712,N_9355);
and UO_836 (O_836,N_9203,N_9018);
nand UO_837 (O_837,N_9315,N_9163);
nand UO_838 (O_838,N_9797,N_9717);
and UO_839 (O_839,N_9118,N_9160);
or UO_840 (O_840,N_9341,N_9929);
or UO_841 (O_841,N_9012,N_9121);
or UO_842 (O_842,N_9052,N_9508);
nand UO_843 (O_843,N_9424,N_9111);
or UO_844 (O_844,N_9531,N_9293);
nand UO_845 (O_845,N_9164,N_9559);
nand UO_846 (O_846,N_9470,N_9513);
and UO_847 (O_847,N_9583,N_9419);
and UO_848 (O_848,N_9814,N_9323);
nand UO_849 (O_849,N_9425,N_9733);
and UO_850 (O_850,N_9224,N_9838);
nor UO_851 (O_851,N_9334,N_9192);
nor UO_852 (O_852,N_9641,N_9245);
or UO_853 (O_853,N_9815,N_9906);
and UO_854 (O_854,N_9750,N_9561);
xnor UO_855 (O_855,N_9777,N_9140);
xnor UO_856 (O_856,N_9209,N_9543);
nor UO_857 (O_857,N_9426,N_9038);
nor UO_858 (O_858,N_9532,N_9098);
or UO_859 (O_859,N_9411,N_9171);
nor UO_860 (O_860,N_9880,N_9762);
or UO_861 (O_861,N_9552,N_9508);
and UO_862 (O_862,N_9057,N_9275);
and UO_863 (O_863,N_9876,N_9628);
or UO_864 (O_864,N_9865,N_9229);
or UO_865 (O_865,N_9435,N_9571);
nor UO_866 (O_866,N_9404,N_9549);
nor UO_867 (O_867,N_9499,N_9027);
xor UO_868 (O_868,N_9486,N_9975);
and UO_869 (O_869,N_9897,N_9456);
and UO_870 (O_870,N_9315,N_9752);
and UO_871 (O_871,N_9684,N_9141);
and UO_872 (O_872,N_9034,N_9540);
nor UO_873 (O_873,N_9017,N_9819);
or UO_874 (O_874,N_9379,N_9581);
and UO_875 (O_875,N_9632,N_9451);
and UO_876 (O_876,N_9804,N_9354);
nor UO_877 (O_877,N_9918,N_9323);
nor UO_878 (O_878,N_9510,N_9779);
or UO_879 (O_879,N_9137,N_9948);
and UO_880 (O_880,N_9622,N_9298);
nand UO_881 (O_881,N_9426,N_9064);
and UO_882 (O_882,N_9608,N_9943);
nand UO_883 (O_883,N_9084,N_9745);
nor UO_884 (O_884,N_9268,N_9384);
nand UO_885 (O_885,N_9966,N_9121);
and UO_886 (O_886,N_9868,N_9630);
nor UO_887 (O_887,N_9259,N_9970);
or UO_888 (O_888,N_9120,N_9243);
or UO_889 (O_889,N_9273,N_9417);
and UO_890 (O_890,N_9263,N_9601);
nor UO_891 (O_891,N_9252,N_9020);
and UO_892 (O_892,N_9436,N_9738);
nand UO_893 (O_893,N_9714,N_9048);
and UO_894 (O_894,N_9549,N_9833);
or UO_895 (O_895,N_9546,N_9342);
and UO_896 (O_896,N_9523,N_9126);
nor UO_897 (O_897,N_9310,N_9989);
nand UO_898 (O_898,N_9518,N_9584);
nor UO_899 (O_899,N_9371,N_9069);
or UO_900 (O_900,N_9784,N_9320);
nor UO_901 (O_901,N_9954,N_9600);
and UO_902 (O_902,N_9199,N_9341);
nand UO_903 (O_903,N_9358,N_9950);
or UO_904 (O_904,N_9707,N_9930);
nor UO_905 (O_905,N_9607,N_9191);
and UO_906 (O_906,N_9130,N_9286);
or UO_907 (O_907,N_9687,N_9229);
and UO_908 (O_908,N_9256,N_9036);
nor UO_909 (O_909,N_9501,N_9844);
or UO_910 (O_910,N_9309,N_9740);
and UO_911 (O_911,N_9790,N_9802);
or UO_912 (O_912,N_9608,N_9115);
nor UO_913 (O_913,N_9975,N_9464);
and UO_914 (O_914,N_9407,N_9001);
and UO_915 (O_915,N_9077,N_9008);
nand UO_916 (O_916,N_9968,N_9228);
nand UO_917 (O_917,N_9817,N_9614);
nor UO_918 (O_918,N_9654,N_9152);
and UO_919 (O_919,N_9687,N_9363);
and UO_920 (O_920,N_9826,N_9118);
or UO_921 (O_921,N_9936,N_9719);
or UO_922 (O_922,N_9467,N_9284);
nand UO_923 (O_923,N_9079,N_9030);
and UO_924 (O_924,N_9291,N_9942);
or UO_925 (O_925,N_9940,N_9000);
nor UO_926 (O_926,N_9996,N_9918);
nor UO_927 (O_927,N_9568,N_9737);
or UO_928 (O_928,N_9652,N_9353);
nor UO_929 (O_929,N_9655,N_9691);
nor UO_930 (O_930,N_9030,N_9389);
nor UO_931 (O_931,N_9434,N_9658);
or UO_932 (O_932,N_9703,N_9711);
nand UO_933 (O_933,N_9551,N_9029);
or UO_934 (O_934,N_9445,N_9382);
or UO_935 (O_935,N_9273,N_9856);
and UO_936 (O_936,N_9689,N_9432);
nand UO_937 (O_937,N_9707,N_9612);
nand UO_938 (O_938,N_9072,N_9852);
and UO_939 (O_939,N_9091,N_9057);
nor UO_940 (O_940,N_9140,N_9241);
or UO_941 (O_941,N_9353,N_9972);
nor UO_942 (O_942,N_9307,N_9917);
nand UO_943 (O_943,N_9713,N_9309);
nor UO_944 (O_944,N_9755,N_9413);
nor UO_945 (O_945,N_9941,N_9928);
nand UO_946 (O_946,N_9147,N_9226);
nor UO_947 (O_947,N_9213,N_9740);
and UO_948 (O_948,N_9139,N_9838);
nor UO_949 (O_949,N_9728,N_9592);
nor UO_950 (O_950,N_9494,N_9584);
and UO_951 (O_951,N_9127,N_9166);
nand UO_952 (O_952,N_9249,N_9457);
or UO_953 (O_953,N_9102,N_9808);
and UO_954 (O_954,N_9996,N_9862);
and UO_955 (O_955,N_9984,N_9291);
nor UO_956 (O_956,N_9802,N_9576);
nand UO_957 (O_957,N_9026,N_9775);
and UO_958 (O_958,N_9040,N_9055);
or UO_959 (O_959,N_9477,N_9510);
nand UO_960 (O_960,N_9410,N_9936);
nor UO_961 (O_961,N_9661,N_9048);
nor UO_962 (O_962,N_9061,N_9819);
and UO_963 (O_963,N_9013,N_9206);
nor UO_964 (O_964,N_9483,N_9116);
nand UO_965 (O_965,N_9016,N_9276);
nand UO_966 (O_966,N_9492,N_9175);
nand UO_967 (O_967,N_9964,N_9038);
and UO_968 (O_968,N_9527,N_9691);
or UO_969 (O_969,N_9206,N_9248);
nand UO_970 (O_970,N_9699,N_9802);
nor UO_971 (O_971,N_9176,N_9042);
nor UO_972 (O_972,N_9828,N_9962);
and UO_973 (O_973,N_9000,N_9503);
nand UO_974 (O_974,N_9256,N_9096);
or UO_975 (O_975,N_9674,N_9324);
nor UO_976 (O_976,N_9267,N_9611);
and UO_977 (O_977,N_9308,N_9247);
and UO_978 (O_978,N_9335,N_9980);
nand UO_979 (O_979,N_9513,N_9053);
nand UO_980 (O_980,N_9309,N_9006);
xnor UO_981 (O_981,N_9985,N_9932);
or UO_982 (O_982,N_9339,N_9095);
nand UO_983 (O_983,N_9132,N_9996);
xnor UO_984 (O_984,N_9556,N_9783);
and UO_985 (O_985,N_9265,N_9457);
and UO_986 (O_986,N_9522,N_9290);
and UO_987 (O_987,N_9582,N_9336);
nand UO_988 (O_988,N_9506,N_9599);
nand UO_989 (O_989,N_9173,N_9814);
nand UO_990 (O_990,N_9810,N_9661);
or UO_991 (O_991,N_9866,N_9786);
and UO_992 (O_992,N_9967,N_9169);
nand UO_993 (O_993,N_9257,N_9189);
and UO_994 (O_994,N_9332,N_9673);
nor UO_995 (O_995,N_9471,N_9404);
or UO_996 (O_996,N_9349,N_9213);
and UO_997 (O_997,N_9528,N_9327);
nand UO_998 (O_998,N_9765,N_9708);
nand UO_999 (O_999,N_9186,N_9507);
and UO_1000 (O_1000,N_9532,N_9127);
nand UO_1001 (O_1001,N_9157,N_9280);
nand UO_1002 (O_1002,N_9733,N_9512);
or UO_1003 (O_1003,N_9125,N_9752);
or UO_1004 (O_1004,N_9187,N_9509);
nand UO_1005 (O_1005,N_9753,N_9626);
nand UO_1006 (O_1006,N_9598,N_9735);
nor UO_1007 (O_1007,N_9903,N_9648);
nor UO_1008 (O_1008,N_9551,N_9513);
and UO_1009 (O_1009,N_9024,N_9288);
nor UO_1010 (O_1010,N_9133,N_9995);
nand UO_1011 (O_1011,N_9996,N_9897);
and UO_1012 (O_1012,N_9192,N_9228);
xor UO_1013 (O_1013,N_9198,N_9844);
or UO_1014 (O_1014,N_9690,N_9755);
nor UO_1015 (O_1015,N_9581,N_9214);
nand UO_1016 (O_1016,N_9357,N_9634);
or UO_1017 (O_1017,N_9667,N_9718);
or UO_1018 (O_1018,N_9047,N_9074);
and UO_1019 (O_1019,N_9697,N_9054);
nand UO_1020 (O_1020,N_9047,N_9045);
and UO_1021 (O_1021,N_9223,N_9463);
and UO_1022 (O_1022,N_9277,N_9534);
nand UO_1023 (O_1023,N_9118,N_9139);
and UO_1024 (O_1024,N_9672,N_9888);
nor UO_1025 (O_1025,N_9665,N_9061);
nor UO_1026 (O_1026,N_9165,N_9857);
nand UO_1027 (O_1027,N_9602,N_9408);
nor UO_1028 (O_1028,N_9376,N_9874);
nand UO_1029 (O_1029,N_9390,N_9398);
nand UO_1030 (O_1030,N_9373,N_9329);
or UO_1031 (O_1031,N_9104,N_9117);
nand UO_1032 (O_1032,N_9865,N_9427);
nor UO_1033 (O_1033,N_9350,N_9977);
nor UO_1034 (O_1034,N_9949,N_9076);
nand UO_1035 (O_1035,N_9813,N_9856);
or UO_1036 (O_1036,N_9637,N_9478);
nand UO_1037 (O_1037,N_9938,N_9320);
nor UO_1038 (O_1038,N_9411,N_9960);
nand UO_1039 (O_1039,N_9966,N_9652);
and UO_1040 (O_1040,N_9153,N_9370);
nor UO_1041 (O_1041,N_9823,N_9830);
nor UO_1042 (O_1042,N_9693,N_9482);
and UO_1043 (O_1043,N_9627,N_9933);
or UO_1044 (O_1044,N_9025,N_9912);
and UO_1045 (O_1045,N_9789,N_9690);
or UO_1046 (O_1046,N_9456,N_9648);
nor UO_1047 (O_1047,N_9001,N_9635);
nand UO_1048 (O_1048,N_9298,N_9660);
nand UO_1049 (O_1049,N_9582,N_9537);
nand UO_1050 (O_1050,N_9325,N_9122);
nand UO_1051 (O_1051,N_9980,N_9983);
or UO_1052 (O_1052,N_9168,N_9836);
nand UO_1053 (O_1053,N_9977,N_9990);
or UO_1054 (O_1054,N_9951,N_9191);
nand UO_1055 (O_1055,N_9269,N_9123);
and UO_1056 (O_1056,N_9787,N_9126);
nor UO_1057 (O_1057,N_9402,N_9083);
nand UO_1058 (O_1058,N_9796,N_9604);
or UO_1059 (O_1059,N_9874,N_9066);
or UO_1060 (O_1060,N_9018,N_9474);
and UO_1061 (O_1061,N_9969,N_9506);
nand UO_1062 (O_1062,N_9244,N_9756);
or UO_1063 (O_1063,N_9795,N_9547);
or UO_1064 (O_1064,N_9384,N_9304);
nand UO_1065 (O_1065,N_9812,N_9603);
nor UO_1066 (O_1066,N_9562,N_9652);
nor UO_1067 (O_1067,N_9154,N_9198);
and UO_1068 (O_1068,N_9319,N_9223);
or UO_1069 (O_1069,N_9933,N_9506);
xnor UO_1070 (O_1070,N_9991,N_9018);
nand UO_1071 (O_1071,N_9213,N_9183);
nand UO_1072 (O_1072,N_9467,N_9444);
nor UO_1073 (O_1073,N_9711,N_9298);
or UO_1074 (O_1074,N_9484,N_9573);
or UO_1075 (O_1075,N_9134,N_9266);
nor UO_1076 (O_1076,N_9179,N_9678);
or UO_1077 (O_1077,N_9833,N_9065);
nand UO_1078 (O_1078,N_9969,N_9498);
nand UO_1079 (O_1079,N_9549,N_9249);
and UO_1080 (O_1080,N_9857,N_9830);
or UO_1081 (O_1081,N_9794,N_9804);
nor UO_1082 (O_1082,N_9354,N_9341);
nand UO_1083 (O_1083,N_9215,N_9145);
and UO_1084 (O_1084,N_9775,N_9727);
and UO_1085 (O_1085,N_9197,N_9094);
nand UO_1086 (O_1086,N_9718,N_9810);
nand UO_1087 (O_1087,N_9462,N_9053);
and UO_1088 (O_1088,N_9747,N_9688);
nor UO_1089 (O_1089,N_9351,N_9394);
nand UO_1090 (O_1090,N_9526,N_9138);
nand UO_1091 (O_1091,N_9428,N_9710);
nor UO_1092 (O_1092,N_9844,N_9487);
and UO_1093 (O_1093,N_9615,N_9147);
and UO_1094 (O_1094,N_9746,N_9315);
nor UO_1095 (O_1095,N_9559,N_9824);
nand UO_1096 (O_1096,N_9194,N_9778);
nor UO_1097 (O_1097,N_9436,N_9671);
and UO_1098 (O_1098,N_9011,N_9587);
nand UO_1099 (O_1099,N_9723,N_9169);
and UO_1100 (O_1100,N_9736,N_9769);
nor UO_1101 (O_1101,N_9175,N_9387);
nor UO_1102 (O_1102,N_9620,N_9784);
nand UO_1103 (O_1103,N_9072,N_9117);
and UO_1104 (O_1104,N_9364,N_9495);
or UO_1105 (O_1105,N_9064,N_9618);
and UO_1106 (O_1106,N_9686,N_9169);
nor UO_1107 (O_1107,N_9229,N_9877);
and UO_1108 (O_1108,N_9689,N_9915);
nor UO_1109 (O_1109,N_9001,N_9996);
or UO_1110 (O_1110,N_9482,N_9010);
or UO_1111 (O_1111,N_9638,N_9088);
and UO_1112 (O_1112,N_9907,N_9748);
or UO_1113 (O_1113,N_9796,N_9230);
nor UO_1114 (O_1114,N_9089,N_9383);
nand UO_1115 (O_1115,N_9573,N_9190);
and UO_1116 (O_1116,N_9766,N_9577);
and UO_1117 (O_1117,N_9420,N_9436);
nand UO_1118 (O_1118,N_9626,N_9953);
nand UO_1119 (O_1119,N_9242,N_9071);
and UO_1120 (O_1120,N_9097,N_9952);
xnor UO_1121 (O_1121,N_9476,N_9492);
nand UO_1122 (O_1122,N_9891,N_9460);
nand UO_1123 (O_1123,N_9105,N_9702);
nand UO_1124 (O_1124,N_9384,N_9668);
or UO_1125 (O_1125,N_9092,N_9479);
or UO_1126 (O_1126,N_9312,N_9406);
and UO_1127 (O_1127,N_9510,N_9569);
nor UO_1128 (O_1128,N_9302,N_9915);
or UO_1129 (O_1129,N_9241,N_9813);
or UO_1130 (O_1130,N_9665,N_9556);
and UO_1131 (O_1131,N_9316,N_9557);
and UO_1132 (O_1132,N_9332,N_9731);
and UO_1133 (O_1133,N_9585,N_9347);
and UO_1134 (O_1134,N_9125,N_9190);
nor UO_1135 (O_1135,N_9345,N_9208);
or UO_1136 (O_1136,N_9853,N_9332);
nand UO_1137 (O_1137,N_9449,N_9973);
nor UO_1138 (O_1138,N_9439,N_9066);
nand UO_1139 (O_1139,N_9664,N_9865);
nor UO_1140 (O_1140,N_9375,N_9756);
nor UO_1141 (O_1141,N_9641,N_9800);
nor UO_1142 (O_1142,N_9008,N_9409);
and UO_1143 (O_1143,N_9700,N_9523);
or UO_1144 (O_1144,N_9739,N_9323);
and UO_1145 (O_1145,N_9339,N_9696);
nand UO_1146 (O_1146,N_9880,N_9597);
or UO_1147 (O_1147,N_9290,N_9002);
and UO_1148 (O_1148,N_9084,N_9444);
and UO_1149 (O_1149,N_9045,N_9217);
nand UO_1150 (O_1150,N_9849,N_9663);
and UO_1151 (O_1151,N_9133,N_9451);
or UO_1152 (O_1152,N_9354,N_9769);
or UO_1153 (O_1153,N_9072,N_9115);
nand UO_1154 (O_1154,N_9270,N_9910);
nor UO_1155 (O_1155,N_9922,N_9561);
or UO_1156 (O_1156,N_9883,N_9747);
or UO_1157 (O_1157,N_9582,N_9129);
nor UO_1158 (O_1158,N_9780,N_9685);
nand UO_1159 (O_1159,N_9105,N_9290);
or UO_1160 (O_1160,N_9894,N_9892);
nand UO_1161 (O_1161,N_9972,N_9615);
nand UO_1162 (O_1162,N_9142,N_9272);
and UO_1163 (O_1163,N_9921,N_9145);
nor UO_1164 (O_1164,N_9268,N_9241);
and UO_1165 (O_1165,N_9227,N_9086);
nor UO_1166 (O_1166,N_9619,N_9320);
xor UO_1167 (O_1167,N_9593,N_9934);
or UO_1168 (O_1168,N_9087,N_9109);
or UO_1169 (O_1169,N_9791,N_9277);
nor UO_1170 (O_1170,N_9351,N_9110);
and UO_1171 (O_1171,N_9836,N_9076);
nor UO_1172 (O_1172,N_9986,N_9717);
nor UO_1173 (O_1173,N_9279,N_9448);
nand UO_1174 (O_1174,N_9007,N_9518);
or UO_1175 (O_1175,N_9208,N_9168);
or UO_1176 (O_1176,N_9595,N_9498);
or UO_1177 (O_1177,N_9207,N_9591);
nand UO_1178 (O_1178,N_9150,N_9194);
nand UO_1179 (O_1179,N_9633,N_9731);
or UO_1180 (O_1180,N_9133,N_9311);
or UO_1181 (O_1181,N_9900,N_9825);
or UO_1182 (O_1182,N_9462,N_9335);
nor UO_1183 (O_1183,N_9353,N_9548);
or UO_1184 (O_1184,N_9646,N_9566);
or UO_1185 (O_1185,N_9591,N_9026);
nand UO_1186 (O_1186,N_9905,N_9699);
or UO_1187 (O_1187,N_9303,N_9152);
nor UO_1188 (O_1188,N_9241,N_9303);
nand UO_1189 (O_1189,N_9804,N_9978);
and UO_1190 (O_1190,N_9423,N_9884);
and UO_1191 (O_1191,N_9679,N_9250);
and UO_1192 (O_1192,N_9923,N_9390);
or UO_1193 (O_1193,N_9537,N_9825);
nand UO_1194 (O_1194,N_9114,N_9692);
and UO_1195 (O_1195,N_9690,N_9327);
nand UO_1196 (O_1196,N_9720,N_9130);
nor UO_1197 (O_1197,N_9532,N_9372);
nand UO_1198 (O_1198,N_9909,N_9715);
nand UO_1199 (O_1199,N_9158,N_9489);
nor UO_1200 (O_1200,N_9330,N_9115);
nand UO_1201 (O_1201,N_9468,N_9278);
nor UO_1202 (O_1202,N_9976,N_9274);
and UO_1203 (O_1203,N_9518,N_9429);
nand UO_1204 (O_1204,N_9801,N_9845);
and UO_1205 (O_1205,N_9020,N_9043);
nand UO_1206 (O_1206,N_9937,N_9943);
nor UO_1207 (O_1207,N_9263,N_9771);
nand UO_1208 (O_1208,N_9745,N_9606);
nor UO_1209 (O_1209,N_9268,N_9549);
or UO_1210 (O_1210,N_9060,N_9111);
nand UO_1211 (O_1211,N_9978,N_9063);
nand UO_1212 (O_1212,N_9084,N_9268);
nand UO_1213 (O_1213,N_9463,N_9815);
nand UO_1214 (O_1214,N_9396,N_9821);
nand UO_1215 (O_1215,N_9282,N_9902);
nor UO_1216 (O_1216,N_9107,N_9066);
nand UO_1217 (O_1217,N_9600,N_9538);
and UO_1218 (O_1218,N_9933,N_9780);
nor UO_1219 (O_1219,N_9135,N_9724);
nor UO_1220 (O_1220,N_9340,N_9107);
nand UO_1221 (O_1221,N_9756,N_9921);
nand UO_1222 (O_1222,N_9815,N_9682);
nor UO_1223 (O_1223,N_9146,N_9159);
or UO_1224 (O_1224,N_9684,N_9783);
nand UO_1225 (O_1225,N_9811,N_9680);
nand UO_1226 (O_1226,N_9146,N_9437);
nand UO_1227 (O_1227,N_9980,N_9046);
and UO_1228 (O_1228,N_9300,N_9120);
nand UO_1229 (O_1229,N_9845,N_9894);
or UO_1230 (O_1230,N_9162,N_9643);
nor UO_1231 (O_1231,N_9889,N_9633);
nand UO_1232 (O_1232,N_9065,N_9323);
nor UO_1233 (O_1233,N_9567,N_9771);
nand UO_1234 (O_1234,N_9894,N_9712);
and UO_1235 (O_1235,N_9300,N_9347);
nor UO_1236 (O_1236,N_9223,N_9067);
and UO_1237 (O_1237,N_9234,N_9837);
nand UO_1238 (O_1238,N_9354,N_9834);
and UO_1239 (O_1239,N_9777,N_9661);
nand UO_1240 (O_1240,N_9357,N_9139);
and UO_1241 (O_1241,N_9844,N_9169);
or UO_1242 (O_1242,N_9794,N_9458);
nor UO_1243 (O_1243,N_9648,N_9466);
and UO_1244 (O_1244,N_9761,N_9812);
or UO_1245 (O_1245,N_9282,N_9153);
nand UO_1246 (O_1246,N_9687,N_9593);
nand UO_1247 (O_1247,N_9061,N_9742);
nand UO_1248 (O_1248,N_9309,N_9175);
nand UO_1249 (O_1249,N_9912,N_9623);
or UO_1250 (O_1250,N_9339,N_9673);
nand UO_1251 (O_1251,N_9482,N_9140);
nand UO_1252 (O_1252,N_9645,N_9498);
and UO_1253 (O_1253,N_9410,N_9832);
nor UO_1254 (O_1254,N_9804,N_9928);
and UO_1255 (O_1255,N_9646,N_9409);
or UO_1256 (O_1256,N_9021,N_9066);
or UO_1257 (O_1257,N_9182,N_9198);
and UO_1258 (O_1258,N_9451,N_9325);
nor UO_1259 (O_1259,N_9256,N_9042);
or UO_1260 (O_1260,N_9009,N_9754);
or UO_1261 (O_1261,N_9767,N_9198);
nor UO_1262 (O_1262,N_9314,N_9697);
nor UO_1263 (O_1263,N_9306,N_9952);
nor UO_1264 (O_1264,N_9663,N_9399);
nor UO_1265 (O_1265,N_9912,N_9392);
and UO_1266 (O_1266,N_9240,N_9633);
and UO_1267 (O_1267,N_9066,N_9397);
or UO_1268 (O_1268,N_9942,N_9753);
nor UO_1269 (O_1269,N_9135,N_9361);
nor UO_1270 (O_1270,N_9608,N_9901);
or UO_1271 (O_1271,N_9958,N_9282);
or UO_1272 (O_1272,N_9638,N_9045);
nor UO_1273 (O_1273,N_9653,N_9691);
nor UO_1274 (O_1274,N_9555,N_9783);
nor UO_1275 (O_1275,N_9436,N_9114);
or UO_1276 (O_1276,N_9694,N_9372);
nand UO_1277 (O_1277,N_9896,N_9516);
xnor UO_1278 (O_1278,N_9443,N_9039);
and UO_1279 (O_1279,N_9840,N_9300);
or UO_1280 (O_1280,N_9308,N_9386);
or UO_1281 (O_1281,N_9661,N_9674);
nor UO_1282 (O_1282,N_9059,N_9176);
nand UO_1283 (O_1283,N_9726,N_9938);
or UO_1284 (O_1284,N_9319,N_9093);
or UO_1285 (O_1285,N_9777,N_9689);
and UO_1286 (O_1286,N_9247,N_9254);
and UO_1287 (O_1287,N_9779,N_9157);
nand UO_1288 (O_1288,N_9342,N_9332);
or UO_1289 (O_1289,N_9561,N_9604);
or UO_1290 (O_1290,N_9371,N_9240);
or UO_1291 (O_1291,N_9304,N_9640);
and UO_1292 (O_1292,N_9534,N_9334);
and UO_1293 (O_1293,N_9788,N_9561);
or UO_1294 (O_1294,N_9271,N_9612);
and UO_1295 (O_1295,N_9611,N_9755);
nand UO_1296 (O_1296,N_9689,N_9608);
nor UO_1297 (O_1297,N_9068,N_9258);
or UO_1298 (O_1298,N_9586,N_9925);
nand UO_1299 (O_1299,N_9024,N_9881);
nor UO_1300 (O_1300,N_9316,N_9584);
nand UO_1301 (O_1301,N_9403,N_9463);
or UO_1302 (O_1302,N_9175,N_9336);
or UO_1303 (O_1303,N_9201,N_9196);
nand UO_1304 (O_1304,N_9922,N_9454);
and UO_1305 (O_1305,N_9317,N_9869);
or UO_1306 (O_1306,N_9293,N_9442);
nor UO_1307 (O_1307,N_9141,N_9055);
nand UO_1308 (O_1308,N_9712,N_9213);
nand UO_1309 (O_1309,N_9364,N_9560);
or UO_1310 (O_1310,N_9319,N_9126);
nand UO_1311 (O_1311,N_9669,N_9501);
nor UO_1312 (O_1312,N_9428,N_9796);
nor UO_1313 (O_1313,N_9046,N_9963);
nor UO_1314 (O_1314,N_9610,N_9123);
nor UO_1315 (O_1315,N_9851,N_9681);
nand UO_1316 (O_1316,N_9795,N_9898);
and UO_1317 (O_1317,N_9318,N_9732);
nand UO_1318 (O_1318,N_9284,N_9404);
nor UO_1319 (O_1319,N_9264,N_9399);
or UO_1320 (O_1320,N_9780,N_9679);
or UO_1321 (O_1321,N_9232,N_9170);
nor UO_1322 (O_1322,N_9621,N_9541);
nor UO_1323 (O_1323,N_9447,N_9702);
or UO_1324 (O_1324,N_9617,N_9913);
and UO_1325 (O_1325,N_9668,N_9429);
or UO_1326 (O_1326,N_9307,N_9539);
and UO_1327 (O_1327,N_9170,N_9804);
nor UO_1328 (O_1328,N_9568,N_9456);
and UO_1329 (O_1329,N_9835,N_9444);
nor UO_1330 (O_1330,N_9158,N_9798);
nor UO_1331 (O_1331,N_9595,N_9548);
nor UO_1332 (O_1332,N_9200,N_9115);
or UO_1333 (O_1333,N_9488,N_9079);
nand UO_1334 (O_1334,N_9479,N_9280);
nand UO_1335 (O_1335,N_9417,N_9624);
nand UO_1336 (O_1336,N_9469,N_9246);
nand UO_1337 (O_1337,N_9415,N_9266);
nor UO_1338 (O_1338,N_9979,N_9579);
nor UO_1339 (O_1339,N_9839,N_9093);
nand UO_1340 (O_1340,N_9959,N_9607);
or UO_1341 (O_1341,N_9977,N_9452);
or UO_1342 (O_1342,N_9010,N_9552);
nand UO_1343 (O_1343,N_9113,N_9705);
and UO_1344 (O_1344,N_9754,N_9646);
or UO_1345 (O_1345,N_9302,N_9932);
and UO_1346 (O_1346,N_9793,N_9045);
and UO_1347 (O_1347,N_9108,N_9185);
and UO_1348 (O_1348,N_9999,N_9726);
nand UO_1349 (O_1349,N_9449,N_9304);
and UO_1350 (O_1350,N_9531,N_9750);
nor UO_1351 (O_1351,N_9094,N_9976);
nand UO_1352 (O_1352,N_9726,N_9338);
nand UO_1353 (O_1353,N_9999,N_9322);
and UO_1354 (O_1354,N_9477,N_9496);
nor UO_1355 (O_1355,N_9389,N_9453);
and UO_1356 (O_1356,N_9786,N_9745);
or UO_1357 (O_1357,N_9808,N_9497);
nand UO_1358 (O_1358,N_9805,N_9422);
and UO_1359 (O_1359,N_9409,N_9700);
nor UO_1360 (O_1360,N_9288,N_9768);
or UO_1361 (O_1361,N_9146,N_9801);
nand UO_1362 (O_1362,N_9666,N_9011);
or UO_1363 (O_1363,N_9400,N_9715);
or UO_1364 (O_1364,N_9795,N_9486);
and UO_1365 (O_1365,N_9849,N_9975);
and UO_1366 (O_1366,N_9184,N_9802);
nor UO_1367 (O_1367,N_9835,N_9647);
nor UO_1368 (O_1368,N_9361,N_9786);
nor UO_1369 (O_1369,N_9963,N_9155);
or UO_1370 (O_1370,N_9987,N_9619);
nand UO_1371 (O_1371,N_9083,N_9087);
and UO_1372 (O_1372,N_9089,N_9054);
and UO_1373 (O_1373,N_9033,N_9124);
or UO_1374 (O_1374,N_9941,N_9429);
and UO_1375 (O_1375,N_9471,N_9804);
and UO_1376 (O_1376,N_9268,N_9661);
or UO_1377 (O_1377,N_9373,N_9000);
nor UO_1378 (O_1378,N_9343,N_9707);
nor UO_1379 (O_1379,N_9989,N_9210);
and UO_1380 (O_1380,N_9299,N_9129);
nor UO_1381 (O_1381,N_9721,N_9016);
nand UO_1382 (O_1382,N_9127,N_9347);
and UO_1383 (O_1383,N_9595,N_9832);
nor UO_1384 (O_1384,N_9155,N_9886);
xnor UO_1385 (O_1385,N_9855,N_9402);
nor UO_1386 (O_1386,N_9475,N_9169);
nand UO_1387 (O_1387,N_9209,N_9328);
nand UO_1388 (O_1388,N_9610,N_9623);
and UO_1389 (O_1389,N_9482,N_9312);
nand UO_1390 (O_1390,N_9929,N_9247);
or UO_1391 (O_1391,N_9884,N_9644);
nor UO_1392 (O_1392,N_9189,N_9278);
nand UO_1393 (O_1393,N_9349,N_9931);
or UO_1394 (O_1394,N_9640,N_9137);
nand UO_1395 (O_1395,N_9611,N_9183);
and UO_1396 (O_1396,N_9526,N_9680);
nor UO_1397 (O_1397,N_9966,N_9497);
nand UO_1398 (O_1398,N_9718,N_9400);
nand UO_1399 (O_1399,N_9021,N_9776);
nand UO_1400 (O_1400,N_9394,N_9493);
and UO_1401 (O_1401,N_9114,N_9003);
nor UO_1402 (O_1402,N_9042,N_9531);
nor UO_1403 (O_1403,N_9312,N_9993);
nor UO_1404 (O_1404,N_9036,N_9293);
nand UO_1405 (O_1405,N_9341,N_9100);
or UO_1406 (O_1406,N_9123,N_9274);
nor UO_1407 (O_1407,N_9736,N_9777);
or UO_1408 (O_1408,N_9729,N_9595);
nand UO_1409 (O_1409,N_9581,N_9320);
or UO_1410 (O_1410,N_9908,N_9311);
and UO_1411 (O_1411,N_9026,N_9444);
or UO_1412 (O_1412,N_9511,N_9213);
nor UO_1413 (O_1413,N_9847,N_9650);
and UO_1414 (O_1414,N_9418,N_9295);
nand UO_1415 (O_1415,N_9510,N_9576);
or UO_1416 (O_1416,N_9118,N_9986);
and UO_1417 (O_1417,N_9375,N_9535);
or UO_1418 (O_1418,N_9945,N_9219);
or UO_1419 (O_1419,N_9637,N_9756);
or UO_1420 (O_1420,N_9854,N_9106);
nand UO_1421 (O_1421,N_9523,N_9120);
and UO_1422 (O_1422,N_9942,N_9182);
or UO_1423 (O_1423,N_9635,N_9126);
nand UO_1424 (O_1424,N_9853,N_9618);
xnor UO_1425 (O_1425,N_9099,N_9389);
nor UO_1426 (O_1426,N_9515,N_9728);
and UO_1427 (O_1427,N_9881,N_9160);
nand UO_1428 (O_1428,N_9812,N_9355);
nor UO_1429 (O_1429,N_9761,N_9142);
and UO_1430 (O_1430,N_9225,N_9789);
and UO_1431 (O_1431,N_9173,N_9499);
nand UO_1432 (O_1432,N_9889,N_9849);
nor UO_1433 (O_1433,N_9532,N_9121);
or UO_1434 (O_1434,N_9135,N_9147);
nand UO_1435 (O_1435,N_9827,N_9789);
and UO_1436 (O_1436,N_9185,N_9568);
nor UO_1437 (O_1437,N_9316,N_9649);
or UO_1438 (O_1438,N_9200,N_9887);
nand UO_1439 (O_1439,N_9967,N_9109);
nor UO_1440 (O_1440,N_9001,N_9694);
nand UO_1441 (O_1441,N_9940,N_9049);
and UO_1442 (O_1442,N_9684,N_9422);
and UO_1443 (O_1443,N_9880,N_9050);
or UO_1444 (O_1444,N_9457,N_9762);
and UO_1445 (O_1445,N_9459,N_9317);
and UO_1446 (O_1446,N_9606,N_9413);
nor UO_1447 (O_1447,N_9227,N_9391);
nor UO_1448 (O_1448,N_9502,N_9339);
or UO_1449 (O_1449,N_9568,N_9552);
or UO_1450 (O_1450,N_9972,N_9569);
nor UO_1451 (O_1451,N_9145,N_9717);
nand UO_1452 (O_1452,N_9603,N_9031);
nor UO_1453 (O_1453,N_9928,N_9019);
nor UO_1454 (O_1454,N_9317,N_9440);
and UO_1455 (O_1455,N_9061,N_9859);
nor UO_1456 (O_1456,N_9582,N_9343);
or UO_1457 (O_1457,N_9008,N_9519);
nand UO_1458 (O_1458,N_9862,N_9327);
nand UO_1459 (O_1459,N_9872,N_9666);
nand UO_1460 (O_1460,N_9224,N_9365);
and UO_1461 (O_1461,N_9758,N_9009);
nand UO_1462 (O_1462,N_9020,N_9527);
or UO_1463 (O_1463,N_9443,N_9535);
or UO_1464 (O_1464,N_9158,N_9535);
nand UO_1465 (O_1465,N_9558,N_9801);
nand UO_1466 (O_1466,N_9128,N_9220);
or UO_1467 (O_1467,N_9771,N_9111);
nand UO_1468 (O_1468,N_9548,N_9521);
and UO_1469 (O_1469,N_9662,N_9222);
and UO_1470 (O_1470,N_9975,N_9030);
and UO_1471 (O_1471,N_9409,N_9945);
and UO_1472 (O_1472,N_9414,N_9787);
nor UO_1473 (O_1473,N_9103,N_9515);
nand UO_1474 (O_1474,N_9076,N_9699);
and UO_1475 (O_1475,N_9326,N_9764);
nand UO_1476 (O_1476,N_9751,N_9039);
and UO_1477 (O_1477,N_9795,N_9389);
nor UO_1478 (O_1478,N_9014,N_9061);
nand UO_1479 (O_1479,N_9853,N_9895);
nand UO_1480 (O_1480,N_9065,N_9948);
or UO_1481 (O_1481,N_9425,N_9620);
and UO_1482 (O_1482,N_9300,N_9476);
and UO_1483 (O_1483,N_9087,N_9239);
nor UO_1484 (O_1484,N_9249,N_9748);
or UO_1485 (O_1485,N_9276,N_9848);
or UO_1486 (O_1486,N_9461,N_9663);
or UO_1487 (O_1487,N_9621,N_9821);
nor UO_1488 (O_1488,N_9911,N_9288);
nand UO_1489 (O_1489,N_9851,N_9696);
nor UO_1490 (O_1490,N_9549,N_9068);
and UO_1491 (O_1491,N_9101,N_9959);
nand UO_1492 (O_1492,N_9676,N_9463);
nor UO_1493 (O_1493,N_9583,N_9959);
nor UO_1494 (O_1494,N_9214,N_9324);
nand UO_1495 (O_1495,N_9022,N_9770);
nor UO_1496 (O_1496,N_9174,N_9581);
nor UO_1497 (O_1497,N_9851,N_9142);
xnor UO_1498 (O_1498,N_9984,N_9694);
nand UO_1499 (O_1499,N_9071,N_9398);
endmodule