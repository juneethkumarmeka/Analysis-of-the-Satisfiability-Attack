module basic_500_3000_500_6_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_42,In_317);
or U1 (N_1,In_427,In_55);
nand U2 (N_2,In_145,In_378);
nor U3 (N_3,In_494,In_220);
nand U4 (N_4,In_355,In_298);
nor U5 (N_5,In_177,In_375);
and U6 (N_6,In_80,In_58);
nor U7 (N_7,In_96,In_283);
or U8 (N_8,In_37,In_117);
and U9 (N_9,In_361,In_119);
and U10 (N_10,In_280,In_10);
and U11 (N_11,In_471,In_174);
nor U12 (N_12,In_473,In_67);
nor U13 (N_13,In_12,In_325);
or U14 (N_14,In_402,In_82);
nand U15 (N_15,In_141,In_104);
nand U16 (N_16,In_328,In_321);
and U17 (N_17,In_28,In_159);
nand U18 (N_18,In_374,In_423);
and U19 (N_19,In_386,In_17);
and U20 (N_20,In_199,In_138);
or U21 (N_21,In_105,In_201);
or U22 (N_22,In_435,In_163);
nor U23 (N_23,In_384,In_343);
or U24 (N_24,In_115,In_479);
nand U25 (N_25,In_33,In_20);
nor U26 (N_26,In_172,In_287);
nand U27 (N_27,In_327,In_196);
or U28 (N_28,In_120,In_26);
or U29 (N_29,In_225,In_249);
and U30 (N_30,In_106,In_292);
and U31 (N_31,In_164,In_38);
and U32 (N_32,In_468,In_122);
and U33 (N_33,In_417,In_493);
or U34 (N_34,In_244,In_185);
or U35 (N_35,In_478,In_277);
or U36 (N_36,In_459,In_0);
nand U37 (N_37,In_415,In_202);
and U38 (N_38,In_245,In_475);
nand U39 (N_39,In_359,In_416);
nor U40 (N_40,In_306,In_31);
nand U41 (N_41,In_438,In_226);
nor U42 (N_42,In_125,In_397);
nand U43 (N_43,In_456,In_398);
nand U44 (N_44,In_383,In_482);
or U45 (N_45,In_276,In_440);
or U46 (N_46,In_318,In_83);
and U47 (N_47,In_144,In_345);
nor U48 (N_48,In_360,In_186);
or U49 (N_49,In_218,In_68);
nand U50 (N_50,In_480,In_235);
or U51 (N_51,In_78,In_29);
or U52 (N_52,In_200,In_162);
nand U53 (N_53,In_319,In_166);
nand U54 (N_54,In_338,In_3);
nand U55 (N_55,In_380,In_123);
or U56 (N_56,In_103,In_279);
nand U57 (N_57,In_290,In_194);
nand U58 (N_58,In_266,In_254);
or U59 (N_59,In_56,In_34);
nor U60 (N_60,In_430,In_93);
or U61 (N_61,In_382,In_87);
nor U62 (N_62,In_333,In_214);
nand U63 (N_63,In_44,In_323);
and U64 (N_64,In_264,In_442);
and U65 (N_65,In_453,In_489);
or U66 (N_66,In_25,In_19);
nor U67 (N_67,In_134,In_448);
or U68 (N_68,In_227,In_248);
xor U69 (N_69,In_498,In_59);
and U70 (N_70,In_253,In_14);
nand U71 (N_71,In_392,In_91);
or U72 (N_72,In_484,In_446);
or U73 (N_73,In_161,In_414);
nand U74 (N_74,In_110,In_272);
nand U75 (N_75,In_45,In_296);
and U76 (N_76,In_242,In_350);
nor U77 (N_77,In_326,In_128);
and U78 (N_78,In_307,In_77);
nor U79 (N_79,In_358,In_195);
or U80 (N_80,In_173,In_90);
and U81 (N_81,In_289,In_140);
nand U82 (N_82,In_499,In_262);
nor U83 (N_83,In_455,In_314);
nor U84 (N_84,In_250,In_267);
nand U85 (N_85,In_39,In_458);
or U86 (N_86,In_63,In_291);
nand U87 (N_87,In_109,In_270);
nand U88 (N_88,In_233,In_5);
nand U89 (N_89,In_370,In_396);
or U90 (N_90,In_6,In_373);
or U91 (N_91,In_139,In_452);
and U92 (N_92,In_352,In_234);
or U93 (N_93,In_488,In_303);
nand U94 (N_94,In_222,In_313);
or U95 (N_95,In_183,In_401);
xnor U96 (N_96,In_192,In_481);
and U97 (N_97,In_189,In_27);
and U98 (N_98,In_1,In_21);
or U99 (N_99,In_36,In_219);
nand U100 (N_100,In_221,In_239);
nor U101 (N_101,In_2,In_454);
nor U102 (N_102,In_205,In_238);
nand U103 (N_103,In_330,In_111);
nand U104 (N_104,In_433,In_335);
nor U105 (N_105,In_15,In_432);
or U106 (N_106,In_50,In_190);
and U107 (N_107,In_76,In_217);
and U108 (N_108,In_390,In_408);
and U109 (N_109,In_278,In_342);
nor U110 (N_110,In_403,In_142);
and U111 (N_111,In_465,In_40);
or U112 (N_112,In_150,In_395);
nor U113 (N_113,In_419,In_208);
or U114 (N_114,In_132,In_391);
or U115 (N_115,In_247,In_348);
or U116 (N_116,In_236,In_477);
and U117 (N_117,In_320,In_75);
and U118 (N_118,In_344,In_170);
or U119 (N_119,In_85,In_153);
or U120 (N_120,In_255,In_400);
nor U121 (N_121,In_223,In_310);
nand U122 (N_122,In_89,In_241);
and U123 (N_123,In_4,In_337);
or U124 (N_124,In_30,In_260);
nand U125 (N_125,In_169,In_47);
and U126 (N_126,In_389,In_197);
nor U127 (N_127,In_251,In_444);
and U128 (N_128,In_116,In_288);
and U129 (N_129,In_347,In_127);
or U130 (N_130,In_193,In_175);
xor U131 (N_131,In_357,In_315);
or U132 (N_132,In_246,In_441);
nand U133 (N_133,In_381,In_450);
and U134 (N_134,In_421,In_469);
or U135 (N_135,In_304,In_215);
nor U136 (N_136,In_377,In_336);
or U137 (N_137,In_302,In_86);
nor U138 (N_138,In_79,In_451);
nor U139 (N_139,In_351,In_213);
and U140 (N_140,In_496,In_439);
nand U141 (N_141,In_486,In_7);
nor U142 (N_142,In_461,In_113);
or U143 (N_143,In_102,In_228);
and U144 (N_144,In_467,In_420);
nor U145 (N_145,In_369,In_230);
and U146 (N_146,In_407,In_346);
nand U147 (N_147,In_284,In_340);
or U148 (N_148,In_273,In_309);
and U149 (N_149,In_495,In_299);
or U150 (N_150,In_387,In_275);
or U151 (N_151,In_457,In_154);
nor U152 (N_152,In_88,In_107);
nor U153 (N_153,In_155,In_112);
nor U154 (N_154,In_70,In_269);
and U155 (N_155,In_41,In_371);
nor U156 (N_156,In_294,In_129);
or U157 (N_157,In_379,In_232);
nor U158 (N_158,In_256,In_43);
xor U159 (N_159,In_312,In_341);
or U160 (N_160,In_405,In_365);
and U161 (N_161,In_472,In_464);
nor U162 (N_162,In_188,In_434);
nand U163 (N_163,In_368,In_490);
nand U164 (N_164,In_274,In_372);
or U165 (N_165,In_148,In_388);
and U166 (N_166,In_470,In_334);
and U167 (N_167,In_206,In_412);
nor U168 (N_168,In_49,In_426);
nand U169 (N_169,In_285,In_62);
nor U170 (N_170,In_331,In_376);
nor U171 (N_171,In_293,In_108);
and U172 (N_172,In_460,In_60);
nor U173 (N_173,In_497,In_353);
and U174 (N_174,In_101,In_257);
nand U175 (N_175,In_11,In_73);
nand U176 (N_176,In_261,In_137);
xnor U177 (N_177,In_363,In_135);
nand U178 (N_178,In_243,In_133);
nand U179 (N_179,In_316,In_210);
or U180 (N_180,In_126,In_281);
nor U181 (N_181,In_124,In_362);
or U182 (N_182,In_176,In_66);
nand U183 (N_183,In_297,In_443);
or U184 (N_184,In_394,In_366);
and U185 (N_185,In_84,In_354);
nand U186 (N_186,In_118,In_425);
and U187 (N_187,In_268,In_385);
or U188 (N_188,In_237,In_259);
nor U189 (N_189,In_178,In_52);
and U190 (N_190,In_436,In_413);
or U191 (N_191,In_282,In_179);
nand U192 (N_192,In_447,In_411);
or U193 (N_193,In_187,In_18);
nand U194 (N_194,In_209,In_157);
nor U195 (N_195,In_212,In_171);
nor U196 (N_196,In_466,In_393);
or U197 (N_197,In_81,In_305);
and U198 (N_198,In_329,In_224);
nand U199 (N_199,In_9,In_308);
and U200 (N_200,In_152,In_399);
and U201 (N_201,In_474,In_130);
or U202 (N_202,In_485,In_445);
nor U203 (N_203,In_53,In_74);
nor U204 (N_204,In_182,In_492);
or U205 (N_205,In_286,In_32);
or U206 (N_206,In_160,In_191);
nand U207 (N_207,In_24,In_198);
and U208 (N_208,In_143,In_311);
nand U209 (N_209,In_146,In_491);
or U210 (N_210,In_165,In_449);
and U211 (N_211,In_356,In_211);
nand U212 (N_212,In_48,In_72);
and U213 (N_213,In_240,In_184);
nor U214 (N_214,In_339,In_424);
xnor U215 (N_215,In_149,In_35);
nor U216 (N_216,In_13,In_151);
nor U217 (N_217,In_406,In_94);
or U218 (N_218,In_462,In_367);
or U219 (N_219,In_156,In_295);
and U220 (N_220,In_69,In_332);
or U221 (N_221,In_168,In_410);
or U222 (N_222,In_61,In_100);
or U223 (N_223,In_437,In_54);
nor U224 (N_224,In_180,In_231);
or U225 (N_225,In_64,In_463);
or U226 (N_226,In_324,In_349);
or U227 (N_227,In_98,In_258);
nand U228 (N_228,In_229,In_99);
or U229 (N_229,In_114,In_428);
nand U230 (N_230,In_121,In_23);
and U231 (N_231,In_487,In_476);
nor U232 (N_232,In_216,In_95);
nor U233 (N_233,In_271,In_300);
nor U234 (N_234,In_46,In_422);
nand U235 (N_235,In_51,In_92);
or U236 (N_236,In_97,In_147);
nor U237 (N_237,In_483,In_207);
or U238 (N_238,In_204,In_322);
nand U239 (N_239,In_71,In_409);
nor U240 (N_240,In_131,In_16);
nand U241 (N_241,In_431,In_418);
nor U242 (N_242,In_252,In_158);
or U243 (N_243,In_22,In_429);
nor U244 (N_244,In_181,In_404);
nor U245 (N_245,In_8,In_65);
or U246 (N_246,In_263,In_265);
or U247 (N_247,In_203,In_364);
nor U248 (N_248,In_301,In_167);
nand U249 (N_249,In_136,In_57);
and U250 (N_250,In_385,In_412);
nand U251 (N_251,In_93,In_362);
or U252 (N_252,In_230,In_3);
or U253 (N_253,In_248,In_123);
or U254 (N_254,In_374,In_425);
xor U255 (N_255,In_452,In_396);
or U256 (N_256,In_453,In_320);
and U257 (N_257,In_317,In_331);
nor U258 (N_258,In_61,In_384);
nor U259 (N_259,In_466,In_404);
nand U260 (N_260,In_199,In_320);
nand U261 (N_261,In_367,In_357);
nand U262 (N_262,In_335,In_110);
nand U263 (N_263,In_327,In_250);
nand U264 (N_264,In_427,In_72);
or U265 (N_265,In_154,In_236);
nor U266 (N_266,In_379,In_82);
and U267 (N_267,In_295,In_497);
nor U268 (N_268,In_457,In_19);
nor U269 (N_269,In_0,In_475);
or U270 (N_270,In_182,In_391);
xnor U271 (N_271,In_48,In_492);
nand U272 (N_272,In_247,In_134);
nor U273 (N_273,In_230,In_363);
nand U274 (N_274,In_24,In_61);
and U275 (N_275,In_100,In_341);
nand U276 (N_276,In_13,In_454);
nor U277 (N_277,In_210,In_9);
or U278 (N_278,In_255,In_265);
nand U279 (N_279,In_252,In_476);
nor U280 (N_280,In_273,In_397);
and U281 (N_281,In_370,In_12);
and U282 (N_282,In_315,In_64);
nand U283 (N_283,In_72,In_339);
nor U284 (N_284,In_35,In_252);
or U285 (N_285,In_264,In_118);
and U286 (N_286,In_138,In_477);
or U287 (N_287,In_24,In_393);
and U288 (N_288,In_410,In_256);
nor U289 (N_289,In_260,In_304);
or U290 (N_290,In_141,In_41);
or U291 (N_291,In_24,In_362);
or U292 (N_292,In_399,In_432);
or U293 (N_293,In_429,In_279);
or U294 (N_294,In_101,In_494);
nand U295 (N_295,In_422,In_343);
and U296 (N_296,In_88,In_458);
or U297 (N_297,In_280,In_374);
or U298 (N_298,In_145,In_150);
nand U299 (N_299,In_174,In_203);
xnor U300 (N_300,In_44,In_281);
or U301 (N_301,In_8,In_459);
nand U302 (N_302,In_469,In_245);
nor U303 (N_303,In_75,In_19);
or U304 (N_304,In_278,In_213);
and U305 (N_305,In_125,In_37);
nor U306 (N_306,In_260,In_347);
and U307 (N_307,In_182,In_397);
and U308 (N_308,In_107,In_158);
and U309 (N_309,In_358,In_343);
and U310 (N_310,In_271,In_177);
or U311 (N_311,In_417,In_451);
and U312 (N_312,In_5,In_471);
or U313 (N_313,In_93,In_329);
and U314 (N_314,In_166,In_316);
and U315 (N_315,In_399,In_424);
nand U316 (N_316,In_197,In_491);
nand U317 (N_317,In_468,In_56);
nor U318 (N_318,In_307,In_342);
xnor U319 (N_319,In_72,In_304);
and U320 (N_320,In_288,In_181);
or U321 (N_321,In_215,In_270);
nand U322 (N_322,In_314,In_442);
nand U323 (N_323,In_311,In_338);
nor U324 (N_324,In_280,In_59);
and U325 (N_325,In_402,In_249);
nand U326 (N_326,In_497,In_345);
nand U327 (N_327,In_381,In_278);
or U328 (N_328,In_261,In_230);
and U329 (N_329,In_370,In_369);
nand U330 (N_330,In_212,In_267);
nor U331 (N_331,In_298,In_427);
and U332 (N_332,In_252,In_391);
and U333 (N_333,In_427,In_211);
or U334 (N_334,In_49,In_293);
and U335 (N_335,In_104,In_258);
nand U336 (N_336,In_129,In_356);
and U337 (N_337,In_472,In_8);
xnor U338 (N_338,In_90,In_248);
and U339 (N_339,In_270,In_318);
nor U340 (N_340,In_131,In_339);
or U341 (N_341,In_287,In_276);
or U342 (N_342,In_3,In_169);
and U343 (N_343,In_387,In_226);
nand U344 (N_344,In_228,In_300);
nor U345 (N_345,In_228,In_339);
and U346 (N_346,In_256,In_104);
and U347 (N_347,In_412,In_310);
and U348 (N_348,In_430,In_378);
and U349 (N_349,In_280,In_58);
nor U350 (N_350,In_89,In_156);
nor U351 (N_351,In_341,In_6);
and U352 (N_352,In_3,In_240);
or U353 (N_353,In_383,In_325);
nand U354 (N_354,In_45,In_189);
xor U355 (N_355,In_295,In_239);
nor U356 (N_356,In_186,In_385);
xor U357 (N_357,In_377,In_497);
nand U358 (N_358,In_4,In_309);
nor U359 (N_359,In_443,In_427);
and U360 (N_360,In_415,In_317);
nor U361 (N_361,In_179,In_481);
and U362 (N_362,In_190,In_480);
nor U363 (N_363,In_367,In_454);
or U364 (N_364,In_167,In_140);
nand U365 (N_365,In_483,In_338);
nand U366 (N_366,In_16,In_452);
or U367 (N_367,In_210,In_393);
or U368 (N_368,In_279,In_434);
or U369 (N_369,In_496,In_448);
nand U370 (N_370,In_389,In_38);
and U371 (N_371,In_281,In_286);
nand U372 (N_372,In_186,In_275);
and U373 (N_373,In_331,In_499);
and U374 (N_374,In_385,In_254);
nand U375 (N_375,In_81,In_381);
nand U376 (N_376,In_323,In_95);
or U377 (N_377,In_232,In_54);
or U378 (N_378,In_52,In_21);
or U379 (N_379,In_202,In_345);
and U380 (N_380,In_394,In_432);
or U381 (N_381,In_45,In_53);
and U382 (N_382,In_183,In_301);
or U383 (N_383,In_267,In_328);
nor U384 (N_384,In_201,In_196);
and U385 (N_385,In_140,In_494);
nand U386 (N_386,In_490,In_472);
nand U387 (N_387,In_82,In_419);
and U388 (N_388,In_276,In_80);
nor U389 (N_389,In_52,In_207);
nor U390 (N_390,In_418,In_61);
nand U391 (N_391,In_461,In_132);
or U392 (N_392,In_294,In_282);
or U393 (N_393,In_354,In_122);
or U394 (N_394,In_142,In_166);
nor U395 (N_395,In_319,In_164);
or U396 (N_396,In_159,In_24);
or U397 (N_397,In_315,In_270);
or U398 (N_398,In_336,In_309);
and U399 (N_399,In_357,In_124);
and U400 (N_400,In_344,In_490);
nand U401 (N_401,In_364,In_285);
and U402 (N_402,In_426,In_420);
or U403 (N_403,In_200,In_74);
and U404 (N_404,In_286,In_343);
nand U405 (N_405,In_354,In_487);
nor U406 (N_406,In_93,In_152);
nor U407 (N_407,In_151,In_186);
or U408 (N_408,In_368,In_202);
nand U409 (N_409,In_355,In_82);
nor U410 (N_410,In_168,In_418);
nand U411 (N_411,In_319,In_91);
and U412 (N_412,In_408,In_258);
and U413 (N_413,In_267,In_92);
or U414 (N_414,In_459,In_279);
nor U415 (N_415,In_303,In_193);
or U416 (N_416,In_422,In_355);
nand U417 (N_417,In_104,In_180);
nor U418 (N_418,In_0,In_249);
nor U419 (N_419,In_104,In_17);
xnor U420 (N_420,In_171,In_83);
nor U421 (N_421,In_190,In_346);
nand U422 (N_422,In_374,In_329);
nand U423 (N_423,In_439,In_282);
or U424 (N_424,In_445,In_336);
nor U425 (N_425,In_186,In_121);
and U426 (N_426,In_43,In_71);
or U427 (N_427,In_455,In_285);
or U428 (N_428,In_155,In_98);
nor U429 (N_429,In_484,In_478);
or U430 (N_430,In_440,In_182);
or U431 (N_431,In_5,In_100);
or U432 (N_432,In_398,In_454);
nand U433 (N_433,In_175,In_404);
or U434 (N_434,In_297,In_35);
nand U435 (N_435,In_450,In_21);
or U436 (N_436,In_256,In_333);
or U437 (N_437,In_461,In_112);
or U438 (N_438,In_126,In_382);
or U439 (N_439,In_295,In_35);
nor U440 (N_440,In_369,In_379);
nor U441 (N_441,In_421,In_383);
nand U442 (N_442,In_432,In_474);
and U443 (N_443,In_466,In_418);
or U444 (N_444,In_341,In_323);
nand U445 (N_445,In_155,In_18);
and U446 (N_446,In_381,In_413);
nand U447 (N_447,In_223,In_463);
nor U448 (N_448,In_239,In_40);
or U449 (N_449,In_408,In_386);
and U450 (N_450,In_349,In_219);
nor U451 (N_451,In_38,In_287);
and U452 (N_452,In_16,In_127);
or U453 (N_453,In_446,In_196);
nand U454 (N_454,In_250,In_197);
nor U455 (N_455,In_193,In_288);
or U456 (N_456,In_1,In_99);
and U457 (N_457,In_346,In_37);
and U458 (N_458,In_110,In_284);
and U459 (N_459,In_148,In_461);
nor U460 (N_460,In_414,In_328);
and U461 (N_461,In_396,In_332);
and U462 (N_462,In_216,In_219);
or U463 (N_463,In_364,In_212);
nand U464 (N_464,In_448,In_201);
or U465 (N_465,In_209,In_40);
nor U466 (N_466,In_412,In_480);
nand U467 (N_467,In_449,In_68);
nor U468 (N_468,In_30,In_85);
nand U469 (N_469,In_128,In_448);
or U470 (N_470,In_20,In_200);
and U471 (N_471,In_265,In_32);
or U472 (N_472,In_196,In_384);
or U473 (N_473,In_218,In_344);
and U474 (N_474,In_90,In_357);
and U475 (N_475,In_219,In_443);
xor U476 (N_476,In_186,In_487);
and U477 (N_477,In_99,In_18);
or U478 (N_478,In_454,In_355);
nor U479 (N_479,In_485,In_193);
and U480 (N_480,In_132,In_92);
or U481 (N_481,In_323,In_250);
nor U482 (N_482,In_120,In_236);
nand U483 (N_483,In_350,In_217);
nand U484 (N_484,In_448,In_288);
nor U485 (N_485,In_60,In_91);
and U486 (N_486,In_259,In_452);
nor U487 (N_487,In_88,In_97);
nand U488 (N_488,In_95,In_58);
and U489 (N_489,In_107,In_23);
and U490 (N_490,In_141,In_469);
and U491 (N_491,In_215,In_201);
nor U492 (N_492,In_317,In_214);
or U493 (N_493,In_73,In_4);
or U494 (N_494,In_483,In_488);
nor U495 (N_495,In_379,In_244);
nor U496 (N_496,In_346,In_72);
and U497 (N_497,In_3,In_403);
nand U498 (N_498,In_348,In_448);
nand U499 (N_499,In_195,In_203);
nor U500 (N_500,N_382,N_137);
nor U501 (N_501,N_442,N_205);
or U502 (N_502,N_84,N_39);
nand U503 (N_503,N_269,N_30);
and U504 (N_504,N_206,N_149);
nand U505 (N_505,N_289,N_15);
nor U506 (N_506,N_241,N_257);
or U507 (N_507,N_83,N_409);
xnor U508 (N_508,N_325,N_316);
nand U509 (N_509,N_197,N_450);
or U510 (N_510,N_247,N_422);
nand U511 (N_511,N_35,N_377);
and U512 (N_512,N_102,N_48);
nand U513 (N_513,N_100,N_221);
or U514 (N_514,N_421,N_473);
nand U515 (N_515,N_98,N_152);
nand U516 (N_516,N_435,N_375);
and U517 (N_517,N_5,N_181);
or U518 (N_518,N_90,N_55);
or U519 (N_519,N_267,N_348);
nand U520 (N_520,N_82,N_238);
nor U521 (N_521,N_258,N_327);
or U522 (N_522,N_338,N_309);
and U523 (N_523,N_346,N_331);
nor U524 (N_524,N_185,N_79);
nor U525 (N_525,N_232,N_352);
and U526 (N_526,N_158,N_318);
and U527 (N_527,N_298,N_337);
nand U528 (N_528,N_488,N_16);
and U529 (N_529,N_339,N_68);
nor U530 (N_530,N_196,N_191);
nor U531 (N_531,N_203,N_417);
nor U532 (N_532,N_198,N_193);
and U533 (N_533,N_343,N_307);
nor U534 (N_534,N_391,N_460);
nand U535 (N_535,N_493,N_277);
nor U536 (N_536,N_118,N_109);
nor U537 (N_537,N_256,N_385);
nor U538 (N_538,N_264,N_380);
or U539 (N_539,N_4,N_354);
nand U540 (N_540,N_73,N_296);
nand U541 (N_541,N_487,N_312);
nand U542 (N_542,N_93,N_279);
nor U543 (N_543,N_92,N_263);
nand U544 (N_544,N_456,N_373);
or U545 (N_545,N_495,N_379);
and U546 (N_546,N_46,N_461);
nand U547 (N_547,N_411,N_472);
and U548 (N_548,N_47,N_266);
or U549 (N_549,N_103,N_278);
nand U550 (N_550,N_283,N_475);
xnor U551 (N_551,N_321,N_174);
nor U552 (N_552,N_175,N_433);
or U553 (N_553,N_58,N_349);
and U554 (N_554,N_42,N_313);
or U555 (N_555,N_280,N_177);
nor U556 (N_556,N_317,N_288);
nand U557 (N_557,N_243,N_392);
nor U558 (N_558,N_437,N_222);
nand U559 (N_559,N_11,N_482);
nand U560 (N_560,N_228,N_169);
nand U561 (N_561,N_53,N_301);
nor U562 (N_562,N_453,N_388);
and U563 (N_563,N_115,N_110);
and U564 (N_564,N_432,N_335);
and U565 (N_565,N_308,N_397);
nand U566 (N_566,N_81,N_50);
or U567 (N_567,N_399,N_424);
and U568 (N_568,N_201,N_129);
nor U569 (N_569,N_220,N_416);
nand U570 (N_570,N_239,N_101);
nor U571 (N_571,N_297,N_275);
nor U572 (N_572,N_31,N_124);
and U573 (N_573,N_383,N_237);
or U574 (N_574,N_489,N_390);
and U575 (N_575,N_326,N_368);
nand U576 (N_576,N_479,N_80);
and U577 (N_577,N_12,N_230);
nand U578 (N_578,N_272,N_187);
or U579 (N_579,N_131,N_125);
and U580 (N_580,N_95,N_150);
or U581 (N_581,N_414,N_29);
and U582 (N_582,N_104,N_28);
or U583 (N_583,N_134,N_285);
nand U584 (N_584,N_86,N_358);
and U585 (N_585,N_67,N_140);
and U586 (N_586,N_260,N_434);
nor U587 (N_587,N_65,N_351);
nand U588 (N_588,N_404,N_440);
nand U589 (N_589,N_347,N_345);
or U590 (N_590,N_387,N_319);
nand U591 (N_591,N_133,N_180);
nor U592 (N_592,N_499,N_464);
and U593 (N_593,N_492,N_393);
nand U594 (N_594,N_142,N_448);
and U595 (N_595,N_21,N_369);
or U596 (N_596,N_71,N_1);
nand U597 (N_597,N_324,N_76);
or U598 (N_598,N_240,N_9);
nand U599 (N_599,N_2,N_136);
nor U600 (N_600,N_211,N_216);
nor U601 (N_601,N_171,N_74);
nor U602 (N_602,N_215,N_334);
xor U603 (N_603,N_480,N_412);
or U604 (N_604,N_213,N_362);
and U605 (N_605,N_294,N_406);
or U606 (N_606,N_159,N_281);
or U607 (N_607,N_157,N_8);
xnor U608 (N_608,N_227,N_378);
or U609 (N_609,N_66,N_160);
or U610 (N_610,N_359,N_374);
and U611 (N_611,N_372,N_57);
nor U612 (N_612,N_184,N_415);
nand U613 (N_613,N_188,N_395);
nor U614 (N_614,N_13,N_43);
nor U615 (N_615,N_481,N_20);
nor U616 (N_616,N_259,N_407);
nor U617 (N_617,N_202,N_428);
nor U618 (N_618,N_165,N_418);
or U619 (N_619,N_56,N_386);
nor U620 (N_620,N_250,N_491);
and U621 (N_621,N_145,N_329);
nand U622 (N_622,N_320,N_291);
nand U623 (N_623,N_94,N_328);
nand U624 (N_624,N_295,N_381);
and U625 (N_625,N_420,N_14);
and U626 (N_626,N_49,N_25);
nand U627 (N_627,N_75,N_154);
and U628 (N_628,N_244,N_311);
nor U629 (N_629,N_225,N_286);
nand U630 (N_630,N_128,N_26);
and U631 (N_631,N_78,N_462);
nor U632 (N_632,N_431,N_126);
nand U633 (N_633,N_340,N_151);
nor U634 (N_634,N_61,N_322);
or U635 (N_635,N_490,N_408);
or U636 (N_636,N_179,N_342);
or U637 (N_637,N_0,N_18);
and U638 (N_638,N_371,N_356);
or U639 (N_639,N_245,N_62);
and U640 (N_640,N_40,N_192);
nor U641 (N_641,N_182,N_189);
or U642 (N_642,N_146,N_376);
or U643 (N_643,N_284,N_156);
nand U644 (N_644,N_344,N_141);
nor U645 (N_645,N_451,N_208);
nor U646 (N_646,N_261,N_224);
nand U647 (N_647,N_452,N_425);
and U648 (N_648,N_106,N_314);
xor U649 (N_649,N_200,N_223);
or U650 (N_650,N_365,N_268);
or U651 (N_651,N_99,N_443);
nor U652 (N_652,N_400,N_252);
nor U653 (N_653,N_107,N_468);
nor U654 (N_654,N_486,N_255);
nor U655 (N_655,N_52,N_226);
nand U656 (N_656,N_130,N_274);
nand U657 (N_657,N_233,N_17);
and U658 (N_658,N_300,N_242);
nor U659 (N_659,N_389,N_370);
or U660 (N_660,N_477,N_168);
nor U661 (N_661,N_463,N_231);
and U662 (N_662,N_60,N_249);
or U663 (N_663,N_176,N_91);
nand U664 (N_664,N_147,N_282);
or U665 (N_665,N_465,N_427);
nand U666 (N_666,N_51,N_85);
nor U667 (N_667,N_302,N_429);
nor U668 (N_668,N_305,N_113);
nand U669 (N_669,N_162,N_323);
and U670 (N_670,N_34,N_436);
or U671 (N_671,N_366,N_271);
nand U672 (N_672,N_253,N_361);
or U673 (N_673,N_310,N_398);
or U674 (N_674,N_87,N_273);
nand U675 (N_675,N_276,N_235);
nand U676 (N_676,N_497,N_293);
or U677 (N_677,N_246,N_24);
or U678 (N_678,N_405,N_350);
or U679 (N_679,N_367,N_114);
xor U680 (N_680,N_117,N_445);
nor U681 (N_681,N_360,N_444);
nor U682 (N_682,N_467,N_248);
nor U683 (N_683,N_54,N_270);
nand U684 (N_684,N_336,N_299);
or U685 (N_685,N_265,N_330);
nand U686 (N_686,N_164,N_483);
or U687 (N_687,N_6,N_207);
nor U688 (N_688,N_97,N_290);
nor U689 (N_689,N_186,N_363);
nor U690 (N_690,N_469,N_132);
nor U691 (N_691,N_139,N_37);
nand U692 (N_692,N_471,N_121);
and U693 (N_693,N_22,N_476);
and U694 (N_694,N_120,N_167);
nor U695 (N_695,N_96,N_199);
nor U696 (N_696,N_172,N_69);
nor U697 (N_697,N_105,N_59);
nor U698 (N_698,N_112,N_163);
or U699 (N_699,N_122,N_3);
or U700 (N_700,N_254,N_166);
nor U701 (N_701,N_143,N_384);
and U702 (N_702,N_148,N_209);
nand U703 (N_703,N_401,N_108);
and U704 (N_704,N_161,N_212);
nand U705 (N_705,N_36,N_396);
or U706 (N_706,N_419,N_315);
or U707 (N_707,N_251,N_426);
nor U708 (N_708,N_485,N_123);
nand U709 (N_709,N_446,N_138);
and U710 (N_710,N_496,N_292);
nand U711 (N_711,N_364,N_218);
and U712 (N_712,N_304,N_498);
nor U713 (N_713,N_195,N_234);
nor U714 (N_714,N_441,N_219);
or U715 (N_715,N_183,N_10);
nand U716 (N_716,N_127,N_457);
or U717 (N_717,N_194,N_64);
or U718 (N_718,N_38,N_341);
nor U719 (N_719,N_77,N_439);
or U720 (N_720,N_88,N_262);
and U721 (N_721,N_303,N_423);
nand U722 (N_722,N_236,N_229);
and U723 (N_723,N_430,N_72);
or U724 (N_724,N_449,N_287);
or U725 (N_725,N_470,N_353);
nor U726 (N_726,N_410,N_153);
nor U727 (N_727,N_178,N_27);
and U728 (N_728,N_402,N_23);
nor U729 (N_729,N_474,N_144);
nor U730 (N_730,N_116,N_70);
and U731 (N_731,N_111,N_210);
nor U732 (N_732,N_494,N_19);
nand U733 (N_733,N_306,N_455);
and U734 (N_734,N_413,N_173);
and U735 (N_735,N_190,N_466);
nand U736 (N_736,N_459,N_217);
and U737 (N_737,N_32,N_458);
nand U738 (N_738,N_355,N_403);
or U739 (N_739,N_357,N_119);
nand U740 (N_740,N_33,N_170);
nor U741 (N_741,N_478,N_484);
nor U742 (N_742,N_454,N_45);
nand U743 (N_743,N_44,N_155);
or U744 (N_744,N_63,N_7);
and U745 (N_745,N_447,N_204);
and U746 (N_746,N_41,N_394);
or U747 (N_747,N_332,N_89);
and U748 (N_748,N_438,N_333);
or U749 (N_749,N_135,N_214);
or U750 (N_750,N_409,N_227);
nor U751 (N_751,N_402,N_123);
nor U752 (N_752,N_172,N_432);
nor U753 (N_753,N_313,N_50);
and U754 (N_754,N_108,N_150);
and U755 (N_755,N_338,N_418);
nand U756 (N_756,N_46,N_478);
and U757 (N_757,N_285,N_204);
or U758 (N_758,N_13,N_118);
xnor U759 (N_759,N_243,N_447);
nor U760 (N_760,N_50,N_23);
or U761 (N_761,N_477,N_176);
and U762 (N_762,N_35,N_438);
or U763 (N_763,N_376,N_213);
nand U764 (N_764,N_274,N_198);
nor U765 (N_765,N_161,N_287);
or U766 (N_766,N_307,N_365);
xnor U767 (N_767,N_173,N_322);
xor U768 (N_768,N_363,N_375);
nand U769 (N_769,N_93,N_154);
and U770 (N_770,N_13,N_86);
and U771 (N_771,N_169,N_181);
or U772 (N_772,N_201,N_457);
or U773 (N_773,N_474,N_209);
or U774 (N_774,N_424,N_102);
or U775 (N_775,N_368,N_62);
nor U776 (N_776,N_183,N_268);
or U777 (N_777,N_441,N_33);
and U778 (N_778,N_248,N_245);
nand U779 (N_779,N_111,N_150);
nor U780 (N_780,N_274,N_367);
and U781 (N_781,N_150,N_290);
nor U782 (N_782,N_471,N_377);
and U783 (N_783,N_217,N_494);
or U784 (N_784,N_177,N_466);
or U785 (N_785,N_288,N_141);
and U786 (N_786,N_458,N_392);
nand U787 (N_787,N_386,N_352);
nand U788 (N_788,N_438,N_322);
nand U789 (N_789,N_43,N_423);
nand U790 (N_790,N_410,N_330);
and U791 (N_791,N_410,N_127);
or U792 (N_792,N_474,N_451);
nor U793 (N_793,N_209,N_282);
nor U794 (N_794,N_167,N_408);
nand U795 (N_795,N_303,N_170);
nand U796 (N_796,N_439,N_331);
or U797 (N_797,N_71,N_400);
or U798 (N_798,N_127,N_189);
or U799 (N_799,N_134,N_179);
nand U800 (N_800,N_269,N_229);
nor U801 (N_801,N_489,N_283);
or U802 (N_802,N_287,N_284);
and U803 (N_803,N_245,N_454);
nand U804 (N_804,N_63,N_273);
or U805 (N_805,N_316,N_111);
nand U806 (N_806,N_151,N_494);
and U807 (N_807,N_145,N_110);
nand U808 (N_808,N_195,N_337);
or U809 (N_809,N_362,N_454);
and U810 (N_810,N_254,N_244);
or U811 (N_811,N_252,N_489);
nand U812 (N_812,N_415,N_245);
and U813 (N_813,N_286,N_410);
nor U814 (N_814,N_338,N_120);
or U815 (N_815,N_185,N_41);
or U816 (N_816,N_13,N_29);
or U817 (N_817,N_138,N_313);
or U818 (N_818,N_355,N_407);
nand U819 (N_819,N_459,N_68);
nand U820 (N_820,N_187,N_473);
and U821 (N_821,N_445,N_418);
nand U822 (N_822,N_203,N_454);
nand U823 (N_823,N_314,N_310);
and U824 (N_824,N_84,N_135);
or U825 (N_825,N_463,N_268);
and U826 (N_826,N_344,N_438);
and U827 (N_827,N_228,N_209);
and U828 (N_828,N_482,N_486);
and U829 (N_829,N_117,N_317);
nand U830 (N_830,N_219,N_12);
nand U831 (N_831,N_293,N_149);
xnor U832 (N_832,N_302,N_465);
or U833 (N_833,N_388,N_283);
and U834 (N_834,N_232,N_284);
nand U835 (N_835,N_490,N_94);
or U836 (N_836,N_495,N_265);
nor U837 (N_837,N_481,N_201);
or U838 (N_838,N_161,N_40);
nand U839 (N_839,N_177,N_44);
and U840 (N_840,N_16,N_42);
nand U841 (N_841,N_97,N_169);
and U842 (N_842,N_444,N_491);
nor U843 (N_843,N_406,N_152);
nor U844 (N_844,N_372,N_438);
nor U845 (N_845,N_438,N_29);
nor U846 (N_846,N_143,N_198);
nand U847 (N_847,N_137,N_128);
or U848 (N_848,N_489,N_347);
or U849 (N_849,N_363,N_9);
or U850 (N_850,N_17,N_408);
nor U851 (N_851,N_359,N_279);
nor U852 (N_852,N_119,N_426);
and U853 (N_853,N_316,N_402);
nand U854 (N_854,N_264,N_44);
nand U855 (N_855,N_258,N_381);
and U856 (N_856,N_29,N_41);
or U857 (N_857,N_125,N_290);
nor U858 (N_858,N_249,N_371);
nand U859 (N_859,N_100,N_411);
and U860 (N_860,N_314,N_101);
nand U861 (N_861,N_401,N_383);
nand U862 (N_862,N_310,N_175);
nand U863 (N_863,N_337,N_189);
or U864 (N_864,N_0,N_465);
nor U865 (N_865,N_478,N_123);
or U866 (N_866,N_65,N_78);
nor U867 (N_867,N_42,N_399);
or U868 (N_868,N_277,N_395);
nor U869 (N_869,N_206,N_320);
and U870 (N_870,N_392,N_346);
and U871 (N_871,N_395,N_157);
nand U872 (N_872,N_100,N_245);
and U873 (N_873,N_61,N_444);
xor U874 (N_874,N_301,N_205);
or U875 (N_875,N_386,N_300);
or U876 (N_876,N_187,N_238);
nand U877 (N_877,N_377,N_95);
or U878 (N_878,N_219,N_42);
nand U879 (N_879,N_452,N_319);
nand U880 (N_880,N_124,N_367);
nor U881 (N_881,N_80,N_165);
nand U882 (N_882,N_148,N_104);
nand U883 (N_883,N_6,N_433);
nor U884 (N_884,N_151,N_389);
or U885 (N_885,N_345,N_380);
nand U886 (N_886,N_273,N_19);
and U887 (N_887,N_194,N_150);
nor U888 (N_888,N_47,N_58);
or U889 (N_889,N_398,N_438);
xnor U890 (N_890,N_443,N_174);
or U891 (N_891,N_41,N_9);
or U892 (N_892,N_496,N_217);
nor U893 (N_893,N_64,N_212);
nor U894 (N_894,N_175,N_271);
or U895 (N_895,N_481,N_233);
and U896 (N_896,N_354,N_272);
nor U897 (N_897,N_12,N_161);
or U898 (N_898,N_389,N_100);
or U899 (N_899,N_318,N_174);
and U900 (N_900,N_157,N_463);
and U901 (N_901,N_215,N_261);
nand U902 (N_902,N_498,N_446);
nor U903 (N_903,N_158,N_445);
nand U904 (N_904,N_199,N_309);
and U905 (N_905,N_466,N_406);
or U906 (N_906,N_477,N_161);
nand U907 (N_907,N_163,N_444);
and U908 (N_908,N_432,N_371);
and U909 (N_909,N_47,N_107);
nand U910 (N_910,N_454,N_321);
and U911 (N_911,N_74,N_469);
and U912 (N_912,N_27,N_453);
or U913 (N_913,N_378,N_261);
nand U914 (N_914,N_165,N_495);
nor U915 (N_915,N_340,N_184);
or U916 (N_916,N_477,N_58);
and U917 (N_917,N_230,N_347);
or U918 (N_918,N_155,N_418);
nor U919 (N_919,N_445,N_453);
and U920 (N_920,N_172,N_56);
or U921 (N_921,N_334,N_186);
or U922 (N_922,N_431,N_397);
nor U923 (N_923,N_245,N_133);
nand U924 (N_924,N_233,N_456);
or U925 (N_925,N_106,N_470);
nand U926 (N_926,N_323,N_496);
and U927 (N_927,N_293,N_211);
xnor U928 (N_928,N_99,N_16);
xor U929 (N_929,N_256,N_343);
and U930 (N_930,N_384,N_18);
nor U931 (N_931,N_310,N_492);
nand U932 (N_932,N_141,N_401);
nand U933 (N_933,N_13,N_205);
nand U934 (N_934,N_415,N_129);
nor U935 (N_935,N_231,N_125);
nor U936 (N_936,N_230,N_444);
or U937 (N_937,N_420,N_244);
nand U938 (N_938,N_235,N_49);
and U939 (N_939,N_460,N_88);
nand U940 (N_940,N_72,N_184);
nor U941 (N_941,N_490,N_119);
nand U942 (N_942,N_24,N_128);
xnor U943 (N_943,N_434,N_331);
nor U944 (N_944,N_312,N_264);
nor U945 (N_945,N_496,N_472);
or U946 (N_946,N_234,N_370);
or U947 (N_947,N_447,N_1);
nor U948 (N_948,N_436,N_328);
and U949 (N_949,N_14,N_248);
and U950 (N_950,N_246,N_235);
nand U951 (N_951,N_365,N_350);
nand U952 (N_952,N_56,N_325);
nor U953 (N_953,N_43,N_263);
nor U954 (N_954,N_191,N_208);
nor U955 (N_955,N_196,N_38);
nor U956 (N_956,N_137,N_28);
nor U957 (N_957,N_425,N_98);
nor U958 (N_958,N_213,N_430);
and U959 (N_959,N_299,N_349);
nand U960 (N_960,N_306,N_434);
or U961 (N_961,N_82,N_68);
nand U962 (N_962,N_241,N_372);
or U963 (N_963,N_11,N_332);
nor U964 (N_964,N_31,N_70);
nand U965 (N_965,N_29,N_97);
nor U966 (N_966,N_41,N_174);
or U967 (N_967,N_65,N_267);
or U968 (N_968,N_273,N_179);
or U969 (N_969,N_412,N_474);
nor U970 (N_970,N_306,N_420);
and U971 (N_971,N_311,N_73);
or U972 (N_972,N_175,N_217);
nor U973 (N_973,N_409,N_97);
or U974 (N_974,N_371,N_324);
nand U975 (N_975,N_147,N_447);
nor U976 (N_976,N_456,N_38);
nor U977 (N_977,N_46,N_325);
nand U978 (N_978,N_5,N_283);
or U979 (N_979,N_184,N_417);
and U980 (N_980,N_380,N_234);
xnor U981 (N_981,N_6,N_232);
nand U982 (N_982,N_173,N_4);
nand U983 (N_983,N_363,N_397);
or U984 (N_984,N_110,N_499);
and U985 (N_985,N_428,N_360);
nand U986 (N_986,N_11,N_237);
nor U987 (N_987,N_315,N_493);
or U988 (N_988,N_184,N_275);
nand U989 (N_989,N_427,N_485);
and U990 (N_990,N_29,N_50);
or U991 (N_991,N_53,N_369);
nor U992 (N_992,N_20,N_369);
nand U993 (N_993,N_195,N_435);
nor U994 (N_994,N_443,N_472);
nand U995 (N_995,N_252,N_49);
or U996 (N_996,N_129,N_317);
and U997 (N_997,N_0,N_176);
and U998 (N_998,N_400,N_456);
nor U999 (N_999,N_296,N_81);
and U1000 (N_1000,N_877,N_929);
nor U1001 (N_1001,N_660,N_831);
nor U1002 (N_1002,N_849,N_815);
or U1003 (N_1003,N_691,N_694);
nor U1004 (N_1004,N_595,N_969);
nor U1005 (N_1005,N_986,N_973);
nand U1006 (N_1006,N_822,N_914);
nand U1007 (N_1007,N_601,N_571);
nand U1008 (N_1008,N_897,N_912);
and U1009 (N_1009,N_667,N_866);
nor U1010 (N_1010,N_952,N_880);
and U1011 (N_1011,N_656,N_616);
and U1012 (N_1012,N_637,N_670);
and U1013 (N_1013,N_545,N_547);
nand U1014 (N_1014,N_573,N_847);
nand U1015 (N_1015,N_625,N_920);
nor U1016 (N_1016,N_610,N_928);
or U1017 (N_1017,N_874,N_621);
nand U1018 (N_1018,N_555,N_622);
nand U1019 (N_1019,N_664,N_905);
xnor U1020 (N_1020,N_825,N_592);
or U1021 (N_1021,N_565,N_506);
and U1022 (N_1022,N_716,N_774);
or U1023 (N_1023,N_628,N_553);
nor U1024 (N_1024,N_557,N_517);
nand U1025 (N_1025,N_665,N_518);
or U1026 (N_1026,N_927,N_567);
and U1027 (N_1027,N_881,N_712);
and U1028 (N_1028,N_790,N_587);
and U1029 (N_1029,N_735,N_942);
nand U1030 (N_1030,N_793,N_629);
and U1031 (N_1031,N_870,N_540);
nand U1032 (N_1032,N_875,N_584);
or U1033 (N_1033,N_820,N_839);
and U1034 (N_1034,N_908,N_792);
nand U1035 (N_1035,N_998,N_980);
nor U1036 (N_1036,N_626,N_674);
nor U1037 (N_1037,N_562,N_534);
and U1038 (N_1038,N_802,N_583);
or U1039 (N_1039,N_701,N_549);
nand U1040 (N_1040,N_860,N_863);
and U1041 (N_1041,N_844,N_972);
or U1042 (N_1042,N_685,N_639);
nand U1043 (N_1043,N_641,N_703);
nor U1044 (N_1044,N_541,N_684);
and U1045 (N_1045,N_807,N_865);
or U1046 (N_1046,N_732,N_982);
and U1047 (N_1047,N_538,N_892);
or U1048 (N_1048,N_653,N_556);
nor U1049 (N_1049,N_944,N_711);
xnor U1050 (N_1050,N_672,N_924);
nor U1051 (N_1051,N_605,N_819);
nor U1052 (N_1052,N_948,N_967);
or U1053 (N_1053,N_649,N_683);
nand U1054 (N_1054,N_657,N_604);
nand U1055 (N_1055,N_654,N_662);
nor U1056 (N_1056,N_658,N_544);
nand U1057 (N_1057,N_514,N_718);
or U1058 (N_1058,N_725,N_743);
and U1059 (N_1059,N_976,N_795);
nor U1060 (N_1060,N_835,N_834);
nor U1061 (N_1061,N_681,N_650);
nor U1062 (N_1062,N_569,N_526);
and U1063 (N_1063,N_776,N_975);
nor U1064 (N_1064,N_726,N_669);
or U1065 (N_1065,N_615,N_960);
and U1066 (N_1066,N_894,N_964);
or U1067 (N_1067,N_590,N_559);
nor U1068 (N_1068,N_680,N_821);
or U1069 (N_1069,N_891,N_777);
and U1070 (N_1070,N_833,N_501);
or U1071 (N_1071,N_539,N_933);
and U1072 (N_1072,N_823,N_751);
and U1073 (N_1073,N_581,N_682);
and U1074 (N_1074,N_638,N_676);
xor U1075 (N_1075,N_773,N_558);
nor U1076 (N_1076,N_500,N_560);
nand U1077 (N_1077,N_736,N_748);
nor U1078 (N_1078,N_630,N_935);
and U1079 (N_1079,N_546,N_698);
nor U1080 (N_1080,N_926,N_572);
nand U1081 (N_1081,N_537,N_826);
and U1082 (N_1082,N_745,N_661);
and U1083 (N_1083,N_854,N_603);
and U1084 (N_1084,N_754,N_841);
nor U1085 (N_1085,N_634,N_575);
and U1086 (N_1086,N_886,N_542);
nand U1087 (N_1087,N_524,N_800);
nor U1088 (N_1088,N_678,N_806);
nor U1089 (N_1089,N_871,N_989);
and U1090 (N_1090,N_692,N_919);
nor U1091 (N_1091,N_816,N_809);
and U1092 (N_1092,N_940,N_530);
and U1093 (N_1093,N_668,N_607);
and U1094 (N_1094,N_750,N_963);
nand U1095 (N_1095,N_861,N_786);
and U1096 (N_1096,N_582,N_700);
or U1097 (N_1097,N_591,N_686);
nor U1098 (N_1098,N_999,N_580);
and U1099 (N_1099,N_768,N_752);
and U1100 (N_1100,N_784,N_695);
and U1101 (N_1101,N_824,N_838);
nand U1102 (N_1102,N_810,N_900);
and U1103 (N_1103,N_859,N_857);
or U1104 (N_1104,N_663,N_950);
nor U1105 (N_1105,N_715,N_708);
nand U1106 (N_1106,N_554,N_947);
and U1107 (N_1107,N_906,N_814);
and U1108 (N_1108,N_525,N_510);
or U1109 (N_1109,N_992,N_991);
nand U1110 (N_1110,N_799,N_643);
nor U1111 (N_1111,N_923,N_535);
nand U1112 (N_1112,N_953,N_761);
or U1113 (N_1113,N_756,N_570);
or U1114 (N_1114,N_918,N_758);
or U1115 (N_1115,N_852,N_746);
nor U1116 (N_1116,N_842,N_652);
nor U1117 (N_1117,N_713,N_946);
and U1118 (N_1118,N_853,N_830);
and U1119 (N_1119,N_627,N_803);
nor U1120 (N_1120,N_633,N_785);
or U1121 (N_1121,N_913,N_837);
nand U1122 (N_1122,N_832,N_878);
xor U1123 (N_1123,N_829,N_943);
or U1124 (N_1124,N_791,N_568);
nand U1125 (N_1125,N_721,N_965);
or U1126 (N_1126,N_884,N_640);
and U1127 (N_1127,N_551,N_729);
or U1128 (N_1128,N_614,N_879);
nand U1129 (N_1129,N_783,N_597);
nand U1130 (N_1130,N_818,N_593);
nand U1131 (N_1131,N_966,N_995);
nand U1132 (N_1132,N_850,N_902);
and U1133 (N_1133,N_502,N_996);
nor U1134 (N_1134,N_903,N_753);
or U1135 (N_1135,N_997,N_951);
or U1136 (N_1136,N_895,N_659);
nor U1137 (N_1137,N_949,N_782);
nor U1138 (N_1138,N_688,N_731);
and U1139 (N_1139,N_631,N_671);
or U1140 (N_1140,N_781,N_666);
nand U1141 (N_1141,N_848,N_939);
nor U1142 (N_1142,N_599,N_981);
or U1143 (N_1143,N_805,N_747);
or U1144 (N_1144,N_602,N_936);
and U1145 (N_1145,N_620,N_520);
and U1146 (N_1146,N_767,N_503);
and U1147 (N_1147,N_741,N_617);
nand U1148 (N_1148,N_679,N_749);
nor U1149 (N_1149,N_907,N_606);
nor U1150 (N_1150,N_722,N_734);
nor U1151 (N_1151,N_646,N_772);
or U1152 (N_1152,N_724,N_521);
nand U1153 (N_1153,N_970,N_873);
or U1154 (N_1154,N_985,N_794);
and U1155 (N_1155,N_704,N_858);
nand U1156 (N_1156,N_645,N_613);
and U1157 (N_1157,N_862,N_804);
xnor U1158 (N_1158,N_687,N_706);
or U1159 (N_1159,N_779,N_608);
xnor U1160 (N_1160,N_910,N_532);
nand U1161 (N_1161,N_988,N_707);
and U1162 (N_1162,N_762,N_720);
and U1163 (N_1163,N_959,N_840);
or U1164 (N_1164,N_755,N_978);
nand U1165 (N_1165,N_778,N_527);
nand U1166 (N_1166,N_655,N_697);
or U1167 (N_1167,N_589,N_522);
or U1168 (N_1168,N_536,N_788);
and U1169 (N_1169,N_512,N_808);
or U1170 (N_1170,N_930,N_885);
and U1171 (N_1171,N_618,N_586);
nor U1172 (N_1172,N_856,N_699);
nand U1173 (N_1173,N_651,N_760);
or U1174 (N_1174,N_855,N_742);
nor U1175 (N_1175,N_515,N_528);
nand U1176 (N_1176,N_828,N_994);
or U1177 (N_1177,N_775,N_909);
or U1178 (N_1178,N_677,N_596);
or U1179 (N_1179,N_843,N_705);
nor U1180 (N_1180,N_673,N_796);
and U1181 (N_1181,N_696,N_588);
and U1182 (N_1182,N_780,N_766);
nand U1183 (N_1183,N_898,N_813);
nand U1184 (N_1184,N_938,N_611);
or U1185 (N_1185,N_523,N_714);
or U1186 (N_1186,N_872,N_513);
and U1187 (N_1187,N_709,N_609);
and U1188 (N_1188,N_723,N_578);
nand U1189 (N_1189,N_864,N_974);
or U1190 (N_1190,N_632,N_757);
nor U1191 (N_1191,N_797,N_533);
or U1192 (N_1192,N_925,N_954);
nor U1193 (N_1193,N_941,N_916);
nand U1194 (N_1194,N_911,N_543);
nor U1195 (N_1195,N_765,N_993);
nor U1196 (N_1196,N_576,N_509);
xor U1197 (N_1197,N_977,N_812);
nor U1198 (N_1198,N_636,N_883);
and U1199 (N_1199,N_887,N_644);
or U1200 (N_1200,N_612,N_552);
and U1201 (N_1201,N_717,N_531);
and U1202 (N_1202,N_739,N_827);
or U1203 (N_1203,N_851,N_769);
and U1204 (N_1204,N_845,N_594);
nand U1205 (N_1205,N_579,N_876);
nor U1206 (N_1206,N_508,N_624);
and U1207 (N_1207,N_869,N_727);
nand U1208 (N_1208,N_836,N_899);
nor U1209 (N_1209,N_619,N_738);
nor U1210 (N_1210,N_600,N_574);
or U1211 (N_1211,N_817,N_759);
nand U1212 (N_1212,N_962,N_566);
and U1213 (N_1213,N_693,N_561);
nor U1214 (N_1214,N_957,N_955);
nor U1215 (N_1215,N_867,N_719);
and U1216 (N_1216,N_598,N_901);
xor U1217 (N_1217,N_789,N_889);
or U1218 (N_1218,N_648,N_763);
nor U1219 (N_1219,N_519,N_917);
nand U1220 (N_1220,N_744,N_529);
nand U1221 (N_1221,N_915,N_798);
or U1222 (N_1222,N_956,N_548);
and U1223 (N_1223,N_507,N_968);
nand U1224 (N_1224,N_893,N_888);
and U1225 (N_1225,N_505,N_764);
and U1226 (N_1226,N_922,N_971);
or U1227 (N_1227,N_730,N_932);
xor U1228 (N_1228,N_771,N_737);
xnor U1229 (N_1229,N_983,N_563);
or U1230 (N_1230,N_934,N_623);
nand U1231 (N_1231,N_511,N_504);
and U1232 (N_1232,N_728,N_516);
nor U1233 (N_1233,N_937,N_890);
nand U1234 (N_1234,N_577,N_787);
nand U1235 (N_1235,N_882,N_958);
and U1236 (N_1236,N_990,N_961);
nand U1237 (N_1237,N_690,N_846);
and U1238 (N_1238,N_733,N_740);
and U1239 (N_1239,N_689,N_675);
or U1240 (N_1240,N_564,N_868);
nor U1241 (N_1241,N_987,N_801);
nor U1242 (N_1242,N_896,N_702);
or U1243 (N_1243,N_635,N_770);
nand U1244 (N_1244,N_642,N_904);
nor U1245 (N_1245,N_550,N_710);
nor U1246 (N_1246,N_984,N_585);
and U1247 (N_1247,N_945,N_979);
and U1248 (N_1248,N_811,N_931);
nand U1249 (N_1249,N_921,N_647);
or U1250 (N_1250,N_966,N_740);
nor U1251 (N_1251,N_560,N_998);
and U1252 (N_1252,N_734,N_579);
nor U1253 (N_1253,N_930,N_566);
and U1254 (N_1254,N_949,N_629);
and U1255 (N_1255,N_830,N_763);
nor U1256 (N_1256,N_685,N_647);
or U1257 (N_1257,N_779,N_973);
xnor U1258 (N_1258,N_629,N_603);
nand U1259 (N_1259,N_662,N_919);
and U1260 (N_1260,N_550,N_840);
nand U1261 (N_1261,N_551,N_563);
nor U1262 (N_1262,N_820,N_829);
nand U1263 (N_1263,N_843,N_525);
nor U1264 (N_1264,N_606,N_585);
nor U1265 (N_1265,N_877,N_656);
or U1266 (N_1266,N_902,N_572);
nor U1267 (N_1267,N_816,N_616);
nor U1268 (N_1268,N_830,N_575);
nand U1269 (N_1269,N_515,N_507);
nor U1270 (N_1270,N_712,N_844);
or U1271 (N_1271,N_920,N_900);
and U1272 (N_1272,N_752,N_774);
and U1273 (N_1273,N_729,N_542);
or U1274 (N_1274,N_949,N_952);
or U1275 (N_1275,N_927,N_760);
xor U1276 (N_1276,N_694,N_617);
nor U1277 (N_1277,N_561,N_515);
and U1278 (N_1278,N_927,N_908);
and U1279 (N_1279,N_871,N_949);
nor U1280 (N_1280,N_814,N_868);
and U1281 (N_1281,N_639,N_895);
xor U1282 (N_1282,N_656,N_849);
nand U1283 (N_1283,N_678,N_916);
or U1284 (N_1284,N_816,N_556);
or U1285 (N_1285,N_811,N_793);
or U1286 (N_1286,N_759,N_930);
nand U1287 (N_1287,N_833,N_942);
and U1288 (N_1288,N_783,N_696);
and U1289 (N_1289,N_955,N_981);
nand U1290 (N_1290,N_501,N_566);
or U1291 (N_1291,N_802,N_862);
nor U1292 (N_1292,N_967,N_938);
nand U1293 (N_1293,N_754,N_775);
nor U1294 (N_1294,N_641,N_841);
nand U1295 (N_1295,N_842,N_853);
and U1296 (N_1296,N_938,N_989);
and U1297 (N_1297,N_755,N_656);
and U1298 (N_1298,N_954,N_997);
nor U1299 (N_1299,N_651,N_525);
or U1300 (N_1300,N_787,N_782);
and U1301 (N_1301,N_885,N_621);
nor U1302 (N_1302,N_589,N_811);
nand U1303 (N_1303,N_636,N_843);
nor U1304 (N_1304,N_793,N_553);
nor U1305 (N_1305,N_983,N_871);
or U1306 (N_1306,N_992,N_654);
nor U1307 (N_1307,N_930,N_988);
or U1308 (N_1308,N_761,N_695);
and U1309 (N_1309,N_862,N_666);
nor U1310 (N_1310,N_682,N_697);
or U1311 (N_1311,N_616,N_626);
nor U1312 (N_1312,N_582,N_807);
and U1313 (N_1313,N_826,N_878);
nor U1314 (N_1314,N_892,N_694);
nand U1315 (N_1315,N_900,N_817);
or U1316 (N_1316,N_852,N_809);
nand U1317 (N_1317,N_947,N_898);
and U1318 (N_1318,N_549,N_839);
and U1319 (N_1319,N_881,N_735);
xnor U1320 (N_1320,N_974,N_525);
xnor U1321 (N_1321,N_670,N_543);
and U1322 (N_1322,N_982,N_678);
and U1323 (N_1323,N_785,N_703);
and U1324 (N_1324,N_520,N_789);
nor U1325 (N_1325,N_525,N_647);
or U1326 (N_1326,N_782,N_956);
or U1327 (N_1327,N_957,N_858);
or U1328 (N_1328,N_540,N_696);
or U1329 (N_1329,N_619,N_880);
nor U1330 (N_1330,N_570,N_924);
or U1331 (N_1331,N_657,N_711);
nor U1332 (N_1332,N_965,N_843);
or U1333 (N_1333,N_748,N_663);
nor U1334 (N_1334,N_882,N_995);
or U1335 (N_1335,N_995,N_998);
nor U1336 (N_1336,N_905,N_507);
nor U1337 (N_1337,N_836,N_988);
or U1338 (N_1338,N_520,N_805);
nand U1339 (N_1339,N_776,N_711);
nand U1340 (N_1340,N_856,N_796);
nand U1341 (N_1341,N_598,N_811);
nor U1342 (N_1342,N_744,N_599);
nor U1343 (N_1343,N_763,N_839);
nor U1344 (N_1344,N_779,N_535);
nor U1345 (N_1345,N_959,N_967);
nand U1346 (N_1346,N_555,N_583);
nand U1347 (N_1347,N_651,N_913);
and U1348 (N_1348,N_723,N_855);
or U1349 (N_1349,N_956,N_591);
and U1350 (N_1350,N_702,N_837);
and U1351 (N_1351,N_649,N_713);
or U1352 (N_1352,N_728,N_781);
nand U1353 (N_1353,N_934,N_614);
nor U1354 (N_1354,N_617,N_827);
and U1355 (N_1355,N_800,N_709);
and U1356 (N_1356,N_688,N_934);
or U1357 (N_1357,N_731,N_681);
nand U1358 (N_1358,N_567,N_879);
or U1359 (N_1359,N_912,N_928);
nor U1360 (N_1360,N_838,N_538);
or U1361 (N_1361,N_880,N_631);
nor U1362 (N_1362,N_563,N_896);
or U1363 (N_1363,N_811,N_918);
and U1364 (N_1364,N_971,N_751);
nand U1365 (N_1365,N_885,N_943);
or U1366 (N_1366,N_992,N_552);
and U1367 (N_1367,N_549,N_996);
and U1368 (N_1368,N_504,N_648);
nor U1369 (N_1369,N_821,N_695);
and U1370 (N_1370,N_692,N_894);
nand U1371 (N_1371,N_939,N_870);
and U1372 (N_1372,N_694,N_510);
nor U1373 (N_1373,N_616,N_921);
nor U1374 (N_1374,N_779,N_669);
or U1375 (N_1375,N_676,N_822);
nand U1376 (N_1376,N_881,N_931);
nor U1377 (N_1377,N_808,N_752);
nor U1378 (N_1378,N_513,N_898);
nor U1379 (N_1379,N_516,N_885);
nand U1380 (N_1380,N_967,N_889);
and U1381 (N_1381,N_790,N_970);
nand U1382 (N_1382,N_727,N_563);
nor U1383 (N_1383,N_611,N_511);
nor U1384 (N_1384,N_939,N_608);
or U1385 (N_1385,N_526,N_933);
or U1386 (N_1386,N_889,N_924);
nor U1387 (N_1387,N_863,N_889);
nand U1388 (N_1388,N_858,N_801);
and U1389 (N_1389,N_664,N_665);
and U1390 (N_1390,N_579,N_877);
and U1391 (N_1391,N_819,N_587);
nor U1392 (N_1392,N_539,N_789);
or U1393 (N_1393,N_965,N_783);
and U1394 (N_1394,N_685,N_577);
and U1395 (N_1395,N_988,N_947);
and U1396 (N_1396,N_516,N_968);
nand U1397 (N_1397,N_757,N_532);
and U1398 (N_1398,N_876,N_606);
nand U1399 (N_1399,N_618,N_812);
and U1400 (N_1400,N_864,N_801);
nand U1401 (N_1401,N_605,N_833);
nor U1402 (N_1402,N_621,N_512);
and U1403 (N_1403,N_566,N_923);
and U1404 (N_1404,N_730,N_672);
nand U1405 (N_1405,N_991,N_611);
nor U1406 (N_1406,N_515,N_818);
and U1407 (N_1407,N_755,N_961);
or U1408 (N_1408,N_767,N_964);
and U1409 (N_1409,N_629,N_620);
nand U1410 (N_1410,N_933,N_741);
or U1411 (N_1411,N_625,N_898);
nor U1412 (N_1412,N_891,N_867);
or U1413 (N_1413,N_826,N_988);
and U1414 (N_1414,N_860,N_918);
nor U1415 (N_1415,N_763,N_557);
nand U1416 (N_1416,N_730,N_972);
nor U1417 (N_1417,N_599,N_886);
or U1418 (N_1418,N_945,N_704);
nor U1419 (N_1419,N_697,N_657);
nor U1420 (N_1420,N_849,N_555);
and U1421 (N_1421,N_812,N_579);
and U1422 (N_1422,N_639,N_665);
and U1423 (N_1423,N_823,N_621);
nand U1424 (N_1424,N_883,N_935);
or U1425 (N_1425,N_748,N_976);
nor U1426 (N_1426,N_842,N_958);
nand U1427 (N_1427,N_765,N_922);
nor U1428 (N_1428,N_856,N_878);
nand U1429 (N_1429,N_994,N_524);
nand U1430 (N_1430,N_978,N_614);
or U1431 (N_1431,N_807,N_975);
nor U1432 (N_1432,N_670,N_617);
nand U1433 (N_1433,N_588,N_932);
nand U1434 (N_1434,N_734,N_968);
and U1435 (N_1435,N_828,N_734);
nor U1436 (N_1436,N_893,N_755);
and U1437 (N_1437,N_527,N_669);
or U1438 (N_1438,N_925,N_911);
nor U1439 (N_1439,N_655,N_918);
nand U1440 (N_1440,N_529,N_541);
nor U1441 (N_1441,N_933,N_723);
and U1442 (N_1442,N_528,N_612);
nor U1443 (N_1443,N_666,N_948);
nand U1444 (N_1444,N_917,N_848);
or U1445 (N_1445,N_510,N_820);
and U1446 (N_1446,N_841,N_521);
and U1447 (N_1447,N_529,N_829);
and U1448 (N_1448,N_717,N_625);
nand U1449 (N_1449,N_646,N_635);
or U1450 (N_1450,N_959,N_817);
or U1451 (N_1451,N_692,N_763);
nor U1452 (N_1452,N_674,N_727);
and U1453 (N_1453,N_531,N_744);
and U1454 (N_1454,N_991,N_569);
or U1455 (N_1455,N_711,N_671);
or U1456 (N_1456,N_781,N_853);
xor U1457 (N_1457,N_961,N_571);
nor U1458 (N_1458,N_712,N_636);
and U1459 (N_1459,N_928,N_669);
nand U1460 (N_1460,N_934,N_567);
nor U1461 (N_1461,N_536,N_640);
nor U1462 (N_1462,N_829,N_860);
and U1463 (N_1463,N_876,N_668);
nor U1464 (N_1464,N_938,N_613);
nand U1465 (N_1465,N_570,N_824);
and U1466 (N_1466,N_638,N_762);
xnor U1467 (N_1467,N_753,N_938);
nand U1468 (N_1468,N_624,N_807);
nor U1469 (N_1469,N_636,N_935);
and U1470 (N_1470,N_813,N_591);
nor U1471 (N_1471,N_993,N_709);
or U1472 (N_1472,N_735,N_552);
or U1473 (N_1473,N_655,N_837);
or U1474 (N_1474,N_835,N_758);
and U1475 (N_1475,N_818,N_836);
or U1476 (N_1476,N_778,N_959);
nor U1477 (N_1477,N_684,N_799);
nand U1478 (N_1478,N_623,N_827);
or U1479 (N_1479,N_713,N_997);
nand U1480 (N_1480,N_711,N_862);
nand U1481 (N_1481,N_651,N_748);
nor U1482 (N_1482,N_567,N_658);
nand U1483 (N_1483,N_515,N_885);
nor U1484 (N_1484,N_823,N_645);
and U1485 (N_1485,N_695,N_610);
nand U1486 (N_1486,N_845,N_751);
and U1487 (N_1487,N_631,N_579);
nor U1488 (N_1488,N_657,N_737);
or U1489 (N_1489,N_581,N_731);
nand U1490 (N_1490,N_610,N_615);
nor U1491 (N_1491,N_781,N_928);
nand U1492 (N_1492,N_624,N_902);
or U1493 (N_1493,N_812,N_793);
and U1494 (N_1494,N_540,N_615);
or U1495 (N_1495,N_843,N_546);
and U1496 (N_1496,N_775,N_732);
nor U1497 (N_1497,N_793,N_562);
or U1498 (N_1498,N_945,N_563);
nand U1499 (N_1499,N_514,N_990);
nand U1500 (N_1500,N_1125,N_1260);
nand U1501 (N_1501,N_1352,N_1332);
nor U1502 (N_1502,N_1297,N_1002);
and U1503 (N_1503,N_1448,N_1270);
and U1504 (N_1504,N_1320,N_1254);
or U1505 (N_1505,N_1455,N_1167);
and U1506 (N_1506,N_1075,N_1006);
and U1507 (N_1507,N_1113,N_1216);
nor U1508 (N_1508,N_1308,N_1048);
xnor U1509 (N_1509,N_1283,N_1482);
and U1510 (N_1510,N_1192,N_1400);
nand U1511 (N_1511,N_1305,N_1007);
nor U1512 (N_1512,N_1241,N_1279);
and U1513 (N_1513,N_1151,N_1214);
or U1514 (N_1514,N_1295,N_1128);
nor U1515 (N_1515,N_1474,N_1083);
nor U1516 (N_1516,N_1120,N_1028);
xnor U1517 (N_1517,N_1029,N_1406);
nand U1518 (N_1518,N_1430,N_1424);
nand U1519 (N_1519,N_1186,N_1240);
and U1520 (N_1520,N_1379,N_1336);
and U1521 (N_1521,N_1215,N_1107);
nand U1522 (N_1522,N_1287,N_1203);
or U1523 (N_1523,N_1257,N_1184);
nor U1524 (N_1524,N_1047,N_1087);
nor U1525 (N_1525,N_1431,N_1085);
nand U1526 (N_1526,N_1372,N_1210);
nor U1527 (N_1527,N_1014,N_1217);
and U1528 (N_1528,N_1414,N_1088);
nand U1529 (N_1529,N_1312,N_1326);
nand U1530 (N_1530,N_1017,N_1265);
nor U1531 (N_1531,N_1137,N_1280);
nor U1532 (N_1532,N_1288,N_1110);
nand U1533 (N_1533,N_1416,N_1053);
nor U1534 (N_1534,N_1129,N_1324);
nor U1535 (N_1535,N_1469,N_1180);
nand U1536 (N_1536,N_1080,N_1106);
nand U1537 (N_1537,N_1383,N_1093);
nor U1538 (N_1538,N_1481,N_1237);
nor U1539 (N_1539,N_1378,N_1025);
nor U1540 (N_1540,N_1425,N_1489);
or U1541 (N_1541,N_1174,N_1330);
and U1542 (N_1542,N_1057,N_1452);
or U1543 (N_1543,N_1478,N_1247);
or U1544 (N_1544,N_1496,N_1126);
or U1545 (N_1545,N_1109,N_1323);
nor U1546 (N_1546,N_1438,N_1294);
and U1547 (N_1547,N_1197,N_1401);
and U1548 (N_1548,N_1410,N_1321);
and U1549 (N_1549,N_1310,N_1419);
nand U1550 (N_1550,N_1204,N_1169);
or U1551 (N_1551,N_1069,N_1050);
and U1552 (N_1552,N_1233,N_1255);
nand U1553 (N_1553,N_1470,N_1038);
nor U1554 (N_1554,N_1189,N_1380);
or U1555 (N_1555,N_1355,N_1181);
or U1556 (N_1556,N_1223,N_1395);
nand U1557 (N_1557,N_1155,N_1306);
or U1558 (N_1558,N_1150,N_1117);
nand U1559 (N_1559,N_1396,N_1073);
nor U1560 (N_1560,N_1039,N_1060);
and U1561 (N_1561,N_1008,N_1198);
xor U1562 (N_1562,N_1300,N_1256);
nand U1563 (N_1563,N_1461,N_1315);
nor U1564 (N_1564,N_1079,N_1421);
nor U1565 (N_1565,N_1072,N_1345);
or U1566 (N_1566,N_1480,N_1148);
nand U1567 (N_1567,N_1479,N_1331);
nor U1568 (N_1568,N_1052,N_1175);
nor U1569 (N_1569,N_1230,N_1092);
nand U1570 (N_1570,N_1311,N_1018);
nor U1571 (N_1571,N_1056,N_1076);
nand U1572 (N_1572,N_1468,N_1339);
nand U1573 (N_1573,N_1037,N_1358);
nor U1574 (N_1574,N_1211,N_1281);
nand U1575 (N_1575,N_1170,N_1182);
nand U1576 (N_1576,N_1185,N_1365);
nand U1577 (N_1577,N_1201,N_1134);
or U1578 (N_1578,N_1229,N_1033);
or U1579 (N_1579,N_1232,N_1221);
and U1580 (N_1580,N_1023,N_1141);
and U1581 (N_1581,N_1486,N_1423);
and U1582 (N_1582,N_1194,N_1413);
nor U1583 (N_1583,N_1245,N_1154);
nand U1584 (N_1584,N_1304,N_1451);
xor U1585 (N_1585,N_1160,N_1034);
nor U1586 (N_1586,N_1049,N_1462);
or U1587 (N_1587,N_1271,N_1450);
nor U1588 (N_1588,N_1131,N_1449);
xor U1589 (N_1589,N_1407,N_1477);
nor U1590 (N_1590,N_1382,N_1368);
nand U1591 (N_1591,N_1001,N_1004);
nor U1592 (N_1592,N_1444,N_1231);
or U1593 (N_1593,N_1242,N_1374);
and U1594 (N_1594,N_1114,N_1096);
or U1595 (N_1595,N_1021,N_1065);
and U1596 (N_1596,N_1370,N_1173);
or U1597 (N_1597,N_1317,N_1222);
and U1598 (N_1598,N_1176,N_1139);
or U1599 (N_1599,N_1082,N_1354);
nand U1600 (N_1600,N_1152,N_1149);
or U1601 (N_1601,N_1268,N_1492);
and U1602 (N_1602,N_1435,N_1196);
nand U1603 (N_1603,N_1070,N_1301);
and U1604 (N_1604,N_1328,N_1195);
or U1605 (N_1605,N_1224,N_1341);
and U1606 (N_1606,N_1101,N_1097);
and U1607 (N_1607,N_1136,N_1031);
or U1608 (N_1608,N_1393,N_1409);
and U1609 (N_1609,N_1377,N_1010);
nor U1610 (N_1610,N_1307,N_1135);
or U1611 (N_1611,N_1266,N_1103);
nor U1612 (N_1612,N_1293,N_1043);
nand U1613 (N_1613,N_1228,N_1249);
nand U1614 (N_1614,N_1188,N_1165);
or U1615 (N_1615,N_1439,N_1239);
nor U1616 (N_1616,N_1346,N_1394);
nor U1617 (N_1617,N_1334,N_1145);
or U1618 (N_1618,N_1497,N_1289);
nand U1619 (N_1619,N_1115,N_1402);
or U1620 (N_1620,N_1314,N_1178);
nand U1621 (N_1621,N_1344,N_1303);
nor U1622 (N_1622,N_1420,N_1463);
nor U1623 (N_1623,N_1251,N_1313);
nand U1624 (N_1624,N_1363,N_1142);
or U1625 (N_1625,N_1465,N_1153);
nand U1626 (N_1626,N_1278,N_1191);
or U1627 (N_1627,N_1291,N_1360);
nand U1628 (N_1628,N_1389,N_1022);
or U1629 (N_1629,N_1200,N_1207);
or U1630 (N_1630,N_1030,N_1067);
nand U1631 (N_1631,N_1099,N_1364);
or U1632 (N_1632,N_1162,N_1166);
nand U1633 (N_1633,N_1071,N_1081);
xor U1634 (N_1634,N_1219,N_1243);
and U1635 (N_1635,N_1392,N_1027);
and U1636 (N_1636,N_1375,N_1227);
or U1637 (N_1637,N_1246,N_1164);
nor U1638 (N_1638,N_1285,N_1112);
and U1639 (N_1639,N_1422,N_1074);
nand U1640 (N_1640,N_1456,N_1353);
nand U1641 (N_1641,N_1398,N_1090);
nand U1642 (N_1642,N_1473,N_1108);
nor U1643 (N_1643,N_1493,N_1272);
nand U1644 (N_1644,N_1361,N_1498);
or U1645 (N_1645,N_1138,N_1284);
nor U1646 (N_1646,N_1475,N_1124);
nor U1647 (N_1647,N_1397,N_1411);
xor U1648 (N_1648,N_1019,N_1143);
nand U1649 (N_1649,N_1376,N_1467);
and U1650 (N_1650,N_1459,N_1051);
nor U1651 (N_1651,N_1234,N_1055);
nand U1652 (N_1652,N_1263,N_1292);
nand U1653 (N_1653,N_1205,N_1133);
or U1654 (N_1654,N_1236,N_1244);
nand U1655 (N_1655,N_1220,N_1041);
or U1656 (N_1656,N_1367,N_1046);
nor U1657 (N_1657,N_1054,N_1362);
nand U1658 (N_1658,N_1427,N_1277);
and U1659 (N_1659,N_1491,N_1369);
nor U1660 (N_1660,N_1333,N_1385);
or U1661 (N_1661,N_1045,N_1111);
nand U1662 (N_1662,N_1453,N_1309);
and U1663 (N_1663,N_1206,N_1168);
or U1664 (N_1664,N_1429,N_1161);
nand U1665 (N_1665,N_1121,N_1040);
nand U1666 (N_1666,N_1086,N_1349);
nand U1667 (N_1667,N_1253,N_1172);
and U1668 (N_1668,N_1248,N_1488);
or U1669 (N_1669,N_1457,N_1144);
nand U1670 (N_1670,N_1011,N_1187);
or U1671 (N_1671,N_1003,N_1009);
or U1672 (N_1672,N_1286,N_1490);
and U1673 (N_1673,N_1381,N_1005);
or U1674 (N_1674,N_1476,N_1259);
or U1675 (N_1675,N_1366,N_1252);
nor U1676 (N_1676,N_1179,N_1499);
nor U1677 (N_1677,N_1102,N_1208);
or U1678 (N_1678,N_1122,N_1171);
nand U1679 (N_1679,N_1212,N_1446);
nor U1680 (N_1680,N_1262,N_1318);
or U1681 (N_1681,N_1238,N_1013);
and U1682 (N_1682,N_1347,N_1066);
and U1683 (N_1683,N_1091,N_1275);
and U1684 (N_1684,N_1209,N_1020);
xnor U1685 (N_1685,N_1322,N_1418);
nand U1686 (N_1686,N_1351,N_1337);
and U1687 (N_1687,N_1348,N_1391);
or U1688 (N_1688,N_1495,N_1442);
nand U1689 (N_1689,N_1032,N_1454);
nand U1690 (N_1690,N_1015,N_1428);
xnor U1691 (N_1691,N_1044,N_1062);
xnor U1692 (N_1692,N_1471,N_1276);
or U1693 (N_1693,N_1258,N_1193);
nor U1694 (N_1694,N_1077,N_1000);
nor U1695 (N_1695,N_1094,N_1024);
nor U1696 (N_1696,N_1436,N_1036);
nand U1697 (N_1697,N_1441,N_1329);
nand U1698 (N_1698,N_1460,N_1123);
nor U1699 (N_1699,N_1388,N_1432);
nor U1700 (N_1700,N_1373,N_1156);
nand U1701 (N_1701,N_1447,N_1359);
or U1702 (N_1702,N_1132,N_1342);
nand U1703 (N_1703,N_1068,N_1302);
nor U1704 (N_1704,N_1177,N_1466);
and U1705 (N_1705,N_1325,N_1035);
nand U1706 (N_1706,N_1319,N_1338);
nor U1707 (N_1707,N_1118,N_1494);
nor U1708 (N_1708,N_1464,N_1440);
and U1709 (N_1709,N_1327,N_1371);
or U1710 (N_1710,N_1434,N_1399);
and U1711 (N_1711,N_1012,N_1403);
nor U1712 (N_1712,N_1226,N_1218);
nor U1713 (N_1713,N_1290,N_1485);
or U1714 (N_1714,N_1274,N_1163);
or U1715 (N_1715,N_1408,N_1095);
or U1716 (N_1716,N_1089,N_1140);
xor U1717 (N_1717,N_1119,N_1084);
nand U1718 (N_1718,N_1404,N_1343);
nor U1719 (N_1719,N_1386,N_1483);
nor U1720 (N_1720,N_1225,N_1104);
nand U1721 (N_1721,N_1437,N_1261);
nand U1722 (N_1722,N_1100,N_1061);
or U1723 (N_1723,N_1157,N_1250);
and U1724 (N_1724,N_1064,N_1146);
nor U1725 (N_1725,N_1130,N_1445);
nand U1726 (N_1726,N_1357,N_1158);
or U1727 (N_1727,N_1190,N_1078);
nor U1728 (N_1728,N_1387,N_1433);
nor U1729 (N_1729,N_1199,N_1299);
nand U1730 (N_1730,N_1472,N_1267);
and U1731 (N_1731,N_1183,N_1016);
nor U1732 (N_1732,N_1340,N_1026);
nor U1733 (N_1733,N_1059,N_1159);
nor U1734 (N_1734,N_1443,N_1415);
or U1735 (N_1735,N_1063,N_1316);
or U1736 (N_1736,N_1412,N_1426);
nor U1737 (N_1737,N_1273,N_1264);
or U1738 (N_1738,N_1458,N_1296);
nand U1739 (N_1739,N_1202,N_1147);
nor U1740 (N_1740,N_1335,N_1417);
or U1741 (N_1741,N_1105,N_1298);
xnor U1742 (N_1742,N_1098,N_1042);
or U1743 (N_1743,N_1350,N_1282);
or U1744 (N_1744,N_1384,N_1390);
nand U1745 (N_1745,N_1269,N_1356);
nand U1746 (N_1746,N_1116,N_1405);
nand U1747 (N_1747,N_1487,N_1235);
nand U1748 (N_1748,N_1213,N_1127);
xor U1749 (N_1749,N_1484,N_1058);
nor U1750 (N_1750,N_1273,N_1261);
nor U1751 (N_1751,N_1348,N_1318);
or U1752 (N_1752,N_1291,N_1263);
or U1753 (N_1753,N_1118,N_1301);
nand U1754 (N_1754,N_1006,N_1020);
and U1755 (N_1755,N_1141,N_1309);
or U1756 (N_1756,N_1474,N_1472);
and U1757 (N_1757,N_1412,N_1382);
and U1758 (N_1758,N_1472,N_1326);
nand U1759 (N_1759,N_1035,N_1458);
nand U1760 (N_1760,N_1058,N_1216);
nor U1761 (N_1761,N_1114,N_1162);
and U1762 (N_1762,N_1204,N_1137);
nand U1763 (N_1763,N_1265,N_1191);
nand U1764 (N_1764,N_1151,N_1230);
nand U1765 (N_1765,N_1054,N_1304);
nor U1766 (N_1766,N_1096,N_1136);
or U1767 (N_1767,N_1136,N_1109);
nor U1768 (N_1768,N_1160,N_1091);
nor U1769 (N_1769,N_1128,N_1169);
nand U1770 (N_1770,N_1236,N_1457);
nor U1771 (N_1771,N_1465,N_1426);
or U1772 (N_1772,N_1326,N_1145);
and U1773 (N_1773,N_1060,N_1306);
or U1774 (N_1774,N_1386,N_1421);
and U1775 (N_1775,N_1029,N_1400);
or U1776 (N_1776,N_1441,N_1003);
nor U1777 (N_1777,N_1124,N_1306);
nand U1778 (N_1778,N_1092,N_1320);
nor U1779 (N_1779,N_1429,N_1071);
or U1780 (N_1780,N_1041,N_1444);
or U1781 (N_1781,N_1497,N_1021);
or U1782 (N_1782,N_1180,N_1201);
xor U1783 (N_1783,N_1346,N_1262);
or U1784 (N_1784,N_1019,N_1012);
xor U1785 (N_1785,N_1256,N_1332);
nand U1786 (N_1786,N_1324,N_1152);
or U1787 (N_1787,N_1381,N_1194);
or U1788 (N_1788,N_1098,N_1494);
nand U1789 (N_1789,N_1310,N_1055);
nand U1790 (N_1790,N_1387,N_1267);
nor U1791 (N_1791,N_1272,N_1426);
nand U1792 (N_1792,N_1099,N_1308);
or U1793 (N_1793,N_1098,N_1364);
nand U1794 (N_1794,N_1240,N_1035);
or U1795 (N_1795,N_1321,N_1345);
nor U1796 (N_1796,N_1291,N_1098);
nand U1797 (N_1797,N_1444,N_1264);
nor U1798 (N_1798,N_1226,N_1473);
xor U1799 (N_1799,N_1020,N_1309);
nor U1800 (N_1800,N_1371,N_1169);
nor U1801 (N_1801,N_1137,N_1347);
and U1802 (N_1802,N_1079,N_1017);
and U1803 (N_1803,N_1118,N_1273);
nand U1804 (N_1804,N_1073,N_1121);
and U1805 (N_1805,N_1480,N_1216);
and U1806 (N_1806,N_1009,N_1229);
nand U1807 (N_1807,N_1203,N_1305);
nor U1808 (N_1808,N_1260,N_1163);
or U1809 (N_1809,N_1041,N_1110);
xor U1810 (N_1810,N_1079,N_1477);
nor U1811 (N_1811,N_1223,N_1070);
nor U1812 (N_1812,N_1156,N_1117);
or U1813 (N_1813,N_1196,N_1422);
and U1814 (N_1814,N_1097,N_1287);
and U1815 (N_1815,N_1258,N_1362);
and U1816 (N_1816,N_1209,N_1190);
or U1817 (N_1817,N_1204,N_1291);
nand U1818 (N_1818,N_1038,N_1037);
nand U1819 (N_1819,N_1443,N_1181);
or U1820 (N_1820,N_1234,N_1126);
nor U1821 (N_1821,N_1075,N_1364);
nor U1822 (N_1822,N_1363,N_1377);
or U1823 (N_1823,N_1410,N_1085);
and U1824 (N_1824,N_1287,N_1168);
and U1825 (N_1825,N_1447,N_1255);
nand U1826 (N_1826,N_1326,N_1074);
or U1827 (N_1827,N_1007,N_1087);
nor U1828 (N_1828,N_1494,N_1255);
or U1829 (N_1829,N_1177,N_1357);
or U1830 (N_1830,N_1074,N_1330);
nor U1831 (N_1831,N_1131,N_1241);
nand U1832 (N_1832,N_1134,N_1117);
nand U1833 (N_1833,N_1123,N_1075);
nand U1834 (N_1834,N_1476,N_1418);
or U1835 (N_1835,N_1219,N_1251);
nand U1836 (N_1836,N_1255,N_1093);
or U1837 (N_1837,N_1387,N_1407);
or U1838 (N_1838,N_1323,N_1261);
and U1839 (N_1839,N_1380,N_1108);
or U1840 (N_1840,N_1343,N_1369);
or U1841 (N_1841,N_1408,N_1353);
nor U1842 (N_1842,N_1194,N_1421);
nand U1843 (N_1843,N_1229,N_1199);
nor U1844 (N_1844,N_1399,N_1093);
nor U1845 (N_1845,N_1208,N_1008);
nor U1846 (N_1846,N_1427,N_1015);
nor U1847 (N_1847,N_1239,N_1063);
nand U1848 (N_1848,N_1376,N_1454);
and U1849 (N_1849,N_1064,N_1038);
and U1850 (N_1850,N_1386,N_1482);
and U1851 (N_1851,N_1227,N_1317);
or U1852 (N_1852,N_1336,N_1157);
nand U1853 (N_1853,N_1283,N_1147);
nor U1854 (N_1854,N_1287,N_1194);
and U1855 (N_1855,N_1144,N_1461);
nor U1856 (N_1856,N_1335,N_1249);
and U1857 (N_1857,N_1440,N_1365);
or U1858 (N_1858,N_1206,N_1036);
or U1859 (N_1859,N_1264,N_1075);
nor U1860 (N_1860,N_1366,N_1317);
nor U1861 (N_1861,N_1092,N_1420);
or U1862 (N_1862,N_1373,N_1258);
or U1863 (N_1863,N_1400,N_1229);
or U1864 (N_1864,N_1284,N_1459);
and U1865 (N_1865,N_1412,N_1056);
or U1866 (N_1866,N_1009,N_1167);
or U1867 (N_1867,N_1311,N_1421);
nand U1868 (N_1868,N_1104,N_1240);
or U1869 (N_1869,N_1311,N_1275);
or U1870 (N_1870,N_1289,N_1156);
and U1871 (N_1871,N_1387,N_1150);
nand U1872 (N_1872,N_1312,N_1234);
nand U1873 (N_1873,N_1032,N_1415);
nor U1874 (N_1874,N_1379,N_1149);
nor U1875 (N_1875,N_1262,N_1491);
nand U1876 (N_1876,N_1057,N_1017);
and U1877 (N_1877,N_1030,N_1366);
or U1878 (N_1878,N_1118,N_1256);
and U1879 (N_1879,N_1407,N_1229);
nand U1880 (N_1880,N_1350,N_1298);
xor U1881 (N_1881,N_1307,N_1123);
and U1882 (N_1882,N_1265,N_1362);
or U1883 (N_1883,N_1024,N_1422);
nor U1884 (N_1884,N_1161,N_1387);
and U1885 (N_1885,N_1336,N_1013);
nand U1886 (N_1886,N_1050,N_1197);
or U1887 (N_1887,N_1079,N_1483);
nand U1888 (N_1888,N_1211,N_1371);
or U1889 (N_1889,N_1411,N_1242);
and U1890 (N_1890,N_1459,N_1046);
nand U1891 (N_1891,N_1260,N_1349);
and U1892 (N_1892,N_1367,N_1369);
and U1893 (N_1893,N_1188,N_1039);
nand U1894 (N_1894,N_1413,N_1480);
nand U1895 (N_1895,N_1286,N_1114);
and U1896 (N_1896,N_1176,N_1249);
nand U1897 (N_1897,N_1314,N_1119);
nand U1898 (N_1898,N_1394,N_1179);
or U1899 (N_1899,N_1155,N_1138);
nand U1900 (N_1900,N_1251,N_1291);
nor U1901 (N_1901,N_1442,N_1396);
and U1902 (N_1902,N_1272,N_1325);
nor U1903 (N_1903,N_1492,N_1063);
and U1904 (N_1904,N_1306,N_1079);
nor U1905 (N_1905,N_1402,N_1047);
nand U1906 (N_1906,N_1285,N_1459);
nor U1907 (N_1907,N_1180,N_1383);
and U1908 (N_1908,N_1244,N_1168);
and U1909 (N_1909,N_1228,N_1135);
and U1910 (N_1910,N_1399,N_1318);
and U1911 (N_1911,N_1383,N_1487);
nand U1912 (N_1912,N_1074,N_1316);
and U1913 (N_1913,N_1440,N_1265);
and U1914 (N_1914,N_1137,N_1140);
and U1915 (N_1915,N_1240,N_1262);
nand U1916 (N_1916,N_1256,N_1281);
and U1917 (N_1917,N_1493,N_1404);
nand U1918 (N_1918,N_1193,N_1274);
and U1919 (N_1919,N_1196,N_1220);
nor U1920 (N_1920,N_1080,N_1149);
and U1921 (N_1921,N_1299,N_1048);
nor U1922 (N_1922,N_1010,N_1343);
or U1923 (N_1923,N_1483,N_1283);
nor U1924 (N_1924,N_1189,N_1028);
or U1925 (N_1925,N_1371,N_1060);
or U1926 (N_1926,N_1242,N_1020);
and U1927 (N_1927,N_1102,N_1101);
nand U1928 (N_1928,N_1208,N_1155);
and U1929 (N_1929,N_1286,N_1077);
and U1930 (N_1930,N_1039,N_1453);
or U1931 (N_1931,N_1373,N_1135);
and U1932 (N_1932,N_1293,N_1232);
nand U1933 (N_1933,N_1387,N_1411);
and U1934 (N_1934,N_1104,N_1224);
nor U1935 (N_1935,N_1407,N_1456);
and U1936 (N_1936,N_1352,N_1361);
and U1937 (N_1937,N_1027,N_1400);
nand U1938 (N_1938,N_1390,N_1009);
nand U1939 (N_1939,N_1208,N_1286);
nand U1940 (N_1940,N_1212,N_1448);
nand U1941 (N_1941,N_1466,N_1068);
nor U1942 (N_1942,N_1064,N_1116);
nand U1943 (N_1943,N_1363,N_1134);
and U1944 (N_1944,N_1238,N_1084);
and U1945 (N_1945,N_1306,N_1497);
or U1946 (N_1946,N_1409,N_1155);
or U1947 (N_1947,N_1296,N_1383);
nor U1948 (N_1948,N_1184,N_1099);
or U1949 (N_1949,N_1006,N_1178);
nand U1950 (N_1950,N_1459,N_1250);
and U1951 (N_1951,N_1352,N_1071);
nor U1952 (N_1952,N_1265,N_1495);
or U1953 (N_1953,N_1470,N_1194);
nand U1954 (N_1954,N_1230,N_1128);
and U1955 (N_1955,N_1490,N_1050);
and U1956 (N_1956,N_1251,N_1325);
nand U1957 (N_1957,N_1364,N_1349);
and U1958 (N_1958,N_1259,N_1336);
nand U1959 (N_1959,N_1228,N_1355);
nor U1960 (N_1960,N_1341,N_1476);
nor U1961 (N_1961,N_1358,N_1223);
nand U1962 (N_1962,N_1239,N_1354);
or U1963 (N_1963,N_1297,N_1062);
and U1964 (N_1964,N_1356,N_1172);
nor U1965 (N_1965,N_1075,N_1034);
nand U1966 (N_1966,N_1300,N_1134);
nor U1967 (N_1967,N_1410,N_1401);
or U1968 (N_1968,N_1348,N_1380);
nor U1969 (N_1969,N_1319,N_1082);
and U1970 (N_1970,N_1176,N_1135);
nand U1971 (N_1971,N_1276,N_1188);
or U1972 (N_1972,N_1284,N_1185);
and U1973 (N_1973,N_1432,N_1177);
nor U1974 (N_1974,N_1068,N_1252);
nor U1975 (N_1975,N_1179,N_1485);
and U1976 (N_1976,N_1459,N_1064);
nor U1977 (N_1977,N_1126,N_1236);
and U1978 (N_1978,N_1363,N_1119);
or U1979 (N_1979,N_1376,N_1105);
xnor U1980 (N_1980,N_1119,N_1004);
or U1981 (N_1981,N_1281,N_1484);
and U1982 (N_1982,N_1404,N_1043);
nand U1983 (N_1983,N_1020,N_1236);
nor U1984 (N_1984,N_1299,N_1419);
and U1985 (N_1985,N_1476,N_1173);
and U1986 (N_1986,N_1101,N_1498);
and U1987 (N_1987,N_1011,N_1303);
nor U1988 (N_1988,N_1262,N_1122);
or U1989 (N_1989,N_1487,N_1131);
and U1990 (N_1990,N_1321,N_1327);
and U1991 (N_1991,N_1036,N_1261);
nor U1992 (N_1992,N_1298,N_1068);
nand U1993 (N_1993,N_1184,N_1446);
nand U1994 (N_1994,N_1050,N_1317);
nand U1995 (N_1995,N_1107,N_1494);
nor U1996 (N_1996,N_1347,N_1318);
nand U1997 (N_1997,N_1367,N_1136);
and U1998 (N_1998,N_1112,N_1117);
nor U1999 (N_1999,N_1364,N_1392);
nor U2000 (N_2000,N_1963,N_1987);
nand U2001 (N_2001,N_1514,N_1622);
nor U2002 (N_2002,N_1841,N_1685);
or U2003 (N_2003,N_1783,N_1529);
nand U2004 (N_2004,N_1637,N_1960);
or U2005 (N_2005,N_1923,N_1997);
nand U2006 (N_2006,N_1786,N_1628);
nor U2007 (N_2007,N_1870,N_1608);
nand U2008 (N_2008,N_1555,N_1597);
and U2009 (N_2009,N_1598,N_1545);
and U2010 (N_2010,N_1862,N_1928);
xor U2011 (N_2011,N_1775,N_1701);
nand U2012 (N_2012,N_1669,N_1714);
nor U2013 (N_2013,N_1889,N_1611);
nor U2014 (N_2014,N_1770,N_1906);
nor U2015 (N_2015,N_1694,N_1926);
nand U2016 (N_2016,N_1808,N_1869);
and U2017 (N_2017,N_1682,N_1924);
nand U2018 (N_2018,N_1740,N_1919);
nor U2019 (N_2019,N_1686,N_1765);
xor U2020 (N_2020,N_1847,N_1848);
nor U2021 (N_2021,N_1874,N_1959);
nor U2022 (N_2022,N_1935,N_1780);
nor U2023 (N_2023,N_1717,N_1534);
and U2024 (N_2024,N_1993,N_1867);
and U2025 (N_2025,N_1676,N_1502);
nor U2026 (N_2026,N_1724,N_1991);
nor U2027 (N_2027,N_1737,N_1704);
nand U2028 (N_2028,N_1673,N_1544);
nor U2029 (N_2029,N_1679,N_1976);
and U2030 (N_2030,N_1984,N_1699);
nor U2031 (N_2031,N_1722,N_1553);
nor U2032 (N_2032,N_1500,N_1620);
nand U2033 (N_2033,N_1680,N_1633);
or U2034 (N_2034,N_1695,N_1768);
or U2035 (N_2035,N_1910,N_1515);
nor U2036 (N_2036,N_1785,N_1845);
and U2037 (N_2037,N_1618,N_1658);
and U2038 (N_2038,N_1754,N_1512);
nand U2039 (N_2039,N_1812,N_1944);
nand U2040 (N_2040,N_1942,N_1784);
or U2041 (N_2041,N_1904,N_1798);
or U2042 (N_2042,N_1882,N_1829);
or U2043 (N_2043,N_1858,N_1623);
nand U2044 (N_2044,N_1833,N_1816);
nand U2045 (N_2045,N_1805,N_1814);
or U2046 (N_2046,N_1751,N_1966);
nand U2047 (N_2047,N_1563,N_1764);
nand U2048 (N_2048,N_1716,N_1688);
nor U2049 (N_2049,N_1649,N_1953);
and U2050 (N_2050,N_1871,N_1659);
nand U2051 (N_2051,N_1605,N_1771);
or U2052 (N_2052,N_1762,N_1840);
nand U2053 (N_2053,N_1733,N_1773);
nor U2054 (N_2054,N_1913,N_1731);
and U2055 (N_2055,N_1647,N_1550);
nand U2056 (N_2056,N_1666,N_1962);
nor U2057 (N_2057,N_1799,N_1629);
nand U2058 (N_2058,N_1908,N_1978);
nor U2059 (N_2059,N_1547,N_1895);
nand U2060 (N_2060,N_1901,N_1561);
or U2061 (N_2061,N_1789,N_1711);
nand U2062 (N_2062,N_1982,N_1892);
or U2063 (N_2063,N_1571,N_1943);
and U2064 (N_2064,N_1807,N_1549);
nand U2065 (N_2065,N_1811,N_1893);
or U2066 (N_2066,N_1533,N_1619);
nor U2067 (N_2067,N_1590,N_1505);
and U2068 (N_2068,N_1625,N_1579);
nor U2069 (N_2069,N_1653,N_1661);
and U2070 (N_2070,N_1902,N_1715);
and U2071 (N_2071,N_1802,N_1531);
and U2072 (N_2072,N_1756,N_1885);
and U2073 (N_2073,N_1994,N_1678);
and U2074 (N_2074,N_1918,N_1983);
or U2075 (N_2075,N_1872,N_1951);
nor U2076 (N_2076,N_1850,N_1566);
and U2077 (N_2077,N_1965,N_1738);
and U2078 (N_2078,N_1543,N_1856);
and U2079 (N_2079,N_1873,N_1638);
and U2080 (N_2080,N_1890,N_1725);
nor U2081 (N_2081,N_1642,N_1650);
or U2082 (N_2082,N_1996,N_1909);
and U2083 (N_2083,N_1745,N_1831);
and U2084 (N_2084,N_1552,N_1970);
or U2085 (N_2085,N_1956,N_1761);
nand U2086 (N_2086,N_1538,N_1684);
or U2087 (N_2087,N_1662,N_1578);
nand U2088 (N_2088,N_1851,N_1922);
or U2089 (N_2089,N_1930,N_1528);
nor U2090 (N_2090,N_1648,N_1532);
and U2091 (N_2091,N_1536,N_1655);
and U2092 (N_2092,N_1573,N_1739);
or U2093 (N_2093,N_1884,N_1626);
nand U2094 (N_2094,N_1986,N_1583);
nand U2095 (N_2095,N_1757,N_1779);
and U2096 (N_2096,N_1792,N_1506);
or U2097 (N_2097,N_1830,N_1663);
or U2098 (N_2098,N_1636,N_1689);
and U2099 (N_2099,N_1957,N_1881);
nor U2100 (N_2100,N_1593,N_1601);
xor U2101 (N_2101,N_1769,N_1972);
nand U2102 (N_2102,N_1609,N_1835);
and U2103 (N_2103,N_1513,N_1946);
nor U2104 (N_2104,N_1582,N_1572);
or U2105 (N_2105,N_1778,N_1866);
nand U2106 (N_2106,N_1511,N_1743);
nor U2107 (N_2107,N_1999,N_1592);
nor U2108 (N_2108,N_1646,N_1879);
and U2109 (N_2109,N_1794,N_1947);
and U2110 (N_2110,N_1693,N_1574);
nor U2111 (N_2111,N_1788,N_1595);
or U2112 (N_2112,N_1969,N_1599);
nand U2113 (N_2113,N_1624,N_1971);
and U2114 (N_2114,N_1846,N_1720);
nor U2115 (N_2115,N_1767,N_1613);
nand U2116 (N_2116,N_1985,N_1735);
or U2117 (N_2117,N_1643,N_1916);
or U2118 (N_2118,N_1558,N_1979);
nand U2119 (N_2119,N_1749,N_1857);
nor U2120 (N_2120,N_1907,N_1824);
nand U2121 (N_2121,N_1782,N_1632);
or U2122 (N_2122,N_1793,N_1995);
or U2123 (N_2123,N_1883,N_1729);
nor U2124 (N_2124,N_1617,N_1852);
or U2125 (N_2125,N_1600,N_1507);
nor U2126 (N_2126,N_1791,N_1570);
or U2127 (N_2127,N_1700,N_1839);
and U2128 (N_2128,N_1774,N_1865);
and U2129 (N_2129,N_1668,N_1980);
or U2130 (N_2130,N_1554,N_1690);
nand U2131 (N_2131,N_1838,N_1525);
xor U2132 (N_2132,N_1569,N_1763);
nand U2133 (N_2133,N_1880,N_1821);
nand U2134 (N_2134,N_1974,N_1886);
nor U2135 (N_2135,N_1567,N_1758);
and U2136 (N_2136,N_1897,N_1925);
nand U2137 (N_2137,N_1940,N_1530);
nor U2138 (N_2138,N_1557,N_1990);
and U2139 (N_2139,N_1713,N_1508);
nand U2140 (N_2140,N_1568,N_1967);
nor U2141 (N_2141,N_1501,N_1518);
and U2142 (N_2142,N_1546,N_1896);
and U2143 (N_2143,N_1683,N_1988);
nand U2144 (N_2144,N_1681,N_1527);
nand U2145 (N_2145,N_1651,N_1698);
nor U2146 (N_2146,N_1702,N_1521);
nand U2147 (N_2147,N_1836,N_1900);
and U2148 (N_2148,N_1864,N_1610);
nand U2149 (N_2149,N_1520,N_1750);
nand U2150 (N_2150,N_1721,N_1730);
or U2151 (N_2151,N_1576,N_1759);
nor U2152 (N_2152,N_1992,N_1644);
nor U2153 (N_2153,N_1586,N_1732);
and U2154 (N_2154,N_1596,N_1975);
nand U2155 (N_2155,N_1818,N_1652);
or U2156 (N_2156,N_1815,N_1604);
nor U2157 (N_2157,N_1559,N_1888);
or U2158 (N_2158,N_1958,N_1674);
or U2159 (N_2159,N_1823,N_1706);
nand U2160 (N_2160,N_1937,N_1667);
or U2161 (N_2161,N_1664,N_1849);
nor U2162 (N_2162,N_1863,N_1854);
nand U2163 (N_2163,N_1710,N_1998);
nand U2164 (N_2164,N_1938,N_1627);
and U2165 (N_2165,N_1537,N_1645);
or U2166 (N_2166,N_1927,N_1606);
or U2167 (N_2167,N_1542,N_1726);
nor U2168 (N_2168,N_1934,N_1719);
nand U2169 (N_2169,N_1703,N_1800);
or U2170 (N_2170,N_1709,N_1898);
nand U2171 (N_2171,N_1837,N_1548);
or U2172 (N_2172,N_1950,N_1932);
and U2173 (N_2173,N_1585,N_1760);
xnor U2174 (N_2174,N_1822,N_1656);
or U2175 (N_2175,N_1945,N_1630);
and U2176 (N_2176,N_1868,N_1806);
and U2177 (N_2177,N_1591,N_1936);
nor U2178 (N_2178,N_1587,N_1781);
or U2179 (N_2179,N_1708,N_1891);
nor U2180 (N_2180,N_1671,N_1861);
nand U2181 (N_2181,N_1660,N_1589);
nand U2182 (N_2182,N_1878,N_1968);
nor U2183 (N_2183,N_1640,N_1921);
nor U2184 (N_2184,N_1635,N_1657);
nand U2185 (N_2185,N_1817,N_1539);
and U2186 (N_2186,N_1639,N_1809);
nand U2187 (N_2187,N_1577,N_1772);
nand U2188 (N_2188,N_1672,N_1594);
and U2189 (N_2189,N_1939,N_1931);
nand U2190 (N_2190,N_1955,N_1556);
nand U2191 (N_2191,N_1575,N_1551);
and U2192 (N_2192,N_1755,N_1920);
or U2193 (N_2193,N_1712,N_1826);
or U2194 (N_2194,N_1853,N_1941);
or U2195 (N_2195,N_1813,N_1894);
nand U2196 (N_2196,N_1753,N_1790);
and U2197 (N_2197,N_1981,N_1509);
nand U2198 (N_2198,N_1564,N_1616);
nor U2199 (N_2199,N_1977,N_1696);
nand U2200 (N_2200,N_1752,N_1746);
and U2201 (N_2201,N_1631,N_1949);
or U2202 (N_2202,N_1670,N_1584);
nand U2203 (N_2203,N_1522,N_1825);
or U2204 (N_2204,N_1634,N_1804);
or U2205 (N_2205,N_1607,N_1948);
or U2206 (N_2206,N_1675,N_1517);
and U2207 (N_2207,N_1503,N_1766);
nand U2208 (N_2208,N_1929,N_1819);
or U2209 (N_2209,N_1723,N_1614);
and U2210 (N_2210,N_1526,N_1603);
and U2211 (N_2211,N_1843,N_1615);
nand U2212 (N_2212,N_1828,N_1973);
and U2213 (N_2213,N_1787,N_1727);
nor U2214 (N_2214,N_1860,N_1887);
nor U2215 (N_2215,N_1560,N_1621);
nor U2216 (N_2216,N_1795,N_1803);
and U2217 (N_2217,N_1734,N_1535);
and U2218 (N_2218,N_1899,N_1612);
or U2219 (N_2219,N_1796,N_1912);
nand U2220 (N_2220,N_1705,N_1915);
nor U2221 (N_2221,N_1504,N_1580);
nand U2222 (N_2222,N_1832,N_1641);
and U2223 (N_2223,N_1961,N_1741);
or U2224 (N_2224,N_1728,N_1540);
or U2225 (N_2225,N_1933,N_1744);
or U2226 (N_2226,N_1516,N_1523);
nand U2227 (N_2227,N_1827,N_1964);
nor U2228 (N_2228,N_1602,N_1718);
or U2229 (N_2229,N_1677,N_1687);
nand U2230 (N_2230,N_1581,N_1665);
nor U2231 (N_2231,N_1911,N_1844);
and U2232 (N_2232,N_1776,N_1707);
nor U2233 (N_2233,N_1777,N_1859);
nand U2234 (N_2234,N_1742,N_1692);
and U2235 (N_2235,N_1565,N_1654);
or U2236 (N_2236,N_1562,N_1917);
nand U2237 (N_2237,N_1736,N_1541);
or U2238 (N_2238,N_1748,N_1820);
xor U2239 (N_2239,N_1747,N_1876);
or U2240 (N_2240,N_1989,N_1524);
or U2241 (N_2241,N_1842,N_1905);
nor U2242 (N_2242,N_1697,N_1510);
nor U2243 (N_2243,N_1952,N_1914);
or U2244 (N_2244,N_1903,N_1797);
and U2245 (N_2245,N_1877,N_1691);
nor U2246 (N_2246,N_1875,N_1810);
xor U2247 (N_2247,N_1801,N_1834);
nor U2248 (N_2248,N_1855,N_1519);
nand U2249 (N_2249,N_1588,N_1954);
and U2250 (N_2250,N_1760,N_1641);
nand U2251 (N_2251,N_1865,N_1863);
or U2252 (N_2252,N_1990,N_1994);
nor U2253 (N_2253,N_1839,N_1637);
nand U2254 (N_2254,N_1763,N_1523);
or U2255 (N_2255,N_1862,N_1665);
nand U2256 (N_2256,N_1688,N_1517);
xor U2257 (N_2257,N_1543,N_1714);
nand U2258 (N_2258,N_1973,N_1673);
or U2259 (N_2259,N_1652,N_1953);
nor U2260 (N_2260,N_1640,N_1521);
and U2261 (N_2261,N_1886,N_1676);
nor U2262 (N_2262,N_1749,N_1742);
or U2263 (N_2263,N_1791,N_1775);
nand U2264 (N_2264,N_1974,N_1937);
or U2265 (N_2265,N_1673,N_1607);
or U2266 (N_2266,N_1801,N_1777);
or U2267 (N_2267,N_1873,N_1990);
and U2268 (N_2268,N_1757,N_1535);
and U2269 (N_2269,N_1829,N_1926);
nor U2270 (N_2270,N_1708,N_1906);
and U2271 (N_2271,N_1512,N_1605);
or U2272 (N_2272,N_1819,N_1888);
nand U2273 (N_2273,N_1955,N_1960);
nand U2274 (N_2274,N_1622,N_1535);
or U2275 (N_2275,N_1690,N_1761);
nor U2276 (N_2276,N_1671,N_1954);
or U2277 (N_2277,N_1623,N_1509);
or U2278 (N_2278,N_1955,N_1641);
and U2279 (N_2279,N_1845,N_1667);
or U2280 (N_2280,N_1858,N_1876);
or U2281 (N_2281,N_1866,N_1911);
nor U2282 (N_2282,N_1801,N_1534);
nor U2283 (N_2283,N_1679,N_1999);
or U2284 (N_2284,N_1822,N_1549);
nand U2285 (N_2285,N_1721,N_1925);
or U2286 (N_2286,N_1577,N_1878);
or U2287 (N_2287,N_1956,N_1669);
and U2288 (N_2288,N_1823,N_1527);
or U2289 (N_2289,N_1591,N_1612);
nor U2290 (N_2290,N_1637,N_1693);
nand U2291 (N_2291,N_1708,N_1635);
or U2292 (N_2292,N_1685,N_1620);
nor U2293 (N_2293,N_1633,N_1509);
nand U2294 (N_2294,N_1841,N_1750);
nor U2295 (N_2295,N_1538,N_1566);
nand U2296 (N_2296,N_1577,N_1634);
and U2297 (N_2297,N_1601,N_1909);
or U2298 (N_2298,N_1888,N_1782);
nand U2299 (N_2299,N_1958,N_1983);
nand U2300 (N_2300,N_1925,N_1805);
nand U2301 (N_2301,N_1613,N_1805);
nor U2302 (N_2302,N_1950,N_1590);
nand U2303 (N_2303,N_1551,N_1857);
and U2304 (N_2304,N_1600,N_1646);
or U2305 (N_2305,N_1874,N_1924);
nand U2306 (N_2306,N_1503,N_1990);
nand U2307 (N_2307,N_1813,N_1553);
nor U2308 (N_2308,N_1662,N_1995);
nand U2309 (N_2309,N_1620,N_1900);
and U2310 (N_2310,N_1888,N_1715);
or U2311 (N_2311,N_1951,N_1745);
nor U2312 (N_2312,N_1691,N_1749);
or U2313 (N_2313,N_1643,N_1636);
nor U2314 (N_2314,N_1663,N_1696);
nand U2315 (N_2315,N_1964,N_1911);
or U2316 (N_2316,N_1897,N_1759);
or U2317 (N_2317,N_1679,N_1600);
nand U2318 (N_2318,N_1858,N_1733);
or U2319 (N_2319,N_1827,N_1997);
nand U2320 (N_2320,N_1911,N_1975);
or U2321 (N_2321,N_1724,N_1596);
and U2322 (N_2322,N_1745,N_1869);
or U2323 (N_2323,N_1614,N_1524);
nand U2324 (N_2324,N_1850,N_1565);
and U2325 (N_2325,N_1646,N_1662);
and U2326 (N_2326,N_1799,N_1706);
nor U2327 (N_2327,N_1595,N_1672);
or U2328 (N_2328,N_1544,N_1618);
and U2329 (N_2329,N_1960,N_1864);
or U2330 (N_2330,N_1762,N_1622);
or U2331 (N_2331,N_1960,N_1828);
or U2332 (N_2332,N_1662,N_1828);
and U2333 (N_2333,N_1558,N_1598);
xor U2334 (N_2334,N_1978,N_1773);
nand U2335 (N_2335,N_1822,N_1943);
nor U2336 (N_2336,N_1848,N_1509);
nand U2337 (N_2337,N_1758,N_1726);
or U2338 (N_2338,N_1832,N_1651);
nor U2339 (N_2339,N_1938,N_1954);
or U2340 (N_2340,N_1739,N_1895);
nor U2341 (N_2341,N_1812,N_1693);
nand U2342 (N_2342,N_1756,N_1795);
nand U2343 (N_2343,N_1536,N_1987);
or U2344 (N_2344,N_1856,N_1936);
nor U2345 (N_2345,N_1518,N_1530);
or U2346 (N_2346,N_1544,N_1617);
or U2347 (N_2347,N_1973,N_1842);
and U2348 (N_2348,N_1716,N_1844);
nor U2349 (N_2349,N_1711,N_1767);
nand U2350 (N_2350,N_1556,N_1555);
or U2351 (N_2351,N_1713,N_1632);
or U2352 (N_2352,N_1524,N_1666);
and U2353 (N_2353,N_1940,N_1716);
nand U2354 (N_2354,N_1606,N_1995);
nor U2355 (N_2355,N_1685,N_1821);
nor U2356 (N_2356,N_1534,N_1787);
and U2357 (N_2357,N_1674,N_1775);
nand U2358 (N_2358,N_1891,N_1514);
xnor U2359 (N_2359,N_1707,N_1819);
nand U2360 (N_2360,N_1843,N_1589);
xor U2361 (N_2361,N_1783,N_1770);
or U2362 (N_2362,N_1754,N_1723);
and U2363 (N_2363,N_1957,N_1528);
nand U2364 (N_2364,N_1805,N_1915);
nand U2365 (N_2365,N_1771,N_1523);
and U2366 (N_2366,N_1531,N_1844);
nor U2367 (N_2367,N_1686,N_1741);
and U2368 (N_2368,N_1690,N_1862);
nand U2369 (N_2369,N_1637,N_1707);
nand U2370 (N_2370,N_1586,N_1891);
or U2371 (N_2371,N_1546,N_1948);
and U2372 (N_2372,N_1561,N_1752);
nor U2373 (N_2373,N_1522,N_1746);
nor U2374 (N_2374,N_1743,N_1774);
or U2375 (N_2375,N_1974,N_1817);
or U2376 (N_2376,N_1722,N_1570);
nand U2377 (N_2377,N_1756,N_1767);
and U2378 (N_2378,N_1719,N_1769);
or U2379 (N_2379,N_1561,N_1637);
or U2380 (N_2380,N_1873,N_1848);
nor U2381 (N_2381,N_1996,N_1535);
or U2382 (N_2382,N_1970,N_1701);
and U2383 (N_2383,N_1580,N_1617);
nand U2384 (N_2384,N_1718,N_1697);
xor U2385 (N_2385,N_1732,N_1927);
nor U2386 (N_2386,N_1888,N_1910);
or U2387 (N_2387,N_1870,N_1733);
and U2388 (N_2388,N_1624,N_1680);
or U2389 (N_2389,N_1761,N_1531);
nand U2390 (N_2390,N_1869,N_1978);
and U2391 (N_2391,N_1774,N_1800);
nor U2392 (N_2392,N_1512,N_1574);
nor U2393 (N_2393,N_1990,N_1616);
and U2394 (N_2394,N_1851,N_1639);
nand U2395 (N_2395,N_1536,N_1503);
nand U2396 (N_2396,N_1752,N_1509);
or U2397 (N_2397,N_1778,N_1635);
nand U2398 (N_2398,N_1833,N_1795);
or U2399 (N_2399,N_1955,N_1842);
xor U2400 (N_2400,N_1554,N_1880);
and U2401 (N_2401,N_1906,N_1919);
and U2402 (N_2402,N_1911,N_1847);
nand U2403 (N_2403,N_1881,N_1738);
nand U2404 (N_2404,N_1784,N_1988);
or U2405 (N_2405,N_1573,N_1603);
nor U2406 (N_2406,N_1994,N_1755);
xor U2407 (N_2407,N_1508,N_1562);
nand U2408 (N_2408,N_1942,N_1524);
and U2409 (N_2409,N_1610,N_1620);
nor U2410 (N_2410,N_1934,N_1670);
nand U2411 (N_2411,N_1636,N_1522);
or U2412 (N_2412,N_1660,N_1595);
or U2413 (N_2413,N_1558,N_1938);
nor U2414 (N_2414,N_1591,N_1815);
or U2415 (N_2415,N_1858,N_1973);
nand U2416 (N_2416,N_1552,N_1955);
nor U2417 (N_2417,N_1717,N_1764);
nand U2418 (N_2418,N_1648,N_1542);
and U2419 (N_2419,N_1909,N_1617);
xnor U2420 (N_2420,N_1932,N_1775);
xor U2421 (N_2421,N_1756,N_1848);
or U2422 (N_2422,N_1706,N_1813);
or U2423 (N_2423,N_1868,N_1628);
and U2424 (N_2424,N_1645,N_1670);
nand U2425 (N_2425,N_1999,N_1822);
or U2426 (N_2426,N_1534,N_1759);
nand U2427 (N_2427,N_1618,N_1500);
nor U2428 (N_2428,N_1739,N_1937);
and U2429 (N_2429,N_1898,N_1537);
and U2430 (N_2430,N_1716,N_1946);
or U2431 (N_2431,N_1720,N_1732);
nor U2432 (N_2432,N_1519,N_1860);
nor U2433 (N_2433,N_1920,N_1982);
or U2434 (N_2434,N_1554,N_1934);
nor U2435 (N_2435,N_1605,N_1696);
and U2436 (N_2436,N_1577,N_1678);
nor U2437 (N_2437,N_1537,N_1787);
nor U2438 (N_2438,N_1885,N_1781);
nand U2439 (N_2439,N_1655,N_1816);
or U2440 (N_2440,N_1672,N_1664);
xor U2441 (N_2441,N_1887,N_1894);
and U2442 (N_2442,N_1995,N_1776);
or U2443 (N_2443,N_1586,N_1775);
and U2444 (N_2444,N_1531,N_1674);
or U2445 (N_2445,N_1644,N_1645);
nor U2446 (N_2446,N_1890,N_1537);
nand U2447 (N_2447,N_1506,N_1810);
or U2448 (N_2448,N_1937,N_1862);
nand U2449 (N_2449,N_1967,N_1962);
or U2450 (N_2450,N_1562,N_1851);
nand U2451 (N_2451,N_1515,N_1898);
and U2452 (N_2452,N_1500,N_1528);
xnor U2453 (N_2453,N_1956,N_1821);
nor U2454 (N_2454,N_1946,N_1693);
nor U2455 (N_2455,N_1991,N_1528);
or U2456 (N_2456,N_1807,N_1751);
nand U2457 (N_2457,N_1838,N_1522);
and U2458 (N_2458,N_1538,N_1768);
nor U2459 (N_2459,N_1920,N_1687);
nand U2460 (N_2460,N_1983,N_1960);
nor U2461 (N_2461,N_1870,N_1589);
nor U2462 (N_2462,N_1812,N_1531);
nor U2463 (N_2463,N_1531,N_1847);
or U2464 (N_2464,N_1630,N_1861);
nor U2465 (N_2465,N_1803,N_1531);
nor U2466 (N_2466,N_1633,N_1833);
or U2467 (N_2467,N_1803,N_1619);
and U2468 (N_2468,N_1969,N_1589);
and U2469 (N_2469,N_1991,N_1888);
nor U2470 (N_2470,N_1765,N_1976);
or U2471 (N_2471,N_1666,N_1675);
or U2472 (N_2472,N_1845,N_1883);
nand U2473 (N_2473,N_1551,N_1825);
or U2474 (N_2474,N_1989,N_1781);
or U2475 (N_2475,N_1520,N_1661);
and U2476 (N_2476,N_1902,N_1644);
nor U2477 (N_2477,N_1966,N_1653);
or U2478 (N_2478,N_1993,N_1885);
xor U2479 (N_2479,N_1586,N_1857);
or U2480 (N_2480,N_1526,N_1922);
nor U2481 (N_2481,N_1612,N_1553);
nand U2482 (N_2482,N_1872,N_1836);
or U2483 (N_2483,N_1926,N_1892);
nor U2484 (N_2484,N_1779,N_1928);
nand U2485 (N_2485,N_1864,N_1609);
and U2486 (N_2486,N_1521,N_1656);
nor U2487 (N_2487,N_1736,N_1725);
or U2488 (N_2488,N_1774,N_1763);
nor U2489 (N_2489,N_1801,N_1643);
nand U2490 (N_2490,N_1581,N_1691);
nor U2491 (N_2491,N_1788,N_1688);
and U2492 (N_2492,N_1574,N_1543);
and U2493 (N_2493,N_1863,N_1762);
nand U2494 (N_2494,N_1698,N_1947);
xor U2495 (N_2495,N_1805,N_1858);
nand U2496 (N_2496,N_1533,N_1807);
nand U2497 (N_2497,N_1506,N_1764);
nand U2498 (N_2498,N_1560,N_1937);
nor U2499 (N_2499,N_1648,N_1618);
nor U2500 (N_2500,N_2331,N_2101);
nor U2501 (N_2501,N_2151,N_2223);
nor U2502 (N_2502,N_2181,N_2452);
xnor U2503 (N_2503,N_2036,N_2350);
or U2504 (N_2504,N_2116,N_2005);
and U2505 (N_2505,N_2374,N_2209);
and U2506 (N_2506,N_2106,N_2333);
and U2507 (N_2507,N_2395,N_2236);
nand U2508 (N_2508,N_2024,N_2413);
nor U2509 (N_2509,N_2100,N_2021);
and U2510 (N_2510,N_2004,N_2317);
and U2511 (N_2511,N_2433,N_2414);
or U2512 (N_2512,N_2308,N_2407);
nor U2513 (N_2513,N_2427,N_2282);
and U2514 (N_2514,N_2243,N_2474);
nand U2515 (N_2515,N_2097,N_2307);
nand U2516 (N_2516,N_2208,N_2083);
nand U2517 (N_2517,N_2439,N_2325);
and U2518 (N_2518,N_2330,N_2456);
and U2519 (N_2519,N_2276,N_2000);
nand U2520 (N_2520,N_2309,N_2112);
or U2521 (N_2521,N_2258,N_2498);
and U2522 (N_2522,N_2271,N_2008);
nand U2523 (N_2523,N_2445,N_2047);
nand U2524 (N_2524,N_2312,N_2486);
nand U2525 (N_2525,N_2449,N_2465);
xnor U2526 (N_2526,N_2180,N_2094);
nand U2527 (N_2527,N_2175,N_2038);
nor U2528 (N_2528,N_2461,N_2107);
or U2529 (N_2529,N_2394,N_2377);
nor U2530 (N_2530,N_2313,N_2393);
or U2531 (N_2531,N_2168,N_2206);
nand U2532 (N_2532,N_2251,N_2010);
and U2533 (N_2533,N_2370,N_2196);
nor U2534 (N_2534,N_2262,N_2401);
nor U2535 (N_2535,N_2037,N_2027);
and U2536 (N_2536,N_2074,N_2232);
nand U2537 (N_2537,N_2314,N_2332);
nor U2538 (N_2538,N_2230,N_2275);
and U2539 (N_2539,N_2158,N_2020);
and U2540 (N_2540,N_2475,N_2328);
nand U2541 (N_2541,N_2029,N_2466);
and U2542 (N_2542,N_2219,N_2227);
and U2543 (N_2543,N_2342,N_2199);
nand U2544 (N_2544,N_2316,N_2381);
or U2545 (N_2545,N_2244,N_2139);
nand U2546 (N_2546,N_2354,N_2338);
or U2547 (N_2547,N_2120,N_2458);
nand U2548 (N_2548,N_2075,N_2015);
nand U2549 (N_2549,N_2294,N_2185);
nor U2550 (N_2550,N_2143,N_2025);
nand U2551 (N_2551,N_2174,N_2007);
or U2552 (N_2552,N_2216,N_2238);
nor U2553 (N_2553,N_2051,N_2079);
or U2554 (N_2554,N_2135,N_2272);
nor U2555 (N_2555,N_2059,N_2121);
xor U2556 (N_2556,N_2281,N_2299);
nor U2557 (N_2557,N_2039,N_2469);
xor U2558 (N_2558,N_2419,N_2129);
nand U2559 (N_2559,N_2428,N_2453);
or U2560 (N_2560,N_2416,N_2434);
nor U2561 (N_2561,N_2493,N_2013);
and U2562 (N_2562,N_2494,N_2470);
or U2563 (N_2563,N_2249,N_2431);
and U2564 (N_2564,N_2357,N_2399);
or U2565 (N_2565,N_2390,N_2489);
or U2566 (N_2566,N_2435,N_2321);
nor U2567 (N_2567,N_2454,N_2149);
and U2568 (N_2568,N_2193,N_2257);
and U2569 (N_2569,N_2422,N_2256);
or U2570 (N_2570,N_2204,N_2405);
or U2571 (N_2571,N_2081,N_2103);
nor U2572 (N_2572,N_2347,N_2064);
and U2573 (N_2573,N_2341,N_2063);
nand U2574 (N_2574,N_2173,N_2468);
nand U2575 (N_2575,N_2187,N_2166);
nand U2576 (N_2576,N_2011,N_2348);
nor U2577 (N_2577,N_2283,N_2300);
nor U2578 (N_2578,N_2162,N_2177);
nor U2579 (N_2579,N_2072,N_2085);
nor U2580 (N_2580,N_2440,N_2268);
nand U2581 (N_2581,N_2183,N_2473);
nand U2582 (N_2582,N_2319,N_2387);
nand U2583 (N_2583,N_2457,N_2197);
nor U2584 (N_2584,N_2302,N_2030);
and U2585 (N_2585,N_2455,N_2369);
nor U2586 (N_2586,N_2430,N_2014);
and U2587 (N_2587,N_2144,N_2136);
nor U2588 (N_2588,N_2046,N_2250);
or U2589 (N_2589,N_2156,N_2436);
nand U2590 (N_2590,N_2049,N_2084);
nand U2591 (N_2591,N_2442,N_2198);
and U2592 (N_2592,N_2484,N_2202);
nor U2593 (N_2593,N_2362,N_2483);
nor U2594 (N_2594,N_2337,N_2041);
nand U2595 (N_2595,N_2190,N_2218);
nor U2596 (N_2596,N_2087,N_2360);
nor U2597 (N_2597,N_2404,N_2071);
and U2598 (N_2598,N_2496,N_2363);
nor U2599 (N_2599,N_2495,N_2217);
xnor U2600 (N_2600,N_2491,N_2476);
or U2601 (N_2601,N_2001,N_2392);
and U2602 (N_2602,N_2095,N_2346);
nor U2603 (N_2603,N_2421,N_2044);
nor U2604 (N_2604,N_2311,N_2022);
nor U2605 (N_2605,N_2032,N_2248);
nor U2606 (N_2606,N_2189,N_2420);
and U2607 (N_2607,N_2142,N_2327);
or U2608 (N_2608,N_2203,N_2479);
or U2609 (N_2609,N_2304,N_2114);
nand U2610 (N_2610,N_2161,N_2228);
nor U2611 (N_2611,N_2205,N_2090);
and U2612 (N_2612,N_2418,N_2165);
and U2613 (N_2613,N_2380,N_2066);
nand U2614 (N_2614,N_2226,N_2211);
and U2615 (N_2615,N_2225,N_2006);
nor U2616 (N_2616,N_2355,N_2176);
nand U2617 (N_2617,N_2270,N_2126);
nor U2618 (N_2618,N_2229,N_2086);
nand U2619 (N_2619,N_2222,N_2012);
or U2620 (N_2620,N_2295,N_2409);
or U2621 (N_2621,N_2368,N_2343);
or U2622 (N_2622,N_2289,N_2105);
or U2623 (N_2623,N_2061,N_2154);
or U2624 (N_2624,N_2091,N_2115);
and U2625 (N_2625,N_2467,N_2089);
nor U2626 (N_2626,N_2220,N_2118);
or U2627 (N_2627,N_2157,N_2048);
and U2628 (N_2628,N_2246,N_2367);
and U2629 (N_2629,N_2386,N_2212);
nor U2630 (N_2630,N_2371,N_2125);
nand U2631 (N_2631,N_2134,N_2352);
or U2632 (N_2632,N_2245,N_2293);
nor U2633 (N_2633,N_2376,N_2096);
nand U2634 (N_2634,N_2344,N_2122);
nor U2635 (N_2635,N_2358,N_2067);
nand U2636 (N_2636,N_2318,N_2102);
and U2637 (N_2637,N_2159,N_2372);
nor U2638 (N_2638,N_2266,N_2057);
nand U2639 (N_2639,N_2378,N_2045);
nor U2640 (N_2640,N_2278,N_2412);
nand U2641 (N_2641,N_2138,N_2373);
or U2642 (N_2642,N_2073,N_2462);
nand U2643 (N_2643,N_2234,N_2028);
nor U2644 (N_2644,N_2402,N_2297);
nand U2645 (N_2645,N_2425,N_2472);
nor U2646 (N_2646,N_2265,N_2329);
and U2647 (N_2647,N_2252,N_2448);
and U2648 (N_2648,N_2303,N_2411);
nand U2649 (N_2649,N_2060,N_2172);
or U2650 (N_2650,N_2026,N_2108);
xnor U2651 (N_2651,N_2273,N_2137);
or U2652 (N_2652,N_2323,N_2443);
nor U2653 (N_2653,N_2379,N_2043);
and U2654 (N_2654,N_2191,N_2023);
and U2655 (N_2655,N_2365,N_2444);
nor U2656 (N_2656,N_2253,N_2383);
or U2657 (N_2657,N_2356,N_2082);
xor U2658 (N_2658,N_2451,N_2147);
nand U2659 (N_2659,N_2153,N_2132);
and U2660 (N_2660,N_2182,N_2396);
or U2661 (N_2661,N_2408,N_2167);
and U2662 (N_2662,N_2235,N_2259);
and U2663 (N_2663,N_2301,N_2429);
nor U2664 (N_2664,N_2305,N_2340);
nor U2665 (N_2665,N_2018,N_2069);
nand U2666 (N_2666,N_2210,N_2195);
nand U2667 (N_2667,N_2133,N_2160);
nor U2668 (N_2668,N_2128,N_2035);
nand U2669 (N_2669,N_2042,N_2123);
or U2670 (N_2670,N_2184,N_2237);
nor U2671 (N_2671,N_2447,N_2109);
and U2672 (N_2672,N_2056,N_2423);
or U2673 (N_2673,N_2099,N_2277);
and U2674 (N_2674,N_2291,N_2214);
xor U2675 (N_2675,N_2279,N_2070);
nor U2676 (N_2676,N_2088,N_2098);
and U2677 (N_2677,N_2076,N_2213);
or U2678 (N_2678,N_2117,N_2002);
or U2679 (N_2679,N_2441,N_2092);
and U2680 (N_2680,N_2391,N_2382);
and U2681 (N_2681,N_2438,N_2009);
nand U2682 (N_2682,N_2364,N_2058);
and U2683 (N_2683,N_2460,N_2388);
or U2684 (N_2684,N_2055,N_2326);
or U2685 (N_2685,N_2155,N_2178);
or U2686 (N_2686,N_2127,N_2334);
and U2687 (N_2687,N_2463,N_2487);
nand U2688 (N_2688,N_2261,N_2034);
nand U2689 (N_2689,N_2192,N_2224);
and U2690 (N_2690,N_2306,N_2003);
nand U2691 (N_2691,N_2287,N_2110);
and U2692 (N_2692,N_2169,N_2062);
and U2693 (N_2693,N_2398,N_2194);
and U2694 (N_2694,N_2446,N_2285);
nor U2695 (N_2695,N_2384,N_2499);
nor U2696 (N_2696,N_2152,N_2339);
xnor U2697 (N_2697,N_2310,N_2324);
or U2698 (N_2698,N_2389,N_2290);
or U2699 (N_2699,N_2078,N_2497);
nand U2700 (N_2700,N_2017,N_2481);
nand U2701 (N_2701,N_2240,N_2437);
and U2702 (N_2702,N_2478,N_2397);
nor U2703 (N_2703,N_2130,N_2410);
nand U2704 (N_2704,N_2280,N_2241);
nand U2705 (N_2705,N_2403,N_2119);
nand U2706 (N_2706,N_2264,N_2322);
and U2707 (N_2707,N_2490,N_2170);
or U2708 (N_2708,N_2488,N_2124);
and U2709 (N_2709,N_2233,N_2267);
or U2710 (N_2710,N_2146,N_2298);
nand U2711 (N_2711,N_2349,N_2335);
and U2712 (N_2712,N_2140,N_2432);
nand U2713 (N_2713,N_2141,N_2288);
nand U2714 (N_2714,N_2315,N_2179);
nor U2715 (N_2715,N_2359,N_2345);
nor U2716 (N_2716,N_2221,N_2186);
nor U2717 (N_2717,N_2415,N_2296);
nor U2718 (N_2718,N_2477,N_2485);
nor U2719 (N_2719,N_2215,N_2093);
or U2720 (N_2720,N_2260,N_2033);
and U2721 (N_2721,N_2482,N_2113);
and U2722 (N_2722,N_2052,N_2050);
nor U2723 (N_2723,N_2320,N_2417);
nand U2724 (N_2724,N_2366,N_2077);
and U2725 (N_2725,N_2426,N_2054);
nand U2726 (N_2726,N_2450,N_2200);
nand U2727 (N_2727,N_2263,N_2459);
and U2728 (N_2728,N_2104,N_2231);
or U2729 (N_2729,N_2286,N_2284);
nor U2730 (N_2730,N_2361,N_2148);
or U2731 (N_2731,N_2019,N_2375);
and U2732 (N_2732,N_2351,N_2040);
xor U2733 (N_2733,N_2080,N_2145);
or U2734 (N_2734,N_2247,N_2053);
nand U2735 (N_2735,N_2171,N_2239);
or U2736 (N_2736,N_2164,N_2188);
or U2737 (N_2737,N_2207,N_2255);
and U2738 (N_2738,N_2400,N_2016);
and U2739 (N_2739,N_2150,N_2406);
and U2740 (N_2740,N_2336,N_2068);
nand U2741 (N_2741,N_2471,N_2385);
nor U2742 (N_2742,N_2163,N_2464);
and U2743 (N_2743,N_2353,N_2492);
nor U2744 (N_2744,N_2274,N_2254);
and U2745 (N_2745,N_2242,N_2269);
nor U2746 (N_2746,N_2480,N_2201);
nor U2747 (N_2747,N_2131,N_2111);
and U2748 (N_2748,N_2031,N_2065);
or U2749 (N_2749,N_2292,N_2424);
nand U2750 (N_2750,N_2198,N_2461);
nor U2751 (N_2751,N_2215,N_2497);
or U2752 (N_2752,N_2106,N_2431);
and U2753 (N_2753,N_2278,N_2038);
nor U2754 (N_2754,N_2173,N_2280);
nand U2755 (N_2755,N_2228,N_2224);
and U2756 (N_2756,N_2121,N_2000);
nor U2757 (N_2757,N_2257,N_2065);
nor U2758 (N_2758,N_2088,N_2400);
nor U2759 (N_2759,N_2185,N_2006);
nor U2760 (N_2760,N_2051,N_2437);
nor U2761 (N_2761,N_2346,N_2056);
and U2762 (N_2762,N_2359,N_2116);
nand U2763 (N_2763,N_2000,N_2138);
nand U2764 (N_2764,N_2252,N_2022);
nor U2765 (N_2765,N_2268,N_2269);
nor U2766 (N_2766,N_2411,N_2498);
and U2767 (N_2767,N_2260,N_2177);
nor U2768 (N_2768,N_2137,N_2461);
and U2769 (N_2769,N_2268,N_2043);
and U2770 (N_2770,N_2033,N_2036);
xnor U2771 (N_2771,N_2283,N_2428);
nand U2772 (N_2772,N_2342,N_2402);
or U2773 (N_2773,N_2131,N_2412);
nand U2774 (N_2774,N_2325,N_2336);
and U2775 (N_2775,N_2456,N_2051);
nand U2776 (N_2776,N_2434,N_2177);
and U2777 (N_2777,N_2490,N_2428);
and U2778 (N_2778,N_2345,N_2062);
and U2779 (N_2779,N_2122,N_2325);
or U2780 (N_2780,N_2336,N_2129);
nor U2781 (N_2781,N_2125,N_2137);
and U2782 (N_2782,N_2166,N_2123);
nand U2783 (N_2783,N_2173,N_2363);
or U2784 (N_2784,N_2450,N_2383);
or U2785 (N_2785,N_2088,N_2421);
nand U2786 (N_2786,N_2067,N_2028);
and U2787 (N_2787,N_2371,N_2290);
nand U2788 (N_2788,N_2248,N_2345);
xor U2789 (N_2789,N_2447,N_2278);
nand U2790 (N_2790,N_2335,N_2060);
nand U2791 (N_2791,N_2466,N_2311);
or U2792 (N_2792,N_2143,N_2218);
or U2793 (N_2793,N_2425,N_2417);
and U2794 (N_2794,N_2125,N_2129);
and U2795 (N_2795,N_2112,N_2279);
or U2796 (N_2796,N_2179,N_2135);
nand U2797 (N_2797,N_2269,N_2029);
nand U2798 (N_2798,N_2400,N_2471);
nand U2799 (N_2799,N_2060,N_2176);
and U2800 (N_2800,N_2318,N_2229);
nand U2801 (N_2801,N_2236,N_2120);
nand U2802 (N_2802,N_2195,N_2483);
nor U2803 (N_2803,N_2498,N_2402);
or U2804 (N_2804,N_2079,N_2455);
nand U2805 (N_2805,N_2122,N_2356);
nand U2806 (N_2806,N_2048,N_2152);
nor U2807 (N_2807,N_2348,N_2105);
or U2808 (N_2808,N_2133,N_2013);
nand U2809 (N_2809,N_2365,N_2260);
and U2810 (N_2810,N_2247,N_2062);
nor U2811 (N_2811,N_2068,N_2331);
and U2812 (N_2812,N_2158,N_2252);
or U2813 (N_2813,N_2133,N_2227);
and U2814 (N_2814,N_2195,N_2352);
or U2815 (N_2815,N_2116,N_2234);
nor U2816 (N_2816,N_2079,N_2327);
and U2817 (N_2817,N_2488,N_2268);
nor U2818 (N_2818,N_2266,N_2092);
and U2819 (N_2819,N_2127,N_2308);
nor U2820 (N_2820,N_2475,N_2343);
or U2821 (N_2821,N_2181,N_2312);
nor U2822 (N_2822,N_2439,N_2340);
nor U2823 (N_2823,N_2156,N_2270);
nand U2824 (N_2824,N_2473,N_2242);
and U2825 (N_2825,N_2209,N_2025);
nand U2826 (N_2826,N_2170,N_2400);
nor U2827 (N_2827,N_2496,N_2147);
and U2828 (N_2828,N_2144,N_2127);
nand U2829 (N_2829,N_2478,N_2283);
nand U2830 (N_2830,N_2418,N_2111);
nand U2831 (N_2831,N_2336,N_2314);
nand U2832 (N_2832,N_2211,N_2389);
nor U2833 (N_2833,N_2365,N_2355);
nand U2834 (N_2834,N_2371,N_2085);
or U2835 (N_2835,N_2148,N_2261);
nor U2836 (N_2836,N_2015,N_2174);
nand U2837 (N_2837,N_2305,N_2005);
or U2838 (N_2838,N_2184,N_2022);
and U2839 (N_2839,N_2332,N_2169);
nor U2840 (N_2840,N_2217,N_2407);
and U2841 (N_2841,N_2001,N_2036);
nor U2842 (N_2842,N_2348,N_2326);
or U2843 (N_2843,N_2259,N_2080);
nor U2844 (N_2844,N_2470,N_2229);
or U2845 (N_2845,N_2142,N_2237);
and U2846 (N_2846,N_2009,N_2422);
or U2847 (N_2847,N_2137,N_2422);
or U2848 (N_2848,N_2326,N_2108);
or U2849 (N_2849,N_2486,N_2098);
and U2850 (N_2850,N_2231,N_2143);
nor U2851 (N_2851,N_2013,N_2095);
and U2852 (N_2852,N_2348,N_2087);
nand U2853 (N_2853,N_2024,N_2169);
and U2854 (N_2854,N_2318,N_2365);
and U2855 (N_2855,N_2104,N_2425);
nand U2856 (N_2856,N_2012,N_2415);
or U2857 (N_2857,N_2100,N_2181);
and U2858 (N_2858,N_2394,N_2359);
xor U2859 (N_2859,N_2365,N_2129);
nand U2860 (N_2860,N_2328,N_2495);
and U2861 (N_2861,N_2488,N_2199);
nand U2862 (N_2862,N_2015,N_2283);
nand U2863 (N_2863,N_2190,N_2109);
and U2864 (N_2864,N_2311,N_2297);
or U2865 (N_2865,N_2323,N_2377);
nand U2866 (N_2866,N_2077,N_2250);
nand U2867 (N_2867,N_2251,N_2033);
or U2868 (N_2868,N_2453,N_2438);
nor U2869 (N_2869,N_2475,N_2094);
nor U2870 (N_2870,N_2060,N_2437);
or U2871 (N_2871,N_2091,N_2237);
nor U2872 (N_2872,N_2045,N_2074);
and U2873 (N_2873,N_2109,N_2403);
xnor U2874 (N_2874,N_2010,N_2478);
and U2875 (N_2875,N_2012,N_2257);
nand U2876 (N_2876,N_2496,N_2138);
nand U2877 (N_2877,N_2176,N_2356);
and U2878 (N_2878,N_2171,N_2306);
or U2879 (N_2879,N_2177,N_2499);
nor U2880 (N_2880,N_2414,N_2391);
or U2881 (N_2881,N_2449,N_2166);
or U2882 (N_2882,N_2241,N_2474);
nand U2883 (N_2883,N_2193,N_2407);
and U2884 (N_2884,N_2374,N_2186);
nand U2885 (N_2885,N_2149,N_2473);
or U2886 (N_2886,N_2359,N_2024);
and U2887 (N_2887,N_2078,N_2276);
or U2888 (N_2888,N_2046,N_2068);
nor U2889 (N_2889,N_2232,N_2238);
or U2890 (N_2890,N_2273,N_2439);
or U2891 (N_2891,N_2391,N_2279);
or U2892 (N_2892,N_2228,N_2499);
nor U2893 (N_2893,N_2127,N_2035);
and U2894 (N_2894,N_2090,N_2451);
and U2895 (N_2895,N_2024,N_2053);
and U2896 (N_2896,N_2226,N_2228);
nor U2897 (N_2897,N_2066,N_2219);
or U2898 (N_2898,N_2147,N_2399);
nor U2899 (N_2899,N_2004,N_2029);
and U2900 (N_2900,N_2161,N_2198);
nor U2901 (N_2901,N_2311,N_2489);
or U2902 (N_2902,N_2325,N_2052);
nor U2903 (N_2903,N_2381,N_2160);
and U2904 (N_2904,N_2325,N_2400);
nand U2905 (N_2905,N_2136,N_2159);
nor U2906 (N_2906,N_2436,N_2180);
and U2907 (N_2907,N_2036,N_2202);
and U2908 (N_2908,N_2471,N_2384);
and U2909 (N_2909,N_2191,N_2177);
nor U2910 (N_2910,N_2461,N_2006);
xor U2911 (N_2911,N_2193,N_2304);
xor U2912 (N_2912,N_2211,N_2493);
nor U2913 (N_2913,N_2033,N_2418);
nand U2914 (N_2914,N_2303,N_2394);
and U2915 (N_2915,N_2176,N_2334);
nor U2916 (N_2916,N_2289,N_2020);
nand U2917 (N_2917,N_2293,N_2207);
xnor U2918 (N_2918,N_2006,N_2094);
and U2919 (N_2919,N_2068,N_2172);
nor U2920 (N_2920,N_2459,N_2351);
nand U2921 (N_2921,N_2286,N_2189);
nor U2922 (N_2922,N_2169,N_2089);
nand U2923 (N_2923,N_2103,N_2168);
nand U2924 (N_2924,N_2475,N_2044);
or U2925 (N_2925,N_2485,N_2085);
nand U2926 (N_2926,N_2469,N_2379);
or U2927 (N_2927,N_2381,N_2392);
nor U2928 (N_2928,N_2333,N_2346);
nor U2929 (N_2929,N_2235,N_2283);
and U2930 (N_2930,N_2074,N_2244);
and U2931 (N_2931,N_2312,N_2402);
and U2932 (N_2932,N_2218,N_2146);
and U2933 (N_2933,N_2059,N_2112);
or U2934 (N_2934,N_2054,N_2101);
or U2935 (N_2935,N_2238,N_2436);
nor U2936 (N_2936,N_2380,N_2283);
nand U2937 (N_2937,N_2131,N_2407);
and U2938 (N_2938,N_2347,N_2014);
and U2939 (N_2939,N_2070,N_2328);
nand U2940 (N_2940,N_2002,N_2473);
or U2941 (N_2941,N_2209,N_2462);
xor U2942 (N_2942,N_2068,N_2087);
nand U2943 (N_2943,N_2360,N_2472);
nand U2944 (N_2944,N_2438,N_2273);
or U2945 (N_2945,N_2230,N_2089);
and U2946 (N_2946,N_2004,N_2150);
nor U2947 (N_2947,N_2263,N_2170);
nand U2948 (N_2948,N_2343,N_2366);
nand U2949 (N_2949,N_2412,N_2188);
and U2950 (N_2950,N_2046,N_2290);
and U2951 (N_2951,N_2390,N_2069);
nand U2952 (N_2952,N_2455,N_2093);
nor U2953 (N_2953,N_2261,N_2227);
and U2954 (N_2954,N_2126,N_2391);
nor U2955 (N_2955,N_2199,N_2461);
xor U2956 (N_2956,N_2360,N_2116);
and U2957 (N_2957,N_2484,N_2058);
nor U2958 (N_2958,N_2033,N_2262);
or U2959 (N_2959,N_2242,N_2049);
and U2960 (N_2960,N_2391,N_2187);
or U2961 (N_2961,N_2277,N_2437);
or U2962 (N_2962,N_2296,N_2433);
nand U2963 (N_2963,N_2079,N_2476);
or U2964 (N_2964,N_2146,N_2421);
nand U2965 (N_2965,N_2029,N_2217);
and U2966 (N_2966,N_2457,N_2259);
nand U2967 (N_2967,N_2099,N_2338);
or U2968 (N_2968,N_2316,N_2166);
nor U2969 (N_2969,N_2492,N_2003);
and U2970 (N_2970,N_2416,N_2053);
nor U2971 (N_2971,N_2271,N_2122);
nand U2972 (N_2972,N_2064,N_2250);
and U2973 (N_2973,N_2235,N_2059);
nor U2974 (N_2974,N_2218,N_2487);
or U2975 (N_2975,N_2118,N_2385);
nor U2976 (N_2976,N_2459,N_2332);
nor U2977 (N_2977,N_2488,N_2240);
nor U2978 (N_2978,N_2355,N_2354);
and U2979 (N_2979,N_2489,N_2259);
or U2980 (N_2980,N_2376,N_2146);
nor U2981 (N_2981,N_2285,N_2357);
and U2982 (N_2982,N_2411,N_2032);
nand U2983 (N_2983,N_2255,N_2391);
nand U2984 (N_2984,N_2497,N_2438);
nor U2985 (N_2985,N_2026,N_2447);
or U2986 (N_2986,N_2184,N_2382);
nand U2987 (N_2987,N_2120,N_2191);
or U2988 (N_2988,N_2073,N_2411);
nor U2989 (N_2989,N_2129,N_2132);
or U2990 (N_2990,N_2411,N_2013);
or U2991 (N_2991,N_2247,N_2428);
nor U2992 (N_2992,N_2283,N_2061);
xnor U2993 (N_2993,N_2382,N_2433);
nand U2994 (N_2994,N_2154,N_2071);
nand U2995 (N_2995,N_2010,N_2142);
xor U2996 (N_2996,N_2027,N_2362);
or U2997 (N_2997,N_2229,N_2366);
nor U2998 (N_2998,N_2199,N_2454);
and U2999 (N_2999,N_2289,N_2324);
or UO_0 (O_0,N_2534,N_2914);
or UO_1 (O_1,N_2814,N_2788);
or UO_2 (O_2,N_2838,N_2915);
nand UO_3 (O_3,N_2620,N_2904);
nand UO_4 (O_4,N_2727,N_2679);
nand UO_5 (O_5,N_2592,N_2665);
nand UO_6 (O_6,N_2930,N_2943);
or UO_7 (O_7,N_2673,N_2526);
or UO_8 (O_8,N_2618,N_2846);
nor UO_9 (O_9,N_2567,N_2580);
nand UO_10 (O_10,N_2529,N_2722);
and UO_11 (O_11,N_2571,N_2530);
nor UO_12 (O_12,N_2718,N_2994);
nor UO_13 (O_13,N_2608,N_2664);
or UO_14 (O_14,N_2570,N_2585);
or UO_15 (O_15,N_2503,N_2968);
nand UO_16 (O_16,N_2791,N_2746);
and UO_17 (O_17,N_2985,N_2852);
nor UO_18 (O_18,N_2751,N_2825);
nor UO_19 (O_19,N_2785,N_2729);
or UO_20 (O_20,N_2697,N_2986);
or UO_21 (O_21,N_2675,N_2654);
or UO_22 (O_22,N_2525,N_2945);
or UO_23 (O_23,N_2861,N_2980);
and UO_24 (O_24,N_2738,N_2784);
and UO_25 (O_25,N_2623,N_2647);
nand UO_26 (O_26,N_2900,N_2541);
or UO_27 (O_27,N_2556,N_2715);
and UO_28 (O_28,N_2912,N_2781);
nand UO_29 (O_29,N_2737,N_2828);
nor UO_30 (O_30,N_2750,N_2509);
and UO_31 (O_31,N_2759,N_2822);
and UO_32 (O_32,N_2579,N_2857);
or UO_33 (O_33,N_2917,N_2682);
nand UO_34 (O_34,N_2862,N_2535);
nor UO_35 (O_35,N_2764,N_2850);
or UO_36 (O_36,N_2868,N_2504);
nand UO_37 (O_37,N_2680,N_2650);
nor UO_38 (O_38,N_2616,N_2820);
or UO_39 (O_39,N_2954,N_2991);
nor UO_40 (O_40,N_2979,N_2905);
nor UO_41 (O_41,N_2578,N_2693);
and UO_42 (O_42,N_2907,N_2593);
xnor UO_43 (O_43,N_2990,N_2925);
xor UO_44 (O_44,N_2830,N_2835);
or UO_45 (O_45,N_2829,N_2603);
and UO_46 (O_46,N_2753,N_2630);
xnor UO_47 (O_47,N_2500,N_2543);
nor UO_48 (O_48,N_2709,N_2842);
or UO_49 (O_49,N_2783,N_2634);
nand UO_50 (O_50,N_2841,N_2872);
or UO_51 (O_51,N_2600,N_2644);
and UO_52 (O_52,N_2594,N_2720);
and UO_53 (O_53,N_2707,N_2596);
nor UO_54 (O_54,N_2811,N_2839);
nor UO_55 (O_55,N_2663,N_2652);
nor UO_56 (O_56,N_2812,N_2807);
nor UO_57 (O_57,N_2657,N_2798);
nor UO_58 (O_58,N_2695,N_2642);
or UO_59 (O_59,N_2937,N_2649);
and UO_60 (O_60,N_2810,N_2893);
or UO_61 (O_61,N_2996,N_2517);
and UO_62 (O_62,N_2871,N_2877);
nor UO_63 (O_63,N_2993,N_2684);
or UO_64 (O_64,N_2884,N_2779);
or UO_65 (O_65,N_2794,N_2774);
nand UO_66 (O_66,N_2832,N_2882);
nor UO_67 (O_67,N_2876,N_2554);
nand UO_68 (O_68,N_2523,N_2888);
and UO_69 (O_69,N_2683,N_2982);
nor UO_70 (O_70,N_2643,N_2706);
nor UO_71 (O_71,N_2582,N_2813);
or UO_72 (O_72,N_2598,N_2632);
and UO_73 (O_73,N_2628,N_2955);
or UO_74 (O_74,N_2676,N_2566);
nor UO_75 (O_75,N_2796,N_2615);
nand UO_76 (O_76,N_2799,N_2797);
nor UO_77 (O_77,N_2749,N_2855);
nor UO_78 (O_78,N_2723,N_2866);
nand UO_79 (O_79,N_2613,N_2671);
nand UO_80 (O_80,N_2775,N_2716);
xnor UO_81 (O_81,N_2790,N_2890);
and UO_82 (O_82,N_2919,N_2983);
and UO_83 (O_83,N_2694,N_2935);
nor UO_84 (O_84,N_2989,N_2896);
or UO_85 (O_85,N_2806,N_2653);
nor UO_86 (O_86,N_2562,N_2621);
and UO_87 (O_87,N_2553,N_2711);
nand UO_88 (O_88,N_2843,N_2856);
nor UO_89 (O_89,N_2988,N_2899);
or UO_90 (O_90,N_2924,N_2953);
nand UO_91 (O_91,N_2879,N_2769);
or UO_92 (O_92,N_2700,N_2538);
and UO_93 (O_93,N_2923,N_2815);
nand UO_94 (O_94,N_2655,N_2740);
nor UO_95 (O_95,N_2854,N_2560);
nor UO_96 (O_96,N_2837,N_2770);
nor UO_97 (O_97,N_2987,N_2959);
and UO_98 (O_98,N_2932,N_2974);
or UO_99 (O_99,N_2678,N_2635);
nor UO_100 (O_100,N_2691,N_2589);
nor UO_101 (O_101,N_2981,N_2966);
nand UO_102 (O_102,N_2614,N_2865);
or UO_103 (O_103,N_2817,N_2777);
nand UO_104 (O_104,N_2858,N_2913);
and UO_105 (O_105,N_2931,N_2920);
nand UO_106 (O_106,N_2611,N_2565);
nor UO_107 (O_107,N_2626,N_2548);
or UO_108 (O_108,N_2662,N_2631);
nor UO_109 (O_109,N_2638,N_2977);
xor UO_110 (O_110,N_2677,N_2940);
nor UO_111 (O_111,N_2909,N_2557);
nand UO_112 (O_112,N_2969,N_2995);
nor UO_113 (O_113,N_2933,N_2745);
or UO_114 (O_114,N_2659,N_2587);
and UO_115 (O_115,N_2946,N_2860);
and UO_116 (O_116,N_2629,N_2514);
and UO_117 (O_117,N_2942,N_2926);
nor UO_118 (O_118,N_2763,N_2533);
or UO_119 (O_119,N_2748,N_2586);
nor UO_120 (O_120,N_2521,N_2725);
xor UO_121 (O_121,N_2511,N_2771);
and UO_122 (O_122,N_2513,N_2941);
xor UO_123 (O_123,N_2609,N_2546);
nand UO_124 (O_124,N_2772,N_2658);
and UO_125 (O_125,N_2574,N_2801);
nor UO_126 (O_126,N_2692,N_2863);
nor UO_127 (O_127,N_2549,N_2532);
nand UO_128 (O_128,N_2961,N_2818);
nor UO_129 (O_129,N_2583,N_2809);
and UO_130 (O_130,N_2625,N_2767);
or UO_131 (O_131,N_2577,N_2889);
nor UO_132 (O_132,N_2765,N_2636);
xnor UO_133 (O_133,N_2536,N_2816);
nor UO_134 (O_134,N_2870,N_2540);
nor UO_135 (O_135,N_2502,N_2936);
or UO_136 (O_136,N_2528,N_2802);
or UO_137 (O_137,N_2964,N_2755);
nand UO_138 (O_138,N_2851,N_2610);
and UO_139 (O_139,N_2927,N_2756);
or UO_140 (O_140,N_2717,N_2782);
or UO_141 (O_141,N_2967,N_2522);
and UO_142 (O_142,N_2505,N_2833);
nand UO_143 (O_143,N_2681,N_2952);
and UO_144 (O_144,N_2508,N_2639);
nand UO_145 (O_145,N_2847,N_2708);
nand UO_146 (O_146,N_2510,N_2520);
nand UO_147 (O_147,N_2962,N_2971);
nor UO_148 (O_148,N_2768,N_2963);
nor UO_149 (O_149,N_2808,N_2958);
or UO_150 (O_150,N_2537,N_2997);
nor UO_151 (O_151,N_2805,N_2637);
or UO_152 (O_152,N_2702,N_2766);
nor UO_153 (O_153,N_2552,N_2688);
nor UO_154 (O_154,N_2894,N_2895);
nor UO_155 (O_155,N_2761,N_2878);
or UO_156 (O_156,N_2826,N_2595);
nand UO_157 (O_157,N_2827,N_2778);
and UO_158 (O_158,N_2760,N_2602);
nor UO_159 (O_159,N_2699,N_2823);
and UO_160 (O_160,N_2668,N_2640);
and UO_161 (O_161,N_2713,N_2624);
nor UO_162 (O_162,N_2641,N_2646);
and UO_163 (O_163,N_2892,N_2627);
and UO_164 (O_164,N_2864,N_2886);
nor UO_165 (O_165,N_2844,N_2800);
and UO_166 (O_166,N_2612,N_2950);
and UO_167 (O_167,N_2550,N_2922);
nor UO_168 (O_168,N_2859,N_2719);
nor UO_169 (O_169,N_2539,N_2795);
and UO_170 (O_170,N_2834,N_2992);
and UO_171 (O_171,N_2883,N_2617);
nand UO_172 (O_172,N_2584,N_2734);
or UO_173 (O_173,N_2604,N_2739);
nand UO_174 (O_174,N_2569,N_2531);
and UO_175 (O_175,N_2885,N_2726);
and UO_176 (O_176,N_2645,N_2733);
nor UO_177 (O_177,N_2921,N_2916);
and UO_178 (O_178,N_2696,N_2633);
or UO_179 (O_179,N_2831,N_2575);
nand UO_180 (O_180,N_2887,N_2527);
nand UO_181 (O_181,N_2910,N_2724);
nor UO_182 (O_182,N_2741,N_2948);
and UO_183 (O_183,N_2588,N_2545);
nor UO_184 (O_184,N_2880,N_2898);
nor UO_185 (O_185,N_2728,N_2957);
and UO_186 (O_186,N_2757,N_2901);
nand UO_187 (O_187,N_2564,N_2787);
and UO_188 (O_188,N_2978,N_2605);
or UO_189 (O_189,N_2874,N_2515);
nor UO_190 (O_190,N_2661,N_2558);
nand UO_191 (O_191,N_2845,N_2911);
nor UO_192 (O_192,N_2803,N_2929);
nor UO_193 (O_193,N_2875,N_2559);
nand UO_194 (O_194,N_2848,N_2591);
or UO_195 (O_195,N_2735,N_2999);
and UO_196 (O_196,N_2572,N_2918);
nor UO_197 (O_197,N_2908,N_2998);
and UO_198 (O_198,N_2744,N_2551);
nor UO_199 (O_199,N_2840,N_2732);
or UO_200 (O_200,N_2747,N_2576);
or UO_201 (O_201,N_2789,N_2542);
nor UO_202 (O_202,N_2975,N_2712);
nor UO_203 (O_203,N_2524,N_2824);
or UO_204 (O_204,N_2599,N_2573);
or UO_205 (O_205,N_2601,N_2849);
nand UO_206 (O_206,N_2897,N_2970);
or UO_207 (O_207,N_2731,N_2786);
nor UO_208 (O_208,N_2506,N_2972);
and UO_209 (O_209,N_2867,N_2973);
nor UO_210 (O_210,N_2976,N_2891);
or UO_211 (O_211,N_2581,N_2698);
nor UO_212 (O_212,N_2721,N_2780);
and UO_213 (O_213,N_2518,N_2561);
nand UO_214 (O_214,N_2701,N_2516);
or UO_215 (O_215,N_2507,N_2776);
nand UO_216 (O_216,N_2519,N_2821);
nand UO_217 (O_217,N_2666,N_2686);
nor UO_218 (O_218,N_2705,N_2669);
and UO_219 (O_219,N_2674,N_2793);
and UO_220 (O_220,N_2670,N_2689);
and UO_221 (O_221,N_2944,N_2906);
nor UO_222 (O_222,N_2881,N_2710);
nand UO_223 (O_223,N_2902,N_2622);
or UO_224 (O_224,N_2597,N_2730);
or UO_225 (O_225,N_2547,N_2960);
xor UO_226 (O_226,N_2690,N_2934);
nand UO_227 (O_227,N_2853,N_2949);
nand UO_228 (O_228,N_2714,N_2965);
and UO_229 (O_229,N_2687,N_2555);
and UO_230 (O_230,N_2568,N_2754);
or UO_231 (O_231,N_2869,N_2752);
nand UO_232 (O_232,N_2736,N_2607);
and UO_233 (O_233,N_2656,N_2704);
or UO_234 (O_234,N_2951,N_2563);
nand UO_235 (O_235,N_2619,N_2873);
and UO_236 (O_236,N_2956,N_2743);
or UO_237 (O_237,N_2939,N_2651);
nand UO_238 (O_238,N_2544,N_2938);
or UO_239 (O_239,N_2660,N_2947);
or UO_240 (O_240,N_2685,N_2742);
nor UO_241 (O_241,N_2590,N_2819);
and UO_242 (O_242,N_2903,N_2792);
or UO_243 (O_243,N_2667,N_2928);
nand UO_244 (O_244,N_2758,N_2606);
or UO_245 (O_245,N_2836,N_2762);
and UO_246 (O_246,N_2984,N_2773);
nor UO_247 (O_247,N_2501,N_2672);
or UO_248 (O_248,N_2703,N_2804);
and UO_249 (O_249,N_2648,N_2512);
xnor UO_250 (O_250,N_2792,N_2800);
nand UO_251 (O_251,N_2517,N_2727);
and UO_252 (O_252,N_2865,N_2676);
or UO_253 (O_253,N_2612,N_2609);
nand UO_254 (O_254,N_2689,N_2758);
nor UO_255 (O_255,N_2805,N_2986);
xnor UO_256 (O_256,N_2503,N_2932);
and UO_257 (O_257,N_2745,N_2621);
or UO_258 (O_258,N_2802,N_2702);
and UO_259 (O_259,N_2581,N_2575);
and UO_260 (O_260,N_2919,N_2623);
nor UO_261 (O_261,N_2777,N_2583);
and UO_262 (O_262,N_2782,N_2999);
nand UO_263 (O_263,N_2629,N_2651);
and UO_264 (O_264,N_2517,N_2512);
nor UO_265 (O_265,N_2672,N_2990);
and UO_266 (O_266,N_2553,N_2870);
nor UO_267 (O_267,N_2633,N_2712);
and UO_268 (O_268,N_2726,N_2796);
nand UO_269 (O_269,N_2748,N_2735);
or UO_270 (O_270,N_2921,N_2551);
xor UO_271 (O_271,N_2662,N_2873);
nor UO_272 (O_272,N_2871,N_2924);
or UO_273 (O_273,N_2825,N_2652);
or UO_274 (O_274,N_2877,N_2825);
nor UO_275 (O_275,N_2677,N_2844);
nor UO_276 (O_276,N_2965,N_2908);
or UO_277 (O_277,N_2820,N_2954);
and UO_278 (O_278,N_2584,N_2515);
and UO_279 (O_279,N_2573,N_2541);
or UO_280 (O_280,N_2875,N_2880);
and UO_281 (O_281,N_2943,N_2884);
xnor UO_282 (O_282,N_2959,N_2531);
or UO_283 (O_283,N_2661,N_2557);
or UO_284 (O_284,N_2856,N_2846);
nand UO_285 (O_285,N_2890,N_2827);
nor UO_286 (O_286,N_2613,N_2944);
or UO_287 (O_287,N_2814,N_2865);
and UO_288 (O_288,N_2999,N_2998);
or UO_289 (O_289,N_2676,N_2635);
or UO_290 (O_290,N_2867,N_2548);
nand UO_291 (O_291,N_2512,N_2788);
xnor UO_292 (O_292,N_2600,N_2678);
nand UO_293 (O_293,N_2976,N_2580);
nand UO_294 (O_294,N_2532,N_2739);
nor UO_295 (O_295,N_2852,N_2799);
nand UO_296 (O_296,N_2795,N_2635);
xor UO_297 (O_297,N_2852,N_2862);
nor UO_298 (O_298,N_2771,N_2646);
and UO_299 (O_299,N_2854,N_2911);
nor UO_300 (O_300,N_2957,N_2725);
and UO_301 (O_301,N_2934,N_2616);
xnor UO_302 (O_302,N_2994,N_2719);
nor UO_303 (O_303,N_2529,N_2787);
xnor UO_304 (O_304,N_2504,N_2991);
nor UO_305 (O_305,N_2761,N_2774);
or UO_306 (O_306,N_2537,N_2526);
or UO_307 (O_307,N_2664,N_2846);
or UO_308 (O_308,N_2567,N_2535);
xor UO_309 (O_309,N_2535,N_2863);
and UO_310 (O_310,N_2649,N_2993);
nor UO_311 (O_311,N_2811,N_2616);
nor UO_312 (O_312,N_2717,N_2729);
and UO_313 (O_313,N_2903,N_2861);
or UO_314 (O_314,N_2935,N_2696);
nand UO_315 (O_315,N_2892,N_2684);
and UO_316 (O_316,N_2744,N_2913);
nor UO_317 (O_317,N_2873,N_2909);
or UO_318 (O_318,N_2859,N_2799);
nor UO_319 (O_319,N_2587,N_2730);
or UO_320 (O_320,N_2616,N_2544);
nor UO_321 (O_321,N_2818,N_2697);
nor UO_322 (O_322,N_2620,N_2872);
or UO_323 (O_323,N_2719,N_2955);
or UO_324 (O_324,N_2617,N_2714);
nand UO_325 (O_325,N_2661,N_2984);
or UO_326 (O_326,N_2804,N_2814);
nor UO_327 (O_327,N_2971,N_2918);
nor UO_328 (O_328,N_2645,N_2668);
nand UO_329 (O_329,N_2969,N_2832);
nand UO_330 (O_330,N_2763,N_2899);
and UO_331 (O_331,N_2754,N_2592);
and UO_332 (O_332,N_2922,N_2873);
or UO_333 (O_333,N_2769,N_2639);
or UO_334 (O_334,N_2618,N_2674);
nand UO_335 (O_335,N_2757,N_2730);
nand UO_336 (O_336,N_2693,N_2800);
or UO_337 (O_337,N_2999,N_2909);
nand UO_338 (O_338,N_2773,N_2715);
and UO_339 (O_339,N_2532,N_2577);
nand UO_340 (O_340,N_2965,N_2547);
or UO_341 (O_341,N_2929,N_2602);
or UO_342 (O_342,N_2841,N_2530);
nand UO_343 (O_343,N_2669,N_2652);
nand UO_344 (O_344,N_2729,N_2851);
or UO_345 (O_345,N_2918,N_2864);
nor UO_346 (O_346,N_2918,N_2639);
nor UO_347 (O_347,N_2859,N_2618);
nand UO_348 (O_348,N_2985,N_2776);
and UO_349 (O_349,N_2842,N_2523);
nor UO_350 (O_350,N_2802,N_2690);
nand UO_351 (O_351,N_2776,N_2789);
and UO_352 (O_352,N_2834,N_2709);
nand UO_353 (O_353,N_2788,N_2851);
nand UO_354 (O_354,N_2541,N_2733);
nor UO_355 (O_355,N_2802,N_2607);
or UO_356 (O_356,N_2705,N_2535);
nand UO_357 (O_357,N_2711,N_2754);
and UO_358 (O_358,N_2559,N_2737);
nor UO_359 (O_359,N_2508,N_2919);
nand UO_360 (O_360,N_2911,N_2877);
or UO_361 (O_361,N_2929,N_2795);
nor UO_362 (O_362,N_2515,N_2607);
or UO_363 (O_363,N_2902,N_2655);
nand UO_364 (O_364,N_2713,N_2812);
nand UO_365 (O_365,N_2878,N_2959);
and UO_366 (O_366,N_2811,N_2556);
nand UO_367 (O_367,N_2521,N_2914);
and UO_368 (O_368,N_2944,N_2544);
nor UO_369 (O_369,N_2754,N_2694);
or UO_370 (O_370,N_2697,N_2946);
or UO_371 (O_371,N_2504,N_2765);
nand UO_372 (O_372,N_2609,N_2936);
and UO_373 (O_373,N_2636,N_2808);
nand UO_374 (O_374,N_2593,N_2870);
or UO_375 (O_375,N_2551,N_2945);
nor UO_376 (O_376,N_2936,N_2875);
nand UO_377 (O_377,N_2658,N_2728);
and UO_378 (O_378,N_2884,N_2601);
nor UO_379 (O_379,N_2690,N_2610);
nor UO_380 (O_380,N_2515,N_2780);
and UO_381 (O_381,N_2768,N_2502);
or UO_382 (O_382,N_2524,N_2745);
nor UO_383 (O_383,N_2858,N_2787);
or UO_384 (O_384,N_2893,N_2638);
nor UO_385 (O_385,N_2706,N_2578);
nor UO_386 (O_386,N_2571,N_2583);
nand UO_387 (O_387,N_2624,N_2696);
and UO_388 (O_388,N_2925,N_2648);
or UO_389 (O_389,N_2800,N_2736);
or UO_390 (O_390,N_2509,N_2932);
nor UO_391 (O_391,N_2959,N_2619);
and UO_392 (O_392,N_2897,N_2504);
nand UO_393 (O_393,N_2800,N_2510);
and UO_394 (O_394,N_2764,N_2986);
xor UO_395 (O_395,N_2970,N_2760);
or UO_396 (O_396,N_2710,N_2627);
and UO_397 (O_397,N_2655,N_2939);
nand UO_398 (O_398,N_2822,N_2912);
or UO_399 (O_399,N_2510,N_2947);
and UO_400 (O_400,N_2818,N_2899);
or UO_401 (O_401,N_2977,N_2664);
or UO_402 (O_402,N_2938,N_2553);
nand UO_403 (O_403,N_2731,N_2887);
or UO_404 (O_404,N_2916,N_2558);
nand UO_405 (O_405,N_2767,N_2882);
nor UO_406 (O_406,N_2624,N_2682);
nand UO_407 (O_407,N_2594,N_2529);
and UO_408 (O_408,N_2510,N_2637);
and UO_409 (O_409,N_2585,N_2734);
nor UO_410 (O_410,N_2965,N_2639);
and UO_411 (O_411,N_2645,N_2933);
and UO_412 (O_412,N_2794,N_2711);
nor UO_413 (O_413,N_2726,N_2713);
and UO_414 (O_414,N_2577,N_2746);
or UO_415 (O_415,N_2867,N_2921);
and UO_416 (O_416,N_2670,N_2671);
nand UO_417 (O_417,N_2914,N_2855);
or UO_418 (O_418,N_2946,N_2809);
nor UO_419 (O_419,N_2980,N_2519);
and UO_420 (O_420,N_2550,N_2647);
and UO_421 (O_421,N_2925,N_2680);
nor UO_422 (O_422,N_2628,N_2992);
or UO_423 (O_423,N_2763,N_2907);
and UO_424 (O_424,N_2892,N_2569);
and UO_425 (O_425,N_2974,N_2961);
xor UO_426 (O_426,N_2999,N_2917);
and UO_427 (O_427,N_2728,N_2644);
nand UO_428 (O_428,N_2726,N_2540);
or UO_429 (O_429,N_2740,N_2861);
nor UO_430 (O_430,N_2505,N_2572);
and UO_431 (O_431,N_2983,N_2788);
and UO_432 (O_432,N_2876,N_2799);
nand UO_433 (O_433,N_2539,N_2634);
nor UO_434 (O_434,N_2870,N_2601);
or UO_435 (O_435,N_2559,N_2967);
nor UO_436 (O_436,N_2572,N_2812);
nand UO_437 (O_437,N_2988,N_2808);
nand UO_438 (O_438,N_2696,N_2625);
and UO_439 (O_439,N_2555,N_2533);
or UO_440 (O_440,N_2603,N_2595);
and UO_441 (O_441,N_2898,N_2837);
nor UO_442 (O_442,N_2967,N_2744);
nor UO_443 (O_443,N_2784,N_2934);
nand UO_444 (O_444,N_2527,N_2896);
nor UO_445 (O_445,N_2728,N_2742);
and UO_446 (O_446,N_2916,N_2630);
nand UO_447 (O_447,N_2873,N_2750);
and UO_448 (O_448,N_2974,N_2846);
and UO_449 (O_449,N_2816,N_2833);
nand UO_450 (O_450,N_2851,N_2594);
nand UO_451 (O_451,N_2918,N_2949);
nor UO_452 (O_452,N_2798,N_2855);
nand UO_453 (O_453,N_2932,N_2870);
and UO_454 (O_454,N_2890,N_2721);
nor UO_455 (O_455,N_2731,N_2895);
and UO_456 (O_456,N_2631,N_2526);
or UO_457 (O_457,N_2856,N_2748);
nand UO_458 (O_458,N_2603,N_2553);
nand UO_459 (O_459,N_2707,N_2870);
nor UO_460 (O_460,N_2792,N_2664);
and UO_461 (O_461,N_2938,N_2955);
and UO_462 (O_462,N_2793,N_2527);
and UO_463 (O_463,N_2748,N_2514);
nor UO_464 (O_464,N_2655,N_2774);
nor UO_465 (O_465,N_2946,N_2626);
and UO_466 (O_466,N_2805,N_2748);
xor UO_467 (O_467,N_2985,N_2987);
and UO_468 (O_468,N_2702,N_2989);
or UO_469 (O_469,N_2841,N_2824);
nand UO_470 (O_470,N_2522,N_2850);
and UO_471 (O_471,N_2868,N_2513);
nand UO_472 (O_472,N_2664,N_2748);
or UO_473 (O_473,N_2883,N_2518);
and UO_474 (O_474,N_2719,N_2925);
nand UO_475 (O_475,N_2635,N_2870);
or UO_476 (O_476,N_2587,N_2958);
and UO_477 (O_477,N_2943,N_2979);
nor UO_478 (O_478,N_2843,N_2522);
or UO_479 (O_479,N_2537,N_2916);
nor UO_480 (O_480,N_2569,N_2528);
and UO_481 (O_481,N_2617,N_2600);
nor UO_482 (O_482,N_2943,N_2987);
or UO_483 (O_483,N_2661,N_2631);
and UO_484 (O_484,N_2629,N_2821);
nand UO_485 (O_485,N_2602,N_2861);
and UO_486 (O_486,N_2791,N_2830);
or UO_487 (O_487,N_2663,N_2639);
nor UO_488 (O_488,N_2875,N_2634);
or UO_489 (O_489,N_2820,N_2749);
and UO_490 (O_490,N_2904,N_2962);
and UO_491 (O_491,N_2613,N_2691);
and UO_492 (O_492,N_2675,N_2806);
or UO_493 (O_493,N_2921,N_2909);
xor UO_494 (O_494,N_2618,N_2796);
nand UO_495 (O_495,N_2861,N_2608);
nor UO_496 (O_496,N_2976,N_2876);
and UO_497 (O_497,N_2912,N_2747);
nand UO_498 (O_498,N_2652,N_2922);
and UO_499 (O_499,N_2980,N_2578);
endmodule