module basic_1000_10000_1500_4_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_517,In_87);
or U1 (N_1,In_146,In_625);
nor U2 (N_2,In_643,In_954);
nand U3 (N_3,In_333,In_201);
nor U4 (N_4,In_335,In_642);
nand U5 (N_5,In_327,In_399);
nor U6 (N_6,In_733,In_186);
nand U7 (N_7,In_614,In_840);
and U8 (N_8,In_653,In_216);
nand U9 (N_9,In_727,In_210);
nor U10 (N_10,In_279,In_801);
and U11 (N_11,In_139,In_77);
and U12 (N_12,In_332,In_483);
or U13 (N_13,In_376,In_773);
or U14 (N_14,In_678,In_549);
or U15 (N_15,In_97,In_177);
and U16 (N_16,In_401,In_853);
or U17 (N_17,In_930,In_35);
or U18 (N_18,In_408,In_121);
nand U19 (N_19,In_405,In_809);
or U20 (N_20,In_576,In_786);
or U21 (N_21,In_981,In_771);
or U22 (N_22,In_388,In_346);
or U23 (N_23,In_626,In_822);
and U24 (N_24,In_639,In_808);
and U25 (N_25,In_648,In_235);
nand U26 (N_26,In_334,In_63);
nand U27 (N_27,In_607,In_212);
nor U28 (N_28,In_883,In_416);
or U29 (N_29,In_652,In_925);
nand U30 (N_30,In_159,In_852);
nand U31 (N_31,In_932,In_162);
nor U32 (N_32,In_444,In_238);
and U33 (N_33,In_963,In_385);
nor U34 (N_34,In_606,In_454);
xnor U35 (N_35,In_521,In_857);
or U36 (N_36,In_179,In_716);
nor U37 (N_37,In_326,In_762);
nor U38 (N_38,In_738,In_861);
nor U39 (N_39,In_383,In_609);
nor U40 (N_40,In_403,In_116);
nand U41 (N_41,In_537,In_126);
nand U42 (N_42,In_310,In_608);
or U43 (N_43,In_95,In_331);
and U44 (N_44,In_568,In_158);
nor U45 (N_45,In_353,In_223);
and U46 (N_46,In_338,In_236);
nor U47 (N_47,In_898,In_93);
nand U48 (N_48,In_835,In_191);
and U49 (N_49,In_205,In_390);
or U50 (N_50,In_277,In_770);
and U51 (N_51,In_763,In_344);
nand U52 (N_52,In_305,In_661);
xnor U53 (N_53,In_410,In_24);
or U54 (N_54,In_744,In_800);
nand U55 (N_55,In_303,In_511);
nand U56 (N_56,In_708,In_970);
or U57 (N_57,In_739,In_50);
nor U58 (N_58,In_219,In_623);
and U59 (N_59,In_990,In_402);
xnor U60 (N_60,In_151,In_282);
nand U61 (N_61,In_718,In_90);
nor U62 (N_62,In_681,In_544);
xnor U63 (N_63,In_901,In_688);
nand U64 (N_64,In_315,In_47);
and U65 (N_65,In_182,In_971);
nor U66 (N_66,In_847,In_479);
nor U67 (N_67,In_664,In_547);
or U68 (N_68,In_706,In_381);
and U69 (N_69,In_319,In_41);
or U70 (N_70,In_977,In_695);
nor U71 (N_71,In_539,In_843);
nor U72 (N_72,In_314,In_341);
nor U73 (N_73,In_92,In_942);
nor U74 (N_74,In_972,In_580);
nor U75 (N_75,In_567,In_407);
nor U76 (N_76,In_218,In_839);
and U77 (N_77,In_197,In_409);
or U78 (N_78,In_188,In_468);
and U79 (N_79,In_329,In_0);
nor U80 (N_80,In_495,In_964);
xor U81 (N_81,In_730,In_242);
nor U82 (N_82,In_339,In_506);
nand U83 (N_83,In_306,In_968);
and U84 (N_84,In_224,In_435);
and U85 (N_85,In_293,In_904);
nand U86 (N_86,In_778,In_816);
and U87 (N_87,In_641,In_621);
and U88 (N_88,In_637,In_690);
and U89 (N_89,In_230,In_906);
nor U90 (N_90,In_138,In_507);
nand U91 (N_91,In_260,In_308);
or U92 (N_92,In_601,In_336);
nor U93 (N_93,In_854,In_119);
or U94 (N_94,In_307,In_784);
nand U95 (N_95,In_591,In_252);
nand U96 (N_96,In_464,In_323);
and U97 (N_97,In_328,In_848);
or U98 (N_98,In_802,In_991);
or U99 (N_99,In_161,In_225);
or U100 (N_100,In_792,In_183);
nand U101 (N_101,In_616,In_589);
nand U102 (N_102,In_562,In_470);
nor U103 (N_103,In_69,In_382);
nor U104 (N_104,In_714,In_190);
nand U105 (N_105,In_394,In_657);
or U106 (N_106,In_76,In_994);
nand U107 (N_107,In_553,In_206);
nor U108 (N_108,In_888,In_458);
nand U109 (N_109,In_819,In_563);
nand U110 (N_110,In_415,In_789);
or U111 (N_111,In_80,In_463);
nand U112 (N_112,In_987,In_540);
nand U113 (N_113,In_634,In_966);
nand U114 (N_114,In_115,In_742);
and U115 (N_115,In_4,In_747);
nor U116 (N_116,In_363,In_3);
or U117 (N_117,In_632,In_620);
or U118 (N_118,In_559,In_810);
nand U119 (N_119,In_500,In_665);
or U120 (N_120,In_297,In_579);
nand U121 (N_121,In_509,In_445);
and U122 (N_122,In_60,In_866);
or U123 (N_123,In_378,In_320);
or U124 (N_124,In_91,In_992);
or U125 (N_125,In_871,In_924);
xor U126 (N_126,In_68,In_803);
and U127 (N_127,In_174,In_325);
or U128 (N_128,In_476,In_575);
or U129 (N_129,In_952,In_419);
nand U130 (N_130,In_349,In_745);
and U131 (N_131,In_743,In_996);
and U132 (N_132,In_294,In_812);
nand U133 (N_133,In_831,In_268);
nand U134 (N_134,In_411,In_168);
nor U135 (N_135,In_550,In_709);
nor U136 (N_136,In_798,In_248);
or U137 (N_137,In_751,In_1);
and U138 (N_138,In_560,In_732);
and U139 (N_139,In_387,In_98);
or U140 (N_140,In_581,In_909);
or U141 (N_141,In_369,In_542);
and U142 (N_142,In_428,In_868);
nor U143 (N_143,In_937,In_460);
nand U144 (N_144,In_286,In_986);
or U145 (N_145,In_702,In_881);
nor U146 (N_146,In_112,In_176);
nor U147 (N_147,In_769,In_675);
nor U148 (N_148,In_25,In_102);
and U149 (N_149,In_828,In_259);
nor U150 (N_150,In_194,In_752);
nor U151 (N_151,In_392,In_198);
or U152 (N_152,In_185,In_720);
and U153 (N_153,In_100,In_489);
and U154 (N_154,In_467,In_677);
nor U155 (N_155,In_70,In_783);
nor U156 (N_156,In_42,In_239);
nor U157 (N_157,In_880,In_203);
and U158 (N_158,In_917,In_291);
nor U159 (N_159,In_75,In_719);
nor U160 (N_160,In_396,In_951);
xnor U161 (N_161,In_624,In_440);
nor U162 (N_162,In_271,In_955);
or U163 (N_163,In_113,In_322);
or U164 (N_164,In_189,In_250);
xnor U165 (N_165,In_241,In_572);
and U166 (N_166,In_386,In_790);
or U167 (N_167,In_377,In_967);
nand U168 (N_168,In_895,In_192);
and U169 (N_169,In_257,In_697);
and U170 (N_170,In_529,In_694);
or U171 (N_171,In_827,In_178);
or U172 (N_172,In_79,In_53);
or U173 (N_173,In_17,In_96);
nand U174 (N_174,In_753,In_232);
or U175 (N_175,In_525,In_358);
and U176 (N_176,In_842,In_873);
and U177 (N_177,In_469,In_774);
nor U178 (N_178,In_103,In_528);
nor U179 (N_179,In_958,In_214);
or U180 (N_180,In_820,In_143);
and U181 (N_181,In_131,In_81);
xor U182 (N_182,In_270,In_950);
or U183 (N_183,In_787,In_170);
and U184 (N_184,In_421,In_86);
or U185 (N_185,In_145,In_109);
xor U186 (N_186,In_56,In_599);
nor U187 (N_187,In_533,In_321);
and U188 (N_188,In_380,In_136);
and U189 (N_189,In_251,In_368);
nor U190 (N_190,In_582,In_947);
or U191 (N_191,In_459,In_863);
or U192 (N_192,In_826,In_106);
nand U193 (N_193,In_207,In_765);
nand U194 (N_194,In_748,In_775);
and U195 (N_195,In_493,In_518);
nor U196 (N_196,In_939,In_361);
or U197 (N_197,In_813,In_573);
or U198 (N_198,In_557,In_595);
and U199 (N_199,In_287,In_974);
nand U200 (N_200,In_299,In_920);
nand U201 (N_201,In_858,In_228);
nand U202 (N_202,In_759,In_619);
nand U203 (N_203,In_375,In_940);
nand U204 (N_204,In_788,In_655);
or U205 (N_205,In_683,In_737);
or U206 (N_206,In_267,In_202);
or U207 (N_207,In_477,In_125);
or U208 (N_208,In_348,In_546);
nand U209 (N_209,In_768,In_833);
or U210 (N_210,In_135,In_172);
or U211 (N_211,In_522,In_276);
nor U212 (N_212,In_806,In_215);
or U213 (N_213,In_141,In_622);
nand U214 (N_214,In_749,In_498);
nand U215 (N_215,In_905,In_231);
xor U216 (N_216,In_88,In_534);
and U217 (N_217,In_636,In_46);
or U218 (N_218,In_997,In_261);
and U219 (N_219,In_611,In_340);
or U220 (N_220,In_284,In_74);
or U221 (N_221,In_29,In_497);
or U222 (N_222,In_603,In_795);
and U223 (N_223,In_379,In_896);
nor U224 (N_224,In_275,In_903);
and U225 (N_225,In_5,In_957);
and U226 (N_226,In_564,In_627);
and U227 (N_227,In_577,In_233);
nand U228 (N_228,In_548,In_649);
and U229 (N_229,In_638,In_437);
and U230 (N_230,In_22,In_300);
nor U231 (N_231,In_443,In_501);
or U232 (N_232,In_911,In_860);
or U233 (N_233,In_628,In_561);
or U234 (N_234,In_961,In_82);
nand U235 (N_235,In_59,In_980);
nor U236 (N_236,In_384,In_166);
and U237 (N_237,In_650,In_587);
nand U238 (N_238,In_864,In_588);
or U239 (N_239,In_108,In_478);
nor U240 (N_240,In_885,In_360);
nand U241 (N_241,In_772,In_26);
nand U242 (N_242,In_491,In_89);
nand U243 (N_243,In_703,In_805);
or U244 (N_244,In_780,In_285);
nor U245 (N_245,In_44,In_845);
nor U246 (N_246,In_701,In_945);
nor U247 (N_247,In_565,In_395);
nor U248 (N_248,In_593,In_612);
and U249 (N_249,In_31,In_137);
nand U250 (N_250,In_566,In_21);
nand U251 (N_251,In_735,In_938);
nand U252 (N_252,In_696,In_281);
or U253 (N_253,In_6,In_691);
nand U254 (N_254,In_910,In_872);
and U255 (N_255,In_280,In_295);
or U256 (N_256,In_503,In_721);
or U257 (N_257,In_596,In_117);
or U258 (N_258,In_462,In_457);
nor U259 (N_259,In_400,In_269);
and U260 (N_260,In_58,In_640);
or U261 (N_261,In_631,In_766);
or U262 (N_262,In_337,In_584);
and U263 (N_263,In_290,In_508);
or U264 (N_264,In_309,In_258);
and U265 (N_265,In_425,In_555);
nor U266 (N_266,In_764,In_240);
and U267 (N_267,In_600,In_551);
or U268 (N_268,In_13,In_304);
nor U269 (N_269,In_935,In_273);
nand U270 (N_270,In_715,In_57);
nand U271 (N_271,In_776,In_254);
nor U272 (N_272,In_351,In_465);
nor U273 (N_273,In_558,In_374);
nand U274 (N_274,In_393,In_229);
nand U275 (N_275,In_645,In_148);
xnor U276 (N_276,In_510,In_931);
nand U277 (N_277,In_618,In_617);
and U278 (N_278,In_527,In_169);
and U279 (N_279,In_943,In_647);
nand U280 (N_280,In_278,In_919);
nor U281 (N_281,In_908,In_899);
and U282 (N_282,In_855,In_244);
nor U283 (N_283,In_673,In_480);
nand U284 (N_284,In_887,In_243);
or U285 (N_285,In_874,In_867);
or U286 (N_286,In_359,In_11);
or U287 (N_287,In_249,In_461);
or U288 (N_288,In_512,In_882);
nor U289 (N_289,In_36,In_760);
nor U290 (N_290,In_679,In_122);
nand U291 (N_291,In_536,In_976);
or U292 (N_292,In_959,In_513);
nand U293 (N_293,In_422,In_38);
nor U294 (N_294,In_700,In_797);
and U295 (N_295,In_844,In_756);
or U296 (N_296,In_451,In_571);
and U297 (N_297,In_535,In_123);
xnor U298 (N_298,In_181,In_414);
nor U299 (N_299,In_670,In_633);
and U300 (N_300,In_644,In_302);
nand U301 (N_301,In_757,In_111);
or U302 (N_302,In_916,In_605);
and U303 (N_303,In_418,In_133);
nor U304 (N_304,In_471,In_144);
and U305 (N_305,In_777,In_921);
or U306 (N_306,In_127,In_283);
nor U307 (N_307,In_167,In_61);
nor U308 (N_308,In_84,In_592);
nor U309 (N_309,In_2,In_985);
and U310 (N_310,In_902,In_312);
or U311 (N_311,In_496,In_362);
or U312 (N_312,In_372,In_472);
and U313 (N_313,In_825,In_175);
nand U314 (N_314,In_791,In_8);
nand U315 (N_315,In_318,In_693);
nor U316 (N_316,In_105,In_504);
nor U317 (N_317,In_978,In_492);
or U318 (N_318,In_519,In_481);
and U319 (N_319,In_204,In_969);
nand U320 (N_320,In_62,In_120);
and U321 (N_321,In_20,In_878);
nor U322 (N_322,In_484,In_729);
nor U323 (N_323,In_746,In_711);
or U324 (N_324,In_417,In_453);
nand U325 (N_325,In_824,In_545);
and U326 (N_326,In_707,In_862);
or U327 (N_327,In_10,In_33);
xnor U328 (N_328,In_993,In_66);
and U329 (N_329,In_934,In_473);
and U330 (N_330,In_629,In_264);
or U331 (N_331,In_211,In_12);
or U332 (N_332,In_821,In_505);
nand U333 (N_333,In_34,In_487);
nor U334 (N_334,In_686,In_823);
or U335 (N_335,In_953,In_927);
nand U336 (N_336,In_705,In_452);
and U337 (N_337,In_660,In_829);
xnor U338 (N_338,In_946,In_253);
or U339 (N_339,In_879,In_900);
nor U340 (N_340,In_962,In_274);
and U341 (N_341,In_54,In_973);
nand U342 (N_342,In_208,In_114);
nor U343 (N_343,In_171,In_30);
or U344 (N_344,In_893,In_140);
and U345 (N_345,In_865,In_32);
nand U346 (N_346,In_195,In_288);
nor U347 (N_347,In_569,In_897);
and U348 (N_348,In_779,In_884);
nand U349 (N_349,In_578,In_72);
nand U350 (N_350,In_814,In_134);
nand U351 (N_351,In_929,In_523);
nor U352 (N_352,In_687,In_907);
and U353 (N_353,In_941,In_441);
and U354 (N_354,In_426,In_193);
nor U355 (N_355,In_213,In_343);
xor U356 (N_356,In_164,In_439);
nand U357 (N_357,In_446,In_838);
and U358 (N_358,In_556,In_311);
nand U359 (N_359,In_658,In_153);
or U360 (N_360,In_289,In_364);
nor U361 (N_361,In_152,In_685);
or U362 (N_362,In_494,In_347);
and U363 (N_363,In_728,In_265);
nor U364 (N_364,In_846,In_9);
nand U365 (N_365,In_811,In_604);
and U366 (N_366,In_263,In_67);
nor U367 (N_367,In_350,In_531);
nand U368 (N_368,In_51,In_815);
nor U369 (N_369,In_856,In_796);
and U370 (N_370,In_52,In_936);
and U371 (N_371,In_45,In_667);
nor U372 (N_372,In_431,In_890);
nand U373 (N_373,In_914,In_710);
nor U374 (N_374,In_316,In_731);
nor U375 (N_375,In_433,In_324);
and U376 (N_376,In_982,In_704);
nor U377 (N_377,In_447,In_226);
and U378 (N_378,In_404,In_684);
or U379 (N_379,In_538,In_173);
nand U380 (N_380,In_94,In_196);
nor U381 (N_381,In_354,In_220);
nand U382 (N_382,In_163,In_16);
or U383 (N_383,In_654,In_948);
nand U384 (N_384,In_662,In_28);
and U385 (N_385,In_237,In_432);
nand U386 (N_386,In_656,In_761);
or U387 (N_387,In_64,In_412);
or U388 (N_388,In_984,In_398);
or U389 (N_389,In_184,In_357);
nand U390 (N_390,In_55,In_39);
nand U391 (N_391,In_475,In_317);
nor U392 (N_392,In_876,In_554);
or U393 (N_393,In_165,In_245);
xor U394 (N_394,In_574,In_912);
nand U395 (N_395,In_132,In_755);
or U396 (N_396,In_834,In_292);
and U397 (N_397,In_448,In_726);
nand U398 (N_398,In_541,In_875);
xor U399 (N_399,In_532,In_597);
nand U400 (N_400,In_246,In_296);
or U401 (N_401,In_692,In_486);
and U402 (N_402,In_758,In_150);
or U403 (N_403,In_222,In_355);
and U404 (N_404,In_7,In_983);
or U405 (N_405,In_723,In_979);
nor U406 (N_406,In_570,In_48);
nand U407 (N_407,In_998,In_602);
and U408 (N_408,In_502,In_147);
or U409 (N_409,In_450,In_869);
or U410 (N_410,In_836,In_23);
nand U411 (N_411,In_668,In_423);
nand U412 (N_412,In_156,In_674);
and U413 (N_413,In_850,In_712);
nand U414 (N_414,In_43,In_83);
and U415 (N_415,In_613,In_717);
or U416 (N_416,In_651,In_442);
and U417 (N_417,In_110,In_155);
xor U418 (N_418,In_741,In_157);
or U419 (N_419,In_19,In_975);
nand U420 (N_420,In_65,In_859);
nor U421 (N_421,In_73,In_734);
nand U422 (N_422,In_130,In_722);
nand U423 (N_423,In_27,In_516);
xnor U424 (N_424,In_988,In_200);
nor U425 (N_425,In_832,In_782);
and U426 (N_426,In_849,In_725);
and U427 (N_427,In_530,In_817);
nor U428 (N_428,In_799,In_456);
nand U429 (N_429,In_272,In_129);
nor U430 (N_430,In_365,In_101);
nor U431 (N_431,In_740,In_552);
and U432 (N_432,In_526,In_180);
nand U433 (N_433,In_913,In_750);
nor U434 (N_434,In_256,In_807);
nand U435 (N_435,In_71,In_352);
nor U436 (N_436,In_672,In_515);
or U437 (N_437,In_313,In_841);
and U438 (N_438,In_49,In_124);
and U439 (N_439,In_342,In_118);
nor U440 (N_440,In_520,In_995);
nand U441 (N_441,In_598,In_793);
and U442 (N_442,In_892,In_889);
or U443 (N_443,In_490,In_671);
nand U444 (N_444,In_37,In_666);
and U445 (N_445,In_356,In_713);
nand U446 (N_446,In_466,In_960);
or U447 (N_447,In_794,In_818);
nor U448 (N_448,In_999,In_455);
or U449 (N_449,In_676,In_370);
or U450 (N_450,In_754,In_199);
and U451 (N_451,In_221,In_434);
or U452 (N_452,In_689,In_965);
nor U453 (N_453,In_669,In_104);
and U454 (N_454,In_449,In_429);
or U455 (N_455,In_524,In_923);
or U456 (N_456,In_301,In_298);
nor U457 (N_457,In_956,In_18);
and U458 (N_458,In_78,In_781);
nand U459 (N_459,In_698,In_918);
or U460 (N_460,In_891,In_438);
or U461 (N_461,In_485,In_682);
nor U462 (N_462,In_989,In_590);
and U463 (N_463,In_851,In_262);
nand U464 (N_464,In_420,In_610);
or U465 (N_465,In_630,In_926);
nor U466 (N_466,In_474,In_85);
nand U467 (N_467,In_785,In_149);
nor U468 (N_468,In_870,In_389);
nor U469 (N_469,In_514,In_583);
nor U470 (N_470,In_436,In_40);
nand U471 (N_471,In_886,In_915);
nand U472 (N_472,In_837,In_736);
nor U473 (N_473,In_391,In_255);
and U474 (N_474,In_944,In_424);
or U475 (N_475,In_659,In_15);
nand U476 (N_476,In_767,In_949);
or U477 (N_477,In_877,In_594);
nand U478 (N_478,In_128,In_427);
or U479 (N_479,In_615,In_373);
nand U480 (N_480,In_894,In_247);
or U481 (N_481,In_830,In_406);
or U482 (N_482,In_724,In_266);
nor U483 (N_483,In_345,In_371);
nand U484 (N_484,In_160,In_699);
nand U485 (N_485,In_209,In_922);
nor U486 (N_486,In_585,In_154);
and U487 (N_487,In_635,In_234);
or U488 (N_488,In_330,In_663);
or U489 (N_489,In_107,In_366);
and U490 (N_490,In_367,In_499);
nor U491 (N_491,In_14,In_482);
nand U492 (N_492,In_99,In_413);
or U493 (N_493,In_804,In_488);
nand U494 (N_494,In_646,In_543);
and U495 (N_495,In_142,In_933);
or U496 (N_496,In_397,In_187);
nand U497 (N_497,In_217,In_928);
nand U498 (N_498,In_227,In_680);
or U499 (N_499,In_430,In_586);
nand U500 (N_500,In_419,In_92);
nand U501 (N_501,In_579,In_543);
nor U502 (N_502,In_868,In_304);
nor U503 (N_503,In_400,In_631);
nand U504 (N_504,In_526,In_745);
nand U505 (N_505,In_421,In_31);
nor U506 (N_506,In_627,In_135);
nand U507 (N_507,In_178,In_698);
nand U508 (N_508,In_958,In_346);
nand U509 (N_509,In_146,In_640);
and U510 (N_510,In_526,In_247);
nor U511 (N_511,In_665,In_156);
nand U512 (N_512,In_168,In_554);
and U513 (N_513,In_570,In_984);
nor U514 (N_514,In_960,In_144);
nand U515 (N_515,In_207,In_491);
and U516 (N_516,In_898,In_437);
nand U517 (N_517,In_407,In_965);
xor U518 (N_518,In_642,In_676);
and U519 (N_519,In_329,In_545);
or U520 (N_520,In_320,In_605);
and U521 (N_521,In_233,In_466);
or U522 (N_522,In_366,In_628);
nor U523 (N_523,In_886,In_933);
nand U524 (N_524,In_998,In_752);
and U525 (N_525,In_516,In_24);
nand U526 (N_526,In_938,In_181);
nand U527 (N_527,In_567,In_988);
or U528 (N_528,In_708,In_820);
and U529 (N_529,In_882,In_340);
nand U530 (N_530,In_495,In_913);
nor U531 (N_531,In_0,In_980);
nor U532 (N_532,In_360,In_660);
nand U533 (N_533,In_577,In_94);
or U534 (N_534,In_136,In_755);
and U535 (N_535,In_918,In_453);
and U536 (N_536,In_702,In_723);
nand U537 (N_537,In_95,In_935);
xor U538 (N_538,In_829,In_481);
or U539 (N_539,In_606,In_770);
nor U540 (N_540,In_871,In_978);
nor U541 (N_541,In_910,In_633);
nor U542 (N_542,In_943,In_37);
nor U543 (N_543,In_250,In_349);
and U544 (N_544,In_196,In_911);
or U545 (N_545,In_362,In_129);
nor U546 (N_546,In_606,In_536);
and U547 (N_547,In_960,In_283);
or U548 (N_548,In_705,In_325);
nor U549 (N_549,In_207,In_295);
nand U550 (N_550,In_97,In_981);
nand U551 (N_551,In_605,In_98);
nor U552 (N_552,In_798,In_134);
and U553 (N_553,In_810,In_362);
or U554 (N_554,In_24,In_651);
nor U555 (N_555,In_94,In_197);
nand U556 (N_556,In_234,In_725);
or U557 (N_557,In_823,In_185);
or U558 (N_558,In_487,In_763);
nand U559 (N_559,In_844,In_614);
and U560 (N_560,In_259,In_697);
or U561 (N_561,In_414,In_109);
and U562 (N_562,In_743,In_296);
nor U563 (N_563,In_387,In_220);
or U564 (N_564,In_440,In_179);
or U565 (N_565,In_24,In_565);
nor U566 (N_566,In_72,In_199);
or U567 (N_567,In_142,In_776);
nor U568 (N_568,In_277,In_823);
or U569 (N_569,In_258,In_431);
and U570 (N_570,In_982,In_277);
and U571 (N_571,In_960,In_494);
or U572 (N_572,In_94,In_850);
nand U573 (N_573,In_234,In_357);
or U574 (N_574,In_746,In_973);
nand U575 (N_575,In_633,In_512);
nor U576 (N_576,In_775,In_383);
nand U577 (N_577,In_921,In_545);
nand U578 (N_578,In_58,In_79);
nand U579 (N_579,In_300,In_509);
or U580 (N_580,In_723,In_892);
and U581 (N_581,In_245,In_378);
nand U582 (N_582,In_428,In_240);
or U583 (N_583,In_479,In_617);
xnor U584 (N_584,In_604,In_351);
or U585 (N_585,In_249,In_977);
nand U586 (N_586,In_812,In_549);
and U587 (N_587,In_874,In_945);
nand U588 (N_588,In_284,In_83);
and U589 (N_589,In_742,In_824);
or U590 (N_590,In_647,In_725);
or U591 (N_591,In_993,In_10);
and U592 (N_592,In_857,In_801);
and U593 (N_593,In_504,In_605);
or U594 (N_594,In_253,In_607);
and U595 (N_595,In_153,In_336);
or U596 (N_596,In_356,In_738);
and U597 (N_597,In_860,In_667);
and U598 (N_598,In_790,In_268);
or U599 (N_599,In_343,In_491);
nand U600 (N_600,In_298,In_139);
nor U601 (N_601,In_813,In_50);
nor U602 (N_602,In_564,In_804);
nor U603 (N_603,In_552,In_381);
and U604 (N_604,In_493,In_564);
and U605 (N_605,In_936,In_107);
or U606 (N_606,In_773,In_411);
or U607 (N_607,In_168,In_343);
or U608 (N_608,In_384,In_882);
nor U609 (N_609,In_821,In_724);
nor U610 (N_610,In_135,In_648);
nor U611 (N_611,In_351,In_28);
nand U612 (N_612,In_599,In_453);
nor U613 (N_613,In_908,In_672);
nor U614 (N_614,In_488,In_507);
nand U615 (N_615,In_938,In_820);
nor U616 (N_616,In_668,In_110);
or U617 (N_617,In_54,In_749);
nor U618 (N_618,In_543,In_252);
nand U619 (N_619,In_231,In_145);
or U620 (N_620,In_15,In_443);
nand U621 (N_621,In_465,In_314);
and U622 (N_622,In_822,In_951);
nand U623 (N_623,In_780,In_111);
nor U624 (N_624,In_361,In_12);
or U625 (N_625,In_843,In_842);
or U626 (N_626,In_578,In_213);
and U627 (N_627,In_62,In_931);
nor U628 (N_628,In_404,In_944);
nand U629 (N_629,In_904,In_810);
and U630 (N_630,In_12,In_792);
nand U631 (N_631,In_733,In_607);
nor U632 (N_632,In_296,In_700);
nand U633 (N_633,In_233,In_740);
and U634 (N_634,In_649,In_318);
or U635 (N_635,In_144,In_400);
and U636 (N_636,In_300,In_47);
and U637 (N_637,In_417,In_943);
nand U638 (N_638,In_618,In_897);
nand U639 (N_639,In_509,In_767);
and U640 (N_640,In_973,In_378);
nor U641 (N_641,In_398,In_721);
nand U642 (N_642,In_569,In_182);
or U643 (N_643,In_618,In_834);
nor U644 (N_644,In_240,In_619);
nand U645 (N_645,In_640,In_833);
and U646 (N_646,In_29,In_611);
nor U647 (N_647,In_990,In_413);
nor U648 (N_648,In_484,In_16);
nand U649 (N_649,In_739,In_983);
nand U650 (N_650,In_849,In_991);
nor U651 (N_651,In_470,In_574);
and U652 (N_652,In_194,In_628);
or U653 (N_653,In_386,In_399);
and U654 (N_654,In_200,In_890);
nand U655 (N_655,In_714,In_294);
nand U656 (N_656,In_407,In_937);
nor U657 (N_657,In_13,In_268);
or U658 (N_658,In_938,In_145);
nand U659 (N_659,In_594,In_124);
nor U660 (N_660,In_68,In_958);
nor U661 (N_661,In_664,In_727);
nor U662 (N_662,In_528,In_704);
or U663 (N_663,In_586,In_41);
nand U664 (N_664,In_1,In_916);
nand U665 (N_665,In_378,In_869);
and U666 (N_666,In_605,In_535);
or U667 (N_667,In_806,In_753);
nor U668 (N_668,In_796,In_447);
nor U669 (N_669,In_336,In_571);
nor U670 (N_670,In_331,In_152);
or U671 (N_671,In_741,In_252);
nand U672 (N_672,In_422,In_592);
nand U673 (N_673,In_45,In_165);
nand U674 (N_674,In_11,In_634);
nor U675 (N_675,In_934,In_904);
nor U676 (N_676,In_786,In_21);
nand U677 (N_677,In_324,In_346);
nand U678 (N_678,In_784,In_8);
or U679 (N_679,In_211,In_43);
nand U680 (N_680,In_690,In_635);
nor U681 (N_681,In_600,In_523);
nor U682 (N_682,In_306,In_659);
and U683 (N_683,In_315,In_74);
and U684 (N_684,In_639,In_217);
xnor U685 (N_685,In_652,In_717);
nor U686 (N_686,In_802,In_658);
and U687 (N_687,In_556,In_227);
nand U688 (N_688,In_29,In_934);
nand U689 (N_689,In_955,In_47);
nor U690 (N_690,In_840,In_911);
and U691 (N_691,In_773,In_986);
xnor U692 (N_692,In_215,In_181);
or U693 (N_693,In_792,In_400);
and U694 (N_694,In_562,In_944);
and U695 (N_695,In_138,In_64);
nor U696 (N_696,In_155,In_246);
nand U697 (N_697,In_772,In_38);
nand U698 (N_698,In_173,In_378);
nor U699 (N_699,In_216,In_268);
nor U700 (N_700,In_164,In_244);
and U701 (N_701,In_188,In_0);
or U702 (N_702,In_66,In_377);
or U703 (N_703,In_774,In_28);
and U704 (N_704,In_105,In_777);
and U705 (N_705,In_29,In_499);
and U706 (N_706,In_37,In_908);
nand U707 (N_707,In_757,In_986);
nor U708 (N_708,In_973,In_142);
and U709 (N_709,In_475,In_293);
or U710 (N_710,In_644,In_737);
and U711 (N_711,In_145,In_159);
xor U712 (N_712,In_215,In_646);
or U713 (N_713,In_11,In_388);
and U714 (N_714,In_756,In_868);
and U715 (N_715,In_682,In_137);
xor U716 (N_716,In_706,In_79);
or U717 (N_717,In_668,In_878);
and U718 (N_718,In_188,In_9);
xor U719 (N_719,In_265,In_863);
nor U720 (N_720,In_612,In_85);
and U721 (N_721,In_289,In_537);
and U722 (N_722,In_969,In_938);
nand U723 (N_723,In_902,In_911);
nor U724 (N_724,In_304,In_607);
and U725 (N_725,In_342,In_840);
nand U726 (N_726,In_193,In_806);
and U727 (N_727,In_557,In_553);
or U728 (N_728,In_589,In_901);
nor U729 (N_729,In_600,In_279);
nor U730 (N_730,In_211,In_680);
and U731 (N_731,In_109,In_937);
or U732 (N_732,In_513,In_625);
or U733 (N_733,In_817,In_440);
nand U734 (N_734,In_159,In_200);
nor U735 (N_735,In_514,In_533);
and U736 (N_736,In_874,In_60);
or U737 (N_737,In_460,In_688);
nand U738 (N_738,In_381,In_932);
or U739 (N_739,In_639,In_369);
nor U740 (N_740,In_559,In_709);
nand U741 (N_741,In_594,In_806);
or U742 (N_742,In_758,In_495);
nor U743 (N_743,In_339,In_327);
nand U744 (N_744,In_950,In_139);
nor U745 (N_745,In_697,In_401);
or U746 (N_746,In_309,In_743);
nand U747 (N_747,In_236,In_864);
nand U748 (N_748,In_82,In_866);
or U749 (N_749,In_68,In_960);
xnor U750 (N_750,In_633,In_258);
nor U751 (N_751,In_716,In_777);
or U752 (N_752,In_482,In_838);
and U753 (N_753,In_45,In_98);
nor U754 (N_754,In_806,In_274);
xnor U755 (N_755,In_243,In_616);
and U756 (N_756,In_703,In_344);
nand U757 (N_757,In_83,In_339);
nand U758 (N_758,In_233,In_198);
or U759 (N_759,In_534,In_964);
nor U760 (N_760,In_590,In_347);
and U761 (N_761,In_256,In_538);
or U762 (N_762,In_172,In_919);
nor U763 (N_763,In_517,In_355);
nand U764 (N_764,In_104,In_808);
nand U765 (N_765,In_36,In_872);
or U766 (N_766,In_736,In_232);
and U767 (N_767,In_586,In_29);
and U768 (N_768,In_877,In_343);
and U769 (N_769,In_947,In_99);
nor U770 (N_770,In_346,In_918);
or U771 (N_771,In_401,In_886);
nand U772 (N_772,In_230,In_713);
nand U773 (N_773,In_214,In_41);
and U774 (N_774,In_299,In_639);
and U775 (N_775,In_318,In_899);
and U776 (N_776,In_568,In_862);
and U777 (N_777,In_731,In_396);
or U778 (N_778,In_296,In_667);
or U779 (N_779,In_113,In_411);
nor U780 (N_780,In_50,In_596);
nor U781 (N_781,In_989,In_897);
and U782 (N_782,In_305,In_797);
nor U783 (N_783,In_930,In_47);
nand U784 (N_784,In_700,In_510);
nor U785 (N_785,In_801,In_446);
or U786 (N_786,In_309,In_660);
nor U787 (N_787,In_232,In_524);
or U788 (N_788,In_112,In_934);
nand U789 (N_789,In_33,In_983);
nor U790 (N_790,In_623,In_222);
nand U791 (N_791,In_860,In_626);
nor U792 (N_792,In_160,In_967);
nor U793 (N_793,In_893,In_240);
and U794 (N_794,In_701,In_209);
nor U795 (N_795,In_305,In_722);
nor U796 (N_796,In_483,In_693);
nand U797 (N_797,In_392,In_16);
nor U798 (N_798,In_707,In_997);
nor U799 (N_799,In_430,In_153);
or U800 (N_800,In_112,In_711);
xnor U801 (N_801,In_336,In_488);
nor U802 (N_802,In_935,In_50);
and U803 (N_803,In_159,In_169);
nor U804 (N_804,In_720,In_161);
nand U805 (N_805,In_278,In_259);
nor U806 (N_806,In_702,In_203);
nand U807 (N_807,In_112,In_190);
nand U808 (N_808,In_300,In_486);
or U809 (N_809,In_111,In_334);
nand U810 (N_810,In_300,In_170);
and U811 (N_811,In_986,In_326);
nor U812 (N_812,In_976,In_89);
or U813 (N_813,In_461,In_780);
nor U814 (N_814,In_218,In_587);
or U815 (N_815,In_861,In_130);
nor U816 (N_816,In_207,In_860);
nor U817 (N_817,In_99,In_379);
and U818 (N_818,In_744,In_673);
and U819 (N_819,In_467,In_11);
and U820 (N_820,In_333,In_633);
or U821 (N_821,In_384,In_682);
and U822 (N_822,In_656,In_938);
or U823 (N_823,In_480,In_136);
nand U824 (N_824,In_247,In_486);
and U825 (N_825,In_994,In_90);
nor U826 (N_826,In_805,In_593);
nor U827 (N_827,In_316,In_520);
and U828 (N_828,In_880,In_185);
and U829 (N_829,In_993,In_952);
nand U830 (N_830,In_235,In_306);
nand U831 (N_831,In_858,In_128);
nand U832 (N_832,In_823,In_933);
nand U833 (N_833,In_845,In_778);
xor U834 (N_834,In_746,In_431);
and U835 (N_835,In_590,In_237);
and U836 (N_836,In_302,In_828);
or U837 (N_837,In_650,In_525);
nand U838 (N_838,In_164,In_417);
nor U839 (N_839,In_731,In_362);
nor U840 (N_840,In_814,In_528);
nand U841 (N_841,In_625,In_294);
nand U842 (N_842,In_838,In_174);
and U843 (N_843,In_846,In_444);
or U844 (N_844,In_585,In_86);
nand U845 (N_845,In_97,In_568);
and U846 (N_846,In_167,In_56);
nand U847 (N_847,In_947,In_704);
nor U848 (N_848,In_502,In_847);
nand U849 (N_849,In_779,In_633);
or U850 (N_850,In_192,In_368);
nor U851 (N_851,In_342,In_853);
and U852 (N_852,In_57,In_712);
nand U853 (N_853,In_318,In_900);
nand U854 (N_854,In_878,In_585);
nand U855 (N_855,In_95,In_629);
nand U856 (N_856,In_813,In_344);
or U857 (N_857,In_469,In_64);
or U858 (N_858,In_506,In_525);
and U859 (N_859,In_908,In_380);
nand U860 (N_860,In_557,In_824);
nand U861 (N_861,In_348,In_748);
nor U862 (N_862,In_915,In_147);
nand U863 (N_863,In_310,In_125);
nand U864 (N_864,In_164,In_661);
or U865 (N_865,In_357,In_942);
or U866 (N_866,In_188,In_329);
nand U867 (N_867,In_599,In_156);
and U868 (N_868,In_531,In_211);
or U869 (N_869,In_603,In_25);
and U870 (N_870,In_938,In_966);
nand U871 (N_871,In_546,In_65);
and U872 (N_872,In_72,In_258);
nand U873 (N_873,In_416,In_603);
or U874 (N_874,In_797,In_367);
or U875 (N_875,In_664,In_55);
or U876 (N_876,In_231,In_48);
nand U877 (N_877,In_809,In_467);
or U878 (N_878,In_146,In_289);
or U879 (N_879,In_609,In_164);
nor U880 (N_880,In_767,In_861);
nand U881 (N_881,In_223,In_206);
and U882 (N_882,In_628,In_858);
nor U883 (N_883,In_886,In_234);
and U884 (N_884,In_625,In_615);
nand U885 (N_885,In_927,In_419);
nor U886 (N_886,In_895,In_824);
nand U887 (N_887,In_680,In_6);
nand U888 (N_888,In_606,In_187);
or U889 (N_889,In_252,In_255);
nor U890 (N_890,In_407,In_782);
nor U891 (N_891,In_74,In_335);
and U892 (N_892,In_360,In_758);
and U893 (N_893,In_639,In_134);
xnor U894 (N_894,In_44,In_957);
xnor U895 (N_895,In_777,In_883);
or U896 (N_896,In_671,In_274);
nor U897 (N_897,In_896,In_237);
nand U898 (N_898,In_832,In_628);
xor U899 (N_899,In_534,In_771);
or U900 (N_900,In_558,In_122);
or U901 (N_901,In_376,In_568);
nand U902 (N_902,In_805,In_777);
or U903 (N_903,In_20,In_574);
nand U904 (N_904,In_265,In_384);
or U905 (N_905,In_984,In_489);
nor U906 (N_906,In_205,In_811);
and U907 (N_907,In_196,In_229);
nor U908 (N_908,In_519,In_171);
and U909 (N_909,In_878,In_867);
and U910 (N_910,In_174,In_29);
nor U911 (N_911,In_827,In_350);
nor U912 (N_912,In_953,In_36);
nor U913 (N_913,In_962,In_312);
nor U914 (N_914,In_401,In_313);
and U915 (N_915,In_187,In_651);
and U916 (N_916,In_408,In_261);
nand U917 (N_917,In_278,In_225);
or U918 (N_918,In_52,In_100);
and U919 (N_919,In_214,In_91);
nand U920 (N_920,In_691,In_918);
or U921 (N_921,In_459,In_813);
or U922 (N_922,In_818,In_515);
nand U923 (N_923,In_615,In_850);
nand U924 (N_924,In_472,In_777);
or U925 (N_925,In_879,In_225);
or U926 (N_926,In_155,In_786);
nand U927 (N_927,In_90,In_523);
nor U928 (N_928,In_861,In_319);
nand U929 (N_929,In_639,In_356);
nor U930 (N_930,In_446,In_862);
xnor U931 (N_931,In_967,In_781);
nor U932 (N_932,In_394,In_813);
nand U933 (N_933,In_873,In_392);
and U934 (N_934,In_922,In_38);
or U935 (N_935,In_946,In_77);
or U936 (N_936,In_934,In_983);
nand U937 (N_937,In_877,In_747);
or U938 (N_938,In_144,In_795);
and U939 (N_939,In_635,In_143);
nand U940 (N_940,In_272,In_506);
nor U941 (N_941,In_199,In_994);
nand U942 (N_942,In_282,In_756);
and U943 (N_943,In_934,In_53);
or U944 (N_944,In_103,In_339);
and U945 (N_945,In_501,In_728);
and U946 (N_946,In_22,In_600);
or U947 (N_947,In_850,In_706);
or U948 (N_948,In_407,In_223);
nor U949 (N_949,In_649,In_33);
nand U950 (N_950,In_895,In_381);
nor U951 (N_951,In_480,In_38);
xnor U952 (N_952,In_680,In_647);
and U953 (N_953,In_922,In_251);
nor U954 (N_954,In_804,In_439);
or U955 (N_955,In_847,In_628);
nand U956 (N_956,In_239,In_809);
and U957 (N_957,In_608,In_454);
and U958 (N_958,In_676,In_314);
or U959 (N_959,In_485,In_856);
or U960 (N_960,In_384,In_527);
and U961 (N_961,In_748,In_383);
nor U962 (N_962,In_355,In_210);
or U963 (N_963,In_646,In_8);
nor U964 (N_964,In_851,In_586);
nor U965 (N_965,In_239,In_934);
nand U966 (N_966,In_490,In_62);
nor U967 (N_967,In_718,In_620);
nand U968 (N_968,In_927,In_286);
nand U969 (N_969,In_597,In_951);
nand U970 (N_970,In_175,In_183);
nor U971 (N_971,In_65,In_539);
or U972 (N_972,In_670,In_89);
nor U973 (N_973,In_525,In_147);
nor U974 (N_974,In_75,In_324);
nor U975 (N_975,In_532,In_700);
and U976 (N_976,In_113,In_268);
and U977 (N_977,In_722,In_598);
and U978 (N_978,In_957,In_617);
nor U979 (N_979,In_464,In_904);
and U980 (N_980,In_875,In_539);
and U981 (N_981,In_276,In_67);
nand U982 (N_982,In_343,In_408);
or U983 (N_983,In_2,In_956);
nor U984 (N_984,In_681,In_827);
nor U985 (N_985,In_142,In_983);
nand U986 (N_986,In_743,In_432);
and U987 (N_987,In_583,In_651);
or U988 (N_988,In_129,In_230);
nor U989 (N_989,In_703,In_951);
nand U990 (N_990,In_323,In_378);
nand U991 (N_991,In_44,In_407);
and U992 (N_992,In_805,In_413);
nand U993 (N_993,In_562,In_109);
nor U994 (N_994,In_900,In_357);
nand U995 (N_995,In_682,In_290);
or U996 (N_996,In_20,In_136);
and U997 (N_997,In_316,In_606);
or U998 (N_998,In_738,In_333);
nor U999 (N_999,In_713,In_500);
and U1000 (N_1000,In_461,In_674);
nor U1001 (N_1001,In_442,In_933);
and U1002 (N_1002,In_492,In_747);
and U1003 (N_1003,In_100,In_575);
and U1004 (N_1004,In_643,In_949);
nor U1005 (N_1005,In_957,In_142);
nand U1006 (N_1006,In_962,In_110);
nand U1007 (N_1007,In_516,In_195);
and U1008 (N_1008,In_468,In_155);
nand U1009 (N_1009,In_563,In_198);
nor U1010 (N_1010,In_177,In_183);
or U1011 (N_1011,In_50,In_23);
nor U1012 (N_1012,In_119,In_614);
and U1013 (N_1013,In_525,In_769);
and U1014 (N_1014,In_321,In_995);
nand U1015 (N_1015,In_699,In_15);
and U1016 (N_1016,In_160,In_384);
xor U1017 (N_1017,In_932,In_784);
nor U1018 (N_1018,In_533,In_741);
nor U1019 (N_1019,In_956,In_280);
xnor U1020 (N_1020,In_385,In_599);
nor U1021 (N_1021,In_882,In_791);
or U1022 (N_1022,In_122,In_196);
and U1023 (N_1023,In_825,In_678);
nor U1024 (N_1024,In_305,In_842);
nand U1025 (N_1025,In_417,In_456);
nand U1026 (N_1026,In_313,In_732);
and U1027 (N_1027,In_913,In_136);
nand U1028 (N_1028,In_162,In_658);
nand U1029 (N_1029,In_324,In_341);
nor U1030 (N_1030,In_16,In_666);
and U1031 (N_1031,In_318,In_716);
or U1032 (N_1032,In_871,In_549);
nor U1033 (N_1033,In_87,In_100);
and U1034 (N_1034,In_297,In_298);
and U1035 (N_1035,In_299,In_761);
and U1036 (N_1036,In_864,In_606);
and U1037 (N_1037,In_802,In_147);
or U1038 (N_1038,In_352,In_910);
nor U1039 (N_1039,In_374,In_375);
nor U1040 (N_1040,In_137,In_706);
or U1041 (N_1041,In_933,In_199);
nand U1042 (N_1042,In_725,In_968);
or U1043 (N_1043,In_942,In_963);
nand U1044 (N_1044,In_790,In_343);
and U1045 (N_1045,In_443,In_871);
or U1046 (N_1046,In_118,In_173);
or U1047 (N_1047,In_842,In_283);
or U1048 (N_1048,In_830,In_937);
nand U1049 (N_1049,In_376,In_426);
or U1050 (N_1050,In_531,In_308);
nand U1051 (N_1051,In_893,In_317);
nand U1052 (N_1052,In_935,In_397);
or U1053 (N_1053,In_480,In_525);
nand U1054 (N_1054,In_789,In_22);
nor U1055 (N_1055,In_237,In_393);
nand U1056 (N_1056,In_252,In_389);
and U1057 (N_1057,In_702,In_374);
or U1058 (N_1058,In_525,In_761);
or U1059 (N_1059,In_598,In_502);
and U1060 (N_1060,In_853,In_320);
nor U1061 (N_1061,In_727,In_648);
xnor U1062 (N_1062,In_869,In_836);
nor U1063 (N_1063,In_778,In_841);
or U1064 (N_1064,In_255,In_109);
nor U1065 (N_1065,In_219,In_755);
nand U1066 (N_1066,In_915,In_584);
nor U1067 (N_1067,In_432,In_599);
and U1068 (N_1068,In_493,In_636);
nand U1069 (N_1069,In_916,In_956);
nand U1070 (N_1070,In_207,In_836);
or U1071 (N_1071,In_956,In_315);
nand U1072 (N_1072,In_934,In_424);
and U1073 (N_1073,In_336,In_344);
nand U1074 (N_1074,In_929,In_279);
nor U1075 (N_1075,In_286,In_398);
nand U1076 (N_1076,In_347,In_23);
nand U1077 (N_1077,In_913,In_455);
nor U1078 (N_1078,In_952,In_527);
nand U1079 (N_1079,In_553,In_627);
and U1080 (N_1080,In_332,In_95);
or U1081 (N_1081,In_441,In_537);
or U1082 (N_1082,In_681,In_968);
and U1083 (N_1083,In_809,In_341);
nor U1084 (N_1084,In_65,In_578);
nand U1085 (N_1085,In_724,In_239);
nor U1086 (N_1086,In_775,In_464);
nand U1087 (N_1087,In_937,In_676);
nor U1088 (N_1088,In_399,In_833);
or U1089 (N_1089,In_493,In_933);
nand U1090 (N_1090,In_996,In_314);
or U1091 (N_1091,In_245,In_350);
nand U1092 (N_1092,In_143,In_908);
or U1093 (N_1093,In_897,In_129);
nand U1094 (N_1094,In_415,In_91);
nand U1095 (N_1095,In_628,In_271);
and U1096 (N_1096,In_315,In_589);
nand U1097 (N_1097,In_240,In_503);
or U1098 (N_1098,In_83,In_209);
nand U1099 (N_1099,In_390,In_487);
nor U1100 (N_1100,In_489,In_667);
nand U1101 (N_1101,In_257,In_213);
nor U1102 (N_1102,In_819,In_69);
and U1103 (N_1103,In_758,In_673);
nor U1104 (N_1104,In_738,In_446);
nor U1105 (N_1105,In_899,In_498);
or U1106 (N_1106,In_972,In_84);
nand U1107 (N_1107,In_168,In_110);
and U1108 (N_1108,In_847,In_25);
xor U1109 (N_1109,In_980,In_561);
nor U1110 (N_1110,In_323,In_286);
nor U1111 (N_1111,In_562,In_454);
nand U1112 (N_1112,In_582,In_358);
nand U1113 (N_1113,In_453,In_370);
nor U1114 (N_1114,In_170,In_426);
or U1115 (N_1115,In_33,In_685);
or U1116 (N_1116,In_357,In_925);
nand U1117 (N_1117,In_728,In_665);
nor U1118 (N_1118,In_684,In_145);
or U1119 (N_1119,In_886,In_78);
and U1120 (N_1120,In_969,In_608);
nor U1121 (N_1121,In_912,In_533);
or U1122 (N_1122,In_271,In_256);
nand U1123 (N_1123,In_72,In_120);
or U1124 (N_1124,In_180,In_732);
nor U1125 (N_1125,In_511,In_106);
or U1126 (N_1126,In_684,In_902);
nor U1127 (N_1127,In_379,In_133);
and U1128 (N_1128,In_862,In_606);
nand U1129 (N_1129,In_174,In_457);
or U1130 (N_1130,In_443,In_726);
or U1131 (N_1131,In_210,In_299);
nand U1132 (N_1132,In_815,In_206);
nand U1133 (N_1133,In_497,In_424);
nor U1134 (N_1134,In_216,In_766);
and U1135 (N_1135,In_350,In_653);
or U1136 (N_1136,In_257,In_987);
nor U1137 (N_1137,In_495,In_709);
nor U1138 (N_1138,In_753,In_732);
nand U1139 (N_1139,In_376,In_519);
nor U1140 (N_1140,In_810,In_561);
nor U1141 (N_1141,In_274,In_954);
or U1142 (N_1142,In_875,In_225);
nand U1143 (N_1143,In_282,In_399);
and U1144 (N_1144,In_574,In_741);
nand U1145 (N_1145,In_557,In_691);
and U1146 (N_1146,In_20,In_5);
or U1147 (N_1147,In_882,In_838);
or U1148 (N_1148,In_734,In_623);
and U1149 (N_1149,In_898,In_970);
nor U1150 (N_1150,In_18,In_33);
or U1151 (N_1151,In_582,In_943);
nand U1152 (N_1152,In_26,In_705);
or U1153 (N_1153,In_946,In_246);
nor U1154 (N_1154,In_823,In_709);
or U1155 (N_1155,In_350,In_540);
or U1156 (N_1156,In_669,In_150);
nor U1157 (N_1157,In_820,In_350);
xnor U1158 (N_1158,In_797,In_32);
nor U1159 (N_1159,In_203,In_943);
and U1160 (N_1160,In_249,In_960);
nand U1161 (N_1161,In_213,In_542);
nand U1162 (N_1162,In_727,In_478);
and U1163 (N_1163,In_744,In_944);
or U1164 (N_1164,In_291,In_876);
and U1165 (N_1165,In_431,In_920);
or U1166 (N_1166,In_910,In_515);
nor U1167 (N_1167,In_338,In_264);
or U1168 (N_1168,In_873,In_826);
nand U1169 (N_1169,In_465,In_295);
or U1170 (N_1170,In_318,In_538);
nand U1171 (N_1171,In_738,In_361);
or U1172 (N_1172,In_36,In_825);
and U1173 (N_1173,In_176,In_179);
or U1174 (N_1174,In_40,In_782);
or U1175 (N_1175,In_271,In_456);
and U1176 (N_1176,In_519,In_146);
nand U1177 (N_1177,In_342,In_21);
nand U1178 (N_1178,In_622,In_329);
or U1179 (N_1179,In_851,In_486);
or U1180 (N_1180,In_556,In_555);
nor U1181 (N_1181,In_365,In_400);
or U1182 (N_1182,In_835,In_645);
or U1183 (N_1183,In_908,In_722);
nand U1184 (N_1184,In_965,In_903);
xor U1185 (N_1185,In_208,In_522);
or U1186 (N_1186,In_460,In_213);
nor U1187 (N_1187,In_914,In_372);
and U1188 (N_1188,In_718,In_697);
or U1189 (N_1189,In_954,In_738);
nor U1190 (N_1190,In_940,In_943);
nor U1191 (N_1191,In_349,In_635);
and U1192 (N_1192,In_315,In_547);
or U1193 (N_1193,In_54,In_66);
or U1194 (N_1194,In_978,In_176);
or U1195 (N_1195,In_386,In_53);
nor U1196 (N_1196,In_476,In_114);
nor U1197 (N_1197,In_844,In_773);
nor U1198 (N_1198,In_502,In_644);
and U1199 (N_1199,In_499,In_297);
and U1200 (N_1200,In_386,In_573);
or U1201 (N_1201,In_182,In_753);
and U1202 (N_1202,In_14,In_811);
or U1203 (N_1203,In_802,In_524);
and U1204 (N_1204,In_811,In_690);
and U1205 (N_1205,In_103,In_407);
nand U1206 (N_1206,In_573,In_948);
nand U1207 (N_1207,In_887,In_230);
nor U1208 (N_1208,In_248,In_984);
nor U1209 (N_1209,In_207,In_194);
nor U1210 (N_1210,In_936,In_22);
and U1211 (N_1211,In_471,In_743);
or U1212 (N_1212,In_316,In_242);
nand U1213 (N_1213,In_785,In_573);
nor U1214 (N_1214,In_737,In_850);
and U1215 (N_1215,In_419,In_31);
nor U1216 (N_1216,In_454,In_907);
or U1217 (N_1217,In_959,In_317);
or U1218 (N_1218,In_941,In_381);
nor U1219 (N_1219,In_962,In_455);
nand U1220 (N_1220,In_517,In_399);
nand U1221 (N_1221,In_266,In_781);
nor U1222 (N_1222,In_453,In_921);
nand U1223 (N_1223,In_533,In_563);
nand U1224 (N_1224,In_34,In_398);
and U1225 (N_1225,In_761,In_35);
or U1226 (N_1226,In_853,In_798);
nor U1227 (N_1227,In_750,In_356);
nor U1228 (N_1228,In_227,In_904);
nand U1229 (N_1229,In_384,In_976);
or U1230 (N_1230,In_965,In_210);
and U1231 (N_1231,In_626,In_435);
nor U1232 (N_1232,In_198,In_69);
nand U1233 (N_1233,In_590,In_377);
and U1234 (N_1234,In_866,In_153);
nor U1235 (N_1235,In_37,In_778);
nand U1236 (N_1236,In_443,In_703);
and U1237 (N_1237,In_272,In_544);
or U1238 (N_1238,In_502,In_552);
or U1239 (N_1239,In_62,In_337);
nand U1240 (N_1240,In_865,In_388);
or U1241 (N_1241,In_951,In_605);
nand U1242 (N_1242,In_292,In_41);
and U1243 (N_1243,In_710,In_71);
and U1244 (N_1244,In_294,In_319);
and U1245 (N_1245,In_529,In_344);
and U1246 (N_1246,In_206,In_915);
xnor U1247 (N_1247,In_76,In_804);
xor U1248 (N_1248,In_40,In_617);
or U1249 (N_1249,In_554,In_590);
and U1250 (N_1250,In_919,In_309);
nor U1251 (N_1251,In_757,In_941);
and U1252 (N_1252,In_82,In_752);
and U1253 (N_1253,In_340,In_425);
nand U1254 (N_1254,In_375,In_600);
nor U1255 (N_1255,In_872,In_9);
nor U1256 (N_1256,In_106,In_169);
nor U1257 (N_1257,In_825,In_44);
nand U1258 (N_1258,In_440,In_933);
and U1259 (N_1259,In_6,In_68);
or U1260 (N_1260,In_478,In_997);
and U1261 (N_1261,In_744,In_770);
and U1262 (N_1262,In_465,In_766);
nand U1263 (N_1263,In_232,In_202);
nand U1264 (N_1264,In_990,In_579);
nor U1265 (N_1265,In_146,In_620);
and U1266 (N_1266,In_779,In_79);
nor U1267 (N_1267,In_564,In_323);
xor U1268 (N_1268,In_416,In_586);
and U1269 (N_1269,In_889,In_375);
and U1270 (N_1270,In_907,In_60);
nand U1271 (N_1271,In_424,In_874);
and U1272 (N_1272,In_104,In_151);
and U1273 (N_1273,In_545,In_895);
or U1274 (N_1274,In_156,In_641);
nand U1275 (N_1275,In_970,In_749);
and U1276 (N_1276,In_355,In_796);
or U1277 (N_1277,In_678,In_996);
and U1278 (N_1278,In_321,In_882);
and U1279 (N_1279,In_32,In_161);
nor U1280 (N_1280,In_616,In_249);
and U1281 (N_1281,In_748,In_690);
or U1282 (N_1282,In_458,In_901);
nor U1283 (N_1283,In_737,In_379);
nand U1284 (N_1284,In_34,In_862);
and U1285 (N_1285,In_14,In_350);
or U1286 (N_1286,In_464,In_478);
nand U1287 (N_1287,In_329,In_559);
and U1288 (N_1288,In_114,In_447);
nand U1289 (N_1289,In_211,In_201);
nor U1290 (N_1290,In_453,In_685);
xnor U1291 (N_1291,In_889,In_825);
nand U1292 (N_1292,In_331,In_797);
nand U1293 (N_1293,In_488,In_290);
and U1294 (N_1294,In_750,In_925);
and U1295 (N_1295,In_885,In_504);
and U1296 (N_1296,In_107,In_342);
nor U1297 (N_1297,In_358,In_324);
or U1298 (N_1298,In_563,In_790);
nand U1299 (N_1299,In_414,In_792);
nor U1300 (N_1300,In_183,In_669);
nor U1301 (N_1301,In_558,In_818);
nand U1302 (N_1302,In_968,In_385);
nand U1303 (N_1303,In_866,In_268);
nor U1304 (N_1304,In_530,In_750);
or U1305 (N_1305,In_385,In_138);
and U1306 (N_1306,In_753,In_144);
nand U1307 (N_1307,In_290,In_104);
or U1308 (N_1308,In_639,In_324);
nand U1309 (N_1309,In_272,In_15);
nor U1310 (N_1310,In_88,In_435);
or U1311 (N_1311,In_712,In_34);
nand U1312 (N_1312,In_415,In_421);
and U1313 (N_1313,In_479,In_144);
nor U1314 (N_1314,In_303,In_632);
and U1315 (N_1315,In_94,In_893);
nand U1316 (N_1316,In_999,In_576);
or U1317 (N_1317,In_409,In_207);
nand U1318 (N_1318,In_707,In_364);
nand U1319 (N_1319,In_490,In_306);
nand U1320 (N_1320,In_124,In_710);
xor U1321 (N_1321,In_382,In_539);
nand U1322 (N_1322,In_44,In_395);
nand U1323 (N_1323,In_409,In_874);
nand U1324 (N_1324,In_32,In_584);
nor U1325 (N_1325,In_818,In_666);
and U1326 (N_1326,In_10,In_236);
and U1327 (N_1327,In_58,In_833);
xor U1328 (N_1328,In_343,In_229);
or U1329 (N_1329,In_636,In_575);
or U1330 (N_1330,In_550,In_791);
and U1331 (N_1331,In_789,In_816);
and U1332 (N_1332,In_82,In_68);
and U1333 (N_1333,In_344,In_965);
nand U1334 (N_1334,In_421,In_423);
and U1335 (N_1335,In_409,In_910);
and U1336 (N_1336,In_244,In_538);
or U1337 (N_1337,In_446,In_325);
or U1338 (N_1338,In_689,In_961);
or U1339 (N_1339,In_56,In_250);
nor U1340 (N_1340,In_618,In_465);
nand U1341 (N_1341,In_506,In_211);
nand U1342 (N_1342,In_506,In_131);
nand U1343 (N_1343,In_301,In_333);
or U1344 (N_1344,In_894,In_410);
or U1345 (N_1345,In_967,In_209);
nor U1346 (N_1346,In_768,In_981);
and U1347 (N_1347,In_885,In_503);
or U1348 (N_1348,In_674,In_108);
nand U1349 (N_1349,In_658,In_799);
nand U1350 (N_1350,In_665,In_1);
nand U1351 (N_1351,In_78,In_368);
nor U1352 (N_1352,In_710,In_893);
and U1353 (N_1353,In_979,In_540);
or U1354 (N_1354,In_895,In_860);
and U1355 (N_1355,In_145,In_768);
and U1356 (N_1356,In_183,In_333);
and U1357 (N_1357,In_973,In_732);
or U1358 (N_1358,In_426,In_637);
xnor U1359 (N_1359,In_106,In_905);
or U1360 (N_1360,In_325,In_609);
nor U1361 (N_1361,In_216,In_539);
nor U1362 (N_1362,In_974,In_347);
nand U1363 (N_1363,In_254,In_169);
nand U1364 (N_1364,In_931,In_118);
nor U1365 (N_1365,In_951,In_562);
nand U1366 (N_1366,In_948,In_55);
and U1367 (N_1367,In_242,In_724);
nor U1368 (N_1368,In_233,In_993);
nand U1369 (N_1369,In_684,In_634);
nor U1370 (N_1370,In_213,In_259);
nor U1371 (N_1371,In_18,In_643);
or U1372 (N_1372,In_412,In_542);
or U1373 (N_1373,In_363,In_96);
and U1374 (N_1374,In_506,In_65);
nor U1375 (N_1375,In_172,In_385);
xnor U1376 (N_1376,In_179,In_978);
and U1377 (N_1377,In_953,In_2);
and U1378 (N_1378,In_251,In_62);
nand U1379 (N_1379,In_449,In_368);
and U1380 (N_1380,In_329,In_935);
or U1381 (N_1381,In_977,In_568);
and U1382 (N_1382,In_404,In_549);
or U1383 (N_1383,In_693,In_395);
nor U1384 (N_1384,In_700,In_530);
nand U1385 (N_1385,In_235,In_381);
nor U1386 (N_1386,In_475,In_425);
or U1387 (N_1387,In_336,In_664);
and U1388 (N_1388,In_546,In_614);
and U1389 (N_1389,In_593,In_935);
nor U1390 (N_1390,In_91,In_521);
and U1391 (N_1391,In_812,In_356);
or U1392 (N_1392,In_240,In_564);
or U1393 (N_1393,In_380,In_9);
nand U1394 (N_1394,In_305,In_891);
and U1395 (N_1395,In_517,In_224);
and U1396 (N_1396,In_958,In_347);
and U1397 (N_1397,In_772,In_858);
and U1398 (N_1398,In_878,In_959);
nor U1399 (N_1399,In_885,In_441);
nand U1400 (N_1400,In_798,In_820);
nor U1401 (N_1401,In_989,In_236);
nor U1402 (N_1402,In_528,In_115);
and U1403 (N_1403,In_363,In_607);
nand U1404 (N_1404,In_31,In_535);
and U1405 (N_1405,In_356,In_504);
and U1406 (N_1406,In_834,In_161);
or U1407 (N_1407,In_256,In_341);
nand U1408 (N_1408,In_749,In_727);
and U1409 (N_1409,In_691,In_309);
and U1410 (N_1410,In_274,In_79);
and U1411 (N_1411,In_481,In_262);
nand U1412 (N_1412,In_738,In_694);
or U1413 (N_1413,In_754,In_745);
nor U1414 (N_1414,In_41,In_421);
nor U1415 (N_1415,In_347,In_460);
nor U1416 (N_1416,In_528,In_751);
or U1417 (N_1417,In_359,In_527);
nor U1418 (N_1418,In_47,In_771);
and U1419 (N_1419,In_366,In_556);
nor U1420 (N_1420,In_507,In_528);
nand U1421 (N_1421,In_833,In_907);
nand U1422 (N_1422,In_213,In_679);
and U1423 (N_1423,In_611,In_565);
or U1424 (N_1424,In_906,In_548);
and U1425 (N_1425,In_660,In_219);
nor U1426 (N_1426,In_231,In_325);
or U1427 (N_1427,In_87,In_176);
nor U1428 (N_1428,In_250,In_420);
nor U1429 (N_1429,In_909,In_677);
or U1430 (N_1430,In_789,In_976);
or U1431 (N_1431,In_529,In_7);
nand U1432 (N_1432,In_330,In_805);
and U1433 (N_1433,In_646,In_513);
or U1434 (N_1434,In_792,In_360);
nor U1435 (N_1435,In_834,In_386);
nor U1436 (N_1436,In_606,In_310);
nand U1437 (N_1437,In_545,In_657);
nand U1438 (N_1438,In_623,In_982);
or U1439 (N_1439,In_186,In_304);
nand U1440 (N_1440,In_426,In_420);
nor U1441 (N_1441,In_709,In_426);
nor U1442 (N_1442,In_67,In_807);
nor U1443 (N_1443,In_568,In_323);
or U1444 (N_1444,In_803,In_73);
nand U1445 (N_1445,In_558,In_246);
nor U1446 (N_1446,In_902,In_593);
or U1447 (N_1447,In_54,In_815);
or U1448 (N_1448,In_66,In_323);
and U1449 (N_1449,In_568,In_342);
nand U1450 (N_1450,In_663,In_564);
and U1451 (N_1451,In_110,In_573);
nor U1452 (N_1452,In_839,In_468);
nand U1453 (N_1453,In_75,In_803);
nand U1454 (N_1454,In_450,In_120);
and U1455 (N_1455,In_264,In_30);
nand U1456 (N_1456,In_547,In_630);
and U1457 (N_1457,In_432,In_246);
and U1458 (N_1458,In_888,In_191);
nand U1459 (N_1459,In_33,In_671);
or U1460 (N_1460,In_614,In_101);
and U1461 (N_1461,In_789,In_782);
nor U1462 (N_1462,In_882,In_281);
nor U1463 (N_1463,In_387,In_509);
nor U1464 (N_1464,In_642,In_175);
and U1465 (N_1465,In_618,In_384);
nand U1466 (N_1466,In_395,In_267);
xnor U1467 (N_1467,In_390,In_374);
nor U1468 (N_1468,In_274,In_516);
nand U1469 (N_1469,In_341,In_826);
or U1470 (N_1470,In_226,In_362);
nand U1471 (N_1471,In_505,In_167);
and U1472 (N_1472,In_155,In_156);
and U1473 (N_1473,In_255,In_322);
or U1474 (N_1474,In_703,In_972);
nand U1475 (N_1475,In_208,In_504);
or U1476 (N_1476,In_309,In_341);
nor U1477 (N_1477,In_490,In_891);
nor U1478 (N_1478,In_667,In_647);
nor U1479 (N_1479,In_993,In_241);
or U1480 (N_1480,In_608,In_990);
nor U1481 (N_1481,In_45,In_706);
and U1482 (N_1482,In_446,In_542);
nand U1483 (N_1483,In_410,In_879);
and U1484 (N_1484,In_860,In_732);
nor U1485 (N_1485,In_582,In_218);
xor U1486 (N_1486,In_381,In_354);
nor U1487 (N_1487,In_600,In_353);
or U1488 (N_1488,In_893,In_156);
and U1489 (N_1489,In_114,In_389);
or U1490 (N_1490,In_299,In_759);
and U1491 (N_1491,In_405,In_836);
or U1492 (N_1492,In_708,In_232);
nor U1493 (N_1493,In_271,In_896);
nand U1494 (N_1494,In_964,In_981);
or U1495 (N_1495,In_549,In_232);
and U1496 (N_1496,In_327,In_177);
nor U1497 (N_1497,In_747,In_649);
nor U1498 (N_1498,In_695,In_717);
or U1499 (N_1499,In_594,In_527);
nor U1500 (N_1500,In_938,In_179);
nor U1501 (N_1501,In_232,In_582);
and U1502 (N_1502,In_938,In_300);
or U1503 (N_1503,In_655,In_329);
or U1504 (N_1504,In_956,In_782);
nand U1505 (N_1505,In_783,In_944);
nor U1506 (N_1506,In_796,In_950);
or U1507 (N_1507,In_659,In_18);
nand U1508 (N_1508,In_585,In_13);
nand U1509 (N_1509,In_748,In_651);
or U1510 (N_1510,In_642,In_708);
nor U1511 (N_1511,In_766,In_913);
or U1512 (N_1512,In_479,In_877);
nand U1513 (N_1513,In_484,In_717);
or U1514 (N_1514,In_1,In_699);
nor U1515 (N_1515,In_89,In_746);
or U1516 (N_1516,In_326,In_579);
nand U1517 (N_1517,In_254,In_74);
or U1518 (N_1518,In_40,In_916);
nand U1519 (N_1519,In_210,In_60);
nor U1520 (N_1520,In_162,In_846);
or U1521 (N_1521,In_537,In_458);
xnor U1522 (N_1522,In_371,In_570);
or U1523 (N_1523,In_525,In_232);
and U1524 (N_1524,In_206,In_712);
nor U1525 (N_1525,In_718,In_705);
and U1526 (N_1526,In_38,In_754);
nand U1527 (N_1527,In_710,In_662);
nand U1528 (N_1528,In_284,In_440);
nand U1529 (N_1529,In_851,In_583);
and U1530 (N_1530,In_752,In_518);
nand U1531 (N_1531,In_71,In_136);
nand U1532 (N_1532,In_754,In_632);
or U1533 (N_1533,In_99,In_677);
nand U1534 (N_1534,In_585,In_441);
and U1535 (N_1535,In_315,In_808);
or U1536 (N_1536,In_733,In_818);
nand U1537 (N_1537,In_3,In_159);
nor U1538 (N_1538,In_358,In_462);
and U1539 (N_1539,In_872,In_5);
nand U1540 (N_1540,In_75,In_226);
xor U1541 (N_1541,In_667,In_525);
or U1542 (N_1542,In_422,In_624);
or U1543 (N_1543,In_474,In_867);
and U1544 (N_1544,In_354,In_765);
xor U1545 (N_1545,In_58,In_160);
nor U1546 (N_1546,In_725,In_262);
or U1547 (N_1547,In_400,In_185);
nand U1548 (N_1548,In_94,In_332);
or U1549 (N_1549,In_593,In_963);
nand U1550 (N_1550,In_437,In_676);
nand U1551 (N_1551,In_290,In_579);
and U1552 (N_1552,In_63,In_44);
and U1553 (N_1553,In_390,In_235);
or U1554 (N_1554,In_499,In_787);
nand U1555 (N_1555,In_454,In_354);
and U1556 (N_1556,In_733,In_72);
and U1557 (N_1557,In_692,In_16);
or U1558 (N_1558,In_192,In_718);
or U1559 (N_1559,In_799,In_796);
nor U1560 (N_1560,In_669,In_630);
and U1561 (N_1561,In_412,In_226);
and U1562 (N_1562,In_376,In_456);
and U1563 (N_1563,In_54,In_388);
or U1564 (N_1564,In_627,In_366);
xor U1565 (N_1565,In_584,In_567);
or U1566 (N_1566,In_543,In_831);
and U1567 (N_1567,In_287,In_678);
nand U1568 (N_1568,In_950,In_15);
nor U1569 (N_1569,In_106,In_524);
nor U1570 (N_1570,In_501,In_708);
nand U1571 (N_1571,In_538,In_105);
or U1572 (N_1572,In_878,In_993);
nor U1573 (N_1573,In_18,In_283);
and U1574 (N_1574,In_958,In_566);
or U1575 (N_1575,In_804,In_458);
nand U1576 (N_1576,In_614,In_847);
nor U1577 (N_1577,In_296,In_210);
or U1578 (N_1578,In_591,In_356);
and U1579 (N_1579,In_554,In_908);
nand U1580 (N_1580,In_240,In_899);
nand U1581 (N_1581,In_230,In_245);
nand U1582 (N_1582,In_79,In_107);
nor U1583 (N_1583,In_372,In_646);
or U1584 (N_1584,In_275,In_475);
nor U1585 (N_1585,In_285,In_720);
and U1586 (N_1586,In_611,In_789);
xnor U1587 (N_1587,In_540,In_696);
nand U1588 (N_1588,In_992,In_349);
xnor U1589 (N_1589,In_281,In_30);
nor U1590 (N_1590,In_817,In_596);
or U1591 (N_1591,In_507,In_762);
and U1592 (N_1592,In_981,In_709);
or U1593 (N_1593,In_368,In_489);
and U1594 (N_1594,In_800,In_820);
or U1595 (N_1595,In_386,In_544);
and U1596 (N_1596,In_873,In_165);
xnor U1597 (N_1597,In_318,In_879);
and U1598 (N_1598,In_908,In_177);
and U1599 (N_1599,In_650,In_500);
or U1600 (N_1600,In_458,In_266);
and U1601 (N_1601,In_729,In_228);
nor U1602 (N_1602,In_56,In_681);
xnor U1603 (N_1603,In_583,In_370);
or U1604 (N_1604,In_805,In_848);
nor U1605 (N_1605,In_198,In_15);
or U1606 (N_1606,In_878,In_916);
or U1607 (N_1607,In_709,In_544);
nand U1608 (N_1608,In_443,In_585);
nand U1609 (N_1609,In_172,In_97);
and U1610 (N_1610,In_883,In_101);
nor U1611 (N_1611,In_317,In_905);
nand U1612 (N_1612,In_34,In_775);
nand U1613 (N_1613,In_700,In_845);
xor U1614 (N_1614,In_321,In_967);
and U1615 (N_1615,In_441,In_8);
nand U1616 (N_1616,In_79,In_191);
nand U1617 (N_1617,In_600,In_651);
nand U1618 (N_1618,In_9,In_455);
nand U1619 (N_1619,In_635,In_749);
nand U1620 (N_1620,In_832,In_208);
nand U1621 (N_1621,In_718,In_446);
nor U1622 (N_1622,In_616,In_511);
nor U1623 (N_1623,In_140,In_362);
nor U1624 (N_1624,In_603,In_929);
nand U1625 (N_1625,In_119,In_40);
nor U1626 (N_1626,In_558,In_699);
or U1627 (N_1627,In_161,In_476);
nand U1628 (N_1628,In_713,In_927);
or U1629 (N_1629,In_409,In_978);
and U1630 (N_1630,In_312,In_564);
nor U1631 (N_1631,In_956,In_268);
nand U1632 (N_1632,In_498,In_483);
nor U1633 (N_1633,In_639,In_883);
nand U1634 (N_1634,In_948,In_744);
nor U1635 (N_1635,In_135,In_52);
or U1636 (N_1636,In_951,In_137);
nand U1637 (N_1637,In_509,In_548);
and U1638 (N_1638,In_771,In_593);
and U1639 (N_1639,In_725,In_235);
and U1640 (N_1640,In_777,In_208);
nand U1641 (N_1641,In_911,In_177);
nor U1642 (N_1642,In_874,In_13);
nor U1643 (N_1643,In_953,In_786);
or U1644 (N_1644,In_124,In_212);
nor U1645 (N_1645,In_423,In_876);
xor U1646 (N_1646,In_601,In_130);
nor U1647 (N_1647,In_747,In_989);
nand U1648 (N_1648,In_195,In_803);
nor U1649 (N_1649,In_82,In_327);
nor U1650 (N_1650,In_750,In_846);
nor U1651 (N_1651,In_147,In_581);
or U1652 (N_1652,In_558,In_75);
nor U1653 (N_1653,In_43,In_249);
and U1654 (N_1654,In_488,In_906);
nor U1655 (N_1655,In_76,In_416);
and U1656 (N_1656,In_572,In_588);
and U1657 (N_1657,In_523,In_482);
and U1658 (N_1658,In_248,In_689);
nand U1659 (N_1659,In_371,In_419);
nor U1660 (N_1660,In_12,In_780);
or U1661 (N_1661,In_163,In_572);
nand U1662 (N_1662,In_931,In_933);
nor U1663 (N_1663,In_327,In_653);
and U1664 (N_1664,In_710,In_245);
nor U1665 (N_1665,In_361,In_873);
or U1666 (N_1666,In_374,In_147);
or U1667 (N_1667,In_426,In_735);
or U1668 (N_1668,In_814,In_238);
or U1669 (N_1669,In_542,In_11);
nor U1670 (N_1670,In_239,In_8);
nor U1671 (N_1671,In_366,In_436);
nand U1672 (N_1672,In_995,In_615);
and U1673 (N_1673,In_112,In_591);
nand U1674 (N_1674,In_260,In_3);
nor U1675 (N_1675,In_417,In_995);
nor U1676 (N_1676,In_466,In_814);
nand U1677 (N_1677,In_208,In_97);
or U1678 (N_1678,In_405,In_628);
and U1679 (N_1679,In_276,In_605);
and U1680 (N_1680,In_290,In_439);
or U1681 (N_1681,In_982,In_668);
and U1682 (N_1682,In_673,In_41);
nand U1683 (N_1683,In_692,In_240);
nand U1684 (N_1684,In_323,In_546);
nand U1685 (N_1685,In_641,In_622);
and U1686 (N_1686,In_999,In_631);
and U1687 (N_1687,In_77,In_464);
or U1688 (N_1688,In_268,In_226);
nor U1689 (N_1689,In_313,In_854);
or U1690 (N_1690,In_353,In_680);
nor U1691 (N_1691,In_18,In_402);
or U1692 (N_1692,In_809,In_51);
and U1693 (N_1693,In_437,In_497);
or U1694 (N_1694,In_113,In_988);
or U1695 (N_1695,In_478,In_64);
nor U1696 (N_1696,In_498,In_829);
nand U1697 (N_1697,In_866,In_708);
xnor U1698 (N_1698,In_679,In_461);
or U1699 (N_1699,In_147,In_128);
and U1700 (N_1700,In_628,In_965);
nor U1701 (N_1701,In_938,In_477);
nand U1702 (N_1702,In_248,In_782);
or U1703 (N_1703,In_351,In_634);
nor U1704 (N_1704,In_856,In_57);
or U1705 (N_1705,In_878,In_965);
and U1706 (N_1706,In_967,In_266);
nand U1707 (N_1707,In_519,In_123);
nor U1708 (N_1708,In_490,In_123);
nor U1709 (N_1709,In_51,In_812);
nand U1710 (N_1710,In_215,In_429);
or U1711 (N_1711,In_280,In_762);
nor U1712 (N_1712,In_373,In_729);
and U1713 (N_1713,In_517,In_405);
and U1714 (N_1714,In_594,In_783);
or U1715 (N_1715,In_228,In_955);
and U1716 (N_1716,In_495,In_526);
nand U1717 (N_1717,In_178,In_533);
nor U1718 (N_1718,In_397,In_402);
and U1719 (N_1719,In_920,In_728);
nor U1720 (N_1720,In_88,In_464);
or U1721 (N_1721,In_574,In_315);
and U1722 (N_1722,In_606,In_124);
nand U1723 (N_1723,In_760,In_294);
nand U1724 (N_1724,In_878,In_553);
nor U1725 (N_1725,In_766,In_806);
or U1726 (N_1726,In_721,In_35);
or U1727 (N_1727,In_179,In_897);
and U1728 (N_1728,In_629,In_283);
or U1729 (N_1729,In_370,In_103);
and U1730 (N_1730,In_350,In_870);
nor U1731 (N_1731,In_530,In_338);
nand U1732 (N_1732,In_988,In_790);
and U1733 (N_1733,In_289,In_918);
nand U1734 (N_1734,In_532,In_391);
nand U1735 (N_1735,In_571,In_789);
nand U1736 (N_1736,In_575,In_176);
nor U1737 (N_1737,In_292,In_900);
and U1738 (N_1738,In_259,In_990);
nand U1739 (N_1739,In_125,In_945);
or U1740 (N_1740,In_447,In_925);
nor U1741 (N_1741,In_262,In_201);
nand U1742 (N_1742,In_823,In_309);
or U1743 (N_1743,In_475,In_919);
nand U1744 (N_1744,In_947,In_425);
or U1745 (N_1745,In_467,In_763);
nand U1746 (N_1746,In_543,In_142);
nand U1747 (N_1747,In_606,In_638);
xor U1748 (N_1748,In_270,In_99);
or U1749 (N_1749,In_35,In_647);
nor U1750 (N_1750,In_247,In_754);
and U1751 (N_1751,In_92,In_447);
nand U1752 (N_1752,In_218,In_683);
nor U1753 (N_1753,In_277,In_803);
nand U1754 (N_1754,In_607,In_816);
and U1755 (N_1755,In_288,In_541);
or U1756 (N_1756,In_485,In_574);
or U1757 (N_1757,In_429,In_576);
nand U1758 (N_1758,In_314,In_23);
or U1759 (N_1759,In_352,In_528);
and U1760 (N_1760,In_534,In_233);
nor U1761 (N_1761,In_731,In_426);
and U1762 (N_1762,In_189,In_304);
nand U1763 (N_1763,In_7,In_903);
and U1764 (N_1764,In_468,In_417);
xor U1765 (N_1765,In_332,In_852);
nor U1766 (N_1766,In_297,In_274);
nor U1767 (N_1767,In_891,In_485);
or U1768 (N_1768,In_785,In_929);
nor U1769 (N_1769,In_323,In_740);
and U1770 (N_1770,In_57,In_551);
and U1771 (N_1771,In_198,In_591);
nand U1772 (N_1772,In_399,In_246);
nor U1773 (N_1773,In_235,In_595);
nand U1774 (N_1774,In_571,In_421);
nor U1775 (N_1775,In_830,In_870);
nand U1776 (N_1776,In_908,In_804);
and U1777 (N_1777,In_257,In_746);
nor U1778 (N_1778,In_212,In_31);
or U1779 (N_1779,In_895,In_43);
and U1780 (N_1780,In_723,In_482);
nor U1781 (N_1781,In_338,In_323);
nand U1782 (N_1782,In_912,In_601);
nor U1783 (N_1783,In_898,In_653);
nand U1784 (N_1784,In_145,In_69);
nor U1785 (N_1785,In_405,In_302);
and U1786 (N_1786,In_428,In_38);
xnor U1787 (N_1787,In_197,In_478);
and U1788 (N_1788,In_734,In_175);
nor U1789 (N_1789,In_653,In_37);
or U1790 (N_1790,In_500,In_202);
nand U1791 (N_1791,In_663,In_233);
or U1792 (N_1792,In_487,In_143);
nor U1793 (N_1793,In_377,In_490);
xor U1794 (N_1794,In_262,In_303);
nor U1795 (N_1795,In_381,In_683);
nand U1796 (N_1796,In_469,In_577);
nand U1797 (N_1797,In_505,In_834);
nand U1798 (N_1798,In_457,In_340);
nand U1799 (N_1799,In_344,In_483);
or U1800 (N_1800,In_839,In_367);
nor U1801 (N_1801,In_43,In_956);
nand U1802 (N_1802,In_142,In_411);
nor U1803 (N_1803,In_283,In_166);
nor U1804 (N_1804,In_717,In_538);
nand U1805 (N_1805,In_848,In_403);
and U1806 (N_1806,In_918,In_457);
and U1807 (N_1807,In_112,In_192);
and U1808 (N_1808,In_770,In_471);
and U1809 (N_1809,In_688,In_790);
and U1810 (N_1810,In_813,In_167);
nand U1811 (N_1811,In_53,In_603);
and U1812 (N_1812,In_295,In_268);
nand U1813 (N_1813,In_44,In_539);
and U1814 (N_1814,In_406,In_851);
or U1815 (N_1815,In_549,In_400);
nor U1816 (N_1816,In_537,In_584);
nand U1817 (N_1817,In_79,In_773);
nor U1818 (N_1818,In_256,In_44);
nand U1819 (N_1819,In_200,In_367);
or U1820 (N_1820,In_377,In_236);
or U1821 (N_1821,In_48,In_961);
nor U1822 (N_1822,In_334,In_189);
and U1823 (N_1823,In_281,In_571);
and U1824 (N_1824,In_69,In_726);
nand U1825 (N_1825,In_614,In_193);
and U1826 (N_1826,In_93,In_13);
or U1827 (N_1827,In_328,In_197);
and U1828 (N_1828,In_861,In_263);
or U1829 (N_1829,In_864,In_951);
or U1830 (N_1830,In_924,In_130);
nor U1831 (N_1831,In_766,In_832);
nor U1832 (N_1832,In_770,In_519);
or U1833 (N_1833,In_273,In_10);
or U1834 (N_1834,In_242,In_777);
or U1835 (N_1835,In_139,In_2);
nor U1836 (N_1836,In_718,In_685);
or U1837 (N_1837,In_112,In_717);
nor U1838 (N_1838,In_555,In_756);
and U1839 (N_1839,In_403,In_929);
nor U1840 (N_1840,In_895,In_687);
nor U1841 (N_1841,In_87,In_243);
nor U1842 (N_1842,In_351,In_851);
nand U1843 (N_1843,In_116,In_171);
nand U1844 (N_1844,In_959,In_198);
nand U1845 (N_1845,In_333,In_765);
nand U1846 (N_1846,In_284,In_781);
nand U1847 (N_1847,In_810,In_568);
nand U1848 (N_1848,In_128,In_305);
nor U1849 (N_1849,In_108,In_863);
or U1850 (N_1850,In_999,In_70);
nand U1851 (N_1851,In_24,In_642);
nand U1852 (N_1852,In_122,In_194);
and U1853 (N_1853,In_902,In_113);
nor U1854 (N_1854,In_774,In_742);
nand U1855 (N_1855,In_51,In_487);
nor U1856 (N_1856,In_998,In_769);
or U1857 (N_1857,In_53,In_96);
and U1858 (N_1858,In_17,In_816);
nor U1859 (N_1859,In_408,In_376);
or U1860 (N_1860,In_790,In_167);
or U1861 (N_1861,In_653,In_603);
nand U1862 (N_1862,In_386,In_287);
nor U1863 (N_1863,In_395,In_355);
or U1864 (N_1864,In_658,In_14);
or U1865 (N_1865,In_991,In_719);
nand U1866 (N_1866,In_890,In_441);
or U1867 (N_1867,In_598,In_973);
nand U1868 (N_1868,In_108,In_206);
nand U1869 (N_1869,In_909,In_886);
or U1870 (N_1870,In_907,In_126);
and U1871 (N_1871,In_852,In_777);
nor U1872 (N_1872,In_668,In_308);
nor U1873 (N_1873,In_789,In_7);
nand U1874 (N_1874,In_33,In_917);
xor U1875 (N_1875,In_572,In_379);
nor U1876 (N_1876,In_582,In_819);
nand U1877 (N_1877,In_996,In_197);
and U1878 (N_1878,In_12,In_502);
and U1879 (N_1879,In_738,In_951);
xor U1880 (N_1880,In_960,In_274);
and U1881 (N_1881,In_733,In_288);
or U1882 (N_1882,In_681,In_625);
or U1883 (N_1883,In_304,In_636);
nor U1884 (N_1884,In_72,In_851);
and U1885 (N_1885,In_991,In_950);
and U1886 (N_1886,In_562,In_444);
or U1887 (N_1887,In_994,In_332);
nand U1888 (N_1888,In_653,In_677);
or U1889 (N_1889,In_159,In_331);
or U1890 (N_1890,In_81,In_932);
or U1891 (N_1891,In_198,In_956);
or U1892 (N_1892,In_154,In_283);
or U1893 (N_1893,In_661,In_595);
nand U1894 (N_1894,In_740,In_378);
or U1895 (N_1895,In_298,In_883);
and U1896 (N_1896,In_203,In_982);
and U1897 (N_1897,In_803,In_403);
and U1898 (N_1898,In_427,In_62);
and U1899 (N_1899,In_176,In_317);
and U1900 (N_1900,In_834,In_513);
nor U1901 (N_1901,In_852,In_563);
and U1902 (N_1902,In_622,In_339);
and U1903 (N_1903,In_563,In_729);
or U1904 (N_1904,In_464,In_779);
nand U1905 (N_1905,In_289,In_975);
or U1906 (N_1906,In_460,In_20);
or U1907 (N_1907,In_665,In_453);
xor U1908 (N_1908,In_425,In_176);
xnor U1909 (N_1909,In_904,In_646);
or U1910 (N_1910,In_828,In_301);
and U1911 (N_1911,In_164,In_452);
nand U1912 (N_1912,In_228,In_177);
nand U1913 (N_1913,In_13,In_634);
and U1914 (N_1914,In_654,In_832);
and U1915 (N_1915,In_192,In_994);
and U1916 (N_1916,In_811,In_477);
and U1917 (N_1917,In_689,In_392);
nor U1918 (N_1918,In_299,In_186);
nand U1919 (N_1919,In_769,In_347);
nor U1920 (N_1920,In_159,In_528);
and U1921 (N_1921,In_109,In_354);
or U1922 (N_1922,In_700,In_998);
xor U1923 (N_1923,In_993,In_277);
and U1924 (N_1924,In_522,In_844);
nand U1925 (N_1925,In_857,In_920);
nor U1926 (N_1926,In_247,In_728);
nand U1927 (N_1927,In_562,In_948);
nor U1928 (N_1928,In_887,In_408);
or U1929 (N_1929,In_818,In_302);
and U1930 (N_1930,In_19,In_715);
nor U1931 (N_1931,In_118,In_768);
or U1932 (N_1932,In_872,In_932);
or U1933 (N_1933,In_29,In_212);
and U1934 (N_1934,In_588,In_332);
nor U1935 (N_1935,In_392,In_507);
and U1936 (N_1936,In_30,In_810);
and U1937 (N_1937,In_588,In_987);
or U1938 (N_1938,In_496,In_680);
or U1939 (N_1939,In_212,In_51);
nor U1940 (N_1940,In_804,In_843);
nor U1941 (N_1941,In_140,In_872);
nor U1942 (N_1942,In_201,In_503);
nor U1943 (N_1943,In_300,In_80);
nand U1944 (N_1944,In_265,In_904);
and U1945 (N_1945,In_190,In_308);
nand U1946 (N_1946,In_587,In_639);
nor U1947 (N_1947,In_41,In_754);
and U1948 (N_1948,In_475,In_403);
nand U1949 (N_1949,In_231,In_121);
or U1950 (N_1950,In_729,In_149);
nor U1951 (N_1951,In_705,In_978);
nand U1952 (N_1952,In_208,In_923);
or U1953 (N_1953,In_569,In_661);
nand U1954 (N_1954,In_827,In_362);
nand U1955 (N_1955,In_480,In_735);
and U1956 (N_1956,In_827,In_371);
nand U1957 (N_1957,In_422,In_101);
and U1958 (N_1958,In_584,In_363);
nand U1959 (N_1959,In_664,In_158);
nand U1960 (N_1960,In_639,In_961);
nor U1961 (N_1961,In_629,In_808);
and U1962 (N_1962,In_312,In_248);
or U1963 (N_1963,In_535,In_118);
nor U1964 (N_1964,In_9,In_643);
and U1965 (N_1965,In_568,In_661);
nand U1966 (N_1966,In_485,In_45);
and U1967 (N_1967,In_957,In_513);
and U1968 (N_1968,In_818,In_253);
nand U1969 (N_1969,In_587,In_598);
or U1970 (N_1970,In_774,In_312);
or U1971 (N_1971,In_53,In_293);
nand U1972 (N_1972,In_220,In_489);
nor U1973 (N_1973,In_461,In_62);
or U1974 (N_1974,In_960,In_90);
or U1975 (N_1975,In_881,In_582);
nor U1976 (N_1976,In_962,In_879);
or U1977 (N_1977,In_197,In_7);
or U1978 (N_1978,In_844,In_883);
nand U1979 (N_1979,In_998,In_691);
xnor U1980 (N_1980,In_360,In_553);
or U1981 (N_1981,In_568,In_963);
and U1982 (N_1982,In_561,In_908);
or U1983 (N_1983,In_764,In_551);
nor U1984 (N_1984,In_745,In_203);
or U1985 (N_1985,In_653,In_747);
nor U1986 (N_1986,In_24,In_876);
or U1987 (N_1987,In_417,In_366);
and U1988 (N_1988,In_295,In_891);
nor U1989 (N_1989,In_949,In_175);
nand U1990 (N_1990,In_897,In_223);
nand U1991 (N_1991,In_359,In_489);
nand U1992 (N_1992,In_761,In_617);
nand U1993 (N_1993,In_685,In_224);
or U1994 (N_1994,In_35,In_554);
nand U1995 (N_1995,In_32,In_955);
nor U1996 (N_1996,In_720,In_226);
nand U1997 (N_1997,In_246,In_438);
and U1998 (N_1998,In_29,In_993);
nor U1999 (N_1999,In_505,In_215);
nand U2000 (N_2000,In_67,In_687);
nor U2001 (N_2001,In_46,In_818);
and U2002 (N_2002,In_974,In_97);
nor U2003 (N_2003,In_112,In_343);
or U2004 (N_2004,In_216,In_965);
nor U2005 (N_2005,In_729,In_998);
nand U2006 (N_2006,In_584,In_423);
or U2007 (N_2007,In_166,In_830);
or U2008 (N_2008,In_774,In_978);
nor U2009 (N_2009,In_177,In_912);
or U2010 (N_2010,In_800,In_146);
or U2011 (N_2011,In_686,In_836);
nand U2012 (N_2012,In_33,In_969);
or U2013 (N_2013,In_282,In_554);
nand U2014 (N_2014,In_485,In_775);
nor U2015 (N_2015,In_227,In_135);
nand U2016 (N_2016,In_513,In_939);
nand U2017 (N_2017,In_535,In_326);
nor U2018 (N_2018,In_160,In_991);
and U2019 (N_2019,In_157,In_301);
nand U2020 (N_2020,In_244,In_176);
or U2021 (N_2021,In_938,In_512);
nor U2022 (N_2022,In_898,In_974);
and U2023 (N_2023,In_838,In_414);
and U2024 (N_2024,In_310,In_925);
nand U2025 (N_2025,In_10,In_336);
nand U2026 (N_2026,In_173,In_910);
nand U2027 (N_2027,In_603,In_883);
and U2028 (N_2028,In_788,In_610);
and U2029 (N_2029,In_19,In_420);
and U2030 (N_2030,In_852,In_681);
nor U2031 (N_2031,In_968,In_882);
or U2032 (N_2032,In_937,In_213);
and U2033 (N_2033,In_370,In_545);
nor U2034 (N_2034,In_444,In_136);
nand U2035 (N_2035,In_750,In_180);
and U2036 (N_2036,In_995,In_310);
and U2037 (N_2037,In_229,In_159);
xor U2038 (N_2038,In_98,In_76);
and U2039 (N_2039,In_370,In_600);
and U2040 (N_2040,In_279,In_150);
nand U2041 (N_2041,In_256,In_742);
or U2042 (N_2042,In_142,In_971);
and U2043 (N_2043,In_642,In_729);
or U2044 (N_2044,In_986,In_521);
nor U2045 (N_2045,In_103,In_163);
and U2046 (N_2046,In_233,In_753);
or U2047 (N_2047,In_577,In_675);
nand U2048 (N_2048,In_807,In_318);
and U2049 (N_2049,In_584,In_848);
nor U2050 (N_2050,In_187,In_381);
nor U2051 (N_2051,In_461,In_872);
nand U2052 (N_2052,In_667,In_432);
nor U2053 (N_2053,In_127,In_139);
nor U2054 (N_2054,In_63,In_766);
nor U2055 (N_2055,In_352,In_654);
or U2056 (N_2056,In_499,In_551);
nand U2057 (N_2057,In_214,In_766);
nand U2058 (N_2058,In_571,In_737);
or U2059 (N_2059,In_301,In_374);
nor U2060 (N_2060,In_936,In_266);
nor U2061 (N_2061,In_239,In_245);
nor U2062 (N_2062,In_252,In_917);
and U2063 (N_2063,In_509,In_741);
or U2064 (N_2064,In_981,In_720);
nand U2065 (N_2065,In_146,In_0);
xor U2066 (N_2066,In_55,In_435);
nor U2067 (N_2067,In_64,In_796);
and U2068 (N_2068,In_271,In_94);
or U2069 (N_2069,In_785,In_832);
nor U2070 (N_2070,In_16,In_858);
or U2071 (N_2071,In_885,In_950);
and U2072 (N_2072,In_507,In_625);
or U2073 (N_2073,In_419,In_152);
nor U2074 (N_2074,In_253,In_16);
nand U2075 (N_2075,In_307,In_947);
or U2076 (N_2076,In_458,In_98);
and U2077 (N_2077,In_879,In_860);
nand U2078 (N_2078,In_77,In_990);
or U2079 (N_2079,In_785,In_538);
xnor U2080 (N_2080,In_996,In_131);
nand U2081 (N_2081,In_332,In_342);
and U2082 (N_2082,In_770,In_647);
and U2083 (N_2083,In_823,In_510);
and U2084 (N_2084,In_128,In_734);
or U2085 (N_2085,In_599,In_968);
nor U2086 (N_2086,In_387,In_775);
or U2087 (N_2087,In_251,In_951);
or U2088 (N_2088,In_223,In_409);
nand U2089 (N_2089,In_609,In_447);
and U2090 (N_2090,In_903,In_687);
nand U2091 (N_2091,In_461,In_691);
xnor U2092 (N_2092,In_275,In_157);
or U2093 (N_2093,In_884,In_899);
and U2094 (N_2094,In_484,In_656);
nor U2095 (N_2095,In_926,In_146);
nand U2096 (N_2096,In_284,In_883);
xor U2097 (N_2097,In_175,In_264);
and U2098 (N_2098,In_905,In_12);
nand U2099 (N_2099,In_166,In_633);
or U2100 (N_2100,In_756,In_817);
nor U2101 (N_2101,In_733,In_462);
nand U2102 (N_2102,In_631,In_549);
nor U2103 (N_2103,In_466,In_307);
nor U2104 (N_2104,In_151,In_775);
and U2105 (N_2105,In_892,In_103);
nand U2106 (N_2106,In_883,In_397);
nand U2107 (N_2107,In_207,In_1);
xor U2108 (N_2108,In_235,In_26);
nor U2109 (N_2109,In_57,In_65);
and U2110 (N_2110,In_816,In_118);
nor U2111 (N_2111,In_413,In_261);
and U2112 (N_2112,In_74,In_490);
and U2113 (N_2113,In_587,In_665);
and U2114 (N_2114,In_2,In_83);
and U2115 (N_2115,In_289,In_817);
nor U2116 (N_2116,In_576,In_695);
nor U2117 (N_2117,In_281,In_745);
nor U2118 (N_2118,In_393,In_198);
nor U2119 (N_2119,In_831,In_169);
or U2120 (N_2120,In_927,In_160);
nand U2121 (N_2121,In_396,In_541);
nor U2122 (N_2122,In_784,In_398);
and U2123 (N_2123,In_860,In_798);
nand U2124 (N_2124,In_190,In_987);
and U2125 (N_2125,In_424,In_582);
nor U2126 (N_2126,In_588,In_855);
and U2127 (N_2127,In_312,In_632);
nor U2128 (N_2128,In_328,In_586);
nand U2129 (N_2129,In_951,In_422);
or U2130 (N_2130,In_648,In_30);
nand U2131 (N_2131,In_784,In_283);
nor U2132 (N_2132,In_637,In_19);
and U2133 (N_2133,In_621,In_906);
and U2134 (N_2134,In_807,In_161);
nor U2135 (N_2135,In_384,In_575);
or U2136 (N_2136,In_2,In_257);
or U2137 (N_2137,In_235,In_343);
and U2138 (N_2138,In_439,In_677);
and U2139 (N_2139,In_135,In_168);
nand U2140 (N_2140,In_531,In_139);
nor U2141 (N_2141,In_257,In_672);
nor U2142 (N_2142,In_247,In_403);
or U2143 (N_2143,In_361,In_295);
or U2144 (N_2144,In_530,In_58);
nand U2145 (N_2145,In_518,In_147);
or U2146 (N_2146,In_223,In_581);
nor U2147 (N_2147,In_851,In_776);
and U2148 (N_2148,In_463,In_372);
nor U2149 (N_2149,In_871,In_467);
nand U2150 (N_2150,In_145,In_751);
nor U2151 (N_2151,In_568,In_330);
and U2152 (N_2152,In_843,In_979);
or U2153 (N_2153,In_969,In_71);
xnor U2154 (N_2154,In_325,In_477);
or U2155 (N_2155,In_537,In_156);
nor U2156 (N_2156,In_744,In_84);
nand U2157 (N_2157,In_386,In_816);
or U2158 (N_2158,In_453,In_872);
nor U2159 (N_2159,In_464,In_862);
nand U2160 (N_2160,In_157,In_782);
or U2161 (N_2161,In_393,In_459);
and U2162 (N_2162,In_798,In_895);
nand U2163 (N_2163,In_799,In_405);
or U2164 (N_2164,In_183,In_102);
nand U2165 (N_2165,In_144,In_672);
nand U2166 (N_2166,In_1,In_697);
or U2167 (N_2167,In_65,In_5);
and U2168 (N_2168,In_383,In_90);
or U2169 (N_2169,In_586,In_941);
nor U2170 (N_2170,In_354,In_389);
and U2171 (N_2171,In_886,In_724);
and U2172 (N_2172,In_390,In_450);
nor U2173 (N_2173,In_806,In_434);
nor U2174 (N_2174,In_390,In_100);
and U2175 (N_2175,In_841,In_235);
nand U2176 (N_2176,In_549,In_418);
or U2177 (N_2177,In_132,In_266);
and U2178 (N_2178,In_497,In_947);
nor U2179 (N_2179,In_686,In_942);
and U2180 (N_2180,In_531,In_543);
or U2181 (N_2181,In_93,In_789);
or U2182 (N_2182,In_880,In_352);
and U2183 (N_2183,In_231,In_510);
nor U2184 (N_2184,In_181,In_336);
or U2185 (N_2185,In_285,In_823);
and U2186 (N_2186,In_61,In_484);
or U2187 (N_2187,In_31,In_694);
nand U2188 (N_2188,In_548,In_448);
nand U2189 (N_2189,In_650,In_369);
and U2190 (N_2190,In_528,In_186);
and U2191 (N_2191,In_755,In_164);
and U2192 (N_2192,In_547,In_837);
or U2193 (N_2193,In_927,In_726);
nor U2194 (N_2194,In_206,In_266);
nor U2195 (N_2195,In_382,In_944);
nor U2196 (N_2196,In_211,In_880);
nor U2197 (N_2197,In_833,In_166);
xnor U2198 (N_2198,In_125,In_43);
nor U2199 (N_2199,In_949,In_211);
xnor U2200 (N_2200,In_466,In_170);
or U2201 (N_2201,In_657,In_612);
nand U2202 (N_2202,In_478,In_448);
and U2203 (N_2203,In_935,In_879);
nand U2204 (N_2204,In_875,In_262);
nand U2205 (N_2205,In_397,In_766);
xor U2206 (N_2206,In_714,In_601);
nand U2207 (N_2207,In_203,In_986);
and U2208 (N_2208,In_586,In_770);
nor U2209 (N_2209,In_145,In_685);
nor U2210 (N_2210,In_87,In_92);
and U2211 (N_2211,In_962,In_873);
nand U2212 (N_2212,In_107,In_106);
nand U2213 (N_2213,In_66,In_626);
or U2214 (N_2214,In_386,In_240);
nor U2215 (N_2215,In_168,In_568);
xor U2216 (N_2216,In_532,In_468);
or U2217 (N_2217,In_675,In_878);
and U2218 (N_2218,In_555,In_45);
nand U2219 (N_2219,In_984,In_848);
or U2220 (N_2220,In_483,In_894);
nor U2221 (N_2221,In_359,In_216);
or U2222 (N_2222,In_347,In_586);
nor U2223 (N_2223,In_483,In_17);
and U2224 (N_2224,In_742,In_745);
and U2225 (N_2225,In_31,In_109);
nor U2226 (N_2226,In_617,In_860);
nor U2227 (N_2227,In_858,In_778);
nor U2228 (N_2228,In_528,In_998);
or U2229 (N_2229,In_684,In_610);
and U2230 (N_2230,In_34,In_602);
nor U2231 (N_2231,In_107,In_842);
and U2232 (N_2232,In_526,In_24);
nand U2233 (N_2233,In_337,In_9);
nand U2234 (N_2234,In_182,In_230);
nor U2235 (N_2235,In_204,In_333);
nor U2236 (N_2236,In_155,In_437);
or U2237 (N_2237,In_624,In_977);
nor U2238 (N_2238,In_13,In_213);
nor U2239 (N_2239,In_259,In_74);
and U2240 (N_2240,In_434,In_684);
nor U2241 (N_2241,In_725,In_856);
and U2242 (N_2242,In_352,In_637);
nand U2243 (N_2243,In_639,In_749);
nand U2244 (N_2244,In_533,In_671);
or U2245 (N_2245,In_330,In_958);
nand U2246 (N_2246,In_15,In_591);
and U2247 (N_2247,In_62,In_183);
nor U2248 (N_2248,In_187,In_348);
nand U2249 (N_2249,In_426,In_757);
nand U2250 (N_2250,In_648,In_473);
nand U2251 (N_2251,In_624,In_399);
nor U2252 (N_2252,In_393,In_818);
nand U2253 (N_2253,In_874,In_32);
and U2254 (N_2254,In_678,In_733);
xor U2255 (N_2255,In_228,In_855);
xnor U2256 (N_2256,In_181,In_470);
nor U2257 (N_2257,In_328,In_243);
or U2258 (N_2258,In_101,In_914);
nand U2259 (N_2259,In_547,In_553);
nor U2260 (N_2260,In_315,In_799);
nand U2261 (N_2261,In_177,In_304);
and U2262 (N_2262,In_719,In_595);
or U2263 (N_2263,In_465,In_632);
nand U2264 (N_2264,In_153,In_213);
and U2265 (N_2265,In_303,In_453);
and U2266 (N_2266,In_422,In_678);
and U2267 (N_2267,In_434,In_683);
xor U2268 (N_2268,In_234,In_34);
xor U2269 (N_2269,In_728,In_577);
nand U2270 (N_2270,In_579,In_696);
nor U2271 (N_2271,In_18,In_516);
and U2272 (N_2272,In_118,In_249);
nand U2273 (N_2273,In_682,In_681);
nand U2274 (N_2274,In_345,In_828);
xnor U2275 (N_2275,In_726,In_11);
nand U2276 (N_2276,In_130,In_812);
nand U2277 (N_2277,In_983,In_299);
and U2278 (N_2278,In_74,In_896);
and U2279 (N_2279,In_866,In_266);
nor U2280 (N_2280,In_769,In_813);
and U2281 (N_2281,In_176,In_840);
or U2282 (N_2282,In_951,In_543);
nand U2283 (N_2283,In_14,In_161);
and U2284 (N_2284,In_473,In_518);
and U2285 (N_2285,In_30,In_273);
nand U2286 (N_2286,In_829,In_822);
and U2287 (N_2287,In_43,In_524);
or U2288 (N_2288,In_971,In_243);
or U2289 (N_2289,In_86,In_171);
nor U2290 (N_2290,In_467,In_691);
nor U2291 (N_2291,In_383,In_315);
or U2292 (N_2292,In_401,In_610);
or U2293 (N_2293,In_993,In_489);
nor U2294 (N_2294,In_979,In_154);
nand U2295 (N_2295,In_255,In_650);
or U2296 (N_2296,In_532,In_858);
nand U2297 (N_2297,In_946,In_395);
nand U2298 (N_2298,In_879,In_763);
nor U2299 (N_2299,In_363,In_467);
or U2300 (N_2300,In_299,In_866);
or U2301 (N_2301,In_653,In_950);
and U2302 (N_2302,In_32,In_527);
and U2303 (N_2303,In_570,In_893);
nor U2304 (N_2304,In_146,In_272);
and U2305 (N_2305,In_604,In_229);
nor U2306 (N_2306,In_591,In_253);
and U2307 (N_2307,In_496,In_319);
and U2308 (N_2308,In_506,In_260);
nand U2309 (N_2309,In_331,In_264);
nor U2310 (N_2310,In_334,In_820);
nand U2311 (N_2311,In_934,In_191);
nor U2312 (N_2312,In_789,In_672);
nand U2313 (N_2313,In_158,In_905);
and U2314 (N_2314,In_379,In_66);
nand U2315 (N_2315,In_833,In_425);
and U2316 (N_2316,In_584,In_922);
or U2317 (N_2317,In_237,In_451);
nand U2318 (N_2318,In_681,In_378);
nor U2319 (N_2319,In_467,In_621);
or U2320 (N_2320,In_324,In_649);
and U2321 (N_2321,In_254,In_541);
and U2322 (N_2322,In_18,In_994);
or U2323 (N_2323,In_777,In_123);
nand U2324 (N_2324,In_595,In_894);
and U2325 (N_2325,In_964,In_56);
nor U2326 (N_2326,In_67,In_379);
nand U2327 (N_2327,In_819,In_625);
nand U2328 (N_2328,In_873,In_140);
nand U2329 (N_2329,In_822,In_754);
nand U2330 (N_2330,In_817,In_854);
or U2331 (N_2331,In_836,In_424);
nand U2332 (N_2332,In_132,In_76);
and U2333 (N_2333,In_436,In_262);
nand U2334 (N_2334,In_626,In_636);
nand U2335 (N_2335,In_671,In_897);
and U2336 (N_2336,In_637,In_793);
nor U2337 (N_2337,In_230,In_280);
nor U2338 (N_2338,In_574,In_179);
nor U2339 (N_2339,In_364,In_757);
nor U2340 (N_2340,In_600,In_74);
nor U2341 (N_2341,In_940,In_905);
xor U2342 (N_2342,In_921,In_869);
nor U2343 (N_2343,In_305,In_756);
nor U2344 (N_2344,In_754,In_55);
nand U2345 (N_2345,In_276,In_774);
nor U2346 (N_2346,In_660,In_49);
or U2347 (N_2347,In_20,In_1);
or U2348 (N_2348,In_365,In_657);
nand U2349 (N_2349,In_448,In_365);
nor U2350 (N_2350,In_121,In_453);
nor U2351 (N_2351,In_68,In_239);
or U2352 (N_2352,In_575,In_243);
nand U2353 (N_2353,In_648,In_751);
or U2354 (N_2354,In_639,In_424);
nor U2355 (N_2355,In_111,In_770);
or U2356 (N_2356,In_882,In_538);
or U2357 (N_2357,In_179,In_721);
nand U2358 (N_2358,In_285,In_849);
and U2359 (N_2359,In_161,In_362);
and U2360 (N_2360,In_280,In_308);
nand U2361 (N_2361,In_256,In_196);
or U2362 (N_2362,In_287,In_989);
nand U2363 (N_2363,In_357,In_564);
nor U2364 (N_2364,In_442,In_544);
xor U2365 (N_2365,In_125,In_260);
nor U2366 (N_2366,In_216,In_637);
or U2367 (N_2367,In_870,In_406);
or U2368 (N_2368,In_326,In_451);
nor U2369 (N_2369,In_914,In_797);
nor U2370 (N_2370,In_619,In_730);
or U2371 (N_2371,In_708,In_318);
nor U2372 (N_2372,In_129,In_801);
or U2373 (N_2373,In_694,In_595);
xnor U2374 (N_2374,In_313,In_962);
nor U2375 (N_2375,In_174,In_206);
xor U2376 (N_2376,In_835,In_699);
or U2377 (N_2377,In_617,In_939);
or U2378 (N_2378,In_748,In_730);
nor U2379 (N_2379,In_592,In_161);
nor U2380 (N_2380,In_130,In_626);
or U2381 (N_2381,In_767,In_282);
and U2382 (N_2382,In_282,In_325);
nor U2383 (N_2383,In_0,In_918);
nor U2384 (N_2384,In_318,In_773);
and U2385 (N_2385,In_226,In_445);
nand U2386 (N_2386,In_846,In_784);
nand U2387 (N_2387,In_687,In_4);
or U2388 (N_2388,In_628,In_47);
nand U2389 (N_2389,In_185,In_709);
nand U2390 (N_2390,In_235,In_584);
nand U2391 (N_2391,In_301,In_492);
nand U2392 (N_2392,In_507,In_323);
nor U2393 (N_2393,In_367,In_724);
nand U2394 (N_2394,In_360,In_535);
nand U2395 (N_2395,In_621,In_633);
nand U2396 (N_2396,In_525,In_592);
nor U2397 (N_2397,In_962,In_112);
nand U2398 (N_2398,In_7,In_886);
or U2399 (N_2399,In_624,In_709);
xnor U2400 (N_2400,In_832,In_43);
or U2401 (N_2401,In_571,In_143);
and U2402 (N_2402,In_858,In_971);
nor U2403 (N_2403,In_211,In_202);
and U2404 (N_2404,In_776,In_102);
nand U2405 (N_2405,In_399,In_197);
or U2406 (N_2406,In_92,In_710);
nor U2407 (N_2407,In_681,In_836);
and U2408 (N_2408,In_23,In_275);
or U2409 (N_2409,In_689,In_959);
nor U2410 (N_2410,In_452,In_246);
nand U2411 (N_2411,In_462,In_835);
nand U2412 (N_2412,In_847,In_786);
nor U2413 (N_2413,In_661,In_636);
xor U2414 (N_2414,In_156,In_381);
and U2415 (N_2415,In_824,In_97);
nand U2416 (N_2416,In_175,In_255);
nand U2417 (N_2417,In_425,In_81);
nor U2418 (N_2418,In_48,In_531);
or U2419 (N_2419,In_400,In_425);
nand U2420 (N_2420,In_666,In_790);
and U2421 (N_2421,In_795,In_324);
and U2422 (N_2422,In_963,In_761);
nor U2423 (N_2423,In_209,In_458);
and U2424 (N_2424,In_825,In_349);
nand U2425 (N_2425,In_521,In_823);
nor U2426 (N_2426,In_812,In_520);
or U2427 (N_2427,In_633,In_898);
and U2428 (N_2428,In_227,In_46);
and U2429 (N_2429,In_928,In_702);
xnor U2430 (N_2430,In_69,In_142);
or U2431 (N_2431,In_593,In_733);
nor U2432 (N_2432,In_973,In_195);
and U2433 (N_2433,In_297,In_555);
nor U2434 (N_2434,In_32,In_128);
nor U2435 (N_2435,In_235,In_11);
or U2436 (N_2436,In_118,In_165);
or U2437 (N_2437,In_40,In_420);
or U2438 (N_2438,In_963,In_434);
xnor U2439 (N_2439,In_394,In_121);
and U2440 (N_2440,In_531,In_895);
nor U2441 (N_2441,In_115,In_676);
nand U2442 (N_2442,In_0,In_486);
or U2443 (N_2443,In_602,In_290);
and U2444 (N_2444,In_668,In_567);
nor U2445 (N_2445,In_461,In_548);
or U2446 (N_2446,In_379,In_95);
nand U2447 (N_2447,In_210,In_450);
or U2448 (N_2448,In_604,In_928);
and U2449 (N_2449,In_307,In_792);
and U2450 (N_2450,In_457,In_242);
or U2451 (N_2451,In_277,In_885);
and U2452 (N_2452,In_696,In_998);
or U2453 (N_2453,In_212,In_474);
nor U2454 (N_2454,In_447,In_781);
or U2455 (N_2455,In_883,In_304);
or U2456 (N_2456,In_140,In_458);
or U2457 (N_2457,In_977,In_637);
or U2458 (N_2458,In_729,In_995);
nor U2459 (N_2459,In_617,In_947);
nand U2460 (N_2460,In_294,In_828);
nand U2461 (N_2461,In_957,In_351);
nand U2462 (N_2462,In_789,In_243);
nor U2463 (N_2463,In_715,In_51);
nand U2464 (N_2464,In_822,In_647);
nor U2465 (N_2465,In_819,In_851);
or U2466 (N_2466,In_5,In_863);
or U2467 (N_2467,In_26,In_728);
and U2468 (N_2468,In_546,In_633);
nor U2469 (N_2469,In_650,In_223);
and U2470 (N_2470,In_620,In_553);
or U2471 (N_2471,In_861,In_153);
or U2472 (N_2472,In_52,In_871);
nand U2473 (N_2473,In_562,In_136);
nand U2474 (N_2474,In_563,In_513);
and U2475 (N_2475,In_90,In_527);
nand U2476 (N_2476,In_421,In_591);
xor U2477 (N_2477,In_5,In_618);
or U2478 (N_2478,In_476,In_487);
or U2479 (N_2479,In_45,In_302);
nand U2480 (N_2480,In_295,In_13);
or U2481 (N_2481,In_334,In_157);
nand U2482 (N_2482,In_738,In_344);
and U2483 (N_2483,In_441,In_53);
nand U2484 (N_2484,In_34,In_548);
or U2485 (N_2485,In_247,In_523);
and U2486 (N_2486,In_502,In_414);
or U2487 (N_2487,In_612,In_651);
or U2488 (N_2488,In_222,In_373);
nor U2489 (N_2489,In_590,In_635);
nor U2490 (N_2490,In_677,In_16);
nor U2491 (N_2491,In_624,In_852);
and U2492 (N_2492,In_988,In_22);
or U2493 (N_2493,In_965,In_575);
or U2494 (N_2494,In_187,In_357);
nand U2495 (N_2495,In_580,In_744);
nor U2496 (N_2496,In_994,In_696);
nor U2497 (N_2497,In_605,In_283);
nor U2498 (N_2498,In_246,In_44);
xor U2499 (N_2499,In_561,In_947);
and U2500 (N_2500,N_677,N_1610);
or U2501 (N_2501,N_37,N_168);
nand U2502 (N_2502,N_652,N_1499);
or U2503 (N_2503,N_854,N_115);
and U2504 (N_2504,N_1150,N_351);
and U2505 (N_2505,N_29,N_1240);
and U2506 (N_2506,N_1720,N_553);
nand U2507 (N_2507,N_1501,N_998);
nor U2508 (N_2508,N_1817,N_1505);
nor U2509 (N_2509,N_446,N_2164);
or U2510 (N_2510,N_188,N_147);
nand U2511 (N_2511,N_9,N_2107);
nand U2512 (N_2512,N_692,N_629);
and U2513 (N_2513,N_693,N_1);
and U2514 (N_2514,N_1184,N_559);
and U2515 (N_2515,N_1483,N_745);
nor U2516 (N_2516,N_1762,N_2313);
xor U2517 (N_2517,N_2077,N_1271);
nor U2518 (N_2518,N_2443,N_2275);
and U2519 (N_2519,N_1074,N_1747);
and U2520 (N_2520,N_1084,N_2398);
xor U2521 (N_2521,N_782,N_2475);
nor U2522 (N_2522,N_2427,N_1173);
nand U2523 (N_2523,N_1392,N_490);
nor U2524 (N_2524,N_1915,N_483);
or U2525 (N_2525,N_752,N_2408);
nand U2526 (N_2526,N_1045,N_1268);
nand U2527 (N_2527,N_1162,N_665);
nor U2528 (N_2528,N_2252,N_915);
and U2529 (N_2529,N_1295,N_167);
and U2530 (N_2530,N_2191,N_1220);
and U2531 (N_2531,N_2158,N_2295);
and U2532 (N_2532,N_2261,N_638);
nor U2533 (N_2533,N_862,N_2325);
and U2534 (N_2534,N_277,N_981);
nor U2535 (N_2535,N_697,N_1124);
or U2536 (N_2536,N_384,N_1684);
xor U2537 (N_2537,N_1893,N_2260);
or U2538 (N_2538,N_56,N_1207);
nor U2539 (N_2539,N_1116,N_1164);
and U2540 (N_2540,N_314,N_1971);
or U2541 (N_2541,N_1721,N_294);
xor U2542 (N_2542,N_235,N_17);
and U2543 (N_2543,N_511,N_2355);
nor U2544 (N_2544,N_2076,N_794);
nand U2545 (N_2545,N_1859,N_1813);
or U2546 (N_2546,N_518,N_2240);
and U2547 (N_2547,N_419,N_2133);
nor U2548 (N_2548,N_229,N_1427);
and U2549 (N_2549,N_424,N_1448);
or U2550 (N_2550,N_1515,N_2119);
and U2551 (N_2551,N_208,N_1791);
nor U2552 (N_2552,N_1739,N_2470);
and U2553 (N_2553,N_416,N_513);
nor U2554 (N_2554,N_20,N_1899);
and U2555 (N_2555,N_1956,N_868);
or U2556 (N_2556,N_1870,N_1988);
nor U2557 (N_2557,N_1619,N_703);
and U2558 (N_2558,N_2364,N_2236);
nand U2559 (N_2559,N_1790,N_1396);
or U2560 (N_2560,N_841,N_427);
nand U2561 (N_2561,N_1100,N_80);
xor U2562 (N_2562,N_1047,N_2173);
nor U2563 (N_2563,N_1332,N_939);
and U2564 (N_2564,N_395,N_1337);
nand U2565 (N_2565,N_1193,N_1259);
and U2566 (N_2566,N_1303,N_546);
or U2567 (N_2567,N_1649,N_273);
or U2568 (N_2568,N_564,N_1951);
or U2569 (N_2569,N_1874,N_1068);
nor U2570 (N_2570,N_912,N_334);
nor U2571 (N_2571,N_1981,N_690);
nor U2572 (N_2572,N_724,N_313);
and U2573 (N_2573,N_1211,N_775);
nand U2574 (N_2574,N_1954,N_886);
nor U2575 (N_2575,N_1135,N_820);
and U2576 (N_2576,N_1546,N_1522);
nand U2577 (N_2577,N_337,N_1370);
nand U2578 (N_2578,N_1149,N_287);
and U2579 (N_2579,N_89,N_741);
xor U2580 (N_2580,N_1907,N_2457);
and U2581 (N_2581,N_1103,N_2485);
or U2582 (N_2582,N_1117,N_1190);
or U2583 (N_2583,N_2310,N_1882);
nand U2584 (N_2584,N_73,N_2347);
nor U2585 (N_2585,N_1452,N_2346);
nand U2586 (N_2586,N_1247,N_975);
and U2587 (N_2587,N_1022,N_925);
nand U2588 (N_2588,N_2218,N_1051);
nand U2589 (N_2589,N_986,N_2028);
nand U2590 (N_2590,N_1126,N_1182);
xnor U2591 (N_2591,N_520,N_1714);
and U2592 (N_2592,N_2352,N_1895);
nand U2593 (N_2593,N_2014,N_579);
nand U2594 (N_2594,N_1146,N_1189);
and U2595 (N_2595,N_1717,N_1434);
nand U2596 (N_2596,N_2009,N_696);
nor U2597 (N_2597,N_1786,N_2113);
or U2598 (N_2598,N_792,N_270);
nand U2599 (N_2599,N_525,N_1497);
nand U2600 (N_2600,N_339,N_207);
nand U2601 (N_2601,N_620,N_1857);
nor U2602 (N_2602,N_461,N_736);
nand U2603 (N_2603,N_828,N_285);
nor U2604 (N_2604,N_815,N_2029);
or U2605 (N_2605,N_327,N_711);
nand U2606 (N_2606,N_2353,N_492);
nor U2607 (N_2607,N_2154,N_1287);
nand U2608 (N_2608,N_876,N_684);
nand U2609 (N_2609,N_2084,N_81);
or U2610 (N_2610,N_1770,N_1498);
xnor U2611 (N_2611,N_945,N_2401);
nor U2612 (N_2612,N_284,N_1925);
nor U2613 (N_2613,N_1234,N_421);
and U2614 (N_2614,N_1968,N_420);
nand U2615 (N_2615,N_197,N_1647);
nor U2616 (N_2616,N_642,N_305);
and U2617 (N_2617,N_1157,N_1339);
or U2618 (N_2618,N_1627,N_226);
nand U2619 (N_2619,N_1379,N_122);
nor U2620 (N_2620,N_687,N_1687);
or U2621 (N_2621,N_1447,N_2195);
nand U2622 (N_2622,N_1403,N_162);
or U2623 (N_2623,N_558,N_738);
and U2624 (N_2624,N_1300,N_1740);
or U2625 (N_2625,N_866,N_1322);
nand U2626 (N_2626,N_1722,N_163);
nand U2627 (N_2627,N_2375,N_2373);
or U2628 (N_2628,N_2326,N_1838);
nor U2629 (N_2629,N_1024,N_491);
nand U2630 (N_2630,N_1897,N_1556);
nor U2631 (N_2631,N_2230,N_2008);
nand U2632 (N_2632,N_610,N_364);
nor U2633 (N_2633,N_574,N_2016);
nand U2634 (N_2634,N_2374,N_917);
and U2635 (N_2635,N_2189,N_402);
xor U2636 (N_2636,N_1602,N_2114);
and U2637 (N_2637,N_465,N_1911);
nand U2638 (N_2638,N_1436,N_1884);
or U2639 (N_2639,N_1382,N_1186);
nand U2640 (N_2640,N_845,N_799);
or U2641 (N_2641,N_1005,N_1282);
xor U2642 (N_2642,N_476,N_173);
nand U2643 (N_2643,N_904,N_2468);
or U2644 (N_2644,N_1554,N_398);
nand U2645 (N_2645,N_643,N_1594);
or U2646 (N_2646,N_2022,N_451);
nand U2647 (N_2647,N_2495,N_2391);
or U2648 (N_2648,N_1773,N_158);
nor U2649 (N_2649,N_460,N_808);
nand U2650 (N_2650,N_1690,N_1168);
or U2651 (N_2651,N_1523,N_1570);
and U2652 (N_2652,N_406,N_1187);
or U2653 (N_2653,N_869,N_1577);
and U2654 (N_2654,N_408,N_2176);
nor U2655 (N_2655,N_2273,N_437);
and U2656 (N_2656,N_457,N_189);
and U2657 (N_2657,N_706,N_341);
or U2658 (N_2658,N_2227,N_1469);
or U2659 (N_2659,N_1652,N_261);
nor U2660 (N_2660,N_219,N_35);
nor U2661 (N_2661,N_2099,N_1131);
nor U2662 (N_2662,N_2038,N_1534);
and U2663 (N_2663,N_463,N_1650);
or U2664 (N_2664,N_137,N_2472);
nand U2665 (N_2665,N_1997,N_1355);
and U2666 (N_2666,N_361,N_1945);
xnor U2667 (N_2667,N_433,N_1365);
nor U2668 (N_2668,N_654,N_681);
or U2669 (N_2669,N_621,N_119);
or U2670 (N_2670,N_443,N_2423);
or U2671 (N_2671,N_2212,N_963);
or U2672 (N_2672,N_1450,N_2267);
or U2673 (N_2673,N_99,N_2349);
nor U2674 (N_2674,N_1063,N_771);
nand U2675 (N_2675,N_24,N_1584);
or U2676 (N_2676,N_1004,N_2378);
and U2677 (N_2677,N_1357,N_565);
nor U2678 (N_2678,N_829,N_425);
nand U2679 (N_2679,N_2024,N_2106);
or U2680 (N_2680,N_1194,N_107);
nor U2681 (N_2681,N_383,N_2455);
nor U2682 (N_2682,N_1175,N_2416);
and U2683 (N_2683,N_399,N_1449);
or U2684 (N_2684,N_202,N_2396);
nand U2685 (N_2685,N_2220,N_1973);
and U2686 (N_2686,N_1031,N_573);
nor U2687 (N_2687,N_2226,N_267);
nand U2688 (N_2688,N_589,N_851);
and U2689 (N_2689,N_781,N_220);
nand U2690 (N_2690,N_1703,N_1646);
and U2691 (N_2691,N_1206,N_861);
or U2692 (N_2692,N_1408,N_2318);
nor U2693 (N_2693,N_744,N_69);
or U2694 (N_2694,N_946,N_787);
or U2695 (N_2695,N_1625,N_2307);
and U2696 (N_2696,N_1623,N_166);
nor U2697 (N_2697,N_153,N_2377);
or U2698 (N_2698,N_502,N_801);
nand U2699 (N_2699,N_1655,N_1353);
and U2700 (N_2700,N_2049,N_1604);
or U2701 (N_2701,N_675,N_8);
nor U2702 (N_2702,N_2225,N_836);
and U2703 (N_2703,N_682,N_1334);
and U2704 (N_2704,N_2253,N_1842);
and U2705 (N_2705,N_892,N_1454);
nand U2706 (N_2706,N_1112,N_2241);
nand U2707 (N_2707,N_901,N_536);
and U2708 (N_2708,N_822,N_250);
and U2709 (N_2709,N_2291,N_2388);
and U2710 (N_2710,N_499,N_2392);
and U2711 (N_2711,N_1597,N_1613);
or U2712 (N_2712,N_342,N_1261);
nor U2713 (N_2713,N_1136,N_2449);
nor U2714 (N_2714,N_1167,N_2292);
nor U2715 (N_2715,N_2342,N_2075);
nand U2716 (N_2716,N_805,N_10);
and U2717 (N_2717,N_1744,N_432);
and U2718 (N_2718,N_2451,N_846);
nand U2719 (N_2719,N_1503,N_1344);
nand U2720 (N_2720,N_345,N_1772);
nor U2721 (N_2721,N_2209,N_193);
nand U2722 (N_2722,N_1735,N_903);
nand U2723 (N_2723,N_1886,N_1587);
nor U2724 (N_2724,N_1305,N_1072);
nand U2725 (N_2725,N_1672,N_1667);
and U2726 (N_2726,N_1898,N_428);
nor U2727 (N_2727,N_1089,N_2067);
and U2728 (N_2728,N_616,N_1768);
and U2729 (N_2729,N_462,N_108);
nor U2730 (N_2730,N_377,N_2040);
nand U2731 (N_2731,N_210,N_1306);
nand U2732 (N_2732,N_375,N_1196);
and U2733 (N_2733,N_369,N_2183);
and U2734 (N_2734,N_271,N_1576);
and U2735 (N_2735,N_1432,N_1979);
and U2736 (N_2736,N_512,N_30);
or U2737 (N_2737,N_709,N_1866);
nand U2738 (N_2738,N_391,N_1535);
or U2739 (N_2739,N_1977,N_1351);
nand U2740 (N_2740,N_1742,N_647);
and U2741 (N_2741,N_130,N_410);
or U2742 (N_2742,N_2320,N_1926);
and U2743 (N_2743,N_1476,N_2399);
nand U2744 (N_2744,N_1118,N_947);
and U2745 (N_2745,N_1170,N_883);
or U2746 (N_2746,N_57,N_544);
and U2747 (N_2747,N_730,N_1950);
or U2748 (N_2748,N_2414,N_1707);
or U2749 (N_2749,N_548,N_1317);
and U2750 (N_2750,N_1413,N_1709);
nand U2751 (N_2751,N_1308,N_1481);
nand U2752 (N_2752,N_1525,N_1936);
nand U2753 (N_2753,N_206,N_774);
nand U2754 (N_2754,N_1976,N_1127);
and U2755 (N_2755,N_485,N_1388);
nor U2756 (N_2756,N_1280,N_1151);
or U2757 (N_2757,N_1083,N_1283);
nand U2758 (N_2758,N_458,N_2324);
and U2759 (N_2759,N_877,N_2441);
and U2760 (N_2760,N_218,N_1488);
and U2761 (N_2761,N_940,N_2498);
or U2762 (N_2762,N_177,N_387);
nand U2763 (N_2763,N_603,N_454);
xnor U2764 (N_2764,N_2034,N_1502);
nand U2765 (N_2765,N_409,N_2413);
or U2766 (N_2766,N_1257,N_1991);
nor U2767 (N_2767,N_117,N_810);
or U2768 (N_2768,N_326,N_749);
nand U2769 (N_2769,N_1464,N_1374);
and U2770 (N_2770,N_2315,N_2163);
nor U2771 (N_2771,N_2434,N_1209);
nor U2772 (N_2772,N_870,N_186);
nor U2773 (N_2773,N_411,N_1037);
or U2774 (N_2774,N_816,N_1730);
or U2775 (N_2775,N_1508,N_129);
and U2776 (N_2776,N_832,N_98);
nor U2777 (N_2777,N_32,N_660);
nand U2778 (N_2778,N_2060,N_386);
or U2779 (N_2779,N_2115,N_2234);
or U2780 (N_2780,N_1021,N_1957);
or U2781 (N_2781,N_1201,N_1756);
xor U2782 (N_2782,N_2268,N_1301);
or U2783 (N_2783,N_614,N_1643);
nor U2784 (N_2784,N_1548,N_1656);
or U2785 (N_2785,N_2361,N_389);
nand U2786 (N_2786,N_545,N_679);
nand U2787 (N_2787,N_255,N_560);
nor U2788 (N_2788,N_97,N_2281);
and U2789 (N_2789,N_1949,N_1266);
or U2790 (N_2790,N_160,N_1496);
nor U2791 (N_2791,N_2190,N_254);
or U2792 (N_2792,N_1273,N_849);
xor U2793 (N_2793,N_2116,N_101);
nor U2794 (N_2794,N_1941,N_2161);
nor U2795 (N_2795,N_817,N_1964);
nor U2796 (N_2796,N_2004,N_1539);
or U2797 (N_2797,N_2358,N_127);
or U2798 (N_2798,N_2186,N_2322);
nor U2799 (N_2799,N_1439,N_1329);
and U2800 (N_2800,N_1485,N_1837);
or U2801 (N_2801,N_65,N_954);
nor U2802 (N_2802,N_2258,N_2194);
nor U2803 (N_2803,N_1142,N_2323);
and U2804 (N_2804,N_655,N_1676);
and U2805 (N_2805,N_2270,N_23);
nand U2806 (N_2806,N_936,N_2182);
and U2807 (N_2807,N_2211,N_2152);
nor U2808 (N_2808,N_215,N_2277);
nor U2809 (N_2809,N_6,N_2370);
and U2810 (N_2810,N_1620,N_312);
nand U2811 (N_2811,N_648,N_456);
or U2812 (N_2812,N_62,N_2006);
nor U2813 (N_2813,N_1120,N_1137);
or U2814 (N_2814,N_1461,N_1455);
nand U2815 (N_2815,N_2481,N_1671);
nor U2816 (N_2816,N_1494,N_282);
and U2817 (N_2817,N_2052,N_174);
nor U2818 (N_2818,N_1575,N_960);
and U2819 (N_2819,N_1460,N_2274);
nand U2820 (N_2820,N_2136,N_1122);
nor U2821 (N_2821,N_1012,N_1512);
or U2822 (N_2822,N_1519,N_1585);
nor U2823 (N_2823,N_2365,N_713);
xor U2824 (N_2824,N_987,N_990);
xor U2825 (N_2825,N_691,N_2096);
nand U2826 (N_2826,N_1718,N_1477);
or U2827 (N_2827,N_673,N_2493);
nand U2828 (N_2828,N_723,N_796);
nand U2829 (N_2829,N_113,N_1996);
or U2830 (N_2830,N_1631,N_2108);
and U2831 (N_2831,N_2012,N_1390);
or U2832 (N_2832,N_1727,N_786);
nor U2833 (N_2833,N_628,N_2421);
or U2834 (N_2834,N_258,N_2184);
or U2835 (N_2835,N_1737,N_1542);
nand U2836 (N_2836,N_1028,N_2490);
or U2837 (N_2837,N_125,N_2231);
nand U2838 (N_2838,N_973,N_916);
nor U2839 (N_2839,N_1389,N_145);
or U2840 (N_2840,N_1098,N_2003);
or U2841 (N_2841,N_957,N_1299);
or U2842 (N_2842,N_1563,N_1386);
or U2843 (N_2843,N_1087,N_529);
and U2844 (N_2844,N_2185,N_809);
nor U2845 (N_2845,N_216,N_1807);
and U2846 (N_2846,N_1891,N_1352);
and U2847 (N_2847,N_1090,N_1759);
nor U2848 (N_2848,N_1480,N_1555);
and U2849 (N_2849,N_1376,N_76);
nand U2850 (N_2850,N_445,N_1212);
nand U2851 (N_2851,N_155,N_1075);
nand U2852 (N_2852,N_134,N_847);
or U2853 (N_2853,N_171,N_328);
and U2854 (N_2854,N_2299,N_1179);
nand U2855 (N_2855,N_2444,N_2247);
and U2856 (N_2856,N_2263,N_1139);
or U2857 (N_2857,N_1743,N_121);
or U2858 (N_2858,N_169,N_2197);
or U2859 (N_2859,N_279,N_1222);
nor U2860 (N_2860,N_1582,N_31);
xnor U2861 (N_2861,N_622,N_2426);
nor U2862 (N_2862,N_1350,N_2025);
and U2863 (N_2863,N_2351,N_1492);
nor U2864 (N_2864,N_1517,N_1583);
nand U2865 (N_2865,N_2249,N_209);
or U2866 (N_2866,N_349,N_1158);
or U2867 (N_2867,N_1552,N_898);
nor U2868 (N_2868,N_13,N_2193);
nand U2869 (N_2869,N_1433,N_2178);
and U2870 (N_2870,N_2327,N_355);
nor U2871 (N_2871,N_2105,N_1110);
nand U2872 (N_2872,N_467,N_1890);
nor U2873 (N_2873,N_1990,N_1699);
or U2874 (N_2874,N_2201,N_600);
and U2875 (N_2875,N_1387,N_1532);
or U2876 (N_2876,N_2454,N_1061);
and U2877 (N_2877,N_299,N_2089);
nand U2878 (N_2878,N_1446,N_1705);
and U2879 (N_2879,N_561,N_950);
nor U2880 (N_2880,N_430,N_1046);
xor U2881 (N_2881,N_2438,N_1441);
nor U2882 (N_2882,N_840,N_2149);
nor U2883 (N_2883,N_2330,N_1260);
and U2884 (N_2884,N_140,N_1371);
and U2885 (N_2885,N_434,N_1984);
and U2886 (N_2886,N_2479,N_602);
and U2887 (N_2887,N_2476,N_199);
or U2888 (N_2888,N_1040,N_2050);
nand U2889 (N_2889,N_1787,N_1632);
or U2890 (N_2890,N_1798,N_754);
or U2891 (N_2891,N_857,N_949);
and U2892 (N_2892,N_1783,N_984);
or U2893 (N_2893,N_2367,N_2376);
and U2894 (N_2894,N_790,N_1733);
nand U2895 (N_2895,N_1141,N_783);
and U2896 (N_2896,N_1873,N_1020);
or U2897 (N_2897,N_1358,N_758);
nand U2898 (N_2898,N_1549,N_2290);
nand U2899 (N_2899,N_1589,N_1816);
nand U2900 (N_2900,N_595,N_1169);
nand U2901 (N_2901,N_1777,N_1292);
and U2902 (N_2902,N_2257,N_1054);
nor U2903 (N_2903,N_1825,N_615);
and U2904 (N_2904,N_370,N_2222);
nand U2905 (N_2905,N_2354,N_860);
nand U2906 (N_2906,N_1385,N_767);
and U2907 (N_2907,N_1393,N_569);
and U2908 (N_2908,N_47,N_1581);
nor U2909 (N_2909,N_380,N_1682);
or U2910 (N_2910,N_2357,N_1302);
nor U2911 (N_2911,N_1239,N_1741);
or U2912 (N_2912,N_42,N_248);
nor U2913 (N_2913,N_373,N_934);
and U2914 (N_2914,N_1797,N_2272);
nand U2915 (N_2915,N_2420,N_1147);
or U2916 (N_2916,N_1152,N_138);
or U2917 (N_2917,N_2360,N_2435);
and U2918 (N_2918,N_367,N_2098);
and U2919 (N_2919,N_2289,N_1654);
or U2920 (N_2920,N_930,N_1544);
or U2921 (N_2921,N_1442,N_286);
or U2922 (N_2922,N_1562,N_606);
nand U2923 (N_2923,N_1011,N_2037);
and U2924 (N_2924,N_1263,N_1067);
and U2925 (N_2925,N_1466,N_1105);
or U2926 (N_2926,N_2431,N_952);
nor U2927 (N_2927,N_2035,N_1509);
nor U2928 (N_2928,N_444,N_2350);
and U2929 (N_2929,N_196,N_944);
nand U2930 (N_2930,N_1608,N_1368);
and U2931 (N_2931,N_2255,N_830);
and U2932 (N_2932,N_969,N_797);
nor U2933 (N_2933,N_888,N_1799);
and U2934 (N_2934,N_1989,N_1923);
and U2935 (N_2935,N_422,N_1865);
nor U2936 (N_2936,N_92,N_2418);
or U2937 (N_2937,N_769,N_539);
nor U2938 (N_2938,N_1943,N_1789);
or U2939 (N_2939,N_1500,N_228);
nor U2940 (N_2940,N_268,N_532);
and U2941 (N_2941,N_1177,N_149);
or U2942 (N_2942,N_203,N_322);
nand U2943 (N_2943,N_612,N_1086);
xor U2944 (N_2944,N_1267,N_70);
and U2945 (N_2945,N_1250,N_2244);
nor U2946 (N_2946,N_743,N_566);
nand U2947 (N_2947,N_1041,N_996);
and U2948 (N_2948,N_1114,N_1644);
nand U2949 (N_2949,N_720,N_1414);
xor U2950 (N_2950,N_1993,N_1806);
nor U2951 (N_2951,N_236,N_114);
nor U2952 (N_2952,N_1121,N_1888);
nor U2953 (N_2953,N_1119,N_2169);
and U2954 (N_2954,N_187,N_534);
and U2955 (N_2955,N_198,N_2065);
xnor U2956 (N_2956,N_2074,N_2316);
nand U2957 (N_2957,N_415,N_1073);
nand U2958 (N_2958,N_404,N_1183);
nand U2959 (N_2959,N_1291,N_2440);
nor U2960 (N_2960,N_2338,N_686);
or U2961 (N_2961,N_1590,N_2429);
or U2962 (N_2962,N_1198,N_2382);
or U2963 (N_2963,N_1420,N_1043);
nor U2964 (N_2964,N_85,N_2132);
and U2965 (N_2965,N_161,N_213);
nand U2966 (N_2966,N_897,N_1948);
and U2967 (N_2967,N_748,N_503);
nor U2968 (N_2968,N_727,N_1543);
nor U2969 (N_2969,N_2135,N_972);
and U2970 (N_2970,N_1814,N_568);
and U2971 (N_2971,N_1285,N_1077);
and U2972 (N_2972,N_1896,N_2469);
nor U2973 (N_2973,N_2383,N_1930);
or U2974 (N_2974,N_1680,N_78);
or U2975 (N_2975,N_1504,N_1975);
nand U2976 (N_2976,N_1421,N_110);
or U2977 (N_2977,N_133,N_2127);
nand U2978 (N_2978,N_1484,N_1960);
or U2979 (N_2979,N_1210,N_227);
or U2980 (N_2980,N_1635,N_14);
nor U2981 (N_2981,N_2073,N_1309);
nand U2982 (N_2982,N_357,N_626);
nor U2983 (N_2983,N_1673,N_1757);
and U2984 (N_2984,N_1140,N_2278);
or U2985 (N_2985,N_292,N_685);
nor U2986 (N_2986,N_1326,N_1881);
xnor U2987 (N_2987,N_2056,N_1732);
or U2988 (N_2988,N_1457,N_481);
nor U2989 (N_2989,N_935,N_1592);
and U2990 (N_2990,N_1846,N_1966);
or U2991 (N_2991,N_1629,N_195);
or U2992 (N_2992,N_1617,N_672);
or U2993 (N_2993,N_1324,N_19);
or U2994 (N_2994,N_1883,N_1172);
nor U2995 (N_2995,N_977,N_459);
or U2996 (N_2996,N_311,N_689);
nand U2997 (N_2997,N_699,N_895);
and U2998 (N_2998,N_2486,N_151);
and U2999 (N_2999,N_1033,N_1661);
xnor U3000 (N_3000,N_927,N_819);
and U3001 (N_3001,N_1223,N_750);
nor U3002 (N_3002,N_15,N_1998);
or U3003 (N_3003,N_838,N_1462);
or U3004 (N_3004,N_721,N_1758);
nand U3005 (N_3005,N_704,N_2117);
nand U3006 (N_3006,N_880,N_1510);
or U3007 (N_3007,N_701,N_1148);
nor U3008 (N_3008,N_2464,N_397);
or U3009 (N_3009,N_1363,N_496);
or U3010 (N_3010,N_575,N_1565);
and U3011 (N_3011,N_1176,N_111);
and U3012 (N_3012,N_1858,N_1224);
nor U3013 (N_3013,N_2057,N_1373);
nor U3014 (N_3014,N_494,N_2199);
nand U3015 (N_3015,N_1161,N_429);
or U3016 (N_3016,N_1475,N_1834);
and U3017 (N_3017,N_757,N_1252);
xnor U3018 (N_3018,N_1754,N_2344);
nor U3019 (N_3019,N_2140,N_1079);
and U3020 (N_3020,N_656,N_1228);
nor U3021 (N_3021,N_1713,N_359);
and U3022 (N_3022,N_1875,N_1335);
and U3023 (N_3023,N_994,N_2482);
and U3024 (N_3024,N_1013,N_1286);
or U3025 (N_3025,N_1264,N_298);
or U3026 (N_3026,N_2083,N_2109);
nand U3027 (N_3027,N_1346,N_2433);
or U3028 (N_3028,N_530,N_666);
or U3029 (N_3029,N_1249,N_453);
nor U3030 (N_3030,N_1793,N_1006);
nor U3031 (N_3031,N_2062,N_2203);
nor U3032 (N_3032,N_1430,N_2013);
and U3033 (N_3033,N_863,N_2243);
and U3034 (N_3034,N_2000,N_584);
nand U3035 (N_3035,N_1014,N_853);
nor U3036 (N_3036,N_1571,N_1422);
nand U3037 (N_3037,N_2393,N_142);
nand U3038 (N_3038,N_617,N_1812);
and U3039 (N_3039,N_1708,N_2412);
or U3040 (N_3040,N_1924,N_242);
and U3041 (N_3041,N_2110,N_1513);
or U3042 (N_3042,N_551,N_1218);
nor U3043 (N_3043,N_1561,N_906);
nand U3044 (N_3044,N_1236,N_1288);
or U3045 (N_3045,N_1204,N_1809);
and U3046 (N_3046,N_1165,N_2410);
nand U3047 (N_3047,N_1628,N_442);
nor U3048 (N_3048,N_1001,N_2445);
and U3049 (N_3049,N_247,N_205);
nor U3050 (N_3050,N_2229,N_976);
nand U3051 (N_3051,N_1202,N_894);
and U3052 (N_3052,N_1530,N_1688);
or U3053 (N_3053,N_580,N_577);
or U3054 (N_3054,N_874,N_2285);
nor U3055 (N_3055,N_1066,N_61);
or U3056 (N_3056,N_1801,N_1569);
xnor U3057 (N_3057,N_105,N_1987);
nor U3058 (N_3058,N_761,N_1641);
nand U3059 (N_3059,N_321,N_478);
nand U3060 (N_3060,N_1974,N_1579);
nor U3061 (N_3061,N_265,N_2174);
and U3062 (N_3062,N_1251,N_1036);
and U3063 (N_3063,N_609,N_317);
nand U3064 (N_3064,N_2095,N_2343);
or U3065 (N_3065,N_651,N_953);
nand U3066 (N_3066,N_2124,N_583);
or U3067 (N_3067,N_2180,N_607);
and U3068 (N_3068,N_48,N_439);
and U3069 (N_3069,N_959,N_507);
and U3070 (N_3070,N_649,N_1419);
and U3071 (N_3071,N_150,N_765);
nand U3072 (N_3072,N_368,N_1440);
nand U3073 (N_3073,N_1319,N_1290);
nand U3074 (N_3074,N_505,N_394);
nand U3075 (N_3075,N_1473,N_143);
nor U3076 (N_3076,N_2463,N_1241);
or U3077 (N_3077,N_403,N_519);
nor U3078 (N_3078,N_928,N_477);
or U3079 (N_3079,N_1779,N_309);
and U3080 (N_3080,N_1701,N_1929);
or U3081 (N_3081,N_2088,N_1908);
or U3082 (N_3082,N_2499,N_1153);
nand U3083 (N_3083,N_962,N_238);
or U3084 (N_3084,N_346,N_1609);
nand U3085 (N_3085,N_1681,N_75);
nand U3086 (N_3086,N_135,N_1664);
or U3087 (N_3087,N_1944,N_96);
nor U3088 (N_3088,N_1685,N_1482);
and U3089 (N_3089,N_112,N_1521);
nand U3090 (N_3090,N_1640,N_1657);
nor U3091 (N_3091,N_1871,N_770);
nor U3092 (N_3092,N_2128,N_1231);
and U3093 (N_3093,N_448,N_588);
nor U3094 (N_3094,N_729,N_2092);
or U3095 (N_3095,N_438,N_1233);
and U3096 (N_3096,N_2415,N_2147);
or U3097 (N_3097,N_785,N_2284);
and U3098 (N_3098,N_2202,N_2172);
nand U3099 (N_3099,N_1246,N_2005);
or U3100 (N_3100,N_471,N_1428);
or U3101 (N_3101,N_1429,N_1861);
or U3102 (N_3102,N_1312,N_1424);
nand U3103 (N_3103,N_663,N_567);
and U3104 (N_3104,N_1443,N_1191);
or U3105 (N_3105,N_1621,N_126);
nand U3106 (N_3106,N_2453,N_72);
and U3107 (N_3107,N_2177,N_2337);
nor U3108 (N_3108,N_431,N_2080);
nor U3109 (N_3109,N_350,N_1227);
or U3110 (N_3110,N_807,N_1645);
or U3111 (N_3111,N_1918,N_995);
or U3112 (N_3112,N_1695,N_1614);
or U3113 (N_3113,N_979,N_964);
or U3114 (N_3114,N_181,N_683);
nand U3115 (N_3115,N_632,N_1827);
nand U3116 (N_3116,N_204,N_2221);
or U3117 (N_3117,N_1321,N_1174);
nor U3118 (N_3118,N_2122,N_831);
nand U3119 (N_3119,N_1524,N_777);
nand U3120 (N_3120,N_194,N_1533);
nand U3121 (N_3121,N_708,N_289);
or U3122 (N_3122,N_855,N_132);
and U3123 (N_3123,N_1106,N_1724);
and U3124 (N_3124,N_929,N_231);
nor U3125 (N_3125,N_224,N_902);
or U3126 (N_3126,N_1995,N_1712);
nor U3127 (N_3127,N_515,N_2126);
nor U3128 (N_3128,N_2321,N_93);
or U3129 (N_3129,N_1913,N_338);
and U3130 (N_3130,N_1912,N_637);
or U3131 (N_3131,N_1281,N_144);
or U3132 (N_3132,N_2042,N_909);
nor U3133 (N_3133,N_1205,N_372);
nand U3134 (N_3134,N_2015,N_2181);
or U3135 (N_3135,N_374,N_1885);
or U3136 (N_3136,N_1125,N_243);
and U3137 (N_3137,N_1752,N_1160);
nand U3138 (N_3138,N_1795,N_1983);
or U3139 (N_3139,N_2303,N_2026);
nor U3140 (N_3140,N_2264,N_154);
nor U3141 (N_3141,N_1381,N_1596);
and U3142 (N_3142,N_253,N_2217);
or U3143 (N_3143,N_2419,N_1145);
nor U3144 (N_3144,N_1289,N_378);
or U3145 (N_3145,N_966,N_1804);
or U3146 (N_3146,N_1573,N_867);
or U3147 (N_3147,N_39,N_2153);
or U3148 (N_3148,N_1719,N_1902);
or U3149 (N_3149,N_795,N_2093);
or U3150 (N_3150,N_232,N_657);
nor U3151 (N_3151,N_64,N_585);
or U3152 (N_3152,N_382,N_1959);
or U3153 (N_3153,N_234,N_2059);
and U3154 (N_3154,N_223,N_2130);
nor U3155 (N_3155,N_2452,N_1314);
nand U3156 (N_3156,N_2079,N_1972);
and U3157 (N_3157,N_535,N_1185);
nor U3158 (N_3158,N_1366,N_601);
nand U3159 (N_3159,N_2150,N_1316);
nand U3160 (N_3160,N_586,N_1952);
or U3161 (N_3161,N_1490,N_79);
or U3162 (N_3162,N_2379,N_734);
and U3163 (N_3163,N_733,N_594);
or U3164 (N_3164,N_1668,N_2145);
nor U3165 (N_3165,N_591,N_2385);
xor U3166 (N_3166,N_1270,N_1000);
and U3167 (N_3167,N_1683,N_1238);
and U3168 (N_3168,N_2348,N_1855);
nand U3169 (N_3169,N_1493,N_1256);
nand U3170 (N_3170,N_66,N_821);
and U3171 (N_3171,N_1788,N_1637);
and U3172 (N_3172,N_2069,N_2216);
nor U3173 (N_3173,N_988,N_2171);
or U3174 (N_3174,N_581,N_318);
nand U3175 (N_3175,N_2123,N_1670);
and U3176 (N_3176,N_760,N_2129);
nor U3177 (N_3177,N_44,N_1361);
nand U3178 (N_3178,N_2246,N_1438);
and U3179 (N_3179,N_2085,N_2033);
xnor U3180 (N_3180,N_641,N_1130);
nand U3181 (N_3181,N_435,N_1841);
and U3182 (N_3182,N_800,N_908);
and U3183 (N_3183,N_41,N_658);
and U3184 (N_3184,N_997,N_2047);
nand U3185 (N_3185,N_340,N_332);
or U3186 (N_3186,N_180,N_1085);
nand U3187 (N_3187,N_2087,N_1038);
or U3188 (N_3188,N_1808,N_393);
or U3189 (N_3189,N_94,N_2121);
nand U3190 (N_3190,N_379,N_71);
or U3191 (N_3191,N_1404,N_493);
nand U3192 (N_3192,N_1946,N_401);
or U3193 (N_3193,N_768,N_217);
nand U3194 (N_3194,N_1572,N_2064);
nand U3195 (N_3195,N_1489,N_1564);
or U3196 (N_3196,N_653,N_784);
and U3197 (N_3197,N_618,N_2125);
nand U3198 (N_3198,N_331,N_1113);
and U3199 (N_3199,N_2167,N_74);
nand U3200 (N_3200,N_1900,N_1134);
nor U3201 (N_3201,N_90,N_500);
and U3202 (N_3202,N_1965,N_170);
and U3203 (N_3203,N_1262,N_2245);
or U3204 (N_3204,N_1541,N_806);
nor U3205 (N_3205,N_1293,N_662);
and U3206 (N_3206,N_1402,N_1364);
nor U3207 (N_3207,N_1666,N_2428);
or U3208 (N_3208,N_27,N_2157);
xnor U3209 (N_3209,N_1731,N_598);
or U3210 (N_3210,N_864,N_630);
and U3211 (N_3211,N_1599,N_1296);
or U3212 (N_3212,N_526,N_83);
or U3213 (N_3213,N_671,N_885);
nand U3214 (N_3214,N_676,N_636);
nand U3215 (N_3215,N_710,N_1694);
or U3216 (N_3216,N_1518,N_192);
and U3217 (N_3217,N_184,N_1274);
nand U3218 (N_3218,N_755,N_2432);
nand U3219 (N_3219,N_1691,N_678);
or U3220 (N_3220,N_1495,N_1761);
nand U3221 (N_3221,N_1359,N_405);
and U3222 (N_3222,N_2137,N_249);
nand U3223 (N_3223,N_926,N_244);
nor U3224 (N_3224,N_2402,N_2465);
and U3225 (N_3225,N_879,N_905);
nor U3226 (N_3226,N_2151,N_22);
xnor U3227 (N_3227,N_1395,N_1338);
nor U3228 (N_3228,N_88,N_214);
nand U3229 (N_3229,N_2460,N_932);
nor U3230 (N_3230,N_543,N_2390);
and U3231 (N_3231,N_722,N_726);
nor U3232 (N_3232,N_1229,N_2200);
nor U3233 (N_3233,N_918,N_53);
and U3234 (N_3234,N_850,N_59);
or U3235 (N_3235,N_449,N_522);
and U3236 (N_3236,N_1869,N_582);
or U3237 (N_3237,N_1425,N_523);
or U3238 (N_3238,N_1163,N_376);
nor U3239 (N_3239,N_1076,N_538);
and U3240 (N_3240,N_52,N_837);
and U3241 (N_3241,N_2010,N_914);
or U3242 (N_3242,N_504,N_2404);
nor U3243 (N_3243,N_872,N_2492);
and U3244 (N_3244,N_1697,N_1080);
nand U3245 (N_3245,N_1560,N_527);
or U3246 (N_3246,N_1651,N_1578);
or U3247 (N_3247,N_2162,N_2232);
or U3248 (N_3248,N_1070,N_106);
nor U3249 (N_3249,N_842,N_633);
and U3250 (N_3250,N_739,N_1819);
nand U3251 (N_3251,N_635,N_0);
or U3252 (N_3252,N_571,N_468);
nor U3253 (N_3253,N_1397,N_275);
xor U3254 (N_3254,N_1967,N_2146);
or U3255 (N_3255,N_646,N_714);
and U3256 (N_3256,N_1860,N_2494);
and U3257 (N_3257,N_2228,N_2448);
or U3258 (N_3258,N_631,N_1529);
and U3259 (N_3259,N_2456,N_2461);
nand U3260 (N_3260,N_1133,N_222);
nand U3261 (N_3261,N_1029,N_164);
and U3262 (N_3262,N_848,N_2044);
nor U3263 (N_3263,N_469,N_34);
nand U3264 (N_3264,N_1940,N_2051);
nor U3265 (N_3265,N_45,N_1007);
nand U3266 (N_3266,N_1313,N_967);
and U3267 (N_3267,N_715,N_1889);
nor U3268 (N_3268,N_746,N_890);
or U3269 (N_3269,N_1771,N_2175);
xnor U3270 (N_3270,N_1197,N_2442);
nor U3271 (N_3271,N_2447,N_1829);
nand U3272 (N_3272,N_1994,N_1275);
and U3273 (N_3273,N_452,N_84);
nand U3274 (N_3274,N_365,N_178);
or U3275 (N_3275,N_347,N_993);
or U3276 (N_3276,N_1903,N_426);
and U3277 (N_3277,N_407,N_246);
and U3278 (N_3278,N_2417,N_1824);
or U3279 (N_3279,N_2138,N_1144);
nor U3280 (N_3280,N_1465,N_1803);
nor U3281 (N_3281,N_1111,N_2437);
xnor U3282 (N_3282,N_1961,N_1765);
or U3283 (N_3283,N_303,N_1221);
or U3284 (N_3284,N_956,N_2223);
nor U3285 (N_3285,N_1766,N_2224);
or U3286 (N_3286,N_1491,N_51);
and U3287 (N_3287,N_1630,N_2235);
and U3288 (N_3288,N_251,N_274);
nor U3289 (N_3289,N_937,N_2271);
nand U3290 (N_3290,N_392,N_1278);
nor U3291 (N_3291,N_1216,N_549);
or U3292 (N_3292,N_2131,N_123);
nor U3293 (N_3293,N_1180,N_2387);
and U3294 (N_3294,N_627,N_1642);
or U3295 (N_3295,N_2111,N_1528);
nand U3296 (N_3296,N_751,N_301);
or U3297 (N_3297,N_971,N_670);
or U3298 (N_3298,N_1566,N_1349);
nand U3299 (N_3299,N_2066,N_1624);
and U3300 (N_3300,N_1003,N_354);
and U3301 (N_3301,N_2293,N_680);
or U3302 (N_3302,N_2280,N_2054);
and U3303 (N_3303,N_2366,N_688);
or U3304 (N_3304,N_1094,N_1053);
nand U3305 (N_3305,N_2317,N_2430);
nand U3306 (N_3306,N_1879,N_1243);
nand U3307 (N_3307,N_1605,N_1017);
nand U3308 (N_3308,N_2422,N_1934);
nor U3309 (N_3309,N_1958,N_2395);
or U3310 (N_3310,N_308,N_288);
nor U3311 (N_3311,N_1909,N_858);
xor U3312 (N_3312,N_659,N_212);
and U3313 (N_3313,N_498,N_778);
nand U3314 (N_3314,N_2306,N_1776);
nor U3315 (N_3315,N_40,N_1760);
nand U3316 (N_3316,N_728,N_1600);
or U3317 (N_3317,N_1342,N_798);
nand U3318 (N_3318,N_2208,N_165);
nand U3319 (N_3319,N_991,N_2248);
xor U3320 (N_3320,N_1155,N_1774);
nor U3321 (N_3321,N_2356,N_756);
or U3322 (N_3322,N_1417,N_362);
and U3323 (N_3323,N_1904,N_1055);
or U3324 (N_3324,N_1784,N_826);
and U3325 (N_3325,N_766,N_613);
nand U3326 (N_3326,N_211,N_2450);
and U3327 (N_3327,N_540,N_136);
and U3328 (N_3328,N_1537,N_1423);
and U3329 (N_3329,N_1805,N_2046);
or U3330 (N_3330,N_1318,N_3);
nor U3331 (N_3331,N_381,N_366);
nor U3332 (N_3332,N_1336,N_1279);
and U3333 (N_3333,N_2254,N_2242);
or U3334 (N_3334,N_2238,N_509);
and U3335 (N_3335,N_1553,N_982);
or U3336 (N_3336,N_1375,N_1736);
and U3337 (N_3337,N_2296,N_1527);
and U3338 (N_3338,N_1880,N_695);
nor U3339 (N_3339,N_725,N_1822);
or U3340 (N_3340,N_645,N_418);
nor U3341 (N_3341,N_1910,N_2031);
or U3342 (N_3342,N_919,N_1426);
or U3343 (N_3343,N_922,N_2336);
and U3344 (N_3344,N_1023,N_1343);
xor U3345 (N_3345,N_555,N_2112);
nand U3346 (N_3346,N_1059,N_1854);
nor U3347 (N_3347,N_2287,N_1725);
nand U3348 (N_3348,N_881,N_1297);
nor U3349 (N_3349,N_495,N_1459);
or U3350 (N_3350,N_141,N_2400);
nor U3351 (N_3351,N_2251,N_102);
and U3352 (N_3352,N_1982,N_371);
or U3353 (N_3353,N_1108,N_528);
and U3354 (N_3354,N_875,N_2166);
nor U3355 (N_3355,N_116,N_1409);
nand U3356 (N_3356,N_2474,N_1058);
nand U3357 (N_3357,N_82,N_2328);
or U3358 (N_3358,N_2333,N_674);
or U3359 (N_3359,N_1401,N_1341);
nor U3360 (N_3360,N_2090,N_604);
nor U3361 (N_3361,N_835,N_295);
and U3362 (N_3362,N_455,N_2250);
and U3363 (N_3363,N_802,N_1018);
nor U3364 (N_3364,N_281,N_1586);
and U3365 (N_3365,N_156,N_414);
or U3366 (N_3366,N_1178,N_1700);
nand U3367 (N_3367,N_2497,N_735);
nor U3368 (N_3368,N_1123,N_1611);
nor U3369 (N_3369,N_1258,N_1195);
or U3370 (N_3370,N_501,N_938);
nand U3371 (N_3371,N_951,N_1932);
nor U3372 (N_3372,N_2389,N_852);
or U3373 (N_3373,N_2160,N_1969);
nor U3374 (N_3374,N_2491,N_2213);
or U3375 (N_3375,N_968,N_896);
nand U3376 (N_3376,N_533,N_1056);
nor U3377 (N_3377,N_38,N_884);
nand U3378 (N_3378,N_510,N_2341);
nor U3379 (N_3379,N_1836,N_570);
and U3380 (N_3380,N_18,N_1914);
and U3381 (N_3381,N_737,N_554);
and U3382 (N_3382,N_1588,N_913);
and U3383 (N_3383,N_2332,N_1323);
nor U3384 (N_3384,N_2082,N_593);
and U3385 (N_3385,N_297,N_978);
nor U3386 (N_3386,N_1901,N_2368);
and U3387 (N_3387,N_2384,N_2017);
nand U3388 (N_3388,N_1612,N_2168);
nor U3389 (N_3389,N_1378,N_336);
and U3390 (N_3390,N_183,N_1686);
nor U3391 (N_3391,N_2397,N_557);
and U3392 (N_3392,N_2282,N_2239);
xor U3393 (N_3393,N_531,N_702);
nor U3394 (N_3394,N_1892,N_974);
nor U3395 (N_3395,N_1962,N_1674);
nor U3396 (N_3396,N_263,N_95);
nand U3397 (N_3397,N_2134,N_1255);
or U3398 (N_3398,N_1905,N_1750);
and U3399 (N_3399,N_1792,N_1591);
nand U3400 (N_3400,N_2380,N_1015);
and U3401 (N_3401,N_12,N_1800);
nand U3402 (N_3402,N_2142,N_2297);
nand U3403 (N_3403,N_49,N_1511);
or U3404 (N_3404,N_2144,N_1027);
nand U3405 (N_3405,N_1156,N_390);
or U3406 (N_3406,N_2266,N_120);
or U3407 (N_3407,N_1531,N_1603);
and U3408 (N_3408,N_958,N_514);
nor U3409 (N_3409,N_2496,N_1580);
nand U3410 (N_3410,N_572,N_2002);
nand U3411 (N_3411,N_1254,N_221);
nor U3412 (N_3412,N_475,N_1648);
or U3413 (N_3413,N_2262,N_2483);
and U3414 (N_3414,N_2027,N_1734);
nor U3415 (N_3415,N_970,N_587);
nand U3416 (N_3416,N_605,N_2359);
or U3417 (N_3417,N_644,N_547);
or U3418 (N_3418,N_753,N_712);
nand U3419 (N_3419,N_1781,N_1867);
and U3420 (N_3420,N_1823,N_747);
nand U3421 (N_3421,N_139,N_873);
nor U3422 (N_3422,N_882,N_290);
nor U3423 (N_3423,N_1748,N_2036);
or U3424 (N_3424,N_623,N_2489);
nor U3425 (N_3425,N_2458,N_2219);
nor U3426 (N_3426,N_961,N_1844);
or U3427 (N_3427,N_1002,N_176);
nor U3428 (N_3428,N_1380,N_310);
nand U3429 (N_3429,N_2045,N_396);
or U3430 (N_3430,N_664,N_1916);
nand U3431 (N_3431,N_2102,N_300);
and U3432 (N_3432,N_1864,N_1849);
nand U3433 (N_3433,N_2462,N_1486);
or U3434 (N_3434,N_447,N_1778);
nand U3435 (N_3435,N_1693,N_1035);
or U3436 (N_3436,N_764,N_146);
nor U3437 (N_3437,N_1764,N_360);
xor U3438 (N_3438,N_480,N_1607);
nand U3439 (N_3439,N_2118,N_473);
or U3440 (N_3440,N_2103,N_2011);
and U3441 (N_3441,N_175,N_86);
nand U3442 (N_3442,N_2156,N_1276);
and U3443 (N_3443,N_36,N_2070);
and U3444 (N_3444,N_965,N_1815);
or U3445 (N_3445,N_1675,N_2188);
and U3446 (N_3446,N_2386,N_780);
nand U3447 (N_3447,N_307,N_1277);
or U3448 (N_3448,N_1832,N_2019);
nand U3449 (N_3449,N_1986,N_1796);
and U3450 (N_3450,N_152,N_2078);
or U3451 (N_3451,N_1831,N_1821);
or U3452 (N_3452,N_1706,N_256);
nand U3453 (N_3453,N_992,N_694);
nor U3454 (N_3454,N_1171,N_7);
nand U3455 (N_3455,N_2312,N_1669);
nand U3456 (N_3456,N_1935,N_625);
and U3457 (N_3457,N_2265,N_1042);
and U3458 (N_3458,N_2068,N_2288);
or U3459 (N_3459,N_1633,N_296);
nand U3460 (N_3460,N_252,N_100);
nand U3461 (N_3461,N_2039,N_2021);
nand U3462 (N_3462,N_1019,N_1315);
nor U3463 (N_3463,N_2314,N_788);
nand U3464 (N_3464,N_1060,N_323);
or U3465 (N_3465,N_1520,N_280);
nand U3466 (N_3466,N_1230,N_1852);
nor U3467 (N_3467,N_266,N_1999);
and U3468 (N_3468,N_60,N_1711);
and U3469 (N_3469,N_2148,N_1845);
nand U3470 (N_3470,N_624,N_486);
or U3471 (N_3471,N_1658,N_989);
nand U3472 (N_3472,N_776,N_1356);
or U3473 (N_3473,N_1692,N_824);
and U3474 (N_3474,N_599,N_1032);
or U3475 (N_3475,N_1159,N_1938);
and U3476 (N_3476,N_1025,N_2407);
and U3477 (N_3477,N_804,N_1933);
or U3478 (N_3478,N_2055,N_2466);
nand U3479 (N_3479,N_942,N_1129);
nand U3480 (N_3480,N_1753,N_302);
or U3481 (N_3481,N_1242,N_43);
and U3482 (N_3482,N_2269,N_1557);
and U3483 (N_3483,N_1853,N_487);
nand U3484 (N_3484,N_2,N_324);
and U3485 (N_3485,N_319,N_1547);
nand U3486 (N_3486,N_1863,N_2425);
nor U3487 (N_3487,N_58,N_1010);
and U3488 (N_3488,N_2478,N_1064);
nand U3489 (N_3489,N_1558,N_185);
nand U3490 (N_3490,N_698,N_1310);
and U3491 (N_3491,N_878,N_2319);
nand U3492 (N_3492,N_172,N_1593);
nand U3493 (N_3493,N_891,N_1104);
nand U3494 (N_3494,N_1008,N_1636);
and U3495 (N_3495,N_1416,N_293);
nand U3496 (N_3496,N_2259,N_237);
or U3497 (N_3497,N_1487,N_1203);
nand U3498 (N_3498,N_1097,N_1253);
nor U3499 (N_3499,N_1638,N_2210);
and U3500 (N_3500,N_1016,N_556);
or U3501 (N_3501,N_1616,N_1639);
nand U3502 (N_3502,N_1679,N_1850);
and U3503 (N_3503,N_1039,N_320);
and U3504 (N_3504,N_262,N_1213);
nor U3505 (N_3505,N_661,N_793);
nand U3506 (N_3506,N_1559,N_464);
nand U3507 (N_3507,N_1478,N_179);
nor U3508 (N_3508,N_2339,N_488);
nor U3509 (N_3509,N_2204,N_1567);
nand U3510 (N_3510,N_1219,N_276);
and U3511 (N_3511,N_1833,N_844);
or U3512 (N_3512,N_1348,N_1052);
and U3513 (N_3513,N_1154,N_2405);
or U3514 (N_3514,N_1835,N_1065);
or U3515 (N_3515,N_1062,N_1856);
and U3516 (N_3516,N_1226,N_506);
nand U3517 (N_3517,N_1606,N_2139);
and U3518 (N_3518,N_1410,N_562);
or U3519 (N_3519,N_669,N_2467);
and U3520 (N_3520,N_201,N_1947);
nor U3521 (N_3521,N_2372,N_542);
and U3522 (N_3522,N_1877,N_1601);
nand U3523 (N_3523,N_1307,N_11);
and U3524 (N_3524,N_1467,N_1921);
or U3525 (N_3525,N_1372,N_1071);
and U3526 (N_3526,N_1181,N_1872);
nand U3527 (N_3527,N_482,N_413);
nor U3528 (N_3528,N_611,N_1763);
and U3529 (N_3529,N_1755,N_260);
nand U3530 (N_3530,N_484,N_1431);
nand U3531 (N_3531,N_440,N_2334);
or U3532 (N_3532,N_2165,N_2198);
nor U3533 (N_3533,N_1826,N_1615);
nand U3534 (N_3534,N_2179,N_1369);
and U3535 (N_3535,N_2205,N_812);
xor U3536 (N_3536,N_1360,N_1868);
or U3537 (N_3537,N_233,N_1399);
and U3538 (N_3538,N_740,N_2048);
nor U3539 (N_3539,N_441,N_1479);
nand U3540 (N_3540,N_1470,N_245);
and U3541 (N_3541,N_388,N_1769);
nand U3542 (N_3542,N_667,N_1330);
or U3543 (N_3543,N_2362,N_1092);
nor U3544 (N_3544,N_343,N_1696);
nor U3545 (N_3545,N_563,N_1340);
nor U3546 (N_3546,N_306,N_541);
or U3547 (N_3547,N_1626,N_823);
and U3548 (N_3548,N_67,N_1143);
and U3549 (N_3549,N_1746,N_412);
xor U3550 (N_3550,N_330,N_1780);
nand U3551 (N_3551,N_1507,N_1354);
nand U3552 (N_3552,N_1138,N_552);
nor U3553 (N_3553,N_608,N_2381);
and U3554 (N_3554,N_2298,N_474);
and U3555 (N_3555,N_128,N_1331);
or U3556 (N_3556,N_1704,N_28);
or U3557 (N_3557,N_931,N_200);
or U3558 (N_3558,N_1463,N_363);
or U3559 (N_3559,N_1811,N_1200);
or U3560 (N_3560,N_1506,N_1917);
nand U3561 (N_3561,N_1311,N_148);
or U3562 (N_3562,N_1471,N_813);
or U3563 (N_3563,N_1785,N_2283);
nor U3564 (N_3564,N_825,N_2369);
or U3565 (N_3565,N_1101,N_576);
nand U3566 (N_3566,N_2394,N_1840);
nand U3567 (N_3567,N_2100,N_1199);
or U3568 (N_3568,N_1362,N_472);
nand U3569 (N_3569,N_1985,N_1906);
nor U3570 (N_3570,N_16,N_2406);
nand U3571 (N_3571,N_759,N_1810);
nor U3572 (N_3572,N_1568,N_889);
or U3573 (N_3573,N_1445,N_1096);
nor U3574 (N_3574,N_2233,N_2487);
nand U3575 (N_3575,N_240,N_335);
nand U3576 (N_3576,N_1265,N_1715);
nand U3577 (N_3577,N_834,N_700);
and U3578 (N_3578,N_272,N_417);
and U3579 (N_3579,N_731,N_2304);
nand U3580 (N_3580,N_77,N_2308);
nand U3581 (N_3581,N_814,N_1444);
nor U3582 (N_3582,N_2424,N_230);
nor U3583 (N_3583,N_68,N_2101);
xor U3584 (N_3584,N_241,N_1942);
nor U3585 (N_3585,N_1225,N_333);
or U3586 (N_3586,N_1034,N_257);
nand U3587 (N_3587,N_1294,N_1333);
nor U3588 (N_3588,N_436,N_1660);
xnor U3589 (N_3589,N_1920,N_46);
or U3590 (N_3590,N_2043,N_190);
nand U3591 (N_3591,N_1405,N_1848);
nor U3592 (N_3592,N_2007,N_1049);
or U3593 (N_3593,N_1109,N_2411);
nand U3594 (N_3594,N_118,N_1030);
and U3595 (N_3595,N_1978,N_2071);
nor U3596 (N_3596,N_1928,N_1662);
nand U3597 (N_3597,N_1115,N_1435);
nand U3598 (N_3598,N_1723,N_2279);
nand U3599 (N_3599,N_1345,N_921);
nand U3600 (N_3600,N_191,N_264);
nand U3601 (N_3601,N_1550,N_1411);
nor U3602 (N_3602,N_1050,N_348);
and U3603 (N_3603,N_772,N_1128);
or U3604 (N_3604,N_856,N_933);
and U3605 (N_3605,N_1598,N_1437);
nand U3606 (N_3606,N_1088,N_2459);
and U3607 (N_3607,N_1468,N_87);
nand U3608 (N_3608,N_2143,N_1304);
or U3609 (N_3609,N_353,N_63);
or U3610 (N_3610,N_1248,N_2309);
and U3611 (N_3611,N_1400,N_104);
nand U3612 (N_3612,N_634,N_1927);
and U3613 (N_3613,N_1751,N_2305);
or U3614 (N_3614,N_1818,N_1048);
and U3615 (N_3615,N_827,N_283);
and U3616 (N_3616,N_1794,N_25);
nand U3617 (N_3617,N_2192,N_1232);
nor U3618 (N_3618,N_1217,N_1698);
nand U3619 (N_3619,N_900,N_2207);
and U3620 (N_3620,N_1665,N_1418);
nor U3621 (N_3621,N_239,N_2120);
or U3622 (N_3622,N_941,N_1081);
and U3623 (N_3623,N_2196,N_2331);
and U3624 (N_3624,N_592,N_1618);
nor U3625 (N_3625,N_983,N_2081);
or U3626 (N_3626,N_818,N_1325);
or U3627 (N_3627,N_1451,N_1828);
or U3628 (N_3628,N_489,N_705);
nand U3629 (N_3629,N_910,N_2345);
or U3630 (N_3630,N_2471,N_1887);
or U3631 (N_3631,N_1843,N_316);
nand U3632 (N_3632,N_789,N_2403);
or U3633 (N_3633,N_2141,N_1406);
or U3634 (N_3634,N_1093,N_2302);
xor U3635 (N_3635,N_893,N_1516);
or U3636 (N_3636,N_1091,N_1970);
and U3637 (N_3637,N_1862,N_1574);
and U3638 (N_3638,N_2480,N_352);
nand U3639 (N_3639,N_1245,N_1992);
nor U3640 (N_3640,N_590,N_1456);
and U3641 (N_3641,N_1595,N_2058);
nor U3642 (N_3642,N_1939,N_717);
or U3643 (N_3643,N_2097,N_1710);
nand U3644 (N_3644,N_2001,N_2086);
nand U3645 (N_3645,N_1099,N_517);
nand U3646 (N_3646,N_2187,N_2072);
nor U3647 (N_3647,N_1407,N_157);
or U3648 (N_3648,N_999,N_2214);
xnor U3649 (N_3649,N_1102,N_773);
nand U3650 (N_3650,N_2091,N_479);
nand U3651 (N_3651,N_1415,N_1689);
nand U3652 (N_3652,N_50,N_639);
nand U3653 (N_3653,N_4,N_521);
nand U3654 (N_3654,N_619,N_1069);
or U3655 (N_3655,N_1269,N_2020);
nor U3656 (N_3656,N_578,N_1384);
nor U3657 (N_3657,N_2041,N_5);
and U3658 (N_3658,N_943,N_1095);
and U3659 (N_3659,N_54,N_423);
nand U3660 (N_3660,N_1188,N_1208);
nor U3661 (N_3661,N_803,N_1078);
nand U3662 (N_3662,N_1244,N_2276);
and U3663 (N_3663,N_109,N_1327);
nand U3664 (N_3664,N_1678,N_1775);
or U3665 (N_3665,N_762,N_955);
and U3666 (N_3666,N_1026,N_1215);
or U3667 (N_3667,N_707,N_1272);
nor U3668 (N_3668,N_550,N_871);
and U3669 (N_3669,N_1820,N_2477);
or U3670 (N_3670,N_650,N_508);
or U3671 (N_3671,N_887,N_1919);
and U3672 (N_3672,N_833,N_470);
or U3673 (N_3673,N_1538,N_159);
and U3674 (N_3674,N_2256,N_1536);
nand U3675 (N_3675,N_2363,N_2409);
or U3676 (N_3676,N_1383,N_1551);
and U3677 (N_3677,N_466,N_400);
nand U3678 (N_3678,N_356,N_2301);
nor U3679 (N_3679,N_843,N_1284);
nor U3680 (N_3680,N_923,N_269);
or U3681 (N_3681,N_225,N_1044);
and U3682 (N_3682,N_811,N_537);
xor U3683 (N_3683,N_920,N_1847);
nor U3684 (N_3684,N_1545,N_2294);
and U3685 (N_3685,N_2030,N_865);
or U3686 (N_3686,N_779,N_742);
and U3687 (N_3687,N_2032,N_2286);
nand U3688 (N_3688,N_55,N_1745);
or U3689 (N_3689,N_1953,N_1922);
and U3690 (N_3690,N_1937,N_2436);
nor U3691 (N_3691,N_2215,N_1663);
nor U3692 (N_3692,N_718,N_596);
and U3693 (N_3693,N_26,N_1622);
nor U3694 (N_3694,N_182,N_2488);
or U3695 (N_3695,N_1367,N_385);
and U3696 (N_3696,N_839,N_1132);
nand U3697 (N_3697,N_497,N_1377);
or U3698 (N_3698,N_1830,N_1398);
or U3699 (N_3699,N_2023,N_1749);
nand U3700 (N_3700,N_2053,N_1677);
and U3701 (N_3701,N_1702,N_1767);
or U3702 (N_3702,N_859,N_1347);
nor U3703 (N_3703,N_716,N_1653);
and U3704 (N_3704,N_668,N_1235);
or U3705 (N_3705,N_1782,N_2206);
nand U3706 (N_3706,N_719,N_2018);
or U3707 (N_3707,N_524,N_597);
and U3708 (N_3708,N_329,N_2170);
and U3709 (N_3709,N_1458,N_1391);
xor U3710 (N_3710,N_980,N_1540);
nor U3711 (N_3711,N_1057,N_1980);
or U3712 (N_3712,N_948,N_1634);
or U3713 (N_3713,N_1728,N_907);
and U3714 (N_3714,N_1716,N_2484);
or U3715 (N_3715,N_2063,N_924);
or U3716 (N_3716,N_2094,N_2329);
nor U3717 (N_3717,N_131,N_1192);
nor U3718 (N_3718,N_1166,N_791);
and U3719 (N_3719,N_1453,N_103);
and U3720 (N_3720,N_2300,N_1298);
nor U3721 (N_3721,N_640,N_911);
and U3722 (N_3722,N_259,N_763);
nor U3723 (N_3723,N_2335,N_1851);
nor U3724 (N_3724,N_1726,N_91);
or U3725 (N_3725,N_2473,N_1328);
nor U3726 (N_3726,N_124,N_304);
nor U3727 (N_3727,N_2155,N_1839);
and U3728 (N_3728,N_1931,N_1214);
or U3729 (N_3729,N_1802,N_21);
nand U3730 (N_3730,N_2446,N_1237);
or U3731 (N_3731,N_1082,N_33);
nor U3732 (N_3732,N_450,N_1472);
nand U3733 (N_3733,N_732,N_2311);
nor U3734 (N_3734,N_2237,N_1412);
and U3735 (N_3735,N_1878,N_2439);
nor U3736 (N_3736,N_2061,N_315);
or U3737 (N_3737,N_1474,N_1738);
and U3738 (N_3738,N_985,N_325);
nand U3739 (N_3739,N_1729,N_1514);
nand U3740 (N_3740,N_1394,N_2340);
nand U3741 (N_3741,N_1876,N_899);
nor U3742 (N_3742,N_1955,N_1107);
nor U3743 (N_3743,N_1009,N_2159);
nor U3744 (N_3744,N_278,N_1659);
and U3745 (N_3745,N_2104,N_291);
and U3746 (N_3746,N_1894,N_344);
and U3747 (N_3747,N_2371,N_516);
or U3748 (N_3748,N_1320,N_1963);
nand U3749 (N_3749,N_358,N_1526);
nand U3750 (N_3750,N_1302,N_561);
nand U3751 (N_3751,N_1641,N_26);
nand U3752 (N_3752,N_1339,N_320);
nand U3753 (N_3753,N_749,N_1143);
nand U3754 (N_3754,N_749,N_154);
or U3755 (N_3755,N_2233,N_1449);
and U3756 (N_3756,N_2456,N_1506);
nand U3757 (N_3757,N_2100,N_1190);
nor U3758 (N_3758,N_934,N_1114);
nand U3759 (N_3759,N_1727,N_2053);
nand U3760 (N_3760,N_1944,N_1873);
nand U3761 (N_3761,N_1179,N_1194);
nor U3762 (N_3762,N_1490,N_854);
and U3763 (N_3763,N_2129,N_54);
and U3764 (N_3764,N_1368,N_179);
nand U3765 (N_3765,N_84,N_1383);
and U3766 (N_3766,N_1791,N_1696);
and U3767 (N_3767,N_1285,N_1570);
or U3768 (N_3768,N_2008,N_1983);
nor U3769 (N_3769,N_2209,N_929);
and U3770 (N_3770,N_1934,N_987);
nand U3771 (N_3771,N_1582,N_1618);
or U3772 (N_3772,N_579,N_2098);
nor U3773 (N_3773,N_1811,N_1463);
and U3774 (N_3774,N_405,N_590);
nand U3775 (N_3775,N_532,N_154);
nor U3776 (N_3776,N_246,N_609);
and U3777 (N_3777,N_794,N_1286);
nor U3778 (N_3778,N_1239,N_1226);
nand U3779 (N_3779,N_812,N_1057);
or U3780 (N_3780,N_1918,N_1133);
nor U3781 (N_3781,N_1981,N_1282);
and U3782 (N_3782,N_262,N_264);
and U3783 (N_3783,N_1614,N_371);
or U3784 (N_3784,N_1925,N_601);
or U3785 (N_3785,N_1412,N_625);
or U3786 (N_3786,N_2089,N_857);
or U3787 (N_3787,N_1030,N_1566);
or U3788 (N_3788,N_1434,N_1417);
and U3789 (N_3789,N_470,N_784);
nor U3790 (N_3790,N_274,N_113);
and U3791 (N_3791,N_167,N_88);
or U3792 (N_3792,N_2059,N_578);
nor U3793 (N_3793,N_736,N_574);
or U3794 (N_3794,N_1415,N_1260);
nor U3795 (N_3795,N_2452,N_1612);
or U3796 (N_3796,N_290,N_348);
nor U3797 (N_3797,N_1025,N_684);
or U3798 (N_3798,N_1560,N_889);
nor U3799 (N_3799,N_1403,N_2365);
nor U3800 (N_3800,N_1440,N_1070);
and U3801 (N_3801,N_1701,N_758);
nand U3802 (N_3802,N_705,N_1756);
and U3803 (N_3803,N_998,N_865);
nand U3804 (N_3804,N_1472,N_528);
and U3805 (N_3805,N_2264,N_1214);
nand U3806 (N_3806,N_905,N_1013);
and U3807 (N_3807,N_1414,N_2401);
nor U3808 (N_3808,N_2036,N_2444);
nor U3809 (N_3809,N_1859,N_1068);
or U3810 (N_3810,N_1495,N_1604);
and U3811 (N_3811,N_1041,N_929);
and U3812 (N_3812,N_1332,N_2204);
or U3813 (N_3813,N_675,N_1189);
and U3814 (N_3814,N_2439,N_278);
and U3815 (N_3815,N_726,N_961);
and U3816 (N_3816,N_1491,N_1039);
and U3817 (N_3817,N_2077,N_890);
nor U3818 (N_3818,N_975,N_209);
and U3819 (N_3819,N_2008,N_914);
nor U3820 (N_3820,N_403,N_244);
or U3821 (N_3821,N_2389,N_97);
nand U3822 (N_3822,N_1022,N_1881);
or U3823 (N_3823,N_2269,N_459);
nor U3824 (N_3824,N_311,N_2064);
nand U3825 (N_3825,N_1758,N_1662);
or U3826 (N_3826,N_1454,N_1424);
nand U3827 (N_3827,N_554,N_12);
and U3828 (N_3828,N_2170,N_1072);
nor U3829 (N_3829,N_1408,N_1035);
nand U3830 (N_3830,N_1747,N_6);
or U3831 (N_3831,N_1895,N_424);
or U3832 (N_3832,N_453,N_302);
nor U3833 (N_3833,N_1215,N_851);
and U3834 (N_3834,N_1230,N_190);
nor U3835 (N_3835,N_927,N_1075);
and U3836 (N_3836,N_209,N_966);
nand U3837 (N_3837,N_1247,N_2289);
or U3838 (N_3838,N_128,N_1902);
or U3839 (N_3839,N_799,N_1971);
or U3840 (N_3840,N_2165,N_911);
xnor U3841 (N_3841,N_722,N_2228);
xnor U3842 (N_3842,N_2024,N_1990);
or U3843 (N_3843,N_2069,N_790);
nor U3844 (N_3844,N_1484,N_2271);
nand U3845 (N_3845,N_646,N_433);
or U3846 (N_3846,N_1308,N_2066);
nand U3847 (N_3847,N_2284,N_586);
xor U3848 (N_3848,N_2294,N_1445);
or U3849 (N_3849,N_1352,N_2293);
or U3850 (N_3850,N_619,N_2257);
and U3851 (N_3851,N_1582,N_1464);
and U3852 (N_3852,N_513,N_362);
xnor U3853 (N_3853,N_618,N_612);
or U3854 (N_3854,N_488,N_1695);
or U3855 (N_3855,N_592,N_1699);
nor U3856 (N_3856,N_853,N_1260);
nor U3857 (N_3857,N_1292,N_206);
nor U3858 (N_3858,N_679,N_118);
nor U3859 (N_3859,N_1428,N_978);
and U3860 (N_3860,N_1372,N_1734);
and U3861 (N_3861,N_2109,N_623);
xnor U3862 (N_3862,N_601,N_9);
nand U3863 (N_3863,N_2192,N_283);
nor U3864 (N_3864,N_1993,N_328);
nor U3865 (N_3865,N_131,N_575);
nand U3866 (N_3866,N_1578,N_152);
or U3867 (N_3867,N_1779,N_1214);
nand U3868 (N_3868,N_2126,N_50);
nor U3869 (N_3869,N_2315,N_1744);
nand U3870 (N_3870,N_1580,N_2448);
and U3871 (N_3871,N_571,N_277);
or U3872 (N_3872,N_101,N_1736);
nand U3873 (N_3873,N_645,N_1473);
nand U3874 (N_3874,N_76,N_345);
xnor U3875 (N_3875,N_409,N_1580);
nand U3876 (N_3876,N_1891,N_644);
nand U3877 (N_3877,N_559,N_1421);
nand U3878 (N_3878,N_2072,N_1277);
nand U3879 (N_3879,N_646,N_1661);
or U3880 (N_3880,N_383,N_1614);
nand U3881 (N_3881,N_505,N_1039);
nor U3882 (N_3882,N_2062,N_176);
nor U3883 (N_3883,N_679,N_777);
nor U3884 (N_3884,N_1134,N_1292);
and U3885 (N_3885,N_981,N_415);
nand U3886 (N_3886,N_2064,N_1975);
nand U3887 (N_3887,N_1229,N_355);
or U3888 (N_3888,N_995,N_1728);
nor U3889 (N_3889,N_441,N_1699);
and U3890 (N_3890,N_2355,N_1886);
xnor U3891 (N_3891,N_1554,N_436);
xnor U3892 (N_3892,N_1634,N_290);
nor U3893 (N_3893,N_655,N_379);
and U3894 (N_3894,N_2235,N_292);
or U3895 (N_3895,N_1587,N_694);
nand U3896 (N_3896,N_293,N_2113);
and U3897 (N_3897,N_1939,N_991);
and U3898 (N_3898,N_335,N_695);
and U3899 (N_3899,N_2224,N_699);
or U3900 (N_3900,N_1865,N_938);
and U3901 (N_3901,N_470,N_2378);
nand U3902 (N_3902,N_2129,N_701);
and U3903 (N_3903,N_615,N_1786);
or U3904 (N_3904,N_1442,N_1804);
or U3905 (N_3905,N_904,N_310);
nor U3906 (N_3906,N_1665,N_593);
xnor U3907 (N_3907,N_2117,N_603);
nand U3908 (N_3908,N_1222,N_417);
and U3909 (N_3909,N_2201,N_796);
nand U3910 (N_3910,N_1370,N_1915);
nor U3911 (N_3911,N_676,N_930);
and U3912 (N_3912,N_1841,N_427);
nor U3913 (N_3913,N_1132,N_733);
and U3914 (N_3914,N_1111,N_1289);
nor U3915 (N_3915,N_685,N_468);
nor U3916 (N_3916,N_122,N_862);
or U3917 (N_3917,N_1120,N_2442);
nor U3918 (N_3918,N_112,N_1660);
xnor U3919 (N_3919,N_2305,N_1009);
or U3920 (N_3920,N_1770,N_974);
or U3921 (N_3921,N_1220,N_1069);
nor U3922 (N_3922,N_2426,N_2405);
and U3923 (N_3923,N_2148,N_1801);
and U3924 (N_3924,N_2074,N_1670);
nand U3925 (N_3925,N_376,N_1123);
or U3926 (N_3926,N_2031,N_2254);
nor U3927 (N_3927,N_409,N_643);
or U3928 (N_3928,N_1997,N_1727);
or U3929 (N_3929,N_1434,N_235);
and U3930 (N_3930,N_1677,N_232);
nor U3931 (N_3931,N_1045,N_2287);
and U3932 (N_3932,N_609,N_1885);
or U3933 (N_3933,N_609,N_1926);
nor U3934 (N_3934,N_657,N_343);
and U3935 (N_3935,N_1533,N_502);
and U3936 (N_3936,N_151,N_1096);
and U3937 (N_3937,N_2497,N_407);
nand U3938 (N_3938,N_2292,N_484);
nor U3939 (N_3939,N_109,N_1043);
or U3940 (N_3940,N_1445,N_1529);
and U3941 (N_3941,N_988,N_2100);
and U3942 (N_3942,N_2074,N_437);
nor U3943 (N_3943,N_1204,N_1254);
nand U3944 (N_3944,N_1978,N_1077);
nand U3945 (N_3945,N_1903,N_343);
or U3946 (N_3946,N_305,N_1495);
nand U3947 (N_3947,N_930,N_213);
nor U3948 (N_3948,N_629,N_218);
nor U3949 (N_3949,N_1830,N_257);
nor U3950 (N_3950,N_1390,N_1147);
nor U3951 (N_3951,N_2200,N_2181);
or U3952 (N_3952,N_2387,N_874);
nor U3953 (N_3953,N_2056,N_12);
or U3954 (N_3954,N_891,N_1124);
xnor U3955 (N_3955,N_828,N_2388);
or U3956 (N_3956,N_1871,N_1530);
or U3957 (N_3957,N_504,N_700);
nand U3958 (N_3958,N_336,N_1590);
and U3959 (N_3959,N_2123,N_432);
and U3960 (N_3960,N_368,N_2403);
and U3961 (N_3961,N_801,N_1410);
nor U3962 (N_3962,N_34,N_916);
nor U3963 (N_3963,N_1054,N_921);
nand U3964 (N_3964,N_2014,N_1537);
nand U3965 (N_3965,N_2165,N_649);
and U3966 (N_3966,N_173,N_1656);
nor U3967 (N_3967,N_1067,N_1421);
nor U3968 (N_3968,N_2290,N_297);
nor U3969 (N_3969,N_1046,N_1937);
nand U3970 (N_3970,N_1970,N_1431);
and U3971 (N_3971,N_2458,N_535);
or U3972 (N_3972,N_749,N_2337);
nor U3973 (N_3973,N_98,N_2472);
nor U3974 (N_3974,N_91,N_1942);
nor U3975 (N_3975,N_2395,N_2272);
or U3976 (N_3976,N_133,N_2153);
nor U3977 (N_3977,N_1413,N_798);
or U3978 (N_3978,N_2303,N_747);
nor U3979 (N_3979,N_1891,N_820);
and U3980 (N_3980,N_1958,N_50);
nand U3981 (N_3981,N_32,N_1591);
or U3982 (N_3982,N_947,N_681);
or U3983 (N_3983,N_1864,N_1246);
nor U3984 (N_3984,N_2068,N_686);
and U3985 (N_3985,N_973,N_1101);
and U3986 (N_3986,N_868,N_198);
or U3987 (N_3987,N_0,N_2199);
and U3988 (N_3988,N_1239,N_554);
and U3989 (N_3989,N_277,N_1643);
xor U3990 (N_3990,N_1710,N_402);
or U3991 (N_3991,N_901,N_558);
nor U3992 (N_3992,N_1933,N_322);
nor U3993 (N_3993,N_335,N_432);
nor U3994 (N_3994,N_1552,N_1946);
nand U3995 (N_3995,N_310,N_1456);
nand U3996 (N_3996,N_2154,N_311);
nor U3997 (N_3997,N_1846,N_1624);
or U3998 (N_3998,N_1506,N_1028);
or U3999 (N_3999,N_684,N_1564);
nand U4000 (N_4000,N_576,N_1676);
nand U4001 (N_4001,N_842,N_2193);
and U4002 (N_4002,N_1592,N_1894);
and U4003 (N_4003,N_740,N_64);
nand U4004 (N_4004,N_454,N_1093);
or U4005 (N_4005,N_914,N_2475);
nand U4006 (N_4006,N_1214,N_730);
and U4007 (N_4007,N_2205,N_473);
and U4008 (N_4008,N_2318,N_702);
nor U4009 (N_4009,N_1333,N_284);
and U4010 (N_4010,N_161,N_1185);
and U4011 (N_4011,N_1068,N_1474);
nand U4012 (N_4012,N_2196,N_1293);
nand U4013 (N_4013,N_2132,N_1911);
nor U4014 (N_4014,N_1588,N_699);
and U4015 (N_4015,N_835,N_135);
nor U4016 (N_4016,N_1700,N_346);
and U4017 (N_4017,N_1375,N_1080);
or U4018 (N_4018,N_2180,N_1138);
nor U4019 (N_4019,N_1689,N_2046);
or U4020 (N_4020,N_63,N_2394);
nand U4021 (N_4021,N_608,N_1046);
nor U4022 (N_4022,N_761,N_1017);
or U4023 (N_4023,N_951,N_1647);
nor U4024 (N_4024,N_967,N_905);
and U4025 (N_4025,N_311,N_2177);
nor U4026 (N_4026,N_344,N_1482);
or U4027 (N_4027,N_1544,N_2314);
nand U4028 (N_4028,N_1092,N_304);
or U4029 (N_4029,N_2000,N_625);
nand U4030 (N_4030,N_1789,N_2492);
nand U4031 (N_4031,N_2117,N_1406);
and U4032 (N_4032,N_1553,N_289);
nand U4033 (N_4033,N_1943,N_1185);
and U4034 (N_4034,N_2408,N_2026);
nor U4035 (N_4035,N_524,N_2428);
nor U4036 (N_4036,N_1798,N_371);
or U4037 (N_4037,N_640,N_1737);
xor U4038 (N_4038,N_1209,N_2020);
and U4039 (N_4039,N_2391,N_1874);
nand U4040 (N_4040,N_1448,N_1020);
and U4041 (N_4041,N_458,N_2184);
nor U4042 (N_4042,N_1419,N_298);
nand U4043 (N_4043,N_729,N_1360);
or U4044 (N_4044,N_1300,N_1525);
nor U4045 (N_4045,N_303,N_2356);
nand U4046 (N_4046,N_1392,N_1021);
nand U4047 (N_4047,N_1136,N_882);
or U4048 (N_4048,N_1278,N_2290);
or U4049 (N_4049,N_657,N_1569);
and U4050 (N_4050,N_369,N_1739);
or U4051 (N_4051,N_1770,N_261);
or U4052 (N_4052,N_1660,N_1779);
and U4053 (N_4053,N_2162,N_840);
and U4054 (N_4054,N_61,N_208);
and U4055 (N_4055,N_2422,N_1393);
nand U4056 (N_4056,N_1323,N_1003);
or U4057 (N_4057,N_1872,N_604);
and U4058 (N_4058,N_395,N_1441);
and U4059 (N_4059,N_2462,N_1948);
nand U4060 (N_4060,N_1240,N_676);
nand U4061 (N_4061,N_503,N_1693);
xnor U4062 (N_4062,N_1469,N_406);
and U4063 (N_4063,N_1331,N_668);
nor U4064 (N_4064,N_2387,N_682);
nand U4065 (N_4065,N_2043,N_887);
or U4066 (N_4066,N_2143,N_337);
or U4067 (N_4067,N_1713,N_33);
nand U4068 (N_4068,N_1672,N_2422);
nor U4069 (N_4069,N_1218,N_1386);
or U4070 (N_4070,N_1247,N_655);
and U4071 (N_4071,N_1923,N_555);
and U4072 (N_4072,N_746,N_2244);
and U4073 (N_4073,N_639,N_2124);
nor U4074 (N_4074,N_392,N_326);
and U4075 (N_4075,N_1674,N_981);
and U4076 (N_4076,N_147,N_613);
xor U4077 (N_4077,N_1813,N_570);
nand U4078 (N_4078,N_407,N_669);
nand U4079 (N_4079,N_509,N_2464);
or U4080 (N_4080,N_2132,N_1138);
nor U4081 (N_4081,N_1680,N_1978);
nor U4082 (N_4082,N_61,N_322);
or U4083 (N_4083,N_1461,N_252);
nor U4084 (N_4084,N_1350,N_71);
or U4085 (N_4085,N_2475,N_499);
or U4086 (N_4086,N_412,N_1489);
nor U4087 (N_4087,N_885,N_1541);
and U4088 (N_4088,N_1484,N_11);
nor U4089 (N_4089,N_2307,N_2110);
nand U4090 (N_4090,N_475,N_773);
nor U4091 (N_4091,N_2451,N_127);
and U4092 (N_4092,N_715,N_2063);
nor U4093 (N_4093,N_974,N_1957);
nand U4094 (N_4094,N_1188,N_2421);
and U4095 (N_4095,N_44,N_105);
nand U4096 (N_4096,N_422,N_2138);
and U4097 (N_4097,N_1834,N_1866);
nand U4098 (N_4098,N_2167,N_1289);
and U4099 (N_4099,N_1756,N_2093);
or U4100 (N_4100,N_699,N_947);
nand U4101 (N_4101,N_1576,N_1289);
nor U4102 (N_4102,N_2426,N_1387);
and U4103 (N_4103,N_2274,N_1);
nor U4104 (N_4104,N_1111,N_2430);
or U4105 (N_4105,N_1736,N_38);
nand U4106 (N_4106,N_2385,N_2266);
nor U4107 (N_4107,N_969,N_545);
and U4108 (N_4108,N_1905,N_2489);
nand U4109 (N_4109,N_1936,N_1085);
nor U4110 (N_4110,N_22,N_1720);
nor U4111 (N_4111,N_626,N_15);
nand U4112 (N_4112,N_492,N_572);
or U4113 (N_4113,N_994,N_745);
nand U4114 (N_4114,N_1002,N_1763);
or U4115 (N_4115,N_155,N_719);
or U4116 (N_4116,N_158,N_63);
nand U4117 (N_4117,N_1295,N_371);
nand U4118 (N_4118,N_914,N_1748);
and U4119 (N_4119,N_2219,N_455);
or U4120 (N_4120,N_102,N_173);
or U4121 (N_4121,N_1658,N_2395);
or U4122 (N_4122,N_1142,N_1344);
nand U4123 (N_4123,N_2479,N_1604);
nor U4124 (N_4124,N_2229,N_856);
or U4125 (N_4125,N_2014,N_377);
or U4126 (N_4126,N_316,N_2020);
and U4127 (N_4127,N_574,N_1180);
and U4128 (N_4128,N_311,N_2139);
and U4129 (N_4129,N_2003,N_1876);
or U4130 (N_4130,N_682,N_545);
and U4131 (N_4131,N_1482,N_687);
nor U4132 (N_4132,N_2412,N_2094);
and U4133 (N_4133,N_2398,N_465);
nor U4134 (N_4134,N_1313,N_2367);
nor U4135 (N_4135,N_1330,N_473);
nor U4136 (N_4136,N_373,N_1674);
nor U4137 (N_4137,N_447,N_282);
nand U4138 (N_4138,N_1480,N_1784);
xor U4139 (N_4139,N_875,N_2148);
nand U4140 (N_4140,N_2300,N_1889);
or U4141 (N_4141,N_1340,N_106);
or U4142 (N_4142,N_330,N_1605);
and U4143 (N_4143,N_519,N_612);
nand U4144 (N_4144,N_1447,N_960);
and U4145 (N_4145,N_2471,N_1991);
nor U4146 (N_4146,N_2277,N_2042);
nand U4147 (N_4147,N_1929,N_2218);
nor U4148 (N_4148,N_2459,N_997);
and U4149 (N_4149,N_898,N_1428);
or U4150 (N_4150,N_1622,N_196);
or U4151 (N_4151,N_1706,N_626);
nand U4152 (N_4152,N_2066,N_2349);
nand U4153 (N_4153,N_983,N_800);
nand U4154 (N_4154,N_1476,N_2143);
or U4155 (N_4155,N_1135,N_1740);
and U4156 (N_4156,N_1428,N_2123);
nand U4157 (N_4157,N_646,N_2458);
and U4158 (N_4158,N_1884,N_1285);
nor U4159 (N_4159,N_2179,N_931);
or U4160 (N_4160,N_537,N_86);
nand U4161 (N_4161,N_74,N_957);
nor U4162 (N_4162,N_116,N_1032);
and U4163 (N_4163,N_1811,N_2292);
or U4164 (N_4164,N_1086,N_1365);
and U4165 (N_4165,N_289,N_1645);
xor U4166 (N_4166,N_1386,N_1321);
nor U4167 (N_4167,N_314,N_1316);
or U4168 (N_4168,N_359,N_2240);
nand U4169 (N_4169,N_1830,N_873);
and U4170 (N_4170,N_482,N_1824);
and U4171 (N_4171,N_1549,N_2388);
nor U4172 (N_4172,N_1215,N_2489);
nand U4173 (N_4173,N_1366,N_463);
and U4174 (N_4174,N_546,N_341);
nand U4175 (N_4175,N_1208,N_444);
or U4176 (N_4176,N_1377,N_266);
or U4177 (N_4177,N_2173,N_2055);
nor U4178 (N_4178,N_19,N_1071);
or U4179 (N_4179,N_1077,N_357);
or U4180 (N_4180,N_2064,N_848);
or U4181 (N_4181,N_2121,N_989);
nor U4182 (N_4182,N_1277,N_1970);
nor U4183 (N_4183,N_1777,N_1878);
and U4184 (N_4184,N_1546,N_752);
or U4185 (N_4185,N_2434,N_1809);
nor U4186 (N_4186,N_97,N_1417);
or U4187 (N_4187,N_213,N_1184);
nor U4188 (N_4188,N_2021,N_1467);
or U4189 (N_4189,N_370,N_82);
nand U4190 (N_4190,N_1540,N_1910);
and U4191 (N_4191,N_670,N_560);
or U4192 (N_4192,N_754,N_1716);
or U4193 (N_4193,N_789,N_1796);
or U4194 (N_4194,N_1470,N_726);
nor U4195 (N_4195,N_534,N_2065);
or U4196 (N_4196,N_2326,N_1935);
or U4197 (N_4197,N_1062,N_971);
or U4198 (N_4198,N_2425,N_1303);
nor U4199 (N_4199,N_1968,N_1073);
or U4200 (N_4200,N_872,N_1518);
nor U4201 (N_4201,N_2439,N_489);
nand U4202 (N_4202,N_208,N_17);
or U4203 (N_4203,N_1079,N_791);
xnor U4204 (N_4204,N_1170,N_1762);
nor U4205 (N_4205,N_2495,N_2410);
and U4206 (N_4206,N_920,N_107);
nand U4207 (N_4207,N_392,N_594);
and U4208 (N_4208,N_559,N_1241);
and U4209 (N_4209,N_338,N_1706);
nand U4210 (N_4210,N_2045,N_165);
xor U4211 (N_4211,N_2034,N_569);
and U4212 (N_4212,N_2398,N_463);
and U4213 (N_4213,N_974,N_1131);
nor U4214 (N_4214,N_1746,N_2496);
nand U4215 (N_4215,N_1455,N_360);
nand U4216 (N_4216,N_2041,N_234);
nand U4217 (N_4217,N_1383,N_438);
nand U4218 (N_4218,N_637,N_2176);
or U4219 (N_4219,N_1928,N_488);
or U4220 (N_4220,N_635,N_416);
or U4221 (N_4221,N_166,N_580);
and U4222 (N_4222,N_90,N_1535);
nor U4223 (N_4223,N_614,N_910);
and U4224 (N_4224,N_669,N_1799);
and U4225 (N_4225,N_1179,N_2230);
or U4226 (N_4226,N_1812,N_1169);
nor U4227 (N_4227,N_321,N_48);
nor U4228 (N_4228,N_1633,N_612);
nor U4229 (N_4229,N_2213,N_1542);
nand U4230 (N_4230,N_223,N_1539);
nor U4231 (N_4231,N_2456,N_104);
and U4232 (N_4232,N_810,N_653);
nand U4233 (N_4233,N_1586,N_1907);
nand U4234 (N_4234,N_1579,N_799);
or U4235 (N_4235,N_2370,N_923);
nand U4236 (N_4236,N_112,N_620);
xnor U4237 (N_4237,N_1873,N_550);
nor U4238 (N_4238,N_1606,N_1711);
nand U4239 (N_4239,N_1591,N_2328);
nand U4240 (N_4240,N_54,N_475);
and U4241 (N_4241,N_2208,N_2223);
nor U4242 (N_4242,N_379,N_1584);
nand U4243 (N_4243,N_122,N_1313);
nor U4244 (N_4244,N_974,N_758);
and U4245 (N_4245,N_2163,N_231);
or U4246 (N_4246,N_1047,N_228);
and U4247 (N_4247,N_1673,N_98);
and U4248 (N_4248,N_84,N_2098);
and U4249 (N_4249,N_2336,N_595);
nor U4250 (N_4250,N_1093,N_1907);
or U4251 (N_4251,N_1020,N_1632);
nand U4252 (N_4252,N_1016,N_322);
and U4253 (N_4253,N_2001,N_439);
nor U4254 (N_4254,N_2087,N_525);
nor U4255 (N_4255,N_1239,N_1391);
or U4256 (N_4256,N_2072,N_952);
nor U4257 (N_4257,N_2035,N_464);
and U4258 (N_4258,N_1795,N_2393);
nor U4259 (N_4259,N_1009,N_2409);
and U4260 (N_4260,N_1944,N_2433);
and U4261 (N_4261,N_1355,N_712);
nand U4262 (N_4262,N_228,N_1289);
nand U4263 (N_4263,N_91,N_2036);
and U4264 (N_4264,N_56,N_1208);
and U4265 (N_4265,N_1931,N_2117);
nand U4266 (N_4266,N_1715,N_413);
nand U4267 (N_4267,N_2112,N_251);
xnor U4268 (N_4268,N_414,N_1381);
or U4269 (N_4269,N_1859,N_1280);
or U4270 (N_4270,N_882,N_1263);
or U4271 (N_4271,N_262,N_2331);
nand U4272 (N_4272,N_1210,N_951);
or U4273 (N_4273,N_1707,N_2224);
nand U4274 (N_4274,N_2072,N_938);
nand U4275 (N_4275,N_1352,N_1278);
and U4276 (N_4276,N_1229,N_1821);
nand U4277 (N_4277,N_1177,N_1887);
or U4278 (N_4278,N_1117,N_2077);
nand U4279 (N_4279,N_2323,N_1765);
or U4280 (N_4280,N_2229,N_314);
and U4281 (N_4281,N_576,N_1780);
nor U4282 (N_4282,N_748,N_1972);
nand U4283 (N_4283,N_2202,N_1353);
and U4284 (N_4284,N_717,N_2123);
nand U4285 (N_4285,N_2327,N_1361);
and U4286 (N_4286,N_1590,N_1532);
or U4287 (N_4287,N_31,N_1670);
and U4288 (N_4288,N_66,N_2467);
and U4289 (N_4289,N_1016,N_207);
or U4290 (N_4290,N_1073,N_2473);
or U4291 (N_4291,N_336,N_2177);
nand U4292 (N_4292,N_1575,N_1496);
nor U4293 (N_4293,N_491,N_566);
nand U4294 (N_4294,N_2343,N_936);
or U4295 (N_4295,N_585,N_1226);
nor U4296 (N_4296,N_1328,N_397);
or U4297 (N_4297,N_1993,N_1109);
nand U4298 (N_4298,N_2125,N_680);
xor U4299 (N_4299,N_1762,N_1216);
or U4300 (N_4300,N_1648,N_1056);
nor U4301 (N_4301,N_70,N_468);
nor U4302 (N_4302,N_1297,N_143);
and U4303 (N_4303,N_1589,N_2288);
or U4304 (N_4304,N_2320,N_1209);
nor U4305 (N_4305,N_403,N_198);
or U4306 (N_4306,N_449,N_2280);
nor U4307 (N_4307,N_262,N_950);
or U4308 (N_4308,N_1016,N_2345);
and U4309 (N_4309,N_78,N_242);
or U4310 (N_4310,N_1456,N_43);
nand U4311 (N_4311,N_191,N_1706);
or U4312 (N_4312,N_1767,N_2340);
nor U4313 (N_4313,N_2490,N_847);
nor U4314 (N_4314,N_177,N_1856);
or U4315 (N_4315,N_1133,N_2461);
and U4316 (N_4316,N_801,N_717);
or U4317 (N_4317,N_1873,N_801);
and U4318 (N_4318,N_650,N_528);
nor U4319 (N_4319,N_699,N_1131);
and U4320 (N_4320,N_1446,N_1617);
nor U4321 (N_4321,N_2043,N_2273);
or U4322 (N_4322,N_937,N_1466);
nand U4323 (N_4323,N_2465,N_1334);
and U4324 (N_4324,N_1865,N_333);
or U4325 (N_4325,N_819,N_738);
or U4326 (N_4326,N_842,N_338);
nor U4327 (N_4327,N_1362,N_1187);
nand U4328 (N_4328,N_573,N_1846);
nor U4329 (N_4329,N_59,N_901);
nor U4330 (N_4330,N_893,N_147);
and U4331 (N_4331,N_1433,N_2037);
or U4332 (N_4332,N_820,N_158);
nor U4333 (N_4333,N_2044,N_2096);
or U4334 (N_4334,N_2342,N_1024);
nand U4335 (N_4335,N_1176,N_835);
nand U4336 (N_4336,N_2381,N_737);
nand U4337 (N_4337,N_1393,N_1921);
or U4338 (N_4338,N_1876,N_938);
xor U4339 (N_4339,N_1492,N_1239);
and U4340 (N_4340,N_1779,N_2177);
or U4341 (N_4341,N_418,N_1867);
or U4342 (N_4342,N_1706,N_1593);
nor U4343 (N_4343,N_1872,N_254);
nor U4344 (N_4344,N_348,N_1570);
and U4345 (N_4345,N_2024,N_1690);
nor U4346 (N_4346,N_1932,N_778);
and U4347 (N_4347,N_1484,N_1531);
or U4348 (N_4348,N_411,N_1634);
and U4349 (N_4349,N_526,N_2433);
and U4350 (N_4350,N_804,N_1956);
and U4351 (N_4351,N_639,N_1828);
nor U4352 (N_4352,N_1609,N_984);
or U4353 (N_4353,N_1139,N_1115);
or U4354 (N_4354,N_72,N_318);
or U4355 (N_4355,N_884,N_865);
or U4356 (N_4356,N_1656,N_794);
or U4357 (N_4357,N_52,N_1699);
and U4358 (N_4358,N_2316,N_1320);
and U4359 (N_4359,N_1449,N_1044);
nand U4360 (N_4360,N_1009,N_2321);
nand U4361 (N_4361,N_321,N_874);
or U4362 (N_4362,N_2200,N_714);
nand U4363 (N_4363,N_293,N_181);
nand U4364 (N_4364,N_223,N_1057);
xnor U4365 (N_4365,N_1149,N_2265);
nand U4366 (N_4366,N_258,N_537);
nor U4367 (N_4367,N_1775,N_1210);
nand U4368 (N_4368,N_1827,N_1096);
nand U4369 (N_4369,N_742,N_2079);
nand U4370 (N_4370,N_1833,N_1852);
xnor U4371 (N_4371,N_2267,N_79);
or U4372 (N_4372,N_1460,N_700);
and U4373 (N_4373,N_1349,N_904);
and U4374 (N_4374,N_2189,N_1885);
nor U4375 (N_4375,N_1657,N_2286);
nor U4376 (N_4376,N_2363,N_919);
or U4377 (N_4377,N_2284,N_1316);
nor U4378 (N_4378,N_769,N_1378);
nor U4379 (N_4379,N_1420,N_2448);
nand U4380 (N_4380,N_1716,N_600);
or U4381 (N_4381,N_1483,N_165);
or U4382 (N_4382,N_1983,N_282);
or U4383 (N_4383,N_838,N_444);
nand U4384 (N_4384,N_2031,N_1167);
nor U4385 (N_4385,N_1479,N_1627);
nor U4386 (N_4386,N_1271,N_258);
or U4387 (N_4387,N_1672,N_1444);
nor U4388 (N_4388,N_2461,N_611);
or U4389 (N_4389,N_1659,N_1859);
nand U4390 (N_4390,N_1009,N_1377);
nand U4391 (N_4391,N_2485,N_437);
and U4392 (N_4392,N_420,N_160);
nor U4393 (N_4393,N_539,N_837);
or U4394 (N_4394,N_2335,N_1424);
nor U4395 (N_4395,N_219,N_1362);
and U4396 (N_4396,N_923,N_441);
nand U4397 (N_4397,N_2175,N_944);
xnor U4398 (N_4398,N_1088,N_1596);
nand U4399 (N_4399,N_280,N_2485);
nor U4400 (N_4400,N_814,N_194);
nand U4401 (N_4401,N_628,N_876);
and U4402 (N_4402,N_763,N_891);
nor U4403 (N_4403,N_216,N_1890);
nor U4404 (N_4404,N_2409,N_332);
and U4405 (N_4405,N_914,N_2277);
nor U4406 (N_4406,N_1741,N_453);
or U4407 (N_4407,N_1508,N_2094);
and U4408 (N_4408,N_1193,N_1492);
nor U4409 (N_4409,N_2298,N_1559);
or U4410 (N_4410,N_1945,N_197);
or U4411 (N_4411,N_1443,N_1346);
nand U4412 (N_4412,N_2237,N_1575);
and U4413 (N_4413,N_1640,N_2085);
nor U4414 (N_4414,N_2077,N_13);
and U4415 (N_4415,N_1123,N_1234);
and U4416 (N_4416,N_1270,N_722);
and U4417 (N_4417,N_621,N_2347);
and U4418 (N_4418,N_172,N_2117);
nand U4419 (N_4419,N_1621,N_2390);
and U4420 (N_4420,N_2038,N_2056);
xor U4421 (N_4421,N_143,N_2080);
or U4422 (N_4422,N_1048,N_680);
nand U4423 (N_4423,N_1387,N_1570);
and U4424 (N_4424,N_1904,N_2138);
nand U4425 (N_4425,N_1185,N_1022);
nand U4426 (N_4426,N_159,N_567);
and U4427 (N_4427,N_232,N_2406);
or U4428 (N_4428,N_1116,N_106);
nor U4429 (N_4429,N_41,N_1125);
or U4430 (N_4430,N_1917,N_1131);
nand U4431 (N_4431,N_969,N_353);
nor U4432 (N_4432,N_2146,N_555);
or U4433 (N_4433,N_2112,N_1091);
or U4434 (N_4434,N_2459,N_1794);
nor U4435 (N_4435,N_2027,N_86);
and U4436 (N_4436,N_1659,N_347);
and U4437 (N_4437,N_2075,N_345);
nand U4438 (N_4438,N_2324,N_1054);
nand U4439 (N_4439,N_1484,N_1581);
and U4440 (N_4440,N_1711,N_1157);
xor U4441 (N_4441,N_1136,N_759);
and U4442 (N_4442,N_2454,N_522);
nor U4443 (N_4443,N_1755,N_1965);
or U4444 (N_4444,N_954,N_224);
and U4445 (N_4445,N_2211,N_1479);
and U4446 (N_4446,N_1281,N_610);
or U4447 (N_4447,N_1512,N_888);
xnor U4448 (N_4448,N_281,N_497);
nor U4449 (N_4449,N_1527,N_1617);
or U4450 (N_4450,N_785,N_1024);
nor U4451 (N_4451,N_1758,N_955);
or U4452 (N_4452,N_377,N_80);
and U4453 (N_4453,N_1695,N_1121);
nor U4454 (N_4454,N_1289,N_1196);
and U4455 (N_4455,N_1529,N_1499);
nor U4456 (N_4456,N_2157,N_497);
nand U4457 (N_4457,N_1990,N_423);
nor U4458 (N_4458,N_2368,N_2045);
or U4459 (N_4459,N_440,N_2329);
and U4460 (N_4460,N_2316,N_1263);
and U4461 (N_4461,N_1518,N_601);
nor U4462 (N_4462,N_1206,N_1353);
nor U4463 (N_4463,N_350,N_358);
nand U4464 (N_4464,N_568,N_2324);
or U4465 (N_4465,N_1953,N_524);
nand U4466 (N_4466,N_406,N_1677);
and U4467 (N_4467,N_609,N_118);
or U4468 (N_4468,N_422,N_1703);
and U4469 (N_4469,N_88,N_1984);
nor U4470 (N_4470,N_1973,N_467);
or U4471 (N_4471,N_1145,N_709);
and U4472 (N_4472,N_90,N_2092);
or U4473 (N_4473,N_127,N_2289);
xor U4474 (N_4474,N_2497,N_1764);
nor U4475 (N_4475,N_279,N_1677);
or U4476 (N_4476,N_1904,N_929);
nand U4477 (N_4477,N_1606,N_241);
nand U4478 (N_4478,N_2253,N_1243);
and U4479 (N_4479,N_923,N_1644);
and U4480 (N_4480,N_2031,N_1362);
and U4481 (N_4481,N_1038,N_250);
nor U4482 (N_4482,N_2195,N_61);
nand U4483 (N_4483,N_1982,N_2378);
and U4484 (N_4484,N_1573,N_822);
or U4485 (N_4485,N_1174,N_1825);
nor U4486 (N_4486,N_1034,N_1225);
xnor U4487 (N_4487,N_2345,N_2099);
nor U4488 (N_4488,N_540,N_481);
nand U4489 (N_4489,N_1290,N_1081);
and U4490 (N_4490,N_1691,N_911);
nand U4491 (N_4491,N_484,N_2354);
nor U4492 (N_4492,N_2254,N_1970);
nand U4493 (N_4493,N_2341,N_11);
and U4494 (N_4494,N_1518,N_250);
and U4495 (N_4495,N_103,N_49);
and U4496 (N_4496,N_560,N_431);
nand U4497 (N_4497,N_707,N_847);
nand U4498 (N_4498,N_2150,N_2);
nor U4499 (N_4499,N_1645,N_306);
or U4500 (N_4500,N_291,N_1641);
nand U4501 (N_4501,N_256,N_1280);
nor U4502 (N_4502,N_2366,N_1836);
nand U4503 (N_4503,N_360,N_41);
nand U4504 (N_4504,N_1666,N_638);
or U4505 (N_4505,N_941,N_2480);
nor U4506 (N_4506,N_1763,N_189);
nor U4507 (N_4507,N_677,N_1709);
nand U4508 (N_4508,N_1126,N_1348);
nand U4509 (N_4509,N_1076,N_147);
nand U4510 (N_4510,N_1086,N_2204);
or U4511 (N_4511,N_2352,N_10);
nor U4512 (N_4512,N_258,N_2465);
or U4513 (N_4513,N_867,N_1584);
and U4514 (N_4514,N_2271,N_1014);
xnor U4515 (N_4515,N_1345,N_778);
nor U4516 (N_4516,N_1648,N_832);
nor U4517 (N_4517,N_923,N_525);
and U4518 (N_4518,N_283,N_1338);
nor U4519 (N_4519,N_1902,N_2133);
and U4520 (N_4520,N_658,N_222);
or U4521 (N_4521,N_1716,N_1545);
and U4522 (N_4522,N_1178,N_1249);
xor U4523 (N_4523,N_139,N_2335);
nor U4524 (N_4524,N_158,N_1244);
or U4525 (N_4525,N_906,N_793);
nand U4526 (N_4526,N_1547,N_807);
nor U4527 (N_4527,N_1890,N_1016);
and U4528 (N_4528,N_1227,N_1974);
nor U4529 (N_4529,N_1228,N_1500);
nand U4530 (N_4530,N_1193,N_556);
nand U4531 (N_4531,N_693,N_1483);
nor U4532 (N_4532,N_2023,N_2141);
and U4533 (N_4533,N_1478,N_1224);
and U4534 (N_4534,N_1392,N_357);
xor U4535 (N_4535,N_1570,N_813);
or U4536 (N_4536,N_2128,N_706);
nor U4537 (N_4537,N_1383,N_141);
or U4538 (N_4538,N_195,N_369);
nor U4539 (N_4539,N_1467,N_1370);
or U4540 (N_4540,N_1850,N_1081);
nand U4541 (N_4541,N_1946,N_1219);
or U4542 (N_4542,N_2380,N_1131);
or U4543 (N_4543,N_2305,N_1711);
nand U4544 (N_4544,N_2216,N_1740);
or U4545 (N_4545,N_2158,N_31);
nor U4546 (N_4546,N_1446,N_218);
nand U4547 (N_4547,N_449,N_650);
nand U4548 (N_4548,N_2229,N_2143);
nor U4549 (N_4549,N_961,N_403);
nor U4550 (N_4550,N_1373,N_2237);
nor U4551 (N_4551,N_2142,N_55);
or U4552 (N_4552,N_342,N_156);
or U4553 (N_4553,N_293,N_668);
nor U4554 (N_4554,N_2016,N_2093);
nand U4555 (N_4555,N_430,N_958);
nor U4556 (N_4556,N_756,N_396);
nand U4557 (N_4557,N_2455,N_592);
nand U4558 (N_4558,N_546,N_780);
nor U4559 (N_4559,N_1167,N_274);
or U4560 (N_4560,N_2287,N_1840);
nand U4561 (N_4561,N_1454,N_532);
nor U4562 (N_4562,N_2087,N_823);
nor U4563 (N_4563,N_876,N_1404);
and U4564 (N_4564,N_693,N_377);
or U4565 (N_4565,N_250,N_319);
or U4566 (N_4566,N_1139,N_1014);
nand U4567 (N_4567,N_1930,N_653);
or U4568 (N_4568,N_391,N_1681);
nor U4569 (N_4569,N_2232,N_1392);
or U4570 (N_4570,N_2136,N_2383);
nor U4571 (N_4571,N_722,N_1561);
or U4572 (N_4572,N_214,N_868);
nor U4573 (N_4573,N_1512,N_1684);
nor U4574 (N_4574,N_803,N_2406);
and U4575 (N_4575,N_1678,N_1750);
nor U4576 (N_4576,N_1471,N_859);
nor U4577 (N_4577,N_1164,N_1452);
and U4578 (N_4578,N_1769,N_1896);
and U4579 (N_4579,N_1403,N_787);
and U4580 (N_4580,N_1455,N_1104);
nor U4581 (N_4581,N_1763,N_1276);
nor U4582 (N_4582,N_554,N_1013);
or U4583 (N_4583,N_1497,N_1255);
and U4584 (N_4584,N_227,N_244);
nor U4585 (N_4585,N_1740,N_1829);
and U4586 (N_4586,N_1398,N_1079);
and U4587 (N_4587,N_47,N_2435);
or U4588 (N_4588,N_1638,N_258);
or U4589 (N_4589,N_1530,N_304);
nand U4590 (N_4590,N_944,N_132);
nand U4591 (N_4591,N_1358,N_1860);
nor U4592 (N_4592,N_1583,N_478);
and U4593 (N_4593,N_2126,N_1727);
or U4594 (N_4594,N_515,N_617);
nand U4595 (N_4595,N_184,N_1055);
xnor U4596 (N_4596,N_768,N_1579);
and U4597 (N_4597,N_809,N_288);
or U4598 (N_4598,N_2474,N_203);
nor U4599 (N_4599,N_1296,N_2025);
or U4600 (N_4600,N_2351,N_826);
nor U4601 (N_4601,N_2014,N_39);
or U4602 (N_4602,N_160,N_604);
xor U4603 (N_4603,N_2432,N_436);
and U4604 (N_4604,N_1906,N_635);
nor U4605 (N_4605,N_934,N_597);
nor U4606 (N_4606,N_1535,N_1520);
nor U4607 (N_4607,N_623,N_603);
and U4608 (N_4608,N_875,N_1780);
or U4609 (N_4609,N_1125,N_610);
and U4610 (N_4610,N_486,N_1803);
nand U4611 (N_4611,N_77,N_2432);
nand U4612 (N_4612,N_352,N_397);
and U4613 (N_4613,N_286,N_1911);
or U4614 (N_4614,N_1500,N_34);
or U4615 (N_4615,N_1622,N_199);
nor U4616 (N_4616,N_1838,N_2306);
nor U4617 (N_4617,N_246,N_414);
and U4618 (N_4618,N_1475,N_1645);
nor U4619 (N_4619,N_1690,N_2076);
nor U4620 (N_4620,N_1400,N_709);
xor U4621 (N_4621,N_1376,N_2191);
nand U4622 (N_4622,N_52,N_744);
nor U4623 (N_4623,N_1052,N_2124);
nand U4624 (N_4624,N_760,N_1225);
and U4625 (N_4625,N_534,N_1673);
or U4626 (N_4626,N_928,N_2147);
nand U4627 (N_4627,N_1281,N_2317);
nand U4628 (N_4628,N_106,N_1325);
or U4629 (N_4629,N_1083,N_1577);
or U4630 (N_4630,N_1666,N_1274);
nor U4631 (N_4631,N_653,N_1075);
nor U4632 (N_4632,N_83,N_2281);
nor U4633 (N_4633,N_2395,N_2399);
nand U4634 (N_4634,N_539,N_81);
nand U4635 (N_4635,N_774,N_2285);
nand U4636 (N_4636,N_579,N_38);
or U4637 (N_4637,N_2214,N_733);
or U4638 (N_4638,N_1536,N_1692);
or U4639 (N_4639,N_2253,N_2393);
or U4640 (N_4640,N_1370,N_1738);
or U4641 (N_4641,N_22,N_1351);
or U4642 (N_4642,N_2312,N_1041);
nand U4643 (N_4643,N_2369,N_932);
or U4644 (N_4644,N_887,N_1475);
and U4645 (N_4645,N_1931,N_2296);
xnor U4646 (N_4646,N_2252,N_1180);
and U4647 (N_4647,N_484,N_2002);
and U4648 (N_4648,N_1642,N_2446);
or U4649 (N_4649,N_657,N_2147);
or U4650 (N_4650,N_891,N_1858);
or U4651 (N_4651,N_917,N_1460);
nand U4652 (N_4652,N_3,N_1351);
nor U4653 (N_4653,N_651,N_2477);
and U4654 (N_4654,N_1061,N_1253);
nand U4655 (N_4655,N_372,N_934);
and U4656 (N_4656,N_932,N_2236);
and U4657 (N_4657,N_1354,N_680);
nand U4658 (N_4658,N_902,N_1916);
and U4659 (N_4659,N_399,N_268);
nand U4660 (N_4660,N_702,N_543);
nand U4661 (N_4661,N_610,N_2476);
and U4662 (N_4662,N_2150,N_637);
nand U4663 (N_4663,N_1862,N_1503);
and U4664 (N_4664,N_668,N_1279);
or U4665 (N_4665,N_318,N_2079);
nand U4666 (N_4666,N_390,N_2130);
or U4667 (N_4667,N_442,N_2096);
and U4668 (N_4668,N_2251,N_339);
or U4669 (N_4669,N_434,N_2019);
nor U4670 (N_4670,N_210,N_1451);
nand U4671 (N_4671,N_1802,N_929);
and U4672 (N_4672,N_4,N_2165);
and U4673 (N_4673,N_969,N_1607);
nand U4674 (N_4674,N_2019,N_130);
nand U4675 (N_4675,N_873,N_2327);
nand U4676 (N_4676,N_1242,N_1138);
nand U4677 (N_4677,N_463,N_216);
xnor U4678 (N_4678,N_610,N_167);
nor U4679 (N_4679,N_667,N_472);
nand U4680 (N_4680,N_260,N_1406);
nor U4681 (N_4681,N_1601,N_2070);
or U4682 (N_4682,N_1699,N_1861);
nor U4683 (N_4683,N_272,N_901);
nand U4684 (N_4684,N_1005,N_2371);
and U4685 (N_4685,N_1430,N_315);
or U4686 (N_4686,N_1167,N_1702);
nor U4687 (N_4687,N_2461,N_199);
nor U4688 (N_4688,N_2293,N_2294);
nor U4689 (N_4689,N_1765,N_1250);
or U4690 (N_4690,N_210,N_2008);
and U4691 (N_4691,N_654,N_1042);
and U4692 (N_4692,N_1506,N_144);
and U4693 (N_4693,N_556,N_2406);
and U4694 (N_4694,N_1914,N_432);
nand U4695 (N_4695,N_1362,N_885);
and U4696 (N_4696,N_2071,N_1905);
or U4697 (N_4697,N_2325,N_842);
xnor U4698 (N_4698,N_2057,N_166);
or U4699 (N_4699,N_2133,N_1322);
or U4700 (N_4700,N_1979,N_1013);
and U4701 (N_4701,N_908,N_2159);
nor U4702 (N_4702,N_2120,N_908);
nor U4703 (N_4703,N_2323,N_1962);
nor U4704 (N_4704,N_972,N_1420);
nor U4705 (N_4705,N_425,N_2431);
nor U4706 (N_4706,N_176,N_1676);
nor U4707 (N_4707,N_1967,N_1418);
nor U4708 (N_4708,N_1065,N_1368);
and U4709 (N_4709,N_1762,N_588);
or U4710 (N_4710,N_1911,N_925);
or U4711 (N_4711,N_1954,N_412);
or U4712 (N_4712,N_2193,N_2423);
and U4713 (N_4713,N_1974,N_1049);
or U4714 (N_4714,N_776,N_1903);
or U4715 (N_4715,N_90,N_125);
and U4716 (N_4716,N_2337,N_1369);
nand U4717 (N_4717,N_908,N_586);
nand U4718 (N_4718,N_796,N_563);
nand U4719 (N_4719,N_1161,N_1358);
nand U4720 (N_4720,N_83,N_2048);
xor U4721 (N_4721,N_1184,N_1679);
or U4722 (N_4722,N_1786,N_2343);
and U4723 (N_4723,N_1248,N_734);
nand U4724 (N_4724,N_399,N_840);
nor U4725 (N_4725,N_615,N_627);
and U4726 (N_4726,N_700,N_712);
nor U4727 (N_4727,N_565,N_1337);
nand U4728 (N_4728,N_184,N_951);
nand U4729 (N_4729,N_1011,N_1757);
nand U4730 (N_4730,N_2278,N_2251);
nor U4731 (N_4731,N_1548,N_2414);
or U4732 (N_4732,N_1614,N_1805);
nor U4733 (N_4733,N_1909,N_632);
and U4734 (N_4734,N_2277,N_2330);
nand U4735 (N_4735,N_2291,N_751);
and U4736 (N_4736,N_62,N_213);
or U4737 (N_4737,N_1994,N_1101);
or U4738 (N_4738,N_644,N_1171);
nor U4739 (N_4739,N_868,N_1702);
nand U4740 (N_4740,N_2434,N_2489);
nor U4741 (N_4741,N_719,N_2388);
nand U4742 (N_4742,N_1454,N_1658);
nand U4743 (N_4743,N_2004,N_1173);
or U4744 (N_4744,N_2227,N_2485);
and U4745 (N_4745,N_98,N_1556);
or U4746 (N_4746,N_597,N_993);
or U4747 (N_4747,N_1156,N_1084);
and U4748 (N_4748,N_1002,N_2082);
and U4749 (N_4749,N_982,N_882);
or U4750 (N_4750,N_677,N_1220);
nand U4751 (N_4751,N_2147,N_1309);
and U4752 (N_4752,N_2028,N_1547);
or U4753 (N_4753,N_867,N_1603);
and U4754 (N_4754,N_468,N_2227);
nor U4755 (N_4755,N_693,N_1718);
nor U4756 (N_4756,N_1643,N_163);
and U4757 (N_4757,N_205,N_2156);
or U4758 (N_4758,N_1543,N_2110);
or U4759 (N_4759,N_1692,N_2269);
or U4760 (N_4760,N_1515,N_2422);
xor U4761 (N_4761,N_2262,N_1948);
or U4762 (N_4762,N_2354,N_1077);
nand U4763 (N_4763,N_675,N_2044);
and U4764 (N_4764,N_1246,N_338);
nand U4765 (N_4765,N_1821,N_1348);
nand U4766 (N_4766,N_1941,N_328);
xnor U4767 (N_4767,N_1177,N_611);
nand U4768 (N_4768,N_80,N_2486);
or U4769 (N_4769,N_616,N_1299);
or U4770 (N_4770,N_2205,N_1356);
and U4771 (N_4771,N_1149,N_2493);
nor U4772 (N_4772,N_416,N_397);
or U4773 (N_4773,N_614,N_1143);
and U4774 (N_4774,N_403,N_610);
nand U4775 (N_4775,N_1802,N_721);
and U4776 (N_4776,N_1004,N_870);
nand U4777 (N_4777,N_2188,N_1466);
nand U4778 (N_4778,N_1432,N_1354);
nand U4779 (N_4779,N_1400,N_792);
nor U4780 (N_4780,N_1225,N_1020);
nor U4781 (N_4781,N_1536,N_2452);
or U4782 (N_4782,N_1288,N_114);
nand U4783 (N_4783,N_147,N_2189);
or U4784 (N_4784,N_1648,N_579);
or U4785 (N_4785,N_2270,N_1075);
nand U4786 (N_4786,N_990,N_363);
and U4787 (N_4787,N_343,N_1874);
nor U4788 (N_4788,N_1109,N_1880);
and U4789 (N_4789,N_980,N_1242);
nand U4790 (N_4790,N_643,N_1483);
nor U4791 (N_4791,N_964,N_1835);
xnor U4792 (N_4792,N_1686,N_655);
or U4793 (N_4793,N_2107,N_440);
nand U4794 (N_4794,N_545,N_650);
or U4795 (N_4795,N_1600,N_1703);
and U4796 (N_4796,N_1269,N_2208);
and U4797 (N_4797,N_1253,N_1152);
nor U4798 (N_4798,N_1940,N_882);
or U4799 (N_4799,N_2473,N_327);
or U4800 (N_4800,N_1131,N_904);
nand U4801 (N_4801,N_1524,N_1291);
or U4802 (N_4802,N_845,N_503);
nand U4803 (N_4803,N_516,N_1426);
nor U4804 (N_4804,N_844,N_2050);
nor U4805 (N_4805,N_1890,N_270);
and U4806 (N_4806,N_601,N_1317);
or U4807 (N_4807,N_1037,N_1519);
and U4808 (N_4808,N_1878,N_29);
nor U4809 (N_4809,N_356,N_1029);
and U4810 (N_4810,N_1551,N_534);
or U4811 (N_4811,N_996,N_2003);
or U4812 (N_4812,N_1591,N_331);
nand U4813 (N_4813,N_1331,N_2135);
or U4814 (N_4814,N_1668,N_550);
or U4815 (N_4815,N_2491,N_1257);
and U4816 (N_4816,N_2404,N_47);
or U4817 (N_4817,N_659,N_141);
nand U4818 (N_4818,N_1306,N_11);
nor U4819 (N_4819,N_1776,N_176);
and U4820 (N_4820,N_1742,N_742);
nor U4821 (N_4821,N_1644,N_2216);
or U4822 (N_4822,N_2347,N_1018);
and U4823 (N_4823,N_1971,N_489);
nor U4824 (N_4824,N_733,N_129);
nor U4825 (N_4825,N_2087,N_1654);
xor U4826 (N_4826,N_1593,N_1002);
nand U4827 (N_4827,N_1288,N_655);
nor U4828 (N_4828,N_684,N_959);
and U4829 (N_4829,N_282,N_981);
and U4830 (N_4830,N_1374,N_1206);
and U4831 (N_4831,N_1486,N_396);
nand U4832 (N_4832,N_886,N_1410);
or U4833 (N_4833,N_2302,N_587);
or U4834 (N_4834,N_1799,N_1097);
or U4835 (N_4835,N_2422,N_1338);
nand U4836 (N_4836,N_2048,N_24);
nand U4837 (N_4837,N_1248,N_2453);
or U4838 (N_4838,N_525,N_1062);
and U4839 (N_4839,N_960,N_2354);
nor U4840 (N_4840,N_1173,N_2283);
nor U4841 (N_4841,N_1059,N_2255);
or U4842 (N_4842,N_387,N_579);
nand U4843 (N_4843,N_365,N_1425);
or U4844 (N_4844,N_582,N_1974);
or U4845 (N_4845,N_975,N_2064);
and U4846 (N_4846,N_1657,N_1433);
and U4847 (N_4847,N_1299,N_1675);
nand U4848 (N_4848,N_679,N_2397);
and U4849 (N_4849,N_408,N_2366);
and U4850 (N_4850,N_1957,N_1267);
and U4851 (N_4851,N_632,N_2454);
nor U4852 (N_4852,N_331,N_2497);
nand U4853 (N_4853,N_229,N_1891);
or U4854 (N_4854,N_220,N_2177);
nand U4855 (N_4855,N_2327,N_2163);
xnor U4856 (N_4856,N_849,N_84);
nor U4857 (N_4857,N_608,N_983);
nand U4858 (N_4858,N_1693,N_538);
nor U4859 (N_4859,N_2282,N_1029);
nor U4860 (N_4860,N_276,N_765);
and U4861 (N_4861,N_318,N_204);
nand U4862 (N_4862,N_809,N_1316);
and U4863 (N_4863,N_211,N_1586);
nor U4864 (N_4864,N_1482,N_2412);
or U4865 (N_4865,N_1001,N_1785);
nand U4866 (N_4866,N_351,N_2265);
or U4867 (N_4867,N_1214,N_2183);
and U4868 (N_4868,N_563,N_124);
nor U4869 (N_4869,N_2196,N_26);
nor U4870 (N_4870,N_14,N_1529);
nor U4871 (N_4871,N_1344,N_417);
or U4872 (N_4872,N_1204,N_434);
nand U4873 (N_4873,N_2140,N_1006);
and U4874 (N_4874,N_2487,N_549);
nand U4875 (N_4875,N_814,N_2410);
and U4876 (N_4876,N_931,N_2054);
nand U4877 (N_4877,N_411,N_1730);
nor U4878 (N_4878,N_2486,N_2018);
nand U4879 (N_4879,N_2076,N_1849);
and U4880 (N_4880,N_1700,N_972);
or U4881 (N_4881,N_1108,N_1575);
nand U4882 (N_4882,N_2397,N_2005);
nand U4883 (N_4883,N_1814,N_1859);
nand U4884 (N_4884,N_218,N_481);
nand U4885 (N_4885,N_238,N_1844);
nor U4886 (N_4886,N_1840,N_106);
and U4887 (N_4887,N_1211,N_710);
xor U4888 (N_4888,N_1440,N_2438);
or U4889 (N_4889,N_2142,N_83);
and U4890 (N_4890,N_2378,N_892);
or U4891 (N_4891,N_440,N_1784);
or U4892 (N_4892,N_1145,N_1766);
or U4893 (N_4893,N_1202,N_267);
or U4894 (N_4894,N_1884,N_2135);
nor U4895 (N_4895,N_2126,N_161);
nor U4896 (N_4896,N_1499,N_1165);
and U4897 (N_4897,N_46,N_804);
or U4898 (N_4898,N_883,N_1255);
nor U4899 (N_4899,N_9,N_2395);
and U4900 (N_4900,N_2145,N_2154);
or U4901 (N_4901,N_2480,N_744);
nand U4902 (N_4902,N_1521,N_2422);
and U4903 (N_4903,N_154,N_1094);
xnor U4904 (N_4904,N_818,N_2143);
or U4905 (N_4905,N_1252,N_2432);
and U4906 (N_4906,N_2073,N_971);
nand U4907 (N_4907,N_724,N_38);
nand U4908 (N_4908,N_892,N_1735);
nor U4909 (N_4909,N_610,N_1394);
nor U4910 (N_4910,N_1135,N_2243);
nor U4911 (N_4911,N_18,N_1912);
nand U4912 (N_4912,N_1006,N_650);
or U4913 (N_4913,N_2349,N_867);
nor U4914 (N_4914,N_2106,N_1318);
xnor U4915 (N_4915,N_1160,N_1808);
nor U4916 (N_4916,N_303,N_2059);
nand U4917 (N_4917,N_1920,N_756);
nand U4918 (N_4918,N_1281,N_1583);
and U4919 (N_4919,N_2268,N_1381);
or U4920 (N_4920,N_1026,N_1671);
nor U4921 (N_4921,N_1263,N_87);
or U4922 (N_4922,N_1194,N_955);
nor U4923 (N_4923,N_118,N_1022);
and U4924 (N_4924,N_1533,N_1750);
nand U4925 (N_4925,N_264,N_878);
nand U4926 (N_4926,N_1363,N_885);
nand U4927 (N_4927,N_502,N_1032);
nand U4928 (N_4928,N_1647,N_1527);
or U4929 (N_4929,N_867,N_1678);
and U4930 (N_4930,N_404,N_1073);
or U4931 (N_4931,N_1757,N_1908);
nand U4932 (N_4932,N_1603,N_1567);
or U4933 (N_4933,N_1864,N_1158);
or U4934 (N_4934,N_961,N_199);
or U4935 (N_4935,N_402,N_278);
xnor U4936 (N_4936,N_2468,N_2301);
nor U4937 (N_4937,N_1513,N_2060);
nand U4938 (N_4938,N_685,N_1401);
and U4939 (N_4939,N_176,N_1064);
or U4940 (N_4940,N_2296,N_2435);
nand U4941 (N_4941,N_988,N_7);
nand U4942 (N_4942,N_501,N_2335);
nand U4943 (N_4943,N_228,N_1002);
or U4944 (N_4944,N_231,N_1402);
and U4945 (N_4945,N_1484,N_500);
nor U4946 (N_4946,N_124,N_178);
and U4947 (N_4947,N_1612,N_1466);
or U4948 (N_4948,N_677,N_1891);
or U4949 (N_4949,N_876,N_1527);
or U4950 (N_4950,N_819,N_40);
nand U4951 (N_4951,N_989,N_1901);
and U4952 (N_4952,N_2097,N_1602);
nand U4953 (N_4953,N_1969,N_1904);
nand U4954 (N_4954,N_2145,N_1771);
and U4955 (N_4955,N_1832,N_2354);
nor U4956 (N_4956,N_183,N_552);
and U4957 (N_4957,N_10,N_589);
nor U4958 (N_4958,N_264,N_1503);
or U4959 (N_4959,N_843,N_247);
nand U4960 (N_4960,N_1214,N_1685);
nor U4961 (N_4961,N_956,N_2261);
nor U4962 (N_4962,N_1496,N_2248);
nand U4963 (N_4963,N_220,N_2370);
nor U4964 (N_4964,N_1513,N_1946);
nor U4965 (N_4965,N_1186,N_2168);
nand U4966 (N_4966,N_334,N_1745);
or U4967 (N_4967,N_1905,N_2436);
and U4968 (N_4968,N_1543,N_2401);
and U4969 (N_4969,N_2052,N_2016);
or U4970 (N_4970,N_2084,N_126);
and U4971 (N_4971,N_2215,N_210);
xor U4972 (N_4972,N_1537,N_1181);
xnor U4973 (N_4973,N_1397,N_1778);
and U4974 (N_4974,N_694,N_395);
nand U4975 (N_4975,N_2443,N_1538);
nor U4976 (N_4976,N_1769,N_14);
nor U4977 (N_4977,N_2359,N_551);
or U4978 (N_4978,N_2187,N_1979);
nand U4979 (N_4979,N_1808,N_2255);
or U4980 (N_4980,N_2038,N_1796);
nor U4981 (N_4981,N_858,N_2094);
nand U4982 (N_4982,N_2392,N_2065);
nor U4983 (N_4983,N_771,N_757);
nor U4984 (N_4984,N_509,N_1455);
and U4985 (N_4985,N_2378,N_1118);
and U4986 (N_4986,N_1243,N_389);
xnor U4987 (N_4987,N_2396,N_964);
nor U4988 (N_4988,N_426,N_336);
nor U4989 (N_4989,N_1417,N_48);
or U4990 (N_4990,N_659,N_905);
nand U4991 (N_4991,N_2128,N_570);
and U4992 (N_4992,N_1796,N_1556);
nand U4993 (N_4993,N_827,N_2198);
nand U4994 (N_4994,N_2190,N_861);
or U4995 (N_4995,N_1407,N_437);
nor U4996 (N_4996,N_1974,N_29);
and U4997 (N_4997,N_659,N_1142);
nor U4998 (N_4998,N_2176,N_1605);
and U4999 (N_4999,N_474,N_1410);
nor U5000 (N_5000,N_2675,N_3966);
or U5001 (N_5001,N_3311,N_3965);
or U5002 (N_5002,N_3833,N_3324);
nor U5003 (N_5003,N_4010,N_4987);
nand U5004 (N_5004,N_3782,N_3267);
nor U5005 (N_5005,N_3089,N_3905);
nor U5006 (N_5006,N_3795,N_4089);
nor U5007 (N_5007,N_3422,N_2924);
or U5008 (N_5008,N_4992,N_2953);
or U5009 (N_5009,N_3605,N_2745);
or U5010 (N_5010,N_3657,N_4384);
or U5011 (N_5011,N_2648,N_4977);
nand U5012 (N_5012,N_4473,N_3265);
and U5013 (N_5013,N_4410,N_4158);
nand U5014 (N_5014,N_3395,N_2578);
and U5015 (N_5015,N_4446,N_3524);
nor U5016 (N_5016,N_2714,N_4948);
nand U5017 (N_5017,N_2504,N_4394);
nand U5018 (N_5018,N_3456,N_3356);
nand U5019 (N_5019,N_4487,N_4896);
nor U5020 (N_5020,N_2593,N_3203);
or U5021 (N_5021,N_2758,N_3945);
nor U5022 (N_5022,N_4703,N_3835);
nand U5023 (N_5023,N_4404,N_4940);
nand U5024 (N_5024,N_4579,N_4848);
or U5025 (N_5025,N_4436,N_4715);
nand U5026 (N_5026,N_2694,N_2958);
nor U5027 (N_5027,N_3042,N_4317);
and U5028 (N_5028,N_3298,N_4538);
nand U5029 (N_5029,N_2582,N_3986);
xor U5030 (N_5030,N_4254,N_4248);
and U5031 (N_5031,N_2802,N_3277);
and U5032 (N_5032,N_4002,N_4878);
and U5033 (N_5033,N_4300,N_4998);
or U5034 (N_5034,N_4282,N_4706);
or U5035 (N_5035,N_3704,N_2641);
nand U5036 (N_5036,N_3645,N_3115);
xor U5037 (N_5037,N_4116,N_3116);
and U5038 (N_5038,N_4418,N_2570);
or U5039 (N_5039,N_4834,N_2643);
nand U5040 (N_5040,N_3652,N_2552);
nand U5041 (N_5041,N_3666,N_3280);
nor U5042 (N_5042,N_4079,N_3545);
xnor U5043 (N_5043,N_2742,N_3948);
nand U5044 (N_5044,N_2936,N_2638);
nor U5045 (N_5045,N_4048,N_3838);
nor U5046 (N_5046,N_3473,N_3174);
or U5047 (N_5047,N_2514,N_4947);
and U5048 (N_5048,N_3005,N_3815);
and U5049 (N_5049,N_3175,N_4063);
nand U5050 (N_5050,N_4392,N_2654);
and U5051 (N_5051,N_2910,N_2780);
and U5052 (N_5052,N_4698,N_3253);
nor U5053 (N_5053,N_4680,N_4910);
nand U5054 (N_5054,N_4453,N_2577);
nor U5055 (N_5055,N_2863,N_3332);
and U5056 (N_5056,N_3960,N_4534);
or U5057 (N_5057,N_4731,N_3262);
nand U5058 (N_5058,N_3104,N_4200);
nor U5059 (N_5059,N_3728,N_3114);
nor U5060 (N_5060,N_3228,N_4800);
or U5061 (N_5061,N_3400,N_3740);
or U5062 (N_5062,N_2815,N_4628);
and U5063 (N_5063,N_3940,N_3839);
and U5064 (N_5064,N_3235,N_2972);
or U5065 (N_5065,N_4000,N_3003);
or U5066 (N_5066,N_2679,N_4806);
nand U5067 (N_5067,N_3661,N_2533);
or U5068 (N_5068,N_4799,N_2833);
nand U5069 (N_5069,N_3390,N_3387);
nor U5070 (N_5070,N_3197,N_4169);
and U5071 (N_5071,N_3901,N_3149);
or U5072 (N_5072,N_3367,N_4832);
and U5073 (N_5073,N_3732,N_3669);
and U5074 (N_5074,N_4699,N_4614);
nand U5075 (N_5075,N_2746,N_2683);
or U5076 (N_5076,N_4865,N_4695);
xnor U5077 (N_5077,N_3075,N_2580);
and U5078 (N_5078,N_4576,N_3096);
and U5079 (N_5079,N_4011,N_4841);
or U5080 (N_5080,N_3542,N_3199);
and U5081 (N_5081,N_4221,N_3920);
or U5082 (N_5082,N_3218,N_4636);
or U5083 (N_5083,N_4855,N_4259);
or U5084 (N_5084,N_4052,N_3240);
or U5085 (N_5085,N_4082,N_3073);
or U5086 (N_5086,N_4463,N_3264);
nor U5087 (N_5087,N_4528,N_4790);
nor U5088 (N_5088,N_4488,N_3018);
or U5089 (N_5089,N_4833,N_4922);
or U5090 (N_5090,N_4499,N_4892);
xnor U5091 (N_5091,N_2724,N_3789);
nand U5092 (N_5092,N_2605,N_2986);
nor U5093 (N_5093,N_3339,N_3787);
nand U5094 (N_5094,N_4816,N_4640);
nor U5095 (N_5095,N_4989,N_2741);
and U5096 (N_5096,N_4038,N_4235);
nor U5097 (N_5097,N_2829,N_3580);
nand U5098 (N_5098,N_3259,N_4592);
nand U5099 (N_5099,N_3141,N_2546);
nor U5100 (N_5100,N_4288,N_2860);
nand U5101 (N_5101,N_4648,N_4752);
nor U5102 (N_5102,N_2579,N_4379);
nand U5103 (N_5103,N_3274,N_4134);
nand U5104 (N_5104,N_4125,N_3284);
nor U5105 (N_5105,N_4130,N_4123);
nor U5106 (N_5106,N_3894,N_3281);
nor U5107 (N_5107,N_4323,N_2681);
or U5108 (N_5108,N_4666,N_4007);
and U5109 (N_5109,N_3824,N_4237);
nand U5110 (N_5110,N_2801,N_4168);
nand U5111 (N_5111,N_3204,N_4705);
nand U5112 (N_5112,N_3779,N_3318);
or U5113 (N_5113,N_4189,N_3739);
or U5114 (N_5114,N_3891,N_3967);
nand U5115 (N_5115,N_3762,N_3229);
or U5116 (N_5116,N_3310,N_3291);
nand U5117 (N_5117,N_2647,N_4956);
and U5118 (N_5118,N_3999,N_3238);
or U5119 (N_5119,N_4805,N_4761);
nand U5120 (N_5120,N_3416,N_2673);
nand U5121 (N_5121,N_3518,N_2666);
and U5122 (N_5122,N_4302,N_3727);
and U5123 (N_5123,N_4146,N_3638);
nor U5124 (N_5124,N_4450,N_4490);
or U5125 (N_5125,N_2528,N_2847);
nor U5126 (N_5126,N_4972,N_3609);
or U5127 (N_5127,N_4916,N_3498);
or U5128 (N_5128,N_3119,N_3176);
or U5129 (N_5129,N_2695,N_4313);
nand U5130 (N_5130,N_3436,N_4193);
and U5131 (N_5131,N_3684,N_4433);
nor U5132 (N_5132,N_2555,N_4264);
or U5133 (N_5133,N_4015,N_3407);
and U5134 (N_5134,N_4988,N_3250);
nand U5135 (N_5135,N_4909,N_3292);
nand U5136 (N_5136,N_2769,N_4687);
or U5137 (N_5137,N_2844,N_2717);
nand U5138 (N_5138,N_2917,N_2756);
nor U5139 (N_5139,N_3365,N_2729);
or U5140 (N_5140,N_4380,N_4004);
nand U5141 (N_5141,N_3523,N_2725);
or U5142 (N_5142,N_3817,N_4206);
and U5143 (N_5143,N_2530,N_3826);
and U5144 (N_5144,N_2612,N_3491);
nor U5145 (N_5145,N_3461,N_2968);
xnor U5146 (N_5146,N_3808,N_2545);
nor U5147 (N_5147,N_3670,N_4965);
nand U5148 (N_5148,N_4926,N_4745);
and U5149 (N_5149,N_2915,N_4420);
and U5150 (N_5150,N_4043,N_3696);
nor U5151 (N_5151,N_3923,N_3431);
or U5152 (N_5152,N_4778,N_3985);
nor U5153 (N_5153,N_3006,N_4293);
nand U5154 (N_5154,N_4406,N_2864);
xnor U5155 (N_5155,N_4567,N_3856);
nor U5156 (N_5156,N_2685,N_3269);
nor U5157 (N_5157,N_4262,N_4190);
nor U5158 (N_5158,N_4162,N_2895);
and U5159 (N_5159,N_2786,N_4588);
and U5160 (N_5160,N_4403,N_3536);
nor U5161 (N_5161,N_3226,N_4794);
nand U5162 (N_5162,N_3902,N_2862);
and U5163 (N_5163,N_2825,N_4961);
or U5164 (N_5164,N_2711,N_3889);
nor U5165 (N_5165,N_3792,N_3336);
and U5166 (N_5166,N_3904,N_3709);
or U5167 (N_5167,N_4586,N_4547);
and U5168 (N_5168,N_3012,N_4722);
nor U5169 (N_5169,N_3463,N_2558);
nand U5170 (N_5170,N_4665,N_3056);
nor U5171 (N_5171,N_2800,N_4818);
xor U5172 (N_5172,N_4257,N_4714);
or U5173 (N_5173,N_4960,N_4654);
or U5174 (N_5174,N_4957,N_3359);
nor U5175 (N_5175,N_3034,N_4887);
or U5176 (N_5176,N_4064,N_4740);
and U5177 (N_5177,N_4198,N_2755);
or U5178 (N_5178,N_3830,N_4419);
and U5179 (N_5179,N_4531,N_2976);
nand U5180 (N_5180,N_4398,N_2965);
or U5181 (N_5181,N_3143,N_3713);
nor U5182 (N_5182,N_3681,N_4175);
nand U5183 (N_5183,N_4311,N_4013);
and U5184 (N_5184,N_4827,N_3249);
or U5185 (N_5185,N_3765,N_4732);
or U5186 (N_5186,N_4545,N_3334);
nor U5187 (N_5187,N_2630,N_3363);
and U5188 (N_5188,N_2640,N_2610);
or U5189 (N_5189,N_3750,N_2871);
or U5190 (N_5190,N_3594,N_2840);
nand U5191 (N_5191,N_3969,N_4735);
nor U5192 (N_5192,N_2571,N_3569);
nor U5193 (N_5193,N_4679,N_2626);
or U5194 (N_5194,N_4611,N_3933);
and U5195 (N_5195,N_4859,N_3330);
nor U5196 (N_5196,N_2880,N_3322);
nor U5197 (N_5197,N_3113,N_3273);
and U5198 (N_5198,N_4966,N_3665);
nand U5199 (N_5199,N_4147,N_3256);
or U5200 (N_5200,N_3624,N_2838);
and U5201 (N_5201,N_3044,N_2914);
nor U5202 (N_5202,N_3368,N_3742);
nand U5203 (N_5203,N_2966,N_3266);
nor U5204 (N_5204,N_3471,N_3447);
nand U5205 (N_5205,N_2993,N_2730);
nand U5206 (N_5206,N_4943,N_4181);
nor U5207 (N_5207,N_3233,N_4774);
nand U5208 (N_5208,N_4728,N_3587);
nand U5209 (N_5209,N_3389,N_3152);
or U5210 (N_5210,N_2969,N_3566);
and U5211 (N_5211,N_2875,N_4641);
nor U5212 (N_5212,N_4782,N_3300);
and U5213 (N_5213,N_2807,N_4622);
nand U5214 (N_5214,N_3351,N_3064);
and U5215 (N_5215,N_4102,N_3917);
or U5216 (N_5216,N_3414,N_2553);
or U5217 (N_5217,N_2889,N_3037);
or U5218 (N_5218,N_2913,N_2524);
nand U5219 (N_5219,N_2943,N_3171);
and U5220 (N_5220,N_4271,N_4937);
or U5221 (N_5221,N_2635,N_3065);
and U5222 (N_5222,N_4194,N_3558);
or U5223 (N_5223,N_3192,N_3213);
nand U5224 (N_5224,N_3385,N_4599);
or U5225 (N_5225,N_2908,N_3305);
or U5226 (N_5226,N_2848,N_4577);
and U5227 (N_5227,N_2731,N_4345);
nor U5228 (N_5228,N_4608,N_3121);
nor U5229 (N_5229,N_3499,N_4391);
nor U5230 (N_5230,N_4569,N_4183);
and U5231 (N_5231,N_3470,N_2602);
or U5232 (N_5232,N_2907,N_2866);
nor U5233 (N_5233,N_4165,N_4858);
nand U5234 (N_5234,N_4938,N_2567);
xnor U5235 (N_5235,N_4651,N_2698);
nor U5236 (N_5236,N_4062,N_4029);
xor U5237 (N_5237,N_3148,N_4372);
nor U5238 (N_5238,N_4967,N_4962);
nor U5239 (N_5239,N_3683,N_4712);
nor U5240 (N_5240,N_3754,N_2657);
or U5241 (N_5241,N_3906,N_4906);
or U5242 (N_5242,N_3723,N_4020);
xor U5243 (N_5243,N_3928,N_4016);
nand U5244 (N_5244,N_3489,N_2781);
or U5245 (N_5245,N_3282,N_2589);
nor U5246 (N_5246,N_3829,N_3621);
nand U5247 (N_5247,N_3800,N_3568);
nand U5248 (N_5248,N_3496,N_2700);
and U5249 (N_5249,N_4104,N_2777);
nor U5250 (N_5250,N_3293,N_4124);
nor U5251 (N_5251,N_3607,N_4874);
nor U5252 (N_5252,N_3929,N_4801);
and U5253 (N_5253,N_4990,N_3790);
and U5254 (N_5254,N_4623,N_4811);
nor U5255 (N_5255,N_3032,N_4822);
and U5256 (N_5256,N_3288,N_2854);
and U5257 (N_5257,N_3751,N_3308);
nand U5258 (N_5258,N_4274,N_3874);
nand U5259 (N_5259,N_3136,N_3964);
or U5260 (N_5260,N_4003,N_3153);
nor U5261 (N_5261,N_3352,N_4660);
and U5262 (N_5262,N_2581,N_4253);
or U5263 (N_5263,N_4905,N_4690);
nor U5264 (N_5264,N_3154,N_4039);
xor U5265 (N_5265,N_3842,N_3731);
nor U5266 (N_5266,N_3878,N_3535);
nor U5267 (N_5267,N_3685,N_2554);
xor U5268 (N_5268,N_4122,N_3514);
or U5269 (N_5269,N_3722,N_4145);
nand U5270 (N_5270,N_4797,N_4668);
nor U5271 (N_5271,N_2713,N_2846);
nand U5272 (N_5272,N_3321,N_4074);
xor U5273 (N_5273,N_4857,N_4299);
and U5274 (N_5274,N_4275,N_3797);
nor U5275 (N_5275,N_3459,N_4566);
nand U5276 (N_5276,N_3675,N_4337);
or U5277 (N_5277,N_2834,N_3510);
and U5278 (N_5278,N_3413,N_4771);
nand U5279 (N_5279,N_4709,N_4040);
nor U5280 (N_5280,N_3531,N_2941);
and U5281 (N_5281,N_4223,N_4921);
or U5282 (N_5282,N_2748,N_4746);
or U5283 (N_5283,N_4726,N_4677);
nand U5284 (N_5284,N_3996,N_4484);
and U5285 (N_5285,N_4369,N_2999);
or U5286 (N_5286,N_4443,N_3563);
nor U5287 (N_5287,N_4787,N_4717);
and U5288 (N_5288,N_4034,N_2988);
nand U5289 (N_5289,N_2808,N_3476);
and U5290 (N_5290,N_2945,N_2734);
nand U5291 (N_5291,N_4914,N_3885);
nand U5292 (N_5292,N_4596,N_4355);
nand U5293 (N_5293,N_2620,N_4343);
nor U5294 (N_5294,N_4021,N_2920);
or U5295 (N_5295,N_4086,N_4642);
nor U5296 (N_5296,N_2811,N_3094);
nor U5297 (N_5297,N_4231,N_4869);
nor U5298 (N_5298,N_4424,N_4796);
and U5299 (N_5299,N_3897,N_4574);
or U5300 (N_5300,N_3737,N_3886);
or U5301 (N_5301,N_2515,N_4481);
and U5302 (N_5302,N_3306,N_2899);
nand U5303 (N_5303,N_3590,N_4144);
and U5304 (N_5304,N_3865,N_2709);
nor U5305 (N_5305,N_4090,N_3887);
nand U5306 (N_5306,N_2989,N_4851);
nor U5307 (N_5307,N_3578,N_2697);
nor U5308 (N_5308,N_2559,N_4336);
nor U5309 (N_5309,N_3924,N_3430);
nand U5310 (N_5310,N_4936,N_2573);
nand U5311 (N_5311,N_3483,N_4526);
nor U5312 (N_5312,N_2703,N_4776);
or U5313 (N_5313,N_4808,N_4121);
or U5314 (N_5314,N_3658,N_4024);
or U5315 (N_5315,N_4929,N_2561);
or U5316 (N_5316,N_3736,N_2728);
nor U5317 (N_5317,N_2757,N_3527);
and U5318 (N_5318,N_2521,N_2896);
or U5319 (N_5319,N_3757,N_2601);
or U5320 (N_5320,N_4456,N_3650);
and U5321 (N_5321,N_2557,N_2835);
nor U5322 (N_5322,N_3724,N_4069);
and U5323 (N_5323,N_3392,N_3972);
or U5324 (N_5324,N_3170,N_3606);
and U5325 (N_5325,N_2609,N_3761);
nand U5326 (N_5326,N_3118,N_4432);
and U5327 (N_5327,N_3002,N_2534);
or U5328 (N_5328,N_4114,N_2735);
or U5329 (N_5329,N_2978,N_2625);
nor U5330 (N_5330,N_4205,N_4331);
nand U5331 (N_5331,N_3433,N_4441);
or U5332 (N_5332,N_4285,N_3268);
nand U5333 (N_5333,N_4460,N_3890);
and U5334 (N_5334,N_2591,N_4843);
or U5335 (N_5335,N_4904,N_4495);
and U5336 (N_5336,N_2588,N_3555);
and U5337 (N_5337,N_3180,N_4604);
or U5338 (N_5338,N_4327,N_4764);
or U5339 (N_5339,N_4609,N_4126);
and U5340 (N_5340,N_3564,N_3185);
nand U5341 (N_5341,N_4058,N_2776);
nand U5342 (N_5342,N_3981,N_4475);
or U5343 (N_5343,N_3221,N_4105);
nand U5344 (N_5344,N_3596,N_4733);
and U5345 (N_5345,N_3690,N_4558);
or U5346 (N_5346,N_4414,N_2510);
and U5347 (N_5347,N_3467,N_2812);
nand U5348 (N_5348,N_2932,N_2660);
and U5349 (N_5349,N_2738,N_4692);
nor U5350 (N_5350,N_4304,N_4853);
nor U5351 (N_5351,N_4543,N_4523);
nand U5352 (N_5352,N_3111,N_4281);
or U5353 (N_5353,N_3546,N_4359);
nand U5354 (N_5354,N_3576,N_3384);
and U5355 (N_5355,N_3845,N_2996);
nor U5356 (N_5356,N_4365,N_3488);
nand U5357 (N_5357,N_3957,N_3343);
and U5358 (N_5358,N_3921,N_4741);
or U5359 (N_5359,N_3011,N_3067);
nor U5360 (N_5360,N_2526,N_4627);
and U5361 (N_5361,N_4584,N_3529);
or U5362 (N_5362,N_4445,N_2865);
or U5363 (N_5363,N_4153,N_4128);
or U5364 (N_5364,N_4537,N_2661);
or U5365 (N_5365,N_3828,N_4397);
nor U5366 (N_5366,N_4232,N_2970);
and U5367 (N_5367,N_4867,N_3585);
and U5368 (N_5368,N_2940,N_2990);
nor U5369 (N_5369,N_3066,N_4141);
or U5370 (N_5370,N_3438,N_3644);
nand U5371 (N_5371,N_4358,N_3078);
or U5372 (N_5372,N_3123,N_2634);
and U5373 (N_5373,N_3107,N_3954);
nor U5374 (N_5374,N_2505,N_3278);
or U5375 (N_5375,N_4767,N_4664);
xnor U5376 (N_5376,N_4439,N_2923);
nand U5377 (N_5377,N_2704,N_2981);
nor U5378 (N_5378,N_4115,N_4291);
nor U5379 (N_5379,N_3486,N_2951);
nor U5380 (N_5380,N_2549,N_2674);
nand U5381 (N_5381,N_2655,N_3870);
and U5382 (N_5382,N_4497,N_3809);
nor U5383 (N_5383,N_4132,N_2747);
nor U5384 (N_5384,N_4001,N_2686);
nand U5385 (N_5385,N_4829,N_4066);
or U5386 (N_5386,N_3677,N_4825);
nor U5387 (N_5387,N_4322,N_3102);
and U5388 (N_5388,N_4762,N_4713);
or U5389 (N_5389,N_3445,N_2952);
and U5390 (N_5390,N_2985,N_4549);
or U5391 (N_5391,N_3883,N_3653);
or U5392 (N_5392,N_2839,N_4129);
and U5393 (N_5393,N_2931,N_2982);
nor U5394 (N_5394,N_4846,N_3942);
nand U5395 (N_5395,N_3232,N_4277);
nor U5396 (N_5396,N_4051,N_3858);
nor U5397 (N_5397,N_4505,N_3840);
nand U5398 (N_5398,N_3798,N_3768);
nor U5399 (N_5399,N_4603,N_3793);
and U5400 (N_5400,N_2603,N_3156);
and U5401 (N_5401,N_4477,N_3021);
or U5402 (N_5402,N_4760,N_2699);
and U5403 (N_5403,N_3866,N_3248);
nor U5404 (N_5404,N_3697,N_4172);
nand U5405 (N_5405,N_2633,N_3245);
and U5406 (N_5406,N_3349,N_3210);
and U5407 (N_5407,N_3672,N_3358);
and U5408 (N_5408,N_4793,N_4585);
nand U5409 (N_5409,N_4081,N_4097);
nor U5410 (N_5410,N_3918,N_3725);
nor U5411 (N_5411,N_4875,N_4931);
and U5412 (N_5412,N_3820,N_4511);
and U5413 (N_5413,N_4440,N_3786);
nand U5414 (N_5414,N_2964,N_2785);
xnor U5415 (N_5415,N_4602,N_4435);
or U5416 (N_5416,N_3922,N_3296);
and U5417 (N_5417,N_4017,N_2876);
nor U5418 (N_5418,N_4199,N_4215);
and U5419 (N_5419,N_3884,N_4661);
and U5420 (N_5420,N_3907,N_2543);
and U5421 (N_5421,N_2874,N_4891);
nor U5422 (N_5422,N_3164,N_4521);
and U5423 (N_5423,N_3505,N_2538);
or U5424 (N_5424,N_2664,N_3515);
or U5425 (N_5425,N_4583,N_3004);
nor U5426 (N_5426,N_4233,N_4898);
nand U5427 (N_5427,N_3374,N_4512);
nor U5428 (N_5428,N_4425,N_3926);
or U5429 (N_5429,N_4630,N_3643);
nand U5430 (N_5430,N_4777,N_3286);
nand U5431 (N_5431,N_2656,N_4492);
nand U5432 (N_5432,N_3843,N_4245);
and U5433 (N_5433,N_2548,N_3756);
or U5434 (N_5434,N_3013,N_4480);
and U5435 (N_5435,N_4634,N_3770);
or U5436 (N_5436,N_3202,N_4619);
and U5437 (N_5437,N_4214,N_4057);
xor U5438 (N_5438,N_3272,N_2564);
nor U5439 (N_5439,N_3802,N_2797);
nor U5440 (N_5440,N_3752,N_4170);
and U5441 (N_5441,N_2754,N_4830);
or U5442 (N_5442,N_3468,N_3200);
and U5443 (N_5443,N_2733,N_3181);
or U5444 (N_5444,N_3452,N_3772);
and U5445 (N_5445,N_4164,N_4580);
nor U5446 (N_5446,N_2706,N_4516);
nand U5447 (N_5447,N_4278,N_4854);
or U5448 (N_5448,N_3335,N_3693);
nor U5449 (N_5449,N_3521,N_4758);
nand U5450 (N_5450,N_3196,N_4819);
nor U5451 (N_5451,N_3589,N_4542);
nand U5452 (N_5452,N_3397,N_3541);
and U5453 (N_5453,N_3773,N_4889);
and U5454 (N_5454,N_4894,N_4031);
nand U5455 (N_5455,N_3297,N_4996);
nor U5456 (N_5456,N_3453,N_3959);
nor U5457 (N_5457,N_4489,N_3909);
or U5458 (N_5458,N_3612,N_4030);
or U5459 (N_5459,N_2677,N_4689);
nand U5460 (N_5460,N_4325,N_4736);
and U5461 (N_5461,N_3161,N_4621);
nand U5462 (N_5462,N_4230,N_2520);
and U5463 (N_5463,N_2804,N_2819);
or U5464 (N_5464,N_2627,N_4286);
nor U5465 (N_5465,N_4416,N_4649);
nor U5466 (N_5466,N_3630,N_2960);
xnor U5467 (N_5467,N_4561,N_3822);
nor U5468 (N_5468,N_3699,N_4658);
and U5469 (N_5469,N_3361,N_3711);
nor U5470 (N_5470,N_3565,N_3207);
nor U5471 (N_5471,N_3425,N_4994);
or U5472 (N_5472,N_4338,N_3559);
nand U5473 (N_5473,N_3216,N_3913);
nor U5474 (N_5474,N_3544,N_4532);
nor U5475 (N_5475,N_4842,N_4785);
or U5476 (N_5476,N_2692,N_4856);
and U5477 (N_5477,N_3759,N_3494);
or U5478 (N_5478,N_2764,N_3026);
and U5479 (N_5479,N_3507,N_4303);
and U5480 (N_5480,N_3561,N_4407);
or U5481 (N_5481,N_4701,N_3504);
or U5482 (N_5482,N_4789,N_4527);
nor U5483 (N_5483,N_3127,N_3304);
nor U5484 (N_5484,N_3968,N_4902);
and U5485 (N_5485,N_2766,N_4413);
nand U5486 (N_5486,N_3420,N_4171);
and U5487 (N_5487,N_3777,N_3070);
nand U5488 (N_5488,N_4804,N_3816);
and U5489 (N_5489,N_3410,N_2830);
and U5490 (N_5490,N_4401,N_2619);
nor U5491 (N_5491,N_4329,N_4018);
and U5492 (N_5492,N_4837,N_4376);
or U5493 (N_5493,N_3910,N_4650);
or U5494 (N_5494,N_2743,N_2737);
and U5495 (N_5495,N_4249,N_4362);
nand U5496 (N_5496,N_2539,N_2905);
nand U5497 (N_5497,N_3105,N_4256);
or U5498 (N_5498,N_3317,N_3059);
and U5499 (N_5499,N_3547,N_3939);
xnor U5500 (N_5500,N_4136,N_3855);
and U5501 (N_5501,N_3602,N_3600);
nor U5502 (N_5502,N_4786,N_3846);
nand U5503 (N_5503,N_4562,N_4041);
nor U5504 (N_5504,N_2859,N_3774);
nand U5505 (N_5505,N_4888,N_3454);
or U5506 (N_5506,N_4341,N_4781);
and U5507 (N_5507,N_4659,N_4110);
nand U5508 (N_5508,N_3687,N_4451);
or U5509 (N_5509,N_3329,N_3001);
or U5510 (N_5510,N_3698,N_4192);
and U5511 (N_5511,N_4975,N_3502);
and U5512 (N_5512,N_4119,N_2678);
nor U5513 (N_5513,N_3497,N_2716);
nor U5514 (N_5514,N_3319,N_3859);
or U5515 (N_5515,N_3487,N_3978);
nand U5516 (N_5516,N_2616,N_2551);
nand U5517 (N_5517,N_2935,N_3464);
and U5518 (N_5518,N_3344,N_3144);
or U5519 (N_5519,N_4087,N_4222);
and U5520 (N_5520,N_3071,N_2994);
and U5521 (N_5521,N_3584,N_3314);
and U5522 (N_5522,N_4616,N_3208);
nand U5523 (N_5523,N_3412,N_2722);
nor U5524 (N_5524,N_4765,N_3261);
and U5525 (N_5525,N_4470,N_3925);
nor U5526 (N_5526,N_2667,N_3571);
nor U5527 (N_5527,N_4072,N_4980);
or U5528 (N_5528,N_4635,N_4838);
and U5529 (N_5529,N_3983,N_4217);
and U5530 (N_5530,N_2849,N_2826);
or U5531 (N_5531,N_2791,N_3540);
nand U5532 (N_5532,N_4201,N_3328);
and U5533 (N_5533,N_4873,N_4840);
nor U5534 (N_5534,N_2921,N_4606);
and U5535 (N_5535,N_3912,N_4113);
and U5536 (N_5536,N_4522,N_2799);
nor U5537 (N_5537,N_2942,N_3603);
and U5538 (N_5538,N_4035,N_3429);
and U5539 (N_5539,N_4226,N_4952);
nor U5540 (N_5540,N_3028,N_3610);
or U5541 (N_5541,N_3206,N_3130);
and U5542 (N_5542,N_3159,N_2901);
or U5543 (N_5543,N_3396,N_3376);
nor U5544 (N_5544,N_3027,N_4252);
nand U5545 (N_5545,N_3382,N_4788);
nor U5546 (N_5546,N_3475,N_3231);
xnor U5547 (N_5547,N_3108,N_4080);
nand U5548 (N_5548,N_3689,N_3557);
or U5549 (N_5549,N_2689,N_2934);
and U5550 (N_5550,N_3092,N_4483);
or U5551 (N_5551,N_3029,N_2947);
nor U5552 (N_5552,N_2869,N_2712);
nor U5553 (N_5553,N_4180,N_4519);
nor U5554 (N_5554,N_2597,N_4229);
or U5555 (N_5555,N_4494,N_4678);
or U5556 (N_5556,N_2512,N_2832);
nor U5557 (N_5557,N_3806,N_3146);
nor U5558 (N_5558,N_4191,N_3348);
or U5559 (N_5559,N_2740,N_3236);
nand U5560 (N_5560,N_4060,N_3799);
nor U5561 (N_5561,N_3827,N_2984);
nand U5562 (N_5562,N_4437,N_3758);
or U5563 (N_5563,N_3850,N_4389);
or U5564 (N_5564,N_2618,N_3533);
nor U5565 (N_5565,N_4321,N_4117);
and U5566 (N_5566,N_3893,N_2763);
or U5567 (N_5567,N_2658,N_3484);
nand U5568 (N_5568,N_2645,N_3719);
and U5569 (N_5569,N_4356,N_2852);
or U5570 (N_5570,N_4022,N_4766);
or U5571 (N_5571,N_3117,N_4294);
and U5572 (N_5572,N_3631,N_3109);
nor U5573 (N_5573,N_2691,N_3528);
and U5574 (N_5574,N_3807,N_4517);
and U5575 (N_5575,N_2979,N_4218);
nand U5576 (N_5576,N_2540,N_4729);
nand U5577 (N_5577,N_2767,N_3030);
nor U5578 (N_5578,N_2576,N_4187);
nor U5579 (N_5579,N_2639,N_3312);
nor U5580 (N_5580,N_2946,N_4400);
nor U5581 (N_5581,N_4696,N_3419);
nand U5582 (N_5582,N_4978,N_2621);
nor U5583 (N_5583,N_2884,N_4601);
nand U5584 (N_5584,N_2980,N_2547);
and U5585 (N_5585,N_3285,N_4826);
or U5586 (N_5586,N_4913,N_4831);
nand U5587 (N_5587,N_4067,N_2696);
nand U5588 (N_5588,N_3898,N_4143);
or U5589 (N_5589,N_2765,N_4240);
and U5590 (N_5590,N_2853,N_3099);
or U5591 (N_5591,N_2822,N_4861);
or U5592 (N_5592,N_2987,N_3963);
nand U5593 (N_5593,N_2890,N_2710);
nand U5594 (N_5594,N_4287,N_3482);
and U5595 (N_5595,N_3183,N_3357);
or U5596 (N_5596,N_3251,N_3962);
or U5597 (N_5597,N_4685,N_4711);
or U5598 (N_5598,N_3949,N_4928);
or U5599 (N_5599,N_4959,N_3217);
or U5600 (N_5600,N_3140,N_3593);
and U5601 (N_5601,N_3646,N_2944);
or U5602 (N_5602,N_4693,N_4319);
or U5603 (N_5603,N_3485,N_4348);
nor U5604 (N_5604,N_4638,N_3294);
nand U5605 (N_5605,N_2671,N_2750);
nor U5606 (N_5606,N_2806,N_4065);
nor U5607 (N_5607,N_3791,N_3526);
or U5608 (N_5608,N_3069,N_2649);
nand U5609 (N_5609,N_4417,N_3147);
and U5610 (N_5610,N_3873,N_3863);
and U5611 (N_5611,N_3053,N_4265);
or U5612 (N_5612,N_3193,N_3342);
nand U5613 (N_5613,N_3686,N_4342);
or U5614 (N_5614,N_4652,N_3313);
nor U5615 (N_5615,N_4054,N_4587);
nand U5616 (N_5616,N_2752,N_3391);
nor U5617 (N_5617,N_4590,N_3090);
nor U5618 (N_5618,N_3745,N_3511);
nor U5619 (N_5619,N_3142,N_4893);
and U5620 (N_5620,N_2550,N_2778);
nor U5621 (N_5621,N_2855,N_3637);
and U5622 (N_5622,N_4591,N_3375);
nand U5623 (N_5623,N_2501,N_3573);
nor U5624 (N_5624,N_3241,N_4320);
nand U5625 (N_5625,N_3706,N_2744);
or U5626 (N_5626,N_3998,N_4812);
or U5627 (N_5627,N_4280,N_4775);
and U5628 (N_5628,N_3493,N_3834);
or U5629 (N_5629,N_3916,N_3371);
nand U5630 (N_5630,N_2774,N_3260);
or U5631 (N_5631,N_4814,N_3441);
or U5632 (N_5632,N_2615,N_3747);
nor U5633 (N_5633,N_2739,N_4371);
nor U5634 (N_5634,N_3674,N_4033);
nor U5635 (N_5635,N_4431,N_4173);
and U5636 (N_5636,N_4077,N_4346);
and U5637 (N_5637,N_4408,N_3879);
or U5638 (N_5638,N_4385,N_3301);
or U5639 (N_5639,N_3340,N_3326);
or U5640 (N_5640,N_4255,N_4289);
or U5641 (N_5641,N_4155,N_3562);
or U5642 (N_5642,N_4915,N_3553);
and U5643 (N_5643,N_4268,N_4298);
nor U5644 (N_5644,N_2954,N_4618);
or U5645 (N_5645,N_4672,N_4879);
xnor U5646 (N_5646,N_3423,N_3333);
or U5647 (N_5647,N_4099,N_4605);
nand U5648 (N_5648,N_3679,N_3844);
and U5649 (N_5649,N_4377,N_3618);
or U5650 (N_5650,N_3854,N_2705);
or U5651 (N_5651,N_3591,N_4780);
nand U5652 (N_5652,N_4997,N_3642);
or U5653 (N_5653,N_3853,N_3355);
or U5654 (N_5654,N_3896,N_3055);
or U5655 (N_5655,N_3081,N_3805);
or U5656 (N_5656,N_2687,N_3673);
or U5657 (N_5657,N_3492,N_3950);
nor U5658 (N_5658,N_4986,N_4349);
or U5659 (N_5659,N_4620,N_4340);
nor U5660 (N_5660,N_4589,N_3796);
nor U5661 (N_5661,N_4629,N_2600);
and U5662 (N_5662,N_2544,N_3263);
nor U5663 (N_5663,N_2587,N_2701);
nor U5664 (N_5664,N_3379,N_2795);
nor U5665 (N_5665,N_3195,N_4228);
and U5666 (N_5666,N_2693,N_3307);
nand U5667 (N_5667,N_2828,N_4290);
or U5668 (N_5668,N_4159,N_2967);
and U5669 (N_5669,N_4491,N_3364);
or U5670 (N_5670,N_4935,N_2841);
nor U5671 (N_5671,N_4045,N_3520);
nor U5672 (N_5672,N_3088,N_4421);
nand U5673 (N_5673,N_4798,N_4813);
nor U5674 (N_5674,N_3597,N_3861);
or U5675 (N_5675,N_2637,N_4088);
and U5676 (N_5676,N_3287,N_4267);
and U5677 (N_5677,N_4510,N_4412);
or U5678 (N_5678,N_2642,N_4598);
and U5679 (N_5679,N_4912,N_4220);
or U5680 (N_5680,N_3785,N_4565);
or U5681 (N_5681,N_4556,N_4507);
nor U5682 (N_5682,N_3474,N_2569);
nor U5683 (N_5683,N_4269,N_4820);
nand U5684 (N_5684,N_2665,N_4925);
nand U5685 (N_5685,N_3583,N_3781);
and U5686 (N_5686,N_4791,N_4261);
nor U5687 (N_5687,N_3575,N_2973);
nor U5688 (N_5688,N_4684,N_3680);
nor U5689 (N_5689,N_3574,N_4266);
nand U5690 (N_5690,N_3350,N_2753);
nor U5691 (N_5691,N_4546,N_3072);
nor U5692 (N_5692,N_3988,N_4127);
nand U5693 (N_5693,N_3191,N_3393);
or U5694 (N_5694,N_3106,N_4920);
and U5695 (N_5695,N_3095,N_3215);
nor U5696 (N_5696,N_2670,N_4946);
nand U5697 (N_5697,N_4457,N_3439);
or U5698 (N_5698,N_4673,N_3255);
nor U5699 (N_5699,N_4409,N_4381);
and U5700 (N_5700,N_3951,N_4390);
nand U5701 (N_5701,N_4387,N_4347);
and U5702 (N_5702,N_4106,N_4708);
or U5703 (N_5703,N_2909,N_2805);
and U5704 (N_5704,N_4933,N_3039);
nor U5705 (N_5705,N_3316,N_3864);
and U5706 (N_5706,N_3060,N_4704);
or U5707 (N_5707,N_4759,N_3290);
and U5708 (N_5708,N_3270,N_4263);
nand U5709 (N_5709,N_2891,N_4817);
or U5710 (N_5710,N_4028,N_3415);
and U5711 (N_5711,N_3362,N_3876);
nand U5712 (N_5712,N_3458,N_3162);
nand U5713 (N_5713,N_4503,N_3599);
and U5714 (N_5714,N_2595,N_3479);
and U5715 (N_5715,N_2636,N_4092);
nor U5716 (N_5716,N_3977,N_3151);
nor U5717 (N_5717,N_3676,N_3303);
nor U5718 (N_5718,N_4328,N_3579);
nor U5719 (N_5719,N_3936,N_4241);
and U5720 (N_5720,N_4139,N_4493);
nand U5721 (N_5721,N_2837,N_2502);
and U5722 (N_5722,N_4836,N_2608);
nand U5723 (N_5723,N_4768,N_4135);
and U5724 (N_5724,N_4163,N_4496);
and U5725 (N_5725,N_4046,N_3662);
or U5726 (N_5726,N_3513,N_3744);
nand U5727 (N_5727,N_3506,N_2991);
nand U5728 (N_5728,N_3048,N_3615);
or U5729 (N_5729,N_4844,N_2933);
nand U5730 (N_5730,N_2784,N_3778);
nand U5731 (N_5731,N_3299,N_4472);
and U5732 (N_5732,N_4881,N_4167);
and U5733 (N_5733,N_4670,N_3862);
or U5734 (N_5734,N_4179,N_3167);
nand U5735 (N_5735,N_3372,N_4008);
nor U5736 (N_5736,N_3046,N_2894);
nand U5737 (N_5737,N_2584,N_2883);
and U5738 (N_5738,N_3900,N_4009);
xnor U5739 (N_5739,N_2529,N_3279);
nand U5740 (N_5740,N_3648,N_3619);
and U5741 (N_5741,N_4908,N_4131);
or U5742 (N_5742,N_2974,N_4025);
nor U5743 (N_5743,N_3077,N_4973);
nor U5744 (N_5744,N_4032,N_3227);
and U5745 (N_5745,N_4430,N_3688);
xnor U5746 (N_5746,N_2813,N_2749);
nor U5747 (N_5747,N_3080,N_2937);
nand U5748 (N_5748,N_4530,N_4663);
nor U5749 (N_5749,N_2598,N_3179);
or U5750 (N_5750,N_3132,N_3083);
and U5751 (N_5751,N_3911,N_2903);
nand U5752 (N_5752,N_2817,N_2782);
or U5753 (N_5753,N_3813,N_2518);
and U5754 (N_5754,N_3427,N_4501);
nor U5755 (N_5755,N_3577,N_3254);
or U5756 (N_5756,N_4753,N_4570);
and U5757 (N_5757,N_3956,N_3038);
nand U5758 (N_5758,N_3009,N_4750);
and U5759 (N_5759,N_2503,N_4529);
nor U5760 (N_5760,N_4197,N_3712);
nor U5761 (N_5761,N_3710,N_4626);
nor U5762 (N_5762,N_4272,N_4444);
or U5763 (N_5763,N_2736,N_4184);
nor U5764 (N_5764,N_3769,N_4118);
nor U5765 (N_5765,N_2594,N_3000);
and U5766 (N_5766,N_3720,N_4950);
or U5767 (N_5767,N_4949,N_2508);
or U5768 (N_5768,N_4027,N_2881);
xor U5769 (N_5769,N_4968,N_4541);
nand U5770 (N_5770,N_4378,N_4610);
xor U5771 (N_5771,N_2922,N_3804);
or U5772 (N_5772,N_3554,N_3927);
nand U5773 (N_5773,N_3692,N_3225);
and U5774 (N_5774,N_3440,N_3025);
nor U5775 (N_5775,N_2949,N_4724);
or U5776 (N_5776,N_2506,N_4559);
nand U5777 (N_5777,N_3997,N_3128);
nand U5778 (N_5778,N_3446,N_3442);
or U5779 (N_5779,N_3360,N_3377);
nor U5780 (N_5780,N_4075,N_2898);
nor U5781 (N_5781,N_2719,N_3801);
nand U5782 (N_5782,N_3047,N_3150);
and U5783 (N_5783,N_2676,N_2575);
nor U5784 (N_5784,N_3755,N_4983);
or U5785 (N_5785,N_4743,N_4447);
or U5786 (N_5786,N_2599,N_3703);
nor U5787 (N_5787,N_3320,N_4270);
nand U5788 (N_5788,N_4415,N_3495);
and U5789 (N_5789,N_3771,N_3871);
nor U5790 (N_5790,N_4876,N_2888);
nor U5791 (N_5791,N_4455,N_4644);
and U5792 (N_5792,N_4907,N_2983);
and U5793 (N_5793,N_2715,N_3641);
and U5794 (N_5794,N_4563,N_3640);
and U5795 (N_5795,N_3930,N_4395);
nor U5796 (N_5796,N_4981,N_4945);
nand U5797 (N_5797,N_4615,N_2542);
and U5798 (N_5798,N_3819,N_3139);
nand U5799 (N_5799,N_3984,N_2566);
nor U5800 (N_5800,N_4754,N_4656);
and U5801 (N_5801,N_4279,N_4485);
or U5802 (N_5802,N_4737,N_2622);
nor U5803 (N_5803,N_3068,N_4779);
nand U5804 (N_5804,N_4366,N_4464);
and U5805 (N_5805,N_3500,N_3671);
nand U5806 (N_5806,N_3378,N_3198);
or U5807 (N_5807,N_2930,N_2523);
or U5808 (N_5808,N_2867,N_3629);
or U5809 (N_5809,N_3509,N_3743);
nor U5810 (N_5810,N_4296,N_3915);
nand U5811 (N_5811,N_3346,N_3417);
and U5812 (N_5812,N_3784,N_4382);
xor U5813 (N_5813,N_4195,N_2861);
nor U5814 (N_5814,N_3007,N_3058);
nor U5815 (N_5815,N_4258,N_2583);
or U5816 (N_5816,N_2879,N_4633);
nand U5817 (N_5817,N_4095,N_3223);
or U5818 (N_5818,N_3126,N_2651);
or U5819 (N_5819,N_3045,N_3230);
and U5820 (N_5820,N_3639,N_3895);
nand U5821 (N_5821,N_4308,N_4339);
nand U5822 (N_5822,N_2793,N_3783);
and U5823 (N_5823,N_2892,N_3098);
nor U5824 (N_5824,N_2886,N_3821);
nand U5825 (N_5825,N_3381,N_4595);
and U5826 (N_5826,N_2770,N_3408);
nor U5827 (N_5827,N_2537,N_3354);
or U5828 (N_5828,N_3803,N_3832);
nand U5829 (N_5829,N_3714,N_3194);
and U5830 (N_5830,N_2720,N_3938);
nand U5831 (N_5831,N_2760,N_3655);
or U5832 (N_5832,N_3383,N_4984);
nand U5833 (N_5833,N_4204,N_4236);
nand U5834 (N_5834,N_2928,N_2507);
and U5835 (N_5835,N_3222,N_4655);
nand U5836 (N_5836,N_3608,N_4225);
or U5837 (N_5837,N_3271,N_3812);
and U5838 (N_5838,N_4763,N_4312);
nand U5839 (N_5839,N_2682,N_3974);
nor U5840 (N_5840,N_2690,N_3405);
nand U5841 (N_5841,N_2851,N_3177);
nand U5842 (N_5842,N_3444,N_3426);
or U5843 (N_5843,N_4895,N_4744);
or U5844 (N_5844,N_4903,N_2798);
and U5845 (N_5845,N_4890,N_2590);
nor U5846 (N_5846,N_3120,N_4725);
and U5847 (N_5847,N_3401,N_2885);
or U5848 (N_5848,N_4053,N_4196);
or U5849 (N_5849,N_2631,N_4211);
nor U5850 (N_5850,N_4361,N_3169);
nand U5851 (N_5851,N_3214,N_4107);
nand U5852 (N_5852,N_4388,N_4963);
and U5853 (N_5853,N_4352,N_4094);
or U5854 (N_5854,N_4955,N_3700);
and U5855 (N_5855,N_4056,N_4970);
or U5856 (N_5856,N_3869,N_3668);
or U5857 (N_5857,N_4239,N_2857);
nor U5858 (N_5858,N_4373,N_3825);
and U5859 (N_5859,N_3212,N_3851);
or U5860 (N_5860,N_4669,N_4213);
and U5861 (N_5861,N_4682,N_4770);
and U5862 (N_5862,N_3570,N_2702);
and U5863 (N_5863,N_3131,N_3289);
nor U5864 (N_5864,N_4076,N_3478);
or U5865 (N_5865,N_4930,N_4544);
and U5866 (N_5866,N_4486,N_4405);
or U5867 (N_5867,N_3187,N_2592);
nor U5868 (N_5868,N_4207,N_3057);
nand U5869 (N_5869,N_4284,N_4368);
and U5870 (N_5870,N_2820,N_3325);
or U5871 (N_5871,N_3403,N_3353);
or U5872 (N_5872,N_3852,N_3539);
or U5873 (N_5873,N_3469,N_3110);
nor U5874 (N_5874,N_3729,N_3020);
and U5875 (N_5875,N_3490,N_3211);
xor U5876 (N_5876,N_3041,N_4462);
xnor U5877 (N_5877,N_4216,N_3122);
nand U5878 (N_5878,N_2522,N_3209);
nor U5879 (N_5879,N_3625,N_4700);
nand U5880 (N_5880,N_4012,N_2975);
nand U5881 (N_5881,N_2632,N_3450);
nand U5882 (N_5882,N_2995,N_4005);
or U5883 (N_5883,N_3257,N_2516);
nor U5884 (N_5884,N_3934,N_2831);
nand U5885 (N_5885,N_4784,N_4548);
nor U5886 (N_5886,N_4260,N_4307);
and U5887 (N_5887,N_4112,N_3847);
and U5888 (N_5888,N_3182,N_4474);
or U5889 (N_5889,N_3386,N_3388);
or U5890 (N_5890,N_4749,N_4314);
nor U5891 (N_5891,N_4354,N_2527);
nor U5892 (N_5892,N_2997,N_4514);
and U5893 (N_5893,N_3788,N_2873);
or U5894 (N_5894,N_3188,N_4646);
and U5895 (N_5895,N_3031,N_3552);
nand U5896 (N_5896,N_3649,N_4810);
and U5897 (N_5897,N_4442,N_2868);
and U5898 (N_5898,N_4539,N_3976);
and U5899 (N_5899,N_2836,N_4234);
nand U5900 (N_5900,N_3867,N_3015);
nor U5901 (N_5901,N_4674,N_4178);
or U5902 (N_5902,N_4295,N_3434);
nor U5903 (N_5903,N_2653,N_2565);
nand U5904 (N_5904,N_4862,N_4632);
and U5905 (N_5905,N_4671,N_2624);
and U5906 (N_5906,N_3345,N_3881);
nand U5907 (N_5907,N_4802,N_2663);
or U5908 (N_5908,N_3971,N_3244);
and U5909 (N_5909,N_4720,N_3085);
and U5910 (N_5910,N_4884,N_3748);
xor U5911 (N_5911,N_3097,N_3309);
and U5912 (N_5912,N_3955,N_3626);
nand U5913 (N_5913,N_4324,N_2536);
nand U5914 (N_5914,N_4718,N_4305);
and U5915 (N_5915,N_3472,N_3008);
nand U5916 (N_5916,N_3993,N_3746);
nand U5917 (N_5917,N_3550,N_3455);
nor U5918 (N_5918,N_3480,N_4186);
nor U5919 (N_5919,N_3708,N_4828);
or U5920 (N_5920,N_3764,N_2525);
nor U5921 (N_5921,N_3428,N_2768);
nand U5922 (N_5922,N_3663,N_3205);
or U5923 (N_5923,N_4919,N_3947);
and U5924 (N_5924,N_3810,N_4969);
or U5925 (N_5925,N_3160,N_4871);
and U5926 (N_5926,N_2721,N_3158);
nand U5927 (N_5927,N_2659,N_3219);
and U5928 (N_5928,N_2916,N_3172);
nand U5929 (N_5929,N_3022,N_4399);
nor U5930 (N_5930,N_4551,N_3477);
nor U5931 (N_5931,N_3234,N_3994);
xnor U5932 (N_5932,N_4219,N_4557);
and U5933 (N_5933,N_3741,N_4974);
and U5934 (N_5934,N_2971,N_4653);
nand U5935 (N_5935,N_4212,N_4924);
and U5936 (N_5936,N_3888,N_3937);
or U5937 (N_5937,N_4571,N_4509);
and U5938 (N_5938,N_3138,N_3133);
nand U5939 (N_5939,N_4852,N_4686);
nand U5940 (N_5940,N_3707,N_4091);
and U5941 (N_5941,N_2906,N_3163);
nor U5942 (N_5942,N_3660,N_2672);
nand U5943 (N_5943,N_4850,N_2560);
or U5944 (N_5944,N_2856,N_3437);
nor U5945 (N_5945,N_3567,N_3165);
or U5946 (N_5946,N_3243,N_4927);
xor U5947 (N_5947,N_2794,N_2959);
or U5948 (N_5948,N_3598,N_4823);
or U5949 (N_5949,N_3016,N_4166);
nor U5950 (N_5950,N_4049,N_2628);
xor U5951 (N_5951,N_4953,N_3462);
or U5952 (N_5952,N_2893,N_4839);
nand U5953 (N_5953,N_4506,N_3035);
or U5954 (N_5954,N_4471,N_4647);
nor U5955 (N_5955,N_3054,N_4364);
and U5956 (N_5956,N_3370,N_4964);
nand U5957 (N_5957,N_2918,N_3033);
nor U5958 (N_5958,N_3448,N_4883);
or U5959 (N_5959,N_2821,N_3076);
nor U5960 (N_5960,N_4553,N_4533);
nor U5961 (N_5961,N_3775,N_4594);
and U5962 (N_5962,N_3811,N_4150);
nand U5963 (N_5963,N_4897,N_4821);
and U5964 (N_5964,N_4939,N_4513);
and U5965 (N_5965,N_4730,N_3019);
nand U5966 (N_5966,N_4694,N_4564);
nand U5967 (N_5967,N_2732,N_3394);
nor U5968 (N_5968,N_3135,N_2668);
nor U5969 (N_5969,N_4315,N_3220);
or U5970 (N_5970,N_4108,N_3620);
or U5971 (N_5971,N_4176,N_4148);
or U5972 (N_5972,N_3242,N_4133);
and U5973 (N_5973,N_2708,N_4036);
nand U5974 (N_5974,N_2511,N_3586);
and U5975 (N_5975,N_4954,N_3932);
nor U5976 (N_5976,N_4468,N_4872);
or U5977 (N_5977,N_3794,N_3633);
nor U5978 (N_5978,N_2650,N_4023);
and U5979 (N_5979,N_2513,N_3678);
nor U5980 (N_5980,N_4613,N_3635);
and U5981 (N_5981,N_4550,N_3953);
or U5982 (N_5982,N_2531,N_2956);
nor U5983 (N_5983,N_2939,N_4860);
nor U5984 (N_5984,N_4182,N_3903);
nand U5985 (N_5985,N_4868,N_2680);
nand U5986 (N_5986,N_4142,N_3125);
or U5987 (N_5987,N_4639,N_3040);
and U5988 (N_5988,N_3129,N_4575);
or U5989 (N_5989,N_2872,N_3062);
nand U5990 (N_5990,N_3952,N_4174);
and U5991 (N_5991,N_3623,N_3636);
and U5992 (N_5992,N_4597,N_4402);
and U5993 (N_5993,N_4283,N_3338);
nor U5994 (N_5994,N_4251,N_4934);
and U5995 (N_5995,N_4809,N_2948);
and U5996 (N_5996,N_2850,N_4334);
and U5997 (N_5997,N_3157,N_4160);
or U5998 (N_5998,N_4637,N_4755);
nor U5999 (N_5999,N_3457,N_3882);
nand U6000 (N_6000,N_2652,N_3246);
nor U6001 (N_6001,N_3537,N_4552);
nor U6002 (N_6002,N_4515,N_4152);
or U6003 (N_6003,N_2858,N_4536);
and U6004 (N_6004,N_2904,N_3617);
nand U6005 (N_6005,N_3868,N_3295);
or U6006 (N_6006,N_2929,N_2727);
nand U6007 (N_6007,N_4845,N_3716);
nand U6008 (N_6008,N_2998,N_4683);
or U6009 (N_6009,N_3451,N_3990);
nor U6010 (N_6010,N_4479,N_4795);
nand U6011 (N_6011,N_3656,N_4276);
nand U6012 (N_6012,N_2843,N_2707);
and U6013 (N_6013,N_3995,N_4448);
nor U6014 (N_6014,N_2723,N_3560);
and U6015 (N_6015,N_2783,N_4466);
nand U6016 (N_6016,N_2925,N_3481);
nor U6017 (N_6017,N_3841,N_2878);
and U6018 (N_6018,N_4985,N_3366);
nor U6019 (N_6019,N_3315,N_4582);
and U6020 (N_6020,N_2787,N_4161);
or U6021 (N_6021,N_4676,N_4151);
nand U6022 (N_6022,N_4078,N_3943);
nand U6023 (N_6023,N_2870,N_2517);
nor U6024 (N_6024,N_3276,N_4877);
nand U6025 (N_6025,N_2613,N_2977);
nand U6026 (N_6026,N_3373,N_4573);
or U6027 (N_6027,N_2818,N_2919);
nor U6028 (N_6028,N_2824,N_4374);
nor U6029 (N_6029,N_4353,N_4297);
nor U6030 (N_6030,N_4427,N_4882);
nor U6031 (N_6031,N_3337,N_4835);
or U6032 (N_6032,N_4520,N_3551);
nand U6033 (N_6033,N_4568,N_4863);
or U6034 (N_6034,N_3875,N_4941);
or U6035 (N_6035,N_4006,N_4944);
and U6036 (N_6036,N_3961,N_4688);
and U6037 (N_6037,N_3979,N_3424);
nor U6038 (N_6038,N_4357,N_3730);
or U6039 (N_6039,N_3435,N_3616);
xnor U6040 (N_6040,N_4560,N_3611);
or U6041 (N_6041,N_3582,N_4995);
nand U6042 (N_6042,N_4508,N_3572);
or U6043 (N_6043,N_4478,N_4310);
and U6044 (N_6044,N_4702,N_3079);
nand U6045 (N_6045,N_4363,N_4157);
nand U6046 (N_6046,N_4498,N_4330);
nor U6047 (N_6047,N_2563,N_4643);
or U6048 (N_6048,N_2556,N_4942);
and U6049 (N_6049,N_2596,N_2519);
nor U6050 (N_6050,N_3892,N_3622);
and U6051 (N_6051,N_2574,N_4044);
and U6052 (N_6052,N_2789,N_3691);
nand U6053 (N_6053,N_3814,N_4951);
nor U6054 (N_6054,N_3549,N_3100);
and U6055 (N_6055,N_4250,N_2803);
or U6056 (N_6056,N_2992,N_3694);
and U6057 (N_6057,N_3418,N_3651);
nand U6058 (N_6058,N_3880,N_4524);
or U6059 (N_6059,N_3776,N_2962);
and U6060 (N_6060,N_4769,N_4572);
or U6061 (N_6061,N_4061,N_4428);
or U6062 (N_6062,N_4815,N_2751);
and U6063 (N_6063,N_2963,N_2809);
or U6064 (N_6064,N_3369,N_2810);
nor U6065 (N_6065,N_4273,N_2957);
or U6066 (N_6066,N_3970,N_3634);
nand U6067 (N_6067,N_3466,N_3512);
nand U6068 (N_6068,N_3734,N_4757);
nor U6069 (N_6069,N_4411,N_2827);
nand U6070 (N_6070,N_2684,N_3604);
nand U6071 (N_6071,N_3763,N_4982);
nor U6072 (N_6072,N_4454,N_4140);
nor U6073 (N_6073,N_2606,N_4423);
nor U6074 (N_6074,N_3931,N_4578);
nor U6075 (N_6075,N_4210,N_3548);
xnor U6076 (N_6076,N_4612,N_4999);
nor U6077 (N_6077,N_3380,N_4866);
nand U6078 (N_6078,N_3849,N_3465);
nand U6079 (N_6079,N_3239,N_2897);
nor U6080 (N_6080,N_3327,N_3899);
and U6081 (N_6081,N_4071,N_2761);
or U6082 (N_6082,N_2568,N_3186);
and U6083 (N_6083,N_4426,N_3101);
or U6084 (N_6084,N_2688,N_3398);
nor U6085 (N_6085,N_4434,N_3189);
nor U6086 (N_6086,N_4593,N_4979);
nor U6087 (N_6087,N_3508,N_3137);
nand U6088 (N_6088,N_4073,N_4899);
and U6089 (N_6089,N_2623,N_4422);
nand U6090 (N_6090,N_3877,N_4864);
nand U6091 (N_6091,N_4203,N_3872);
nand U6092 (N_6092,N_4748,N_4710);
and U6093 (N_6093,N_3049,N_2911);
and U6094 (N_6094,N_2961,N_4792);
and U6095 (N_6095,N_4617,N_2788);
nor U6096 (N_6096,N_4607,N_4370);
nor U6097 (N_6097,N_4535,N_4742);
or U6098 (N_6098,N_4344,N_3190);
or U6099 (N_6099,N_3753,N_4100);
or U6100 (N_6100,N_4227,N_4991);
nand U6101 (N_6101,N_2938,N_4469);
nor U6102 (N_6102,N_3063,N_4675);
nand U6103 (N_6103,N_3404,N_2509);
or U6104 (N_6104,N_4707,N_3831);
and U6105 (N_6105,N_3614,N_3052);
nand U6106 (N_6106,N_4085,N_3975);
and U6107 (N_6107,N_3935,N_3184);
nand U6108 (N_6108,N_2926,N_3103);
nand U6109 (N_6109,N_4723,N_4042);
and U6110 (N_6110,N_3749,N_3036);
xnor U6111 (N_6111,N_3449,N_4209);
and U6112 (N_6112,N_2607,N_4467);
nand U6113 (N_6113,N_4351,N_2669);
nand U6114 (N_6114,N_4482,N_4047);
nand U6115 (N_6115,N_4886,N_3818);
and U6116 (N_6116,N_4137,N_4068);
and U6117 (N_6117,N_4739,N_4309);
nand U6118 (N_6118,N_3155,N_2562);
or U6119 (N_6119,N_3908,N_3980);
and U6120 (N_6120,N_4037,N_3718);
or U6121 (N_6121,N_2535,N_2950);
and U6122 (N_6122,N_3726,N_3023);
nor U6123 (N_6123,N_3982,N_4224);
nand U6124 (N_6124,N_4247,N_3760);
or U6125 (N_6125,N_3406,N_3992);
nor U6126 (N_6126,N_3860,N_4540);
and U6127 (N_6127,N_3588,N_3024);
nor U6128 (N_6128,N_4783,N_3702);
or U6129 (N_6129,N_2614,N_3767);
nor U6130 (N_6130,N_4581,N_4292);
xor U6131 (N_6131,N_3247,N_3275);
nor U6132 (N_6132,N_4803,N_4386);
nor U6133 (N_6133,N_4465,N_4716);
nor U6134 (N_6134,N_4900,N_4518);
and U6135 (N_6135,N_3632,N_4109);
nor U6136 (N_6136,N_2887,N_2842);
nand U6137 (N_6137,N_4625,N_4751);
or U6138 (N_6138,N_4849,N_2585);
nor U6139 (N_6139,N_3168,N_3715);
nor U6140 (N_6140,N_2772,N_3409);
nor U6141 (N_6141,N_3682,N_4070);
nor U6142 (N_6142,N_3421,N_3733);
nor U6143 (N_6143,N_4138,N_3659);
or U6144 (N_6144,N_3919,N_4096);
and U6145 (N_6145,N_3735,N_4697);
and U6146 (N_6146,N_3443,N_4500);
and U6147 (N_6147,N_3857,N_4055);
nor U6148 (N_6148,N_3654,N_2629);
and U6149 (N_6149,N_4932,N_4185);
and U6150 (N_6150,N_3766,N_3224);
nand U6151 (N_6151,N_2792,N_4555);
or U6152 (N_6152,N_3592,N_4242);
nor U6153 (N_6153,N_2644,N_2927);
and U6154 (N_6154,N_4120,N_3086);
nand U6155 (N_6155,N_4525,N_2572);
nor U6156 (N_6156,N_3145,N_3534);
nor U6157 (N_6157,N_3647,N_2955);
nor U6158 (N_6158,N_4093,N_4901);
nor U6159 (N_6159,N_3837,N_4360);
and U6160 (N_6160,N_2646,N_3043);
nand U6161 (N_6161,N_3958,N_4202);
nor U6162 (N_6162,N_4438,N_2912);
nor U6163 (N_6163,N_4301,N_4662);
and U6164 (N_6164,N_4504,N_4918);
nor U6165 (N_6165,N_3399,N_4880);
nor U6166 (N_6166,N_4383,N_3501);
and U6167 (N_6167,N_4429,N_4773);
nand U6168 (N_6168,N_4318,N_3084);
or U6169 (N_6169,N_4208,N_4335);
and U6170 (N_6170,N_3721,N_4971);
nor U6171 (N_6171,N_3201,N_2900);
nor U6172 (N_6172,N_3411,N_3987);
and U6173 (N_6173,N_4756,N_3695);
nand U6174 (N_6174,N_3944,N_3082);
and U6175 (N_6175,N_3134,N_4103);
or U6176 (N_6176,N_3973,N_3667);
or U6177 (N_6177,N_3532,N_2877);
nor U6178 (N_6178,N_4691,N_3061);
or U6179 (N_6179,N_3347,N_2796);
or U6180 (N_6180,N_2500,N_4375);
xnor U6181 (N_6181,N_3595,N_3991);
or U6182 (N_6182,N_3516,N_3823);
or U6183 (N_6183,N_4111,N_3543);
or U6184 (N_6184,N_3050,N_4738);
or U6185 (N_6185,N_2816,N_4156);
xor U6186 (N_6186,N_4917,N_4449);
nand U6187 (N_6187,N_3402,N_3628);
or U6188 (N_6188,N_4747,N_3538);
nand U6189 (N_6189,N_2532,N_4098);
or U6190 (N_6190,N_4976,N_4681);
nand U6191 (N_6191,N_4667,N_3519);
nor U6192 (N_6192,N_4734,N_4993);
nand U6193 (N_6193,N_3432,N_3252);
nand U6194 (N_6194,N_3323,N_4847);
or U6195 (N_6195,N_2775,N_4050);
or U6196 (N_6196,N_2611,N_4084);
nor U6197 (N_6197,N_4326,N_4149);
or U6198 (N_6198,N_4911,N_3780);
nand U6199 (N_6199,N_4600,N_4958);
nor U6200 (N_6200,N_3087,N_3989);
nor U6201 (N_6201,N_2771,N_3664);
nor U6202 (N_6202,N_3166,N_2902);
nand U6203 (N_6203,N_4885,N_4459);
or U6204 (N_6204,N_2779,N_4807);
and U6205 (N_6205,N_4452,N_4059);
nor U6206 (N_6206,N_3091,N_3258);
nor U6207 (N_6207,N_4393,N_2541);
or U6208 (N_6208,N_3717,N_3017);
and U6209 (N_6209,N_4727,N_3124);
nand U6210 (N_6210,N_3613,N_4101);
and U6211 (N_6211,N_4824,N_3460);
or U6212 (N_6212,N_4476,N_4719);
nand U6213 (N_6213,N_2726,N_4350);
and U6214 (N_6214,N_4333,N_4177);
and U6215 (N_6215,N_3581,N_4306);
nand U6216 (N_6216,N_4026,N_3941);
or U6217 (N_6217,N_3738,N_4083);
nor U6218 (N_6218,N_3836,N_4332);
nor U6219 (N_6219,N_4870,N_4243);
xnor U6220 (N_6220,N_2662,N_4244);
and U6221 (N_6221,N_4502,N_3178);
and U6222 (N_6222,N_4923,N_3093);
and U6223 (N_6223,N_2762,N_4772);
nand U6224 (N_6224,N_3517,N_3701);
or U6225 (N_6225,N_2586,N_3556);
and U6226 (N_6226,N_2845,N_4461);
and U6227 (N_6227,N_3705,N_4554);
and U6228 (N_6228,N_3525,N_2759);
nor U6229 (N_6229,N_4458,N_3341);
or U6230 (N_6230,N_3074,N_2882);
nand U6231 (N_6231,N_4631,N_2773);
nand U6232 (N_6232,N_3302,N_3530);
nand U6233 (N_6233,N_4367,N_4019);
nor U6234 (N_6234,N_4316,N_4624);
and U6235 (N_6235,N_3503,N_3601);
nand U6236 (N_6236,N_3627,N_2617);
nor U6237 (N_6237,N_4014,N_3237);
nor U6238 (N_6238,N_3283,N_3010);
nor U6239 (N_6239,N_3173,N_3946);
or U6240 (N_6240,N_3331,N_3051);
and U6241 (N_6241,N_4721,N_3848);
xnor U6242 (N_6242,N_3914,N_3014);
nor U6243 (N_6243,N_4238,N_2823);
nand U6244 (N_6244,N_4188,N_4645);
nand U6245 (N_6245,N_4396,N_3112);
nand U6246 (N_6246,N_2604,N_4154);
nor U6247 (N_6247,N_4657,N_4246);
nand U6248 (N_6248,N_2790,N_2718);
and U6249 (N_6249,N_3522,N_2814);
nand U6250 (N_6250,N_3752,N_3990);
or U6251 (N_6251,N_2819,N_3804);
and U6252 (N_6252,N_4173,N_3916);
and U6253 (N_6253,N_4958,N_4497);
and U6254 (N_6254,N_3975,N_3785);
nand U6255 (N_6255,N_4232,N_3631);
nor U6256 (N_6256,N_3938,N_4516);
and U6257 (N_6257,N_3577,N_4804);
or U6258 (N_6258,N_3217,N_3570);
nand U6259 (N_6259,N_4920,N_3259);
nor U6260 (N_6260,N_4168,N_4218);
or U6261 (N_6261,N_2802,N_3878);
nor U6262 (N_6262,N_3942,N_3465);
and U6263 (N_6263,N_3972,N_3940);
nor U6264 (N_6264,N_4386,N_2786);
or U6265 (N_6265,N_2694,N_2918);
nand U6266 (N_6266,N_3280,N_3675);
nand U6267 (N_6267,N_4548,N_4806);
nand U6268 (N_6268,N_2549,N_4877);
nor U6269 (N_6269,N_4353,N_3657);
or U6270 (N_6270,N_3083,N_4471);
nor U6271 (N_6271,N_2969,N_4563);
nand U6272 (N_6272,N_4865,N_4032);
nor U6273 (N_6273,N_4989,N_4583);
and U6274 (N_6274,N_3549,N_2522);
or U6275 (N_6275,N_3271,N_2502);
nor U6276 (N_6276,N_2774,N_4953);
nor U6277 (N_6277,N_3578,N_2919);
or U6278 (N_6278,N_4263,N_3639);
or U6279 (N_6279,N_3286,N_3338);
xnor U6280 (N_6280,N_3684,N_4183);
nor U6281 (N_6281,N_2947,N_4300);
or U6282 (N_6282,N_4564,N_4247);
and U6283 (N_6283,N_4989,N_4774);
nor U6284 (N_6284,N_3566,N_3899);
and U6285 (N_6285,N_3700,N_3944);
nand U6286 (N_6286,N_3645,N_3569);
or U6287 (N_6287,N_4098,N_3502);
nor U6288 (N_6288,N_3093,N_4286);
nand U6289 (N_6289,N_4158,N_4698);
nor U6290 (N_6290,N_4596,N_2575);
and U6291 (N_6291,N_3039,N_3850);
and U6292 (N_6292,N_2671,N_2969);
nor U6293 (N_6293,N_4957,N_4959);
or U6294 (N_6294,N_3881,N_3177);
and U6295 (N_6295,N_4842,N_4250);
and U6296 (N_6296,N_4298,N_4051);
nor U6297 (N_6297,N_3179,N_2744);
nor U6298 (N_6298,N_3376,N_4363);
and U6299 (N_6299,N_3424,N_3903);
nor U6300 (N_6300,N_4339,N_4182);
nor U6301 (N_6301,N_4336,N_2872);
nor U6302 (N_6302,N_4661,N_4756);
or U6303 (N_6303,N_4493,N_4806);
and U6304 (N_6304,N_4316,N_4063);
nand U6305 (N_6305,N_3201,N_3659);
or U6306 (N_6306,N_3791,N_4854);
and U6307 (N_6307,N_2579,N_2607);
and U6308 (N_6308,N_2636,N_4899);
and U6309 (N_6309,N_3015,N_4936);
or U6310 (N_6310,N_4603,N_3472);
and U6311 (N_6311,N_2912,N_3873);
nand U6312 (N_6312,N_4038,N_2738);
and U6313 (N_6313,N_2843,N_3604);
nor U6314 (N_6314,N_3312,N_4757);
or U6315 (N_6315,N_2823,N_3699);
nor U6316 (N_6316,N_3737,N_4817);
nand U6317 (N_6317,N_2567,N_4447);
and U6318 (N_6318,N_4584,N_3837);
and U6319 (N_6319,N_2729,N_4036);
nor U6320 (N_6320,N_4233,N_2838);
and U6321 (N_6321,N_3417,N_2601);
or U6322 (N_6322,N_3935,N_2900);
nand U6323 (N_6323,N_2804,N_4288);
nand U6324 (N_6324,N_3560,N_3298);
and U6325 (N_6325,N_3453,N_3505);
nand U6326 (N_6326,N_3750,N_2904);
or U6327 (N_6327,N_4709,N_4452);
and U6328 (N_6328,N_4592,N_4550);
nand U6329 (N_6329,N_2737,N_4899);
nor U6330 (N_6330,N_2705,N_2915);
or U6331 (N_6331,N_2855,N_4969);
nor U6332 (N_6332,N_3964,N_3910);
nand U6333 (N_6333,N_4937,N_4920);
or U6334 (N_6334,N_3536,N_4084);
nor U6335 (N_6335,N_2666,N_4260);
and U6336 (N_6336,N_3999,N_2528);
or U6337 (N_6337,N_4904,N_2500);
nand U6338 (N_6338,N_4543,N_3413);
nand U6339 (N_6339,N_3474,N_4377);
or U6340 (N_6340,N_4627,N_4541);
nand U6341 (N_6341,N_3981,N_2756);
and U6342 (N_6342,N_4438,N_4576);
and U6343 (N_6343,N_3130,N_4675);
or U6344 (N_6344,N_4143,N_2957);
nor U6345 (N_6345,N_3328,N_3242);
nor U6346 (N_6346,N_3293,N_2502);
and U6347 (N_6347,N_3241,N_3152);
and U6348 (N_6348,N_4925,N_4772);
nor U6349 (N_6349,N_4600,N_4919);
nand U6350 (N_6350,N_3334,N_4600);
nand U6351 (N_6351,N_3137,N_4841);
or U6352 (N_6352,N_3080,N_2549);
xor U6353 (N_6353,N_4060,N_3407);
or U6354 (N_6354,N_3384,N_3092);
and U6355 (N_6355,N_4427,N_3345);
or U6356 (N_6356,N_4586,N_3691);
xor U6357 (N_6357,N_3226,N_3285);
nor U6358 (N_6358,N_4766,N_4933);
nand U6359 (N_6359,N_3535,N_4158);
nand U6360 (N_6360,N_2659,N_3737);
and U6361 (N_6361,N_3896,N_3180);
or U6362 (N_6362,N_4191,N_4353);
nor U6363 (N_6363,N_4211,N_2957);
and U6364 (N_6364,N_4475,N_3347);
nor U6365 (N_6365,N_3314,N_4666);
nand U6366 (N_6366,N_4192,N_4120);
or U6367 (N_6367,N_3873,N_3556);
nor U6368 (N_6368,N_2630,N_3187);
and U6369 (N_6369,N_3842,N_4864);
and U6370 (N_6370,N_2562,N_4004);
or U6371 (N_6371,N_3868,N_4294);
or U6372 (N_6372,N_2953,N_4367);
nand U6373 (N_6373,N_3114,N_3940);
and U6374 (N_6374,N_4487,N_4888);
nor U6375 (N_6375,N_4528,N_4945);
nor U6376 (N_6376,N_2925,N_4620);
or U6377 (N_6377,N_3139,N_3784);
nand U6378 (N_6378,N_3665,N_4103);
nor U6379 (N_6379,N_4904,N_3109);
and U6380 (N_6380,N_2711,N_3299);
xor U6381 (N_6381,N_3799,N_2836);
nor U6382 (N_6382,N_4017,N_3118);
nand U6383 (N_6383,N_3476,N_4581);
or U6384 (N_6384,N_3754,N_2806);
and U6385 (N_6385,N_3668,N_4232);
or U6386 (N_6386,N_4933,N_4381);
or U6387 (N_6387,N_2873,N_3553);
and U6388 (N_6388,N_3794,N_3016);
and U6389 (N_6389,N_4506,N_3225);
nor U6390 (N_6390,N_4521,N_2675);
or U6391 (N_6391,N_3116,N_2929);
and U6392 (N_6392,N_3542,N_4695);
xor U6393 (N_6393,N_4233,N_4630);
and U6394 (N_6394,N_3658,N_4163);
nand U6395 (N_6395,N_3983,N_3060);
and U6396 (N_6396,N_4413,N_3256);
or U6397 (N_6397,N_2957,N_4971);
nand U6398 (N_6398,N_4501,N_4127);
xor U6399 (N_6399,N_4599,N_4661);
or U6400 (N_6400,N_3941,N_4424);
and U6401 (N_6401,N_3932,N_3484);
or U6402 (N_6402,N_4564,N_2878);
nor U6403 (N_6403,N_4543,N_3591);
nor U6404 (N_6404,N_3933,N_4535);
nor U6405 (N_6405,N_3916,N_4460);
nand U6406 (N_6406,N_3304,N_2810);
and U6407 (N_6407,N_4437,N_3921);
nor U6408 (N_6408,N_4316,N_2822);
or U6409 (N_6409,N_4279,N_4979);
nand U6410 (N_6410,N_4000,N_4128);
nor U6411 (N_6411,N_3479,N_4048);
or U6412 (N_6412,N_4468,N_2674);
xor U6413 (N_6413,N_3950,N_3604);
nor U6414 (N_6414,N_3157,N_4709);
nor U6415 (N_6415,N_3129,N_2741);
or U6416 (N_6416,N_4903,N_4870);
nor U6417 (N_6417,N_4837,N_4234);
and U6418 (N_6418,N_4225,N_4452);
nor U6419 (N_6419,N_3486,N_2867);
nor U6420 (N_6420,N_3429,N_3498);
nor U6421 (N_6421,N_4637,N_3396);
or U6422 (N_6422,N_4357,N_4495);
or U6423 (N_6423,N_4955,N_4904);
nor U6424 (N_6424,N_2941,N_3975);
or U6425 (N_6425,N_3955,N_3720);
or U6426 (N_6426,N_3822,N_4033);
nor U6427 (N_6427,N_3959,N_3964);
nand U6428 (N_6428,N_3965,N_3301);
nor U6429 (N_6429,N_4473,N_2820);
and U6430 (N_6430,N_4784,N_4911);
nor U6431 (N_6431,N_4331,N_2519);
or U6432 (N_6432,N_3392,N_3831);
nand U6433 (N_6433,N_3043,N_4287);
nand U6434 (N_6434,N_4972,N_2915);
or U6435 (N_6435,N_3275,N_2594);
nand U6436 (N_6436,N_2514,N_2532);
nand U6437 (N_6437,N_3068,N_3770);
nand U6438 (N_6438,N_2756,N_3954);
nor U6439 (N_6439,N_2816,N_3532);
nor U6440 (N_6440,N_4268,N_4227);
and U6441 (N_6441,N_3723,N_4590);
nand U6442 (N_6442,N_4726,N_2539);
nor U6443 (N_6443,N_4343,N_4997);
xnor U6444 (N_6444,N_4418,N_4689);
and U6445 (N_6445,N_3785,N_4379);
nand U6446 (N_6446,N_3440,N_4381);
and U6447 (N_6447,N_3782,N_4340);
nor U6448 (N_6448,N_4510,N_2934);
and U6449 (N_6449,N_4643,N_2847);
or U6450 (N_6450,N_3297,N_4078);
nor U6451 (N_6451,N_4411,N_4308);
nand U6452 (N_6452,N_3651,N_4605);
or U6453 (N_6453,N_4699,N_3770);
nor U6454 (N_6454,N_4417,N_2534);
nand U6455 (N_6455,N_4780,N_4644);
nor U6456 (N_6456,N_4700,N_4911);
or U6457 (N_6457,N_4609,N_3059);
nor U6458 (N_6458,N_2512,N_4463);
nor U6459 (N_6459,N_2732,N_3572);
nor U6460 (N_6460,N_2572,N_3281);
or U6461 (N_6461,N_4225,N_3345);
or U6462 (N_6462,N_4988,N_3885);
and U6463 (N_6463,N_3906,N_3740);
nand U6464 (N_6464,N_3630,N_3902);
nor U6465 (N_6465,N_3373,N_2740);
and U6466 (N_6466,N_2655,N_3069);
and U6467 (N_6467,N_4107,N_2831);
and U6468 (N_6468,N_4157,N_2670);
nand U6469 (N_6469,N_3452,N_4974);
nor U6470 (N_6470,N_4357,N_4132);
nand U6471 (N_6471,N_4485,N_2894);
or U6472 (N_6472,N_3625,N_3696);
nor U6473 (N_6473,N_2597,N_2868);
and U6474 (N_6474,N_4774,N_4863);
or U6475 (N_6475,N_2907,N_2501);
nand U6476 (N_6476,N_4967,N_4843);
nand U6477 (N_6477,N_3233,N_3201);
and U6478 (N_6478,N_2841,N_3071);
and U6479 (N_6479,N_4875,N_3133);
or U6480 (N_6480,N_3998,N_4859);
nor U6481 (N_6481,N_3784,N_4080);
nand U6482 (N_6482,N_4260,N_2880);
nand U6483 (N_6483,N_4757,N_2989);
nand U6484 (N_6484,N_4006,N_4226);
nand U6485 (N_6485,N_2934,N_2549);
nand U6486 (N_6486,N_2560,N_4945);
or U6487 (N_6487,N_4684,N_4330);
and U6488 (N_6488,N_3120,N_3260);
nand U6489 (N_6489,N_4633,N_2821);
xor U6490 (N_6490,N_4521,N_3909);
nand U6491 (N_6491,N_2559,N_3274);
and U6492 (N_6492,N_4397,N_3249);
nor U6493 (N_6493,N_4969,N_3662);
nor U6494 (N_6494,N_2935,N_4747);
nor U6495 (N_6495,N_3305,N_3212);
nand U6496 (N_6496,N_2549,N_2641);
and U6497 (N_6497,N_4972,N_3671);
or U6498 (N_6498,N_2868,N_3222);
and U6499 (N_6499,N_4850,N_3308);
nand U6500 (N_6500,N_3231,N_2715);
or U6501 (N_6501,N_3030,N_3028);
and U6502 (N_6502,N_4502,N_4083);
or U6503 (N_6503,N_4535,N_4289);
nor U6504 (N_6504,N_2870,N_4570);
nand U6505 (N_6505,N_4576,N_2507);
xor U6506 (N_6506,N_4983,N_3451);
nor U6507 (N_6507,N_2876,N_4513);
nor U6508 (N_6508,N_4751,N_3550);
and U6509 (N_6509,N_4318,N_2689);
nor U6510 (N_6510,N_2880,N_2597);
nor U6511 (N_6511,N_4922,N_3184);
nor U6512 (N_6512,N_3565,N_3783);
or U6513 (N_6513,N_3097,N_3669);
nor U6514 (N_6514,N_4557,N_3818);
nor U6515 (N_6515,N_2709,N_4023);
and U6516 (N_6516,N_2728,N_4493);
nor U6517 (N_6517,N_4195,N_2744);
and U6518 (N_6518,N_4875,N_4520);
or U6519 (N_6519,N_4487,N_3701);
nor U6520 (N_6520,N_4222,N_2924);
xor U6521 (N_6521,N_3163,N_3037);
and U6522 (N_6522,N_3607,N_3059);
nor U6523 (N_6523,N_3368,N_2983);
or U6524 (N_6524,N_2754,N_2996);
or U6525 (N_6525,N_4357,N_2998);
and U6526 (N_6526,N_4500,N_2914);
and U6527 (N_6527,N_3219,N_2933);
nand U6528 (N_6528,N_3592,N_4130);
and U6529 (N_6529,N_3585,N_2625);
and U6530 (N_6530,N_2578,N_4096);
and U6531 (N_6531,N_4950,N_4738);
or U6532 (N_6532,N_4692,N_3288);
and U6533 (N_6533,N_3670,N_4182);
nand U6534 (N_6534,N_3388,N_3935);
or U6535 (N_6535,N_4769,N_3615);
and U6536 (N_6536,N_3810,N_4436);
xnor U6537 (N_6537,N_4947,N_3486);
nand U6538 (N_6538,N_2769,N_3208);
or U6539 (N_6539,N_4858,N_3262);
nor U6540 (N_6540,N_4129,N_3217);
nor U6541 (N_6541,N_3122,N_4713);
xor U6542 (N_6542,N_4842,N_4571);
or U6543 (N_6543,N_3632,N_4364);
nand U6544 (N_6544,N_4677,N_3969);
or U6545 (N_6545,N_4727,N_2936);
nand U6546 (N_6546,N_4425,N_4410);
or U6547 (N_6547,N_4614,N_4514);
or U6548 (N_6548,N_3118,N_2543);
or U6549 (N_6549,N_3261,N_2550);
and U6550 (N_6550,N_4730,N_4692);
nand U6551 (N_6551,N_4747,N_4148);
nor U6552 (N_6552,N_3370,N_3626);
nor U6553 (N_6553,N_2875,N_4997);
and U6554 (N_6554,N_2816,N_4118);
and U6555 (N_6555,N_3369,N_3361);
or U6556 (N_6556,N_3522,N_3153);
xor U6557 (N_6557,N_4456,N_2953);
nand U6558 (N_6558,N_3244,N_3993);
nand U6559 (N_6559,N_4572,N_4057);
or U6560 (N_6560,N_4891,N_4176);
nand U6561 (N_6561,N_3921,N_4087);
nand U6562 (N_6562,N_3998,N_3088);
or U6563 (N_6563,N_3297,N_3255);
and U6564 (N_6564,N_3050,N_3122);
or U6565 (N_6565,N_4226,N_3650);
nor U6566 (N_6566,N_4652,N_3637);
and U6567 (N_6567,N_3201,N_3285);
and U6568 (N_6568,N_4849,N_3729);
and U6569 (N_6569,N_2912,N_2924);
nor U6570 (N_6570,N_4768,N_3639);
nand U6571 (N_6571,N_4116,N_4423);
nand U6572 (N_6572,N_3300,N_3444);
nor U6573 (N_6573,N_2815,N_3655);
and U6574 (N_6574,N_4254,N_2947);
nand U6575 (N_6575,N_2800,N_3178);
or U6576 (N_6576,N_3778,N_3936);
nor U6577 (N_6577,N_3423,N_2773);
nand U6578 (N_6578,N_3082,N_4008);
nor U6579 (N_6579,N_3925,N_2882);
nand U6580 (N_6580,N_2636,N_3914);
nor U6581 (N_6581,N_3781,N_3424);
and U6582 (N_6582,N_3266,N_2729);
or U6583 (N_6583,N_4506,N_3490);
nor U6584 (N_6584,N_4366,N_2948);
and U6585 (N_6585,N_4973,N_3303);
and U6586 (N_6586,N_3436,N_4184);
or U6587 (N_6587,N_4540,N_2574);
nor U6588 (N_6588,N_2613,N_2754);
nor U6589 (N_6589,N_4605,N_4514);
nand U6590 (N_6590,N_4565,N_3281);
xnor U6591 (N_6591,N_4168,N_3730);
and U6592 (N_6592,N_3801,N_2656);
nand U6593 (N_6593,N_2818,N_4743);
and U6594 (N_6594,N_3004,N_2701);
nor U6595 (N_6595,N_4668,N_3281);
and U6596 (N_6596,N_4013,N_3014);
and U6597 (N_6597,N_2996,N_4955);
or U6598 (N_6598,N_4961,N_4109);
or U6599 (N_6599,N_4845,N_3517);
nand U6600 (N_6600,N_2747,N_3475);
or U6601 (N_6601,N_4254,N_2906);
or U6602 (N_6602,N_4990,N_2533);
or U6603 (N_6603,N_3756,N_3104);
nor U6604 (N_6604,N_3042,N_2621);
nand U6605 (N_6605,N_3205,N_2958);
nand U6606 (N_6606,N_4917,N_3237);
or U6607 (N_6607,N_4029,N_4988);
and U6608 (N_6608,N_2867,N_3033);
or U6609 (N_6609,N_3672,N_4516);
nor U6610 (N_6610,N_4906,N_4020);
or U6611 (N_6611,N_3923,N_2690);
or U6612 (N_6612,N_2975,N_2886);
nor U6613 (N_6613,N_3045,N_2830);
and U6614 (N_6614,N_3973,N_4338);
and U6615 (N_6615,N_3907,N_3972);
and U6616 (N_6616,N_4388,N_3493);
or U6617 (N_6617,N_2755,N_4190);
and U6618 (N_6618,N_2946,N_4585);
or U6619 (N_6619,N_3262,N_2503);
nor U6620 (N_6620,N_4309,N_3212);
and U6621 (N_6621,N_3429,N_4952);
nand U6622 (N_6622,N_3037,N_4029);
and U6623 (N_6623,N_2708,N_4995);
nor U6624 (N_6624,N_4726,N_2915);
nand U6625 (N_6625,N_3453,N_3215);
nand U6626 (N_6626,N_3491,N_3383);
nor U6627 (N_6627,N_3295,N_4919);
or U6628 (N_6628,N_3921,N_4905);
nor U6629 (N_6629,N_4560,N_4478);
nand U6630 (N_6630,N_3843,N_3141);
and U6631 (N_6631,N_2622,N_4593);
and U6632 (N_6632,N_4812,N_3381);
nor U6633 (N_6633,N_4885,N_2682);
nand U6634 (N_6634,N_3861,N_4810);
nor U6635 (N_6635,N_4637,N_4242);
and U6636 (N_6636,N_4783,N_3535);
nand U6637 (N_6637,N_4105,N_4121);
or U6638 (N_6638,N_3800,N_4527);
or U6639 (N_6639,N_4655,N_3360);
and U6640 (N_6640,N_4795,N_4525);
nand U6641 (N_6641,N_2564,N_4001);
and U6642 (N_6642,N_4249,N_2620);
xnor U6643 (N_6643,N_2512,N_4916);
and U6644 (N_6644,N_4470,N_3282);
nand U6645 (N_6645,N_3535,N_3034);
or U6646 (N_6646,N_4298,N_2883);
nor U6647 (N_6647,N_4253,N_2913);
or U6648 (N_6648,N_4734,N_3685);
nand U6649 (N_6649,N_4637,N_4819);
nor U6650 (N_6650,N_3238,N_4731);
nor U6651 (N_6651,N_4872,N_3362);
or U6652 (N_6652,N_4934,N_4673);
nor U6653 (N_6653,N_2806,N_4510);
nand U6654 (N_6654,N_4279,N_3080);
nand U6655 (N_6655,N_3620,N_3146);
nand U6656 (N_6656,N_4044,N_3125);
and U6657 (N_6657,N_4184,N_3420);
nand U6658 (N_6658,N_4187,N_2713);
nand U6659 (N_6659,N_2906,N_3808);
nor U6660 (N_6660,N_2762,N_2807);
or U6661 (N_6661,N_2817,N_3207);
or U6662 (N_6662,N_3983,N_4781);
or U6663 (N_6663,N_3582,N_3211);
or U6664 (N_6664,N_4152,N_3408);
nand U6665 (N_6665,N_3239,N_3955);
and U6666 (N_6666,N_4938,N_2539);
or U6667 (N_6667,N_3716,N_3520);
nor U6668 (N_6668,N_3501,N_3966);
or U6669 (N_6669,N_4919,N_4008);
or U6670 (N_6670,N_3481,N_3568);
nand U6671 (N_6671,N_3258,N_4300);
nand U6672 (N_6672,N_4341,N_2886);
xnor U6673 (N_6673,N_3938,N_3358);
or U6674 (N_6674,N_3848,N_4308);
and U6675 (N_6675,N_3685,N_4905);
or U6676 (N_6676,N_4075,N_4432);
nor U6677 (N_6677,N_4058,N_4435);
or U6678 (N_6678,N_4560,N_4318);
and U6679 (N_6679,N_2729,N_3432);
and U6680 (N_6680,N_4880,N_3674);
and U6681 (N_6681,N_2770,N_2874);
nor U6682 (N_6682,N_3274,N_3966);
and U6683 (N_6683,N_4999,N_3705);
and U6684 (N_6684,N_4848,N_3110);
nor U6685 (N_6685,N_3588,N_3858);
nand U6686 (N_6686,N_3680,N_2886);
or U6687 (N_6687,N_4027,N_2722);
or U6688 (N_6688,N_4833,N_4883);
nor U6689 (N_6689,N_4414,N_3230);
nor U6690 (N_6690,N_4787,N_4038);
nand U6691 (N_6691,N_4488,N_4957);
nor U6692 (N_6692,N_3351,N_4734);
nand U6693 (N_6693,N_2644,N_3046);
or U6694 (N_6694,N_4332,N_3896);
or U6695 (N_6695,N_2911,N_4219);
or U6696 (N_6696,N_2902,N_2558);
or U6697 (N_6697,N_4732,N_3455);
nor U6698 (N_6698,N_3519,N_3654);
nor U6699 (N_6699,N_3556,N_3370);
xor U6700 (N_6700,N_2559,N_3369);
and U6701 (N_6701,N_2690,N_4064);
nor U6702 (N_6702,N_3494,N_4864);
nand U6703 (N_6703,N_2702,N_2587);
or U6704 (N_6704,N_4782,N_3861);
nor U6705 (N_6705,N_3396,N_3964);
xnor U6706 (N_6706,N_4678,N_4005);
or U6707 (N_6707,N_4873,N_3984);
nand U6708 (N_6708,N_4033,N_3673);
or U6709 (N_6709,N_2847,N_3159);
nand U6710 (N_6710,N_2797,N_3552);
nor U6711 (N_6711,N_2803,N_4317);
and U6712 (N_6712,N_3325,N_3806);
or U6713 (N_6713,N_3016,N_2901);
nor U6714 (N_6714,N_2591,N_4006);
nor U6715 (N_6715,N_2866,N_2958);
nand U6716 (N_6716,N_4225,N_3793);
nor U6717 (N_6717,N_2657,N_4040);
and U6718 (N_6718,N_3596,N_2586);
or U6719 (N_6719,N_2658,N_4362);
or U6720 (N_6720,N_4916,N_4834);
or U6721 (N_6721,N_4246,N_2596);
xor U6722 (N_6722,N_2898,N_3079);
or U6723 (N_6723,N_2672,N_4689);
nand U6724 (N_6724,N_4689,N_3025);
or U6725 (N_6725,N_4326,N_2842);
nand U6726 (N_6726,N_4371,N_2913);
or U6727 (N_6727,N_4988,N_2774);
xnor U6728 (N_6728,N_3706,N_4097);
nand U6729 (N_6729,N_4011,N_2881);
nand U6730 (N_6730,N_4654,N_3977);
or U6731 (N_6731,N_4617,N_4228);
nor U6732 (N_6732,N_3630,N_2885);
or U6733 (N_6733,N_4607,N_2690);
or U6734 (N_6734,N_4277,N_3429);
nand U6735 (N_6735,N_4031,N_2763);
and U6736 (N_6736,N_4739,N_2709);
and U6737 (N_6737,N_4168,N_3792);
nor U6738 (N_6738,N_2647,N_4110);
or U6739 (N_6739,N_4922,N_3719);
or U6740 (N_6740,N_3028,N_4898);
or U6741 (N_6741,N_2581,N_4607);
nor U6742 (N_6742,N_4635,N_3942);
or U6743 (N_6743,N_3037,N_4228);
and U6744 (N_6744,N_4623,N_3452);
nand U6745 (N_6745,N_3400,N_3566);
and U6746 (N_6746,N_2774,N_2832);
nand U6747 (N_6747,N_4494,N_3774);
nor U6748 (N_6748,N_4797,N_4211);
or U6749 (N_6749,N_3986,N_4273);
or U6750 (N_6750,N_3903,N_4819);
nand U6751 (N_6751,N_3003,N_2761);
nor U6752 (N_6752,N_3328,N_2749);
xnor U6753 (N_6753,N_4088,N_4008);
or U6754 (N_6754,N_3854,N_2887);
nor U6755 (N_6755,N_4916,N_2903);
or U6756 (N_6756,N_3810,N_3111);
nor U6757 (N_6757,N_3708,N_4400);
nand U6758 (N_6758,N_4050,N_4274);
or U6759 (N_6759,N_3547,N_3932);
or U6760 (N_6760,N_4094,N_2706);
nor U6761 (N_6761,N_4837,N_4834);
or U6762 (N_6762,N_3763,N_4456);
and U6763 (N_6763,N_2581,N_3374);
nor U6764 (N_6764,N_4815,N_3516);
nand U6765 (N_6765,N_4819,N_4884);
nand U6766 (N_6766,N_3779,N_4187);
nand U6767 (N_6767,N_3965,N_2751);
and U6768 (N_6768,N_4554,N_4627);
nor U6769 (N_6769,N_3700,N_3067);
nand U6770 (N_6770,N_3133,N_4033);
and U6771 (N_6771,N_3747,N_4567);
and U6772 (N_6772,N_3719,N_4971);
or U6773 (N_6773,N_3457,N_2795);
and U6774 (N_6774,N_2601,N_4344);
and U6775 (N_6775,N_2698,N_4382);
or U6776 (N_6776,N_4298,N_3857);
or U6777 (N_6777,N_3044,N_2768);
and U6778 (N_6778,N_4253,N_3370);
nor U6779 (N_6779,N_4443,N_4446);
or U6780 (N_6780,N_3489,N_2564);
and U6781 (N_6781,N_4462,N_2738);
and U6782 (N_6782,N_4446,N_4373);
and U6783 (N_6783,N_3929,N_4093);
nand U6784 (N_6784,N_4975,N_4670);
or U6785 (N_6785,N_4829,N_4109);
nor U6786 (N_6786,N_3563,N_3505);
or U6787 (N_6787,N_4251,N_4077);
and U6788 (N_6788,N_3773,N_3582);
or U6789 (N_6789,N_4596,N_3684);
nor U6790 (N_6790,N_4472,N_3928);
nor U6791 (N_6791,N_3159,N_3302);
and U6792 (N_6792,N_4634,N_2584);
and U6793 (N_6793,N_4494,N_3850);
nand U6794 (N_6794,N_4156,N_3271);
and U6795 (N_6795,N_3022,N_2732);
nor U6796 (N_6796,N_2849,N_4073);
or U6797 (N_6797,N_2684,N_3429);
nor U6798 (N_6798,N_4350,N_2658);
xor U6799 (N_6799,N_4956,N_2716);
or U6800 (N_6800,N_4783,N_3827);
or U6801 (N_6801,N_2869,N_3182);
nand U6802 (N_6802,N_4790,N_4629);
and U6803 (N_6803,N_2603,N_3929);
nor U6804 (N_6804,N_3901,N_4811);
nand U6805 (N_6805,N_2614,N_3884);
nand U6806 (N_6806,N_4908,N_4463);
nor U6807 (N_6807,N_4358,N_3470);
nand U6808 (N_6808,N_3036,N_3117);
nor U6809 (N_6809,N_3173,N_3748);
xnor U6810 (N_6810,N_4660,N_4790);
and U6811 (N_6811,N_4011,N_3117);
and U6812 (N_6812,N_2820,N_2907);
and U6813 (N_6813,N_3027,N_3604);
nor U6814 (N_6814,N_3794,N_4449);
or U6815 (N_6815,N_3969,N_3871);
and U6816 (N_6816,N_2982,N_3779);
nand U6817 (N_6817,N_3977,N_2819);
or U6818 (N_6818,N_3131,N_4406);
nand U6819 (N_6819,N_3406,N_3458);
nor U6820 (N_6820,N_2925,N_4941);
nand U6821 (N_6821,N_4077,N_4881);
nand U6822 (N_6822,N_3795,N_4026);
and U6823 (N_6823,N_2684,N_3539);
xnor U6824 (N_6824,N_4010,N_3910);
xor U6825 (N_6825,N_3121,N_4817);
nand U6826 (N_6826,N_4082,N_3525);
or U6827 (N_6827,N_4205,N_4625);
and U6828 (N_6828,N_4879,N_4058);
and U6829 (N_6829,N_2902,N_4490);
or U6830 (N_6830,N_3605,N_4674);
and U6831 (N_6831,N_3949,N_4681);
nand U6832 (N_6832,N_2681,N_3127);
and U6833 (N_6833,N_3363,N_3867);
or U6834 (N_6834,N_3199,N_3561);
or U6835 (N_6835,N_4218,N_3569);
or U6836 (N_6836,N_4629,N_4933);
or U6837 (N_6837,N_3683,N_4072);
and U6838 (N_6838,N_3667,N_2890);
or U6839 (N_6839,N_4718,N_2775);
or U6840 (N_6840,N_2721,N_4143);
nor U6841 (N_6841,N_2783,N_3376);
nand U6842 (N_6842,N_4260,N_2834);
and U6843 (N_6843,N_3208,N_4262);
nand U6844 (N_6844,N_2661,N_3051);
and U6845 (N_6845,N_3089,N_4969);
nand U6846 (N_6846,N_3321,N_4057);
nand U6847 (N_6847,N_4289,N_4300);
nand U6848 (N_6848,N_3995,N_4402);
and U6849 (N_6849,N_4155,N_3389);
nand U6850 (N_6850,N_3861,N_2926);
and U6851 (N_6851,N_4452,N_2779);
and U6852 (N_6852,N_4380,N_4421);
nor U6853 (N_6853,N_3258,N_2912);
nor U6854 (N_6854,N_4787,N_2822);
nor U6855 (N_6855,N_2887,N_2596);
or U6856 (N_6856,N_3529,N_2548);
or U6857 (N_6857,N_3754,N_2951);
nor U6858 (N_6858,N_3581,N_4442);
nor U6859 (N_6859,N_3618,N_3318);
and U6860 (N_6860,N_3804,N_4224);
and U6861 (N_6861,N_4963,N_3277);
nor U6862 (N_6862,N_4445,N_3809);
and U6863 (N_6863,N_4241,N_4741);
and U6864 (N_6864,N_4400,N_4678);
nor U6865 (N_6865,N_4999,N_4707);
and U6866 (N_6866,N_4331,N_3349);
nor U6867 (N_6867,N_2909,N_2874);
nand U6868 (N_6868,N_2752,N_4448);
and U6869 (N_6869,N_3109,N_2809);
and U6870 (N_6870,N_4835,N_4744);
and U6871 (N_6871,N_3641,N_3780);
nand U6872 (N_6872,N_2861,N_2545);
or U6873 (N_6873,N_4178,N_4440);
and U6874 (N_6874,N_4664,N_4258);
or U6875 (N_6875,N_4241,N_2906);
nor U6876 (N_6876,N_4491,N_4535);
nand U6877 (N_6877,N_3477,N_4631);
nand U6878 (N_6878,N_4340,N_2529);
nand U6879 (N_6879,N_3407,N_4012);
xor U6880 (N_6880,N_3421,N_4810);
nand U6881 (N_6881,N_4100,N_4788);
nor U6882 (N_6882,N_4497,N_4227);
or U6883 (N_6883,N_4030,N_2836);
nand U6884 (N_6884,N_4091,N_3369);
and U6885 (N_6885,N_4992,N_4169);
and U6886 (N_6886,N_3580,N_4853);
nand U6887 (N_6887,N_4511,N_4545);
and U6888 (N_6888,N_2979,N_4631);
nor U6889 (N_6889,N_2592,N_4371);
nand U6890 (N_6890,N_3947,N_3867);
nor U6891 (N_6891,N_3381,N_4594);
nand U6892 (N_6892,N_4170,N_4715);
or U6893 (N_6893,N_4895,N_4336);
nand U6894 (N_6894,N_4121,N_3656);
and U6895 (N_6895,N_4432,N_3256);
and U6896 (N_6896,N_3623,N_3179);
nor U6897 (N_6897,N_3279,N_2913);
and U6898 (N_6898,N_3667,N_3429);
or U6899 (N_6899,N_4733,N_4901);
and U6900 (N_6900,N_4416,N_3768);
xor U6901 (N_6901,N_3631,N_3224);
nand U6902 (N_6902,N_2696,N_2521);
nand U6903 (N_6903,N_4326,N_4053);
nor U6904 (N_6904,N_3881,N_2836);
nor U6905 (N_6905,N_4793,N_2815);
or U6906 (N_6906,N_2835,N_2803);
and U6907 (N_6907,N_3454,N_2857);
or U6908 (N_6908,N_2584,N_3060);
nor U6909 (N_6909,N_3359,N_2928);
nor U6910 (N_6910,N_3050,N_4324);
or U6911 (N_6911,N_2795,N_2538);
nand U6912 (N_6912,N_3956,N_4397);
or U6913 (N_6913,N_3124,N_3075);
nand U6914 (N_6914,N_3035,N_4021);
and U6915 (N_6915,N_2793,N_4456);
or U6916 (N_6916,N_4980,N_3885);
or U6917 (N_6917,N_2733,N_2801);
nor U6918 (N_6918,N_4540,N_3570);
or U6919 (N_6919,N_3052,N_4640);
or U6920 (N_6920,N_4804,N_3853);
nor U6921 (N_6921,N_3445,N_3605);
nor U6922 (N_6922,N_4260,N_4570);
and U6923 (N_6923,N_4304,N_2691);
nand U6924 (N_6924,N_3846,N_4601);
and U6925 (N_6925,N_4927,N_3310);
and U6926 (N_6926,N_3420,N_2984);
nand U6927 (N_6927,N_2729,N_4101);
nand U6928 (N_6928,N_2594,N_4460);
and U6929 (N_6929,N_3728,N_3731);
and U6930 (N_6930,N_3000,N_3863);
nand U6931 (N_6931,N_3710,N_2570);
nand U6932 (N_6932,N_4486,N_4166);
or U6933 (N_6933,N_2859,N_2824);
nor U6934 (N_6934,N_3002,N_3058);
nand U6935 (N_6935,N_4240,N_4196);
nor U6936 (N_6936,N_3148,N_4096);
nor U6937 (N_6937,N_4946,N_3137);
and U6938 (N_6938,N_3068,N_3925);
or U6939 (N_6939,N_4380,N_3723);
or U6940 (N_6940,N_3826,N_4700);
or U6941 (N_6941,N_4642,N_4919);
nor U6942 (N_6942,N_4492,N_2850);
and U6943 (N_6943,N_3185,N_4915);
or U6944 (N_6944,N_4084,N_2707);
and U6945 (N_6945,N_3515,N_3659);
and U6946 (N_6946,N_3685,N_2772);
or U6947 (N_6947,N_4002,N_3536);
or U6948 (N_6948,N_4423,N_2575);
nor U6949 (N_6949,N_4461,N_2788);
nor U6950 (N_6950,N_3355,N_3053);
or U6951 (N_6951,N_2876,N_4215);
nor U6952 (N_6952,N_4045,N_3896);
nand U6953 (N_6953,N_2902,N_2629);
or U6954 (N_6954,N_2657,N_3026);
nand U6955 (N_6955,N_2729,N_4312);
nand U6956 (N_6956,N_3105,N_4660);
and U6957 (N_6957,N_3305,N_4774);
nand U6958 (N_6958,N_3445,N_3031);
or U6959 (N_6959,N_3483,N_3058);
xnor U6960 (N_6960,N_2874,N_3855);
and U6961 (N_6961,N_4850,N_3830);
or U6962 (N_6962,N_3587,N_3582);
or U6963 (N_6963,N_4939,N_3779);
or U6964 (N_6964,N_2865,N_3094);
nor U6965 (N_6965,N_3234,N_4011);
or U6966 (N_6966,N_4413,N_2996);
or U6967 (N_6967,N_4090,N_2749);
nand U6968 (N_6968,N_4365,N_3365);
and U6969 (N_6969,N_2812,N_4135);
or U6970 (N_6970,N_2507,N_3867);
nor U6971 (N_6971,N_2963,N_3491);
nor U6972 (N_6972,N_3016,N_2881);
nand U6973 (N_6973,N_2973,N_2576);
nor U6974 (N_6974,N_3319,N_4009);
nand U6975 (N_6975,N_2704,N_2765);
nor U6976 (N_6976,N_3054,N_4552);
or U6977 (N_6977,N_4514,N_4189);
and U6978 (N_6978,N_2712,N_4776);
nor U6979 (N_6979,N_2791,N_3469);
nand U6980 (N_6980,N_2572,N_4644);
or U6981 (N_6981,N_3033,N_4625);
nand U6982 (N_6982,N_4970,N_3615);
and U6983 (N_6983,N_2905,N_4345);
or U6984 (N_6984,N_2753,N_3463);
nor U6985 (N_6985,N_4286,N_2933);
and U6986 (N_6986,N_3672,N_4384);
or U6987 (N_6987,N_4472,N_3331);
nand U6988 (N_6988,N_4607,N_4391);
or U6989 (N_6989,N_3353,N_3448);
nor U6990 (N_6990,N_4077,N_3002);
or U6991 (N_6991,N_2679,N_2613);
nand U6992 (N_6992,N_3332,N_3420);
nor U6993 (N_6993,N_3508,N_3630);
or U6994 (N_6994,N_3624,N_3502);
and U6995 (N_6995,N_2585,N_4640);
and U6996 (N_6996,N_3574,N_2967);
and U6997 (N_6997,N_3214,N_4066);
nand U6998 (N_6998,N_4685,N_3179);
xnor U6999 (N_6999,N_2976,N_3980);
or U7000 (N_7000,N_3039,N_2533);
and U7001 (N_7001,N_4195,N_2704);
nor U7002 (N_7002,N_4609,N_3587);
or U7003 (N_7003,N_4860,N_2732);
or U7004 (N_7004,N_3515,N_3127);
nand U7005 (N_7005,N_4598,N_4601);
and U7006 (N_7006,N_2995,N_2824);
nor U7007 (N_7007,N_3416,N_4655);
and U7008 (N_7008,N_4588,N_3681);
or U7009 (N_7009,N_4460,N_3244);
nand U7010 (N_7010,N_4375,N_3572);
or U7011 (N_7011,N_4128,N_3803);
xor U7012 (N_7012,N_4598,N_4916);
and U7013 (N_7013,N_3282,N_4795);
or U7014 (N_7014,N_3206,N_3560);
nand U7015 (N_7015,N_4801,N_3668);
nor U7016 (N_7016,N_3331,N_3093);
nand U7017 (N_7017,N_4398,N_3315);
and U7018 (N_7018,N_3003,N_3299);
nand U7019 (N_7019,N_4442,N_4177);
nand U7020 (N_7020,N_4165,N_3157);
nand U7021 (N_7021,N_4914,N_4886);
and U7022 (N_7022,N_2916,N_4758);
or U7023 (N_7023,N_4506,N_2741);
and U7024 (N_7024,N_3662,N_3385);
or U7025 (N_7025,N_3717,N_3666);
nand U7026 (N_7026,N_3366,N_4205);
nand U7027 (N_7027,N_2872,N_4393);
nand U7028 (N_7028,N_4429,N_4086);
and U7029 (N_7029,N_2893,N_4252);
and U7030 (N_7030,N_2645,N_3947);
and U7031 (N_7031,N_3023,N_3328);
or U7032 (N_7032,N_4391,N_4707);
and U7033 (N_7033,N_3673,N_3764);
or U7034 (N_7034,N_4056,N_3652);
or U7035 (N_7035,N_3626,N_3975);
and U7036 (N_7036,N_3969,N_2667);
or U7037 (N_7037,N_3177,N_4659);
nand U7038 (N_7038,N_2750,N_4705);
and U7039 (N_7039,N_3952,N_3963);
nand U7040 (N_7040,N_3018,N_3604);
nand U7041 (N_7041,N_3355,N_4116);
nand U7042 (N_7042,N_4927,N_4717);
and U7043 (N_7043,N_4711,N_4303);
nor U7044 (N_7044,N_4414,N_4678);
nand U7045 (N_7045,N_3882,N_2869);
or U7046 (N_7046,N_3078,N_2640);
nand U7047 (N_7047,N_2768,N_3630);
and U7048 (N_7048,N_3766,N_4106);
nor U7049 (N_7049,N_3500,N_3079);
nand U7050 (N_7050,N_4438,N_4098);
or U7051 (N_7051,N_2562,N_2833);
nor U7052 (N_7052,N_3347,N_4484);
and U7053 (N_7053,N_4294,N_4493);
nor U7054 (N_7054,N_3746,N_4484);
and U7055 (N_7055,N_4047,N_2874);
nor U7056 (N_7056,N_3729,N_3479);
or U7057 (N_7057,N_3554,N_2764);
or U7058 (N_7058,N_2643,N_2800);
nor U7059 (N_7059,N_4224,N_3530);
or U7060 (N_7060,N_3096,N_4304);
or U7061 (N_7061,N_3345,N_2862);
or U7062 (N_7062,N_4940,N_4560);
or U7063 (N_7063,N_2651,N_4251);
or U7064 (N_7064,N_4404,N_3698);
nor U7065 (N_7065,N_3031,N_4913);
nor U7066 (N_7066,N_3223,N_3876);
or U7067 (N_7067,N_4403,N_3451);
nor U7068 (N_7068,N_4250,N_4047);
nor U7069 (N_7069,N_4821,N_3728);
or U7070 (N_7070,N_3995,N_4007);
and U7071 (N_7071,N_3204,N_4446);
or U7072 (N_7072,N_3402,N_4006);
xor U7073 (N_7073,N_4989,N_3612);
nand U7074 (N_7074,N_2618,N_2937);
or U7075 (N_7075,N_4928,N_3696);
or U7076 (N_7076,N_3452,N_3093);
and U7077 (N_7077,N_3504,N_4543);
and U7078 (N_7078,N_3124,N_3524);
nand U7079 (N_7079,N_2978,N_3645);
nand U7080 (N_7080,N_3582,N_3482);
nor U7081 (N_7081,N_2558,N_2600);
nand U7082 (N_7082,N_3578,N_2771);
and U7083 (N_7083,N_2633,N_4188);
nand U7084 (N_7084,N_4458,N_4187);
nor U7085 (N_7085,N_2990,N_2995);
nor U7086 (N_7086,N_3346,N_2579);
nor U7087 (N_7087,N_2557,N_4298);
nand U7088 (N_7088,N_4323,N_4263);
xnor U7089 (N_7089,N_3978,N_3441);
nor U7090 (N_7090,N_4275,N_4574);
and U7091 (N_7091,N_4395,N_2502);
nand U7092 (N_7092,N_3842,N_4125);
xor U7093 (N_7093,N_4331,N_2595);
nor U7094 (N_7094,N_4741,N_3988);
nand U7095 (N_7095,N_3681,N_3342);
and U7096 (N_7096,N_4390,N_3084);
or U7097 (N_7097,N_3967,N_4380);
nor U7098 (N_7098,N_2922,N_3850);
and U7099 (N_7099,N_4470,N_3674);
nand U7100 (N_7100,N_2800,N_3246);
or U7101 (N_7101,N_4921,N_3069);
or U7102 (N_7102,N_3054,N_3852);
or U7103 (N_7103,N_4778,N_4107);
nor U7104 (N_7104,N_4422,N_3038);
nand U7105 (N_7105,N_2501,N_3646);
or U7106 (N_7106,N_3951,N_4463);
nand U7107 (N_7107,N_4090,N_3954);
nor U7108 (N_7108,N_3081,N_4716);
or U7109 (N_7109,N_4224,N_2505);
and U7110 (N_7110,N_3175,N_3109);
nor U7111 (N_7111,N_4968,N_4664);
or U7112 (N_7112,N_4087,N_3662);
and U7113 (N_7113,N_4610,N_4666);
nand U7114 (N_7114,N_3524,N_4345);
nor U7115 (N_7115,N_4955,N_3180);
nand U7116 (N_7116,N_3836,N_4290);
or U7117 (N_7117,N_2663,N_2520);
or U7118 (N_7118,N_3337,N_4431);
nand U7119 (N_7119,N_4472,N_3447);
nor U7120 (N_7120,N_2573,N_4090);
nor U7121 (N_7121,N_4784,N_2896);
nand U7122 (N_7122,N_3959,N_3815);
or U7123 (N_7123,N_4678,N_2542);
nand U7124 (N_7124,N_3668,N_3018);
nand U7125 (N_7125,N_2960,N_3163);
nor U7126 (N_7126,N_2734,N_2590);
nand U7127 (N_7127,N_3850,N_3019);
nand U7128 (N_7128,N_3999,N_4641);
and U7129 (N_7129,N_3689,N_3306);
nor U7130 (N_7130,N_3129,N_4513);
nand U7131 (N_7131,N_2855,N_3324);
nor U7132 (N_7132,N_3316,N_2677);
and U7133 (N_7133,N_4845,N_3186);
nand U7134 (N_7134,N_3166,N_2687);
nand U7135 (N_7135,N_4641,N_3438);
or U7136 (N_7136,N_4121,N_4321);
nand U7137 (N_7137,N_4832,N_4131);
and U7138 (N_7138,N_4978,N_3670);
and U7139 (N_7139,N_4377,N_3059);
nor U7140 (N_7140,N_4539,N_4795);
xor U7141 (N_7141,N_3232,N_3888);
or U7142 (N_7142,N_3082,N_4707);
nor U7143 (N_7143,N_4893,N_2745);
nand U7144 (N_7144,N_3840,N_2710);
nor U7145 (N_7145,N_4468,N_3311);
nor U7146 (N_7146,N_3277,N_3835);
or U7147 (N_7147,N_4553,N_4073);
or U7148 (N_7148,N_4817,N_4088);
nand U7149 (N_7149,N_3335,N_4468);
and U7150 (N_7150,N_4076,N_2995);
nand U7151 (N_7151,N_4364,N_3810);
or U7152 (N_7152,N_4040,N_4343);
or U7153 (N_7153,N_2675,N_2868);
or U7154 (N_7154,N_3086,N_3316);
and U7155 (N_7155,N_3185,N_4945);
nand U7156 (N_7156,N_4292,N_4548);
and U7157 (N_7157,N_2903,N_3808);
nor U7158 (N_7158,N_2509,N_3138);
xnor U7159 (N_7159,N_2849,N_3595);
or U7160 (N_7160,N_4370,N_3268);
and U7161 (N_7161,N_2681,N_2848);
or U7162 (N_7162,N_3827,N_2652);
nand U7163 (N_7163,N_2859,N_2800);
or U7164 (N_7164,N_4178,N_4404);
xor U7165 (N_7165,N_2528,N_4897);
and U7166 (N_7166,N_3474,N_4344);
and U7167 (N_7167,N_4032,N_4108);
nor U7168 (N_7168,N_4062,N_3429);
or U7169 (N_7169,N_3137,N_3736);
nand U7170 (N_7170,N_2824,N_4608);
nand U7171 (N_7171,N_4193,N_3633);
or U7172 (N_7172,N_2894,N_3045);
nor U7173 (N_7173,N_4407,N_3695);
or U7174 (N_7174,N_4589,N_3470);
or U7175 (N_7175,N_4628,N_3137);
nand U7176 (N_7176,N_3801,N_3186);
and U7177 (N_7177,N_4477,N_4732);
xnor U7178 (N_7178,N_3056,N_3448);
nand U7179 (N_7179,N_3918,N_3611);
nand U7180 (N_7180,N_4149,N_4371);
and U7181 (N_7181,N_3740,N_4388);
nor U7182 (N_7182,N_3652,N_3780);
or U7183 (N_7183,N_3898,N_4918);
and U7184 (N_7184,N_3926,N_4435);
nor U7185 (N_7185,N_3957,N_2537);
nor U7186 (N_7186,N_3936,N_4866);
nand U7187 (N_7187,N_4074,N_3663);
nand U7188 (N_7188,N_4609,N_3276);
nor U7189 (N_7189,N_2730,N_3201);
or U7190 (N_7190,N_4748,N_3809);
nor U7191 (N_7191,N_4519,N_3072);
nand U7192 (N_7192,N_2730,N_2594);
nand U7193 (N_7193,N_3196,N_4314);
nor U7194 (N_7194,N_3394,N_3549);
nor U7195 (N_7195,N_2526,N_3399);
or U7196 (N_7196,N_3254,N_4240);
and U7197 (N_7197,N_3433,N_2686);
nor U7198 (N_7198,N_3744,N_4660);
xor U7199 (N_7199,N_4684,N_2571);
nand U7200 (N_7200,N_4065,N_3069);
nor U7201 (N_7201,N_2689,N_2978);
xor U7202 (N_7202,N_4499,N_3987);
or U7203 (N_7203,N_3669,N_3172);
nor U7204 (N_7204,N_4104,N_4822);
and U7205 (N_7205,N_2674,N_4936);
or U7206 (N_7206,N_3714,N_3982);
or U7207 (N_7207,N_3506,N_3195);
and U7208 (N_7208,N_4086,N_2910);
or U7209 (N_7209,N_4245,N_4919);
nand U7210 (N_7210,N_4907,N_2659);
nor U7211 (N_7211,N_3771,N_3109);
xor U7212 (N_7212,N_2777,N_4893);
or U7213 (N_7213,N_3717,N_4341);
nor U7214 (N_7214,N_4335,N_4128);
nor U7215 (N_7215,N_3208,N_3729);
and U7216 (N_7216,N_2637,N_3218);
nand U7217 (N_7217,N_2736,N_4246);
nand U7218 (N_7218,N_4568,N_2674);
and U7219 (N_7219,N_4552,N_3459);
and U7220 (N_7220,N_3216,N_3621);
nand U7221 (N_7221,N_3693,N_4863);
and U7222 (N_7222,N_4620,N_3686);
or U7223 (N_7223,N_4438,N_2853);
xnor U7224 (N_7224,N_3666,N_2541);
and U7225 (N_7225,N_3903,N_4902);
nand U7226 (N_7226,N_4287,N_3220);
and U7227 (N_7227,N_2982,N_3400);
xor U7228 (N_7228,N_4534,N_3594);
nand U7229 (N_7229,N_2912,N_4342);
and U7230 (N_7230,N_4657,N_3392);
nand U7231 (N_7231,N_3367,N_2544);
nand U7232 (N_7232,N_2542,N_3159);
nand U7233 (N_7233,N_3152,N_2827);
and U7234 (N_7234,N_2654,N_4520);
and U7235 (N_7235,N_3335,N_3426);
nand U7236 (N_7236,N_4543,N_3287);
nor U7237 (N_7237,N_4193,N_2567);
or U7238 (N_7238,N_2871,N_3587);
nand U7239 (N_7239,N_4983,N_4797);
nor U7240 (N_7240,N_3685,N_2766);
nor U7241 (N_7241,N_3102,N_3834);
nand U7242 (N_7242,N_2756,N_2901);
xor U7243 (N_7243,N_3614,N_3973);
or U7244 (N_7244,N_3099,N_3183);
or U7245 (N_7245,N_2537,N_2744);
and U7246 (N_7246,N_4603,N_4329);
nor U7247 (N_7247,N_2568,N_3216);
nand U7248 (N_7248,N_4886,N_3445);
and U7249 (N_7249,N_3268,N_3994);
nor U7250 (N_7250,N_4430,N_4069);
and U7251 (N_7251,N_4816,N_2722);
or U7252 (N_7252,N_2572,N_2612);
or U7253 (N_7253,N_4874,N_3860);
nor U7254 (N_7254,N_3285,N_2613);
nor U7255 (N_7255,N_2897,N_3203);
xnor U7256 (N_7256,N_3148,N_2943);
nand U7257 (N_7257,N_3315,N_4657);
or U7258 (N_7258,N_4631,N_3459);
nand U7259 (N_7259,N_3975,N_2568);
and U7260 (N_7260,N_4640,N_4438);
nor U7261 (N_7261,N_3617,N_2712);
nand U7262 (N_7262,N_3154,N_4470);
or U7263 (N_7263,N_4615,N_3601);
or U7264 (N_7264,N_3423,N_4392);
or U7265 (N_7265,N_4366,N_2571);
nor U7266 (N_7266,N_3802,N_2835);
or U7267 (N_7267,N_4497,N_3639);
nand U7268 (N_7268,N_3178,N_3576);
and U7269 (N_7269,N_4135,N_4157);
and U7270 (N_7270,N_3480,N_4065);
nand U7271 (N_7271,N_2777,N_3356);
nor U7272 (N_7272,N_2953,N_3876);
nor U7273 (N_7273,N_3926,N_3427);
or U7274 (N_7274,N_3344,N_4088);
nand U7275 (N_7275,N_3823,N_2574);
nor U7276 (N_7276,N_4618,N_3611);
or U7277 (N_7277,N_2582,N_4561);
nor U7278 (N_7278,N_2583,N_2826);
nor U7279 (N_7279,N_2621,N_3620);
and U7280 (N_7280,N_2550,N_3665);
nand U7281 (N_7281,N_4611,N_3853);
and U7282 (N_7282,N_4253,N_4197);
nand U7283 (N_7283,N_4520,N_2559);
nor U7284 (N_7284,N_4819,N_3584);
and U7285 (N_7285,N_3579,N_3099);
nand U7286 (N_7286,N_3363,N_4118);
nor U7287 (N_7287,N_4916,N_4704);
or U7288 (N_7288,N_4049,N_3468);
and U7289 (N_7289,N_4963,N_3077);
nor U7290 (N_7290,N_4554,N_2710);
nand U7291 (N_7291,N_4259,N_3417);
nand U7292 (N_7292,N_3093,N_2750);
or U7293 (N_7293,N_3297,N_4866);
and U7294 (N_7294,N_3413,N_2803);
nand U7295 (N_7295,N_3409,N_3944);
nand U7296 (N_7296,N_3861,N_2522);
or U7297 (N_7297,N_4083,N_4376);
or U7298 (N_7298,N_2701,N_3978);
nor U7299 (N_7299,N_4326,N_4429);
nor U7300 (N_7300,N_2792,N_3285);
nand U7301 (N_7301,N_3454,N_3324);
or U7302 (N_7302,N_4472,N_4909);
and U7303 (N_7303,N_2768,N_3798);
nand U7304 (N_7304,N_4372,N_2800);
nand U7305 (N_7305,N_4634,N_3356);
and U7306 (N_7306,N_4622,N_4338);
nor U7307 (N_7307,N_2529,N_3635);
or U7308 (N_7308,N_2573,N_3682);
nor U7309 (N_7309,N_2616,N_4770);
nand U7310 (N_7310,N_4147,N_3161);
nor U7311 (N_7311,N_4563,N_3239);
nor U7312 (N_7312,N_4224,N_2577);
and U7313 (N_7313,N_4508,N_4944);
nor U7314 (N_7314,N_4305,N_2510);
nor U7315 (N_7315,N_4238,N_3495);
nor U7316 (N_7316,N_3312,N_4044);
nor U7317 (N_7317,N_3166,N_4078);
and U7318 (N_7318,N_4941,N_4729);
or U7319 (N_7319,N_2572,N_4576);
nand U7320 (N_7320,N_3826,N_3709);
and U7321 (N_7321,N_2934,N_4545);
and U7322 (N_7322,N_4624,N_4111);
nor U7323 (N_7323,N_2800,N_3896);
and U7324 (N_7324,N_4530,N_4047);
or U7325 (N_7325,N_4155,N_2998);
and U7326 (N_7326,N_4132,N_4386);
and U7327 (N_7327,N_2504,N_4935);
nand U7328 (N_7328,N_3790,N_3671);
nor U7329 (N_7329,N_3817,N_3455);
nor U7330 (N_7330,N_4580,N_2987);
nor U7331 (N_7331,N_4725,N_3851);
and U7332 (N_7332,N_3343,N_4527);
or U7333 (N_7333,N_3403,N_3175);
xor U7334 (N_7334,N_3222,N_3709);
nand U7335 (N_7335,N_4032,N_3253);
and U7336 (N_7336,N_4874,N_3326);
or U7337 (N_7337,N_4827,N_3512);
and U7338 (N_7338,N_4880,N_3060);
nand U7339 (N_7339,N_4164,N_4255);
or U7340 (N_7340,N_2638,N_2538);
nand U7341 (N_7341,N_4145,N_2583);
and U7342 (N_7342,N_2978,N_2970);
xnor U7343 (N_7343,N_4456,N_2892);
or U7344 (N_7344,N_2707,N_3078);
nor U7345 (N_7345,N_2629,N_3389);
and U7346 (N_7346,N_4654,N_4877);
nor U7347 (N_7347,N_4472,N_3842);
and U7348 (N_7348,N_3174,N_2813);
or U7349 (N_7349,N_3476,N_3454);
nor U7350 (N_7350,N_2508,N_3392);
nor U7351 (N_7351,N_4539,N_4178);
nand U7352 (N_7352,N_2503,N_2956);
nor U7353 (N_7353,N_3113,N_2684);
nor U7354 (N_7354,N_4383,N_4212);
or U7355 (N_7355,N_3300,N_2506);
and U7356 (N_7356,N_2712,N_3907);
nand U7357 (N_7357,N_3914,N_3270);
or U7358 (N_7358,N_3161,N_2842);
and U7359 (N_7359,N_2531,N_3903);
nand U7360 (N_7360,N_4864,N_3214);
and U7361 (N_7361,N_2517,N_4736);
or U7362 (N_7362,N_2506,N_4758);
nand U7363 (N_7363,N_4678,N_3533);
or U7364 (N_7364,N_3122,N_2768);
nand U7365 (N_7365,N_4683,N_4283);
or U7366 (N_7366,N_3753,N_3782);
or U7367 (N_7367,N_2573,N_2514);
and U7368 (N_7368,N_3271,N_2595);
nand U7369 (N_7369,N_3445,N_3572);
and U7370 (N_7370,N_3407,N_4173);
nand U7371 (N_7371,N_3273,N_4622);
nor U7372 (N_7372,N_3194,N_4586);
nand U7373 (N_7373,N_4463,N_4079);
and U7374 (N_7374,N_4575,N_4374);
and U7375 (N_7375,N_4419,N_2907);
and U7376 (N_7376,N_3964,N_4820);
nor U7377 (N_7377,N_3262,N_3154);
nor U7378 (N_7378,N_3978,N_4156);
nand U7379 (N_7379,N_3658,N_4291);
nor U7380 (N_7380,N_3146,N_2884);
nand U7381 (N_7381,N_3618,N_3544);
nor U7382 (N_7382,N_4273,N_4457);
and U7383 (N_7383,N_4889,N_3952);
or U7384 (N_7384,N_4742,N_2985);
nor U7385 (N_7385,N_4660,N_4390);
nor U7386 (N_7386,N_4406,N_3065);
and U7387 (N_7387,N_4947,N_4128);
or U7388 (N_7388,N_4183,N_4083);
or U7389 (N_7389,N_3332,N_4647);
or U7390 (N_7390,N_2961,N_3406);
xnor U7391 (N_7391,N_4956,N_3894);
or U7392 (N_7392,N_4264,N_4439);
xnor U7393 (N_7393,N_3384,N_4570);
nor U7394 (N_7394,N_4332,N_3796);
nor U7395 (N_7395,N_4744,N_3092);
or U7396 (N_7396,N_4718,N_2564);
nor U7397 (N_7397,N_3449,N_4186);
or U7398 (N_7398,N_4912,N_4694);
nand U7399 (N_7399,N_2915,N_2941);
nand U7400 (N_7400,N_4738,N_3667);
or U7401 (N_7401,N_3426,N_2535);
and U7402 (N_7402,N_3406,N_4079);
or U7403 (N_7403,N_4513,N_3141);
or U7404 (N_7404,N_3559,N_2732);
nor U7405 (N_7405,N_2969,N_2977);
nor U7406 (N_7406,N_4236,N_3029);
and U7407 (N_7407,N_2838,N_4859);
and U7408 (N_7408,N_4992,N_4571);
nor U7409 (N_7409,N_3485,N_3849);
and U7410 (N_7410,N_4332,N_4006);
nor U7411 (N_7411,N_3949,N_4160);
nand U7412 (N_7412,N_2608,N_3113);
nor U7413 (N_7413,N_4508,N_2971);
nand U7414 (N_7414,N_4997,N_4717);
and U7415 (N_7415,N_3958,N_3493);
and U7416 (N_7416,N_4707,N_3001);
or U7417 (N_7417,N_3068,N_2532);
nor U7418 (N_7418,N_4245,N_3135);
or U7419 (N_7419,N_3556,N_2589);
and U7420 (N_7420,N_4774,N_3610);
nor U7421 (N_7421,N_2944,N_3968);
nand U7422 (N_7422,N_4664,N_3194);
nand U7423 (N_7423,N_4032,N_4383);
and U7424 (N_7424,N_4029,N_3600);
nand U7425 (N_7425,N_4342,N_2879);
nor U7426 (N_7426,N_2507,N_2990);
nor U7427 (N_7427,N_2725,N_3986);
and U7428 (N_7428,N_4486,N_2974);
nand U7429 (N_7429,N_3827,N_3915);
nor U7430 (N_7430,N_4983,N_2831);
and U7431 (N_7431,N_4655,N_3485);
nand U7432 (N_7432,N_3495,N_4305);
and U7433 (N_7433,N_2706,N_2516);
nor U7434 (N_7434,N_3330,N_2899);
nor U7435 (N_7435,N_3533,N_4472);
nand U7436 (N_7436,N_4092,N_2755);
nand U7437 (N_7437,N_4095,N_3531);
nand U7438 (N_7438,N_4873,N_3147);
or U7439 (N_7439,N_4714,N_2824);
and U7440 (N_7440,N_3123,N_4078);
nor U7441 (N_7441,N_2572,N_3642);
nand U7442 (N_7442,N_3501,N_3368);
or U7443 (N_7443,N_4353,N_3132);
nand U7444 (N_7444,N_4221,N_2974);
and U7445 (N_7445,N_4583,N_3867);
nor U7446 (N_7446,N_3366,N_2594);
nor U7447 (N_7447,N_4119,N_2974);
and U7448 (N_7448,N_4229,N_4385);
and U7449 (N_7449,N_3434,N_4611);
nor U7450 (N_7450,N_3036,N_4710);
and U7451 (N_7451,N_3525,N_3790);
and U7452 (N_7452,N_4798,N_4809);
nor U7453 (N_7453,N_3523,N_4705);
and U7454 (N_7454,N_4202,N_2507);
or U7455 (N_7455,N_2982,N_3227);
xnor U7456 (N_7456,N_4910,N_4897);
and U7457 (N_7457,N_4456,N_2752);
and U7458 (N_7458,N_4789,N_4432);
nand U7459 (N_7459,N_2581,N_4412);
nor U7460 (N_7460,N_3743,N_4483);
nor U7461 (N_7461,N_3401,N_4470);
nor U7462 (N_7462,N_2858,N_2756);
xnor U7463 (N_7463,N_4085,N_2552);
nor U7464 (N_7464,N_3544,N_2862);
xor U7465 (N_7465,N_3672,N_3283);
or U7466 (N_7466,N_4068,N_4733);
nor U7467 (N_7467,N_4788,N_2976);
and U7468 (N_7468,N_3235,N_3673);
nand U7469 (N_7469,N_4016,N_4123);
and U7470 (N_7470,N_3232,N_3760);
nor U7471 (N_7471,N_4102,N_2561);
nor U7472 (N_7472,N_2915,N_3372);
or U7473 (N_7473,N_3434,N_2669);
nand U7474 (N_7474,N_3934,N_3610);
nand U7475 (N_7475,N_3418,N_3946);
nor U7476 (N_7476,N_4578,N_4344);
nor U7477 (N_7477,N_4634,N_4251);
or U7478 (N_7478,N_3935,N_4976);
nor U7479 (N_7479,N_4724,N_3052);
nor U7480 (N_7480,N_3415,N_3566);
nor U7481 (N_7481,N_2666,N_3336);
nor U7482 (N_7482,N_3944,N_4937);
or U7483 (N_7483,N_3065,N_3264);
or U7484 (N_7484,N_4490,N_4563);
or U7485 (N_7485,N_4130,N_3019);
or U7486 (N_7486,N_3876,N_4305);
nand U7487 (N_7487,N_2868,N_2722);
nor U7488 (N_7488,N_4364,N_4686);
and U7489 (N_7489,N_2775,N_3331);
or U7490 (N_7490,N_4546,N_4928);
nor U7491 (N_7491,N_4562,N_4590);
nand U7492 (N_7492,N_2612,N_3887);
or U7493 (N_7493,N_3613,N_2586);
nor U7494 (N_7494,N_4729,N_4804);
nand U7495 (N_7495,N_2697,N_3373);
nand U7496 (N_7496,N_3609,N_2830);
nand U7497 (N_7497,N_4033,N_2958);
nand U7498 (N_7498,N_4592,N_3438);
nand U7499 (N_7499,N_4374,N_4166);
nand U7500 (N_7500,N_5528,N_6581);
and U7501 (N_7501,N_6786,N_5152);
and U7502 (N_7502,N_5042,N_5177);
or U7503 (N_7503,N_7195,N_5360);
or U7504 (N_7504,N_6810,N_7458);
or U7505 (N_7505,N_7491,N_6811);
and U7506 (N_7506,N_5405,N_5126);
or U7507 (N_7507,N_6593,N_5967);
nor U7508 (N_7508,N_7386,N_6288);
nand U7509 (N_7509,N_5899,N_6353);
nand U7510 (N_7510,N_7354,N_5088);
xor U7511 (N_7511,N_5020,N_5320);
nand U7512 (N_7512,N_6013,N_6741);
xor U7513 (N_7513,N_6592,N_7336);
nand U7514 (N_7514,N_7142,N_7008);
and U7515 (N_7515,N_7042,N_6924);
nor U7516 (N_7516,N_5745,N_6470);
and U7517 (N_7517,N_7229,N_5366);
and U7518 (N_7518,N_6688,N_6823);
or U7519 (N_7519,N_7120,N_6402);
and U7520 (N_7520,N_6467,N_6956);
and U7521 (N_7521,N_6083,N_5499);
nand U7522 (N_7522,N_5246,N_5440);
nor U7523 (N_7523,N_5759,N_6619);
or U7524 (N_7524,N_7198,N_7216);
xor U7525 (N_7525,N_6701,N_5812);
or U7526 (N_7526,N_5969,N_5615);
or U7527 (N_7527,N_7275,N_6175);
or U7528 (N_7528,N_5199,N_6395);
nand U7529 (N_7529,N_5879,N_6066);
nand U7530 (N_7530,N_6416,N_6559);
and U7531 (N_7531,N_6617,N_5546);
nor U7532 (N_7532,N_6829,N_5724);
and U7533 (N_7533,N_6469,N_5106);
nor U7534 (N_7534,N_6366,N_5941);
nor U7535 (N_7535,N_5913,N_6448);
or U7536 (N_7536,N_6174,N_6704);
nor U7537 (N_7537,N_6020,N_6135);
nor U7538 (N_7538,N_7424,N_5992);
nor U7539 (N_7539,N_7103,N_6892);
nand U7540 (N_7540,N_5704,N_6106);
nor U7541 (N_7541,N_5024,N_6797);
or U7542 (N_7542,N_7166,N_7095);
nor U7543 (N_7543,N_6684,N_5515);
nand U7544 (N_7544,N_7334,N_5858);
nand U7545 (N_7545,N_6143,N_5776);
or U7546 (N_7546,N_5131,N_7309);
and U7547 (N_7547,N_6382,N_5504);
or U7548 (N_7548,N_6224,N_6550);
or U7549 (N_7549,N_6530,N_5685);
or U7550 (N_7550,N_5006,N_6299);
nand U7551 (N_7551,N_5471,N_5094);
nor U7552 (N_7552,N_5894,N_5557);
nor U7553 (N_7553,N_5313,N_7190);
or U7554 (N_7554,N_6354,N_5204);
nor U7555 (N_7555,N_6942,N_5775);
or U7556 (N_7556,N_6739,N_6386);
nor U7557 (N_7557,N_6928,N_6677);
and U7558 (N_7558,N_5781,N_5558);
nor U7559 (N_7559,N_6180,N_7163);
nor U7560 (N_7560,N_5149,N_5358);
or U7561 (N_7561,N_6052,N_7050);
nand U7562 (N_7562,N_6358,N_7063);
and U7563 (N_7563,N_5770,N_6290);
nand U7564 (N_7564,N_5439,N_7387);
nor U7565 (N_7565,N_7033,N_6461);
and U7566 (N_7566,N_6912,N_5034);
nand U7567 (N_7567,N_5295,N_6867);
and U7568 (N_7568,N_5093,N_6221);
and U7569 (N_7569,N_6766,N_5133);
and U7570 (N_7570,N_5999,N_6310);
and U7571 (N_7571,N_6447,N_5814);
or U7572 (N_7572,N_7162,N_5019);
or U7573 (N_7573,N_7367,N_5827);
nand U7574 (N_7574,N_6239,N_5336);
and U7575 (N_7575,N_5262,N_5198);
nand U7576 (N_7576,N_6674,N_6501);
nand U7577 (N_7577,N_7277,N_5587);
and U7578 (N_7578,N_5692,N_5092);
or U7579 (N_7579,N_6226,N_5514);
and U7580 (N_7580,N_6838,N_6654);
xnor U7581 (N_7581,N_7028,N_5064);
nor U7582 (N_7582,N_5965,N_7327);
and U7583 (N_7583,N_5771,N_6517);
or U7584 (N_7584,N_7058,N_5889);
or U7585 (N_7585,N_5872,N_5184);
and U7586 (N_7586,N_6736,N_7441);
or U7587 (N_7587,N_6719,N_7391);
nor U7588 (N_7588,N_5304,N_6995);
nand U7589 (N_7589,N_6064,N_7023);
nand U7590 (N_7590,N_7171,N_5936);
and U7591 (N_7591,N_5312,N_5388);
nor U7592 (N_7592,N_7179,N_5179);
nor U7593 (N_7593,N_6352,N_6601);
or U7594 (N_7594,N_7081,N_5297);
or U7595 (N_7595,N_6259,N_5810);
nand U7596 (N_7596,N_7437,N_6332);
and U7597 (N_7597,N_5221,N_6941);
and U7598 (N_7598,N_5037,N_6128);
xor U7599 (N_7599,N_6877,N_5891);
nand U7600 (N_7600,N_6258,N_5933);
nand U7601 (N_7601,N_7268,N_5361);
nor U7602 (N_7602,N_6820,N_6391);
or U7603 (N_7603,N_5616,N_6666);
or U7604 (N_7604,N_7046,N_7300);
nand U7605 (N_7605,N_5063,N_5916);
and U7606 (N_7606,N_5857,N_6051);
and U7607 (N_7607,N_6513,N_6854);
nor U7608 (N_7608,N_5637,N_7127);
nor U7609 (N_7609,N_5736,N_7359);
or U7610 (N_7610,N_5619,N_5680);
and U7611 (N_7611,N_7496,N_7096);
nand U7612 (N_7612,N_6860,N_5247);
nand U7613 (N_7613,N_6998,N_5472);
and U7614 (N_7614,N_6847,N_6283);
or U7615 (N_7615,N_6050,N_7168);
nand U7616 (N_7616,N_5169,N_7237);
nor U7617 (N_7617,N_6451,N_6648);
nand U7618 (N_7618,N_5245,N_7251);
nand U7619 (N_7619,N_6527,N_5143);
and U7620 (N_7620,N_7094,N_7423);
nor U7621 (N_7621,N_6111,N_5929);
or U7622 (N_7622,N_5105,N_5310);
nand U7623 (N_7623,N_6148,N_6405);
and U7624 (N_7624,N_6409,N_5322);
nand U7625 (N_7625,N_5720,N_7269);
and U7626 (N_7626,N_5255,N_6240);
nand U7627 (N_7627,N_7146,N_6801);
and U7628 (N_7628,N_7206,N_5280);
and U7629 (N_7629,N_6965,N_5442);
and U7630 (N_7630,N_5039,N_7427);
nand U7631 (N_7631,N_7291,N_5666);
and U7632 (N_7632,N_7211,N_6529);
or U7633 (N_7633,N_6579,N_5686);
or U7634 (N_7634,N_7485,N_7201);
nand U7635 (N_7635,N_6782,N_6967);
and U7636 (N_7636,N_7410,N_5743);
or U7637 (N_7637,N_5506,N_6557);
nand U7638 (N_7638,N_6977,N_5520);
or U7639 (N_7639,N_6113,N_6444);
or U7640 (N_7640,N_6843,N_5017);
nand U7641 (N_7641,N_6780,N_5387);
nor U7642 (N_7642,N_7435,N_7452);
nand U7643 (N_7643,N_5645,N_6993);
and U7644 (N_7644,N_5355,N_6558);
nand U7645 (N_7645,N_6958,N_6039);
nor U7646 (N_7646,N_5371,N_5987);
nor U7647 (N_7647,N_5309,N_7199);
and U7648 (N_7648,N_6777,N_6563);
nand U7649 (N_7649,N_7134,N_6693);
nor U7650 (N_7650,N_5729,N_6207);
or U7651 (N_7651,N_7341,N_5918);
nand U7652 (N_7652,N_6269,N_6033);
and U7653 (N_7653,N_6551,N_5582);
nor U7654 (N_7654,N_5817,N_5267);
or U7655 (N_7655,N_5127,N_7202);
or U7656 (N_7656,N_5239,N_7383);
nand U7657 (N_7657,N_6538,N_6828);
nor U7658 (N_7658,N_5335,N_5279);
nand U7659 (N_7659,N_5290,N_6954);
and U7660 (N_7660,N_6936,N_5975);
or U7661 (N_7661,N_7151,N_5406);
nand U7662 (N_7662,N_6154,N_6479);
or U7663 (N_7663,N_5910,N_5240);
and U7664 (N_7664,N_6534,N_5517);
and U7665 (N_7665,N_5481,N_5624);
or U7666 (N_7666,N_5809,N_5136);
or U7667 (N_7667,N_6834,N_5964);
and U7668 (N_7668,N_5154,N_6940);
nand U7669 (N_7669,N_5926,N_6301);
and U7670 (N_7670,N_5993,N_5328);
nand U7671 (N_7671,N_6464,N_6276);
or U7672 (N_7672,N_5639,N_6983);
and U7673 (N_7673,N_6398,N_6548);
and U7674 (N_7674,N_7082,N_6699);
or U7675 (N_7675,N_5047,N_6636);
or U7676 (N_7676,N_5458,N_6404);
or U7677 (N_7677,N_5392,N_6496);
xor U7678 (N_7678,N_5753,N_6193);
and U7679 (N_7679,N_7333,N_6880);
and U7680 (N_7680,N_6788,N_5207);
nor U7681 (N_7681,N_6562,N_5241);
or U7682 (N_7682,N_5353,N_6298);
or U7683 (N_7683,N_7080,N_6652);
and U7684 (N_7684,N_5869,N_6795);
nor U7685 (N_7685,N_6508,N_6225);
nand U7686 (N_7686,N_5605,N_6709);
or U7687 (N_7687,N_6974,N_7343);
nand U7688 (N_7688,N_7144,N_5176);
nor U7689 (N_7689,N_5762,N_5836);
nand U7690 (N_7690,N_5691,N_6914);
or U7691 (N_7691,N_7061,N_7394);
and U7692 (N_7692,N_5760,N_5581);
and U7693 (N_7693,N_7018,N_6690);
nor U7694 (N_7694,N_6104,N_5378);
or U7695 (N_7695,N_7234,N_6753);
or U7696 (N_7696,N_6089,N_5300);
nor U7697 (N_7697,N_7426,N_5072);
or U7698 (N_7698,N_6884,N_7246);
nor U7699 (N_7699,N_5892,N_6403);
nand U7700 (N_7700,N_5303,N_5139);
nand U7701 (N_7701,N_6608,N_6771);
and U7702 (N_7702,N_5804,N_7340);
or U7703 (N_7703,N_7389,N_5235);
and U7704 (N_7704,N_5545,N_5174);
nand U7705 (N_7705,N_7167,N_5757);
nor U7706 (N_7706,N_5167,N_6500);
or U7707 (N_7707,N_6157,N_5798);
and U7708 (N_7708,N_6026,N_5877);
and U7709 (N_7709,N_7363,N_6660);
or U7710 (N_7710,N_7401,N_7479);
or U7711 (N_7711,N_6244,N_7013);
or U7712 (N_7712,N_6155,N_6726);
or U7713 (N_7713,N_6742,N_5706);
or U7714 (N_7714,N_6948,N_6599);
nand U7715 (N_7715,N_5001,N_5601);
and U7716 (N_7716,N_5473,N_5079);
and U7717 (N_7717,N_6605,N_6423);
and U7718 (N_7718,N_6432,N_5219);
nand U7719 (N_7719,N_5140,N_5432);
nor U7720 (N_7720,N_7481,N_6274);
and U7721 (N_7721,N_6511,N_6337);
nand U7722 (N_7722,N_5529,N_6308);
or U7723 (N_7723,N_7484,N_5652);
or U7724 (N_7724,N_5409,N_6700);
and U7725 (N_7725,N_7271,N_6161);
and U7726 (N_7726,N_5159,N_7430);
or U7727 (N_7727,N_7009,N_5888);
and U7728 (N_7728,N_6902,N_5566);
nand U7729 (N_7729,N_6925,N_6431);
nor U7730 (N_7730,N_6058,N_5045);
nand U7731 (N_7731,N_6278,N_6037);
or U7732 (N_7732,N_5043,N_5611);
and U7733 (N_7733,N_6393,N_6082);
nor U7734 (N_7734,N_6465,N_7098);
nand U7735 (N_7735,N_5897,N_6979);
and U7736 (N_7736,N_6566,N_6069);
and U7737 (N_7737,N_6072,N_5739);
and U7738 (N_7738,N_5732,N_7468);
nand U7739 (N_7739,N_6628,N_6865);
or U7740 (N_7740,N_5026,N_6759);
or U7741 (N_7741,N_6851,N_5486);
or U7742 (N_7742,N_6573,N_6126);
nand U7743 (N_7743,N_5530,N_6241);
and U7744 (N_7744,N_6687,N_6356);
or U7745 (N_7745,N_5098,N_5447);
xor U7746 (N_7746,N_6179,N_6891);
nand U7747 (N_7747,N_7360,N_6105);
nor U7748 (N_7748,N_7257,N_6091);
nor U7749 (N_7749,N_7345,N_5596);
nor U7750 (N_7750,N_7175,N_5828);
nor U7751 (N_7751,N_6365,N_7026);
nor U7752 (N_7752,N_5233,N_7362);
nor U7753 (N_7753,N_6063,N_5062);
nor U7754 (N_7754,N_5172,N_7284);
nor U7755 (N_7755,N_6540,N_5912);
nor U7756 (N_7756,N_5166,N_5423);
nor U7757 (N_7757,N_5697,N_5029);
nand U7758 (N_7758,N_5232,N_5007);
or U7759 (N_7759,N_5372,N_6888);
or U7760 (N_7760,N_6735,N_6515);
nand U7761 (N_7761,N_5212,N_7224);
nor U7762 (N_7762,N_6057,N_6307);
nand U7763 (N_7763,N_6053,N_6947);
nor U7764 (N_7764,N_7226,N_7358);
nand U7765 (N_7765,N_5324,N_6195);
nand U7766 (N_7766,N_6714,N_6087);
or U7767 (N_7767,N_6476,N_7370);
and U7768 (N_7768,N_5206,N_6908);
and U7769 (N_7769,N_5583,N_5896);
nand U7770 (N_7770,N_6981,N_5483);
nand U7771 (N_7771,N_7270,N_6176);
and U7772 (N_7772,N_5868,N_6672);
nor U7773 (N_7773,N_7433,N_7073);
or U7774 (N_7774,N_7189,N_6554);
or U7775 (N_7775,N_5285,N_5027);
and U7776 (N_7776,N_7411,N_7302);
nand U7777 (N_7777,N_5971,N_5821);
or U7778 (N_7778,N_7003,N_5469);
or U7779 (N_7779,N_6305,N_6659);
or U7780 (N_7780,N_6863,N_5428);
and U7781 (N_7781,N_5038,N_5947);
nor U7782 (N_7782,N_6637,N_5348);
nor U7783 (N_7783,N_5180,N_6133);
nor U7784 (N_7784,N_7139,N_5939);
and U7785 (N_7785,N_7316,N_7417);
nand U7786 (N_7786,N_5989,N_6325);
or U7787 (N_7787,N_6896,N_6320);
xor U7788 (N_7788,N_6282,N_5907);
or U7789 (N_7789,N_6218,N_5540);
or U7790 (N_7790,N_5217,N_5973);
nand U7791 (N_7791,N_6616,N_6270);
and U7792 (N_7792,N_7128,N_6236);
nand U7793 (N_7793,N_7295,N_5151);
or U7794 (N_7794,N_7260,N_5856);
nand U7795 (N_7795,N_6591,N_7222);
and U7796 (N_7796,N_6852,N_6080);
nand U7797 (N_7797,N_7005,N_5049);
nor U7798 (N_7798,N_7380,N_6638);
nor U7799 (N_7799,N_5880,N_6302);
nor U7800 (N_7800,N_6519,N_6303);
or U7801 (N_7801,N_5096,N_5460);
nor U7802 (N_7802,N_6696,N_6016);
and U7803 (N_7803,N_5211,N_6446);
nor U7804 (N_7804,N_7010,N_5264);
and U7805 (N_7805,N_5516,N_5002);
nor U7806 (N_7806,N_7322,N_5134);
and U7807 (N_7807,N_5922,N_5044);
nor U7808 (N_7808,N_5824,N_6351);
and U7809 (N_7809,N_7022,N_5494);
xnor U7810 (N_7810,N_6036,N_5751);
nor U7811 (N_7811,N_7407,N_6487);
or U7812 (N_7812,N_5865,N_5847);
nand U7813 (N_7813,N_5925,N_6108);
nor U7814 (N_7814,N_7332,N_7489);
and U7815 (N_7815,N_6243,N_5488);
or U7816 (N_7816,N_6612,N_5915);
nor U7817 (N_7817,N_5153,N_5484);
nor U7818 (N_7818,N_6361,N_5332);
and U7819 (N_7819,N_5905,N_6034);
and U7820 (N_7820,N_6521,N_6440);
nand U7821 (N_7821,N_5369,N_6185);
nor U7822 (N_7822,N_6721,N_6205);
nand U7823 (N_7823,N_6170,N_6065);
and U7824 (N_7824,N_6710,N_5537);
and U7825 (N_7825,N_6043,N_6821);
and U7826 (N_7826,N_6049,N_7111);
and U7827 (N_7827,N_7041,N_5476);
and U7828 (N_7828,N_6536,N_6552);
nor U7829 (N_7829,N_5866,N_6433);
nor U7830 (N_7830,N_5091,N_7155);
nand U7831 (N_7831,N_5761,N_5385);
nand U7832 (N_7832,N_5128,N_5844);
nor U7833 (N_7833,N_7113,N_5287);
and U7834 (N_7834,N_5033,N_7373);
nand U7835 (N_7835,N_7487,N_6056);
nand U7836 (N_7836,N_5025,N_5022);
and U7837 (N_7837,N_6022,N_5725);
and U7838 (N_7838,N_5842,N_7115);
xnor U7839 (N_7839,N_6198,N_6230);
nand U7840 (N_7840,N_7021,N_6632);
nor U7841 (N_7841,N_5508,N_7434);
nand U7842 (N_7842,N_6452,N_5244);
and U7843 (N_7843,N_5884,N_5876);
and U7844 (N_7844,N_6280,N_5521);
and U7845 (N_7845,N_6247,N_6748);
nand U7846 (N_7846,N_7228,N_6492);
and U7847 (N_7847,N_6946,N_5597);
or U7848 (N_7848,N_7196,N_7178);
nor U7849 (N_7849,N_5111,N_6029);
nand U7850 (N_7850,N_6653,N_6856);
and U7851 (N_7851,N_5860,N_6078);
or U7852 (N_7852,N_5782,N_5397);
and U7853 (N_7853,N_6392,N_6328);
and U7854 (N_7854,N_6631,N_7274);
nor U7855 (N_7855,N_6886,N_6943);
nand U7856 (N_7856,N_6061,N_7014);
or U7857 (N_7857,N_5920,N_6643);
nor U7858 (N_7858,N_5323,N_6339);
nand U7859 (N_7859,N_6168,N_5144);
nand U7860 (N_7860,N_7272,N_5855);
and U7861 (N_7861,N_5644,N_6156);
nor U7862 (N_7862,N_7281,N_5364);
xor U7863 (N_7863,N_6134,N_5502);
nand U7864 (N_7864,N_5573,N_6261);
and U7865 (N_7865,N_6397,N_7088);
nor U7866 (N_7866,N_6858,N_6669);
nand U7867 (N_7867,N_5843,N_5393);
xor U7868 (N_7868,N_6761,N_6808);
nor U7869 (N_7869,N_6640,N_7415);
and U7870 (N_7870,N_5069,N_5283);
nand U7871 (N_7871,N_7390,N_5501);
nand U7872 (N_7872,N_7412,N_6215);
or U7873 (N_7873,N_7069,N_7205);
and U7874 (N_7874,N_7244,N_5709);
and U7875 (N_7875,N_5413,N_5742);
nor U7876 (N_7876,N_6642,N_6567);
nand U7877 (N_7877,N_5263,N_6369);
or U7878 (N_7878,N_6260,N_6285);
nor U7879 (N_7879,N_5535,N_6478);
xnor U7880 (N_7880,N_6449,N_6665);
xor U7881 (N_7881,N_6937,N_5946);
and U7882 (N_7882,N_5148,N_5556);
nor U7883 (N_7883,N_7099,N_7482);
xnor U7884 (N_7884,N_5008,N_5259);
and U7885 (N_7885,N_7455,N_5354);
and U7886 (N_7886,N_6149,N_6675);
or U7887 (N_7887,N_5935,N_5617);
and U7888 (N_7888,N_5748,N_5293);
nor U7889 (N_7889,N_6556,N_7393);
and U7890 (N_7890,N_5269,N_6575);
nand U7891 (N_7891,N_6570,N_6312);
nor U7892 (N_7892,N_5851,N_5703);
nand U7893 (N_7893,N_6976,N_7067);
nand U7894 (N_7894,N_6868,N_5383);
nand U7895 (N_7895,N_7293,N_6079);
nor U7896 (N_7896,N_5498,N_6522);
nand U7897 (N_7897,N_7301,N_5822);
and U7898 (N_7898,N_5273,N_7066);
nand U7899 (N_7899,N_6685,N_7121);
and U7900 (N_7900,N_6939,N_7298);
nor U7901 (N_7901,N_5738,N_6035);
and U7902 (N_7902,N_5984,N_7319);
xor U7903 (N_7903,N_7213,N_5667);
nor U7904 (N_7904,N_6495,N_5068);
nor U7905 (N_7905,N_5403,N_6819);
nand U7906 (N_7906,N_5278,N_5115);
nor U7907 (N_7907,N_7068,N_6790);
nor U7908 (N_7908,N_5612,N_5480);
and U7909 (N_7909,N_6263,N_5086);
and U7910 (N_7910,N_6264,N_5189);
nand U7911 (N_7911,N_6614,N_5200);
nor U7912 (N_7912,N_7034,N_5690);
nand U7913 (N_7913,N_7152,N_6773);
nor U7914 (N_7914,N_5630,N_5996);
or U7915 (N_7915,N_7177,N_5023);
and U7916 (N_7916,N_5533,N_6561);
nor U7917 (N_7917,N_7462,N_6765);
nor U7918 (N_7918,N_5650,N_7138);
nand U7919 (N_7919,N_6005,N_5636);
nor U7920 (N_7920,N_7024,N_5839);
and U7921 (N_7921,N_7245,N_5834);
or U7922 (N_7922,N_6737,N_6357);
nand U7923 (N_7923,N_5418,N_6691);
nor U7924 (N_7924,N_6331,N_5150);
nor U7925 (N_7925,N_6641,N_5787);
and U7926 (N_7926,N_6222,N_6295);
xnor U7927 (N_7927,N_5251,N_5252);
and U7928 (N_7928,N_6510,N_5741);
nor U7929 (N_7929,N_6344,N_7065);
or U7930 (N_7930,N_6920,N_6418);
nor U7931 (N_7931,N_6623,N_5818);
nor U7932 (N_7932,N_5651,N_7249);
nor U7933 (N_7933,N_7480,N_7239);
or U7934 (N_7934,N_6122,N_7283);
and U7935 (N_7935,N_6602,N_6103);
nor U7936 (N_7936,N_6438,N_6889);
or U7937 (N_7937,N_7157,N_5945);
and U7938 (N_7938,N_5672,N_5873);
or U7939 (N_7939,N_5988,N_7051);
nand U7940 (N_7940,N_6796,N_7055);
and U7941 (N_7941,N_6480,N_6692);
and U7942 (N_7942,N_5885,N_5223);
nor U7943 (N_7943,N_6070,N_6132);
nor U7944 (N_7944,N_7369,N_6862);
or U7945 (N_7945,N_7338,N_5065);
nor U7946 (N_7946,N_5513,N_5744);
or U7947 (N_7947,N_5800,N_5410);
and U7948 (N_7948,N_7027,N_6102);
and U7949 (N_7949,N_5253,N_6779);
nor U7950 (N_7950,N_7403,N_5379);
and U7951 (N_7951,N_6504,N_6618);
or U7952 (N_7952,N_6147,N_6763);
or U7953 (N_7953,N_5203,N_5076);
or U7954 (N_7954,N_5902,N_6001);
or U7955 (N_7955,N_6425,N_7252);
and U7956 (N_7956,N_6662,N_5503);
nand U7957 (N_7957,N_5389,N_5142);
or U7958 (N_7958,N_5525,N_5914);
xor U7959 (N_7959,N_6262,N_6878);
nand U7960 (N_7960,N_7037,N_6646);
nor U7961 (N_7961,N_6876,N_7215);
and U7962 (N_7962,N_6378,N_7238);
or U7963 (N_7963,N_5934,N_6007);
and U7964 (N_7964,N_7020,N_7477);
and U7965 (N_7965,N_6625,N_7077);
nand U7966 (N_7966,N_7305,N_5077);
or U7967 (N_7967,N_6376,N_5108);
nor U7968 (N_7968,N_7374,N_5436);
nor U7969 (N_7969,N_5845,N_6112);
and U7970 (N_7970,N_6968,N_5549);
or U7971 (N_7971,N_7118,N_6901);
nor U7972 (N_7972,N_6553,N_6927);
nand U7973 (N_7973,N_6966,N_6422);
xor U7974 (N_7974,N_7247,N_6383);
and U7975 (N_7975,N_5437,N_6201);
nor U7976 (N_7976,N_5420,N_6539);
or U7977 (N_7977,N_5979,N_6006);
and U7978 (N_7978,N_6150,N_6749);
and U7979 (N_7979,N_6678,N_6871);
and U7980 (N_7980,N_6384,N_6603);
nor U7981 (N_7981,N_5162,N_6774);
nand U7982 (N_7982,N_6453,N_6297);
or U7983 (N_7983,N_5791,N_6898);
and U7984 (N_7984,N_5548,N_5165);
nand U7985 (N_7985,N_7165,N_7123);
or U7986 (N_7986,N_7158,N_6118);
nand U7987 (N_7987,N_7191,N_5875);
or U7988 (N_7988,N_7255,N_6746);
nor U7989 (N_7989,N_7250,N_7413);
nor U7990 (N_7990,N_5237,N_7308);
nor U7991 (N_7991,N_5185,N_6442);
nor U7992 (N_7992,N_7207,N_6471);
nor U7993 (N_7993,N_5861,N_5841);
nand U7994 (N_7994,N_7337,N_5677);
nand U7995 (N_7995,N_5249,N_5248);
and U7996 (N_7996,N_6987,N_6695);
or U7997 (N_7997,N_6313,N_7012);
nand U7998 (N_7998,N_6864,N_6917);
and U7999 (N_7999,N_6371,N_6523);
nand U8000 (N_8000,N_5874,N_6327);
and U8001 (N_8001,N_6723,N_7349);
and U8002 (N_8002,N_5213,N_6875);
and U8003 (N_8003,N_5270,N_7231);
and U8004 (N_8004,N_6832,N_6913);
and U8005 (N_8005,N_6564,N_7070);
nand U8006 (N_8006,N_6733,N_5256);
nor U8007 (N_8007,N_6997,N_5003);
or U8008 (N_8008,N_6291,N_6526);
and U8009 (N_8009,N_5187,N_7071);
and U8010 (N_8010,N_6210,N_5640);
and U8011 (N_8011,N_7085,N_5399);
and U8012 (N_8012,N_7038,N_5978);
nor U8013 (N_8013,N_6555,N_7031);
or U8014 (N_8014,N_7355,N_5404);
and U8015 (N_8015,N_6805,N_5299);
and U8016 (N_8016,N_6512,N_5056);
and U8017 (N_8017,N_5286,N_6990);
or U8018 (N_8018,N_6489,N_5555);
nor U8019 (N_8019,N_7494,N_7091);
and U8020 (N_8020,N_6783,N_6587);
nor U8021 (N_8021,N_5735,N_5974);
nor U8022 (N_8022,N_5754,N_5591);
and U8023 (N_8023,N_5449,N_7236);
xor U8024 (N_8024,N_5250,N_6081);
nor U8025 (N_8025,N_6474,N_6481);
or U8026 (N_8026,N_6385,N_6324);
nor U8027 (N_8027,N_7395,N_5009);
and U8028 (N_8028,N_6506,N_7241);
nor U8029 (N_8029,N_6869,N_5919);
nand U8030 (N_8030,N_5182,N_5714);
nor U8031 (N_8031,N_7109,N_6368);
or U8032 (N_8032,N_5930,N_6427);
nor U8033 (N_8033,N_5479,N_7451);
nand U8034 (N_8034,N_6075,N_5220);
or U8035 (N_8035,N_6973,N_6933);
and U8036 (N_8036,N_6117,N_6249);
or U8037 (N_8037,N_6798,N_7185);
or U8038 (N_8038,N_6014,N_5347);
and U8039 (N_8039,N_6960,N_5075);
or U8040 (N_8040,N_6857,N_6620);
or U8041 (N_8041,N_5268,N_7266);
and U8042 (N_8042,N_6165,N_7147);
and U8043 (N_8043,N_5658,N_5181);
and U8044 (N_8044,N_5823,N_5156);
or U8045 (N_8045,N_5116,N_5367);
xor U8046 (N_8046,N_5433,N_5696);
and U8047 (N_8047,N_7015,N_7273);
and U8048 (N_8048,N_6343,N_5004);
and U8049 (N_8049,N_6182,N_6437);
nor U8050 (N_8050,N_5158,N_6234);
or U8051 (N_8051,N_5294,N_5276);
and U8052 (N_8052,N_7299,N_5215);
nand U8053 (N_8053,N_5682,N_5794);
and U8054 (N_8054,N_7232,N_5465);
or U8055 (N_8055,N_7079,N_6595);
nor U8056 (N_8056,N_6101,N_6816);
nor U8057 (N_8057,N_5224,N_6219);
nand U8058 (N_8058,N_6518,N_7090);
nand U8059 (N_8059,N_5560,N_5274);
or U8060 (N_8060,N_6074,N_5482);
xor U8061 (N_8061,N_7093,N_5170);
nor U8062 (N_8062,N_5261,N_7422);
nand U8063 (N_8063,N_7170,N_7135);
nor U8064 (N_8064,N_6047,N_6059);
nand U8065 (N_8065,N_6544,N_6528);
nor U8066 (N_8066,N_5496,N_6743);
nor U8067 (N_8067,N_5602,N_6460);
nor U8068 (N_8068,N_5629,N_7208);
nor U8069 (N_8069,N_5173,N_6334);
and U8070 (N_8070,N_5119,N_6188);
and U8071 (N_8071,N_6199,N_5928);
and U8072 (N_8072,N_5500,N_5786);
nand U8073 (N_8073,N_7457,N_5343);
nand U8074 (N_8074,N_5719,N_5577);
and U8075 (N_8075,N_6428,N_5649);
nor U8076 (N_8076,N_5531,N_7447);
nor U8077 (N_8077,N_5684,N_6268);
nand U8078 (N_8078,N_5598,N_5523);
xor U8079 (N_8079,N_7004,N_6842);
or U8080 (N_8080,N_6296,N_7429);
or U8081 (N_8081,N_6836,N_7209);
or U8082 (N_8082,N_5942,N_6009);
or U8083 (N_8083,N_5319,N_5067);
nand U8084 (N_8084,N_5419,N_5631);
or U8085 (N_8085,N_7169,N_6751);
xor U8086 (N_8086,N_5681,N_6085);
or U8087 (N_8087,N_6744,N_7466);
and U8088 (N_8088,N_7161,N_7323);
nand U8089 (N_8089,N_5801,N_7365);
nor U8090 (N_8090,N_5803,N_5468);
nor U8091 (N_8091,N_5848,N_6390);
nand U8092 (N_8092,N_6830,N_5664);
and U8093 (N_8093,N_5507,N_6827);
and U8094 (N_8094,N_5099,N_5589);
or U8095 (N_8095,N_5475,N_6846);
nor U8096 (N_8096,N_5976,N_7353);
and U8097 (N_8097,N_5103,N_7052);
nor U8098 (N_8098,N_5425,N_6068);
nor U8099 (N_8099,N_7325,N_6445);
or U8100 (N_8100,N_7483,N_6650);
or U8101 (N_8101,N_7124,N_6166);
and U8102 (N_8102,N_7285,N_6430);
nor U8103 (N_8103,N_6597,N_5647);
and U8104 (N_8104,N_6238,N_6609);
nand U8105 (N_8105,N_6657,N_6273);
and U8106 (N_8106,N_6237,N_6975);
nor U8107 (N_8107,N_7258,N_6757);
nand U8108 (N_8108,N_6895,N_7405);
and U8109 (N_8109,N_5721,N_7306);
or U8110 (N_8110,N_5994,N_5230);
or U8111 (N_8111,N_6577,N_6340);
or U8112 (N_8112,N_7122,N_5968);
nor U8113 (N_8113,N_5660,N_5613);
or U8114 (N_8114,N_5411,N_5837);
nor U8115 (N_8115,N_6611,N_7210);
nor U8116 (N_8116,N_5850,N_5584);
nor U8117 (N_8117,N_6861,N_6162);
or U8118 (N_8118,N_6728,N_6718);
and U8119 (N_8119,N_6289,N_5305);
or U8120 (N_8120,N_7160,N_5567);
and U8121 (N_8121,N_5222,N_5193);
nand U8122 (N_8122,N_5522,N_6242);
xnor U8123 (N_8123,N_7444,N_5394);
and U8124 (N_8124,N_6750,N_5377);
nand U8125 (N_8125,N_5550,N_6121);
nand U8126 (N_8126,N_6116,N_7056);
or U8127 (N_8127,N_6267,N_5599);
or U8128 (N_8128,N_7385,N_5192);
and U8129 (N_8129,N_6799,N_6590);
nor U8130 (N_8130,N_5307,N_6668);
or U8131 (N_8131,N_5368,N_6099);
and U8132 (N_8132,N_7454,N_6915);
or U8133 (N_8133,N_5564,N_5081);
nand U8134 (N_8134,N_5061,N_5359);
or U8135 (N_8135,N_7192,N_6086);
nand U8136 (N_8136,N_6459,N_5944);
nand U8137 (N_8137,N_5396,N_6844);
or U8138 (N_8138,N_5191,N_5784);
and U8139 (N_8139,N_6985,N_6196);
nand U8140 (N_8140,N_6142,N_5593);
nand U8141 (N_8141,N_6839,N_6963);
and U8142 (N_8142,N_6760,N_6419);
and U8143 (N_8143,N_5429,N_7379);
and U8144 (N_8144,N_7467,N_7408);
and U8145 (N_8145,N_6408,N_5175);
nand U8146 (N_8146,N_5485,N_7075);
nand U8147 (N_8147,N_5575,N_6374);
or U8148 (N_8148,N_5802,N_6477);
nor U8149 (N_8149,N_5057,N_5493);
or U8150 (N_8150,N_6212,N_5339);
nand U8151 (N_8151,N_6944,N_6203);
nor U8152 (N_8152,N_6806,N_6494);
and U8153 (N_8153,N_6883,N_5453);
nand U8154 (N_8154,N_7221,N_6457);
nand U8155 (N_8155,N_6497,N_5713);
nor U8156 (N_8156,N_7442,N_5227);
and U8157 (N_8157,N_5060,N_7154);
and U8158 (N_8158,N_5693,N_6306);
or U8159 (N_8159,N_5321,N_6321);
and U8160 (N_8160,N_6855,N_5750);
nand U8161 (N_8161,N_6163,N_7486);
or U8162 (N_8162,N_7019,N_5132);
and U8163 (N_8163,N_7440,N_7107);
nand U8164 (N_8164,N_5461,N_6062);
and U8165 (N_8165,N_5538,N_5141);
and U8166 (N_8166,N_6809,N_6071);
nand U8167 (N_8167,N_6046,N_5870);
and U8168 (N_8168,N_6767,N_7320);
or U8169 (N_8169,N_6158,N_7261);
nor U8170 (N_8170,N_5534,N_7060);
nand U8171 (N_8171,N_7416,N_5012);
and U8172 (N_8172,N_7409,N_6315);
or U8173 (N_8173,N_6568,N_5160);
nand U8174 (N_8174,N_5793,N_5123);
or U8175 (N_8175,N_5752,N_7072);
and U8176 (N_8176,N_6716,N_6938);
xor U8177 (N_8177,N_6698,N_6475);
nor U8178 (N_8178,N_6769,N_6030);
nor U8179 (N_8179,N_6341,N_5788);
nor U8180 (N_8180,N_5590,N_6778);
and U8181 (N_8181,N_5620,N_6664);
nor U8182 (N_8182,N_6349,N_5318);
nor U8183 (N_8183,N_5078,N_5216);
and U8184 (N_8184,N_6410,N_5035);
or U8185 (N_8185,N_6794,N_7243);
nand U8186 (N_8186,N_5197,N_6707);
and U8187 (N_8187,N_7290,N_5435);
and U8188 (N_8188,N_7493,N_6745);
nor U8189 (N_8189,N_7377,N_5698);
nand U8190 (N_8190,N_6191,N_7347);
nor U8191 (N_8191,N_5627,N_5950);
and U8192 (N_8192,N_5398,N_7102);
nand U8193 (N_8193,N_5670,N_7172);
or U8194 (N_8194,N_7490,N_5606);
and U8195 (N_8195,N_5048,N_6680);
nand U8196 (N_8196,N_6491,N_5559);
nand U8197 (N_8197,N_5570,N_5089);
nand U8198 (N_8198,N_7223,N_6172);
nand U8199 (N_8199,N_6413,N_5659);
nor U8200 (N_8200,N_7180,N_6164);
and U8201 (N_8201,N_5715,N_5292);
or U8202 (N_8202,N_5849,N_6435);
nor U8203 (N_8203,N_6125,N_5120);
or U8204 (N_8204,N_5618,N_5040);
nand U8205 (N_8205,N_6509,N_6715);
nor U8206 (N_8206,N_5391,N_6434);
and U8207 (N_8207,N_6124,N_5298);
xor U8208 (N_8208,N_6904,N_6882);
or U8209 (N_8209,N_6569,N_5853);
nor U8210 (N_8210,N_5960,N_6986);
nor U8211 (N_8211,N_5562,N_5107);
or U8212 (N_8212,N_5317,N_7101);
nor U8213 (N_8213,N_5467,N_6683);
nand U8214 (N_8214,N_5554,N_6897);
nand U8215 (N_8215,N_7086,N_7136);
or U8216 (N_8216,N_6100,N_6932);
nor U8217 (N_8217,N_5755,N_5778);
nor U8218 (N_8218,N_5316,N_6010);
or U8219 (N_8219,N_6945,N_7248);
nor U8220 (N_8220,N_6800,N_6139);
and U8221 (N_8221,N_6817,N_7174);
nand U8222 (N_8222,N_5205,N_6473);
or U8223 (N_8223,N_5395,N_6345);
and U8224 (N_8224,N_5083,N_6824);
xor U8225 (N_8225,N_6254,N_6747);
nand U8226 (N_8226,N_7097,N_6859);
nor U8227 (N_8227,N_7495,N_6275);
nand U8228 (N_8228,N_7421,N_6131);
nand U8229 (N_8229,N_7361,N_7438);
nand U8230 (N_8230,N_7398,N_5553);
nor U8231 (N_8231,N_6837,N_5145);
nor U8232 (N_8232,N_7218,N_5694);
or U8233 (N_8233,N_6645,N_5579);
nand U8234 (N_8234,N_5110,N_6606);
nand U8235 (N_8235,N_7307,N_5032);
nand U8236 (N_8236,N_5415,N_6734);
nand U8237 (N_8237,N_6266,N_7039);
nand U8238 (N_8238,N_6329,N_6572);
or U8239 (N_8239,N_5931,N_5082);
nor U8240 (N_8240,N_6533,N_6999);
nand U8241 (N_8241,N_7461,N_6872);
or U8242 (N_8242,N_7141,N_5337);
and U8243 (N_8243,N_5632,N_5370);
nand U8244 (N_8244,N_7328,N_6493);
nor U8245 (N_8245,N_5655,N_7350);
and U8246 (N_8246,N_5674,N_7463);
nor U8247 (N_8247,N_7313,N_5663);
nand U8248 (N_8248,N_7312,N_5726);
nor U8249 (N_8249,N_5016,N_5635);
or U8250 (N_8250,N_7406,N_6202);
nor U8251 (N_8251,N_6787,N_5109);
nand U8252 (N_8252,N_7025,N_6145);
nor U8253 (N_8253,N_7011,N_6338);
and U8254 (N_8254,N_5532,N_6885);
or U8255 (N_8255,N_6622,N_5813);
and U8256 (N_8256,N_5114,N_5623);
nand U8257 (N_8257,N_6686,N_5137);
nor U8258 (N_8258,N_7078,N_6776);
or U8259 (N_8259,N_5308,N_5764);
xnor U8260 (N_8260,N_7445,N_6373);
and U8261 (N_8261,N_5497,N_6730);
nor U8262 (N_8262,N_5478,N_7368);
nand U8263 (N_8263,N_6845,N_6429);
nor U8264 (N_8264,N_5097,N_6008);
or U8265 (N_8265,N_5161,N_5700);
or U8266 (N_8266,N_6870,N_7212);
xor U8267 (N_8267,N_5265,N_7253);
or U8268 (N_8268,N_5633,N_7254);
or U8269 (N_8269,N_5277,N_5186);
or U8270 (N_8270,N_7242,N_5000);
or U8271 (N_8271,N_5402,N_5923);
nand U8272 (N_8272,N_7472,N_5777);
nor U8273 (N_8273,N_5129,N_6194);
nor U8274 (N_8274,N_5669,N_6420);
nor U8275 (N_8275,N_5422,N_6277);
and U8276 (N_8276,N_6588,N_5226);
nor U8277 (N_8277,N_7287,N_6621);
or U8278 (N_8278,N_7145,N_5955);
nor U8279 (N_8279,N_7372,N_5675);
and U8280 (N_8280,N_6994,N_5662);
nor U8281 (N_8281,N_5628,N_6400);
nand U8282 (N_8282,N_5080,N_5600);
nor U8283 (N_8283,N_7443,N_6535);
nor U8284 (N_8284,N_5058,N_5569);
or U8285 (N_8285,N_5883,N_5164);
and U8286 (N_8286,N_6041,N_6381);
nor U8287 (N_8287,N_5296,N_6722);
or U8288 (N_8288,N_7375,N_5983);
nand U8289 (N_8289,N_7106,N_6209);
xor U8290 (N_8290,N_6853,N_6926);
nor U8291 (N_8291,N_5386,N_6541);
nand U8292 (N_8292,N_6964,N_6411);
nor U8293 (N_8293,N_7076,N_6576);
or U8294 (N_8294,N_5878,N_5864);
nand U8295 (N_8295,N_6090,N_5238);
or U8296 (N_8296,N_6731,N_7007);
or U8297 (N_8297,N_6598,N_5438);
and U8298 (N_8298,N_6962,N_6484);
and U8299 (N_8299,N_5953,N_6173);
nand U8300 (N_8300,N_6814,N_6952);
xor U8301 (N_8301,N_6360,N_6676);
nor U8302 (N_8302,N_5594,N_6292);
nor U8303 (N_8303,N_6812,N_7276);
nand U8304 (N_8304,N_5344,N_7418);
and U8305 (N_8305,N_5459,N_7130);
or U8306 (N_8306,N_5733,N_6919);
nand U8307 (N_8307,N_5005,N_7314);
and U8308 (N_8308,N_5958,N_5763);
xor U8309 (N_8309,N_6524,N_6531);
or U8310 (N_8310,N_6971,N_5608);
or U8311 (N_8311,N_5679,N_5966);
nor U8312 (N_8312,N_5661,N_6996);
nand U8313 (N_8313,N_6387,N_6935);
or U8314 (N_8314,N_6679,N_5349);
xnor U8315 (N_8315,N_5737,N_6129);
and U8316 (N_8316,N_5053,N_5580);
and U8317 (N_8317,N_5731,N_6922);
or U8318 (N_8318,N_5708,N_6803);
or U8319 (N_8319,N_6804,N_6781);
nor U8320 (N_8320,N_7384,N_7156);
nor U8321 (N_8321,N_5610,N_5376);
or U8322 (N_8322,N_7465,N_7132);
and U8323 (N_8323,N_5676,N_6443);
and U8324 (N_8324,N_7381,N_6724);
nand U8325 (N_8325,N_5524,N_7364);
nand U8326 (N_8326,N_6881,N_5071);
nand U8327 (N_8327,N_6729,N_5657);
nand U8328 (N_8328,N_7112,N_5831);
and U8329 (N_8329,N_6583,N_5452);
nand U8330 (N_8330,N_6318,N_6346);
and U8331 (N_8331,N_5511,N_5852);
nand U8332 (N_8332,N_7282,N_5614);
or U8333 (N_8333,N_5774,N_5541);
nand U8334 (N_8334,N_6323,N_5302);
nor U8335 (N_8335,N_6582,N_7084);
or U8336 (N_8336,N_5454,N_5122);
or U8337 (N_8337,N_5416,N_7420);
nand U8338 (N_8338,N_6200,N_6848);
nor U8339 (N_8339,N_6151,N_6094);
nand U8340 (N_8340,N_6525,N_6955);
nand U8341 (N_8341,N_5424,N_5210);
nor U8342 (N_8342,N_7074,N_7100);
or U8343 (N_8343,N_6003,N_5196);
and U8344 (N_8344,N_5272,N_5117);
nand U8345 (N_8345,N_7304,N_7400);
and U8346 (N_8346,N_6472,N_6153);
and U8347 (N_8347,N_7346,N_5641);
nand U8348 (N_8348,N_5797,N_7288);
nor U8349 (N_8349,N_5121,N_6032);
nor U8350 (N_8350,N_5231,N_6004);
nand U8351 (N_8351,N_5734,N_7225);
nand U8352 (N_8352,N_6136,N_5621);
or U8353 (N_8353,N_7294,N_6702);
nand U8354 (N_8354,N_6253,N_6190);
nor U8355 (N_8355,N_5464,N_5168);
or U8356 (N_8356,N_5796,N_7471);
and U8357 (N_8357,N_6849,N_7092);
and U8358 (N_8358,N_6011,N_7404);
nor U8359 (N_8359,N_7016,N_5758);
and U8360 (N_8360,N_6490,N_6144);
nor U8361 (N_8361,N_7497,N_6874);
or U8362 (N_8362,N_5417,N_5816);
or U8363 (N_8363,N_7043,N_5785);
or U8364 (N_8364,N_5986,N_5011);
and U8365 (N_8365,N_6639,N_6031);
nand U8366 (N_8366,N_6178,N_5407);
and U8367 (N_8367,N_6785,N_6309);
nor U8368 (N_8368,N_6520,N_6727);
and U8369 (N_8369,N_7318,N_5728);
or U8370 (N_8370,N_6115,N_6930);
nor U8371 (N_8371,N_6407,N_6835);
nand U8372 (N_8372,N_6507,N_6565);
nand U8373 (N_8373,N_7183,N_7262);
and U8374 (N_8374,N_7193,N_6626);
or U8375 (N_8375,N_6560,N_5526);
nor U8376 (N_8376,N_6681,N_6187);
nand U8377 (N_8377,N_5730,N_7339);
and U8378 (N_8378,N_6019,N_5665);
nand U8379 (N_8379,N_6711,N_6456);
nor U8380 (N_8380,N_5956,N_7045);
and U8381 (N_8381,N_6505,N_6951);
nor U8382 (N_8382,N_6114,N_6092);
and U8383 (N_8383,N_5687,N_6206);
and U8384 (N_8384,N_5927,N_5574);
nor U8385 (N_8385,N_5171,N_5643);
or U8386 (N_8386,N_7396,N_5767);
nor U8387 (N_8387,N_6980,N_5146);
nand U8388 (N_8388,N_5805,N_7469);
and U8389 (N_8389,N_7049,N_7449);
nor U8390 (N_8390,N_7419,N_7425);
or U8391 (N_8391,N_6549,N_6791);
nand U8392 (N_8392,N_5882,N_6705);
nor U8393 (N_8393,N_5375,N_5565);
or U8394 (N_8394,N_6426,N_5477);
nor U8395 (N_8395,N_6615,N_5490);
xor U8396 (N_8396,N_7129,N_6907);
and U8397 (N_8397,N_7197,N_5135);
or U8398 (N_8398,N_5982,N_6152);
or U8399 (N_8399,N_5790,N_5780);
nor U8400 (N_8400,N_6073,N_5938);
and U8401 (N_8401,N_6682,N_5090);
nand U8402 (N_8402,N_7388,N_6159);
nor U8403 (N_8403,N_5825,N_5084);
nor U8404 (N_8404,N_6256,N_5607);
or U8405 (N_8405,N_7414,N_6208);
or U8406 (N_8406,N_5977,N_5489);
or U8407 (N_8407,N_6018,N_7133);
or U8408 (N_8408,N_6098,N_5648);
nand U8409 (N_8409,N_5357,N_5070);
or U8410 (N_8410,N_7256,N_6655);
or U8411 (N_8411,N_7478,N_6792);
or U8412 (N_8412,N_6077,N_6916);
nand U8413 (N_8413,N_6417,N_6350);
and U8414 (N_8414,N_7335,N_6850);
nor U8415 (N_8415,N_5282,N_6793);
nand U8416 (N_8416,N_7267,N_5940);
nor U8417 (N_8417,N_6216,N_5288);
or U8418 (N_8418,N_6545,N_5015);
and U8419 (N_8419,N_5374,N_7029);
or U8420 (N_8420,N_6412,N_5959);
or U8421 (N_8421,N_5163,N_5051);
xor U8422 (N_8422,N_5815,N_5766);
nor U8423 (N_8423,N_7035,N_6284);
and U8424 (N_8424,N_7498,N_6076);
or U8425 (N_8425,N_5578,N_6772);
nand U8426 (N_8426,N_7125,N_5301);
nor U8427 (N_8427,N_6978,N_6486);
nand U8428 (N_8428,N_5028,N_7114);
nor U8429 (N_8429,N_6169,N_6775);
nand U8430 (N_8430,N_6251,N_6969);
and U8431 (N_8431,N_6137,N_5808);
nor U8432 (N_8432,N_6929,N_5995);
nor U8433 (N_8433,N_5710,N_5561);
nor U8434 (N_8434,N_6866,N_7296);
and U8435 (N_8435,N_6028,N_6537);
nor U8436 (N_8436,N_5441,N_5100);
or U8437 (N_8437,N_6415,N_5688);
or U8438 (N_8438,N_6532,N_7448);
nor U8439 (N_8439,N_6367,N_6738);
and U8440 (N_8440,N_5626,N_5178);
or U8441 (N_8441,N_5656,N_6441);
and U8442 (N_8442,N_6580,N_5266);
nand U8443 (N_8443,N_6025,N_7297);
nand U8444 (N_8444,N_7324,N_5073);
and U8445 (N_8445,N_6633,N_5306);
nor U8446 (N_8446,N_5342,N_6414);
xnor U8447 (N_8447,N_5102,N_6097);
nand U8448 (N_8448,N_6712,N_5701);
nand U8449 (N_8449,N_5338,N_7453);
or U8450 (N_8450,N_6911,N_5756);
nor U8451 (N_8451,N_5634,N_5334);
nand U8452 (N_8452,N_7286,N_6463);
and U8453 (N_8453,N_5013,N_7348);
nor U8454 (N_8454,N_5329,N_5746);
nor U8455 (N_8455,N_6213,N_5991);
nand U8456 (N_8456,N_5536,N_6252);
and U8457 (N_8457,N_6503,N_5678);
and U8458 (N_8458,N_7159,N_7402);
nor U8459 (N_8459,N_6910,N_5085);
or U8460 (N_8460,N_6379,N_6055);
xnor U8461 (N_8461,N_5957,N_6084);
or U8462 (N_8462,N_5234,N_7149);
nand U8463 (N_8463,N_7187,N_6953);
nor U8464 (N_8464,N_7148,N_7188);
nor U8465 (N_8465,N_5689,N_6516);
and U8466 (N_8466,N_5401,N_6991);
nand U8467 (N_8467,N_6833,N_5236);
nand U8468 (N_8468,N_5118,N_5052);
and U8469 (N_8469,N_6038,N_7436);
or U8470 (N_8470,N_6498,N_7002);
nand U8471 (N_8471,N_6436,N_6768);
and U8472 (N_8472,N_7315,N_5284);
or U8473 (N_8473,N_5819,N_6272);
nand U8474 (N_8474,N_7397,N_5806);
nand U8475 (N_8475,N_5390,N_6048);
or U8476 (N_8476,N_5543,N_7240);
or U8477 (N_8477,N_5492,N_6054);
nand U8478 (N_8478,N_6784,N_5772);
and U8479 (N_8479,N_5970,N_5948);
xor U8480 (N_8480,N_6725,N_6322);
nor U8481 (N_8481,N_6697,N_7317);
and U8482 (N_8482,N_6547,N_5542);
nand U8483 (N_8483,N_6585,N_6905);
or U8484 (N_8484,N_6394,N_6235);
or U8485 (N_8485,N_5695,N_6197);
nor U8486 (N_8486,N_6293,N_5544);
nand U8487 (N_8487,N_7176,N_7473);
or U8488 (N_8488,N_6708,N_6370);
nand U8489 (N_8489,N_6223,N_7280);
and U8490 (N_8490,N_5202,N_5711);
nand U8491 (N_8491,N_5932,N_7059);
and U8492 (N_8492,N_6589,N_7356);
nor U8493 (N_8493,N_6110,N_5653);
or U8494 (N_8494,N_6713,N_5183);
or U8495 (N_8495,N_5901,N_6988);
or U8496 (N_8496,N_6450,N_7194);
or U8497 (N_8497,N_6903,N_5826);
nand U8498 (N_8498,N_6802,N_5363);
xor U8499 (N_8499,N_6401,N_7143);
nor U8500 (N_8500,N_5924,N_5937);
and U8501 (N_8501,N_6096,N_7450);
nand U8502 (N_8502,N_5654,N_6717);
nand U8503 (N_8503,N_6992,N_6689);
or U8504 (N_8504,N_5887,N_7371);
and U8505 (N_8505,N_7366,N_6286);
nor U8506 (N_8506,N_7432,N_6647);
nor U8507 (N_8507,N_6146,N_6732);
nor U8508 (N_8508,N_7259,N_5833);
nand U8509 (N_8509,N_5673,N_6424);
nor U8510 (N_8510,N_6027,N_7044);
nor U8511 (N_8511,N_6755,N_6214);
nand U8512 (N_8512,N_5949,N_7219);
nor U8513 (N_8513,N_5400,N_5446);
nor U8514 (N_8514,N_6333,N_6347);
and U8515 (N_8515,N_5095,N_7104);
nand U8516 (N_8516,N_6770,N_6211);
xor U8517 (N_8517,N_6873,N_5014);
or U8518 (N_8518,N_5408,N_5046);
or U8519 (N_8519,N_6899,N_5074);
and U8520 (N_8520,N_5208,N_5838);
nand U8521 (N_8521,N_6900,N_5314);
or U8522 (N_8522,N_6934,N_6246);
and U8523 (N_8523,N_5412,N_6000);
or U8524 (N_8524,N_5747,N_5830);
nor U8525 (N_8525,N_6181,N_5642);
nor U8526 (N_8526,N_6826,N_6294);
or U8527 (N_8527,N_6024,N_5125);
nand U8528 (N_8528,N_7054,N_5904);
and U8529 (N_8529,N_5723,N_5209);
nor U8530 (N_8530,N_5194,N_6375);
or U8531 (N_8531,N_7203,N_5683);
and U8532 (N_8532,N_5722,N_6893);
or U8533 (N_8533,N_7439,N_6807);
or U8534 (N_8534,N_6107,N_5462);
xnor U8535 (N_8535,N_7235,N_6362);
or U8536 (N_8536,N_7173,N_6959);
nor U8537 (N_8537,N_6663,N_5990);
or U8538 (N_8538,N_7040,N_6656);
nor U8539 (N_8539,N_5124,N_6281);
nor U8540 (N_8540,N_7064,N_7351);
or U8541 (N_8541,N_5225,N_5113);
nor U8542 (N_8542,N_5041,N_6279);
and U8543 (N_8543,N_5512,N_6594);
nand U8544 (N_8544,N_6250,N_6167);
nor U8545 (N_8545,N_7330,N_6123);
nand U8546 (N_8546,N_6613,N_6044);
and U8547 (N_8547,N_7264,N_5448);
and U8548 (N_8548,N_6488,N_5981);
nand U8549 (N_8549,N_5443,N_5346);
and U8550 (N_8550,N_6227,N_7265);
nor U8551 (N_8551,N_6758,N_5018);
nand U8552 (N_8552,N_5789,N_5331);
nor U8553 (N_8553,N_6177,N_5087);
nand U8554 (N_8554,N_5576,N_5188);
nand U8555 (N_8555,N_5010,N_7357);
nand U8556 (N_8556,N_6336,N_6119);
nor U8557 (N_8557,N_6184,N_6543);
nor U8558 (N_8558,N_6542,N_7310);
or U8559 (N_8559,N_6189,N_6752);
nand U8560 (N_8560,N_6192,N_5820);
nand U8561 (N_8561,N_5551,N_5954);
nand U8562 (N_8562,N_6255,N_5773);
nor U8563 (N_8563,N_7048,N_7342);
nor U8564 (N_8564,N_6970,N_5846);
and U8565 (N_8565,N_5431,N_6607);
nand U8566 (N_8566,N_6245,N_6483);
nand U8567 (N_8567,N_5539,N_6671);
and U8568 (N_8568,N_7220,N_6359);
nand U8569 (N_8569,N_6762,N_7292);
or U8570 (N_8570,N_5491,N_6421);
and U8571 (N_8571,N_6217,N_6228);
or U8572 (N_8572,N_7204,N_5799);
nand U8573 (N_8573,N_5895,N_7001);
or U8574 (N_8574,N_6629,N_5509);
nand U8575 (N_8575,N_6220,N_6231);
nand U8576 (N_8576,N_5963,N_5603);
nand U8577 (N_8577,N_5972,N_6183);
nor U8578 (N_8578,N_6454,N_5505);
nor U8579 (N_8579,N_6740,N_5341);
nor U8580 (N_8580,N_5702,N_5699);
nand U8581 (N_8581,N_5373,N_5951);
or U8582 (N_8582,N_6918,N_7083);
and U8583 (N_8583,N_5054,N_7036);
or U8584 (N_8584,N_7399,N_7289);
nor U8585 (N_8585,N_6673,N_5712);
nor U8586 (N_8586,N_5943,N_5519);
nand U8587 (N_8587,N_7184,N_6822);
or U8588 (N_8588,N_5430,N_7279);
and U8589 (N_8589,N_6160,N_5903);
and U8590 (N_8590,N_6703,N_6909);
nor U8591 (N_8591,N_6088,N_7000);
and U8592 (N_8592,N_7499,N_5021);
nand U8593 (N_8593,N_5426,N_7182);
and U8594 (N_8594,N_7446,N_6485);
nor U8595 (N_8595,N_5961,N_6813);
nand U8596 (N_8596,N_5717,N_7278);
or U8597 (N_8597,N_5138,N_7108);
nand U8598 (N_8598,N_5333,N_5718);
nor U8599 (N_8599,N_6462,N_5330);
nand U8600 (N_8600,N_5195,N_5547);
nor U8601 (N_8601,N_5909,N_5434);
nand U8602 (N_8602,N_6023,N_6311);
and U8603 (N_8603,N_6314,N_6644);
and U8604 (N_8604,N_6694,N_7230);
or U8605 (N_8605,N_5350,N_5886);
nor U8606 (N_8606,N_5130,N_6364);
nor U8607 (N_8607,N_5381,N_6171);
nand U8608 (N_8608,N_5289,N_5281);
nor U8609 (N_8609,N_5740,N_5380);
nand U8610 (N_8610,N_7186,N_5036);
nand U8611 (N_8611,N_6002,N_6265);
or U8612 (N_8612,N_6658,N_6610);
or U8613 (N_8613,N_5588,N_6317);
and U8614 (N_8614,N_7488,N_7105);
nor U8615 (N_8615,N_7428,N_6634);
nor U8616 (N_8616,N_6624,N_6095);
nor U8617 (N_8617,N_5311,N_6466);
or U8618 (N_8618,N_7326,N_5568);
and U8619 (N_8619,N_5859,N_7476);
or U8620 (N_8620,N_7470,N_5201);
and U8621 (N_8621,N_7164,N_6300);
and U8622 (N_8622,N_6502,N_5382);
nand U8623 (N_8623,N_6406,N_5980);
and U8624 (N_8624,N_6204,N_5571);
nor U8625 (N_8625,N_7475,N_6067);
and U8626 (N_8626,N_6389,N_5811);
or U8627 (N_8627,N_6600,N_5456);
nand U8628 (N_8628,N_7087,N_6756);
nor U8629 (N_8629,N_6482,N_7431);
or U8630 (N_8630,N_5059,N_5668);
or U8631 (N_8631,N_5921,N_6229);
nor U8632 (N_8632,N_6109,N_5807);
nand U8633 (N_8633,N_5622,N_5867);
nand U8634 (N_8634,N_7126,N_7459);
and U8635 (N_8635,N_5260,N_5527);
nor U8636 (N_8636,N_5325,N_7047);
and U8637 (N_8637,N_5228,N_5890);
nand U8638 (N_8638,N_6348,N_5275);
and U8639 (N_8639,N_6818,N_6304);
nand U8640 (N_8640,N_5229,N_5055);
or U8641 (N_8641,N_5625,N_5466);
or U8642 (N_8642,N_6989,N_5427);
nand U8643 (N_8643,N_5829,N_7053);
and U8644 (N_8644,N_5362,N_6257);
nor U8645 (N_8645,N_5862,N_5155);
nor U8646 (N_8646,N_5779,N_5768);
and U8647 (N_8647,N_5962,N_5414);
nor U8648 (N_8648,N_5365,N_5470);
and U8649 (N_8649,N_6040,N_6455);
nand U8650 (N_8650,N_6248,N_6815);
and U8651 (N_8651,N_6584,N_7303);
and U8652 (N_8652,N_7137,N_6330);
or U8653 (N_8653,N_5952,N_6335);
or U8654 (N_8654,N_6130,N_6754);
nor U8655 (N_8655,N_6093,N_7140);
nand U8656 (N_8656,N_6377,N_6574);
and U8657 (N_8657,N_7117,N_6319);
or U8658 (N_8658,N_6316,N_5190);
nand U8659 (N_8659,N_6931,N_6380);
nor U8660 (N_8660,N_5595,N_5592);
and U8661 (N_8661,N_5450,N_6399);
nor U8662 (N_8662,N_5050,N_6879);
xnor U8663 (N_8663,N_6764,N_5384);
and U8664 (N_8664,N_6015,N_6949);
or U8665 (N_8665,N_5783,N_6578);
or U8666 (N_8666,N_5487,N_5646);
and U8667 (N_8667,N_5340,N_5609);
or U8668 (N_8668,N_5835,N_6890);
and U8669 (N_8669,N_5351,N_6706);
and U8670 (N_8670,N_6651,N_7344);
nor U8671 (N_8671,N_5997,N_6630);
nand U8672 (N_8672,N_6439,N_5586);
nor U8673 (N_8673,N_7331,N_7200);
or U8674 (N_8674,N_5881,N_7181);
nand U8675 (N_8675,N_5832,N_6825);
and U8676 (N_8676,N_7089,N_5031);
or U8677 (N_8677,N_6950,N_5352);
and U8678 (N_8678,N_6841,N_5474);
nand U8679 (N_8679,N_5218,N_5254);
and U8680 (N_8680,N_7131,N_6546);
nor U8681 (N_8681,N_6138,N_5716);
nand U8682 (N_8682,N_5445,N_7227);
nor U8683 (N_8683,N_5066,N_6326);
and U8684 (N_8684,N_6894,N_5421);
or U8685 (N_8685,N_5563,N_5840);
or U8686 (N_8686,N_6388,N_6060);
nor U8687 (N_8687,N_5749,N_5898);
and U8688 (N_8688,N_5345,N_7062);
and U8689 (N_8689,N_5985,N_6670);
nor U8690 (N_8690,N_5518,N_7153);
nand U8691 (N_8691,N_7329,N_5552);
or U8692 (N_8692,N_7233,N_5243);
nand U8693 (N_8693,N_5157,N_6372);
or U8694 (N_8694,N_7057,N_5242);
or U8695 (N_8695,N_6961,N_7030);
nand U8696 (N_8696,N_6499,N_6661);
nand U8697 (N_8697,N_7378,N_6127);
nor U8698 (N_8698,N_6720,N_6468);
nor U8699 (N_8699,N_6906,N_6012);
or U8700 (N_8700,N_7116,N_6342);
xnor U8701 (N_8701,N_5572,N_5906);
nand U8702 (N_8702,N_6604,N_6355);
nor U8703 (N_8703,N_6840,N_5727);
xnor U8704 (N_8704,N_6887,N_7464);
or U8705 (N_8705,N_5893,N_5765);
and U8706 (N_8706,N_5257,N_5585);
or U8707 (N_8707,N_6789,N_6596);
or U8708 (N_8708,N_6627,N_6017);
nor U8709 (N_8709,N_6649,N_5444);
nor U8710 (N_8710,N_5908,N_7032);
nand U8711 (N_8711,N_5604,N_7352);
and U8712 (N_8712,N_5214,N_6232);
and U8713 (N_8713,N_5854,N_6984);
nand U8714 (N_8714,N_7460,N_5451);
and U8715 (N_8715,N_6045,N_6120);
nor U8716 (N_8716,N_6396,N_6514);
nand U8717 (N_8717,N_5900,N_7217);
nor U8718 (N_8718,N_7311,N_6972);
nand U8719 (N_8719,N_5707,N_6271);
nand U8720 (N_8720,N_5455,N_5147);
nand U8721 (N_8721,N_7376,N_6458);
and U8722 (N_8722,N_5769,N_6586);
and U8723 (N_8723,N_6021,N_5030);
and U8724 (N_8724,N_5315,N_7006);
or U8725 (N_8725,N_6186,N_5112);
and U8726 (N_8726,N_5863,N_5258);
or U8727 (N_8727,N_5104,N_6042);
nand U8728 (N_8728,N_5326,N_7017);
nand U8729 (N_8729,N_5101,N_5510);
and U8730 (N_8730,N_7263,N_6635);
nand U8731 (N_8731,N_6233,N_6140);
nor U8732 (N_8732,N_5998,N_7392);
and U8733 (N_8733,N_6141,N_7382);
or U8734 (N_8734,N_5917,N_5795);
nor U8735 (N_8735,N_6982,N_5792);
nor U8736 (N_8736,N_5871,N_6957);
xnor U8737 (N_8737,N_6921,N_6923);
nand U8738 (N_8738,N_5638,N_5463);
nand U8739 (N_8739,N_6667,N_6287);
and U8740 (N_8740,N_6571,N_5457);
and U8741 (N_8741,N_7110,N_7214);
nand U8742 (N_8742,N_5671,N_7474);
nand U8743 (N_8743,N_7119,N_7150);
and U8744 (N_8744,N_6831,N_7456);
or U8745 (N_8745,N_5327,N_7492);
and U8746 (N_8746,N_5705,N_7321);
and U8747 (N_8747,N_5911,N_6363);
nor U8748 (N_8748,N_5356,N_5291);
nor U8749 (N_8749,N_5495,N_5271);
nand U8750 (N_8750,N_5922,N_5068);
nand U8751 (N_8751,N_6844,N_6865);
nand U8752 (N_8752,N_5412,N_6107);
or U8753 (N_8753,N_5248,N_7485);
nand U8754 (N_8754,N_5192,N_6295);
and U8755 (N_8755,N_7296,N_7009);
and U8756 (N_8756,N_5368,N_5485);
or U8757 (N_8757,N_6891,N_5098);
nand U8758 (N_8758,N_5107,N_6667);
nor U8759 (N_8759,N_5843,N_6990);
or U8760 (N_8760,N_5075,N_5433);
nand U8761 (N_8761,N_5671,N_6947);
and U8762 (N_8762,N_5791,N_5913);
and U8763 (N_8763,N_6460,N_6750);
and U8764 (N_8764,N_6574,N_6515);
nor U8765 (N_8765,N_6587,N_7460);
and U8766 (N_8766,N_7035,N_5841);
nor U8767 (N_8767,N_5227,N_5250);
nand U8768 (N_8768,N_7278,N_5109);
nand U8769 (N_8769,N_5156,N_5149);
nand U8770 (N_8770,N_5000,N_7140);
xnor U8771 (N_8771,N_6126,N_6157);
or U8772 (N_8772,N_5034,N_6974);
nand U8773 (N_8773,N_7236,N_6614);
or U8774 (N_8774,N_6594,N_6679);
xnor U8775 (N_8775,N_6707,N_5876);
or U8776 (N_8776,N_6359,N_5267);
or U8777 (N_8777,N_6274,N_5294);
or U8778 (N_8778,N_6482,N_6338);
or U8779 (N_8779,N_6445,N_6815);
or U8780 (N_8780,N_5771,N_6822);
and U8781 (N_8781,N_5708,N_6216);
or U8782 (N_8782,N_6263,N_5207);
or U8783 (N_8783,N_6061,N_6641);
nor U8784 (N_8784,N_7033,N_5098);
nor U8785 (N_8785,N_6814,N_7351);
and U8786 (N_8786,N_6187,N_7314);
nor U8787 (N_8787,N_7376,N_7310);
or U8788 (N_8788,N_5479,N_7092);
nand U8789 (N_8789,N_6706,N_7205);
or U8790 (N_8790,N_6941,N_6712);
and U8791 (N_8791,N_5214,N_7396);
and U8792 (N_8792,N_5155,N_5331);
nor U8793 (N_8793,N_7433,N_6623);
nor U8794 (N_8794,N_6903,N_6009);
and U8795 (N_8795,N_5570,N_5872);
and U8796 (N_8796,N_6178,N_7249);
nand U8797 (N_8797,N_6778,N_6790);
nand U8798 (N_8798,N_5563,N_7044);
nor U8799 (N_8799,N_5480,N_5463);
nor U8800 (N_8800,N_6613,N_6222);
nor U8801 (N_8801,N_7470,N_5645);
nand U8802 (N_8802,N_5078,N_5943);
xor U8803 (N_8803,N_5697,N_5737);
or U8804 (N_8804,N_5623,N_6783);
nor U8805 (N_8805,N_6514,N_5116);
or U8806 (N_8806,N_5379,N_7229);
xor U8807 (N_8807,N_5598,N_6902);
or U8808 (N_8808,N_5895,N_5107);
and U8809 (N_8809,N_7177,N_7023);
and U8810 (N_8810,N_7278,N_7173);
and U8811 (N_8811,N_7370,N_6197);
nor U8812 (N_8812,N_7248,N_7148);
and U8813 (N_8813,N_6841,N_5480);
or U8814 (N_8814,N_6100,N_5205);
nor U8815 (N_8815,N_5470,N_5265);
or U8816 (N_8816,N_7131,N_7287);
xnor U8817 (N_8817,N_5118,N_5255);
nand U8818 (N_8818,N_7134,N_5561);
and U8819 (N_8819,N_5918,N_6159);
nand U8820 (N_8820,N_6824,N_6849);
or U8821 (N_8821,N_6216,N_6921);
nand U8822 (N_8822,N_6010,N_7473);
nand U8823 (N_8823,N_5048,N_6475);
nor U8824 (N_8824,N_6931,N_7121);
or U8825 (N_8825,N_5697,N_6891);
and U8826 (N_8826,N_6861,N_7254);
nand U8827 (N_8827,N_7033,N_6368);
or U8828 (N_8828,N_6445,N_6400);
nor U8829 (N_8829,N_7237,N_6815);
xnor U8830 (N_8830,N_6669,N_5871);
nand U8831 (N_8831,N_5760,N_6618);
nand U8832 (N_8832,N_6947,N_5060);
or U8833 (N_8833,N_6483,N_6509);
and U8834 (N_8834,N_5973,N_7108);
nand U8835 (N_8835,N_5927,N_5023);
nor U8836 (N_8836,N_5906,N_7335);
and U8837 (N_8837,N_5666,N_7140);
and U8838 (N_8838,N_6006,N_7256);
or U8839 (N_8839,N_6636,N_5664);
and U8840 (N_8840,N_7123,N_6274);
or U8841 (N_8841,N_6875,N_6173);
and U8842 (N_8842,N_7071,N_6584);
and U8843 (N_8843,N_6342,N_5620);
xor U8844 (N_8844,N_6202,N_6033);
or U8845 (N_8845,N_5776,N_5225);
nand U8846 (N_8846,N_7024,N_6522);
or U8847 (N_8847,N_5431,N_6844);
nor U8848 (N_8848,N_7049,N_6575);
nor U8849 (N_8849,N_6198,N_6239);
nor U8850 (N_8850,N_5040,N_7315);
nand U8851 (N_8851,N_7468,N_5381);
nand U8852 (N_8852,N_6396,N_5452);
and U8853 (N_8853,N_7243,N_5433);
or U8854 (N_8854,N_6209,N_5025);
or U8855 (N_8855,N_6392,N_6988);
xor U8856 (N_8856,N_5121,N_5079);
nor U8857 (N_8857,N_6495,N_6947);
or U8858 (N_8858,N_6822,N_6625);
and U8859 (N_8859,N_5194,N_5004);
and U8860 (N_8860,N_6260,N_7427);
nand U8861 (N_8861,N_5297,N_5265);
or U8862 (N_8862,N_6632,N_7133);
and U8863 (N_8863,N_7206,N_7435);
nor U8864 (N_8864,N_5494,N_5375);
or U8865 (N_8865,N_6405,N_7097);
nor U8866 (N_8866,N_5650,N_7304);
or U8867 (N_8867,N_6728,N_5196);
nor U8868 (N_8868,N_5583,N_5201);
or U8869 (N_8869,N_6693,N_5624);
nor U8870 (N_8870,N_5048,N_6221);
nand U8871 (N_8871,N_5932,N_5780);
or U8872 (N_8872,N_5422,N_5219);
nor U8873 (N_8873,N_5414,N_5161);
and U8874 (N_8874,N_6279,N_5879);
nor U8875 (N_8875,N_6606,N_6069);
or U8876 (N_8876,N_5065,N_6456);
and U8877 (N_8877,N_5423,N_6668);
nand U8878 (N_8878,N_6297,N_6292);
xnor U8879 (N_8879,N_5778,N_5455);
and U8880 (N_8880,N_6967,N_6378);
or U8881 (N_8881,N_5903,N_5523);
or U8882 (N_8882,N_5217,N_7112);
xnor U8883 (N_8883,N_7284,N_5663);
and U8884 (N_8884,N_5989,N_5482);
and U8885 (N_8885,N_7082,N_5423);
nand U8886 (N_8886,N_6855,N_5440);
nand U8887 (N_8887,N_5351,N_6059);
or U8888 (N_8888,N_6853,N_7200);
nor U8889 (N_8889,N_6742,N_6171);
and U8890 (N_8890,N_5984,N_7080);
xnor U8891 (N_8891,N_7196,N_6009);
and U8892 (N_8892,N_5138,N_7107);
and U8893 (N_8893,N_6680,N_5382);
or U8894 (N_8894,N_5837,N_6306);
or U8895 (N_8895,N_5604,N_5069);
nand U8896 (N_8896,N_6304,N_5647);
and U8897 (N_8897,N_5331,N_6160);
and U8898 (N_8898,N_6470,N_6523);
nand U8899 (N_8899,N_6563,N_6173);
and U8900 (N_8900,N_5268,N_5165);
nor U8901 (N_8901,N_6990,N_6565);
or U8902 (N_8902,N_5428,N_5784);
nand U8903 (N_8903,N_5803,N_5076);
or U8904 (N_8904,N_7174,N_5396);
or U8905 (N_8905,N_5479,N_6723);
nand U8906 (N_8906,N_5949,N_6141);
or U8907 (N_8907,N_7281,N_7420);
nor U8908 (N_8908,N_5123,N_5005);
nand U8909 (N_8909,N_5206,N_6234);
nand U8910 (N_8910,N_5809,N_7458);
and U8911 (N_8911,N_5234,N_6646);
and U8912 (N_8912,N_7068,N_5125);
and U8913 (N_8913,N_6073,N_5141);
xnor U8914 (N_8914,N_5951,N_5255);
nor U8915 (N_8915,N_5190,N_7325);
nand U8916 (N_8916,N_6030,N_7327);
and U8917 (N_8917,N_6196,N_6242);
or U8918 (N_8918,N_6610,N_7381);
and U8919 (N_8919,N_6063,N_6942);
and U8920 (N_8920,N_5751,N_6430);
nand U8921 (N_8921,N_5016,N_6139);
and U8922 (N_8922,N_6122,N_6912);
and U8923 (N_8923,N_6182,N_5699);
or U8924 (N_8924,N_6150,N_5512);
nand U8925 (N_8925,N_6615,N_6308);
nor U8926 (N_8926,N_6972,N_7147);
nor U8927 (N_8927,N_6730,N_5490);
nand U8928 (N_8928,N_7199,N_7395);
nand U8929 (N_8929,N_7034,N_6085);
nor U8930 (N_8930,N_5646,N_6589);
nand U8931 (N_8931,N_5688,N_5369);
and U8932 (N_8932,N_5141,N_6836);
nand U8933 (N_8933,N_6988,N_6243);
nor U8934 (N_8934,N_6191,N_5371);
and U8935 (N_8935,N_6627,N_5990);
nor U8936 (N_8936,N_5397,N_6247);
or U8937 (N_8937,N_6242,N_6451);
nand U8938 (N_8938,N_7234,N_5296);
xnor U8939 (N_8939,N_6037,N_7172);
and U8940 (N_8940,N_7268,N_7030);
xnor U8941 (N_8941,N_6017,N_5048);
and U8942 (N_8942,N_6925,N_5189);
or U8943 (N_8943,N_7237,N_5642);
nor U8944 (N_8944,N_6770,N_6746);
nand U8945 (N_8945,N_6831,N_7151);
nor U8946 (N_8946,N_5688,N_5516);
and U8947 (N_8947,N_6639,N_5630);
and U8948 (N_8948,N_6799,N_6358);
and U8949 (N_8949,N_5569,N_6161);
nand U8950 (N_8950,N_6947,N_5574);
or U8951 (N_8951,N_7275,N_5859);
nand U8952 (N_8952,N_6419,N_5495);
and U8953 (N_8953,N_6063,N_7183);
nand U8954 (N_8954,N_5029,N_5687);
nor U8955 (N_8955,N_5028,N_7412);
nand U8956 (N_8956,N_6987,N_5924);
or U8957 (N_8957,N_7072,N_6652);
and U8958 (N_8958,N_5656,N_5757);
xor U8959 (N_8959,N_5133,N_6223);
and U8960 (N_8960,N_5187,N_6345);
or U8961 (N_8961,N_5764,N_6258);
nor U8962 (N_8962,N_6964,N_5639);
and U8963 (N_8963,N_5869,N_5954);
nor U8964 (N_8964,N_5286,N_5400);
or U8965 (N_8965,N_6110,N_7417);
or U8966 (N_8966,N_7461,N_7110);
nand U8967 (N_8967,N_7494,N_5221);
nor U8968 (N_8968,N_5904,N_5787);
nand U8969 (N_8969,N_5536,N_5032);
nand U8970 (N_8970,N_6493,N_6929);
nand U8971 (N_8971,N_7164,N_6265);
nor U8972 (N_8972,N_7180,N_5513);
or U8973 (N_8973,N_7394,N_5130);
nor U8974 (N_8974,N_5347,N_5280);
and U8975 (N_8975,N_5870,N_6078);
nor U8976 (N_8976,N_6933,N_6777);
nor U8977 (N_8977,N_5660,N_6088);
or U8978 (N_8978,N_7312,N_6978);
or U8979 (N_8979,N_6936,N_6204);
or U8980 (N_8980,N_7020,N_6177);
or U8981 (N_8981,N_7213,N_6613);
nor U8982 (N_8982,N_5600,N_6035);
or U8983 (N_8983,N_6705,N_5224);
and U8984 (N_8984,N_5169,N_5539);
nor U8985 (N_8985,N_5732,N_5864);
nand U8986 (N_8986,N_5133,N_6295);
nor U8987 (N_8987,N_7465,N_7386);
xor U8988 (N_8988,N_5257,N_5390);
or U8989 (N_8989,N_7030,N_6174);
and U8990 (N_8990,N_7315,N_6428);
nand U8991 (N_8991,N_5988,N_5029);
and U8992 (N_8992,N_5375,N_6730);
and U8993 (N_8993,N_6988,N_6376);
xnor U8994 (N_8994,N_6706,N_5647);
nand U8995 (N_8995,N_6902,N_7327);
nand U8996 (N_8996,N_6914,N_5771);
and U8997 (N_8997,N_6201,N_5025);
nand U8998 (N_8998,N_5523,N_5518);
and U8999 (N_8999,N_7088,N_6284);
nor U9000 (N_9000,N_6668,N_7385);
or U9001 (N_9001,N_7423,N_5372);
nand U9002 (N_9002,N_5688,N_6660);
and U9003 (N_9003,N_6414,N_6609);
xor U9004 (N_9004,N_6278,N_5223);
nor U9005 (N_9005,N_6272,N_6320);
and U9006 (N_9006,N_6621,N_5030);
nor U9007 (N_9007,N_6118,N_5675);
nand U9008 (N_9008,N_5617,N_6083);
and U9009 (N_9009,N_5107,N_6579);
nor U9010 (N_9010,N_5488,N_7152);
and U9011 (N_9011,N_5494,N_6058);
nor U9012 (N_9012,N_5943,N_7310);
and U9013 (N_9013,N_7485,N_6694);
and U9014 (N_9014,N_7221,N_7170);
nand U9015 (N_9015,N_6094,N_5140);
or U9016 (N_9016,N_6877,N_7020);
nor U9017 (N_9017,N_6154,N_6665);
and U9018 (N_9018,N_5255,N_5215);
nand U9019 (N_9019,N_6583,N_7090);
or U9020 (N_9020,N_5960,N_5289);
and U9021 (N_9021,N_5956,N_6648);
nand U9022 (N_9022,N_6246,N_6725);
nor U9023 (N_9023,N_5866,N_5187);
nor U9024 (N_9024,N_6083,N_5057);
or U9025 (N_9025,N_6145,N_7020);
or U9026 (N_9026,N_5506,N_6740);
and U9027 (N_9027,N_6434,N_5981);
nand U9028 (N_9028,N_6096,N_6241);
nor U9029 (N_9029,N_5758,N_5285);
or U9030 (N_9030,N_7195,N_5628);
or U9031 (N_9031,N_5450,N_5329);
or U9032 (N_9032,N_5539,N_6887);
and U9033 (N_9033,N_5039,N_6574);
nand U9034 (N_9034,N_6725,N_5857);
and U9035 (N_9035,N_5403,N_6664);
and U9036 (N_9036,N_6884,N_6174);
nor U9037 (N_9037,N_5973,N_7356);
nand U9038 (N_9038,N_6391,N_7042);
nor U9039 (N_9039,N_5149,N_5093);
xnor U9040 (N_9040,N_5531,N_5775);
or U9041 (N_9041,N_6340,N_6272);
or U9042 (N_9042,N_7228,N_6289);
and U9043 (N_9043,N_6933,N_5843);
or U9044 (N_9044,N_5498,N_5682);
or U9045 (N_9045,N_6958,N_6118);
nor U9046 (N_9046,N_7392,N_5893);
nand U9047 (N_9047,N_5635,N_6585);
nor U9048 (N_9048,N_5527,N_7179);
or U9049 (N_9049,N_6962,N_5845);
and U9050 (N_9050,N_6381,N_6492);
or U9051 (N_9051,N_5679,N_5408);
nor U9052 (N_9052,N_5007,N_6636);
xor U9053 (N_9053,N_5042,N_5076);
and U9054 (N_9054,N_7325,N_5907);
nor U9055 (N_9055,N_6356,N_6340);
and U9056 (N_9056,N_6826,N_6812);
and U9057 (N_9057,N_6875,N_5295);
xor U9058 (N_9058,N_5102,N_6019);
nand U9059 (N_9059,N_6160,N_6892);
nand U9060 (N_9060,N_6207,N_5911);
nor U9061 (N_9061,N_7058,N_6999);
and U9062 (N_9062,N_6239,N_5329);
xnor U9063 (N_9063,N_6035,N_5943);
nand U9064 (N_9064,N_5397,N_5174);
nor U9065 (N_9065,N_6359,N_5046);
and U9066 (N_9066,N_6953,N_6710);
nand U9067 (N_9067,N_5771,N_6779);
nand U9068 (N_9068,N_7226,N_5630);
nor U9069 (N_9069,N_7490,N_5774);
and U9070 (N_9070,N_5953,N_5982);
and U9071 (N_9071,N_6520,N_7374);
or U9072 (N_9072,N_6523,N_5212);
or U9073 (N_9073,N_5957,N_6478);
or U9074 (N_9074,N_5017,N_7135);
or U9075 (N_9075,N_5629,N_6074);
and U9076 (N_9076,N_7106,N_6311);
or U9077 (N_9077,N_5517,N_6750);
or U9078 (N_9078,N_7226,N_6631);
or U9079 (N_9079,N_6318,N_7440);
nor U9080 (N_9080,N_6616,N_5868);
or U9081 (N_9081,N_5370,N_6623);
nor U9082 (N_9082,N_6422,N_7320);
nand U9083 (N_9083,N_7090,N_6346);
or U9084 (N_9084,N_7454,N_5153);
nand U9085 (N_9085,N_7498,N_5581);
nand U9086 (N_9086,N_6346,N_5477);
nor U9087 (N_9087,N_5548,N_6497);
nor U9088 (N_9088,N_6507,N_7349);
nand U9089 (N_9089,N_7313,N_6648);
xnor U9090 (N_9090,N_7490,N_7414);
nor U9091 (N_9091,N_7269,N_5911);
nor U9092 (N_9092,N_6745,N_6789);
or U9093 (N_9093,N_5638,N_7391);
and U9094 (N_9094,N_6662,N_7408);
or U9095 (N_9095,N_6516,N_6169);
nand U9096 (N_9096,N_6921,N_5682);
and U9097 (N_9097,N_6117,N_5106);
and U9098 (N_9098,N_7221,N_5234);
or U9099 (N_9099,N_5868,N_5800);
xor U9100 (N_9100,N_5021,N_5868);
nand U9101 (N_9101,N_7381,N_7274);
nand U9102 (N_9102,N_6528,N_5995);
or U9103 (N_9103,N_5112,N_5152);
nor U9104 (N_9104,N_5281,N_5686);
and U9105 (N_9105,N_5954,N_5063);
xor U9106 (N_9106,N_5176,N_5357);
nand U9107 (N_9107,N_6095,N_7076);
or U9108 (N_9108,N_6662,N_5889);
nand U9109 (N_9109,N_6560,N_6324);
or U9110 (N_9110,N_7327,N_5726);
and U9111 (N_9111,N_7227,N_5897);
or U9112 (N_9112,N_7133,N_5274);
or U9113 (N_9113,N_5630,N_5859);
or U9114 (N_9114,N_6908,N_5168);
nand U9115 (N_9115,N_6707,N_5744);
nor U9116 (N_9116,N_6897,N_6056);
or U9117 (N_9117,N_6003,N_6664);
nand U9118 (N_9118,N_5031,N_6167);
or U9119 (N_9119,N_5347,N_5254);
and U9120 (N_9120,N_5654,N_7325);
nand U9121 (N_9121,N_5862,N_7206);
or U9122 (N_9122,N_7193,N_5828);
and U9123 (N_9123,N_5986,N_6731);
and U9124 (N_9124,N_5442,N_5256);
and U9125 (N_9125,N_5708,N_6320);
and U9126 (N_9126,N_5131,N_7022);
nor U9127 (N_9127,N_7329,N_7040);
or U9128 (N_9128,N_5810,N_5627);
or U9129 (N_9129,N_6890,N_7073);
nor U9130 (N_9130,N_7481,N_6357);
or U9131 (N_9131,N_6959,N_6137);
nor U9132 (N_9132,N_6404,N_6599);
nand U9133 (N_9133,N_6335,N_6942);
nand U9134 (N_9134,N_5488,N_5092);
or U9135 (N_9135,N_5601,N_6912);
and U9136 (N_9136,N_6456,N_5445);
nand U9137 (N_9137,N_6785,N_5799);
and U9138 (N_9138,N_6458,N_6837);
nand U9139 (N_9139,N_6222,N_6813);
xor U9140 (N_9140,N_5800,N_5392);
and U9141 (N_9141,N_6443,N_7328);
and U9142 (N_9142,N_6192,N_5647);
or U9143 (N_9143,N_6353,N_5939);
nor U9144 (N_9144,N_6344,N_5274);
or U9145 (N_9145,N_6572,N_5244);
or U9146 (N_9146,N_6935,N_5211);
nand U9147 (N_9147,N_6904,N_7337);
nand U9148 (N_9148,N_6920,N_6215);
nand U9149 (N_9149,N_5241,N_6108);
nor U9150 (N_9150,N_6268,N_5542);
or U9151 (N_9151,N_5002,N_6002);
and U9152 (N_9152,N_5219,N_7282);
nand U9153 (N_9153,N_6392,N_6333);
and U9154 (N_9154,N_7254,N_6659);
nor U9155 (N_9155,N_6496,N_7463);
nand U9156 (N_9156,N_5096,N_5309);
or U9157 (N_9157,N_5660,N_7489);
and U9158 (N_9158,N_5696,N_7416);
and U9159 (N_9159,N_7158,N_7477);
nand U9160 (N_9160,N_6762,N_6987);
nand U9161 (N_9161,N_5265,N_7483);
nor U9162 (N_9162,N_7357,N_5208);
nor U9163 (N_9163,N_5560,N_6070);
or U9164 (N_9164,N_5703,N_6866);
and U9165 (N_9165,N_5005,N_7228);
nor U9166 (N_9166,N_6430,N_6086);
xnor U9167 (N_9167,N_6589,N_5702);
nor U9168 (N_9168,N_6974,N_6651);
and U9169 (N_9169,N_6592,N_5100);
and U9170 (N_9170,N_7244,N_5950);
or U9171 (N_9171,N_6066,N_7124);
and U9172 (N_9172,N_5396,N_6839);
nor U9173 (N_9173,N_5733,N_5994);
nor U9174 (N_9174,N_5421,N_5286);
nand U9175 (N_9175,N_6892,N_6340);
nand U9176 (N_9176,N_5676,N_6369);
or U9177 (N_9177,N_6456,N_7186);
nor U9178 (N_9178,N_5198,N_7111);
nor U9179 (N_9179,N_5801,N_5808);
nor U9180 (N_9180,N_7348,N_7069);
nand U9181 (N_9181,N_6064,N_7098);
or U9182 (N_9182,N_7199,N_6644);
nor U9183 (N_9183,N_6333,N_7234);
nor U9184 (N_9184,N_6169,N_6080);
and U9185 (N_9185,N_5926,N_6037);
nor U9186 (N_9186,N_5715,N_5747);
nor U9187 (N_9187,N_7141,N_7309);
xor U9188 (N_9188,N_5308,N_5503);
and U9189 (N_9189,N_6309,N_6369);
nand U9190 (N_9190,N_6945,N_7198);
nand U9191 (N_9191,N_5015,N_5116);
or U9192 (N_9192,N_6103,N_5233);
nor U9193 (N_9193,N_6616,N_6612);
nand U9194 (N_9194,N_5383,N_6710);
and U9195 (N_9195,N_6956,N_6089);
and U9196 (N_9196,N_5273,N_7009);
or U9197 (N_9197,N_5454,N_6292);
nand U9198 (N_9198,N_6078,N_5475);
nand U9199 (N_9199,N_6411,N_7238);
or U9200 (N_9200,N_5994,N_6898);
or U9201 (N_9201,N_5421,N_6178);
or U9202 (N_9202,N_5268,N_7184);
nor U9203 (N_9203,N_7075,N_6370);
nand U9204 (N_9204,N_5404,N_5658);
and U9205 (N_9205,N_7437,N_5608);
nand U9206 (N_9206,N_5985,N_7231);
nand U9207 (N_9207,N_7439,N_7382);
nand U9208 (N_9208,N_5099,N_5146);
or U9209 (N_9209,N_5449,N_5139);
nor U9210 (N_9210,N_5326,N_6283);
nor U9211 (N_9211,N_5481,N_5570);
or U9212 (N_9212,N_6151,N_6291);
nor U9213 (N_9213,N_6910,N_6122);
nor U9214 (N_9214,N_6131,N_6877);
or U9215 (N_9215,N_6778,N_5743);
xor U9216 (N_9216,N_5093,N_5525);
or U9217 (N_9217,N_7088,N_7168);
nand U9218 (N_9218,N_6220,N_7361);
or U9219 (N_9219,N_6546,N_5985);
nand U9220 (N_9220,N_6489,N_7272);
and U9221 (N_9221,N_5202,N_6342);
and U9222 (N_9222,N_5445,N_6642);
nor U9223 (N_9223,N_7287,N_6238);
and U9224 (N_9224,N_6407,N_5607);
and U9225 (N_9225,N_7235,N_7258);
or U9226 (N_9226,N_6347,N_5063);
nand U9227 (N_9227,N_6615,N_6639);
nand U9228 (N_9228,N_6117,N_5207);
nor U9229 (N_9229,N_6301,N_5542);
nor U9230 (N_9230,N_5428,N_7070);
or U9231 (N_9231,N_7076,N_5683);
nand U9232 (N_9232,N_6376,N_5347);
nor U9233 (N_9233,N_6646,N_5952);
nor U9234 (N_9234,N_5797,N_6148);
nand U9235 (N_9235,N_6516,N_7208);
nor U9236 (N_9236,N_6821,N_7095);
or U9237 (N_9237,N_5174,N_6672);
and U9238 (N_9238,N_5886,N_6212);
nand U9239 (N_9239,N_5888,N_6510);
nor U9240 (N_9240,N_5054,N_6548);
nor U9241 (N_9241,N_5423,N_6873);
nand U9242 (N_9242,N_6442,N_6160);
xnor U9243 (N_9243,N_5654,N_5687);
nand U9244 (N_9244,N_6122,N_7186);
and U9245 (N_9245,N_5859,N_6523);
and U9246 (N_9246,N_5784,N_5150);
or U9247 (N_9247,N_6966,N_6029);
or U9248 (N_9248,N_6089,N_6304);
nand U9249 (N_9249,N_5129,N_6541);
nand U9250 (N_9250,N_7032,N_5149);
xor U9251 (N_9251,N_6740,N_7130);
xnor U9252 (N_9252,N_7293,N_6658);
nand U9253 (N_9253,N_7070,N_6312);
and U9254 (N_9254,N_5474,N_6896);
nor U9255 (N_9255,N_5000,N_5310);
nor U9256 (N_9256,N_7414,N_5536);
nor U9257 (N_9257,N_6043,N_5783);
or U9258 (N_9258,N_6447,N_7018);
or U9259 (N_9259,N_6902,N_6289);
nor U9260 (N_9260,N_5549,N_6367);
nor U9261 (N_9261,N_5018,N_6839);
or U9262 (N_9262,N_5131,N_7067);
and U9263 (N_9263,N_6888,N_5500);
nand U9264 (N_9264,N_6316,N_6834);
or U9265 (N_9265,N_5679,N_6323);
and U9266 (N_9266,N_5245,N_7025);
and U9267 (N_9267,N_5059,N_6191);
or U9268 (N_9268,N_6637,N_6031);
nand U9269 (N_9269,N_6889,N_5151);
nand U9270 (N_9270,N_6943,N_5661);
or U9271 (N_9271,N_5475,N_6748);
or U9272 (N_9272,N_5654,N_6637);
nand U9273 (N_9273,N_5617,N_5711);
nor U9274 (N_9274,N_6070,N_5043);
and U9275 (N_9275,N_5945,N_5030);
nand U9276 (N_9276,N_5280,N_7292);
and U9277 (N_9277,N_5490,N_5288);
or U9278 (N_9278,N_7053,N_5729);
nor U9279 (N_9279,N_7338,N_5329);
or U9280 (N_9280,N_7075,N_5056);
or U9281 (N_9281,N_5417,N_7479);
and U9282 (N_9282,N_5953,N_5526);
nor U9283 (N_9283,N_6324,N_5250);
or U9284 (N_9284,N_5433,N_5693);
nand U9285 (N_9285,N_7043,N_5330);
or U9286 (N_9286,N_5895,N_5536);
or U9287 (N_9287,N_6229,N_6481);
nor U9288 (N_9288,N_5006,N_6216);
or U9289 (N_9289,N_6358,N_5844);
or U9290 (N_9290,N_6988,N_5794);
nand U9291 (N_9291,N_5349,N_6413);
and U9292 (N_9292,N_5111,N_6471);
and U9293 (N_9293,N_5415,N_6459);
nor U9294 (N_9294,N_5043,N_7344);
nor U9295 (N_9295,N_5062,N_7378);
xor U9296 (N_9296,N_6290,N_5595);
or U9297 (N_9297,N_6164,N_7240);
and U9298 (N_9298,N_5964,N_5638);
nor U9299 (N_9299,N_5342,N_7147);
xnor U9300 (N_9300,N_5526,N_5391);
and U9301 (N_9301,N_7210,N_7238);
and U9302 (N_9302,N_7041,N_5196);
and U9303 (N_9303,N_5099,N_5532);
and U9304 (N_9304,N_6512,N_5228);
nor U9305 (N_9305,N_6992,N_6561);
nor U9306 (N_9306,N_5371,N_5288);
and U9307 (N_9307,N_7484,N_6341);
nor U9308 (N_9308,N_7396,N_6515);
nand U9309 (N_9309,N_5712,N_7025);
and U9310 (N_9310,N_5960,N_5123);
nand U9311 (N_9311,N_5838,N_5854);
and U9312 (N_9312,N_5394,N_6568);
nand U9313 (N_9313,N_5690,N_5405);
or U9314 (N_9314,N_6204,N_6440);
or U9315 (N_9315,N_6707,N_5705);
nor U9316 (N_9316,N_5242,N_5202);
xnor U9317 (N_9317,N_5110,N_5556);
nand U9318 (N_9318,N_7337,N_5412);
nand U9319 (N_9319,N_5406,N_7412);
or U9320 (N_9320,N_7006,N_7130);
xnor U9321 (N_9321,N_6966,N_5474);
or U9322 (N_9322,N_5280,N_6744);
or U9323 (N_9323,N_5449,N_5630);
nor U9324 (N_9324,N_7324,N_5102);
nor U9325 (N_9325,N_5461,N_5102);
or U9326 (N_9326,N_5594,N_6350);
and U9327 (N_9327,N_6601,N_5684);
and U9328 (N_9328,N_7179,N_7036);
nor U9329 (N_9329,N_6683,N_6573);
and U9330 (N_9330,N_7011,N_6303);
and U9331 (N_9331,N_5138,N_5888);
nand U9332 (N_9332,N_6703,N_6277);
or U9333 (N_9333,N_6678,N_7124);
or U9334 (N_9334,N_5441,N_6757);
and U9335 (N_9335,N_6538,N_6365);
nand U9336 (N_9336,N_5051,N_5947);
nor U9337 (N_9337,N_7056,N_7342);
and U9338 (N_9338,N_6626,N_5871);
nor U9339 (N_9339,N_7199,N_6709);
nor U9340 (N_9340,N_7469,N_5072);
xor U9341 (N_9341,N_7428,N_6935);
xnor U9342 (N_9342,N_7272,N_6120);
or U9343 (N_9343,N_7256,N_6454);
or U9344 (N_9344,N_6903,N_5230);
and U9345 (N_9345,N_6950,N_6452);
nand U9346 (N_9346,N_5084,N_5976);
nand U9347 (N_9347,N_7221,N_7313);
and U9348 (N_9348,N_5518,N_5539);
and U9349 (N_9349,N_7415,N_7371);
nor U9350 (N_9350,N_6497,N_7173);
and U9351 (N_9351,N_5519,N_7150);
and U9352 (N_9352,N_5449,N_6828);
nand U9353 (N_9353,N_5169,N_6031);
nand U9354 (N_9354,N_7498,N_6912);
nor U9355 (N_9355,N_7366,N_7028);
and U9356 (N_9356,N_5273,N_6988);
nor U9357 (N_9357,N_6710,N_6806);
or U9358 (N_9358,N_7357,N_5491);
nor U9359 (N_9359,N_6728,N_7310);
and U9360 (N_9360,N_5369,N_7066);
nor U9361 (N_9361,N_5062,N_7306);
nand U9362 (N_9362,N_5139,N_5781);
nor U9363 (N_9363,N_5754,N_6916);
or U9364 (N_9364,N_5026,N_6393);
nor U9365 (N_9365,N_5219,N_6508);
xor U9366 (N_9366,N_6638,N_6469);
or U9367 (N_9367,N_6221,N_6931);
nand U9368 (N_9368,N_6467,N_5025);
nor U9369 (N_9369,N_6451,N_5218);
nor U9370 (N_9370,N_5805,N_6507);
and U9371 (N_9371,N_6785,N_6083);
and U9372 (N_9372,N_5380,N_5711);
or U9373 (N_9373,N_6628,N_5972);
nor U9374 (N_9374,N_6742,N_6728);
nand U9375 (N_9375,N_7253,N_5829);
and U9376 (N_9376,N_6665,N_5556);
or U9377 (N_9377,N_5767,N_5532);
or U9378 (N_9378,N_7252,N_6889);
and U9379 (N_9379,N_7029,N_5743);
and U9380 (N_9380,N_6780,N_7147);
nor U9381 (N_9381,N_5711,N_5099);
nand U9382 (N_9382,N_6766,N_5634);
nand U9383 (N_9383,N_6773,N_5204);
or U9384 (N_9384,N_6770,N_5624);
nand U9385 (N_9385,N_6635,N_5063);
or U9386 (N_9386,N_6408,N_5766);
nand U9387 (N_9387,N_6039,N_5184);
nor U9388 (N_9388,N_7017,N_6016);
nand U9389 (N_9389,N_7348,N_6623);
or U9390 (N_9390,N_6887,N_6869);
or U9391 (N_9391,N_5108,N_7419);
or U9392 (N_9392,N_6627,N_6690);
nand U9393 (N_9393,N_7220,N_5585);
and U9394 (N_9394,N_7061,N_6741);
or U9395 (N_9395,N_5778,N_5954);
and U9396 (N_9396,N_5847,N_6875);
nand U9397 (N_9397,N_5649,N_6115);
or U9398 (N_9398,N_6295,N_5894);
and U9399 (N_9399,N_5433,N_5344);
and U9400 (N_9400,N_7463,N_6251);
and U9401 (N_9401,N_6056,N_5271);
and U9402 (N_9402,N_5307,N_5399);
nor U9403 (N_9403,N_5847,N_5134);
or U9404 (N_9404,N_6797,N_6853);
nand U9405 (N_9405,N_5845,N_7094);
nand U9406 (N_9406,N_6295,N_5447);
or U9407 (N_9407,N_6104,N_5007);
and U9408 (N_9408,N_6854,N_5660);
nand U9409 (N_9409,N_5488,N_6871);
nor U9410 (N_9410,N_6815,N_5138);
or U9411 (N_9411,N_6389,N_5683);
nand U9412 (N_9412,N_7403,N_6888);
nor U9413 (N_9413,N_5843,N_6828);
nor U9414 (N_9414,N_7433,N_7368);
nor U9415 (N_9415,N_5148,N_5495);
and U9416 (N_9416,N_6849,N_6246);
nor U9417 (N_9417,N_5627,N_7035);
and U9418 (N_9418,N_6894,N_6794);
and U9419 (N_9419,N_6857,N_6158);
or U9420 (N_9420,N_5021,N_5002);
and U9421 (N_9421,N_7036,N_6829);
and U9422 (N_9422,N_6630,N_5721);
or U9423 (N_9423,N_6918,N_5387);
and U9424 (N_9424,N_5134,N_6111);
or U9425 (N_9425,N_6735,N_6820);
and U9426 (N_9426,N_5066,N_6339);
or U9427 (N_9427,N_5704,N_5091);
nand U9428 (N_9428,N_5179,N_5259);
nand U9429 (N_9429,N_6208,N_6559);
nand U9430 (N_9430,N_6600,N_6535);
or U9431 (N_9431,N_5776,N_5968);
or U9432 (N_9432,N_6121,N_6087);
nand U9433 (N_9433,N_5119,N_6201);
xor U9434 (N_9434,N_6440,N_6514);
nor U9435 (N_9435,N_5102,N_5958);
nand U9436 (N_9436,N_6446,N_6484);
nand U9437 (N_9437,N_6593,N_5431);
nand U9438 (N_9438,N_6403,N_5106);
nand U9439 (N_9439,N_7086,N_7028);
and U9440 (N_9440,N_6923,N_7073);
or U9441 (N_9441,N_7402,N_5340);
or U9442 (N_9442,N_6566,N_5752);
or U9443 (N_9443,N_6822,N_5491);
and U9444 (N_9444,N_5891,N_5608);
or U9445 (N_9445,N_5100,N_6717);
nor U9446 (N_9446,N_6359,N_5059);
nand U9447 (N_9447,N_5251,N_7375);
nand U9448 (N_9448,N_6398,N_7490);
nand U9449 (N_9449,N_5319,N_6899);
or U9450 (N_9450,N_5173,N_7144);
nand U9451 (N_9451,N_6419,N_5152);
and U9452 (N_9452,N_5062,N_6700);
and U9453 (N_9453,N_6181,N_5620);
and U9454 (N_9454,N_5775,N_5159);
and U9455 (N_9455,N_7238,N_5395);
and U9456 (N_9456,N_6248,N_5610);
nand U9457 (N_9457,N_7458,N_5128);
and U9458 (N_9458,N_5621,N_5778);
nand U9459 (N_9459,N_5584,N_6935);
nor U9460 (N_9460,N_5427,N_5618);
nor U9461 (N_9461,N_6988,N_7041);
or U9462 (N_9462,N_6875,N_5258);
or U9463 (N_9463,N_5754,N_6316);
nand U9464 (N_9464,N_6418,N_6001);
nand U9465 (N_9465,N_6199,N_5142);
nand U9466 (N_9466,N_7408,N_5261);
or U9467 (N_9467,N_6221,N_7446);
xor U9468 (N_9468,N_6630,N_6392);
nand U9469 (N_9469,N_5263,N_6268);
and U9470 (N_9470,N_5895,N_5328);
nand U9471 (N_9471,N_5186,N_5592);
nand U9472 (N_9472,N_5181,N_6159);
nand U9473 (N_9473,N_6485,N_6933);
and U9474 (N_9474,N_6137,N_5880);
or U9475 (N_9475,N_7459,N_5991);
nand U9476 (N_9476,N_5272,N_5664);
and U9477 (N_9477,N_7237,N_6888);
xnor U9478 (N_9478,N_6810,N_6171);
or U9479 (N_9479,N_5195,N_6544);
and U9480 (N_9480,N_6825,N_7238);
xor U9481 (N_9481,N_6921,N_6404);
nor U9482 (N_9482,N_5824,N_6063);
or U9483 (N_9483,N_5353,N_7292);
or U9484 (N_9484,N_5939,N_7003);
nor U9485 (N_9485,N_5551,N_7188);
nor U9486 (N_9486,N_5482,N_5831);
or U9487 (N_9487,N_7103,N_6133);
nand U9488 (N_9488,N_5855,N_6476);
or U9489 (N_9489,N_6106,N_6275);
nor U9490 (N_9490,N_6077,N_6555);
and U9491 (N_9491,N_5437,N_6287);
nor U9492 (N_9492,N_5728,N_6360);
and U9493 (N_9493,N_6640,N_6454);
nor U9494 (N_9494,N_5770,N_6220);
and U9495 (N_9495,N_5903,N_5120);
nor U9496 (N_9496,N_6280,N_7042);
and U9497 (N_9497,N_7113,N_5976);
nor U9498 (N_9498,N_7155,N_5023);
nand U9499 (N_9499,N_5117,N_7426);
and U9500 (N_9500,N_6680,N_6312);
nor U9501 (N_9501,N_5015,N_7115);
nand U9502 (N_9502,N_6915,N_7028);
or U9503 (N_9503,N_5934,N_6435);
nor U9504 (N_9504,N_6485,N_6803);
and U9505 (N_9505,N_6217,N_6614);
and U9506 (N_9506,N_7361,N_5100);
and U9507 (N_9507,N_6064,N_6632);
nand U9508 (N_9508,N_6518,N_5534);
or U9509 (N_9509,N_6828,N_5696);
nand U9510 (N_9510,N_6928,N_7090);
nor U9511 (N_9511,N_5462,N_6154);
nand U9512 (N_9512,N_6373,N_7308);
nand U9513 (N_9513,N_7057,N_6759);
nor U9514 (N_9514,N_5679,N_5337);
and U9515 (N_9515,N_6343,N_6598);
and U9516 (N_9516,N_7014,N_5393);
nand U9517 (N_9517,N_5218,N_6260);
and U9518 (N_9518,N_7470,N_6022);
nor U9519 (N_9519,N_6430,N_5832);
and U9520 (N_9520,N_5114,N_7334);
nor U9521 (N_9521,N_7105,N_5852);
and U9522 (N_9522,N_6412,N_6942);
and U9523 (N_9523,N_5605,N_6419);
or U9524 (N_9524,N_6336,N_6526);
nand U9525 (N_9525,N_5907,N_5659);
nor U9526 (N_9526,N_6485,N_5234);
nor U9527 (N_9527,N_5002,N_6711);
and U9528 (N_9528,N_7094,N_6571);
or U9529 (N_9529,N_6567,N_6630);
nor U9530 (N_9530,N_5159,N_7458);
and U9531 (N_9531,N_5799,N_7116);
nor U9532 (N_9532,N_7319,N_5480);
nand U9533 (N_9533,N_7047,N_5519);
and U9534 (N_9534,N_6137,N_6249);
nand U9535 (N_9535,N_5431,N_7046);
nand U9536 (N_9536,N_7446,N_6036);
nor U9537 (N_9537,N_5193,N_5948);
nor U9538 (N_9538,N_6318,N_6633);
or U9539 (N_9539,N_6349,N_6219);
or U9540 (N_9540,N_6500,N_5249);
or U9541 (N_9541,N_5668,N_7155);
or U9542 (N_9542,N_6897,N_6306);
nor U9543 (N_9543,N_6293,N_6213);
nor U9544 (N_9544,N_5979,N_7047);
nor U9545 (N_9545,N_7416,N_5893);
nand U9546 (N_9546,N_5859,N_6893);
and U9547 (N_9547,N_6268,N_6069);
nand U9548 (N_9548,N_6440,N_6233);
nor U9549 (N_9549,N_5421,N_6966);
and U9550 (N_9550,N_5303,N_7063);
or U9551 (N_9551,N_5771,N_6535);
or U9552 (N_9552,N_6041,N_6850);
nand U9553 (N_9553,N_5596,N_5420);
nand U9554 (N_9554,N_6022,N_5530);
and U9555 (N_9555,N_6574,N_5454);
nand U9556 (N_9556,N_6019,N_6557);
or U9557 (N_9557,N_6569,N_6468);
or U9558 (N_9558,N_7321,N_6889);
and U9559 (N_9559,N_6108,N_6071);
and U9560 (N_9560,N_5827,N_5763);
and U9561 (N_9561,N_6613,N_6203);
or U9562 (N_9562,N_5509,N_5857);
and U9563 (N_9563,N_5399,N_5452);
nor U9564 (N_9564,N_5577,N_7093);
nand U9565 (N_9565,N_7363,N_5696);
xor U9566 (N_9566,N_6968,N_6870);
or U9567 (N_9567,N_7483,N_5315);
xnor U9568 (N_9568,N_7026,N_6820);
or U9569 (N_9569,N_6926,N_5862);
and U9570 (N_9570,N_6421,N_5561);
or U9571 (N_9571,N_7371,N_6547);
and U9572 (N_9572,N_6034,N_5990);
nand U9573 (N_9573,N_6754,N_5698);
nor U9574 (N_9574,N_6281,N_7306);
or U9575 (N_9575,N_6705,N_7386);
nand U9576 (N_9576,N_6816,N_6268);
and U9577 (N_9577,N_6025,N_5959);
nand U9578 (N_9578,N_6640,N_7205);
and U9579 (N_9579,N_7393,N_6506);
nand U9580 (N_9580,N_5884,N_7463);
or U9581 (N_9581,N_5442,N_6514);
nor U9582 (N_9582,N_7056,N_6206);
or U9583 (N_9583,N_7469,N_7398);
nor U9584 (N_9584,N_5315,N_6183);
and U9585 (N_9585,N_5261,N_5698);
nand U9586 (N_9586,N_6676,N_5897);
or U9587 (N_9587,N_6468,N_7111);
or U9588 (N_9588,N_6580,N_5836);
nand U9589 (N_9589,N_5263,N_5751);
and U9590 (N_9590,N_5456,N_7170);
nor U9591 (N_9591,N_5124,N_7069);
or U9592 (N_9592,N_7175,N_6313);
nor U9593 (N_9593,N_5646,N_5677);
and U9594 (N_9594,N_6200,N_5730);
nor U9595 (N_9595,N_5502,N_5152);
or U9596 (N_9596,N_7137,N_6767);
and U9597 (N_9597,N_6893,N_6988);
nand U9598 (N_9598,N_5903,N_6180);
and U9599 (N_9599,N_7289,N_5390);
and U9600 (N_9600,N_6520,N_5822);
or U9601 (N_9601,N_6348,N_5623);
nor U9602 (N_9602,N_6457,N_6167);
or U9603 (N_9603,N_5246,N_7467);
nand U9604 (N_9604,N_5866,N_7119);
nand U9605 (N_9605,N_5920,N_6712);
and U9606 (N_9606,N_6415,N_5952);
or U9607 (N_9607,N_7034,N_5811);
and U9608 (N_9608,N_5620,N_6455);
or U9609 (N_9609,N_6281,N_6664);
nand U9610 (N_9610,N_7311,N_5482);
nand U9611 (N_9611,N_6994,N_5774);
or U9612 (N_9612,N_7260,N_5059);
or U9613 (N_9613,N_5941,N_6753);
nor U9614 (N_9614,N_5062,N_7249);
nand U9615 (N_9615,N_6411,N_5981);
nor U9616 (N_9616,N_6283,N_5334);
or U9617 (N_9617,N_6021,N_6927);
nand U9618 (N_9618,N_5551,N_6380);
nand U9619 (N_9619,N_6780,N_5828);
nand U9620 (N_9620,N_6253,N_6843);
or U9621 (N_9621,N_6110,N_5864);
and U9622 (N_9622,N_6587,N_6797);
or U9623 (N_9623,N_5150,N_6131);
nor U9624 (N_9624,N_6629,N_5740);
and U9625 (N_9625,N_5123,N_5050);
nand U9626 (N_9626,N_5009,N_6784);
and U9627 (N_9627,N_5473,N_6109);
nor U9628 (N_9628,N_6995,N_6415);
xor U9629 (N_9629,N_5643,N_6758);
nor U9630 (N_9630,N_6564,N_5214);
and U9631 (N_9631,N_5231,N_5986);
and U9632 (N_9632,N_6263,N_5168);
and U9633 (N_9633,N_6724,N_5407);
or U9634 (N_9634,N_5405,N_5040);
and U9635 (N_9635,N_7438,N_7117);
nand U9636 (N_9636,N_7464,N_6209);
nand U9637 (N_9637,N_5386,N_5059);
nand U9638 (N_9638,N_7241,N_5605);
and U9639 (N_9639,N_7227,N_7254);
and U9640 (N_9640,N_5850,N_6693);
nand U9641 (N_9641,N_7328,N_5678);
or U9642 (N_9642,N_5728,N_6874);
and U9643 (N_9643,N_6740,N_7239);
nor U9644 (N_9644,N_7016,N_7410);
and U9645 (N_9645,N_5616,N_6792);
nand U9646 (N_9646,N_5603,N_6429);
nand U9647 (N_9647,N_6508,N_5072);
or U9648 (N_9648,N_6833,N_7112);
nor U9649 (N_9649,N_5008,N_5934);
or U9650 (N_9650,N_7114,N_5455);
nor U9651 (N_9651,N_6950,N_6426);
or U9652 (N_9652,N_5273,N_7240);
nand U9653 (N_9653,N_6748,N_5688);
and U9654 (N_9654,N_5118,N_5257);
nand U9655 (N_9655,N_6551,N_6536);
or U9656 (N_9656,N_5791,N_5877);
and U9657 (N_9657,N_6382,N_6602);
nor U9658 (N_9658,N_6116,N_6461);
and U9659 (N_9659,N_5798,N_6566);
nor U9660 (N_9660,N_7022,N_5916);
nor U9661 (N_9661,N_6809,N_7004);
nor U9662 (N_9662,N_5801,N_5233);
or U9663 (N_9663,N_5218,N_5919);
nand U9664 (N_9664,N_6081,N_6923);
nand U9665 (N_9665,N_6063,N_5243);
and U9666 (N_9666,N_6820,N_7319);
and U9667 (N_9667,N_6011,N_7083);
nand U9668 (N_9668,N_5518,N_6816);
or U9669 (N_9669,N_6136,N_5612);
or U9670 (N_9670,N_5772,N_6806);
or U9671 (N_9671,N_7498,N_6752);
and U9672 (N_9672,N_7319,N_5350);
nand U9673 (N_9673,N_6591,N_5948);
or U9674 (N_9674,N_6574,N_7008);
or U9675 (N_9675,N_6036,N_5172);
and U9676 (N_9676,N_7321,N_6502);
nand U9677 (N_9677,N_6802,N_5454);
nand U9678 (N_9678,N_7066,N_5313);
xnor U9679 (N_9679,N_6896,N_7398);
and U9680 (N_9680,N_5646,N_6049);
nand U9681 (N_9681,N_7074,N_6262);
and U9682 (N_9682,N_5449,N_6408);
nand U9683 (N_9683,N_5538,N_6723);
or U9684 (N_9684,N_5751,N_6092);
or U9685 (N_9685,N_6190,N_5853);
xor U9686 (N_9686,N_6826,N_5919);
nor U9687 (N_9687,N_5578,N_5423);
nand U9688 (N_9688,N_7328,N_6466);
nand U9689 (N_9689,N_5019,N_6119);
nor U9690 (N_9690,N_5166,N_5862);
or U9691 (N_9691,N_5924,N_7216);
xnor U9692 (N_9692,N_7449,N_6182);
nand U9693 (N_9693,N_5205,N_6522);
and U9694 (N_9694,N_7364,N_5239);
nor U9695 (N_9695,N_6921,N_6463);
and U9696 (N_9696,N_5678,N_5629);
or U9697 (N_9697,N_5497,N_5712);
nor U9698 (N_9698,N_5782,N_7257);
nand U9699 (N_9699,N_6080,N_6337);
xnor U9700 (N_9700,N_5374,N_5603);
or U9701 (N_9701,N_6326,N_6258);
and U9702 (N_9702,N_5991,N_6853);
nand U9703 (N_9703,N_6729,N_5319);
and U9704 (N_9704,N_7496,N_6965);
nor U9705 (N_9705,N_5838,N_7389);
nand U9706 (N_9706,N_7157,N_6556);
nand U9707 (N_9707,N_6989,N_5179);
nor U9708 (N_9708,N_7225,N_5216);
nand U9709 (N_9709,N_7074,N_5448);
nand U9710 (N_9710,N_5814,N_7143);
or U9711 (N_9711,N_5026,N_6159);
nand U9712 (N_9712,N_7384,N_6013);
and U9713 (N_9713,N_5614,N_5958);
or U9714 (N_9714,N_7477,N_5754);
and U9715 (N_9715,N_5224,N_7376);
nand U9716 (N_9716,N_6590,N_6197);
or U9717 (N_9717,N_5229,N_5803);
or U9718 (N_9718,N_7359,N_5043);
nand U9719 (N_9719,N_7104,N_7202);
and U9720 (N_9720,N_6721,N_5408);
nor U9721 (N_9721,N_5416,N_7065);
or U9722 (N_9722,N_6914,N_6848);
nand U9723 (N_9723,N_6260,N_6879);
and U9724 (N_9724,N_6538,N_6927);
or U9725 (N_9725,N_6292,N_6276);
nor U9726 (N_9726,N_6576,N_5384);
and U9727 (N_9727,N_5553,N_7222);
nand U9728 (N_9728,N_5381,N_5023);
nor U9729 (N_9729,N_6549,N_5862);
nand U9730 (N_9730,N_5284,N_6808);
nand U9731 (N_9731,N_5128,N_7012);
nand U9732 (N_9732,N_5168,N_5919);
xor U9733 (N_9733,N_5244,N_6390);
or U9734 (N_9734,N_6541,N_5786);
nor U9735 (N_9735,N_7042,N_6728);
or U9736 (N_9736,N_7246,N_5328);
nand U9737 (N_9737,N_6970,N_7221);
nor U9738 (N_9738,N_5341,N_6642);
nand U9739 (N_9739,N_7292,N_7295);
nor U9740 (N_9740,N_5841,N_6744);
nand U9741 (N_9741,N_5030,N_7172);
or U9742 (N_9742,N_6252,N_6360);
and U9743 (N_9743,N_6209,N_6627);
nor U9744 (N_9744,N_5639,N_6199);
nor U9745 (N_9745,N_6508,N_5843);
xnor U9746 (N_9746,N_5481,N_6052);
xor U9747 (N_9747,N_6008,N_6940);
or U9748 (N_9748,N_5661,N_5488);
or U9749 (N_9749,N_5019,N_5666);
nand U9750 (N_9750,N_6927,N_5579);
xnor U9751 (N_9751,N_5327,N_5056);
nand U9752 (N_9752,N_6148,N_6359);
nor U9753 (N_9753,N_7238,N_6941);
nor U9754 (N_9754,N_6462,N_7080);
or U9755 (N_9755,N_5046,N_5040);
nor U9756 (N_9756,N_7163,N_5972);
nand U9757 (N_9757,N_5299,N_5858);
and U9758 (N_9758,N_6210,N_7302);
nor U9759 (N_9759,N_6490,N_6839);
nand U9760 (N_9760,N_6664,N_6323);
or U9761 (N_9761,N_6363,N_5653);
nor U9762 (N_9762,N_7224,N_6496);
or U9763 (N_9763,N_7110,N_5287);
and U9764 (N_9764,N_5877,N_6987);
nor U9765 (N_9765,N_6551,N_5275);
and U9766 (N_9766,N_5629,N_6147);
and U9767 (N_9767,N_6108,N_6755);
and U9768 (N_9768,N_6882,N_7178);
or U9769 (N_9769,N_6881,N_5840);
nand U9770 (N_9770,N_5059,N_6829);
and U9771 (N_9771,N_5752,N_6145);
or U9772 (N_9772,N_5393,N_7147);
and U9773 (N_9773,N_6854,N_6251);
nor U9774 (N_9774,N_5938,N_7414);
and U9775 (N_9775,N_6022,N_6939);
or U9776 (N_9776,N_6229,N_7248);
or U9777 (N_9777,N_6701,N_5751);
or U9778 (N_9778,N_6607,N_5087);
and U9779 (N_9779,N_6151,N_6803);
and U9780 (N_9780,N_7136,N_7135);
or U9781 (N_9781,N_7046,N_6620);
and U9782 (N_9782,N_5407,N_5502);
and U9783 (N_9783,N_7471,N_5851);
xor U9784 (N_9784,N_5924,N_5424);
nand U9785 (N_9785,N_5448,N_7300);
nand U9786 (N_9786,N_5231,N_7175);
nor U9787 (N_9787,N_5361,N_7059);
nand U9788 (N_9788,N_5993,N_6402);
nand U9789 (N_9789,N_6844,N_6777);
or U9790 (N_9790,N_6716,N_5364);
nor U9791 (N_9791,N_5797,N_5065);
nand U9792 (N_9792,N_5640,N_6720);
nor U9793 (N_9793,N_6953,N_5603);
nor U9794 (N_9794,N_6864,N_5418);
nor U9795 (N_9795,N_7270,N_5952);
or U9796 (N_9796,N_5264,N_5601);
xnor U9797 (N_9797,N_6026,N_7370);
and U9798 (N_9798,N_5797,N_5073);
nor U9799 (N_9799,N_6984,N_6544);
and U9800 (N_9800,N_7229,N_7432);
and U9801 (N_9801,N_6849,N_6743);
or U9802 (N_9802,N_7107,N_6618);
xor U9803 (N_9803,N_6631,N_5685);
nor U9804 (N_9804,N_6823,N_6700);
and U9805 (N_9805,N_5914,N_5699);
nor U9806 (N_9806,N_5987,N_6755);
xnor U9807 (N_9807,N_7281,N_5288);
nor U9808 (N_9808,N_5220,N_5083);
nor U9809 (N_9809,N_5363,N_5031);
nand U9810 (N_9810,N_5402,N_6523);
nor U9811 (N_9811,N_7126,N_7102);
nand U9812 (N_9812,N_6788,N_5215);
or U9813 (N_9813,N_5657,N_5846);
nor U9814 (N_9814,N_6288,N_7336);
nand U9815 (N_9815,N_5638,N_6695);
and U9816 (N_9816,N_7319,N_6618);
nand U9817 (N_9817,N_6925,N_5735);
and U9818 (N_9818,N_6393,N_6584);
nand U9819 (N_9819,N_6378,N_6599);
xor U9820 (N_9820,N_5090,N_5006);
nand U9821 (N_9821,N_6564,N_5470);
and U9822 (N_9822,N_5412,N_5634);
xnor U9823 (N_9823,N_5649,N_6102);
and U9824 (N_9824,N_6567,N_5846);
nor U9825 (N_9825,N_5213,N_5927);
nor U9826 (N_9826,N_5678,N_7482);
and U9827 (N_9827,N_5549,N_5116);
nand U9828 (N_9828,N_7076,N_7127);
xnor U9829 (N_9829,N_5994,N_5869);
nand U9830 (N_9830,N_6145,N_6293);
nor U9831 (N_9831,N_5761,N_7207);
or U9832 (N_9832,N_7221,N_6904);
nor U9833 (N_9833,N_5561,N_5522);
nor U9834 (N_9834,N_6189,N_7031);
nor U9835 (N_9835,N_5290,N_5912);
and U9836 (N_9836,N_5902,N_5880);
nand U9837 (N_9837,N_5996,N_5722);
or U9838 (N_9838,N_5375,N_5651);
and U9839 (N_9839,N_6657,N_6623);
nand U9840 (N_9840,N_6281,N_5682);
and U9841 (N_9841,N_6873,N_5861);
or U9842 (N_9842,N_5812,N_7238);
nand U9843 (N_9843,N_6186,N_6988);
nand U9844 (N_9844,N_5607,N_5080);
and U9845 (N_9845,N_6415,N_5150);
and U9846 (N_9846,N_5311,N_7110);
or U9847 (N_9847,N_6579,N_6016);
and U9848 (N_9848,N_5714,N_6470);
nor U9849 (N_9849,N_5105,N_5747);
or U9850 (N_9850,N_7489,N_5907);
or U9851 (N_9851,N_7295,N_7138);
nor U9852 (N_9852,N_6061,N_7107);
or U9853 (N_9853,N_7149,N_6280);
nor U9854 (N_9854,N_6670,N_5188);
nor U9855 (N_9855,N_7414,N_5219);
nor U9856 (N_9856,N_6260,N_5933);
or U9857 (N_9857,N_7479,N_6897);
or U9858 (N_9858,N_7429,N_6017);
and U9859 (N_9859,N_6686,N_6268);
or U9860 (N_9860,N_5441,N_5526);
and U9861 (N_9861,N_6834,N_6624);
nand U9862 (N_9862,N_6974,N_5502);
and U9863 (N_9863,N_5514,N_5140);
nand U9864 (N_9864,N_5860,N_6705);
and U9865 (N_9865,N_7259,N_6551);
or U9866 (N_9866,N_6503,N_5100);
and U9867 (N_9867,N_5421,N_6420);
or U9868 (N_9868,N_7302,N_5711);
nor U9869 (N_9869,N_7469,N_6756);
or U9870 (N_9870,N_6371,N_6657);
and U9871 (N_9871,N_5869,N_7248);
and U9872 (N_9872,N_6821,N_7206);
nor U9873 (N_9873,N_7125,N_7153);
and U9874 (N_9874,N_5275,N_6233);
nor U9875 (N_9875,N_6722,N_5243);
nand U9876 (N_9876,N_5590,N_5625);
nor U9877 (N_9877,N_6653,N_6153);
nand U9878 (N_9878,N_7091,N_6639);
nand U9879 (N_9879,N_5772,N_5746);
nor U9880 (N_9880,N_5705,N_5927);
and U9881 (N_9881,N_5893,N_5030);
nand U9882 (N_9882,N_5821,N_5072);
nand U9883 (N_9883,N_7272,N_6487);
xnor U9884 (N_9884,N_7145,N_7454);
nor U9885 (N_9885,N_6150,N_7479);
or U9886 (N_9886,N_5060,N_5871);
nor U9887 (N_9887,N_6832,N_6299);
or U9888 (N_9888,N_6556,N_5632);
nand U9889 (N_9889,N_6392,N_5720);
and U9890 (N_9890,N_7160,N_6688);
nor U9891 (N_9891,N_6373,N_6326);
and U9892 (N_9892,N_6171,N_5225);
or U9893 (N_9893,N_5082,N_7201);
nand U9894 (N_9894,N_5064,N_6205);
xnor U9895 (N_9895,N_6069,N_7138);
nor U9896 (N_9896,N_6772,N_6788);
and U9897 (N_9897,N_7118,N_5613);
or U9898 (N_9898,N_5502,N_7349);
nor U9899 (N_9899,N_6570,N_5375);
or U9900 (N_9900,N_5336,N_6271);
or U9901 (N_9901,N_7465,N_7432);
nor U9902 (N_9902,N_5510,N_5966);
nand U9903 (N_9903,N_6550,N_5814);
or U9904 (N_9904,N_5346,N_7164);
and U9905 (N_9905,N_6356,N_5461);
nor U9906 (N_9906,N_6597,N_7209);
nand U9907 (N_9907,N_7319,N_5750);
nor U9908 (N_9908,N_5939,N_7478);
or U9909 (N_9909,N_5834,N_7256);
nand U9910 (N_9910,N_5867,N_7423);
nand U9911 (N_9911,N_6040,N_6599);
or U9912 (N_9912,N_7483,N_6722);
xor U9913 (N_9913,N_5989,N_5768);
nor U9914 (N_9914,N_6351,N_6727);
nand U9915 (N_9915,N_5445,N_5947);
nand U9916 (N_9916,N_7425,N_6880);
and U9917 (N_9917,N_7081,N_5729);
nand U9918 (N_9918,N_5849,N_5582);
xor U9919 (N_9919,N_7022,N_6143);
and U9920 (N_9920,N_5281,N_5247);
or U9921 (N_9921,N_7260,N_5535);
or U9922 (N_9922,N_5789,N_7313);
and U9923 (N_9923,N_6276,N_5197);
or U9924 (N_9924,N_7109,N_5633);
nor U9925 (N_9925,N_5322,N_5766);
nor U9926 (N_9926,N_5822,N_6600);
nand U9927 (N_9927,N_7466,N_7124);
xor U9928 (N_9928,N_7407,N_6386);
nor U9929 (N_9929,N_7455,N_6108);
and U9930 (N_9930,N_5838,N_5796);
nor U9931 (N_9931,N_5538,N_6059);
or U9932 (N_9932,N_6635,N_6962);
nor U9933 (N_9933,N_5951,N_5598);
nor U9934 (N_9934,N_5261,N_6658);
and U9935 (N_9935,N_5233,N_5678);
and U9936 (N_9936,N_6475,N_7156);
or U9937 (N_9937,N_6156,N_6280);
or U9938 (N_9938,N_5786,N_6140);
nor U9939 (N_9939,N_5425,N_6773);
or U9940 (N_9940,N_6106,N_5867);
and U9941 (N_9941,N_6242,N_5807);
or U9942 (N_9942,N_6818,N_7161);
nor U9943 (N_9943,N_5095,N_7071);
nand U9944 (N_9944,N_6037,N_6191);
xnor U9945 (N_9945,N_6573,N_6639);
or U9946 (N_9946,N_5773,N_6173);
nor U9947 (N_9947,N_5182,N_5692);
nand U9948 (N_9948,N_7201,N_6941);
and U9949 (N_9949,N_5253,N_5951);
nand U9950 (N_9950,N_6724,N_6051);
nor U9951 (N_9951,N_7208,N_6287);
or U9952 (N_9952,N_5594,N_7237);
nor U9953 (N_9953,N_7404,N_6901);
and U9954 (N_9954,N_6820,N_7169);
nand U9955 (N_9955,N_6890,N_5131);
nand U9956 (N_9956,N_5137,N_6642);
or U9957 (N_9957,N_6806,N_6296);
and U9958 (N_9958,N_6030,N_6887);
and U9959 (N_9959,N_5970,N_7186);
or U9960 (N_9960,N_5862,N_6368);
nand U9961 (N_9961,N_5851,N_6116);
nor U9962 (N_9962,N_6160,N_6158);
nand U9963 (N_9963,N_6796,N_7035);
nand U9964 (N_9964,N_5149,N_5650);
nand U9965 (N_9965,N_5100,N_7091);
nor U9966 (N_9966,N_6279,N_6128);
nor U9967 (N_9967,N_7095,N_6468);
nand U9968 (N_9968,N_6586,N_5661);
and U9969 (N_9969,N_7484,N_6787);
and U9970 (N_9970,N_6038,N_6581);
and U9971 (N_9971,N_7170,N_6147);
and U9972 (N_9972,N_7199,N_6894);
nor U9973 (N_9973,N_7010,N_6153);
nor U9974 (N_9974,N_5969,N_5596);
nor U9975 (N_9975,N_6065,N_6786);
nand U9976 (N_9976,N_6708,N_5891);
nor U9977 (N_9977,N_7253,N_7037);
nor U9978 (N_9978,N_6216,N_6666);
nand U9979 (N_9979,N_5557,N_7114);
nand U9980 (N_9980,N_6462,N_6111);
nor U9981 (N_9981,N_5419,N_6695);
nor U9982 (N_9982,N_5561,N_5377);
or U9983 (N_9983,N_5145,N_7150);
and U9984 (N_9984,N_6573,N_6187);
nor U9985 (N_9985,N_5092,N_5382);
and U9986 (N_9986,N_7324,N_5592);
or U9987 (N_9987,N_6097,N_5245);
or U9988 (N_9988,N_5734,N_5779);
xnor U9989 (N_9989,N_7106,N_5019);
or U9990 (N_9990,N_5523,N_6675);
and U9991 (N_9991,N_7293,N_5569);
nand U9992 (N_9992,N_6661,N_7142);
nand U9993 (N_9993,N_6224,N_7281);
nor U9994 (N_9994,N_6903,N_6387);
nand U9995 (N_9995,N_6319,N_5690);
nand U9996 (N_9996,N_7489,N_7316);
nor U9997 (N_9997,N_5606,N_6288);
nand U9998 (N_9998,N_7087,N_6748);
and U9999 (N_9999,N_6085,N_5528);
and UO_0 (O_0,N_7815,N_9553);
nor UO_1 (O_1,N_9048,N_7547);
and UO_2 (O_2,N_7534,N_9689);
or UO_3 (O_3,N_9247,N_7566);
nand UO_4 (O_4,N_9976,N_9390);
nand UO_5 (O_5,N_7631,N_7753);
and UO_6 (O_6,N_7918,N_8359);
nand UO_7 (O_7,N_9192,N_8910);
and UO_8 (O_8,N_7654,N_8968);
nand UO_9 (O_9,N_8828,N_9913);
nor UO_10 (O_10,N_7934,N_9906);
and UO_11 (O_11,N_9452,N_8844);
xnor UO_12 (O_12,N_8084,N_9824);
nor UO_13 (O_13,N_9130,N_8100);
nand UO_14 (O_14,N_8031,N_8788);
and UO_15 (O_15,N_8219,N_8108);
nand UO_16 (O_16,N_8687,N_9015);
nor UO_17 (O_17,N_7866,N_8428);
nor UO_18 (O_18,N_8866,N_7682);
nor UO_19 (O_19,N_8778,N_7587);
nand UO_20 (O_20,N_7892,N_8837);
or UO_21 (O_21,N_8401,N_9091);
nor UO_22 (O_22,N_9672,N_8038);
nor UO_23 (O_23,N_8296,N_7962);
and UO_24 (O_24,N_9308,N_8545);
or UO_25 (O_25,N_8379,N_7997);
or UO_26 (O_26,N_9950,N_7855);
nor UO_27 (O_27,N_9534,N_7707);
and UO_28 (O_28,N_9682,N_7709);
or UO_29 (O_29,N_8135,N_7567);
nand UO_30 (O_30,N_8931,N_9529);
nor UO_31 (O_31,N_8602,N_7910);
or UO_32 (O_32,N_8249,N_8824);
nand UO_33 (O_33,N_7693,N_9416);
and UO_34 (O_34,N_8344,N_9379);
nand UO_35 (O_35,N_7665,N_7965);
or UO_36 (O_36,N_7782,N_8624);
nand UO_37 (O_37,N_8611,N_7519);
or UO_38 (O_38,N_9227,N_7717);
nand UO_39 (O_39,N_8833,N_8520);
nor UO_40 (O_40,N_8391,N_9267);
and UO_41 (O_41,N_8935,N_8403);
or UO_42 (O_42,N_7677,N_9571);
or UO_43 (O_43,N_9386,N_8934);
and UO_44 (O_44,N_8407,N_9068);
or UO_45 (O_45,N_8338,N_8321);
or UO_46 (O_46,N_7669,N_9823);
nor UO_47 (O_47,N_7915,N_7554);
nor UO_48 (O_48,N_9144,N_8144);
nand UO_49 (O_49,N_9791,N_8838);
or UO_50 (O_50,N_8067,N_8522);
and UO_51 (O_51,N_9463,N_8559);
or UO_52 (O_52,N_8238,N_7950);
and UO_53 (O_53,N_9219,N_7886);
nor UO_54 (O_54,N_9148,N_8974);
nor UO_55 (O_55,N_8993,N_9923);
and UO_56 (O_56,N_9900,N_8761);
nor UO_57 (O_57,N_9589,N_8836);
and UO_58 (O_58,N_9440,N_8277);
nand UO_59 (O_59,N_7739,N_9607);
nor UO_60 (O_60,N_7546,N_9320);
nand UO_61 (O_61,N_8731,N_9277);
nand UO_62 (O_62,N_7616,N_8871);
nor UO_63 (O_63,N_9132,N_8620);
and UO_64 (O_64,N_9590,N_8521);
nor UO_65 (O_65,N_9852,N_7964);
nand UO_66 (O_66,N_8926,N_7958);
and UO_67 (O_67,N_9761,N_9565);
nor UO_68 (O_68,N_9433,N_8257);
or UO_69 (O_69,N_9645,N_7561);
or UO_70 (O_70,N_8656,N_7775);
nand UO_71 (O_71,N_9347,N_9254);
and UO_72 (O_72,N_8068,N_9343);
nand UO_73 (O_73,N_9289,N_9972);
nand UO_74 (O_74,N_9635,N_8515);
or UO_75 (O_75,N_8167,N_9202);
and UO_76 (O_76,N_8215,N_8625);
and UO_77 (O_77,N_9973,N_7689);
and UO_78 (O_78,N_7553,N_9818);
or UO_79 (O_79,N_8904,N_9969);
nor UO_80 (O_80,N_9723,N_8468);
and UO_81 (O_81,N_8117,N_9399);
and UO_82 (O_82,N_8216,N_9451);
and UO_83 (O_83,N_8438,N_8819);
nor UO_84 (O_84,N_7933,N_8063);
and UO_85 (O_85,N_9889,N_9070);
nor UO_86 (O_86,N_8448,N_7759);
and UO_87 (O_87,N_8912,N_8231);
nand UO_88 (O_88,N_8193,N_8430);
nor UO_89 (O_89,N_9807,N_8358);
and UO_90 (O_90,N_9816,N_8382);
or UO_91 (O_91,N_9592,N_8812);
nand UO_92 (O_92,N_9510,N_9485);
nand UO_93 (O_93,N_7778,N_7568);
nand UO_94 (O_94,N_7835,N_8504);
nor UO_95 (O_95,N_8503,N_7727);
nand UO_96 (O_96,N_9705,N_9221);
nand UO_97 (O_97,N_9581,N_9491);
xor UO_98 (O_98,N_9321,N_7879);
nand UO_99 (O_99,N_9316,N_9276);
nor UO_100 (O_100,N_7639,N_9191);
nand UO_101 (O_101,N_7578,N_9947);
and UO_102 (O_102,N_9615,N_8032);
and UO_103 (O_103,N_9515,N_8875);
or UO_104 (O_104,N_9763,N_8714);
nand UO_105 (O_105,N_8133,N_8311);
nand UO_106 (O_106,N_9415,N_7819);
and UO_107 (O_107,N_7992,N_9545);
nand UO_108 (O_108,N_8138,N_7668);
and UO_109 (O_109,N_7943,N_9785);
or UO_110 (O_110,N_7684,N_9292);
or UO_111 (O_111,N_7975,N_8813);
nor UO_112 (O_112,N_8886,N_8134);
nand UO_113 (O_113,N_9237,N_7876);
or UO_114 (O_114,N_7661,N_8678);
and UO_115 (O_115,N_7741,N_8347);
nand UO_116 (O_116,N_9480,N_9108);
nor UO_117 (O_117,N_9026,N_8066);
nand UO_118 (O_118,N_7862,N_8431);
nor UO_119 (O_119,N_9685,N_9876);
and UO_120 (O_120,N_9446,N_7941);
xnor UO_121 (O_121,N_9676,N_8738);
nor UO_122 (O_122,N_8684,N_9625);
nand UO_123 (O_123,N_8380,N_8488);
nor UO_124 (O_124,N_9476,N_9945);
nand UO_125 (O_125,N_7514,N_8073);
or UO_126 (O_126,N_7725,N_8682);
xor UO_127 (O_127,N_9483,N_9044);
or UO_128 (O_128,N_9944,N_8252);
or UO_129 (O_129,N_7990,N_8486);
nor UO_130 (O_130,N_7538,N_8023);
nand UO_131 (O_131,N_8809,N_8927);
or UO_132 (O_132,N_9284,N_9879);
or UO_133 (O_133,N_8242,N_8500);
or UO_134 (O_134,N_7909,N_7613);
and UO_135 (O_135,N_9102,N_7721);
and UO_136 (O_136,N_9001,N_9624);
and UO_137 (O_137,N_8473,N_8298);
nor UO_138 (O_138,N_9904,N_8071);
nor UO_139 (O_139,N_7884,N_9438);
nand UO_140 (O_140,N_8537,N_8642);
nor UO_141 (O_141,N_9080,N_9633);
nor UO_142 (O_142,N_9739,N_8578);
and UO_143 (O_143,N_8665,N_9586);
and UO_144 (O_144,N_8889,N_7555);
nor UO_145 (O_145,N_9055,N_9787);
or UO_146 (O_146,N_8777,N_9429);
nor UO_147 (O_147,N_8955,N_7598);
nand UO_148 (O_148,N_9754,N_9346);
nor UO_149 (O_149,N_8436,N_9306);
or UO_150 (O_150,N_9640,N_8739);
nand UO_151 (O_151,N_9465,N_8948);
nor UO_152 (O_152,N_9554,N_9541);
nor UO_153 (O_153,N_8973,N_8363);
nor UO_154 (O_154,N_9502,N_9424);
nand UO_155 (O_155,N_8169,N_8530);
nand UO_156 (O_156,N_8888,N_8165);
nand UO_157 (O_157,N_8322,N_8876);
and UO_158 (O_158,N_9018,N_8471);
or UO_159 (O_159,N_8939,N_8571);
or UO_160 (O_160,N_8799,N_8137);
and UO_161 (O_161,N_8709,N_7698);
nand UO_162 (O_162,N_9870,N_7860);
nor UO_163 (O_163,N_9792,N_8972);
nor UO_164 (O_164,N_7812,N_9370);
xnor UO_165 (O_165,N_9097,N_7895);
and UO_166 (O_166,N_7762,N_9223);
and UO_167 (O_167,N_7742,N_7694);
xnor UO_168 (O_168,N_9993,N_8657);
nor UO_169 (O_169,N_8007,N_8465);
nor UO_170 (O_170,N_8342,N_9008);
or UO_171 (O_171,N_8364,N_9563);
nand UO_172 (O_172,N_8154,N_7969);
and UO_173 (O_173,N_8750,N_9938);
or UO_174 (O_174,N_7829,N_8418);
nand UO_175 (O_175,N_8177,N_7672);
nand UO_176 (O_176,N_9076,N_8985);
and UO_177 (O_177,N_9500,N_9421);
nor UO_178 (O_178,N_7731,N_8148);
or UO_179 (O_179,N_9899,N_9608);
and UO_180 (O_180,N_9060,N_8132);
and UO_181 (O_181,N_8557,N_8028);
nand UO_182 (O_182,N_9569,N_9318);
xnor UO_183 (O_183,N_9867,N_8880);
nor UO_184 (O_184,N_9720,N_9989);
and UO_185 (O_185,N_8383,N_7550);
or UO_186 (O_186,N_8692,N_9755);
nand UO_187 (O_187,N_7501,N_8070);
nand UO_188 (O_188,N_9744,N_9382);
or UO_189 (O_189,N_9146,N_7632);
nand UO_190 (O_190,N_8782,N_9279);
nor UO_191 (O_191,N_9332,N_7692);
and UO_192 (O_192,N_8282,N_9765);
nand UO_193 (O_193,N_7838,N_8923);
nor UO_194 (O_194,N_9393,N_8513);
and UO_195 (O_195,N_8373,N_8981);
nand UO_196 (O_196,N_9134,N_9925);
nand UO_197 (O_197,N_8109,N_9437);
nor UO_198 (O_198,N_8632,N_8289);
nand UO_199 (O_199,N_8958,N_8015);
nor UO_200 (O_200,N_8287,N_7715);
nand UO_201 (O_201,N_8233,N_8176);
or UO_202 (O_202,N_9599,N_8872);
and UO_203 (O_203,N_8369,N_9647);
or UO_204 (O_204,N_9381,N_8111);
nor UO_205 (O_205,N_8098,N_9956);
nor UO_206 (O_206,N_9936,N_7617);
nand UO_207 (O_207,N_9525,N_7521);
nor UO_208 (O_208,N_7635,N_9391);
or UO_209 (O_209,N_8439,N_8114);
or UO_210 (O_210,N_8721,N_8095);
or UO_211 (O_211,N_8495,N_8827);
or UO_212 (O_212,N_8320,N_9588);
nand UO_213 (O_213,N_8519,N_9403);
or UO_214 (O_214,N_9780,N_7618);
or UO_215 (O_215,N_8285,N_8779);
nand UO_216 (O_216,N_9269,N_8618);
nand UO_217 (O_217,N_8808,N_8390);
or UO_218 (O_218,N_7542,N_9115);
nand UO_219 (O_219,N_9136,N_8190);
nand UO_220 (O_220,N_7947,N_7510);
nor UO_221 (O_221,N_8327,N_8697);
nand UO_222 (O_222,N_8646,N_8386);
and UO_223 (O_223,N_9957,N_8938);
nor UO_224 (O_224,N_9698,N_8220);
and UO_225 (O_225,N_8004,N_9329);
xor UO_226 (O_226,N_9622,N_8393);
nand UO_227 (O_227,N_9105,N_9657);
nand UO_228 (O_228,N_9241,N_8535);
and UO_229 (O_229,N_9345,N_7652);
or UO_230 (O_230,N_8275,N_8708);
nand UO_231 (O_231,N_8843,N_7908);
and UO_232 (O_232,N_7904,N_9492);
or UO_233 (O_233,N_8966,N_7802);
xnor UO_234 (O_234,N_9441,N_9022);
or UO_235 (O_235,N_8039,N_8204);
nand UO_236 (O_236,N_8397,N_9988);
nor UO_237 (O_237,N_7795,N_8278);
nor UO_238 (O_238,N_9605,N_7755);
nor UO_239 (O_239,N_9783,N_8641);
nor UO_240 (O_240,N_7922,N_9600);
and UO_241 (O_241,N_7912,N_8351);
nand UO_242 (O_242,N_9142,N_7560);
or UO_243 (O_243,N_8326,N_7705);
or UO_244 (O_244,N_8997,N_8588);
nor UO_245 (O_245,N_9039,N_9653);
nand UO_246 (O_246,N_8952,N_9328);
and UO_247 (O_247,N_7607,N_7834);
and UO_248 (O_248,N_8835,N_7869);
and UO_249 (O_249,N_8821,N_8756);
or UO_250 (O_250,N_8541,N_8614);
nand UO_251 (O_251,N_9781,N_8659);
or UO_252 (O_252,N_8423,N_9776);
nand UO_253 (O_253,N_8470,N_9695);
xnor UO_254 (O_254,N_8865,N_9866);
nand UO_255 (O_255,N_9921,N_8677);
nor UO_256 (O_256,N_9287,N_7936);
and UO_257 (O_257,N_9533,N_8770);
nor UO_258 (O_258,N_8884,N_9639);
or UO_259 (O_259,N_9208,N_9914);
nand UO_260 (O_260,N_9642,N_9244);
nand UO_261 (O_261,N_9021,N_7940);
nand UO_262 (O_262,N_8329,N_8699);
nor UO_263 (O_263,N_8259,N_9771);
nor UO_264 (O_264,N_8455,N_9283);
nand UO_265 (O_265,N_8149,N_9859);
nor UO_266 (O_266,N_8728,N_8054);
and UO_267 (O_267,N_9798,N_8774);
and UO_268 (O_268,N_9729,N_9644);
nand UO_269 (O_269,N_8505,N_8052);
nand UO_270 (O_270,N_8601,N_9074);
or UO_271 (O_271,N_9479,N_7558);
or UO_272 (O_272,N_9195,N_9087);
nand UO_273 (O_273,N_9082,N_8967);
nand UO_274 (O_274,N_8356,N_8897);
nor UO_275 (O_275,N_9246,N_8551);
nand UO_276 (O_276,N_9171,N_9450);
nand UO_277 (O_277,N_8956,N_9718);
or UO_278 (O_278,N_8088,N_8789);
nor UO_279 (O_279,N_9675,N_9673);
and UO_280 (O_280,N_8664,N_7877);
nand UO_281 (O_281,N_7513,N_7574);
nand UO_282 (O_282,N_8826,N_8166);
and UO_283 (O_283,N_8309,N_8757);
or UO_284 (O_284,N_8268,N_8343);
xnor UO_285 (O_285,N_8553,N_8544);
or UO_286 (O_286,N_8203,N_9160);
nor UO_287 (O_287,N_8569,N_7619);
xor UO_288 (O_288,N_9960,N_8570);
and UO_289 (O_289,N_7900,N_9941);
and UO_290 (O_290,N_9669,N_9730);
or UO_291 (O_291,N_7529,N_9487);
nand UO_292 (O_292,N_9325,N_9954);
nand UO_293 (O_293,N_8698,N_7552);
nand UO_294 (O_294,N_9875,N_8053);
and UO_295 (O_295,N_8690,N_8723);
nand UO_296 (O_296,N_9951,N_9499);
and UO_297 (O_297,N_8832,N_9539);
nand UO_298 (O_298,N_8766,N_8603);
nor UO_299 (O_299,N_7984,N_9775);
and UO_300 (O_300,N_8457,N_9892);
nor UO_301 (O_301,N_9069,N_8254);
and UO_302 (O_302,N_7718,N_8726);
or UO_303 (O_303,N_9072,N_8538);
and UO_304 (O_304,N_8310,N_8388);
and UO_305 (O_305,N_9704,N_8925);
nand UO_306 (O_306,N_9457,N_9456);
or UO_307 (O_307,N_9182,N_7946);
or UO_308 (O_308,N_8396,N_9516);
nand UO_309 (O_309,N_7564,N_9757);
and UO_310 (O_310,N_7599,N_9377);
or UO_311 (O_311,N_8971,N_9715);
or UO_312 (O_312,N_8302,N_8691);
and UO_313 (O_313,N_7535,N_8555);
nand UO_314 (O_314,N_8283,N_7852);
or UO_315 (O_315,N_7585,N_8000);
nand UO_316 (O_316,N_9414,N_7633);
or UO_317 (O_317,N_8858,N_8615);
nor UO_318 (O_318,N_8499,N_8501);
or UO_319 (O_319,N_9686,N_9627);
nand UO_320 (O_320,N_7889,N_9595);
nand UO_321 (O_321,N_9507,N_8159);
and UO_322 (O_322,N_7559,N_9305);
nand UO_323 (O_323,N_8341,N_8492);
and UO_324 (O_324,N_9861,N_8335);
and UO_325 (O_325,N_8550,N_9408);
and UO_326 (O_326,N_7624,N_8306);
or UO_327 (O_327,N_8528,N_7512);
and UO_328 (O_328,N_9760,N_7743);
and UO_329 (O_329,N_7994,N_7893);
nor UO_330 (O_330,N_8706,N_7730);
or UO_331 (O_331,N_9339,N_7752);
or UO_332 (O_332,N_8208,N_7785);
or UO_333 (O_333,N_9344,N_7590);
nand UO_334 (O_334,N_9317,N_8362);
nand UO_335 (O_335,N_8506,N_9240);
nor UO_336 (O_336,N_9203,N_8076);
nor UO_337 (O_337,N_9658,N_7985);
nor UO_338 (O_338,N_8724,N_9089);
nor UO_339 (O_339,N_9845,N_9767);
xnor UO_340 (O_340,N_8058,N_8354);
nor UO_341 (O_341,N_9943,N_9519);
and UO_342 (O_342,N_9931,N_9178);
and UO_343 (O_343,N_9295,N_9290);
nor UO_344 (O_344,N_7620,N_8531);
and UO_345 (O_345,N_9612,N_9410);
and UO_346 (O_346,N_9618,N_8083);
nand UO_347 (O_347,N_7569,N_7953);
and UO_348 (O_348,N_9811,N_8147);
and UO_349 (O_349,N_9555,N_8387);
nand UO_350 (O_350,N_9575,N_9073);
or UO_351 (O_351,N_9229,N_9017);
nor UO_352 (O_352,N_8152,N_7971);
nor UO_353 (O_353,N_7858,N_8795);
or UO_354 (O_354,N_9352,N_8930);
and UO_355 (O_355,N_8890,N_7540);
or UO_356 (O_356,N_7736,N_8599);
and UO_357 (O_357,N_7606,N_8785);
or UO_358 (O_358,N_8218,N_9323);
nand UO_359 (O_359,N_8466,N_9453);
nand UO_360 (O_360,N_8862,N_8790);
xor UO_361 (O_361,N_9131,N_8304);
nor UO_362 (O_362,N_8037,N_9409);
or UO_363 (O_363,N_9426,N_9122);
and UO_364 (O_364,N_9610,N_8755);
nand UO_365 (O_365,N_9315,N_8561);
or UO_366 (O_366,N_9172,N_8185);
nand UO_367 (O_367,N_7744,N_9827);
nor UO_368 (O_368,N_7629,N_9817);
nor UO_369 (O_369,N_8671,N_7854);
nor UO_370 (O_370,N_8994,N_9447);
or UO_371 (O_371,N_7848,N_8527);
or UO_372 (O_372,N_7779,N_9762);
or UO_373 (O_373,N_8173,N_7924);
nor UO_374 (O_374,N_7956,N_7667);
or UO_375 (O_375,N_9062,N_9650);
xnor UO_376 (O_376,N_8735,N_7926);
nor UO_377 (O_377,N_9562,N_8831);
nor UO_378 (O_378,N_7737,N_8469);
nor UO_379 (O_379,N_9789,N_9366);
or UO_380 (O_380,N_9979,N_8801);
nor UO_381 (O_381,N_8653,N_8201);
or UO_382 (O_382,N_9819,N_9474);
and UO_383 (O_383,N_7515,N_9140);
nor UO_384 (O_384,N_9919,N_8496);
nand UO_385 (O_385,N_9175,N_7660);
or UO_386 (O_386,N_9559,N_8734);
and UO_387 (O_387,N_8686,N_9693);
nor UO_388 (O_388,N_8957,N_9064);
and UO_389 (O_389,N_9226,N_7604);
nand UO_390 (O_390,N_9768,N_7967);
nor UO_391 (O_391,N_9367,N_9877);
or UO_392 (O_392,N_9782,N_8035);
and UO_393 (O_393,N_9000,N_8020);
nor UO_394 (O_394,N_9712,N_7708);
or UO_395 (O_395,N_9706,N_8415);
or UO_396 (O_396,N_7638,N_8491);
nor UO_397 (O_397,N_7865,N_7827);
or UO_398 (O_398,N_9006,N_8575);
nor UO_399 (O_399,N_8695,N_8759);
nor UO_400 (O_400,N_7563,N_9832);
and UO_401 (O_401,N_9207,N_9585);
nand UO_402 (O_402,N_8370,N_7735);
or UO_403 (O_403,N_8719,N_8552);
or UO_404 (O_404,N_9855,N_9138);
nor UO_405 (O_405,N_7983,N_8893);
nand UO_406 (O_406,N_8003,N_9436);
and UO_407 (O_407,N_8892,N_9112);
nor UO_408 (O_408,N_7581,N_9873);
nor UO_409 (O_409,N_9190,N_7919);
nor UO_410 (O_410,N_9319,N_7653);
or UO_411 (O_411,N_7565,N_9364);
and UO_412 (O_412,N_8284,N_7573);
nor UO_413 (O_413,N_8043,N_8451);
and UO_414 (O_414,N_8946,N_9858);
or UO_415 (O_415,N_9907,N_8034);
or UO_416 (O_416,N_9025,N_9733);
and UO_417 (O_417,N_9667,N_8959);
or UO_418 (O_418,N_8869,N_8404);
and UO_419 (O_419,N_8232,N_9197);
or UO_420 (O_420,N_7504,N_8280);
nand UO_421 (O_421,N_9666,N_9802);
or UO_422 (O_422,N_9854,N_7928);
or UO_423 (O_423,N_8518,N_9580);
nand UO_424 (O_424,N_9684,N_9978);
nor UO_425 (O_425,N_7863,N_9868);
nor UO_426 (O_426,N_9806,N_8881);
and UO_427 (O_427,N_9149,N_8919);
xnor UO_428 (O_428,N_9127,N_8806);
nand UO_429 (O_429,N_8752,N_8915);
and UO_430 (O_430,N_9093,N_8102);
or UO_431 (O_431,N_9997,N_9201);
and UO_432 (O_432,N_7982,N_8896);
nand UO_433 (O_433,N_9081,N_7734);
and UO_434 (O_434,N_8840,N_9309);
nor UO_435 (O_435,N_8211,N_7592);
nor UO_436 (O_436,N_9591,N_9561);
nand UO_437 (O_437,N_9905,N_7981);
and UO_438 (O_438,N_8701,N_9939);
nor UO_439 (O_439,N_8345,N_8863);
nor UO_440 (O_440,N_7676,N_9825);
nand UO_441 (O_441,N_9054,N_8798);
nor UO_442 (O_442,N_9946,N_9238);
nor UO_443 (O_443,N_8247,N_9623);
nor UO_444 (O_444,N_8630,N_8437);
nor UO_445 (O_445,N_8206,N_8803);
nor UO_446 (O_446,N_7516,N_7872);
and UO_447 (O_447,N_8199,N_9294);
or UO_448 (O_448,N_7822,N_8720);
nand UO_449 (O_449,N_8047,N_8125);
xnor UO_450 (O_450,N_7800,N_9641);
or UO_451 (O_451,N_9129,N_9137);
nor UO_452 (O_452,N_9310,N_9740);
nand UO_453 (O_453,N_8334,N_9758);
nor UO_454 (O_454,N_7626,N_8882);
and UO_455 (O_455,N_9020,N_7781);
nand UO_456 (O_456,N_9716,N_9694);
nand UO_457 (O_457,N_9128,N_8508);
or UO_458 (O_458,N_8784,N_9917);
and UO_459 (O_459,N_8086,N_8940);
or UO_460 (O_460,N_8027,N_9752);
nand UO_461 (O_461,N_8754,N_9596);
or UO_462 (O_462,N_8445,N_8652);
and UO_463 (O_463,N_9168,N_7976);
nor UO_464 (O_464,N_8597,N_9119);
nand UO_465 (O_465,N_8577,N_8791);
and UO_466 (O_466,N_7740,N_9540);
or UO_467 (O_467,N_9746,N_9493);
and UO_468 (O_468,N_7646,N_9828);
and UO_469 (O_469,N_8591,N_7843);
nor UO_470 (O_470,N_7760,N_9751);
nor UO_471 (O_471,N_9531,N_9880);
nand UO_472 (O_472,N_8787,N_9501);
nor UO_473 (O_473,N_7771,N_8440);
and UO_474 (O_474,N_8091,N_9745);
nand UO_475 (O_475,N_9503,N_9371);
and UO_476 (O_476,N_9257,N_8769);
and UO_477 (O_477,N_9342,N_7864);
xnor UO_478 (O_478,N_9930,N_9312);
nand UO_479 (O_479,N_9604,N_9544);
and UO_480 (O_480,N_8852,N_7963);
or UO_481 (O_481,N_7615,N_7506);
and UO_482 (O_482,N_9412,N_9714);
or UO_483 (O_483,N_7820,N_7808);
or UO_484 (O_484,N_8617,N_8730);
and UO_485 (O_485,N_8619,N_8540);
or UO_486 (O_486,N_8346,N_9674);
and UO_487 (O_487,N_8303,N_8853);
or UO_488 (O_488,N_8891,N_8947);
or UO_489 (O_489,N_9546,N_8222);
nor UO_490 (O_490,N_8096,N_9103);
nand UO_491 (O_491,N_7888,N_9075);
or UO_492 (O_492,N_7695,N_9630);
or UO_493 (O_493,N_8977,N_9826);
or UO_494 (O_494,N_9844,N_9583);
or UO_495 (O_495,N_7833,N_9123);
or UO_496 (O_496,N_8517,N_8205);
or UO_497 (O_497,N_9111,N_9187);
nor UO_498 (O_498,N_8765,N_8319);
xnor UO_499 (O_499,N_8894,N_8658);
or UO_500 (O_500,N_9461,N_9847);
nand UO_501 (O_501,N_7657,N_8818);
and UO_502 (O_502,N_8604,N_8026);
nand UO_503 (O_503,N_8796,N_8902);
nand UO_504 (O_504,N_8494,N_8006);
or UO_505 (O_505,N_9511,N_9722);
nand UO_506 (O_506,N_9286,N_8516);
nand UO_507 (O_507,N_7749,N_8410);
nor UO_508 (O_508,N_7772,N_8606);
nand UO_509 (O_509,N_9488,N_9737);
nor UO_510 (O_510,N_7898,N_8075);
or UO_511 (O_511,N_9968,N_7720);
or UO_512 (O_512,N_9373,N_9609);
and UO_513 (O_513,N_9690,N_8859);
nor UO_514 (O_514,N_7644,N_7859);
and UO_515 (O_515,N_8136,N_9679);
nand UO_516 (O_516,N_8458,N_8776);
and UO_517 (O_517,N_8005,N_7696);
or UO_518 (O_518,N_9952,N_7656);
nor UO_519 (O_519,N_7831,N_8197);
or UO_520 (O_520,N_9882,N_9402);
nand UO_521 (O_521,N_7750,N_8049);
and UO_522 (O_522,N_8547,N_9724);
nand UO_523 (O_523,N_8638,N_9301);
and UO_524 (O_524,N_9885,N_9363);
or UO_525 (O_525,N_7973,N_8978);
or UO_526 (O_526,N_8767,N_9209);
nor UO_527 (O_527,N_8683,N_8429);
and UO_528 (O_528,N_8583,N_9983);
and UO_529 (O_529,N_8292,N_9547);
and UO_530 (O_530,N_9849,N_8643);
and UO_531 (O_531,N_9655,N_9831);
nor UO_532 (O_532,N_8610,N_8224);
xnor UO_533 (O_533,N_8113,N_9863);
nor UO_534 (O_534,N_8480,N_7610);
nor UO_535 (O_535,N_8463,N_8811);
or UO_536 (O_536,N_8402,N_8945);
nand UO_537 (O_537,N_8077,N_8124);
and UO_538 (O_538,N_9029,N_8061);
nand UO_539 (O_539,N_7745,N_9296);
or UO_540 (O_540,N_9125,N_8584);
or UO_541 (O_541,N_8929,N_8253);
nor UO_542 (O_542,N_7957,N_9005);
and UO_543 (O_543,N_8348,N_8669);
nor UO_544 (O_544,N_9235,N_9794);
nand UO_545 (O_545,N_9728,N_7770);
nor UO_546 (O_546,N_8580,N_9556);
nand UO_547 (O_547,N_8751,N_8857);
nor UO_548 (O_548,N_8667,N_8421);
nor UO_549 (O_549,N_9738,N_9860);
and UO_550 (O_550,N_8195,N_9526);
nor UO_551 (O_551,N_7509,N_8702);
nand UO_552 (O_552,N_8368,N_8793);
nand UO_553 (O_553,N_9193,N_9508);
nor UO_554 (O_554,N_7518,N_9949);
and UO_555 (O_555,N_9948,N_8366);
xor UO_556 (O_556,N_8822,N_7951);
or UO_557 (O_557,N_9986,N_7883);
nand UO_558 (O_558,N_8953,N_9932);
or UO_559 (O_559,N_8024,N_9883);
nor UO_560 (O_560,N_9243,N_9004);
or UO_561 (O_561,N_9509,N_9220);
nor UO_562 (O_562,N_9288,N_7623);
or UO_563 (O_563,N_8961,N_7837);
nand UO_564 (O_564,N_8250,N_8189);
nand UO_565 (O_565,N_8449,N_8243);
nand UO_566 (O_566,N_9846,N_8223);
or UO_567 (O_567,N_9560,N_9330);
nor UO_568 (O_568,N_7641,N_7557);
and UO_569 (O_569,N_9611,N_8841);
or UO_570 (O_570,N_8244,N_9053);
nand UO_571 (O_571,N_8514,N_8014);
nand UO_572 (O_572,N_7505,N_8693);
nand UO_573 (O_573,N_9632,N_9601);
and UO_574 (O_574,N_9378,N_8163);
xnor UO_575 (O_575,N_7671,N_8922);
and UO_576 (O_576,N_8021,N_7856);
and UO_577 (O_577,N_9272,N_8874);
nor UO_578 (O_578,N_8747,N_7916);
or UO_579 (O_579,N_8093,N_8607);
or UO_580 (O_580,N_9460,N_7816);
and UO_581 (O_581,N_9985,N_7897);
nand UO_582 (O_582,N_9638,N_9028);
nor UO_583 (O_583,N_9574,N_7847);
and UO_584 (O_584,N_8908,N_8887);
and UO_585 (O_585,N_9159,N_7970);
nor UO_586 (O_586,N_9059,N_9239);
nand UO_587 (O_587,N_7729,N_8814);
or UO_588 (O_588,N_8427,N_7938);
and UO_589 (O_589,N_8804,N_8210);
nand UO_590 (O_590,N_9063,N_9649);
or UO_591 (O_591,N_8685,N_7959);
xnor UO_592 (O_592,N_7579,N_9741);
nor UO_593 (O_593,N_9908,N_8291);
nor UO_594 (O_594,N_9928,N_8936);
nor UO_595 (O_595,N_9784,N_9701);
nand UO_596 (O_596,N_7930,N_8119);
and UO_597 (O_597,N_9886,N_7783);
nor UO_598 (O_598,N_9537,N_9663);
and UO_599 (O_599,N_9566,N_7679);
or UO_600 (O_600,N_8414,N_9088);
or UO_601 (O_601,N_7666,N_8675);
and UO_602 (O_602,N_9430,N_9890);
or UO_603 (O_603,N_8975,N_9009);
nor UO_604 (O_604,N_9336,N_9445);
or UO_605 (O_605,N_7927,N_9955);
or UO_606 (O_606,N_9839,N_8318);
and UO_607 (O_607,N_7972,N_8526);
or UO_608 (O_608,N_9814,N_7507);
nor UO_609 (O_609,N_8235,N_7921);
and UO_610 (O_610,N_9994,N_9518);
nand UO_611 (O_611,N_8523,N_8140);
or UO_612 (O_612,N_9333,N_9079);
and UO_613 (O_613,N_8905,N_8155);
nor UO_614 (O_614,N_9620,N_9918);
nand UO_615 (O_615,N_7543,N_8272);
nand UO_616 (O_616,N_9857,N_8246);
or UO_617 (O_617,N_9356,N_9582);
nor UO_618 (O_618,N_9587,N_7597);
nand UO_619 (O_619,N_8564,N_9096);
or UO_620 (O_620,N_8405,N_9769);
and UO_621 (O_621,N_9404,N_9405);
or UO_622 (O_622,N_7608,N_8707);
nor UO_623 (O_623,N_8502,N_8025);
nand UO_624 (O_624,N_8670,N_8786);
nor UO_625 (O_625,N_7955,N_9872);
nand UO_626 (O_626,N_9522,N_7747);
or UO_627 (O_627,N_8573,N_9341);
nand UO_628 (O_628,N_9189,N_7524);
nor UO_629 (O_629,N_7769,N_8949);
xnor UO_630 (O_630,N_9617,N_7825);
nor UO_631 (O_631,N_9098,N_8099);
and UO_632 (O_632,N_7651,N_8995);
nand UO_633 (O_633,N_8988,N_8433);
or UO_634 (O_634,N_8758,N_8481);
nor UO_635 (O_635,N_9046,N_8141);
or UO_636 (O_636,N_8637,N_8256);
and UO_637 (O_637,N_8248,N_7589);
nand UO_638 (O_638,N_8122,N_9965);
nand UO_639 (O_639,N_9013,N_7814);
xnor UO_640 (O_640,N_8991,N_9958);
and UO_641 (O_641,N_8273,N_9183);
or UO_642 (O_642,N_7896,N_9637);
nand UO_643 (O_643,N_9250,N_7522);
nor UO_644 (O_644,N_8416,N_7591);
nor UO_645 (O_645,N_7583,N_8183);
xor UO_646 (O_646,N_9735,N_8308);
nor UO_647 (O_647,N_8411,N_8399);
nand UO_648 (O_648,N_9032,N_8916);
nor UO_649 (O_649,N_9790,N_9796);
xnor UO_650 (O_650,N_8426,N_9770);
nor UO_651 (O_651,N_8225,N_8593);
nand UO_652 (O_652,N_8834,N_8258);
or UO_653 (O_653,N_9871,N_9162);
nand UO_654 (O_654,N_8001,N_9278);
and UO_655 (O_655,N_8613,N_7821);
and UO_656 (O_656,N_8775,N_8434);
or UO_657 (O_657,N_9594,N_9517);
nor UO_658 (O_658,N_8172,N_8331);
nand UO_659 (O_659,N_9897,N_7685);
or UO_660 (O_660,N_8542,N_7776);
nand UO_661 (O_661,N_8846,N_8660);
xor UO_662 (O_662,N_8116,N_8554);
nor UO_663 (O_663,N_9466,N_7764);
nor UO_664 (O_664,N_7645,N_8768);
or UO_665 (O_665,N_8576,N_8666);
nor UO_666 (O_666,N_8885,N_8647);
or UO_667 (O_667,N_8030,N_8009);
or UO_668 (O_668,N_9113,N_9477);
nor UO_669 (O_669,N_9448,N_9893);
nand UO_670 (O_670,N_8145,N_8059);
nor UO_671 (O_671,N_8293,N_7508);
nor UO_672 (O_672,N_9829,N_8560);
nor UO_673 (O_673,N_9217,N_8187);
or UO_674 (O_674,N_8164,N_8533);
and UO_675 (O_675,N_7716,N_8568);
and UO_676 (O_676,N_8251,N_9734);
xor UO_677 (O_677,N_8482,N_8816);
and UO_678 (O_678,N_9671,N_9200);
and UO_679 (O_679,N_9139,N_7576);
or UO_680 (O_680,N_8703,N_9271);
nor UO_681 (O_681,N_9083,N_9158);
nor UO_682 (O_682,N_8230,N_7949);
and UO_683 (O_683,N_8722,N_8631);
nand UO_684 (O_684,N_9270,N_8467);
nor UO_685 (O_685,N_8781,N_9214);
and UO_686 (O_686,N_9703,N_8241);
and UO_687 (O_687,N_8679,N_9753);
or UO_688 (O_688,N_8040,N_9169);
nand UO_689 (O_689,N_9420,N_9143);
nand UO_690 (O_690,N_9764,N_7780);
xor UO_691 (O_691,N_7818,N_7944);
nor UO_692 (O_692,N_7625,N_8207);
or UO_693 (O_693,N_8089,N_9114);
nor UO_694 (O_694,N_9224,N_8989);
or UO_695 (O_695,N_9413,N_7528);
nand UO_696 (O_696,N_8493,N_8965);
or UO_697 (O_697,N_7659,N_8115);
nand UO_698 (O_698,N_8944,N_7784);
nor UO_699 (O_699,N_7987,N_7531);
nor UO_700 (O_700,N_9542,N_7798);
or UO_701 (O_701,N_9179,N_7768);
and UO_702 (O_702,N_8228,N_9273);
nor UO_703 (O_703,N_7712,N_8727);
nor UO_704 (O_704,N_8825,N_9443);
and UO_705 (O_705,N_7562,N_9660);
nor UO_706 (O_706,N_9687,N_9304);
and UO_707 (O_707,N_8128,N_8174);
or UO_708 (O_708,N_7907,N_7977);
nor UO_709 (O_709,N_8131,N_9840);
and UO_710 (O_710,N_9929,N_8074);
nand UO_711 (O_711,N_9702,N_8532);
nor UO_712 (O_712,N_8548,N_8688);
or UO_713 (O_713,N_8384,N_8700);
nor UO_714 (O_714,N_8425,N_7887);
xnor UO_715 (O_715,N_9992,N_8198);
nand UO_716 (O_716,N_7690,N_8674);
nand UO_717 (O_717,N_8810,N_9700);
or UO_718 (O_718,N_8717,N_8911);
nand UO_719 (O_719,N_7605,N_7611);
xor UO_720 (O_720,N_9634,N_8105);
and UO_721 (O_721,N_9253,N_9853);
nor UO_722 (O_722,N_8041,N_9154);
or UO_723 (O_723,N_7634,N_9249);
and UO_724 (O_724,N_9793,N_7711);
and UO_725 (O_725,N_7842,N_8337);
or UO_726 (O_726,N_9661,N_7714);
and UO_727 (O_727,N_8171,N_9362);
nand UO_728 (O_728,N_9494,N_9035);
or UO_729 (O_729,N_9709,N_8763);
nand UO_730 (O_730,N_7761,N_8120);
nor UO_731 (O_731,N_8712,N_7797);
nor UO_732 (O_732,N_9444,N_7539);
and UO_733 (O_733,N_8483,N_8389);
nor UO_734 (O_734,N_8168,N_7960);
nand UO_735 (O_735,N_8680,N_9407);
or UO_736 (O_736,N_9800,N_9262);
nor UO_737 (O_737,N_8305,N_8639);
or UO_738 (O_738,N_8033,N_7621);
and UO_739 (O_739,N_9388,N_8651);
nor UO_740 (O_740,N_9198,N_8950);
nor UO_741 (O_741,N_9084,N_8710);
nor UO_742 (O_742,N_9355,N_9212);
or UO_743 (O_743,N_7850,N_8903);
nor UO_744 (O_744,N_8055,N_9052);
and UO_745 (O_745,N_9151,N_7500);
and UO_746 (O_746,N_7813,N_8543);
or UO_747 (O_747,N_8556,N_8336);
nor UO_748 (O_748,N_8312,N_8546);
nand UO_749 (O_749,N_8072,N_9888);
and UO_750 (O_750,N_8281,N_9303);
nor UO_751 (O_751,N_9335,N_8487);
or UO_752 (O_752,N_9225,N_7925);
or UO_753 (O_753,N_8013,N_8510);
or UO_754 (O_754,N_8022,N_9173);
and UO_755 (O_755,N_7637,N_7614);
nand UO_756 (O_756,N_9258,N_8987);
nand UO_757 (O_757,N_9268,N_8572);
and UO_758 (O_758,N_8976,N_9389);
and UO_759 (O_759,N_7758,N_7874);
nand UO_760 (O_760,N_9117,N_7756);
nand UO_761 (O_761,N_9822,N_8654);
or UO_762 (O_762,N_8797,N_9033);
nor UO_763 (O_763,N_7636,N_9161);
or UO_764 (O_764,N_8276,N_8462);
xor UO_765 (O_765,N_9155,N_8877);
nand UO_766 (O_766,N_7674,N_9498);
and UO_767 (O_767,N_9464,N_8549);
or UO_768 (O_768,N_9963,N_8012);
xor UO_769 (O_769,N_8017,N_8815);
nand UO_770 (O_770,N_9417,N_8191);
or UO_771 (O_771,N_8476,N_7999);
or UO_772 (O_772,N_9552,N_7995);
or UO_773 (O_773,N_9530,N_9431);
or UO_774 (O_774,N_9731,N_9281);
and UO_775 (O_775,N_9652,N_9468);
nand UO_776 (O_776,N_8855,N_8325);
nor UO_777 (O_777,N_8590,N_8984);
nor UO_778 (O_778,N_7868,N_9194);
nor UO_779 (O_779,N_8101,N_9656);
xor UO_780 (O_780,N_7939,N_8107);
nor UO_781 (O_781,N_9205,N_8640);
xnor UO_782 (O_782,N_8534,N_8139);
nand UO_783 (O_783,N_8743,N_8442);
nor UO_784 (O_784,N_7658,N_8450);
and UO_785 (O_785,N_9233,N_9895);
nand UO_786 (O_786,N_8044,N_9307);
nor UO_787 (O_787,N_9042,N_8265);
nor UO_788 (O_788,N_9878,N_7595);
or UO_789 (O_789,N_9167,N_8274);
or UO_790 (O_790,N_9265,N_8998);
or UO_791 (O_791,N_9396,N_7902);
nand UO_792 (O_792,N_8616,N_8928);
nand UO_793 (O_793,N_8980,N_9801);
nor UO_794 (O_794,N_9648,N_9245);
and UO_795 (O_795,N_9543,N_9280);
nor UO_796 (O_796,N_9206,N_9864);
or UO_797 (O_797,N_7681,N_8010);
and UO_798 (O_798,N_8933,N_9489);
and UO_799 (O_799,N_9467,N_8008);
nor UO_800 (O_800,N_8713,N_8696);
and UO_801 (O_801,N_9174,N_8097);
xor UO_802 (O_802,N_9916,N_9747);
or UO_803 (O_803,N_8002,N_9538);
nand UO_804 (O_804,N_9470,N_7792);
nand UO_805 (O_805,N_8314,N_9778);
nand UO_806 (O_806,N_8663,N_8477);
and UO_807 (O_807,N_8626,N_8498);
nand UO_808 (O_808,N_7878,N_9099);
and UO_809 (O_809,N_8829,N_9912);
and UO_810 (O_810,N_8447,N_9406);
or UO_811 (O_811,N_8629,N_8294);
nor UO_812 (O_812,N_9380,N_7688);
nor UO_813 (O_813,N_7732,N_8900);
nor UO_814 (O_814,N_8443,N_7582);
nand UO_815 (O_815,N_9505,N_9490);
or UO_816 (O_816,N_9692,N_9971);
nand UO_817 (O_817,N_9260,N_8512);
nand UO_818 (O_818,N_7584,N_8360);
xor UO_819 (O_819,N_7880,N_8269);
or UO_820 (O_820,N_9557,N_7523);
and UO_821 (O_821,N_9598,N_7777);
and UO_822 (O_822,N_9773,N_8954);
or UO_823 (O_823,N_9991,N_8036);
nand UO_824 (O_824,N_7844,N_9248);
nor UO_825 (O_825,N_7670,N_8392);
nor UO_826 (O_826,N_9442,N_7766);
nor UO_827 (O_827,N_9812,N_8802);
nand UO_828 (O_828,N_8842,N_8650);
or UO_829 (O_829,N_7913,N_8595);
or UO_830 (O_830,N_8018,N_9334);
and UO_831 (O_831,N_7687,N_8999);
nand UO_832 (O_832,N_8413,N_9810);
and UO_833 (O_833,N_7602,N_7805);
nor UO_834 (O_834,N_8170,N_9124);
nor UO_835 (O_835,N_9631,N_9815);
and UO_836 (O_836,N_7733,N_7588);
and UO_837 (O_837,N_8864,N_8130);
nor UO_838 (O_838,N_9293,N_7713);
nand UO_839 (O_839,N_9213,N_9432);
and UO_840 (O_840,N_7807,N_7849);
nand UO_841 (O_841,N_8920,N_7942);
or UO_842 (O_842,N_8762,N_9216);
xnor UO_843 (O_843,N_8422,N_9513);
and UO_844 (O_844,N_8484,N_8992);
nand UO_845 (O_845,N_8146,N_9707);
nand UO_846 (O_846,N_7799,N_8741);
nor UO_847 (O_847,N_8725,N_8589);
nand UO_848 (O_848,N_9743,N_9536);
nand UO_849 (O_849,N_7532,N_7748);
nor UO_850 (O_850,N_8563,N_9311);
or UO_851 (O_851,N_9177,N_8419);
or UO_852 (O_852,N_9999,N_8472);
or UO_853 (O_853,N_9572,N_9156);
or UO_854 (O_854,N_7931,N_9646);
or UO_855 (O_855,N_7701,N_9996);
xor UO_856 (O_856,N_8854,N_9593);
or UO_857 (O_857,N_8996,N_8753);
or UO_858 (O_858,N_9713,N_7586);
nand UO_859 (O_859,N_8446,N_8909);
and UO_860 (O_860,N_8158,N_8586);
xor UO_861 (O_861,N_7937,N_9314);
or UO_862 (O_862,N_9067,N_8062);
nor UO_863 (O_863,N_7678,N_7903);
nand UO_864 (O_864,N_7601,N_7851);
nand UO_865 (O_865,N_8895,N_7998);
or UO_866 (O_866,N_9010,N_8381);
or UO_867 (O_867,N_9772,N_7899);
nand UO_868 (O_868,N_7765,N_8060);
or UO_869 (O_869,N_7526,N_9092);
nor UO_870 (O_870,N_9251,N_9681);
and UO_871 (O_871,N_9153,N_9210);
nor UO_872 (O_872,N_8262,N_8878);
or UO_873 (O_873,N_9699,N_9215);
nand UO_874 (O_874,N_9708,N_8350);
nor UO_875 (O_875,N_9567,N_7796);
nand UO_876 (O_876,N_9759,N_9368);
or UO_877 (O_877,N_9266,N_8011);
nor UO_878 (O_878,N_7793,N_9369);
nand UO_879 (O_879,N_9349,N_8085);
or UO_880 (O_880,N_8704,N_7640);
nand UO_881 (O_881,N_9953,N_9659);
nor UO_882 (O_882,N_8983,N_7502);
nand UO_883 (O_883,N_9011,N_8817);
and UO_884 (O_884,N_9397,N_9497);
or UO_885 (O_885,N_8221,N_8378);
and UO_886 (O_886,N_9419,N_8744);
nand UO_887 (O_887,N_7911,N_7609);
and UO_888 (O_888,N_7790,N_8385);
nor UO_889 (O_889,N_9898,N_9394);
or UO_890 (O_890,N_9788,N_8090);
xor UO_891 (O_891,N_9869,N_8970);
or UO_892 (O_892,N_8562,N_7811);
or UO_893 (O_893,N_7664,N_9524);
nor UO_894 (O_894,N_8301,N_7809);
and UO_895 (O_895,N_8565,N_8924);
or UO_896 (O_896,N_7881,N_9078);
nand UO_897 (O_897,N_7788,N_9662);
and UO_898 (O_898,N_9504,N_9398);
or UO_899 (O_899,N_7647,N_8587);
xnor UO_900 (O_900,N_9977,N_9166);
nand UO_901 (O_901,N_8921,N_9967);
or UO_902 (O_902,N_8525,N_8850);
nand UO_903 (O_903,N_7517,N_9049);
or UO_904 (O_904,N_9458,N_8175);
nor UO_905 (O_905,N_8460,N_8056);
and UO_906 (O_906,N_9274,N_7726);
and UO_907 (O_907,N_9469,N_9568);
and UO_908 (O_908,N_8805,N_8715);
nor UO_909 (O_909,N_7751,N_8461);
nand UO_910 (O_910,N_7806,N_9348);
nand UO_911 (O_911,N_7503,N_7870);
nand UO_912 (O_912,N_9891,N_9313);
and UO_913 (O_913,N_7948,N_8628);
and UO_914 (O_914,N_9725,N_7952);
and UO_915 (O_915,N_9066,N_8186);
nand UO_916 (O_916,N_7627,N_9795);
and UO_917 (O_917,N_7914,N_9031);
nor UO_918 (O_918,N_8964,N_7891);
and UO_919 (O_919,N_9106,N_9549);
or UO_920 (O_920,N_8839,N_8694);
and UO_921 (O_921,N_9121,N_7991);
and UO_922 (O_922,N_7691,N_9326);
or UO_923 (O_923,N_7923,N_8456);
nand UO_924 (O_924,N_7832,N_8558);
and UO_925 (O_925,N_8214,N_7548);
nor UO_926 (O_926,N_8943,N_9282);
or UO_927 (O_927,N_8655,N_9427);
nor UO_928 (O_928,N_8184,N_9920);
nand UO_929 (O_929,N_8209,N_7738);
xnor UO_930 (O_930,N_8129,N_7594);
and UO_931 (O_931,N_9454,N_9966);
nand UO_932 (O_932,N_9056,N_9422);
nor UO_933 (O_933,N_7873,N_9573);
xor UO_934 (O_934,N_8474,N_9527);
and UO_935 (O_935,N_9974,N_8408);
nand UO_936 (O_936,N_8367,N_9300);
nor UO_937 (O_937,N_9843,N_9324);
or UO_938 (O_938,N_9838,N_8202);
nand UO_939 (O_939,N_8851,N_8315);
nand UO_940 (O_940,N_9717,N_8412);
nor UO_941 (O_941,N_7826,N_9350);
nand UO_942 (O_942,N_8917,N_9721);
or UO_943 (O_943,N_8106,N_8316);
and UO_944 (O_944,N_8050,N_9881);
nor UO_945 (O_945,N_9100,N_7885);
xnor UO_946 (O_946,N_9696,N_8524);
nand UO_947 (O_947,N_9163,N_9104);
nor UO_948 (O_948,N_9803,N_9629);
nand UO_949 (O_949,N_9400,N_7571);
and UO_950 (O_950,N_9261,N_7662);
or UO_951 (O_951,N_8898,N_7754);
or UO_952 (O_952,N_8596,N_7978);
nand UO_953 (O_953,N_9478,N_8340);
nand UO_954 (O_954,N_9222,N_8377);
or UO_955 (O_955,N_8906,N_9016);
nor UO_956 (O_956,N_8395,N_7917);
and UO_957 (O_957,N_7996,N_9297);
nor UO_958 (O_958,N_9841,N_8636);
nor UO_959 (O_959,N_8432,N_9495);
nor UO_960 (O_960,N_9462,N_9351);
nor UO_961 (O_961,N_8016,N_8574);
and UO_962 (O_962,N_8932,N_8181);
nand UO_963 (O_963,N_9057,N_7980);
nand UO_964 (O_964,N_7840,N_7680);
or UO_965 (O_965,N_9915,N_9813);
nor UO_966 (O_966,N_7663,N_9023);
nor UO_967 (O_967,N_9911,N_9449);
nor UO_968 (O_968,N_8459,N_9392);
nand UO_969 (O_969,N_7841,N_7830);
nand UO_970 (O_970,N_7757,N_9401);
nor UO_971 (O_971,N_7697,N_9896);
or UO_972 (O_972,N_8406,N_9340);
nor UO_973 (O_973,N_8180,N_9514);
or UO_974 (O_974,N_8732,N_8867);
or UO_975 (O_975,N_9749,N_8807);
nor UO_976 (O_976,N_9037,N_9603);
and UO_977 (O_977,N_8245,N_9145);
and UO_978 (O_978,N_9835,N_9181);
and UO_979 (O_979,N_7702,N_9820);
nand UO_980 (O_980,N_9327,N_8942);
or UO_981 (O_981,N_9094,N_8979);
nand UO_982 (O_982,N_9804,N_9164);
and UO_983 (O_983,N_9520,N_9834);
nand UO_984 (O_984,N_9887,N_8267);
nor UO_985 (O_985,N_9779,N_8969);
nor UO_986 (O_986,N_8475,N_9263);
and UO_987 (O_987,N_9434,N_9558);
and UO_988 (O_988,N_9118,N_8760);
nor UO_989 (O_989,N_8182,N_8143);
and UO_990 (O_990,N_7804,N_7643);
or UO_991 (O_991,N_7836,N_7533);
and UO_992 (O_992,N_7710,N_9285);
nand UO_993 (O_993,N_7703,N_9157);
nand UO_994 (O_994,N_9234,N_9964);
and UO_995 (O_995,N_9275,N_9578);
and UO_996 (O_996,N_8594,N_9903);
nand UO_997 (O_997,N_9616,N_8029);
and UO_998 (O_998,N_9435,N_8237);
nand UO_999 (O_999,N_7929,N_8161);
nand UO_1000 (O_1000,N_9120,N_7673);
and UO_1001 (O_1001,N_7724,N_7988);
and UO_1002 (O_1002,N_9742,N_9230);
nor UO_1003 (O_1003,N_9748,N_9109);
and UO_1004 (O_1004,N_8300,N_9302);
nor UO_1005 (O_1005,N_8634,N_7894);
and UO_1006 (O_1006,N_7596,N_9651);
nor UO_1007 (O_1007,N_9664,N_8567);
or UO_1008 (O_1008,N_9579,N_9374);
xnor UO_1009 (O_1009,N_7600,N_8417);
nor UO_1010 (O_1010,N_8200,N_9047);
and UO_1011 (O_1011,N_8156,N_7875);
or UO_1012 (O_1012,N_8676,N_8579);
and UO_1013 (O_1013,N_8941,N_9357);
nor UO_1014 (O_1014,N_8372,N_8112);
or UO_1015 (O_1015,N_8509,N_7556);
or UO_1016 (O_1016,N_9750,N_9626);
or UO_1017 (O_1017,N_8213,N_7839);
nor UO_1018 (O_1018,N_9459,N_8452);
and UO_1019 (O_1019,N_8539,N_8582);
nand UO_1020 (O_1020,N_8937,N_7650);
and UO_1021 (O_1021,N_7871,N_8918);
or UO_1022 (O_1022,N_9484,N_8600);
nor UO_1023 (O_1023,N_7906,N_9331);
or UO_1024 (O_1024,N_9252,N_9036);
and UO_1025 (O_1025,N_9338,N_9030);
nor UO_1026 (O_1026,N_8226,N_9475);
nand UO_1027 (O_1027,N_9836,N_9358);
nand UO_1028 (O_1028,N_8497,N_7525);
and UO_1029 (O_1029,N_8830,N_9959);
nand UO_1030 (O_1030,N_8212,N_9894);
and UO_1031 (O_1031,N_8764,N_9423);
or UO_1032 (O_1032,N_7545,N_8339);
or UO_1033 (O_1033,N_8057,N_8080);
or UO_1034 (O_1034,N_9584,N_9680);
and UO_1035 (O_1035,N_9218,N_8737);
nand UO_1036 (O_1036,N_9186,N_9359);
or UO_1037 (O_1037,N_8907,N_7794);
nand UO_1038 (O_1038,N_7789,N_8681);
and UO_1039 (O_1039,N_9231,N_7648);
nand UO_1040 (O_1040,N_8376,N_8783);
and UO_1041 (O_1041,N_8861,N_7968);
nor UO_1042 (O_1042,N_9670,N_9995);
nor UO_1043 (O_1043,N_9204,N_8623);
or UO_1044 (O_1044,N_7612,N_8879);
nand UO_1045 (O_1045,N_8507,N_9677);
or UO_1046 (O_1046,N_9165,N_8042);
and UO_1047 (O_1047,N_9732,N_9570);
nand UO_1048 (O_1048,N_8153,N_7890);
nand UO_1049 (O_1049,N_9697,N_8566);
or UO_1050 (O_1050,N_9038,N_9909);
or UO_1051 (O_1051,N_9107,N_9051);
or UO_1052 (O_1052,N_7817,N_9848);
xnor UO_1053 (O_1053,N_7857,N_9264);
or UO_1054 (O_1054,N_8069,N_9361);
xnor UO_1055 (O_1055,N_8260,N_7655);
or UO_1056 (O_1056,N_9232,N_8672);
nor UO_1057 (O_1057,N_8773,N_9418);
nand UO_1058 (O_1058,N_8239,N_9147);
nand UO_1059 (O_1059,N_9185,N_9628);
or UO_1060 (O_1060,N_9970,N_9981);
nor UO_1061 (O_1061,N_8196,N_8740);
nor UO_1062 (O_1062,N_9643,N_7824);
and UO_1063 (O_1063,N_7675,N_9188);
nor UO_1064 (O_1064,N_9322,N_9298);
nor UO_1065 (O_1065,N_8121,N_7861);
nor UO_1066 (O_1066,N_9865,N_9535);
or UO_1067 (O_1067,N_9473,N_8435);
and UO_1068 (O_1068,N_8394,N_9085);
or UO_1069 (O_1069,N_8157,N_8266);
nand UO_1070 (O_1070,N_9095,N_9506);
nor UO_1071 (O_1071,N_8820,N_7803);
nor UO_1072 (O_1072,N_8192,N_9472);
or UO_1073 (O_1073,N_9228,N_8771);
nor UO_1074 (O_1074,N_8662,N_8962);
nand UO_1075 (O_1075,N_9045,N_7853);
nand UO_1076 (O_1076,N_9934,N_8986);
nor UO_1077 (O_1077,N_8127,N_8332);
and UO_1078 (O_1078,N_9982,N_9636);
and UO_1079 (O_1079,N_9990,N_8951);
and UO_1080 (O_1080,N_8868,N_8581);
nor UO_1081 (O_1081,N_8264,N_8598);
or UO_1082 (O_1082,N_8092,N_9884);
nand UO_1083 (O_1083,N_7577,N_9058);
and UO_1084 (O_1084,N_9902,N_9799);
nand UO_1085 (O_1085,N_9176,N_8236);
nor UO_1086 (O_1086,N_9041,N_9002);
or UO_1087 (O_1087,N_8489,N_9597);
or UO_1088 (O_1088,N_9668,N_9299);
xnor UO_1089 (O_1089,N_7993,N_9236);
nand UO_1090 (O_1090,N_8179,N_8716);
and UO_1091 (O_1091,N_8286,N_9711);
or UO_1092 (O_1092,N_8800,N_9774);
and UO_1093 (O_1093,N_7642,N_8160);
nand UO_1094 (O_1094,N_7649,N_8194);
and UO_1095 (O_1095,N_8661,N_9077);
nor UO_1096 (O_1096,N_9024,N_9786);
nor UO_1097 (O_1097,N_7763,N_8255);
or UO_1098 (O_1098,N_9564,N_8349);
xor UO_1099 (O_1099,N_8188,N_9766);
or UO_1100 (O_1100,N_8279,N_9521);
or UO_1101 (O_1101,N_7746,N_8772);
and UO_1102 (O_1102,N_8361,N_9576);
nand UO_1103 (O_1103,N_7549,N_8142);
nor UO_1104 (O_1104,N_8365,N_9090);
nand UO_1105 (O_1105,N_7544,N_9180);
and UO_1106 (O_1106,N_8529,N_9141);
and UO_1107 (O_1107,N_9937,N_7954);
or UO_1108 (O_1108,N_9842,N_8087);
or UO_1109 (O_1109,N_9933,N_8126);
and UO_1110 (O_1110,N_9940,N_8371);
nand UO_1111 (O_1111,N_8848,N_8019);
nor UO_1112 (O_1112,N_7767,N_9621);
nand UO_1113 (O_1113,N_8424,N_7986);
nand UO_1114 (O_1114,N_8605,N_9116);
or UO_1115 (O_1115,N_8317,N_9962);
nor UO_1116 (O_1116,N_8847,N_9242);
nand UO_1117 (O_1117,N_9577,N_8845);
and UO_1118 (O_1118,N_8307,N_8780);
nand UO_1119 (O_1119,N_8048,N_8323);
or UO_1120 (O_1120,N_9101,N_8511);
nand UO_1121 (O_1121,N_9797,N_7551);
xnor UO_1122 (O_1122,N_8748,N_8227);
nor UO_1123 (O_1123,N_9532,N_7882);
nand UO_1124 (O_1124,N_9133,N_9512);
or UO_1125 (O_1125,N_8644,N_8357);
nor UO_1126 (O_1126,N_8051,N_8792);
or UO_1127 (O_1127,N_9135,N_9387);
and UO_1128 (O_1128,N_9777,N_8261);
and UO_1129 (O_1129,N_8645,N_9619);
and UO_1130 (O_1130,N_7932,N_8151);
nand UO_1131 (O_1131,N_8478,N_8420);
nand UO_1132 (O_1132,N_7541,N_9411);
and UO_1133 (O_1133,N_8123,N_8178);
nor UO_1134 (O_1134,N_8689,N_8217);
nand UO_1135 (O_1135,N_8352,N_9726);
or UO_1136 (O_1136,N_9678,N_9455);
and UO_1137 (O_1137,N_9372,N_8635);
or UO_1138 (O_1138,N_9550,N_7787);
nand UO_1139 (O_1139,N_9850,N_7728);
or UO_1140 (O_1140,N_8982,N_7536);
or UO_1141 (O_1141,N_8118,N_8263);
nor UO_1142 (O_1142,N_9935,N_8870);
and UO_1143 (O_1143,N_7630,N_9654);
and UO_1144 (O_1144,N_9710,N_9043);
and UO_1145 (O_1145,N_9830,N_9691);
and UO_1146 (O_1146,N_8794,N_7683);
or UO_1147 (O_1147,N_9998,N_8324);
and UO_1148 (O_1148,N_8823,N_9014);
nand UO_1149 (O_1149,N_8081,N_9365);
nor UO_1150 (O_1150,N_9034,N_8400);
or UO_1151 (O_1151,N_7901,N_8398);
nor UO_1152 (O_1152,N_9375,N_9126);
and UO_1153 (O_1153,N_8633,N_8355);
or UO_1154 (O_1154,N_7593,N_8454);
or UO_1155 (O_1155,N_9613,N_8668);
and UO_1156 (O_1156,N_9924,N_9833);
nor UO_1157 (O_1157,N_8229,N_7699);
and UO_1158 (O_1158,N_8960,N_8536);
nand UO_1159 (O_1159,N_8914,N_9439);
nand UO_1160 (O_1160,N_9856,N_8490);
nand UO_1161 (O_1161,N_8240,N_9110);
or UO_1162 (O_1162,N_8873,N_8705);
nand UO_1163 (O_1163,N_8718,N_9975);
nand UO_1164 (O_1164,N_7989,N_9809);
and UO_1165 (O_1165,N_8271,N_9065);
nand UO_1166 (O_1166,N_8612,N_9602);
and UO_1167 (O_1167,N_7786,N_7845);
nor UO_1168 (O_1168,N_7867,N_7706);
nand UO_1169 (O_1169,N_8609,N_8608);
nand UO_1170 (O_1170,N_8234,N_8103);
or UO_1171 (O_1171,N_9425,N_9003);
nor UO_1172 (O_1172,N_8913,N_9061);
or UO_1173 (O_1173,N_9353,N_8270);
nor UO_1174 (O_1174,N_7810,N_8592);
nand UO_1175 (O_1175,N_8328,N_8849);
nand UO_1176 (O_1176,N_9980,N_9384);
nand UO_1177 (O_1177,N_8409,N_9019);
nor UO_1178 (O_1178,N_8585,N_9383);
nor UO_1179 (O_1179,N_9211,N_7974);
or UO_1180 (O_1180,N_9027,N_9688);
and UO_1181 (O_1181,N_9152,N_9927);
nand UO_1182 (O_1182,N_8485,N_8464);
and UO_1183 (O_1183,N_9256,N_9551);
nand UO_1184 (O_1184,N_8899,N_9614);
nor UO_1185 (O_1185,N_9922,N_9606);
and UO_1186 (O_1186,N_8299,N_9808);
nor UO_1187 (O_1187,N_9071,N_8733);
nand UO_1188 (O_1188,N_8353,N_8065);
nand UO_1189 (O_1189,N_9007,N_8104);
and UO_1190 (O_1190,N_9984,N_9170);
and UO_1191 (O_1191,N_9719,N_8330);
xor UO_1192 (O_1192,N_9805,N_8990);
nor UO_1193 (O_1193,N_9683,N_7527);
nor UO_1194 (O_1194,N_8736,N_7961);
nand UO_1195 (O_1195,N_9523,N_8046);
nor UO_1196 (O_1196,N_9987,N_7979);
and UO_1197 (O_1197,N_9756,N_8150);
and UO_1198 (O_1198,N_9255,N_7572);
and UO_1199 (O_1199,N_8622,N_7570);
nor UO_1200 (O_1200,N_9727,N_7905);
and UO_1201 (O_1201,N_9486,N_9360);
xnor UO_1202 (O_1202,N_9150,N_8094);
xor UO_1203 (O_1203,N_8673,N_9376);
nand UO_1204 (O_1204,N_7935,N_9428);
or UO_1205 (O_1205,N_8064,N_9012);
and UO_1206 (O_1206,N_9665,N_7622);
nand UO_1207 (O_1207,N_8479,N_9901);
nor UO_1208 (O_1208,N_9837,N_7704);
and UO_1209 (O_1209,N_7628,N_8453);
and UO_1210 (O_1210,N_7723,N_8621);
nor UO_1211 (O_1211,N_7966,N_8711);
nor UO_1212 (O_1212,N_9471,N_9942);
and UO_1213 (O_1213,N_7686,N_8749);
nand UO_1214 (O_1214,N_7774,N_9736);
nand UO_1215 (O_1215,N_8883,N_8297);
or UO_1216 (O_1216,N_9199,N_9926);
nand UO_1217 (O_1217,N_9481,N_7823);
and UO_1218 (O_1218,N_9040,N_7920);
and UO_1219 (O_1219,N_8648,N_8649);
nor UO_1220 (O_1220,N_9337,N_9851);
xor UO_1221 (O_1221,N_8333,N_8901);
or UO_1222 (O_1222,N_8082,N_7700);
nand UO_1223 (O_1223,N_9395,N_9910);
nor UO_1224 (O_1224,N_7719,N_8290);
or UO_1225 (O_1225,N_9528,N_7801);
or UO_1226 (O_1226,N_9196,N_9874);
nor UO_1227 (O_1227,N_8745,N_7828);
and UO_1228 (O_1228,N_7791,N_9184);
or UO_1229 (O_1229,N_7537,N_8860);
nor UO_1230 (O_1230,N_7575,N_8375);
or UO_1231 (O_1231,N_9961,N_8444);
nand UO_1232 (O_1232,N_9821,N_8627);
or UO_1233 (O_1233,N_8079,N_8162);
or UO_1234 (O_1234,N_7846,N_8078);
nor UO_1235 (O_1235,N_7773,N_9548);
or UO_1236 (O_1236,N_8288,N_9291);
or UO_1237 (O_1237,N_8110,N_8295);
or UO_1238 (O_1238,N_8746,N_9385);
nor UO_1239 (O_1239,N_7511,N_8441);
xnor UO_1240 (O_1240,N_8374,N_7580);
nand UO_1241 (O_1241,N_8045,N_9862);
or UO_1242 (O_1242,N_8313,N_9050);
nor UO_1243 (O_1243,N_9482,N_9354);
nor UO_1244 (O_1244,N_7520,N_8856);
and UO_1245 (O_1245,N_7722,N_8963);
nor UO_1246 (O_1246,N_7530,N_7945);
and UO_1247 (O_1247,N_9086,N_9496);
nor UO_1248 (O_1248,N_7603,N_8729);
and UO_1249 (O_1249,N_9259,N_8742);
or UO_1250 (O_1250,N_9173,N_8280);
and UO_1251 (O_1251,N_7793,N_9224);
nand UO_1252 (O_1252,N_9623,N_9103);
nand UO_1253 (O_1253,N_9684,N_7948);
nand UO_1254 (O_1254,N_8820,N_7920);
nor UO_1255 (O_1255,N_7778,N_9298);
and UO_1256 (O_1256,N_8085,N_8285);
and UO_1257 (O_1257,N_9942,N_9227);
or UO_1258 (O_1258,N_8845,N_9513);
and UO_1259 (O_1259,N_8503,N_9024);
and UO_1260 (O_1260,N_8180,N_7953);
or UO_1261 (O_1261,N_8634,N_8558);
and UO_1262 (O_1262,N_9102,N_9714);
or UO_1263 (O_1263,N_9480,N_9434);
nand UO_1264 (O_1264,N_8467,N_8907);
xor UO_1265 (O_1265,N_8205,N_8174);
nor UO_1266 (O_1266,N_8098,N_9754);
and UO_1267 (O_1267,N_9326,N_8907);
nor UO_1268 (O_1268,N_7684,N_8752);
and UO_1269 (O_1269,N_8875,N_8011);
nor UO_1270 (O_1270,N_7609,N_7845);
nor UO_1271 (O_1271,N_8434,N_8239);
nand UO_1272 (O_1272,N_9268,N_8683);
and UO_1273 (O_1273,N_7757,N_9294);
and UO_1274 (O_1274,N_8912,N_9482);
or UO_1275 (O_1275,N_9755,N_7829);
or UO_1276 (O_1276,N_8234,N_9954);
or UO_1277 (O_1277,N_9778,N_8361);
nor UO_1278 (O_1278,N_9051,N_8253);
or UO_1279 (O_1279,N_9629,N_8337);
nand UO_1280 (O_1280,N_8777,N_9079);
nand UO_1281 (O_1281,N_8113,N_7532);
or UO_1282 (O_1282,N_7696,N_8452);
or UO_1283 (O_1283,N_8918,N_9020);
and UO_1284 (O_1284,N_9923,N_9130);
or UO_1285 (O_1285,N_9917,N_9587);
or UO_1286 (O_1286,N_9002,N_8624);
nor UO_1287 (O_1287,N_8833,N_7730);
and UO_1288 (O_1288,N_9772,N_8627);
or UO_1289 (O_1289,N_8787,N_9476);
nor UO_1290 (O_1290,N_8935,N_9249);
nor UO_1291 (O_1291,N_7596,N_9626);
nor UO_1292 (O_1292,N_7599,N_9553);
or UO_1293 (O_1293,N_8067,N_8787);
or UO_1294 (O_1294,N_8719,N_8255);
nor UO_1295 (O_1295,N_8380,N_7749);
or UO_1296 (O_1296,N_9745,N_8397);
and UO_1297 (O_1297,N_7912,N_9953);
nand UO_1298 (O_1298,N_8701,N_9952);
nor UO_1299 (O_1299,N_9669,N_8045);
or UO_1300 (O_1300,N_8908,N_7655);
and UO_1301 (O_1301,N_9421,N_8868);
or UO_1302 (O_1302,N_8131,N_8008);
or UO_1303 (O_1303,N_7810,N_9482);
nor UO_1304 (O_1304,N_9399,N_8426);
and UO_1305 (O_1305,N_8041,N_8397);
nor UO_1306 (O_1306,N_9323,N_9300);
and UO_1307 (O_1307,N_7624,N_9965);
or UO_1308 (O_1308,N_9560,N_8858);
nand UO_1309 (O_1309,N_9014,N_8454);
nand UO_1310 (O_1310,N_9088,N_9367);
and UO_1311 (O_1311,N_9858,N_8277);
and UO_1312 (O_1312,N_7867,N_8801);
or UO_1313 (O_1313,N_8150,N_9002);
nor UO_1314 (O_1314,N_9240,N_8751);
nand UO_1315 (O_1315,N_7633,N_9536);
or UO_1316 (O_1316,N_9187,N_8021);
nor UO_1317 (O_1317,N_9439,N_8613);
or UO_1318 (O_1318,N_7972,N_8844);
nor UO_1319 (O_1319,N_8025,N_9293);
nand UO_1320 (O_1320,N_9274,N_8078);
nor UO_1321 (O_1321,N_7732,N_9026);
and UO_1322 (O_1322,N_8747,N_9255);
nand UO_1323 (O_1323,N_8526,N_9839);
or UO_1324 (O_1324,N_7989,N_9980);
or UO_1325 (O_1325,N_8429,N_7869);
and UO_1326 (O_1326,N_9170,N_9902);
or UO_1327 (O_1327,N_8966,N_8829);
or UO_1328 (O_1328,N_7638,N_8727);
nor UO_1329 (O_1329,N_8489,N_8657);
or UO_1330 (O_1330,N_8128,N_8978);
xnor UO_1331 (O_1331,N_9017,N_7718);
and UO_1332 (O_1332,N_8779,N_7903);
or UO_1333 (O_1333,N_9575,N_9014);
nand UO_1334 (O_1334,N_9482,N_8934);
nor UO_1335 (O_1335,N_8566,N_9915);
nand UO_1336 (O_1336,N_9167,N_8225);
nand UO_1337 (O_1337,N_9498,N_9651);
or UO_1338 (O_1338,N_9388,N_9455);
or UO_1339 (O_1339,N_8467,N_8221);
and UO_1340 (O_1340,N_8295,N_9757);
nor UO_1341 (O_1341,N_9999,N_9348);
and UO_1342 (O_1342,N_9783,N_9588);
nor UO_1343 (O_1343,N_8321,N_9304);
or UO_1344 (O_1344,N_8403,N_8582);
or UO_1345 (O_1345,N_7942,N_9132);
or UO_1346 (O_1346,N_9141,N_8686);
and UO_1347 (O_1347,N_8502,N_9697);
nand UO_1348 (O_1348,N_8548,N_9064);
nor UO_1349 (O_1349,N_7859,N_9335);
nor UO_1350 (O_1350,N_8856,N_9214);
nor UO_1351 (O_1351,N_9294,N_9553);
nor UO_1352 (O_1352,N_8424,N_9946);
and UO_1353 (O_1353,N_8753,N_9950);
and UO_1354 (O_1354,N_8328,N_8527);
nand UO_1355 (O_1355,N_8313,N_8569);
and UO_1356 (O_1356,N_9538,N_8196);
nand UO_1357 (O_1357,N_9941,N_8585);
or UO_1358 (O_1358,N_8799,N_8761);
or UO_1359 (O_1359,N_9762,N_8904);
nor UO_1360 (O_1360,N_9948,N_8337);
nand UO_1361 (O_1361,N_8713,N_7576);
nor UO_1362 (O_1362,N_7904,N_9796);
and UO_1363 (O_1363,N_8743,N_8410);
and UO_1364 (O_1364,N_9594,N_9645);
nor UO_1365 (O_1365,N_8878,N_8757);
and UO_1366 (O_1366,N_8603,N_7948);
nand UO_1367 (O_1367,N_9310,N_9211);
nor UO_1368 (O_1368,N_9676,N_9352);
nand UO_1369 (O_1369,N_7633,N_9375);
and UO_1370 (O_1370,N_8609,N_9858);
nor UO_1371 (O_1371,N_8293,N_7852);
or UO_1372 (O_1372,N_9482,N_7985);
or UO_1373 (O_1373,N_9392,N_9691);
nand UO_1374 (O_1374,N_8456,N_8613);
and UO_1375 (O_1375,N_8241,N_8585);
or UO_1376 (O_1376,N_7799,N_8463);
nand UO_1377 (O_1377,N_7699,N_9787);
nand UO_1378 (O_1378,N_9271,N_8920);
nor UO_1379 (O_1379,N_7789,N_7902);
nor UO_1380 (O_1380,N_9286,N_9871);
or UO_1381 (O_1381,N_8234,N_8878);
or UO_1382 (O_1382,N_9178,N_9988);
xor UO_1383 (O_1383,N_9938,N_8404);
nand UO_1384 (O_1384,N_8949,N_9243);
nor UO_1385 (O_1385,N_8225,N_9166);
and UO_1386 (O_1386,N_7880,N_9528);
nor UO_1387 (O_1387,N_7840,N_8457);
or UO_1388 (O_1388,N_8666,N_7774);
and UO_1389 (O_1389,N_7848,N_9271);
nor UO_1390 (O_1390,N_8615,N_7672);
xor UO_1391 (O_1391,N_8273,N_7619);
or UO_1392 (O_1392,N_7843,N_9923);
nor UO_1393 (O_1393,N_7731,N_8907);
nand UO_1394 (O_1394,N_9011,N_8913);
nand UO_1395 (O_1395,N_8840,N_7582);
nand UO_1396 (O_1396,N_8662,N_7811);
nor UO_1397 (O_1397,N_7519,N_9196);
nor UO_1398 (O_1398,N_9606,N_7549);
or UO_1399 (O_1399,N_8909,N_9899);
or UO_1400 (O_1400,N_9331,N_9135);
nand UO_1401 (O_1401,N_9477,N_8245);
nand UO_1402 (O_1402,N_9287,N_7870);
or UO_1403 (O_1403,N_8566,N_9598);
nor UO_1404 (O_1404,N_9358,N_9015);
nand UO_1405 (O_1405,N_8946,N_8790);
and UO_1406 (O_1406,N_8690,N_9511);
or UO_1407 (O_1407,N_8599,N_9300);
or UO_1408 (O_1408,N_7878,N_9505);
nor UO_1409 (O_1409,N_8837,N_9185);
and UO_1410 (O_1410,N_9316,N_7742);
nor UO_1411 (O_1411,N_7722,N_9574);
nand UO_1412 (O_1412,N_8436,N_9974);
and UO_1413 (O_1413,N_8786,N_9370);
nand UO_1414 (O_1414,N_9448,N_8568);
and UO_1415 (O_1415,N_8068,N_8444);
nand UO_1416 (O_1416,N_9457,N_9594);
and UO_1417 (O_1417,N_9408,N_9001);
nand UO_1418 (O_1418,N_8630,N_9492);
nor UO_1419 (O_1419,N_8473,N_8063);
or UO_1420 (O_1420,N_8099,N_8806);
and UO_1421 (O_1421,N_7735,N_8164);
nand UO_1422 (O_1422,N_9840,N_7837);
xor UO_1423 (O_1423,N_9386,N_9294);
nor UO_1424 (O_1424,N_7962,N_8213);
and UO_1425 (O_1425,N_9778,N_7589);
nand UO_1426 (O_1426,N_8422,N_8478);
nand UO_1427 (O_1427,N_8530,N_8977);
or UO_1428 (O_1428,N_7915,N_8842);
or UO_1429 (O_1429,N_8392,N_7525);
xnor UO_1430 (O_1430,N_9729,N_8823);
or UO_1431 (O_1431,N_9670,N_8953);
and UO_1432 (O_1432,N_9895,N_8646);
xnor UO_1433 (O_1433,N_9112,N_9206);
or UO_1434 (O_1434,N_9355,N_8132);
or UO_1435 (O_1435,N_9767,N_8711);
or UO_1436 (O_1436,N_9391,N_7724);
nor UO_1437 (O_1437,N_9528,N_8074);
xnor UO_1438 (O_1438,N_8246,N_8299);
or UO_1439 (O_1439,N_9207,N_7831);
nor UO_1440 (O_1440,N_9251,N_9943);
and UO_1441 (O_1441,N_8661,N_8536);
and UO_1442 (O_1442,N_8792,N_7714);
and UO_1443 (O_1443,N_8019,N_8741);
and UO_1444 (O_1444,N_9430,N_7850);
nand UO_1445 (O_1445,N_8007,N_7756);
or UO_1446 (O_1446,N_8040,N_9119);
nand UO_1447 (O_1447,N_8293,N_8144);
nand UO_1448 (O_1448,N_9151,N_9317);
nand UO_1449 (O_1449,N_9453,N_9921);
and UO_1450 (O_1450,N_8132,N_9915);
and UO_1451 (O_1451,N_9593,N_7522);
nand UO_1452 (O_1452,N_8924,N_8952);
nor UO_1453 (O_1453,N_7990,N_8141);
or UO_1454 (O_1454,N_9923,N_8112);
nor UO_1455 (O_1455,N_7761,N_8832);
and UO_1456 (O_1456,N_8399,N_8451);
and UO_1457 (O_1457,N_8037,N_7705);
or UO_1458 (O_1458,N_7986,N_8503);
and UO_1459 (O_1459,N_7854,N_8234);
and UO_1460 (O_1460,N_7685,N_7850);
nor UO_1461 (O_1461,N_9950,N_8488);
and UO_1462 (O_1462,N_8058,N_8456);
nand UO_1463 (O_1463,N_9034,N_8751);
xor UO_1464 (O_1464,N_8731,N_7811);
nor UO_1465 (O_1465,N_7733,N_9359);
and UO_1466 (O_1466,N_9181,N_8071);
nor UO_1467 (O_1467,N_9633,N_7563);
nand UO_1468 (O_1468,N_9678,N_7940);
nor UO_1469 (O_1469,N_8024,N_9210);
xnor UO_1470 (O_1470,N_9828,N_8247);
nor UO_1471 (O_1471,N_9964,N_9216);
nor UO_1472 (O_1472,N_8916,N_7659);
or UO_1473 (O_1473,N_8387,N_8366);
nand UO_1474 (O_1474,N_8661,N_9861);
nand UO_1475 (O_1475,N_7579,N_7572);
and UO_1476 (O_1476,N_7518,N_8479);
xnor UO_1477 (O_1477,N_9525,N_8252);
or UO_1478 (O_1478,N_7932,N_9584);
and UO_1479 (O_1479,N_7612,N_9970);
and UO_1480 (O_1480,N_9518,N_7949);
or UO_1481 (O_1481,N_8536,N_7634);
or UO_1482 (O_1482,N_8744,N_8981);
nand UO_1483 (O_1483,N_9265,N_7613);
nand UO_1484 (O_1484,N_9469,N_9558);
and UO_1485 (O_1485,N_7904,N_8399);
or UO_1486 (O_1486,N_9481,N_7857);
or UO_1487 (O_1487,N_7973,N_8713);
and UO_1488 (O_1488,N_9709,N_8394);
or UO_1489 (O_1489,N_8010,N_8348);
or UO_1490 (O_1490,N_9957,N_8052);
or UO_1491 (O_1491,N_9499,N_9462);
nor UO_1492 (O_1492,N_9374,N_8017);
nand UO_1493 (O_1493,N_9180,N_9147);
nand UO_1494 (O_1494,N_7658,N_8664);
and UO_1495 (O_1495,N_8924,N_7994);
or UO_1496 (O_1496,N_9126,N_7572);
and UO_1497 (O_1497,N_9050,N_9168);
nand UO_1498 (O_1498,N_8396,N_9143);
nand UO_1499 (O_1499,N_9998,N_8130);
endmodule