module basic_750_5000_1000_25_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_735,In_356);
nor U1 (N_1,In_148,In_526);
or U2 (N_2,In_407,In_0);
xnor U3 (N_3,In_1,In_646);
and U4 (N_4,In_524,In_691);
or U5 (N_5,In_465,In_500);
nor U6 (N_6,In_583,In_170);
nand U7 (N_7,In_687,In_121);
or U8 (N_8,In_80,In_554);
and U9 (N_9,In_579,In_580);
or U10 (N_10,In_661,In_479);
or U11 (N_11,In_74,In_634);
nor U12 (N_12,In_701,In_330);
or U13 (N_13,In_532,In_262);
or U14 (N_14,In_671,In_615);
nand U15 (N_15,In_42,In_582);
nand U16 (N_16,In_221,In_313);
nor U17 (N_17,In_567,In_405);
or U18 (N_18,In_429,In_46);
nand U19 (N_19,In_557,In_723);
or U20 (N_20,In_450,In_627);
xor U21 (N_21,In_527,In_112);
or U22 (N_22,In_435,In_499);
or U23 (N_23,In_288,In_252);
nand U24 (N_24,In_54,In_482);
and U25 (N_25,In_133,In_111);
nor U26 (N_26,In_13,In_53);
nand U27 (N_27,In_144,In_726);
nand U28 (N_28,In_572,In_180);
or U29 (N_29,In_529,In_169);
or U30 (N_30,In_394,In_264);
and U31 (N_31,In_707,In_365);
nand U32 (N_32,In_430,In_519);
and U33 (N_33,In_584,In_103);
or U34 (N_34,In_421,In_127);
or U35 (N_35,In_623,In_680);
and U36 (N_36,In_190,In_402);
or U37 (N_37,In_420,In_652);
and U38 (N_38,In_94,In_391);
and U39 (N_39,In_724,In_64);
and U40 (N_40,In_125,In_152);
or U41 (N_41,In_9,In_19);
nor U42 (N_42,In_88,In_145);
nand U43 (N_43,In_534,In_352);
and U44 (N_44,In_236,In_281);
nor U45 (N_45,In_558,In_643);
nor U46 (N_46,In_495,In_697);
or U47 (N_47,In_187,In_101);
and U48 (N_48,In_59,In_569);
nand U49 (N_49,In_209,In_475);
nand U50 (N_50,In_685,In_107);
nand U51 (N_51,In_503,In_740);
or U52 (N_52,In_174,In_415);
and U53 (N_53,In_162,In_681);
or U54 (N_54,In_164,In_630);
and U55 (N_55,In_73,In_218);
and U56 (N_56,In_449,In_275);
nand U57 (N_57,In_538,In_16);
and U58 (N_58,In_361,In_206);
and U59 (N_59,In_219,In_314);
nor U60 (N_60,In_151,In_466);
or U61 (N_61,In_26,In_179);
nand U62 (N_62,In_158,In_291);
nand U63 (N_63,In_292,In_674);
and U64 (N_64,In_709,In_633);
nor U65 (N_65,In_510,In_478);
nor U66 (N_66,In_11,In_22);
or U67 (N_67,In_310,In_416);
and U68 (N_68,In_24,In_381);
or U69 (N_69,In_520,In_290);
nor U70 (N_70,In_531,In_596);
and U71 (N_71,In_181,In_473);
xor U72 (N_72,In_142,In_85);
nor U73 (N_73,In_620,In_120);
nor U74 (N_74,In_703,In_632);
nor U75 (N_75,In_146,In_637);
and U76 (N_76,In_102,In_340);
and U77 (N_77,In_344,In_258);
nor U78 (N_78,In_669,In_679);
nor U79 (N_79,In_114,In_207);
or U80 (N_80,In_182,In_55);
and U81 (N_81,In_624,In_692);
or U82 (N_82,In_476,In_561);
nand U83 (N_83,In_666,In_123);
nor U84 (N_84,In_149,In_617);
nand U85 (N_85,In_303,In_237);
nand U86 (N_86,In_18,In_463);
nand U87 (N_87,In_338,In_300);
nor U88 (N_88,In_548,In_15);
nor U89 (N_89,In_447,In_157);
nand U90 (N_90,In_698,In_48);
nor U91 (N_91,In_193,In_651);
nor U92 (N_92,In_550,In_585);
or U93 (N_93,In_222,In_342);
nor U94 (N_94,In_555,In_660);
nor U95 (N_95,In_382,In_343);
or U96 (N_96,In_571,In_371);
and U97 (N_97,In_368,In_166);
or U98 (N_98,In_460,In_595);
and U99 (N_99,In_270,In_594);
and U100 (N_100,In_605,In_17);
nor U101 (N_101,In_434,In_335);
nor U102 (N_102,In_639,In_433);
nand U103 (N_103,In_717,In_189);
nand U104 (N_104,In_483,In_119);
nand U105 (N_105,In_197,In_325);
and U106 (N_106,In_367,In_665);
and U107 (N_107,In_67,In_250);
or U108 (N_108,In_192,In_204);
or U109 (N_109,In_577,In_556);
and U110 (N_110,In_86,In_686);
nor U111 (N_111,In_84,In_497);
nand U112 (N_112,In_467,In_432);
or U113 (N_113,In_241,In_737);
and U114 (N_114,In_25,In_654);
and U115 (N_115,In_183,In_684);
or U116 (N_116,In_379,In_484);
nand U117 (N_117,In_592,In_663);
nand U118 (N_118,In_372,In_513);
nand U119 (N_119,In_259,In_511);
and U120 (N_120,In_89,In_211);
or U121 (N_121,In_159,In_109);
nor U122 (N_122,In_129,In_688);
nand U123 (N_123,In_140,In_357);
nand U124 (N_124,In_280,In_648);
nand U125 (N_125,In_227,In_235);
nand U126 (N_126,In_456,In_202);
nor U127 (N_127,In_323,In_58);
and U128 (N_128,In_732,In_733);
nor U129 (N_129,In_738,In_441);
nand U130 (N_130,In_619,In_100);
nand U131 (N_131,In_134,In_165);
nor U132 (N_132,In_71,In_494);
nand U133 (N_133,In_150,In_588);
xnor U134 (N_134,In_163,In_366);
nand U135 (N_135,In_44,In_355);
or U136 (N_136,In_505,In_216);
nor U137 (N_137,In_161,In_574);
nand U138 (N_138,In_345,In_5);
or U139 (N_139,In_563,In_12);
nor U140 (N_140,In_198,In_126);
nand U141 (N_141,In_647,In_385);
nand U142 (N_142,In_747,In_535);
nor U143 (N_143,In_279,In_399);
and U144 (N_144,In_650,In_224);
or U145 (N_145,In_72,In_742);
or U146 (N_146,In_283,In_70);
nor U147 (N_147,In_228,In_409);
or U148 (N_148,In_455,In_546);
or U149 (N_149,In_358,In_457);
nor U150 (N_150,In_33,In_502);
or U151 (N_151,In_589,In_454);
or U152 (N_152,In_286,In_676);
nand U153 (N_153,In_570,In_263);
nand U154 (N_154,In_50,In_348);
and U155 (N_155,In_299,In_136);
nand U156 (N_156,In_445,In_746);
nor U157 (N_157,In_4,In_631);
nor U158 (N_158,In_736,In_285);
or U159 (N_159,In_614,In_253);
nand U160 (N_160,In_408,In_506);
nor U161 (N_161,In_400,In_269);
nand U162 (N_162,In_184,In_425);
or U163 (N_163,In_346,In_629);
nand U164 (N_164,In_375,In_451);
and U165 (N_165,In_373,In_79);
and U166 (N_166,In_199,In_251);
or U167 (N_167,In_234,In_390);
and U168 (N_168,In_98,In_131);
nor U169 (N_169,In_316,In_468);
nand U170 (N_170,In_38,In_713);
nand U171 (N_171,In_196,In_522);
nor U172 (N_172,In_370,In_734);
or U173 (N_173,In_745,In_20);
and U174 (N_174,In_641,In_477);
or U175 (N_175,In_124,In_223);
nor U176 (N_176,In_37,In_28);
nor U177 (N_177,In_62,In_139);
nand U178 (N_178,In_712,In_160);
or U179 (N_179,In_312,In_35);
xor U180 (N_180,In_718,In_377);
or U181 (N_181,In_655,In_444);
or U182 (N_182,In_528,In_374);
nor U183 (N_183,In_599,In_256);
nand U184 (N_184,In_530,In_29);
and U185 (N_185,In_81,In_118);
nor U186 (N_186,In_622,In_297);
or U187 (N_187,In_398,In_568);
nand U188 (N_188,In_326,In_353);
and U189 (N_189,In_339,In_99);
and U190 (N_190,In_474,In_659);
and U191 (N_191,In_267,In_135);
or U192 (N_192,In_254,In_683);
nor U193 (N_193,In_284,In_21);
or U194 (N_194,In_308,In_512);
or U195 (N_195,In_39,In_501);
or U196 (N_196,In_294,In_272);
nand U197 (N_197,In_644,In_255);
nand U198 (N_198,In_699,In_591);
and U199 (N_199,In_2,In_7);
or U200 (N_200,N_73,N_65);
or U201 (N_201,In_606,In_489);
nor U202 (N_202,In_231,N_85);
or U203 (N_203,In_401,N_11);
or U204 (N_204,In_56,In_616);
or U205 (N_205,In_113,In_329);
and U206 (N_206,N_189,In_274);
and U207 (N_207,N_135,N_46);
or U208 (N_208,In_387,N_76);
nor U209 (N_209,N_54,In_396);
and U210 (N_210,In_265,N_82);
nand U211 (N_211,In_544,In_682);
or U212 (N_212,N_10,In_298);
nor U213 (N_213,N_112,In_551);
or U214 (N_214,In_66,In_384);
or U215 (N_215,In_191,In_76);
nand U216 (N_216,In_749,N_142);
nand U217 (N_217,In_458,In_741);
or U218 (N_218,N_89,In_731);
nand U219 (N_219,N_184,N_64);
nor U220 (N_220,In_155,In_635);
or U221 (N_221,In_34,In_725);
and U222 (N_222,In_410,In_404);
and U223 (N_223,In_452,In_716);
nand U224 (N_224,N_24,N_134);
nor U225 (N_225,N_186,In_287);
nor U226 (N_226,In_47,N_138);
nor U227 (N_227,N_172,N_106);
nor U228 (N_228,In_257,In_696);
and U229 (N_229,In_156,In_130);
or U230 (N_230,N_192,In_30);
nor U231 (N_231,In_675,In_271);
nor U232 (N_232,N_50,In_436);
nand U233 (N_233,In_645,In_115);
and U234 (N_234,N_109,N_77);
or U235 (N_235,In_657,In_60);
and U236 (N_236,In_293,In_442);
nand U237 (N_237,In_260,N_165);
nand U238 (N_238,In_320,N_70);
and U239 (N_239,In_302,In_273);
or U240 (N_240,In_542,N_16);
nand U241 (N_241,In_453,In_75);
nor U242 (N_242,In_147,In_45);
nor U243 (N_243,In_32,N_79);
and U244 (N_244,In_137,N_68);
nor U245 (N_245,N_183,N_20);
nand U246 (N_246,In_203,In_612);
and U247 (N_247,In_278,In_440);
nand U248 (N_248,N_80,In_87);
nand U249 (N_249,In_498,In_266);
and U250 (N_250,N_93,N_196);
and U251 (N_251,In_277,In_138);
or U252 (N_252,N_181,In_201);
nor U253 (N_253,N_8,N_101);
nand U254 (N_254,N_40,In_743);
nor U255 (N_255,In_406,N_69);
nand U256 (N_256,In_610,N_94);
or U257 (N_257,N_115,In_230);
nand U258 (N_258,In_694,N_177);
nand U259 (N_259,In_350,N_22);
and U260 (N_260,In_378,In_496);
or U261 (N_261,N_168,In_173);
nor U262 (N_262,In_564,In_188);
or U263 (N_263,In_508,N_42);
nor U264 (N_264,N_17,In_347);
nor U265 (N_265,N_125,N_27);
nor U266 (N_266,In_351,In_493);
and U267 (N_267,In_10,In_176);
nor U268 (N_268,N_104,In_448);
or U269 (N_269,In_678,In_491);
and U270 (N_270,In_186,N_30);
nand U271 (N_271,N_75,In_472);
or U272 (N_272,In_178,N_56);
nand U273 (N_273,In_708,In_593);
and U274 (N_274,In_702,In_296);
nor U275 (N_275,In_248,N_136);
or U276 (N_276,In_600,N_72);
and U277 (N_277,In_658,N_170);
or U278 (N_278,N_148,N_57);
nor U279 (N_279,N_151,In_319);
and U280 (N_280,In_249,N_55);
nor U281 (N_281,In_232,In_225);
or U282 (N_282,In_93,N_83);
nand U283 (N_283,N_120,In_462);
nor U284 (N_284,N_92,In_553);
nand U285 (N_285,In_311,N_121);
xor U286 (N_286,In_380,N_132);
and U287 (N_287,In_649,N_139);
nand U288 (N_288,N_71,In_324);
or U289 (N_289,N_0,In_672);
nor U290 (N_290,In_597,In_525);
nand U291 (N_291,In_431,In_705);
or U292 (N_292,In_322,In_744);
or U293 (N_293,In_565,N_4);
nor U294 (N_294,In_306,N_198);
or U295 (N_295,In_172,In_307);
or U296 (N_296,In_559,In_90);
nor U297 (N_297,N_44,N_131);
and U298 (N_298,In_6,In_243);
or U299 (N_299,In_461,In_309);
or U300 (N_300,In_437,N_52);
or U301 (N_301,In_389,N_164);
nor U302 (N_302,In_341,N_23);
or U303 (N_303,In_673,N_188);
nand U304 (N_304,In_586,N_197);
or U305 (N_305,In_562,In_656);
or U306 (N_306,N_36,N_173);
nor U307 (N_307,In_321,In_504);
nand U308 (N_308,N_74,N_111);
or U309 (N_309,In_167,In_486);
or U310 (N_310,In_695,In_573);
and U311 (N_311,N_37,In_383);
nand U312 (N_312,In_68,N_43);
and U313 (N_313,In_194,In_51);
and U314 (N_314,N_147,N_9);
nor U315 (N_315,N_174,N_47);
or U316 (N_316,N_124,In_412);
or U317 (N_317,In_245,In_552);
xor U318 (N_318,In_443,N_150);
nand U319 (N_319,In_560,In_69);
nor U320 (N_320,In_195,In_422);
and U321 (N_321,N_144,N_117);
or U322 (N_322,In_485,In_57);
or U323 (N_323,In_471,In_369);
or U324 (N_324,N_155,In_327);
and U325 (N_325,In_693,N_116);
and U326 (N_326,In_481,In_514);
nor U327 (N_327,In_141,In_185);
or U328 (N_328,In_536,In_719);
nor U329 (N_329,N_166,In_545);
nor U330 (N_330,N_86,In_305);
nor U331 (N_331,In_247,N_32);
or U332 (N_332,In_83,In_690);
nand U333 (N_333,In_14,In_8);
and U334 (N_334,In_428,N_98);
or U335 (N_335,In_268,In_598);
and U336 (N_336,N_193,N_103);
or U337 (N_337,N_38,N_169);
and U338 (N_338,N_108,N_91);
and U339 (N_339,In_419,In_439);
nand U340 (N_340,In_364,N_59);
and U341 (N_341,N_18,In_613);
nor U342 (N_342,In_446,In_41);
nor U343 (N_343,N_58,N_180);
nor U344 (N_344,In_540,N_122);
nand U345 (N_345,N_154,N_195);
nand U346 (N_346,In_168,N_45);
nand U347 (N_347,In_214,N_129);
and U348 (N_348,In_229,N_102);
or U349 (N_349,In_360,In_470);
nor U350 (N_350,N_126,In_464);
or U351 (N_351,In_331,In_132);
nor U352 (N_352,In_547,In_608);
nor U353 (N_353,N_15,In_362);
or U354 (N_354,N_21,N_149);
or U355 (N_355,In_43,In_507);
or U356 (N_356,In_122,In_246);
nand U357 (N_357,N_12,N_113);
and U358 (N_358,N_191,In_618);
and U359 (N_359,In_376,In_244);
and U360 (N_360,In_304,In_77);
and U361 (N_361,In_108,N_97);
and U362 (N_362,In_727,In_226);
nor U363 (N_363,In_337,N_95);
and U364 (N_364,N_123,In_411);
and U365 (N_365,In_541,N_187);
or U366 (N_366,In_576,In_354);
and U367 (N_367,In_233,In_607);
and U368 (N_368,In_700,N_81);
nor U369 (N_369,In_328,In_105);
nand U370 (N_370,N_185,N_175);
or U371 (N_371,In_662,In_143);
or U372 (N_372,In_642,In_636);
nor U373 (N_373,N_35,N_29);
and U374 (N_374,In_480,In_36);
or U375 (N_375,In_609,In_706);
nor U376 (N_376,N_163,In_729);
or U377 (N_377,In_677,In_336);
nor U378 (N_378,In_392,In_213);
nand U379 (N_379,N_84,In_714);
or U380 (N_380,In_578,In_276);
nand U381 (N_381,N_190,In_587);
nand U382 (N_382,N_130,In_239);
or U383 (N_383,N_160,N_162);
and U384 (N_384,N_14,In_533);
and U385 (N_385,In_418,N_176);
nor U386 (N_386,In_516,In_171);
nand U387 (N_387,N_6,N_153);
and U388 (N_388,In_413,In_704);
and U389 (N_389,N_159,In_730);
nand U390 (N_390,In_625,In_549);
nor U391 (N_391,N_105,N_48);
and U392 (N_392,N_100,N_145);
nor U393 (N_393,In_110,N_2);
nor U394 (N_394,In_117,In_317);
and U395 (N_395,N_78,N_152);
nand U396 (N_396,In_363,N_141);
nor U397 (N_397,In_82,N_51);
and U398 (N_398,N_118,In_626);
nand U399 (N_399,N_157,N_60);
or U400 (N_400,N_194,In_739);
nor U401 (N_401,In_515,N_26);
or U402 (N_402,In_91,N_221);
or U403 (N_403,N_372,In_200);
nand U404 (N_404,N_369,In_217);
nand U405 (N_405,N_365,N_363);
and U406 (N_406,N_88,In_96);
nand U407 (N_407,N_167,In_23);
or U408 (N_408,N_99,In_397);
or U409 (N_409,N_326,N_272);
xor U410 (N_410,N_255,In_488);
and U411 (N_411,In_517,N_358);
nand U412 (N_412,In_242,N_41);
or U413 (N_413,N_210,In_469);
nand U414 (N_414,In_359,N_323);
or U415 (N_415,N_220,N_204);
nand U416 (N_416,N_355,N_333);
nor U417 (N_417,N_203,N_302);
nor U418 (N_418,In_52,In_566);
nor U419 (N_419,N_211,In_689);
or U420 (N_420,In_537,N_212);
or U421 (N_421,N_327,N_274);
nand U422 (N_422,In_3,In_175);
or U423 (N_423,In_403,N_291);
and U424 (N_424,N_298,In_590);
nand U425 (N_425,N_354,N_280);
nor U426 (N_426,In_459,N_228);
or U427 (N_427,N_119,N_156);
or U428 (N_428,N_63,N_347);
or U429 (N_429,In_386,N_215);
or U430 (N_430,In_289,In_492);
nand U431 (N_431,N_345,N_143);
and U432 (N_432,N_290,N_205);
nand U433 (N_433,N_246,In_295);
and U434 (N_434,N_178,N_268);
or U435 (N_435,N_305,In_261);
nand U436 (N_436,In_424,N_295);
or U437 (N_437,In_721,N_357);
nor U438 (N_438,In_490,N_262);
or U439 (N_439,N_399,N_110);
nor U440 (N_440,N_337,N_202);
nand U441 (N_441,N_331,N_332);
nand U442 (N_442,N_390,N_224);
and U443 (N_443,N_285,In_116);
nand U444 (N_444,In_334,N_61);
nor U445 (N_445,N_316,N_281);
nor U446 (N_446,N_334,N_360);
nor U447 (N_447,N_229,N_49);
or U448 (N_448,N_361,In_602);
nand U449 (N_449,N_243,In_49);
and U450 (N_450,N_265,In_63);
or U451 (N_451,In_748,N_294);
or U452 (N_452,N_370,N_225);
or U453 (N_453,N_340,N_179);
or U454 (N_454,In_670,N_62);
nor U455 (N_455,N_286,In_711);
nand U456 (N_456,N_397,N_230);
nor U457 (N_457,In_539,In_393);
nor U458 (N_458,In_426,N_379);
and U459 (N_459,N_382,N_227);
nand U460 (N_460,N_306,In_208);
or U461 (N_461,N_90,N_283);
or U462 (N_462,N_259,In_575);
or U463 (N_463,N_312,N_292);
or U464 (N_464,N_256,In_315);
nor U465 (N_465,N_161,N_182);
or U466 (N_466,In_349,N_367);
xnor U467 (N_467,In_640,N_137);
nand U468 (N_468,N_127,N_266);
or U469 (N_469,N_107,N_233);
nor U470 (N_470,In_509,In_523);
and U471 (N_471,N_232,N_33);
nor U472 (N_472,In_282,N_374);
nor U473 (N_473,N_237,N_214);
nand U474 (N_474,N_387,N_322);
and U475 (N_475,N_336,In_427);
or U476 (N_476,In_388,N_315);
nor U477 (N_477,In_668,N_385);
and U478 (N_478,In_61,N_275);
nor U479 (N_479,N_278,N_140);
nor U480 (N_480,N_356,N_353);
nand U481 (N_481,In_521,N_338);
nand U482 (N_482,In_710,In_603);
nor U483 (N_483,N_341,N_271);
nor U484 (N_484,N_261,In_518);
nand U485 (N_485,N_248,N_378);
nor U486 (N_486,N_273,In_210);
or U487 (N_487,In_628,N_279);
nand U488 (N_488,N_267,In_92);
nand U489 (N_489,N_207,N_260);
or U490 (N_490,N_171,In_611);
xor U491 (N_491,In_332,N_200);
nor U492 (N_492,N_366,N_359);
nand U493 (N_493,N_219,N_310);
nand U494 (N_494,N_371,N_304);
and U495 (N_495,In_31,N_342);
nand U496 (N_496,N_314,N_234);
or U497 (N_497,N_87,N_287);
and U498 (N_498,In_220,N_289);
nand U499 (N_499,N_239,N_269);
and U500 (N_500,N_391,N_231);
or U501 (N_501,In_395,N_303);
and U502 (N_502,N_201,In_333);
nor U503 (N_503,N_311,N_320);
nor U504 (N_504,N_350,N_377);
or U505 (N_505,N_31,N_348);
nand U506 (N_506,N_34,In_27);
or U507 (N_507,N_349,N_321);
nor U508 (N_508,In_153,In_720);
nor U509 (N_509,N_67,N_264);
nand U510 (N_510,N_1,N_209);
and U511 (N_511,In_238,N_319);
nor U512 (N_512,N_263,N_344);
nand U513 (N_513,N_395,In_65);
nand U514 (N_514,N_368,In_664);
nor U515 (N_515,N_288,In_414);
and U516 (N_516,N_114,N_309);
or U517 (N_517,N_301,In_621);
and U518 (N_518,N_352,N_392);
and U519 (N_519,N_346,N_324);
nand U520 (N_520,N_375,N_158);
or U521 (N_521,N_282,N_318);
or U522 (N_522,In_667,N_343);
nand U523 (N_523,N_362,N_258);
nor U524 (N_524,In_212,N_381);
nor U525 (N_525,In_78,In_301);
nand U526 (N_526,N_25,N_299);
or U527 (N_527,N_373,N_284);
nand U528 (N_528,N_218,In_318);
nor U529 (N_529,In_154,N_398);
or U530 (N_530,N_270,N_133);
or U531 (N_531,N_236,N_251);
nor U532 (N_532,N_235,N_19);
nor U533 (N_533,In_215,In_722);
and U534 (N_534,N_213,N_253);
and U535 (N_535,In_128,N_3);
and U536 (N_536,In_581,N_244);
or U537 (N_537,N_296,In_423);
or U538 (N_538,N_206,N_242);
nor U539 (N_539,In_604,N_313);
nand U540 (N_540,N_226,N_386);
nor U541 (N_541,N_383,N_39);
or U542 (N_542,In_240,N_217);
and U543 (N_543,N_276,N_335);
nor U544 (N_544,N_238,N_208);
and U545 (N_545,In_106,N_394);
nand U546 (N_546,In_417,N_393);
nand U547 (N_547,In_715,In_543);
or U548 (N_548,In_653,In_40);
nand U549 (N_549,In_487,In_104);
and U550 (N_550,N_249,N_245);
nand U551 (N_551,In_438,N_328);
or U552 (N_552,N_250,N_96);
nand U553 (N_553,In_97,N_293);
nand U554 (N_554,In_95,N_216);
and U555 (N_555,N_128,N_146);
nand U556 (N_556,N_199,N_307);
or U557 (N_557,N_7,N_240);
nor U558 (N_558,In_728,N_376);
nor U559 (N_559,In_177,In_638);
and U560 (N_560,N_247,N_5);
and U561 (N_561,N_257,In_601);
or U562 (N_562,N_222,N_380);
nor U563 (N_563,N_252,N_223);
and U564 (N_564,N_325,N_277);
nor U565 (N_565,N_330,N_13);
and U566 (N_566,N_339,N_53);
and U567 (N_567,N_254,N_66);
or U568 (N_568,N_297,N_28);
nand U569 (N_569,N_388,N_364);
nor U570 (N_570,N_384,In_205);
nand U571 (N_571,N_389,N_300);
nor U572 (N_572,N_329,N_396);
or U573 (N_573,N_308,N_317);
or U574 (N_574,N_351,N_241);
and U575 (N_575,N_369,N_49);
or U576 (N_576,N_41,N_351);
and U577 (N_577,N_327,N_284);
nand U578 (N_578,N_376,N_234);
and U579 (N_579,N_245,N_247);
nor U580 (N_580,In_3,N_387);
or U581 (N_581,N_306,In_575);
nor U582 (N_582,N_365,In_417);
or U583 (N_583,N_340,In_638);
nor U584 (N_584,N_350,In_217);
nand U585 (N_585,In_318,N_262);
nor U586 (N_586,N_238,In_282);
nor U587 (N_587,N_13,N_371);
and U588 (N_588,N_232,In_521);
and U589 (N_589,N_347,N_337);
or U590 (N_590,In_490,In_715);
nor U591 (N_591,N_338,In_200);
and U592 (N_592,N_233,N_26);
nor U593 (N_593,N_110,N_338);
and U594 (N_594,N_53,N_291);
and U595 (N_595,N_379,In_575);
nor U596 (N_596,In_95,In_417);
nor U597 (N_597,N_264,N_305);
nand U598 (N_598,In_653,In_611);
or U599 (N_599,N_233,N_267);
and U600 (N_600,N_458,N_558);
nand U601 (N_601,N_454,N_514);
and U602 (N_602,N_466,N_513);
nand U603 (N_603,N_547,N_530);
or U604 (N_604,N_515,N_533);
nand U605 (N_605,N_542,N_437);
or U606 (N_606,N_519,N_512);
nor U607 (N_607,N_476,N_587);
nand U608 (N_608,N_550,N_579);
nand U609 (N_609,N_598,N_420);
nand U610 (N_610,N_589,N_505);
nor U611 (N_611,N_539,N_578);
nand U612 (N_612,N_583,N_557);
or U613 (N_613,N_592,N_448);
and U614 (N_614,N_510,N_534);
nor U615 (N_615,N_503,N_551);
nor U616 (N_616,N_481,N_541);
and U617 (N_617,N_411,N_544);
nand U618 (N_618,N_426,N_450);
and U619 (N_619,N_455,N_418);
or U620 (N_620,N_472,N_482);
nor U621 (N_621,N_574,N_507);
nand U622 (N_622,N_561,N_500);
xnor U623 (N_623,N_444,N_469);
nor U624 (N_624,N_459,N_492);
or U625 (N_625,N_400,N_532);
or U626 (N_626,N_517,N_494);
nand U627 (N_627,N_453,N_438);
or U628 (N_628,N_461,N_549);
or U629 (N_629,N_478,N_475);
or U630 (N_630,N_566,N_595);
nor U631 (N_631,N_498,N_594);
nand U632 (N_632,N_597,N_467);
or U633 (N_633,N_456,N_548);
nor U634 (N_634,N_483,N_405);
nand U635 (N_635,N_406,N_423);
or U636 (N_636,N_591,N_447);
nand U637 (N_637,N_559,N_402);
nor U638 (N_638,N_429,N_511);
and U639 (N_639,N_445,N_485);
nand U640 (N_640,N_535,N_556);
nor U641 (N_641,N_428,N_486);
or U642 (N_642,N_424,N_401);
nand U643 (N_643,N_590,N_462);
or U644 (N_644,N_442,N_520);
nor U645 (N_645,N_573,N_470);
nand U646 (N_646,N_497,N_523);
or U647 (N_647,N_477,N_493);
nor U648 (N_648,N_540,N_495);
and U649 (N_649,N_436,N_528);
and U650 (N_650,N_584,N_451);
nor U651 (N_651,N_571,N_479);
and U652 (N_652,N_435,N_412);
nand U653 (N_653,N_553,N_552);
or U654 (N_654,N_414,N_518);
or U655 (N_655,N_572,N_487);
nand U656 (N_656,N_516,N_554);
nor U657 (N_657,N_570,N_489);
nor U658 (N_658,N_521,N_567);
and U659 (N_659,N_506,N_427);
nor U660 (N_660,N_504,N_588);
nor U661 (N_661,N_501,N_499);
nand U662 (N_662,N_460,N_491);
or U663 (N_663,N_413,N_465);
and U664 (N_664,N_508,N_522);
nand U665 (N_665,N_509,N_490);
or U666 (N_666,N_471,N_409);
or U667 (N_667,N_526,N_408);
and U668 (N_668,N_431,N_543);
and U669 (N_669,N_531,N_582);
nor U670 (N_670,N_449,N_546);
and U671 (N_671,N_564,N_586);
and U672 (N_672,N_527,N_581);
nand U673 (N_673,N_425,N_502);
nor U674 (N_674,N_457,N_410);
nor U675 (N_675,N_415,N_430);
and U676 (N_676,N_585,N_575);
or U677 (N_677,N_536,N_403);
nor U678 (N_678,N_496,N_404);
or U679 (N_679,N_443,N_545);
nor U680 (N_680,N_441,N_565);
and U681 (N_681,N_568,N_480);
and U682 (N_682,N_488,N_529);
nor U683 (N_683,N_464,N_577);
or U684 (N_684,N_569,N_421);
nand U685 (N_685,N_432,N_484);
or U686 (N_686,N_434,N_580);
nand U687 (N_687,N_468,N_416);
and U688 (N_688,N_452,N_433);
nor U689 (N_689,N_560,N_555);
or U690 (N_690,N_524,N_537);
nand U691 (N_691,N_562,N_538);
and U692 (N_692,N_417,N_463);
or U693 (N_693,N_596,N_474);
and U694 (N_694,N_599,N_473);
nor U695 (N_695,N_563,N_419);
and U696 (N_696,N_525,N_407);
nand U697 (N_697,N_439,N_422);
nand U698 (N_698,N_576,N_446);
or U699 (N_699,N_593,N_440);
and U700 (N_700,N_585,N_483);
or U701 (N_701,N_469,N_590);
or U702 (N_702,N_524,N_564);
and U703 (N_703,N_417,N_543);
or U704 (N_704,N_460,N_484);
nand U705 (N_705,N_565,N_531);
nand U706 (N_706,N_482,N_459);
and U707 (N_707,N_562,N_488);
nand U708 (N_708,N_451,N_416);
nor U709 (N_709,N_501,N_479);
nand U710 (N_710,N_596,N_576);
nand U711 (N_711,N_559,N_594);
and U712 (N_712,N_580,N_537);
and U713 (N_713,N_457,N_424);
or U714 (N_714,N_485,N_452);
or U715 (N_715,N_422,N_536);
or U716 (N_716,N_420,N_437);
and U717 (N_717,N_422,N_528);
or U718 (N_718,N_493,N_453);
or U719 (N_719,N_534,N_526);
or U720 (N_720,N_518,N_536);
nor U721 (N_721,N_421,N_400);
and U722 (N_722,N_472,N_448);
or U723 (N_723,N_401,N_419);
nand U724 (N_724,N_489,N_599);
nor U725 (N_725,N_566,N_515);
or U726 (N_726,N_571,N_511);
nand U727 (N_727,N_455,N_466);
or U728 (N_728,N_596,N_528);
nand U729 (N_729,N_446,N_545);
and U730 (N_730,N_598,N_446);
xnor U731 (N_731,N_538,N_453);
or U732 (N_732,N_414,N_534);
or U733 (N_733,N_409,N_466);
or U734 (N_734,N_542,N_547);
nor U735 (N_735,N_409,N_461);
and U736 (N_736,N_401,N_562);
nor U737 (N_737,N_456,N_594);
nor U738 (N_738,N_423,N_552);
or U739 (N_739,N_543,N_416);
nor U740 (N_740,N_472,N_435);
nor U741 (N_741,N_597,N_446);
nand U742 (N_742,N_431,N_579);
nand U743 (N_743,N_543,N_551);
and U744 (N_744,N_577,N_563);
and U745 (N_745,N_486,N_410);
nand U746 (N_746,N_444,N_460);
nor U747 (N_747,N_593,N_400);
and U748 (N_748,N_470,N_587);
nor U749 (N_749,N_464,N_598);
and U750 (N_750,N_532,N_521);
nor U751 (N_751,N_502,N_595);
or U752 (N_752,N_452,N_500);
or U753 (N_753,N_527,N_577);
and U754 (N_754,N_540,N_461);
nand U755 (N_755,N_568,N_435);
nand U756 (N_756,N_444,N_576);
nor U757 (N_757,N_439,N_416);
nand U758 (N_758,N_535,N_493);
nand U759 (N_759,N_582,N_454);
and U760 (N_760,N_506,N_576);
nand U761 (N_761,N_530,N_434);
or U762 (N_762,N_448,N_590);
nor U763 (N_763,N_452,N_488);
or U764 (N_764,N_521,N_556);
and U765 (N_765,N_479,N_488);
or U766 (N_766,N_463,N_461);
or U767 (N_767,N_436,N_557);
xnor U768 (N_768,N_520,N_428);
or U769 (N_769,N_490,N_579);
and U770 (N_770,N_591,N_430);
nand U771 (N_771,N_424,N_475);
and U772 (N_772,N_580,N_413);
nor U773 (N_773,N_436,N_572);
and U774 (N_774,N_555,N_591);
and U775 (N_775,N_572,N_527);
nor U776 (N_776,N_525,N_553);
nor U777 (N_777,N_407,N_538);
or U778 (N_778,N_467,N_567);
and U779 (N_779,N_508,N_463);
or U780 (N_780,N_568,N_581);
and U781 (N_781,N_529,N_574);
nor U782 (N_782,N_515,N_438);
nand U783 (N_783,N_493,N_520);
nand U784 (N_784,N_503,N_477);
nand U785 (N_785,N_484,N_472);
nor U786 (N_786,N_540,N_464);
and U787 (N_787,N_519,N_415);
nand U788 (N_788,N_563,N_436);
and U789 (N_789,N_524,N_481);
or U790 (N_790,N_442,N_555);
and U791 (N_791,N_407,N_574);
nand U792 (N_792,N_415,N_405);
nand U793 (N_793,N_494,N_489);
nand U794 (N_794,N_406,N_587);
or U795 (N_795,N_528,N_552);
nor U796 (N_796,N_597,N_449);
nor U797 (N_797,N_588,N_471);
nor U798 (N_798,N_578,N_517);
or U799 (N_799,N_565,N_575);
nand U800 (N_800,N_646,N_797);
nand U801 (N_801,N_723,N_717);
nand U802 (N_802,N_708,N_724);
nor U803 (N_803,N_662,N_697);
nor U804 (N_804,N_771,N_690);
and U805 (N_805,N_714,N_600);
or U806 (N_806,N_700,N_788);
nor U807 (N_807,N_673,N_707);
nand U808 (N_808,N_778,N_683);
xor U809 (N_809,N_718,N_686);
nand U810 (N_810,N_668,N_680);
nand U811 (N_811,N_766,N_740);
and U812 (N_812,N_676,N_765);
or U813 (N_813,N_783,N_713);
and U814 (N_814,N_795,N_688);
and U815 (N_815,N_782,N_609);
or U816 (N_816,N_764,N_637);
and U817 (N_817,N_664,N_726);
nor U818 (N_818,N_616,N_739);
or U819 (N_819,N_663,N_665);
and U820 (N_820,N_635,N_636);
and U821 (N_821,N_709,N_704);
nand U822 (N_822,N_622,N_784);
nor U823 (N_823,N_639,N_674);
and U824 (N_824,N_669,N_602);
or U825 (N_825,N_610,N_672);
xnor U826 (N_826,N_691,N_786);
or U827 (N_827,N_762,N_612);
and U828 (N_828,N_745,N_629);
or U829 (N_829,N_747,N_626);
nor U830 (N_830,N_730,N_710);
nor U831 (N_831,N_684,N_647);
nand U832 (N_832,N_623,N_748);
or U833 (N_833,N_632,N_601);
nor U834 (N_834,N_667,N_706);
or U835 (N_835,N_608,N_794);
nor U836 (N_836,N_759,N_789);
and U837 (N_837,N_792,N_793);
and U838 (N_838,N_634,N_781);
or U839 (N_839,N_722,N_640);
or U840 (N_840,N_638,N_620);
and U841 (N_841,N_692,N_657);
and U842 (N_842,N_627,N_621);
and U843 (N_843,N_751,N_643);
and U844 (N_844,N_744,N_687);
nand U845 (N_845,N_698,N_619);
nor U846 (N_846,N_749,N_611);
nor U847 (N_847,N_753,N_727);
nand U848 (N_848,N_716,N_613);
and U849 (N_849,N_628,N_689);
or U850 (N_850,N_725,N_770);
or U851 (N_851,N_768,N_705);
nand U852 (N_852,N_650,N_605);
nor U853 (N_853,N_696,N_767);
nand U854 (N_854,N_607,N_712);
nor U855 (N_855,N_654,N_735);
and U856 (N_856,N_779,N_617);
nor U857 (N_857,N_791,N_741);
nor U858 (N_858,N_677,N_656);
and U859 (N_859,N_750,N_798);
or U860 (N_860,N_757,N_615);
or U861 (N_861,N_652,N_777);
and U862 (N_862,N_760,N_631);
nand U863 (N_863,N_774,N_695);
nor U864 (N_864,N_670,N_699);
or U865 (N_865,N_701,N_651);
and U866 (N_866,N_679,N_702);
nand U867 (N_867,N_658,N_773);
nand U868 (N_868,N_675,N_728);
nor U869 (N_869,N_681,N_653);
and U870 (N_870,N_763,N_743);
nor U871 (N_871,N_787,N_734);
nand U872 (N_872,N_715,N_761);
or U873 (N_873,N_742,N_796);
nor U874 (N_874,N_671,N_729);
and U875 (N_875,N_703,N_754);
or U876 (N_876,N_746,N_666);
and U877 (N_877,N_625,N_694);
nor U878 (N_878,N_678,N_756);
nor U879 (N_879,N_655,N_769);
or U880 (N_880,N_711,N_721);
or U881 (N_881,N_685,N_630);
nand U882 (N_882,N_645,N_644);
nor U883 (N_883,N_736,N_799);
nor U884 (N_884,N_732,N_641);
nand U885 (N_885,N_682,N_733);
and U886 (N_886,N_752,N_758);
or U887 (N_887,N_780,N_633);
nand U888 (N_888,N_606,N_648);
nand U889 (N_889,N_776,N_772);
nor U890 (N_890,N_693,N_661);
or U891 (N_891,N_775,N_659);
nor U892 (N_892,N_642,N_731);
and U893 (N_893,N_649,N_719);
and U894 (N_894,N_755,N_790);
nor U895 (N_895,N_785,N_738);
and U896 (N_896,N_603,N_604);
nor U897 (N_897,N_660,N_614);
and U898 (N_898,N_618,N_737);
or U899 (N_899,N_720,N_624);
or U900 (N_900,N_758,N_680);
or U901 (N_901,N_670,N_646);
and U902 (N_902,N_614,N_678);
nand U903 (N_903,N_787,N_694);
nor U904 (N_904,N_636,N_634);
nor U905 (N_905,N_649,N_610);
or U906 (N_906,N_651,N_638);
and U907 (N_907,N_739,N_617);
and U908 (N_908,N_631,N_695);
nand U909 (N_909,N_735,N_691);
nor U910 (N_910,N_652,N_672);
nand U911 (N_911,N_627,N_655);
nor U912 (N_912,N_753,N_716);
nand U913 (N_913,N_695,N_649);
nor U914 (N_914,N_718,N_707);
and U915 (N_915,N_617,N_726);
and U916 (N_916,N_677,N_638);
and U917 (N_917,N_778,N_755);
and U918 (N_918,N_740,N_779);
nand U919 (N_919,N_707,N_605);
or U920 (N_920,N_722,N_607);
xor U921 (N_921,N_799,N_660);
or U922 (N_922,N_739,N_789);
or U923 (N_923,N_792,N_646);
nand U924 (N_924,N_742,N_658);
or U925 (N_925,N_620,N_680);
nand U926 (N_926,N_607,N_789);
nor U927 (N_927,N_752,N_729);
nand U928 (N_928,N_721,N_682);
nand U929 (N_929,N_729,N_621);
nand U930 (N_930,N_746,N_676);
and U931 (N_931,N_722,N_626);
and U932 (N_932,N_779,N_668);
or U933 (N_933,N_699,N_642);
and U934 (N_934,N_707,N_666);
nand U935 (N_935,N_777,N_685);
or U936 (N_936,N_602,N_616);
or U937 (N_937,N_613,N_650);
nor U938 (N_938,N_670,N_601);
or U939 (N_939,N_612,N_633);
nand U940 (N_940,N_677,N_715);
or U941 (N_941,N_746,N_658);
or U942 (N_942,N_680,N_609);
nand U943 (N_943,N_636,N_622);
or U944 (N_944,N_757,N_792);
nor U945 (N_945,N_736,N_703);
or U946 (N_946,N_648,N_688);
nor U947 (N_947,N_727,N_742);
nor U948 (N_948,N_645,N_730);
nor U949 (N_949,N_710,N_697);
nand U950 (N_950,N_674,N_664);
nand U951 (N_951,N_671,N_711);
nor U952 (N_952,N_714,N_660);
nor U953 (N_953,N_664,N_668);
nand U954 (N_954,N_691,N_762);
nand U955 (N_955,N_670,N_718);
nor U956 (N_956,N_602,N_780);
and U957 (N_957,N_628,N_679);
nand U958 (N_958,N_757,N_764);
and U959 (N_959,N_795,N_738);
and U960 (N_960,N_621,N_770);
and U961 (N_961,N_766,N_739);
nor U962 (N_962,N_640,N_675);
or U963 (N_963,N_753,N_766);
nor U964 (N_964,N_752,N_689);
or U965 (N_965,N_787,N_735);
nor U966 (N_966,N_757,N_742);
and U967 (N_967,N_693,N_699);
and U968 (N_968,N_673,N_768);
nand U969 (N_969,N_652,N_754);
or U970 (N_970,N_717,N_651);
or U971 (N_971,N_703,N_656);
nor U972 (N_972,N_798,N_769);
nand U973 (N_973,N_730,N_797);
and U974 (N_974,N_620,N_654);
and U975 (N_975,N_686,N_721);
nand U976 (N_976,N_714,N_647);
nor U977 (N_977,N_673,N_677);
nand U978 (N_978,N_649,N_652);
and U979 (N_979,N_622,N_772);
and U980 (N_980,N_617,N_678);
nor U981 (N_981,N_625,N_733);
and U982 (N_982,N_633,N_614);
nor U983 (N_983,N_780,N_628);
nand U984 (N_984,N_662,N_725);
nor U985 (N_985,N_717,N_661);
and U986 (N_986,N_727,N_646);
or U987 (N_987,N_690,N_673);
and U988 (N_988,N_771,N_768);
nor U989 (N_989,N_617,N_612);
nor U990 (N_990,N_701,N_758);
nor U991 (N_991,N_769,N_725);
nor U992 (N_992,N_765,N_702);
or U993 (N_993,N_614,N_625);
or U994 (N_994,N_616,N_638);
or U995 (N_995,N_703,N_753);
or U996 (N_996,N_647,N_671);
and U997 (N_997,N_677,N_613);
and U998 (N_998,N_753,N_761);
nor U999 (N_999,N_635,N_638);
and U1000 (N_1000,N_969,N_801);
xnor U1001 (N_1001,N_944,N_940);
or U1002 (N_1002,N_803,N_972);
and U1003 (N_1003,N_996,N_974);
nand U1004 (N_1004,N_946,N_907);
and U1005 (N_1005,N_800,N_950);
and U1006 (N_1006,N_882,N_982);
and U1007 (N_1007,N_839,N_964);
or U1008 (N_1008,N_920,N_929);
or U1009 (N_1009,N_930,N_966);
nand U1010 (N_1010,N_859,N_881);
and U1011 (N_1011,N_921,N_868);
or U1012 (N_1012,N_909,N_955);
or U1013 (N_1013,N_908,N_885);
nor U1014 (N_1014,N_861,N_802);
and U1015 (N_1015,N_806,N_919);
or U1016 (N_1016,N_928,N_834);
or U1017 (N_1017,N_942,N_915);
and U1018 (N_1018,N_887,N_835);
or U1019 (N_1019,N_865,N_918);
and U1020 (N_1020,N_814,N_849);
or U1021 (N_1021,N_995,N_992);
nand U1022 (N_1022,N_979,N_903);
nor U1023 (N_1023,N_988,N_821);
or U1024 (N_1024,N_949,N_855);
and U1025 (N_1025,N_847,N_961);
nor U1026 (N_1026,N_923,N_937);
or U1027 (N_1027,N_963,N_986);
nor U1028 (N_1028,N_926,N_945);
and U1029 (N_1029,N_917,N_993);
or U1030 (N_1030,N_958,N_876);
or U1031 (N_1031,N_828,N_846);
or U1032 (N_1032,N_867,N_932);
or U1033 (N_1033,N_805,N_850);
nand U1034 (N_1034,N_904,N_819);
or U1035 (N_1035,N_948,N_845);
and U1036 (N_1036,N_875,N_816);
and U1037 (N_1037,N_895,N_911);
nand U1038 (N_1038,N_981,N_910);
and U1039 (N_1039,N_874,N_977);
nand U1040 (N_1040,N_815,N_894);
or U1041 (N_1041,N_884,N_990);
nor U1042 (N_1042,N_943,N_860);
nand U1043 (N_1043,N_832,N_858);
or U1044 (N_1044,N_960,N_871);
or U1045 (N_1045,N_879,N_991);
or U1046 (N_1046,N_817,N_888);
nor U1047 (N_1047,N_813,N_864);
nor U1048 (N_1048,N_956,N_826);
nand U1049 (N_1049,N_880,N_938);
nor U1050 (N_1050,N_900,N_983);
or U1051 (N_1051,N_878,N_952);
and U1052 (N_1052,N_978,N_939);
nand U1053 (N_1053,N_840,N_954);
and U1054 (N_1054,N_973,N_916);
nand U1055 (N_1055,N_886,N_931);
or U1056 (N_1056,N_820,N_812);
nor U1057 (N_1057,N_844,N_967);
nand U1058 (N_1058,N_866,N_934);
and U1059 (N_1059,N_851,N_872);
nand U1060 (N_1060,N_856,N_985);
or U1061 (N_1061,N_959,N_975);
and U1062 (N_1062,N_968,N_889);
nor U1063 (N_1063,N_994,N_933);
nor U1064 (N_1064,N_841,N_863);
or U1065 (N_1065,N_925,N_810);
nor U1066 (N_1066,N_902,N_953);
nand U1067 (N_1067,N_825,N_924);
nand U1068 (N_1068,N_852,N_873);
nor U1069 (N_1069,N_890,N_842);
and U1070 (N_1070,N_896,N_989);
or U1071 (N_1071,N_898,N_935);
or U1072 (N_1072,N_807,N_824);
or U1073 (N_1073,N_857,N_854);
nand U1074 (N_1074,N_905,N_912);
nor U1075 (N_1075,N_970,N_999);
nor U1076 (N_1076,N_836,N_901);
or U1077 (N_1077,N_914,N_936);
nor U1078 (N_1078,N_962,N_899);
nor U1079 (N_1079,N_843,N_883);
nand U1080 (N_1080,N_811,N_913);
nor U1081 (N_1081,N_922,N_829);
or U1082 (N_1082,N_941,N_997);
nor U1083 (N_1083,N_893,N_831);
or U1084 (N_1084,N_951,N_869);
or U1085 (N_1085,N_891,N_980);
or U1086 (N_1086,N_804,N_827);
or U1087 (N_1087,N_862,N_971);
and U1088 (N_1088,N_837,N_853);
and U1089 (N_1089,N_830,N_897);
or U1090 (N_1090,N_984,N_822);
or U1091 (N_1091,N_987,N_965);
or U1092 (N_1092,N_998,N_906);
xor U1093 (N_1093,N_809,N_818);
nor U1094 (N_1094,N_877,N_947);
and U1095 (N_1095,N_808,N_870);
nor U1096 (N_1096,N_976,N_927);
and U1097 (N_1097,N_957,N_823);
or U1098 (N_1098,N_833,N_838);
nand U1099 (N_1099,N_848,N_892);
and U1100 (N_1100,N_903,N_906);
or U1101 (N_1101,N_924,N_812);
and U1102 (N_1102,N_977,N_812);
nand U1103 (N_1103,N_838,N_823);
and U1104 (N_1104,N_892,N_958);
or U1105 (N_1105,N_981,N_876);
nor U1106 (N_1106,N_811,N_865);
nor U1107 (N_1107,N_978,N_858);
nand U1108 (N_1108,N_998,N_979);
nand U1109 (N_1109,N_977,N_861);
nor U1110 (N_1110,N_997,N_818);
or U1111 (N_1111,N_902,N_956);
nor U1112 (N_1112,N_912,N_985);
nor U1113 (N_1113,N_816,N_990);
nor U1114 (N_1114,N_848,N_840);
or U1115 (N_1115,N_885,N_956);
nand U1116 (N_1116,N_976,N_995);
and U1117 (N_1117,N_817,N_826);
or U1118 (N_1118,N_929,N_915);
nand U1119 (N_1119,N_995,N_818);
nor U1120 (N_1120,N_921,N_876);
nor U1121 (N_1121,N_970,N_841);
nand U1122 (N_1122,N_996,N_915);
nand U1123 (N_1123,N_977,N_987);
and U1124 (N_1124,N_929,N_844);
or U1125 (N_1125,N_844,N_966);
and U1126 (N_1126,N_804,N_964);
nand U1127 (N_1127,N_997,N_926);
nand U1128 (N_1128,N_966,N_897);
and U1129 (N_1129,N_815,N_956);
or U1130 (N_1130,N_959,N_803);
or U1131 (N_1131,N_943,N_894);
and U1132 (N_1132,N_803,N_940);
nand U1133 (N_1133,N_878,N_867);
or U1134 (N_1134,N_863,N_973);
nor U1135 (N_1135,N_896,N_946);
or U1136 (N_1136,N_922,N_927);
nor U1137 (N_1137,N_851,N_918);
nand U1138 (N_1138,N_835,N_911);
nor U1139 (N_1139,N_857,N_868);
nor U1140 (N_1140,N_807,N_948);
nor U1141 (N_1141,N_952,N_831);
nor U1142 (N_1142,N_899,N_978);
nand U1143 (N_1143,N_889,N_859);
nor U1144 (N_1144,N_829,N_962);
and U1145 (N_1145,N_985,N_983);
or U1146 (N_1146,N_843,N_881);
and U1147 (N_1147,N_885,N_972);
or U1148 (N_1148,N_812,N_874);
nor U1149 (N_1149,N_878,N_965);
nor U1150 (N_1150,N_970,N_920);
nand U1151 (N_1151,N_926,N_998);
or U1152 (N_1152,N_927,N_874);
nand U1153 (N_1153,N_862,N_887);
nand U1154 (N_1154,N_986,N_938);
nor U1155 (N_1155,N_834,N_855);
nand U1156 (N_1156,N_960,N_990);
nor U1157 (N_1157,N_843,N_905);
or U1158 (N_1158,N_865,N_909);
and U1159 (N_1159,N_827,N_886);
and U1160 (N_1160,N_882,N_983);
or U1161 (N_1161,N_800,N_996);
nor U1162 (N_1162,N_860,N_930);
nand U1163 (N_1163,N_966,N_927);
or U1164 (N_1164,N_982,N_986);
or U1165 (N_1165,N_854,N_995);
or U1166 (N_1166,N_858,N_939);
nor U1167 (N_1167,N_958,N_917);
nand U1168 (N_1168,N_981,N_872);
nor U1169 (N_1169,N_805,N_811);
nor U1170 (N_1170,N_853,N_859);
or U1171 (N_1171,N_927,N_994);
nand U1172 (N_1172,N_841,N_899);
nand U1173 (N_1173,N_843,N_973);
and U1174 (N_1174,N_884,N_905);
nand U1175 (N_1175,N_996,N_945);
or U1176 (N_1176,N_976,N_843);
nor U1177 (N_1177,N_836,N_833);
and U1178 (N_1178,N_977,N_899);
nor U1179 (N_1179,N_876,N_945);
nand U1180 (N_1180,N_999,N_842);
nand U1181 (N_1181,N_948,N_873);
or U1182 (N_1182,N_845,N_872);
and U1183 (N_1183,N_988,N_898);
nor U1184 (N_1184,N_909,N_968);
nor U1185 (N_1185,N_875,N_874);
nor U1186 (N_1186,N_839,N_814);
or U1187 (N_1187,N_973,N_932);
nand U1188 (N_1188,N_890,N_906);
and U1189 (N_1189,N_955,N_985);
nand U1190 (N_1190,N_901,N_841);
nor U1191 (N_1191,N_907,N_970);
nor U1192 (N_1192,N_984,N_823);
or U1193 (N_1193,N_921,N_849);
nand U1194 (N_1194,N_859,N_927);
nand U1195 (N_1195,N_908,N_916);
nor U1196 (N_1196,N_908,N_998);
nor U1197 (N_1197,N_832,N_955);
and U1198 (N_1198,N_960,N_884);
and U1199 (N_1199,N_933,N_894);
nand U1200 (N_1200,N_1199,N_1047);
and U1201 (N_1201,N_1167,N_1198);
nand U1202 (N_1202,N_1179,N_1101);
nand U1203 (N_1203,N_1193,N_1010);
and U1204 (N_1204,N_1061,N_1190);
and U1205 (N_1205,N_1065,N_1079);
and U1206 (N_1206,N_1104,N_1036);
nor U1207 (N_1207,N_1168,N_1161);
nor U1208 (N_1208,N_1176,N_1169);
nand U1209 (N_1209,N_1068,N_1125);
nand U1210 (N_1210,N_1120,N_1052);
nand U1211 (N_1211,N_1038,N_1042);
nor U1212 (N_1212,N_1128,N_1013);
nor U1213 (N_1213,N_1126,N_1160);
nor U1214 (N_1214,N_1019,N_1124);
xnor U1215 (N_1215,N_1005,N_1002);
nor U1216 (N_1216,N_1114,N_1166);
nand U1217 (N_1217,N_1064,N_1162);
nand U1218 (N_1218,N_1075,N_1037);
nand U1219 (N_1219,N_1043,N_1122);
nor U1220 (N_1220,N_1194,N_1041);
nand U1221 (N_1221,N_1146,N_1089);
nand U1222 (N_1222,N_1118,N_1185);
and U1223 (N_1223,N_1099,N_1046);
nor U1224 (N_1224,N_1113,N_1196);
nand U1225 (N_1225,N_1136,N_1096);
nor U1226 (N_1226,N_1082,N_1029);
nor U1227 (N_1227,N_1024,N_1111);
and U1228 (N_1228,N_1195,N_1164);
nand U1229 (N_1229,N_1112,N_1008);
xnor U1230 (N_1230,N_1197,N_1015);
nand U1231 (N_1231,N_1181,N_1135);
and U1232 (N_1232,N_1092,N_1009);
nor U1233 (N_1233,N_1186,N_1063);
nor U1234 (N_1234,N_1060,N_1087);
nand U1235 (N_1235,N_1067,N_1070);
nor U1236 (N_1236,N_1182,N_1007);
nand U1237 (N_1237,N_1172,N_1023);
or U1238 (N_1238,N_1192,N_1083);
and U1239 (N_1239,N_1033,N_1137);
and U1240 (N_1240,N_1115,N_1030);
and U1241 (N_1241,N_1027,N_1129);
and U1242 (N_1242,N_1094,N_1093);
and U1243 (N_1243,N_1156,N_1003);
nor U1244 (N_1244,N_1022,N_1175);
and U1245 (N_1245,N_1178,N_1119);
nor U1246 (N_1246,N_1151,N_1116);
nor U1247 (N_1247,N_1088,N_1016);
and U1248 (N_1248,N_1091,N_1143);
nor U1249 (N_1249,N_1012,N_1157);
and U1250 (N_1250,N_1098,N_1174);
or U1251 (N_1251,N_1090,N_1085);
or U1252 (N_1252,N_1057,N_1084);
nand U1253 (N_1253,N_1105,N_1158);
and U1254 (N_1254,N_1055,N_1148);
or U1255 (N_1255,N_1153,N_1140);
nand U1256 (N_1256,N_1159,N_1017);
nor U1257 (N_1257,N_1031,N_1004);
nor U1258 (N_1258,N_1028,N_1142);
nand U1259 (N_1259,N_1134,N_1001);
and U1260 (N_1260,N_1049,N_1006);
nand U1261 (N_1261,N_1020,N_1138);
nand U1262 (N_1262,N_1173,N_1170);
or U1263 (N_1263,N_1149,N_1051);
or U1264 (N_1264,N_1184,N_1107);
nor U1265 (N_1265,N_1177,N_1141);
and U1266 (N_1266,N_1066,N_1011);
nand U1267 (N_1267,N_1133,N_1165);
nand U1268 (N_1268,N_1180,N_1058);
or U1269 (N_1269,N_1102,N_1062);
nor U1270 (N_1270,N_1080,N_1072);
nand U1271 (N_1271,N_1018,N_1077);
nor U1272 (N_1272,N_1097,N_1069);
and U1273 (N_1273,N_1189,N_1191);
nand U1274 (N_1274,N_1152,N_1034);
and U1275 (N_1275,N_1144,N_1000);
or U1276 (N_1276,N_1073,N_1188);
or U1277 (N_1277,N_1127,N_1053);
nor U1278 (N_1278,N_1139,N_1130);
nor U1279 (N_1279,N_1050,N_1095);
nand U1280 (N_1280,N_1048,N_1039);
and U1281 (N_1281,N_1117,N_1076);
or U1282 (N_1282,N_1154,N_1132);
nand U1283 (N_1283,N_1014,N_1187);
and U1284 (N_1284,N_1155,N_1032);
or U1285 (N_1285,N_1171,N_1145);
xor U1286 (N_1286,N_1110,N_1045);
nor U1287 (N_1287,N_1163,N_1131);
nor U1288 (N_1288,N_1044,N_1040);
nor U1289 (N_1289,N_1035,N_1108);
nor U1290 (N_1290,N_1059,N_1103);
or U1291 (N_1291,N_1026,N_1081);
nor U1292 (N_1292,N_1056,N_1121);
nand U1293 (N_1293,N_1086,N_1078);
and U1294 (N_1294,N_1054,N_1183);
nor U1295 (N_1295,N_1109,N_1100);
or U1296 (N_1296,N_1025,N_1123);
nand U1297 (N_1297,N_1074,N_1106);
nand U1298 (N_1298,N_1150,N_1021);
nand U1299 (N_1299,N_1071,N_1147);
nand U1300 (N_1300,N_1119,N_1061);
nand U1301 (N_1301,N_1194,N_1017);
nor U1302 (N_1302,N_1127,N_1123);
nor U1303 (N_1303,N_1000,N_1016);
nor U1304 (N_1304,N_1031,N_1144);
or U1305 (N_1305,N_1158,N_1125);
or U1306 (N_1306,N_1041,N_1102);
nand U1307 (N_1307,N_1146,N_1145);
and U1308 (N_1308,N_1095,N_1037);
and U1309 (N_1309,N_1154,N_1168);
or U1310 (N_1310,N_1038,N_1018);
nand U1311 (N_1311,N_1125,N_1011);
nor U1312 (N_1312,N_1074,N_1048);
nand U1313 (N_1313,N_1097,N_1171);
and U1314 (N_1314,N_1021,N_1125);
or U1315 (N_1315,N_1040,N_1072);
xor U1316 (N_1316,N_1163,N_1140);
and U1317 (N_1317,N_1154,N_1010);
and U1318 (N_1318,N_1196,N_1173);
and U1319 (N_1319,N_1079,N_1026);
nand U1320 (N_1320,N_1025,N_1017);
nand U1321 (N_1321,N_1071,N_1164);
nand U1322 (N_1322,N_1086,N_1104);
nand U1323 (N_1323,N_1118,N_1155);
or U1324 (N_1324,N_1061,N_1039);
or U1325 (N_1325,N_1183,N_1186);
or U1326 (N_1326,N_1111,N_1023);
and U1327 (N_1327,N_1024,N_1169);
or U1328 (N_1328,N_1009,N_1165);
or U1329 (N_1329,N_1178,N_1052);
and U1330 (N_1330,N_1118,N_1109);
and U1331 (N_1331,N_1030,N_1133);
nor U1332 (N_1332,N_1175,N_1011);
and U1333 (N_1333,N_1128,N_1166);
or U1334 (N_1334,N_1017,N_1128);
or U1335 (N_1335,N_1159,N_1090);
nand U1336 (N_1336,N_1012,N_1070);
or U1337 (N_1337,N_1156,N_1108);
nand U1338 (N_1338,N_1050,N_1084);
xnor U1339 (N_1339,N_1046,N_1032);
nand U1340 (N_1340,N_1157,N_1075);
and U1341 (N_1341,N_1018,N_1168);
and U1342 (N_1342,N_1037,N_1101);
or U1343 (N_1343,N_1122,N_1138);
nor U1344 (N_1344,N_1124,N_1162);
or U1345 (N_1345,N_1131,N_1091);
nand U1346 (N_1346,N_1027,N_1022);
and U1347 (N_1347,N_1009,N_1100);
or U1348 (N_1348,N_1080,N_1103);
xor U1349 (N_1349,N_1024,N_1011);
and U1350 (N_1350,N_1140,N_1026);
or U1351 (N_1351,N_1048,N_1128);
or U1352 (N_1352,N_1116,N_1082);
or U1353 (N_1353,N_1030,N_1056);
and U1354 (N_1354,N_1176,N_1092);
and U1355 (N_1355,N_1075,N_1187);
or U1356 (N_1356,N_1098,N_1130);
nor U1357 (N_1357,N_1178,N_1125);
and U1358 (N_1358,N_1170,N_1174);
nand U1359 (N_1359,N_1091,N_1118);
nor U1360 (N_1360,N_1044,N_1008);
nand U1361 (N_1361,N_1101,N_1159);
and U1362 (N_1362,N_1109,N_1056);
or U1363 (N_1363,N_1143,N_1097);
nand U1364 (N_1364,N_1017,N_1003);
nor U1365 (N_1365,N_1037,N_1013);
nand U1366 (N_1366,N_1097,N_1158);
and U1367 (N_1367,N_1044,N_1158);
nor U1368 (N_1368,N_1151,N_1119);
or U1369 (N_1369,N_1022,N_1090);
nand U1370 (N_1370,N_1188,N_1096);
nand U1371 (N_1371,N_1118,N_1140);
nand U1372 (N_1372,N_1152,N_1118);
or U1373 (N_1373,N_1125,N_1160);
nor U1374 (N_1374,N_1027,N_1199);
nor U1375 (N_1375,N_1081,N_1162);
nand U1376 (N_1376,N_1133,N_1004);
or U1377 (N_1377,N_1082,N_1008);
and U1378 (N_1378,N_1167,N_1083);
and U1379 (N_1379,N_1184,N_1150);
nand U1380 (N_1380,N_1183,N_1002);
and U1381 (N_1381,N_1023,N_1057);
or U1382 (N_1382,N_1187,N_1048);
nor U1383 (N_1383,N_1012,N_1072);
or U1384 (N_1384,N_1075,N_1042);
and U1385 (N_1385,N_1103,N_1114);
nor U1386 (N_1386,N_1098,N_1053);
and U1387 (N_1387,N_1005,N_1038);
or U1388 (N_1388,N_1187,N_1041);
or U1389 (N_1389,N_1160,N_1024);
or U1390 (N_1390,N_1087,N_1066);
nand U1391 (N_1391,N_1151,N_1104);
nor U1392 (N_1392,N_1139,N_1112);
nor U1393 (N_1393,N_1101,N_1087);
nand U1394 (N_1394,N_1135,N_1013);
nor U1395 (N_1395,N_1031,N_1095);
nand U1396 (N_1396,N_1126,N_1116);
and U1397 (N_1397,N_1043,N_1129);
and U1398 (N_1398,N_1121,N_1032);
and U1399 (N_1399,N_1063,N_1059);
or U1400 (N_1400,N_1339,N_1323);
and U1401 (N_1401,N_1322,N_1251);
or U1402 (N_1402,N_1319,N_1369);
and U1403 (N_1403,N_1346,N_1201);
and U1404 (N_1404,N_1310,N_1357);
and U1405 (N_1405,N_1326,N_1358);
nor U1406 (N_1406,N_1291,N_1380);
nand U1407 (N_1407,N_1397,N_1315);
nor U1408 (N_1408,N_1231,N_1209);
nor U1409 (N_1409,N_1305,N_1250);
nor U1410 (N_1410,N_1354,N_1371);
and U1411 (N_1411,N_1298,N_1236);
nor U1412 (N_1412,N_1279,N_1327);
nor U1413 (N_1413,N_1259,N_1216);
and U1414 (N_1414,N_1265,N_1263);
nor U1415 (N_1415,N_1246,N_1233);
or U1416 (N_1416,N_1329,N_1321);
or U1417 (N_1417,N_1395,N_1242);
nand U1418 (N_1418,N_1227,N_1278);
and U1419 (N_1419,N_1208,N_1235);
or U1420 (N_1420,N_1283,N_1223);
nand U1421 (N_1421,N_1306,N_1363);
nor U1422 (N_1422,N_1388,N_1337);
nand U1423 (N_1423,N_1325,N_1301);
or U1424 (N_1424,N_1269,N_1333);
and U1425 (N_1425,N_1360,N_1393);
nor U1426 (N_1426,N_1222,N_1331);
nand U1427 (N_1427,N_1232,N_1320);
or U1428 (N_1428,N_1332,N_1334);
nand U1429 (N_1429,N_1200,N_1308);
nor U1430 (N_1430,N_1302,N_1290);
or U1431 (N_1431,N_1318,N_1330);
nand U1432 (N_1432,N_1328,N_1373);
nor U1433 (N_1433,N_1244,N_1273);
or U1434 (N_1434,N_1226,N_1218);
or U1435 (N_1435,N_1314,N_1309);
nor U1436 (N_1436,N_1387,N_1378);
and U1437 (N_1437,N_1258,N_1353);
or U1438 (N_1438,N_1351,N_1381);
nand U1439 (N_1439,N_1238,N_1254);
nor U1440 (N_1440,N_1268,N_1215);
or U1441 (N_1441,N_1344,N_1262);
nor U1442 (N_1442,N_1287,N_1205);
nor U1443 (N_1443,N_1221,N_1288);
nor U1444 (N_1444,N_1240,N_1347);
nand U1445 (N_1445,N_1229,N_1335);
or U1446 (N_1446,N_1261,N_1342);
nor U1447 (N_1447,N_1389,N_1355);
and U1448 (N_1448,N_1361,N_1230);
and U1449 (N_1449,N_1376,N_1362);
nand U1450 (N_1450,N_1202,N_1257);
and U1451 (N_1451,N_1364,N_1300);
and U1452 (N_1452,N_1228,N_1270);
or U1453 (N_1453,N_1281,N_1324);
nand U1454 (N_1454,N_1392,N_1260);
nand U1455 (N_1455,N_1374,N_1255);
nor U1456 (N_1456,N_1352,N_1276);
nand U1457 (N_1457,N_1390,N_1264);
and U1458 (N_1458,N_1241,N_1267);
or U1459 (N_1459,N_1266,N_1292);
nor U1460 (N_1460,N_1365,N_1366);
nand U1461 (N_1461,N_1399,N_1316);
nor U1462 (N_1462,N_1370,N_1275);
nand U1463 (N_1463,N_1396,N_1285);
nor U1464 (N_1464,N_1271,N_1237);
nor U1465 (N_1465,N_1282,N_1304);
nor U1466 (N_1466,N_1296,N_1312);
nand U1467 (N_1467,N_1252,N_1217);
nand U1468 (N_1468,N_1204,N_1343);
or U1469 (N_1469,N_1256,N_1207);
nand U1470 (N_1470,N_1398,N_1224);
and U1471 (N_1471,N_1356,N_1313);
nand U1472 (N_1472,N_1299,N_1294);
or U1473 (N_1473,N_1372,N_1280);
or U1474 (N_1474,N_1211,N_1338);
or U1475 (N_1475,N_1206,N_1317);
nand U1476 (N_1476,N_1350,N_1225);
or U1477 (N_1477,N_1248,N_1394);
xnor U1478 (N_1478,N_1214,N_1386);
nand U1479 (N_1479,N_1272,N_1289);
nand U1480 (N_1480,N_1213,N_1293);
and U1481 (N_1481,N_1249,N_1349);
nor U1482 (N_1482,N_1297,N_1375);
nand U1483 (N_1483,N_1307,N_1212);
and U1484 (N_1484,N_1384,N_1277);
nand U1485 (N_1485,N_1253,N_1311);
nand U1486 (N_1486,N_1367,N_1336);
nand U1487 (N_1487,N_1219,N_1382);
or U1488 (N_1488,N_1385,N_1379);
and U1489 (N_1489,N_1243,N_1377);
nor U1490 (N_1490,N_1247,N_1359);
nor U1491 (N_1491,N_1345,N_1341);
or U1492 (N_1492,N_1303,N_1286);
or U1493 (N_1493,N_1210,N_1391);
nand U1494 (N_1494,N_1368,N_1348);
nand U1495 (N_1495,N_1295,N_1274);
and U1496 (N_1496,N_1284,N_1340);
nand U1497 (N_1497,N_1234,N_1220);
or U1498 (N_1498,N_1239,N_1383);
or U1499 (N_1499,N_1245,N_1203);
nor U1500 (N_1500,N_1308,N_1278);
or U1501 (N_1501,N_1337,N_1251);
nand U1502 (N_1502,N_1207,N_1366);
or U1503 (N_1503,N_1372,N_1315);
or U1504 (N_1504,N_1292,N_1240);
and U1505 (N_1505,N_1346,N_1387);
nand U1506 (N_1506,N_1208,N_1311);
nor U1507 (N_1507,N_1342,N_1244);
nor U1508 (N_1508,N_1312,N_1298);
nand U1509 (N_1509,N_1214,N_1366);
nand U1510 (N_1510,N_1265,N_1215);
nand U1511 (N_1511,N_1204,N_1334);
nand U1512 (N_1512,N_1206,N_1230);
nand U1513 (N_1513,N_1392,N_1243);
nand U1514 (N_1514,N_1379,N_1399);
nor U1515 (N_1515,N_1320,N_1339);
nor U1516 (N_1516,N_1396,N_1309);
or U1517 (N_1517,N_1301,N_1258);
or U1518 (N_1518,N_1375,N_1211);
nand U1519 (N_1519,N_1214,N_1361);
nor U1520 (N_1520,N_1214,N_1354);
nand U1521 (N_1521,N_1390,N_1347);
and U1522 (N_1522,N_1334,N_1233);
nor U1523 (N_1523,N_1361,N_1390);
nor U1524 (N_1524,N_1367,N_1230);
nand U1525 (N_1525,N_1250,N_1397);
nand U1526 (N_1526,N_1231,N_1281);
and U1527 (N_1527,N_1318,N_1376);
nand U1528 (N_1528,N_1216,N_1324);
and U1529 (N_1529,N_1238,N_1347);
nor U1530 (N_1530,N_1374,N_1393);
nor U1531 (N_1531,N_1316,N_1362);
nand U1532 (N_1532,N_1337,N_1347);
nor U1533 (N_1533,N_1232,N_1330);
nand U1534 (N_1534,N_1340,N_1253);
nand U1535 (N_1535,N_1265,N_1354);
or U1536 (N_1536,N_1303,N_1347);
nor U1537 (N_1537,N_1281,N_1329);
and U1538 (N_1538,N_1335,N_1311);
nand U1539 (N_1539,N_1273,N_1345);
nor U1540 (N_1540,N_1361,N_1355);
and U1541 (N_1541,N_1245,N_1249);
and U1542 (N_1542,N_1325,N_1376);
or U1543 (N_1543,N_1222,N_1210);
nor U1544 (N_1544,N_1313,N_1288);
xor U1545 (N_1545,N_1204,N_1361);
and U1546 (N_1546,N_1325,N_1394);
nand U1547 (N_1547,N_1382,N_1256);
or U1548 (N_1548,N_1276,N_1257);
nor U1549 (N_1549,N_1243,N_1289);
and U1550 (N_1550,N_1374,N_1380);
and U1551 (N_1551,N_1211,N_1359);
and U1552 (N_1552,N_1321,N_1356);
and U1553 (N_1553,N_1392,N_1372);
or U1554 (N_1554,N_1369,N_1256);
nand U1555 (N_1555,N_1263,N_1258);
and U1556 (N_1556,N_1340,N_1310);
or U1557 (N_1557,N_1341,N_1212);
nor U1558 (N_1558,N_1345,N_1281);
nor U1559 (N_1559,N_1344,N_1216);
and U1560 (N_1560,N_1256,N_1279);
and U1561 (N_1561,N_1259,N_1388);
nor U1562 (N_1562,N_1257,N_1302);
nand U1563 (N_1563,N_1211,N_1393);
or U1564 (N_1564,N_1295,N_1373);
or U1565 (N_1565,N_1370,N_1247);
and U1566 (N_1566,N_1271,N_1254);
nor U1567 (N_1567,N_1392,N_1258);
and U1568 (N_1568,N_1302,N_1262);
and U1569 (N_1569,N_1316,N_1331);
nor U1570 (N_1570,N_1382,N_1372);
nand U1571 (N_1571,N_1257,N_1201);
or U1572 (N_1572,N_1311,N_1210);
or U1573 (N_1573,N_1325,N_1352);
and U1574 (N_1574,N_1370,N_1386);
nand U1575 (N_1575,N_1247,N_1273);
or U1576 (N_1576,N_1222,N_1220);
nor U1577 (N_1577,N_1359,N_1321);
or U1578 (N_1578,N_1217,N_1259);
or U1579 (N_1579,N_1388,N_1256);
or U1580 (N_1580,N_1214,N_1297);
nor U1581 (N_1581,N_1315,N_1385);
nand U1582 (N_1582,N_1383,N_1262);
nand U1583 (N_1583,N_1263,N_1304);
nor U1584 (N_1584,N_1280,N_1204);
or U1585 (N_1585,N_1268,N_1200);
nand U1586 (N_1586,N_1277,N_1317);
or U1587 (N_1587,N_1342,N_1315);
and U1588 (N_1588,N_1350,N_1384);
nand U1589 (N_1589,N_1380,N_1304);
or U1590 (N_1590,N_1270,N_1254);
nand U1591 (N_1591,N_1353,N_1327);
nor U1592 (N_1592,N_1282,N_1339);
nor U1593 (N_1593,N_1228,N_1305);
and U1594 (N_1594,N_1309,N_1307);
nand U1595 (N_1595,N_1341,N_1394);
or U1596 (N_1596,N_1251,N_1303);
nand U1597 (N_1597,N_1330,N_1349);
nor U1598 (N_1598,N_1374,N_1390);
or U1599 (N_1599,N_1225,N_1286);
nand U1600 (N_1600,N_1521,N_1584);
and U1601 (N_1601,N_1543,N_1428);
and U1602 (N_1602,N_1595,N_1539);
nor U1603 (N_1603,N_1557,N_1503);
nor U1604 (N_1604,N_1413,N_1527);
and U1605 (N_1605,N_1476,N_1488);
and U1606 (N_1606,N_1438,N_1401);
nor U1607 (N_1607,N_1496,N_1422);
nor U1608 (N_1608,N_1437,N_1477);
nor U1609 (N_1609,N_1554,N_1571);
nor U1610 (N_1610,N_1450,N_1564);
nand U1611 (N_1611,N_1485,N_1480);
nand U1612 (N_1612,N_1430,N_1525);
xor U1613 (N_1613,N_1563,N_1502);
or U1614 (N_1614,N_1507,N_1403);
and U1615 (N_1615,N_1552,N_1446);
xnor U1616 (N_1616,N_1528,N_1433);
nor U1617 (N_1617,N_1548,N_1458);
or U1618 (N_1618,N_1593,N_1442);
or U1619 (N_1619,N_1558,N_1483);
nand U1620 (N_1620,N_1501,N_1583);
or U1621 (N_1621,N_1547,N_1463);
nor U1622 (N_1622,N_1466,N_1482);
and U1623 (N_1623,N_1471,N_1455);
nand U1624 (N_1624,N_1504,N_1536);
nand U1625 (N_1625,N_1538,N_1551);
and U1626 (N_1626,N_1578,N_1506);
nor U1627 (N_1627,N_1434,N_1461);
nor U1628 (N_1628,N_1582,N_1418);
nand U1629 (N_1629,N_1491,N_1423);
nor U1630 (N_1630,N_1594,N_1499);
and U1631 (N_1631,N_1472,N_1556);
nor U1632 (N_1632,N_1518,N_1549);
nand U1633 (N_1633,N_1432,N_1529);
and U1634 (N_1634,N_1510,N_1550);
or U1635 (N_1635,N_1524,N_1516);
and U1636 (N_1636,N_1546,N_1440);
nor U1637 (N_1637,N_1407,N_1565);
or U1638 (N_1638,N_1479,N_1405);
nand U1639 (N_1639,N_1452,N_1560);
and U1640 (N_1640,N_1492,N_1589);
and U1641 (N_1641,N_1576,N_1585);
and U1642 (N_1642,N_1526,N_1454);
xnor U1643 (N_1643,N_1400,N_1416);
and U1644 (N_1644,N_1577,N_1460);
nor U1645 (N_1645,N_1481,N_1581);
and U1646 (N_1646,N_1410,N_1498);
or U1647 (N_1647,N_1532,N_1404);
or U1648 (N_1648,N_1459,N_1597);
nor U1649 (N_1649,N_1531,N_1444);
nand U1650 (N_1650,N_1417,N_1569);
nand U1651 (N_1651,N_1530,N_1449);
nor U1652 (N_1652,N_1588,N_1425);
nor U1653 (N_1653,N_1475,N_1535);
nand U1654 (N_1654,N_1505,N_1409);
and U1655 (N_1655,N_1568,N_1462);
nor U1656 (N_1656,N_1533,N_1414);
xor U1657 (N_1657,N_1559,N_1523);
or U1658 (N_1658,N_1443,N_1487);
and U1659 (N_1659,N_1519,N_1453);
or U1660 (N_1660,N_1470,N_1473);
nor U1661 (N_1661,N_1495,N_1415);
nor U1662 (N_1662,N_1579,N_1490);
nor U1663 (N_1663,N_1542,N_1494);
nand U1664 (N_1664,N_1570,N_1591);
nor U1665 (N_1665,N_1464,N_1513);
nand U1666 (N_1666,N_1486,N_1562);
nand U1667 (N_1667,N_1419,N_1587);
or U1668 (N_1668,N_1517,N_1515);
nand U1669 (N_1669,N_1574,N_1599);
and U1670 (N_1670,N_1468,N_1580);
nand U1671 (N_1671,N_1474,N_1408);
or U1672 (N_1672,N_1500,N_1520);
and U1673 (N_1673,N_1447,N_1427);
and U1674 (N_1674,N_1439,N_1411);
and U1675 (N_1675,N_1448,N_1436);
or U1676 (N_1676,N_1435,N_1412);
or U1677 (N_1677,N_1598,N_1402);
nand U1678 (N_1678,N_1572,N_1445);
or U1679 (N_1679,N_1484,N_1426);
or U1680 (N_1680,N_1489,N_1534);
and U1681 (N_1681,N_1586,N_1537);
nor U1682 (N_1682,N_1420,N_1555);
and U1683 (N_1683,N_1573,N_1512);
and U1684 (N_1684,N_1545,N_1596);
nand U1685 (N_1685,N_1590,N_1421);
and U1686 (N_1686,N_1566,N_1509);
nor U1687 (N_1687,N_1429,N_1497);
nand U1688 (N_1688,N_1424,N_1431);
nor U1689 (N_1689,N_1575,N_1451);
or U1690 (N_1690,N_1522,N_1478);
and U1691 (N_1691,N_1467,N_1441);
or U1692 (N_1692,N_1544,N_1508);
nor U1693 (N_1693,N_1567,N_1514);
and U1694 (N_1694,N_1456,N_1561);
and U1695 (N_1695,N_1541,N_1540);
or U1696 (N_1696,N_1406,N_1469);
xnor U1697 (N_1697,N_1553,N_1457);
or U1698 (N_1698,N_1511,N_1465);
nand U1699 (N_1699,N_1592,N_1493);
nor U1700 (N_1700,N_1568,N_1436);
nor U1701 (N_1701,N_1416,N_1524);
or U1702 (N_1702,N_1590,N_1423);
and U1703 (N_1703,N_1481,N_1556);
or U1704 (N_1704,N_1435,N_1551);
and U1705 (N_1705,N_1501,N_1560);
or U1706 (N_1706,N_1488,N_1523);
nand U1707 (N_1707,N_1595,N_1541);
nand U1708 (N_1708,N_1401,N_1551);
nor U1709 (N_1709,N_1408,N_1448);
nor U1710 (N_1710,N_1492,N_1409);
xor U1711 (N_1711,N_1445,N_1520);
and U1712 (N_1712,N_1427,N_1587);
nor U1713 (N_1713,N_1549,N_1406);
or U1714 (N_1714,N_1434,N_1582);
nor U1715 (N_1715,N_1474,N_1421);
nor U1716 (N_1716,N_1577,N_1454);
nor U1717 (N_1717,N_1495,N_1423);
and U1718 (N_1718,N_1539,N_1434);
nand U1719 (N_1719,N_1579,N_1409);
nor U1720 (N_1720,N_1484,N_1489);
and U1721 (N_1721,N_1495,N_1565);
nor U1722 (N_1722,N_1476,N_1403);
nand U1723 (N_1723,N_1514,N_1562);
or U1724 (N_1724,N_1495,N_1419);
nor U1725 (N_1725,N_1482,N_1522);
nand U1726 (N_1726,N_1554,N_1437);
or U1727 (N_1727,N_1545,N_1485);
nand U1728 (N_1728,N_1551,N_1535);
nand U1729 (N_1729,N_1439,N_1537);
nand U1730 (N_1730,N_1439,N_1518);
nor U1731 (N_1731,N_1544,N_1488);
or U1732 (N_1732,N_1566,N_1588);
or U1733 (N_1733,N_1467,N_1573);
and U1734 (N_1734,N_1410,N_1579);
nand U1735 (N_1735,N_1562,N_1591);
nand U1736 (N_1736,N_1407,N_1586);
or U1737 (N_1737,N_1557,N_1587);
or U1738 (N_1738,N_1451,N_1403);
nor U1739 (N_1739,N_1522,N_1400);
nor U1740 (N_1740,N_1439,N_1543);
nand U1741 (N_1741,N_1562,N_1400);
and U1742 (N_1742,N_1403,N_1449);
nor U1743 (N_1743,N_1591,N_1434);
or U1744 (N_1744,N_1503,N_1470);
and U1745 (N_1745,N_1546,N_1568);
nor U1746 (N_1746,N_1501,N_1416);
nor U1747 (N_1747,N_1472,N_1481);
or U1748 (N_1748,N_1456,N_1447);
nor U1749 (N_1749,N_1400,N_1454);
and U1750 (N_1750,N_1407,N_1441);
nand U1751 (N_1751,N_1520,N_1454);
or U1752 (N_1752,N_1593,N_1546);
nor U1753 (N_1753,N_1470,N_1421);
and U1754 (N_1754,N_1439,N_1469);
nor U1755 (N_1755,N_1526,N_1478);
nor U1756 (N_1756,N_1533,N_1563);
nand U1757 (N_1757,N_1482,N_1491);
nor U1758 (N_1758,N_1535,N_1418);
nor U1759 (N_1759,N_1574,N_1555);
nand U1760 (N_1760,N_1541,N_1567);
or U1761 (N_1761,N_1570,N_1412);
nor U1762 (N_1762,N_1599,N_1572);
or U1763 (N_1763,N_1487,N_1517);
and U1764 (N_1764,N_1497,N_1528);
and U1765 (N_1765,N_1457,N_1487);
nor U1766 (N_1766,N_1447,N_1432);
nand U1767 (N_1767,N_1459,N_1551);
or U1768 (N_1768,N_1540,N_1467);
or U1769 (N_1769,N_1533,N_1492);
nand U1770 (N_1770,N_1520,N_1568);
or U1771 (N_1771,N_1570,N_1519);
and U1772 (N_1772,N_1599,N_1486);
nor U1773 (N_1773,N_1455,N_1496);
or U1774 (N_1774,N_1577,N_1422);
or U1775 (N_1775,N_1537,N_1520);
and U1776 (N_1776,N_1457,N_1535);
and U1777 (N_1777,N_1589,N_1590);
nand U1778 (N_1778,N_1558,N_1528);
nor U1779 (N_1779,N_1424,N_1425);
or U1780 (N_1780,N_1456,N_1441);
nor U1781 (N_1781,N_1403,N_1559);
or U1782 (N_1782,N_1598,N_1496);
nand U1783 (N_1783,N_1594,N_1435);
and U1784 (N_1784,N_1457,N_1488);
nor U1785 (N_1785,N_1492,N_1438);
nand U1786 (N_1786,N_1467,N_1501);
and U1787 (N_1787,N_1526,N_1432);
and U1788 (N_1788,N_1473,N_1575);
and U1789 (N_1789,N_1466,N_1527);
and U1790 (N_1790,N_1494,N_1472);
and U1791 (N_1791,N_1400,N_1456);
nor U1792 (N_1792,N_1504,N_1507);
and U1793 (N_1793,N_1448,N_1432);
or U1794 (N_1794,N_1506,N_1512);
nand U1795 (N_1795,N_1515,N_1473);
nand U1796 (N_1796,N_1475,N_1454);
nor U1797 (N_1797,N_1452,N_1483);
nor U1798 (N_1798,N_1481,N_1417);
nor U1799 (N_1799,N_1448,N_1499);
or U1800 (N_1800,N_1767,N_1796);
or U1801 (N_1801,N_1634,N_1783);
nor U1802 (N_1802,N_1797,N_1661);
nand U1803 (N_1803,N_1731,N_1648);
nand U1804 (N_1804,N_1721,N_1624);
or U1805 (N_1805,N_1620,N_1759);
nand U1806 (N_1806,N_1708,N_1679);
nand U1807 (N_1807,N_1752,N_1741);
nor U1808 (N_1808,N_1655,N_1610);
nor U1809 (N_1809,N_1794,N_1725);
nand U1810 (N_1810,N_1615,N_1740);
or U1811 (N_1811,N_1680,N_1652);
and U1812 (N_1812,N_1612,N_1710);
nand U1813 (N_1813,N_1630,N_1674);
and U1814 (N_1814,N_1696,N_1607);
nand U1815 (N_1815,N_1733,N_1686);
nor U1816 (N_1816,N_1753,N_1777);
or U1817 (N_1817,N_1700,N_1750);
and U1818 (N_1818,N_1769,N_1697);
nor U1819 (N_1819,N_1659,N_1699);
nor U1820 (N_1820,N_1606,N_1644);
and U1821 (N_1821,N_1738,N_1685);
nor U1822 (N_1822,N_1760,N_1650);
or U1823 (N_1823,N_1799,N_1706);
or U1824 (N_1824,N_1623,N_1715);
nand U1825 (N_1825,N_1719,N_1614);
or U1826 (N_1826,N_1660,N_1734);
and U1827 (N_1827,N_1773,N_1724);
nor U1828 (N_1828,N_1736,N_1732);
or U1829 (N_1829,N_1601,N_1751);
and U1830 (N_1830,N_1766,N_1691);
or U1831 (N_1831,N_1664,N_1718);
or U1832 (N_1832,N_1657,N_1792);
nand U1833 (N_1833,N_1716,N_1681);
nand U1834 (N_1834,N_1662,N_1742);
or U1835 (N_1835,N_1683,N_1694);
nand U1836 (N_1836,N_1682,N_1621);
and U1837 (N_1837,N_1779,N_1762);
nand U1838 (N_1838,N_1763,N_1778);
or U1839 (N_1839,N_1717,N_1602);
nor U1840 (N_1840,N_1789,N_1647);
nand U1841 (N_1841,N_1771,N_1663);
or U1842 (N_1842,N_1730,N_1653);
nor U1843 (N_1843,N_1635,N_1627);
or U1844 (N_1844,N_1641,N_1656);
or U1845 (N_1845,N_1711,N_1619);
nand U1846 (N_1846,N_1714,N_1654);
or U1847 (N_1847,N_1600,N_1625);
or U1848 (N_1848,N_1622,N_1651);
nor U1849 (N_1849,N_1720,N_1791);
or U1850 (N_1850,N_1688,N_1748);
nand U1851 (N_1851,N_1729,N_1788);
and U1852 (N_1852,N_1605,N_1626);
nor U1853 (N_1853,N_1701,N_1643);
nor U1854 (N_1854,N_1687,N_1629);
or U1855 (N_1855,N_1632,N_1772);
nand U1856 (N_1856,N_1727,N_1709);
nand U1857 (N_1857,N_1678,N_1616);
or U1858 (N_1858,N_1669,N_1705);
and U1859 (N_1859,N_1603,N_1702);
and U1860 (N_1860,N_1722,N_1745);
nor U1861 (N_1861,N_1713,N_1690);
nand U1862 (N_1862,N_1695,N_1786);
or U1863 (N_1863,N_1768,N_1739);
nor U1864 (N_1864,N_1646,N_1746);
or U1865 (N_1865,N_1787,N_1611);
and U1866 (N_1866,N_1780,N_1782);
and U1867 (N_1867,N_1723,N_1761);
and U1868 (N_1868,N_1618,N_1747);
nand U1869 (N_1869,N_1689,N_1617);
nor U1870 (N_1870,N_1665,N_1784);
nor U1871 (N_1871,N_1609,N_1798);
nand U1872 (N_1872,N_1671,N_1672);
nand U1873 (N_1873,N_1636,N_1604);
and U1874 (N_1874,N_1684,N_1675);
nor U1875 (N_1875,N_1639,N_1793);
nor U1876 (N_1876,N_1764,N_1703);
nand U1877 (N_1877,N_1781,N_1785);
nand U1878 (N_1878,N_1638,N_1795);
and U1879 (N_1879,N_1774,N_1667);
xnor U1880 (N_1880,N_1670,N_1668);
and U1881 (N_1881,N_1726,N_1735);
or U1882 (N_1882,N_1770,N_1677);
nand U1883 (N_1883,N_1744,N_1712);
or U1884 (N_1884,N_1633,N_1756);
or U1885 (N_1885,N_1631,N_1776);
or U1886 (N_1886,N_1698,N_1613);
nor U1887 (N_1887,N_1649,N_1754);
nor U1888 (N_1888,N_1743,N_1737);
or U1889 (N_1889,N_1645,N_1658);
nand U1890 (N_1890,N_1765,N_1790);
or U1891 (N_1891,N_1673,N_1707);
nor U1892 (N_1892,N_1637,N_1757);
and U1893 (N_1893,N_1704,N_1755);
and U1894 (N_1894,N_1642,N_1676);
xor U1895 (N_1895,N_1758,N_1749);
or U1896 (N_1896,N_1666,N_1608);
nor U1897 (N_1897,N_1775,N_1692);
xnor U1898 (N_1898,N_1693,N_1628);
and U1899 (N_1899,N_1728,N_1640);
or U1900 (N_1900,N_1605,N_1734);
nor U1901 (N_1901,N_1696,N_1682);
and U1902 (N_1902,N_1623,N_1754);
nor U1903 (N_1903,N_1672,N_1679);
nor U1904 (N_1904,N_1653,N_1736);
nand U1905 (N_1905,N_1670,N_1718);
or U1906 (N_1906,N_1792,N_1750);
or U1907 (N_1907,N_1776,N_1696);
or U1908 (N_1908,N_1688,N_1770);
nand U1909 (N_1909,N_1765,N_1654);
nand U1910 (N_1910,N_1613,N_1763);
or U1911 (N_1911,N_1770,N_1792);
and U1912 (N_1912,N_1712,N_1650);
nor U1913 (N_1913,N_1772,N_1621);
and U1914 (N_1914,N_1790,N_1660);
nor U1915 (N_1915,N_1656,N_1699);
and U1916 (N_1916,N_1601,N_1645);
or U1917 (N_1917,N_1633,N_1733);
and U1918 (N_1918,N_1662,N_1747);
nor U1919 (N_1919,N_1627,N_1612);
and U1920 (N_1920,N_1750,N_1693);
xor U1921 (N_1921,N_1749,N_1689);
and U1922 (N_1922,N_1643,N_1797);
nand U1923 (N_1923,N_1687,N_1764);
or U1924 (N_1924,N_1769,N_1673);
and U1925 (N_1925,N_1664,N_1795);
or U1926 (N_1926,N_1606,N_1607);
and U1927 (N_1927,N_1667,N_1734);
or U1928 (N_1928,N_1749,N_1765);
or U1929 (N_1929,N_1638,N_1620);
nor U1930 (N_1930,N_1607,N_1770);
or U1931 (N_1931,N_1726,N_1697);
and U1932 (N_1932,N_1714,N_1690);
nor U1933 (N_1933,N_1769,N_1614);
nor U1934 (N_1934,N_1782,N_1622);
and U1935 (N_1935,N_1626,N_1710);
nand U1936 (N_1936,N_1680,N_1666);
nand U1937 (N_1937,N_1694,N_1736);
and U1938 (N_1938,N_1667,N_1608);
nand U1939 (N_1939,N_1676,N_1753);
and U1940 (N_1940,N_1704,N_1656);
or U1941 (N_1941,N_1666,N_1743);
or U1942 (N_1942,N_1730,N_1781);
nor U1943 (N_1943,N_1628,N_1606);
nor U1944 (N_1944,N_1713,N_1704);
or U1945 (N_1945,N_1761,N_1766);
nor U1946 (N_1946,N_1658,N_1708);
nand U1947 (N_1947,N_1623,N_1636);
nand U1948 (N_1948,N_1619,N_1640);
nand U1949 (N_1949,N_1658,N_1699);
nor U1950 (N_1950,N_1637,N_1691);
or U1951 (N_1951,N_1660,N_1714);
nand U1952 (N_1952,N_1785,N_1755);
nor U1953 (N_1953,N_1780,N_1682);
or U1954 (N_1954,N_1616,N_1665);
xor U1955 (N_1955,N_1622,N_1737);
xor U1956 (N_1956,N_1796,N_1723);
nor U1957 (N_1957,N_1626,N_1667);
xnor U1958 (N_1958,N_1675,N_1627);
and U1959 (N_1959,N_1660,N_1642);
xor U1960 (N_1960,N_1701,N_1674);
nor U1961 (N_1961,N_1637,N_1736);
or U1962 (N_1962,N_1630,N_1729);
and U1963 (N_1963,N_1630,N_1620);
xor U1964 (N_1964,N_1617,N_1651);
xnor U1965 (N_1965,N_1727,N_1691);
nor U1966 (N_1966,N_1743,N_1732);
nor U1967 (N_1967,N_1646,N_1651);
and U1968 (N_1968,N_1625,N_1643);
nor U1969 (N_1969,N_1685,N_1747);
or U1970 (N_1970,N_1763,N_1620);
nand U1971 (N_1971,N_1625,N_1785);
nand U1972 (N_1972,N_1615,N_1680);
nor U1973 (N_1973,N_1776,N_1761);
nand U1974 (N_1974,N_1707,N_1664);
or U1975 (N_1975,N_1727,N_1734);
and U1976 (N_1976,N_1685,N_1683);
nor U1977 (N_1977,N_1746,N_1661);
or U1978 (N_1978,N_1605,N_1687);
or U1979 (N_1979,N_1640,N_1679);
or U1980 (N_1980,N_1702,N_1764);
or U1981 (N_1981,N_1645,N_1673);
or U1982 (N_1982,N_1606,N_1616);
or U1983 (N_1983,N_1687,N_1700);
and U1984 (N_1984,N_1769,N_1687);
nor U1985 (N_1985,N_1705,N_1736);
or U1986 (N_1986,N_1729,N_1736);
nor U1987 (N_1987,N_1710,N_1728);
nor U1988 (N_1988,N_1741,N_1731);
nor U1989 (N_1989,N_1725,N_1753);
and U1990 (N_1990,N_1601,N_1705);
and U1991 (N_1991,N_1769,N_1753);
or U1992 (N_1992,N_1727,N_1694);
nand U1993 (N_1993,N_1600,N_1679);
nor U1994 (N_1994,N_1744,N_1792);
nand U1995 (N_1995,N_1629,N_1762);
or U1996 (N_1996,N_1776,N_1732);
nand U1997 (N_1997,N_1653,N_1600);
and U1998 (N_1998,N_1788,N_1699);
or U1999 (N_1999,N_1793,N_1682);
or U2000 (N_2000,N_1910,N_1806);
nand U2001 (N_2001,N_1831,N_1982);
and U2002 (N_2002,N_1857,N_1882);
or U2003 (N_2003,N_1977,N_1930);
or U2004 (N_2004,N_1926,N_1864);
nand U2005 (N_2005,N_1959,N_1851);
and U2006 (N_2006,N_1922,N_1802);
nand U2007 (N_2007,N_1804,N_1801);
nor U2008 (N_2008,N_1933,N_1971);
xnor U2009 (N_2009,N_1991,N_1872);
and U2010 (N_2010,N_1875,N_1853);
nand U2011 (N_2011,N_1927,N_1810);
nand U2012 (N_2012,N_1808,N_1989);
nand U2013 (N_2013,N_1805,N_1844);
or U2014 (N_2014,N_1811,N_1845);
or U2015 (N_2015,N_1825,N_1992);
or U2016 (N_2016,N_1894,N_1969);
nand U2017 (N_2017,N_1919,N_1861);
xnor U2018 (N_2018,N_1813,N_1909);
nand U2019 (N_2019,N_1859,N_1812);
or U2020 (N_2020,N_1895,N_1837);
or U2021 (N_2021,N_1877,N_1896);
and U2022 (N_2022,N_1945,N_1914);
or U2023 (N_2023,N_1824,N_1958);
nor U2024 (N_2024,N_1957,N_1905);
nor U2025 (N_2025,N_1954,N_1918);
nor U2026 (N_2026,N_1986,N_1974);
and U2027 (N_2027,N_1803,N_1809);
or U2028 (N_2028,N_1822,N_1807);
or U2029 (N_2029,N_1902,N_1846);
nor U2030 (N_2030,N_1967,N_1978);
or U2031 (N_2031,N_1965,N_1884);
nand U2032 (N_2032,N_1893,N_1998);
nor U2033 (N_2033,N_1976,N_1943);
and U2034 (N_2034,N_1887,N_1862);
and U2035 (N_2035,N_1836,N_1947);
nor U2036 (N_2036,N_1869,N_1953);
nand U2037 (N_2037,N_1913,N_1904);
nor U2038 (N_2038,N_1841,N_1987);
nor U2039 (N_2039,N_1962,N_1979);
nand U2040 (N_2040,N_1983,N_1972);
and U2041 (N_2041,N_1973,N_1963);
and U2042 (N_2042,N_1888,N_1984);
or U2043 (N_2043,N_1815,N_1827);
nor U2044 (N_2044,N_1931,N_1880);
nor U2045 (N_2045,N_1964,N_1871);
or U2046 (N_2046,N_1951,N_1940);
or U2047 (N_2047,N_1906,N_1903);
and U2048 (N_2048,N_1874,N_1800);
nand U2049 (N_2049,N_1900,N_1823);
nand U2050 (N_2050,N_1925,N_1942);
nand U2051 (N_2051,N_1995,N_1936);
or U2052 (N_2052,N_1879,N_1929);
xnor U2053 (N_2053,N_1838,N_1817);
nor U2054 (N_2054,N_1981,N_1941);
nor U2055 (N_2055,N_1826,N_1829);
nor U2056 (N_2056,N_1840,N_1960);
nor U2057 (N_2057,N_1863,N_1821);
nand U2058 (N_2058,N_1816,N_1956);
and U2059 (N_2059,N_1892,N_1849);
nor U2060 (N_2060,N_1867,N_1928);
nand U2061 (N_2061,N_1833,N_1916);
nand U2062 (N_2062,N_1912,N_1876);
or U2063 (N_2063,N_1886,N_1889);
or U2064 (N_2064,N_1949,N_1854);
nor U2065 (N_2065,N_1890,N_1915);
nor U2066 (N_2066,N_1921,N_1938);
and U2067 (N_2067,N_1834,N_1946);
nand U2068 (N_2068,N_1924,N_1897);
or U2069 (N_2069,N_1891,N_1939);
nor U2070 (N_2070,N_1999,N_1856);
and U2071 (N_2071,N_1873,N_1950);
or U2072 (N_2072,N_1866,N_1852);
and U2073 (N_2073,N_1934,N_1980);
or U2074 (N_2074,N_1907,N_1868);
and U2075 (N_2075,N_1988,N_1848);
or U2076 (N_2076,N_1937,N_1885);
nor U2077 (N_2077,N_1835,N_1993);
nor U2078 (N_2078,N_1860,N_1883);
and U2079 (N_2079,N_1911,N_1878);
or U2080 (N_2080,N_1818,N_1948);
or U2081 (N_2081,N_1898,N_1917);
nand U2082 (N_2082,N_1975,N_1966);
nor U2083 (N_2083,N_1843,N_1830);
or U2084 (N_2084,N_1935,N_1908);
or U2085 (N_2085,N_1881,N_1855);
nor U2086 (N_2086,N_1990,N_1955);
and U2087 (N_2087,N_1865,N_1952);
or U2088 (N_2088,N_1994,N_1985);
nand U2089 (N_2089,N_1944,N_1899);
and U2090 (N_2090,N_1839,N_1920);
or U2091 (N_2091,N_1858,N_1847);
nand U2092 (N_2092,N_1828,N_1968);
nand U2093 (N_2093,N_1970,N_1870);
or U2094 (N_2094,N_1901,N_1923);
nand U2095 (N_2095,N_1996,N_1850);
and U2096 (N_2096,N_1932,N_1832);
nor U2097 (N_2097,N_1997,N_1819);
and U2098 (N_2098,N_1814,N_1842);
and U2099 (N_2099,N_1961,N_1820);
or U2100 (N_2100,N_1897,N_1915);
and U2101 (N_2101,N_1952,N_1869);
nand U2102 (N_2102,N_1973,N_1829);
and U2103 (N_2103,N_1959,N_1986);
nor U2104 (N_2104,N_1985,N_1956);
or U2105 (N_2105,N_1904,N_1912);
nor U2106 (N_2106,N_1864,N_1880);
nor U2107 (N_2107,N_1939,N_1831);
or U2108 (N_2108,N_1880,N_1984);
nand U2109 (N_2109,N_1808,N_1868);
nor U2110 (N_2110,N_1841,N_1827);
and U2111 (N_2111,N_1961,N_1868);
or U2112 (N_2112,N_1856,N_1969);
and U2113 (N_2113,N_1801,N_1862);
nand U2114 (N_2114,N_1846,N_1838);
nand U2115 (N_2115,N_1872,N_1839);
or U2116 (N_2116,N_1867,N_1861);
nand U2117 (N_2117,N_1900,N_1996);
and U2118 (N_2118,N_1983,N_1886);
nor U2119 (N_2119,N_1840,N_1891);
or U2120 (N_2120,N_1860,N_1859);
nor U2121 (N_2121,N_1844,N_1884);
and U2122 (N_2122,N_1806,N_1970);
nand U2123 (N_2123,N_1997,N_1839);
or U2124 (N_2124,N_1872,N_1916);
nand U2125 (N_2125,N_1954,N_1905);
or U2126 (N_2126,N_1833,N_1810);
or U2127 (N_2127,N_1819,N_1821);
and U2128 (N_2128,N_1814,N_1966);
nand U2129 (N_2129,N_1996,N_1914);
and U2130 (N_2130,N_1837,N_1982);
nor U2131 (N_2131,N_1802,N_1951);
nor U2132 (N_2132,N_1910,N_1929);
or U2133 (N_2133,N_1825,N_1808);
or U2134 (N_2134,N_1800,N_1883);
or U2135 (N_2135,N_1889,N_1809);
nor U2136 (N_2136,N_1870,N_1997);
or U2137 (N_2137,N_1982,N_1977);
nand U2138 (N_2138,N_1985,N_1841);
nor U2139 (N_2139,N_1948,N_1993);
nand U2140 (N_2140,N_1927,N_1894);
nor U2141 (N_2141,N_1973,N_1890);
or U2142 (N_2142,N_1946,N_1810);
nor U2143 (N_2143,N_1836,N_1821);
or U2144 (N_2144,N_1827,N_1803);
and U2145 (N_2145,N_1992,N_1883);
nand U2146 (N_2146,N_1988,N_1857);
nand U2147 (N_2147,N_1883,N_1871);
or U2148 (N_2148,N_1943,N_1898);
nand U2149 (N_2149,N_1935,N_1815);
nor U2150 (N_2150,N_1929,N_1899);
nand U2151 (N_2151,N_1917,N_1936);
or U2152 (N_2152,N_1832,N_1948);
and U2153 (N_2153,N_1989,N_1964);
nor U2154 (N_2154,N_1894,N_1839);
nand U2155 (N_2155,N_1945,N_1932);
nand U2156 (N_2156,N_1947,N_1987);
and U2157 (N_2157,N_1942,N_1872);
and U2158 (N_2158,N_1937,N_1813);
nand U2159 (N_2159,N_1829,N_1873);
and U2160 (N_2160,N_1806,N_1862);
nor U2161 (N_2161,N_1846,N_1865);
or U2162 (N_2162,N_1888,N_1813);
nand U2163 (N_2163,N_1864,N_1980);
nor U2164 (N_2164,N_1892,N_1813);
nand U2165 (N_2165,N_1985,N_1937);
or U2166 (N_2166,N_1860,N_1809);
nor U2167 (N_2167,N_1990,N_1964);
and U2168 (N_2168,N_1824,N_1833);
or U2169 (N_2169,N_1819,N_1884);
nand U2170 (N_2170,N_1994,N_1872);
nand U2171 (N_2171,N_1801,N_1808);
and U2172 (N_2172,N_1843,N_1815);
or U2173 (N_2173,N_1821,N_1824);
nor U2174 (N_2174,N_1842,N_1942);
and U2175 (N_2175,N_1814,N_1834);
nand U2176 (N_2176,N_1988,N_1844);
and U2177 (N_2177,N_1889,N_1896);
nor U2178 (N_2178,N_1906,N_1962);
and U2179 (N_2179,N_1884,N_1899);
nor U2180 (N_2180,N_1935,N_1829);
nor U2181 (N_2181,N_1855,N_1826);
nand U2182 (N_2182,N_1980,N_1961);
and U2183 (N_2183,N_1988,N_1882);
nor U2184 (N_2184,N_1933,N_1863);
nand U2185 (N_2185,N_1830,N_1880);
nand U2186 (N_2186,N_1850,N_1883);
nor U2187 (N_2187,N_1856,N_1852);
and U2188 (N_2188,N_1922,N_1800);
and U2189 (N_2189,N_1981,N_1901);
nand U2190 (N_2190,N_1849,N_1903);
or U2191 (N_2191,N_1864,N_1822);
nand U2192 (N_2192,N_1957,N_1947);
and U2193 (N_2193,N_1913,N_1915);
nor U2194 (N_2194,N_1839,N_1946);
nor U2195 (N_2195,N_1970,N_1950);
nor U2196 (N_2196,N_1950,N_1907);
nand U2197 (N_2197,N_1856,N_1887);
nand U2198 (N_2198,N_1930,N_1949);
and U2199 (N_2199,N_1879,N_1983);
nand U2200 (N_2200,N_2046,N_2157);
nor U2201 (N_2201,N_2103,N_2057);
nor U2202 (N_2202,N_2129,N_2159);
or U2203 (N_2203,N_2024,N_2147);
and U2204 (N_2204,N_2111,N_2174);
nor U2205 (N_2205,N_2125,N_2079);
and U2206 (N_2206,N_2171,N_2016);
nor U2207 (N_2207,N_2012,N_2176);
or U2208 (N_2208,N_2102,N_2136);
and U2209 (N_2209,N_2052,N_2199);
or U2210 (N_2210,N_2084,N_2184);
or U2211 (N_2211,N_2183,N_2180);
and U2212 (N_2212,N_2143,N_2175);
or U2213 (N_2213,N_2100,N_2077);
nor U2214 (N_2214,N_2163,N_2121);
and U2215 (N_2215,N_2109,N_2044);
nand U2216 (N_2216,N_2127,N_2197);
or U2217 (N_2217,N_2085,N_2075);
and U2218 (N_2218,N_2099,N_2123);
and U2219 (N_2219,N_2006,N_2178);
nand U2220 (N_2220,N_2071,N_2089);
or U2221 (N_2221,N_2078,N_2166);
and U2222 (N_2222,N_2040,N_2132);
and U2223 (N_2223,N_2139,N_2117);
nor U2224 (N_2224,N_2135,N_2060);
nor U2225 (N_2225,N_2005,N_2082);
or U2226 (N_2226,N_2122,N_2058);
nand U2227 (N_2227,N_2134,N_2140);
or U2228 (N_2228,N_2148,N_2039);
nand U2229 (N_2229,N_2104,N_2098);
or U2230 (N_2230,N_2113,N_2149);
nor U2231 (N_2231,N_2061,N_2186);
or U2232 (N_2232,N_2032,N_2120);
and U2233 (N_2233,N_2118,N_2073);
nand U2234 (N_2234,N_2172,N_2086);
or U2235 (N_2235,N_2043,N_2144);
nor U2236 (N_2236,N_2054,N_2170);
nor U2237 (N_2237,N_2145,N_2025);
nand U2238 (N_2238,N_2003,N_2177);
or U2239 (N_2239,N_2094,N_2187);
and U2240 (N_2240,N_2072,N_2126);
or U2241 (N_2241,N_2023,N_2080);
and U2242 (N_2242,N_2000,N_2059);
nor U2243 (N_2243,N_2055,N_2151);
or U2244 (N_2244,N_2188,N_2093);
or U2245 (N_2245,N_2002,N_2069);
and U2246 (N_2246,N_2007,N_2161);
and U2247 (N_2247,N_2115,N_2181);
or U2248 (N_2248,N_2090,N_2088);
nor U2249 (N_2249,N_2001,N_2097);
nor U2250 (N_2250,N_2068,N_2026);
nand U2251 (N_2251,N_2066,N_2105);
or U2252 (N_2252,N_2092,N_2168);
or U2253 (N_2253,N_2138,N_2008);
and U2254 (N_2254,N_2070,N_2156);
or U2255 (N_2255,N_2037,N_2050);
nor U2256 (N_2256,N_2133,N_2033);
nor U2257 (N_2257,N_2164,N_2036);
nor U2258 (N_2258,N_2131,N_2167);
or U2259 (N_2259,N_2116,N_2114);
or U2260 (N_2260,N_2049,N_2194);
or U2261 (N_2261,N_2019,N_2014);
or U2262 (N_2262,N_2190,N_2124);
or U2263 (N_2263,N_2095,N_2027);
nor U2264 (N_2264,N_2196,N_2051);
nor U2265 (N_2265,N_2042,N_2169);
nor U2266 (N_2266,N_2110,N_2022);
nor U2267 (N_2267,N_2021,N_2053);
or U2268 (N_2268,N_2074,N_2153);
and U2269 (N_2269,N_2011,N_2152);
nor U2270 (N_2270,N_2150,N_2063);
or U2271 (N_2271,N_2038,N_2160);
or U2272 (N_2272,N_2018,N_2119);
nand U2273 (N_2273,N_2162,N_2064);
nor U2274 (N_2274,N_2076,N_2004);
and U2275 (N_2275,N_2047,N_2193);
and U2276 (N_2276,N_2045,N_2195);
or U2277 (N_2277,N_2096,N_2137);
or U2278 (N_2278,N_2009,N_2091);
nor U2279 (N_2279,N_2065,N_2031);
and U2280 (N_2280,N_2107,N_2146);
nor U2281 (N_2281,N_2141,N_2142);
nor U2282 (N_2282,N_2048,N_2056);
and U2283 (N_2283,N_2035,N_2112);
nand U2284 (N_2284,N_2020,N_2106);
nor U2285 (N_2285,N_2029,N_2165);
and U2286 (N_2286,N_2185,N_2034);
or U2287 (N_2287,N_2015,N_2154);
nand U2288 (N_2288,N_2158,N_2182);
and U2289 (N_2289,N_2017,N_2191);
or U2290 (N_2290,N_2062,N_2192);
and U2291 (N_2291,N_2041,N_2198);
nand U2292 (N_2292,N_2128,N_2010);
and U2293 (N_2293,N_2083,N_2173);
xnor U2294 (N_2294,N_2081,N_2179);
nand U2295 (N_2295,N_2028,N_2155);
and U2296 (N_2296,N_2189,N_2108);
nor U2297 (N_2297,N_2130,N_2030);
nand U2298 (N_2298,N_2087,N_2067);
or U2299 (N_2299,N_2013,N_2101);
nand U2300 (N_2300,N_2032,N_2173);
or U2301 (N_2301,N_2005,N_2132);
nor U2302 (N_2302,N_2041,N_2036);
nand U2303 (N_2303,N_2118,N_2120);
and U2304 (N_2304,N_2070,N_2167);
and U2305 (N_2305,N_2150,N_2117);
nand U2306 (N_2306,N_2004,N_2033);
or U2307 (N_2307,N_2011,N_2142);
nand U2308 (N_2308,N_2124,N_2191);
nand U2309 (N_2309,N_2176,N_2166);
nand U2310 (N_2310,N_2117,N_2093);
nor U2311 (N_2311,N_2042,N_2161);
nand U2312 (N_2312,N_2160,N_2142);
and U2313 (N_2313,N_2031,N_2112);
nor U2314 (N_2314,N_2075,N_2018);
nor U2315 (N_2315,N_2099,N_2170);
nor U2316 (N_2316,N_2063,N_2011);
nand U2317 (N_2317,N_2157,N_2114);
or U2318 (N_2318,N_2094,N_2183);
nand U2319 (N_2319,N_2187,N_2157);
nor U2320 (N_2320,N_2003,N_2146);
or U2321 (N_2321,N_2092,N_2050);
nand U2322 (N_2322,N_2034,N_2189);
or U2323 (N_2323,N_2045,N_2072);
nand U2324 (N_2324,N_2131,N_2026);
nand U2325 (N_2325,N_2111,N_2159);
nor U2326 (N_2326,N_2009,N_2020);
and U2327 (N_2327,N_2003,N_2072);
nand U2328 (N_2328,N_2038,N_2106);
nor U2329 (N_2329,N_2104,N_2072);
nor U2330 (N_2330,N_2164,N_2146);
and U2331 (N_2331,N_2105,N_2152);
nor U2332 (N_2332,N_2077,N_2106);
nand U2333 (N_2333,N_2177,N_2014);
or U2334 (N_2334,N_2041,N_2131);
nand U2335 (N_2335,N_2187,N_2125);
nand U2336 (N_2336,N_2139,N_2008);
and U2337 (N_2337,N_2111,N_2031);
nand U2338 (N_2338,N_2088,N_2028);
or U2339 (N_2339,N_2127,N_2081);
nand U2340 (N_2340,N_2100,N_2156);
or U2341 (N_2341,N_2000,N_2046);
or U2342 (N_2342,N_2066,N_2142);
or U2343 (N_2343,N_2085,N_2111);
nand U2344 (N_2344,N_2143,N_2156);
nor U2345 (N_2345,N_2061,N_2009);
nand U2346 (N_2346,N_2139,N_2030);
and U2347 (N_2347,N_2111,N_2062);
and U2348 (N_2348,N_2091,N_2066);
nand U2349 (N_2349,N_2071,N_2017);
nor U2350 (N_2350,N_2005,N_2044);
and U2351 (N_2351,N_2071,N_2103);
nand U2352 (N_2352,N_2003,N_2170);
or U2353 (N_2353,N_2114,N_2055);
and U2354 (N_2354,N_2005,N_2138);
or U2355 (N_2355,N_2173,N_2061);
nand U2356 (N_2356,N_2033,N_2145);
and U2357 (N_2357,N_2070,N_2162);
or U2358 (N_2358,N_2010,N_2120);
and U2359 (N_2359,N_2067,N_2170);
or U2360 (N_2360,N_2060,N_2049);
and U2361 (N_2361,N_2125,N_2199);
nor U2362 (N_2362,N_2190,N_2137);
nand U2363 (N_2363,N_2051,N_2068);
nor U2364 (N_2364,N_2011,N_2143);
and U2365 (N_2365,N_2015,N_2159);
or U2366 (N_2366,N_2027,N_2140);
or U2367 (N_2367,N_2112,N_2032);
nand U2368 (N_2368,N_2189,N_2185);
or U2369 (N_2369,N_2098,N_2114);
or U2370 (N_2370,N_2039,N_2073);
nand U2371 (N_2371,N_2119,N_2107);
nor U2372 (N_2372,N_2187,N_2055);
and U2373 (N_2373,N_2173,N_2148);
and U2374 (N_2374,N_2043,N_2089);
and U2375 (N_2375,N_2075,N_2003);
nor U2376 (N_2376,N_2044,N_2062);
nand U2377 (N_2377,N_2041,N_2121);
nor U2378 (N_2378,N_2074,N_2052);
or U2379 (N_2379,N_2196,N_2092);
nor U2380 (N_2380,N_2026,N_2104);
nand U2381 (N_2381,N_2119,N_2136);
nor U2382 (N_2382,N_2060,N_2104);
or U2383 (N_2383,N_2147,N_2107);
nor U2384 (N_2384,N_2090,N_2057);
or U2385 (N_2385,N_2154,N_2127);
and U2386 (N_2386,N_2086,N_2189);
nor U2387 (N_2387,N_2154,N_2066);
nor U2388 (N_2388,N_2124,N_2046);
or U2389 (N_2389,N_2110,N_2175);
and U2390 (N_2390,N_2094,N_2025);
and U2391 (N_2391,N_2187,N_2144);
and U2392 (N_2392,N_2064,N_2052);
nor U2393 (N_2393,N_2199,N_2139);
nand U2394 (N_2394,N_2097,N_2053);
nor U2395 (N_2395,N_2062,N_2090);
nand U2396 (N_2396,N_2194,N_2016);
and U2397 (N_2397,N_2136,N_2025);
and U2398 (N_2398,N_2043,N_2046);
nand U2399 (N_2399,N_2011,N_2111);
or U2400 (N_2400,N_2367,N_2229);
nand U2401 (N_2401,N_2325,N_2362);
or U2402 (N_2402,N_2284,N_2223);
or U2403 (N_2403,N_2300,N_2259);
nand U2404 (N_2404,N_2280,N_2269);
or U2405 (N_2405,N_2270,N_2234);
or U2406 (N_2406,N_2351,N_2309);
nor U2407 (N_2407,N_2294,N_2253);
or U2408 (N_2408,N_2252,N_2208);
and U2409 (N_2409,N_2271,N_2272);
xor U2410 (N_2410,N_2215,N_2239);
or U2411 (N_2411,N_2293,N_2263);
nand U2412 (N_2412,N_2368,N_2345);
and U2413 (N_2413,N_2261,N_2366);
and U2414 (N_2414,N_2307,N_2321);
nor U2415 (N_2415,N_2278,N_2371);
or U2416 (N_2416,N_2361,N_2308);
or U2417 (N_2417,N_2343,N_2224);
nand U2418 (N_2418,N_2295,N_2383);
nor U2419 (N_2419,N_2329,N_2203);
and U2420 (N_2420,N_2274,N_2242);
or U2421 (N_2421,N_2398,N_2357);
nand U2422 (N_2422,N_2227,N_2245);
nor U2423 (N_2423,N_2247,N_2399);
xor U2424 (N_2424,N_2276,N_2216);
or U2425 (N_2425,N_2334,N_2297);
nor U2426 (N_2426,N_2221,N_2249);
nor U2427 (N_2427,N_2290,N_2380);
or U2428 (N_2428,N_2360,N_2205);
nand U2429 (N_2429,N_2246,N_2340);
nand U2430 (N_2430,N_2363,N_2244);
and U2431 (N_2431,N_2265,N_2254);
xnor U2432 (N_2432,N_2299,N_2328);
nor U2433 (N_2433,N_2241,N_2303);
nor U2434 (N_2434,N_2313,N_2291);
nand U2435 (N_2435,N_2317,N_2326);
nand U2436 (N_2436,N_2289,N_2302);
nand U2437 (N_2437,N_2220,N_2304);
nor U2438 (N_2438,N_2267,N_2232);
or U2439 (N_2439,N_2335,N_2288);
nand U2440 (N_2440,N_2332,N_2339);
and U2441 (N_2441,N_2237,N_2238);
nand U2442 (N_2442,N_2320,N_2262);
and U2443 (N_2443,N_2222,N_2354);
nand U2444 (N_2444,N_2369,N_2352);
and U2445 (N_2445,N_2212,N_2201);
nand U2446 (N_2446,N_2217,N_2377);
or U2447 (N_2447,N_2281,N_2250);
and U2448 (N_2448,N_2344,N_2277);
nand U2449 (N_2449,N_2218,N_2268);
nand U2450 (N_2450,N_2266,N_2384);
nor U2451 (N_2451,N_2375,N_2393);
and U2452 (N_2452,N_2347,N_2319);
or U2453 (N_2453,N_2337,N_2349);
and U2454 (N_2454,N_2397,N_2350);
nor U2455 (N_2455,N_2382,N_2260);
and U2456 (N_2456,N_2359,N_2391);
nor U2457 (N_2457,N_2286,N_2327);
or U2458 (N_2458,N_2379,N_2213);
and U2459 (N_2459,N_2228,N_2214);
and U2460 (N_2460,N_2355,N_2318);
nor U2461 (N_2461,N_2386,N_2283);
nor U2462 (N_2462,N_2305,N_2202);
or U2463 (N_2463,N_2285,N_2209);
and U2464 (N_2464,N_2240,N_2396);
nand U2465 (N_2465,N_2353,N_2389);
and U2466 (N_2466,N_2388,N_2275);
and U2467 (N_2467,N_2210,N_2233);
nor U2468 (N_2468,N_2207,N_2374);
or U2469 (N_2469,N_2211,N_2392);
nand U2470 (N_2470,N_2279,N_2292);
nor U2471 (N_2471,N_2230,N_2225);
and U2472 (N_2472,N_2236,N_2231);
or U2473 (N_2473,N_2372,N_2394);
xor U2474 (N_2474,N_2333,N_2257);
nand U2475 (N_2475,N_2316,N_2204);
or U2476 (N_2476,N_2311,N_2356);
or U2477 (N_2477,N_2346,N_2331);
nor U2478 (N_2478,N_2365,N_2336);
xor U2479 (N_2479,N_2251,N_2376);
nor U2480 (N_2480,N_2390,N_2235);
nor U2481 (N_2481,N_2255,N_2373);
and U2482 (N_2482,N_2387,N_2395);
nor U2483 (N_2483,N_2358,N_2342);
xor U2484 (N_2484,N_2323,N_2273);
nand U2485 (N_2485,N_2364,N_2282);
xor U2486 (N_2486,N_2314,N_2310);
or U2487 (N_2487,N_2298,N_2324);
or U2488 (N_2488,N_2312,N_2296);
or U2489 (N_2489,N_2219,N_2248);
nor U2490 (N_2490,N_2330,N_2370);
nor U2491 (N_2491,N_2322,N_2338);
and U2492 (N_2492,N_2378,N_2315);
and U2493 (N_2493,N_2287,N_2306);
or U2494 (N_2494,N_2301,N_2258);
nand U2495 (N_2495,N_2341,N_2200);
nor U2496 (N_2496,N_2264,N_2381);
nand U2497 (N_2497,N_2256,N_2226);
and U2498 (N_2498,N_2385,N_2243);
and U2499 (N_2499,N_2348,N_2206);
nor U2500 (N_2500,N_2223,N_2386);
or U2501 (N_2501,N_2261,N_2207);
nand U2502 (N_2502,N_2227,N_2351);
nor U2503 (N_2503,N_2355,N_2332);
or U2504 (N_2504,N_2237,N_2293);
or U2505 (N_2505,N_2304,N_2236);
nor U2506 (N_2506,N_2251,N_2301);
nand U2507 (N_2507,N_2345,N_2243);
nor U2508 (N_2508,N_2271,N_2264);
or U2509 (N_2509,N_2219,N_2229);
or U2510 (N_2510,N_2248,N_2260);
and U2511 (N_2511,N_2316,N_2347);
nor U2512 (N_2512,N_2341,N_2210);
or U2513 (N_2513,N_2245,N_2341);
and U2514 (N_2514,N_2296,N_2331);
nor U2515 (N_2515,N_2253,N_2238);
nor U2516 (N_2516,N_2337,N_2241);
or U2517 (N_2517,N_2311,N_2368);
nand U2518 (N_2518,N_2273,N_2216);
nand U2519 (N_2519,N_2361,N_2329);
nor U2520 (N_2520,N_2268,N_2220);
nand U2521 (N_2521,N_2209,N_2282);
and U2522 (N_2522,N_2372,N_2351);
and U2523 (N_2523,N_2385,N_2271);
nand U2524 (N_2524,N_2322,N_2217);
nand U2525 (N_2525,N_2396,N_2353);
nand U2526 (N_2526,N_2270,N_2358);
nor U2527 (N_2527,N_2301,N_2325);
nand U2528 (N_2528,N_2223,N_2382);
or U2529 (N_2529,N_2392,N_2225);
nor U2530 (N_2530,N_2390,N_2331);
nor U2531 (N_2531,N_2369,N_2237);
nand U2532 (N_2532,N_2289,N_2288);
and U2533 (N_2533,N_2322,N_2381);
nor U2534 (N_2534,N_2311,N_2245);
or U2535 (N_2535,N_2269,N_2271);
or U2536 (N_2536,N_2332,N_2319);
nand U2537 (N_2537,N_2367,N_2203);
nand U2538 (N_2538,N_2350,N_2227);
or U2539 (N_2539,N_2220,N_2373);
nand U2540 (N_2540,N_2260,N_2322);
and U2541 (N_2541,N_2386,N_2385);
nand U2542 (N_2542,N_2249,N_2316);
and U2543 (N_2543,N_2330,N_2311);
nand U2544 (N_2544,N_2363,N_2321);
or U2545 (N_2545,N_2303,N_2328);
or U2546 (N_2546,N_2212,N_2206);
nand U2547 (N_2547,N_2239,N_2333);
nor U2548 (N_2548,N_2233,N_2310);
nor U2549 (N_2549,N_2391,N_2237);
or U2550 (N_2550,N_2208,N_2325);
nor U2551 (N_2551,N_2287,N_2245);
nor U2552 (N_2552,N_2243,N_2326);
nand U2553 (N_2553,N_2240,N_2235);
nand U2554 (N_2554,N_2221,N_2382);
nand U2555 (N_2555,N_2357,N_2271);
or U2556 (N_2556,N_2329,N_2258);
nand U2557 (N_2557,N_2241,N_2330);
xor U2558 (N_2558,N_2222,N_2277);
and U2559 (N_2559,N_2347,N_2234);
or U2560 (N_2560,N_2202,N_2228);
nand U2561 (N_2561,N_2310,N_2295);
nand U2562 (N_2562,N_2381,N_2291);
nand U2563 (N_2563,N_2220,N_2239);
and U2564 (N_2564,N_2323,N_2387);
nor U2565 (N_2565,N_2260,N_2262);
nand U2566 (N_2566,N_2244,N_2257);
or U2567 (N_2567,N_2266,N_2232);
and U2568 (N_2568,N_2253,N_2345);
and U2569 (N_2569,N_2313,N_2243);
or U2570 (N_2570,N_2281,N_2208);
nor U2571 (N_2571,N_2277,N_2225);
nor U2572 (N_2572,N_2306,N_2381);
nand U2573 (N_2573,N_2211,N_2316);
or U2574 (N_2574,N_2224,N_2276);
nand U2575 (N_2575,N_2329,N_2357);
or U2576 (N_2576,N_2230,N_2370);
nand U2577 (N_2577,N_2304,N_2216);
nand U2578 (N_2578,N_2204,N_2350);
nand U2579 (N_2579,N_2271,N_2225);
and U2580 (N_2580,N_2258,N_2203);
or U2581 (N_2581,N_2351,N_2357);
or U2582 (N_2582,N_2244,N_2291);
or U2583 (N_2583,N_2218,N_2362);
nand U2584 (N_2584,N_2360,N_2217);
nand U2585 (N_2585,N_2289,N_2397);
nor U2586 (N_2586,N_2382,N_2279);
nand U2587 (N_2587,N_2395,N_2246);
or U2588 (N_2588,N_2260,N_2256);
and U2589 (N_2589,N_2242,N_2237);
or U2590 (N_2590,N_2227,N_2287);
and U2591 (N_2591,N_2292,N_2348);
and U2592 (N_2592,N_2352,N_2212);
or U2593 (N_2593,N_2273,N_2382);
nand U2594 (N_2594,N_2375,N_2332);
and U2595 (N_2595,N_2366,N_2397);
and U2596 (N_2596,N_2326,N_2356);
or U2597 (N_2597,N_2225,N_2353);
nor U2598 (N_2598,N_2372,N_2250);
and U2599 (N_2599,N_2337,N_2262);
nand U2600 (N_2600,N_2488,N_2589);
and U2601 (N_2601,N_2549,N_2514);
nand U2602 (N_2602,N_2579,N_2505);
and U2603 (N_2603,N_2440,N_2468);
and U2604 (N_2604,N_2470,N_2525);
nor U2605 (N_2605,N_2567,N_2536);
or U2606 (N_2606,N_2534,N_2432);
nor U2607 (N_2607,N_2489,N_2504);
or U2608 (N_2608,N_2535,N_2582);
nor U2609 (N_2609,N_2403,N_2402);
or U2610 (N_2610,N_2410,N_2598);
and U2611 (N_2611,N_2496,N_2423);
nand U2612 (N_2612,N_2502,N_2583);
nor U2613 (N_2613,N_2543,N_2587);
or U2614 (N_2614,N_2564,N_2561);
or U2615 (N_2615,N_2448,N_2452);
and U2616 (N_2616,N_2434,N_2530);
nand U2617 (N_2617,N_2506,N_2577);
nor U2618 (N_2618,N_2592,N_2517);
and U2619 (N_2619,N_2511,N_2580);
nand U2620 (N_2620,N_2429,N_2510);
nand U2621 (N_2621,N_2466,N_2478);
and U2622 (N_2622,N_2519,N_2487);
nand U2623 (N_2623,N_2435,N_2537);
and U2624 (N_2624,N_2513,N_2586);
or U2625 (N_2625,N_2441,N_2558);
and U2626 (N_2626,N_2411,N_2479);
and U2627 (N_2627,N_2565,N_2526);
and U2628 (N_2628,N_2591,N_2590);
nor U2629 (N_2629,N_2464,N_2493);
nor U2630 (N_2630,N_2424,N_2538);
nor U2631 (N_2631,N_2497,N_2486);
and U2632 (N_2632,N_2548,N_2588);
nor U2633 (N_2633,N_2539,N_2474);
nor U2634 (N_2634,N_2473,N_2422);
nand U2635 (N_2635,N_2557,N_2485);
nor U2636 (N_2636,N_2551,N_2451);
nor U2637 (N_2637,N_2460,N_2472);
or U2638 (N_2638,N_2481,N_2419);
or U2639 (N_2639,N_2584,N_2476);
or U2640 (N_2640,N_2477,N_2457);
nor U2641 (N_2641,N_2544,N_2568);
nand U2642 (N_2642,N_2596,N_2520);
nor U2643 (N_2643,N_2471,N_2401);
or U2644 (N_2644,N_2495,N_2439);
and U2645 (N_2645,N_2599,N_2484);
or U2646 (N_2646,N_2572,N_2503);
nor U2647 (N_2647,N_2461,N_2570);
or U2648 (N_2648,N_2509,N_2450);
and U2649 (N_2649,N_2454,N_2574);
and U2650 (N_2650,N_2566,N_2532);
and U2651 (N_2651,N_2418,N_2542);
or U2652 (N_2652,N_2407,N_2547);
nor U2653 (N_2653,N_2400,N_2420);
xnor U2654 (N_2654,N_2428,N_2508);
nor U2655 (N_2655,N_2545,N_2521);
nor U2656 (N_2656,N_2512,N_2553);
and U2657 (N_2657,N_2430,N_2412);
or U2658 (N_2658,N_2458,N_2500);
nor U2659 (N_2659,N_2524,N_2499);
nor U2660 (N_2660,N_2569,N_2585);
and U2661 (N_2661,N_2527,N_2413);
and U2662 (N_2662,N_2456,N_2404);
and U2663 (N_2663,N_2581,N_2431);
nor U2664 (N_2664,N_2475,N_2406);
nand U2665 (N_2665,N_2453,N_2449);
nand U2666 (N_2666,N_2405,N_2491);
nand U2667 (N_2667,N_2550,N_2507);
or U2668 (N_2668,N_2516,N_2559);
and U2669 (N_2669,N_2546,N_2426);
and U2670 (N_2670,N_2465,N_2409);
and U2671 (N_2671,N_2459,N_2462);
and U2672 (N_2672,N_2552,N_2541);
nand U2673 (N_2673,N_2518,N_2490);
nor U2674 (N_2674,N_2438,N_2563);
or U2675 (N_2675,N_2416,N_2480);
and U2676 (N_2676,N_2522,N_2436);
nor U2677 (N_2677,N_2555,N_2575);
nand U2678 (N_2678,N_2562,N_2576);
nor U2679 (N_2679,N_2501,N_2433);
xor U2680 (N_2680,N_2531,N_2533);
nand U2681 (N_2681,N_2556,N_2425);
and U2682 (N_2682,N_2421,N_2443);
nor U2683 (N_2683,N_2482,N_2554);
and U2684 (N_2684,N_2446,N_2529);
nand U2685 (N_2685,N_2578,N_2437);
nand U2686 (N_2686,N_2445,N_2571);
nor U2687 (N_2687,N_2595,N_2492);
nand U2688 (N_2688,N_2442,N_2463);
or U2689 (N_2689,N_2515,N_2494);
nor U2690 (N_2690,N_2427,N_2447);
nor U2691 (N_2691,N_2444,N_2414);
nor U2692 (N_2692,N_2523,N_2597);
and U2693 (N_2693,N_2593,N_2415);
nor U2694 (N_2694,N_2408,N_2455);
nor U2695 (N_2695,N_2483,N_2498);
and U2696 (N_2696,N_2594,N_2417);
and U2697 (N_2697,N_2540,N_2467);
nor U2698 (N_2698,N_2528,N_2573);
or U2699 (N_2699,N_2560,N_2469);
and U2700 (N_2700,N_2536,N_2512);
nand U2701 (N_2701,N_2580,N_2537);
nor U2702 (N_2702,N_2493,N_2561);
nand U2703 (N_2703,N_2445,N_2429);
nand U2704 (N_2704,N_2570,N_2586);
nand U2705 (N_2705,N_2530,N_2589);
nor U2706 (N_2706,N_2429,N_2590);
or U2707 (N_2707,N_2552,N_2480);
nand U2708 (N_2708,N_2509,N_2514);
and U2709 (N_2709,N_2591,N_2567);
nor U2710 (N_2710,N_2452,N_2586);
nor U2711 (N_2711,N_2511,N_2548);
nand U2712 (N_2712,N_2561,N_2439);
nor U2713 (N_2713,N_2424,N_2541);
and U2714 (N_2714,N_2471,N_2482);
and U2715 (N_2715,N_2425,N_2447);
nor U2716 (N_2716,N_2497,N_2440);
nand U2717 (N_2717,N_2577,N_2515);
nor U2718 (N_2718,N_2421,N_2448);
and U2719 (N_2719,N_2529,N_2561);
nor U2720 (N_2720,N_2427,N_2510);
nor U2721 (N_2721,N_2574,N_2465);
nor U2722 (N_2722,N_2575,N_2448);
and U2723 (N_2723,N_2585,N_2571);
nand U2724 (N_2724,N_2412,N_2551);
and U2725 (N_2725,N_2472,N_2436);
and U2726 (N_2726,N_2462,N_2415);
and U2727 (N_2727,N_2493,N_2468);
nor U2728 (N_2728,N_2552,N_2435);
and U2729 (N_2729,N_2530,N_2475);
nand U2730 (N_2730,N_2579,N_2425);
or U2731 (N_2731,N_2433,N_2403);
or U2732 (N_2732,N_2570,N_2517);
and U2733 (N_2733,N_2579,N_2540);
nor U2734 (N_2734,N_2503,N_2588);
and U2735 (N_2735,N_2540,N_2558);
nor U2736 (N_2736,N_2560,N_2414);
or U2737 (N_2737,N_2527,N_2573);
and U2738 (N_2738,N_2551,N_2484);
or U2739 (N_2739,N_2490,N_2577);
nor U2740 (N_2740,N_2513,N_2572);
or U2741 (N_2741,N_2563,N_2537);
or U2742 (N_2742,N_2596,N_2582);
nand U2743 (N_2743,N_2441,N_2578);
xor U2744 (N_2744,N_2402,N_2430);
or U2745 (N_2745,N_2413,N_2401);
and U2746 (N_2746,N_2506,N_2579);
nand U2747 (N_2747,N_2414,N_2432);
and U2748 (N_2748,N_2423,N_2499);
and U2749 (N_2749,N_2431,N_2487);
and U2750 (N_2750,N_2585,N_2570);
or U2751 (N_2751,N_2420,N_2471);
nand U2752 (N_2752,N_2559,N_2470);
nor U2753 (N_2753,N_2444,N_2404);
or U2754 (N_2754,N_2436,N_2488);
or U2755 (N_2755,N_2571,N_2590);
nor U2756 (N_2756,N_2412,N_2465);
or U2757 (N_2757,N_2541,N_2557);
nor U2758 (N_2758,N_2495,N_2401);
and U2759 (N_2759,N_2434,N_2474);
or U2760 (N_2760,N_2550,N_2578);
nand U2761 (N_2761,N_2431,N_2582);
nand U2762 (N_2762,N_2420,N_2494);
and U2763 (N_2763,N_2552,N_2429);
nor U2764 (N_2764,N_2560,N_2562);
or U2765 (N_2765,N_2478,N_2433);
nor U2766 (N_2766,N_2433,N_2544);
nor U2767 (N_2767,N_2555,N_2427);
or U2768 (N_2768,N_2538,N_2512);
nand U2769 (N_2769,N_2508,N_2432);
nor U2770 (N_2770,N_2514,N_2550);
and U2771 (N_2771,N_2525,N_2463);
nor U2772 (N_2772,N_2530,N_2518);
and U2773 (N_2773,N_2599,N_2590);
nor U2774 (N_2774,N_2496,N_2567);
or U2775 (N_2775,N_2425,N_2467);
nand U2776 (N_2776,N_2494,N_2520);
or U2777 (N_2777,N_2544,N_2503);
or U2778 (N_2778,N_2442,N_2471);
or U2779 (N_2779,N_2490,N_2430);
and U2780 (N_2780,N_2546,N_2404);
or U2781 (N_2781,N_2583,N_2535);
nand U2782 (N_2782,N_2465,N_2592);
nand U2783 (N_2783,N_2415,N_2535);
and U2784 (N_2784,N_2410,N_2539);
and U2785 (N_2785,N_2430,N_2488);
and U2786 (N_2786,N_2591,N_2498);
and U2787 (N_2787,N_2570,N_2437);
nor U2788 (N_2788,N_2493,N_2525);
nand U2789 (N_2789,N_2552,N_2510);
or U2790 (N_2790,N_2473,N_2532);
or U2791 (N_2791,N_2534,N_2431);
nand U2792 (N_2792,N_2449,N_2558);
or U2793 (N_2793,N_2545,N_2482);
nand U2794 (N_2794,N_2527,N_2427);
and U2795 (N_2795,N_2414,N_2448);
and U2796 (N_2796,N_2441,N_2440);
and U2797 (N_2797,N_2437,N_2468);
nor U2798 (N_2798,N_2553,N_2519);
nand U2799 (N_2799,N_2598,N_2576);
or U2800 (N_2800,N_2665,N_2617);
and U2801 (N_2801,N_2711,N_2703);
nor U2802 (N_2802,N_2623,N_2682);
or U2803 (N_2803,N_2693,N_2673);
nand U2804 (N_2804,N_2698,N_2717);
nand U2805 (N_2805,N_2615,N_2742);
nand U2806 (N_2806,N_2733,N_2672);
nand U2807 (N_2807,N_2643,N_2628);
nand U2808 (N_2808,N_2636,N_2605);
and U2809 (N_2809,N_2708,N_2688);
nand U2810 (N_2810,N_2791,N_2757);
or U2811 (N_2811,N_2639,N_2752);
nor U2812 (N_2812,N_2611,N_2724);
or U2813 (N_2813,N_2642,N_2695);
nand U2814 (N_2814,N_2610,N_2762);
and U2815 (N_2815,N_2713,N_2716);
and U2816 (N_2816,N_2771,N_2753);
nor U2817 (N_2817,N_2602,N_2691);
nor U2818 (N_2818,N_2649,N_2741);
or U2819 (N_2819,N_2680,N_2660);
nor U2820 (N_2820,N_2790,N_2766);
or U2821 (N_2821,N_2701,N_2750);
nor U2822 (N_2822,N_2606,N_2777);
and U2823 (N_2823,N_2743,N_2600);
and U2824 (N_2824,N_2630,N_2638);
nand U2825 (N_2825,N_2616,N_2760);
or U2826 (N_2826,N_2761,N_2727);
or U2827 (N_2827,N_2756,N_2629);
nand U2828 (N_2828,N_2645,N_2709);
nand U2829 (N_2829,N_2646,N_2765);
and U2830 (N_2830,N_2626,N_2764);
and U2831 (N_2831,N_2674,N_2787);
and U2832 (N_2832,N_2705,N_2699);
or U2833 (N_2833,N_2782,N_2775);
nand U2834 (N_2834,N_2740,N_2614);
and U2835 (N_2835,N_2671,N_2633);
nor U2836 (N_2836,N_2729,N_2654);
nand U2837 (N_2837,N_2669,N_2748);
or U2838 (N_2838,N_2797,N_2784);
nand U2839 (N_2839,N_2792,N_2655);
nand U2840 (N_2840,N_2613,N_2749);
nor U2841 (N_2841,N_2735,N_2763);
nor U2842 (N_2842,N_2662,N_2624);
and U2843 (N_2843,N_2773,N_2744);
and U2844 (N_2844,N_2607,N_2689);
and U2845 (N_2845,N_2603,N_2641);
nand U2846 (N_2846,N_2650,N_2686);
nand U2847 (N_2847,N_2621,N_2767);
nor U2848 (N_2848,N_2751,N_2786);
or U2849 (N_2849,N_2652,N_2710);
and U2850 (N_2850,N_2653,N_2738);
nor U2851 (N_2851,N_2627,N_2619);
or U2852 (N_2852,N_2685,N_2799);
nand U2853 (N_2853,N_2601,N_2687);
and U2854 (N_2854,N_2656,N_2696);
nand U2855 (N_2855,N_2684,N_2631);
nor U2856 (N_2856,N_2746,N_2759);
nor U2857 (N_2857,N_2768,N_2793);
or U2858 (N_2858,N_2658,N_2651);
nor U2859 (N_2859,N_2676,N_2675);
or U2860 (N_2860,N_2668,N_2620);
and U2861 (N_2861,N_2769,N_2700);
nand U2862 (N_2862,N_2755,N_2778);
and U2863 (N_2863,N_2608,N_2728);
nand U2864 (N_2864,N_2734,N_2795);
nor U2865 (N_2865,N_2697,N_2604);
nand U2866 (N_2866,N_2719,N_2722);
or U2867 (N_2867,N_2702,N_2664);
and U2868 (N_2868,N_2659,N_2657);
and U2869 (N_2869,N_2625,N_2725);
and U2870 (N_2870,N_2788,N_2721);
nand U2871 (N_2871,N_2712,N_2770);
nand U2872 (N_2872,N_2635,N_2681);
nand U2873 (N_2873,N_2715,N_2747);
and U2874 (N_2874,N_2632,N_2723);
or U2875 (N_2875,N_2739,N_2726);
nand U2876 (N_2876,N_2694,N_2634);
nor U2877 (N_2877,N_2720,N_2666);
and U2878 (N_2878,N_2737,N_2647);
and U2879 (N_2879,N_2663,N_2618);
or U2880 (N_2880,N_2683,N_2640);
nand U2881 (N_2881,N_2706,N_2783);
and U2882 (N_2882,N_2718,N_2754);
nand U2883 (N_2883,N_2796,N_2772);
or U2884 (N_2884,N_2678,N_2692);
nor U2885 (N_2885,N_2667,N_2714);
or U2886 (N_2886,N_2731,N_2661);
and U2887 (N_2887,N_2644,N_2707);
and U2888 (N_2888,N_2776,N_2736);
or U2889 (N_2889,N_2612,N_2677);
and U2890 (N_2890,N_2637,N_2704);
and U2891 (N_2891,N_2780,N_2794);
or U2892 (N_2892,N_2774,N_2732);
nand U2893 (N_2893,N_2730,N_2781);
or U2894 (N_2894,N_2798,N_2690);
and U2895 (N_2895,N_2670,N_2789);
xor U2896 (N_2896,N_2679,N_2609);
or U2897 (N_2897,N_2785,N_2745);
nand U2898 (N_2898,N_2758,N_2648);
and U2899 (N_2899,N_2622,N_2779);
nor U2900 (N_2900,N_2684,N_2765);
nand U2901 (N_2901,N_2743,N_2617);
or U2902 (N_2902,N_2708,N_2669);
nor U2903 (N_2903,N_2749,N_2639);
and U2904 (N_2904,N_2745,N_2607);
nor U2905 (N_2905,N_2761,N_2660);
or U2906 (N_2906,N_2732,N_2739);
and U2907 (N_2907,N_2684,N_2648);
or U2908 (N_2908,N_2675,N_2733);
or U2909 (N_2909,N_2693,N_2789);
nand U2910 (N_2910,N_2714,N_2650);
nand U2911 (N_2911,N_2749,N_2665);
or U2912 (N_2912,N_2653,N_2672);
nand U2913 (N_2913,N_2707,N_2663);
or U2914 (N_2914,N_2657,N_2668);
nor U2915 (N_2915,N_2689,N_2731);
nor U2916 (N_2916,N_2643,N_2720);
nand U2917 (N_2917,N_2614,N_2658);
nand U2918 (N_2918,N_2667,N_2662);
or U2919 (N_2919,N_2768,N_2651);
or U2920 (N_2920,N_2623,N_2702);
or U2921 (N_2921,N_2706,N_2787);
nor U2922 (N_2922,N_2726,N_2779);
and U2923 (N_2923,N_2764,N_2630);
and U2924 (N_2924,N_2707,N_2736);
and U2925 (N_2925,N_2641,N_2673);
nand U2926 (N_2926,N_2654,N_2708);
nand U2927 (N_2927,N_2621,N_2772);
or U2928 (N_2928,N_2780,N_2702);
and U2929 (N_2929,N_2624,N_2758);
or U2930 (N_2930,N_2642,N_2612);
nand U2931 (N_2931,N_2686,N_2715);
nand U2932 (N_2932,N_2741,N_2702);
nand U2933 (N_2933,N_2700,N_2705);
and U2934 (N_2934,N_2759,N_2755);
nand U2935 (N_2935,N_2767,N_2684);
nor U2936 (N_2936,N_2715,N_2735);
nor U2937 (N_2937,N_2784,N_2745);
and U2938 (N_2938,N_2693,N_2787);
nand U2939 (N_2939,N_2748,N_2783);
nor U2940 (N_2940,N_2742,N_2709);
nor U2941 (N_2941,N_2658,N_2649);
and U2942 (N_2942,N_2685,N_2741);
and U2943 (N_2943,N_2725,N_2762);
nor U2944 (N_2944,N_2694,N_2740);
or U2945 (N_2945,N_2694,N_2765);
nand U2946 (N_2946,N_2763,N_2679);
and U2947 (N_2947,N_2643,N_2751);
and U2948 (N_2948,N_2745,N_2794);
or U2949 (N_2949,N_2683,N_2764);
and U2950 (N_2950,N_2679,N_2644);
or U2951 (N_2951,N_2677,N_2770);
or U2952 (N_2952,N_2713,N_2680);
or U2953 (N_2953,N_2685,N_2615);
nand U2954 (N_2954,N_2627,N_2655);
nand U2955 (N_2955,N_2642,N_2775);
or U2956 (N_2956,N_2603,N_2647);
nor U2957 (N_2957,N_2796,N_2610);
and U2958 (N_2958,N_2786,N_2699);
nor U2959 (N_2959,N_2630,N_2680);
nand U2960 (N_2960,N_2638,N_2790);
xor U2961 (N_2961,N_2755,N_2796);
nor U2962 (N_2962,N_2700,N_2607);
nand U2963 (N_2963,N_2620,N_2777);
nor U2964 (N_2964,N_2623,N_2649);
nand U2965 (N_2965,N_2719,N_2639);
nand U2966 (N_2966,N_2689,N_2631);
nand U2967 (N_2967,N_2685,N_2706);
and U2968 (N_2968,N_2711,N_2797);
nor U2969 (N_2969,N_2605,N_2679);
or U2970 (N_2970,N_2702,N_2799);
and U2971 (N_2971,N_2637,N_2604);
or U2972 (N_2972,N_2793,N_2749);
nand U2973 (N_2973,N_2663,N_2691);
nor U2974 (N_2974,N_2684,N_2722);
nor U2975 (N_2975,N_2657,N_2727);
nor U2976 (N_2976,N_2657,N_2694);
or U2977 (N_2977,N_2673,N_2633);
or U2978 (N_2978,N_2666,N_2770);
or U2979 (N_2979,N_2606,N_2670);
nand U2980 (N_2980,N_2764,N_2789);
or U2981 (N_2981,N_2632,N_2662);
or U2982 (N_2982,N_2641,N_2694);
and U2983 (N_2983,N_2663,N_2779);
and U2984 (N_2984,N_2772,N_2665);
or U2985 (N_2985,N_2622,N_2743);
nor U2986 (N_2986,N_2717,N_2672);
nor U2987 (N_2987,N_2666,N_2625);
or U2988 (N_2988,N_2780,N_2646);
and U2989 (N_2989,N_2677,N_2726);
or U2990 (N_2990,N_2635,N_2638);
or U2991 (N_2991,N_2756,N_2638);
nand U2992 (N_2992,N_2727,N_2796);
or U2993 (N_2993,N_2619,N_2643);
and U2994 (N_2994,N_2762,N_2686);
nor U2995 (N_2995,N_2789,N_2775);
nand U2996 (N_2996,N_2614,N_2700);
nand U2997 (N_2997,N_2637,N_2682);
nor U2998 (N_2998,N_2738,N_2734);
nor U2999 (N_2999,N_2636,N_2720);
or U3000 (N_3000,N_2951,N_2810);
xnor U3001 (N_3001,N_2923,N_2863);
or U3002 (N_3002,N_2930,N_2904);
nand U3003 (N_3003,N_2932,N_2976);
and U3004 (N_3004,N_2815,N_2903);
nor U3005 (N_3005,N_2895,N_2838);
or U3006 (N_3006,N_2882,N_2966);
and U3007 (N_3007,N_2853,N_2864);
nand U3008 (N_3008,N_2885,N_2816);
and U3009 (N_3009,N_2920,N_2894);
nand U3010 (N_3010,N_2870,N_2841);
or U3011 (N_3011,N_2866,N_2917);
or U3012 (N_3012,N_2948,N_2822);
and U3013 (N_3013,N_2829,N_2813);
nor U3014 (N_3014,N_2846,N_2890);
nor U3015 (N_3015,N_2972,N_2851);
nor U3016 (N_3016,N_2807,N_2985);
or U3017 (N_3017,N_2961,N_2989);
or U3018 (N_3018,N_2913,N_2945);
nor U3019 (N_3019,N_2939,N_2912);
nand U3020 (N_3020,N_2959,N_2995);
or U3021 (N_3021,N_2804,N_2929);
nand U3022 (N_3022,N_2868,N_2955);
nor U3023 (N_3023,N_2861,N_2896);
and U3024 (N_3024,N_2839,N_2997);
nor U3025 (N_3025,N_2935,N_2921);
or U3026 (N_3026,N_2835,N_2879);
nand U3027 (N_3027,N_2978,N_2944);
nand U3028 (N_3028,N_2805,N_2982);
and U3029 (N_3029,N_2949,N_2943);
or U3030 (N_3030,N_2905,N_2821);
nand U3031 (N_3031,N_2899,N_2897);
and U3032 (N_3032,N_2802,N_2809);
nor U3033 (N_3033,N_2991,N_2857);
nor U3034 (N_3034,N_2850,N_2987);
or U3035 (N_3035,N_2918,N_2957);
and U3036 (N_3036,N_2883,N_2862);
and U3037 (N_3037,N_2892,N_2823);
nand U3038 (N_3038,N_2840,N_2977);
nand U3039 (N_3039,N_2963,N_2900);
or U3040 (N_3040,N_2867,N_2849);
nand U3041 (N_3041,N_2832,N_2852);
nand U3042 (N_3042,N_2889,N_2836);
nor U3043 (N_3043,N_2859,N_2884);
nand U3044 (N_3044,N_2803,N_2964);
or U3045 (N_3045,N_2979,N_2937);
or U3046 (N_3046,N_2954,N_2925);
nand U3047 (N_3047,N_2830,N_2993);
or U3048 (N_3048,N_2988,N_2901);
and U3049 (N_3049,N_2916,N_2886);
nand U3050 (N_3050,N_2946,N_2817);
or U3051 (N_3051,N_2994,N_2981);
and U3052 (N_3052,N_2960,N_2927);
and U3053 (N_3053,N_2983,N_2941);
and U3054 (N_3054,N_2953,N_2842);
or U3055 (N_3055,N_2915,N_2996);
nor U3056 (N_3056,N_2940,N_2876);
and U3057 (N_3057,N_2933,N_2888);
and U3058 (N_3058,N_2980,N_2986);
nand U3059 (N_3059,N_2965,N_2924);
nor U3060 (N_3060,N_2818,N_2902);
and U3061 (N_3061,N_2990,N_2906);
or U3062 (N_3062,N_2967,N_2952);
and U3063 (N_3063,N_2909,N_2971);
or U3064 (N_3064,N_2869,N_2812);
nand U3065 (N_3065,N_2898,N_2998);
nand U3066 (N_3066,N_2843,N_2824);
nor U3067 (N_3067,N_2910,N_2828);
nand U3068 (N_3068,N_2936,N_2938);
and U3069 (N_3069,N_2950,N_2992);
and U3070 (N_3070,N_2831,N_2934);
nand U3071 (N_3071,N_2801,N_2922);
nor U3072 (N_3072,N_2865,N_2819);
and U3073 (N_3073,N_2956,N_2947);
nor U3074 (N_3074,N_2928,N_2907);
nor U3075 (N_3075,N_2820,N_2958);
nor U3076 (N_3076,N_2808,N_2825);
nand U3077 (N_3077,N_2962,N_2891);
nor U3078 (N_3078,N_2881,N_2848);
nand U3079 (N_3079,N_2999,N_2860);
nand U3080 (N_3080,N_2834,N_2806);
or U3081 (N_3081,N_2975,N_2814);
nor U3082 (N_3082,N_2837,N_2877);
or U3083 (N_3083,N_2833,N_2873);
nand U3084 (N_3084,N_2969,N_2887);
nand U3085 (N_3085,N_2847,N_2973);
nand U3086 (N_3086,N_2875,N_2893);
and U3087 (N_3087,N_2855,N_2874);
and U3088 (N_3088,N_2974,N_2984);
or U3089 (N_3089,N_2926,N_2800);
nor U3090 (N_3090,N_2871,N_2854);
or U3091 (N_3091,N_2872,N_2811);
and U3092 (N_3092,N_2880,N_2914);
nand U3093 (N_3093,N_2844,N_2931);
and U3094 (N_3094,N_2970,N_2968);
and U3095 (N_3095,N_2826,N_2827);
and U3096 (N_3096,N_2845,N_2942);
and U3097 (N_3097,N_2919,N_2911);
nor U3098 (N_3098,N_2856,N_2878);
nand U3099 (N_3099,N_2908,N_2858);
or U3100 (N_3100,N_2811,N_2861);
nor U3101 (N_3101,N_2823,N_2860);
nand U3102 (N_3102,N_2841,N_2962);
nand U3103 (N_3103,N_2882,N_2824);
and U3104 (N_3104,N_2892,N_2962);
nand U3105 (N_3105,N_2976,N_2830);
nand U3106 (N_3106,N_2854,N_2933);
nor U3107 (N_3107,N_2800,N_2847);
nand U3108 (N_3108,N_2969,N_2808);
and U3109 (N_3109,N_2826,N_2990);
and U3110 (N_3110,N_2833,N_2925);
or U3111 (N_3111,N_2852,N_2889);
nor U3112 (N_3112,N_2813,N_2920);
and U3113 (N_3113,N_2900,N_2983);
and U3114 (N_3114,N_2861,N_2829);
nor U3115 (N_3115,N_2871,N_2868);
and U3116 (N_3116,N_2956,N_2869);
or U3117 (N_3117,N_2989,N_2837);
nand U3118 (N_3118,N_2911,N_2871);
nor U3119 (N_3119,N_2916,N_2907);
nand U3120 (N_3120,N_2865,N_2871);
nor U3121 (N_3121,N_2888,N_2861);
nand U3122 (N_3122,N_2985,N_2951);
nor U3123 (N_3123,N_2839,N_2977);
nor U3124 (N_3124,N_2862,N_2940);
nand U3125 (N_3125,N_2994,N_2941);
or U3126 (N_3126,N_2845,N_2957);
and U3127 (N_3127,N_2958,N_2998);
and U3128 (N_3128,N_2841,N_2974);
nor U3129 (N_3129,N_2957,N_2852);
or U3130 (N_3130,N_2907,N_2978);
and U3131 (N_3131,N_2808,N_2994);
or U3132 (N_3132,N_2823,N_2882);
nor U3133 (N_3133,N_2990,N_2823);
or U3134 (N_3134,N_2806,N_2958);
nor U3135 (N_3135,N_2880,N_2886);
nand U3136 (N_3136,N_2853,N_2921);
nor U3137 (N_3137,N_2800,N_2878);
or U3138 (N_3138,N_2852,N_2951);
nand U3139 (N_3139,N_2890,N_2849);
nand U3140 (N_3140,N_2851,N_2819);
or U3141 (N_3141,N_2972,N_2825);
nor U3142 (N_3142,N_2892,N_2846);
and U3143 (N_3143,N_2881,N_2809);
nor U3144 (N_3144,N_2950,N_2821);
and U3145 (N_3145,N_2905,N_2833);
nor U3146 (N_3146,N_2856,N_2997);
nand U3147 (N_3147,N_2912,N_2943);
and U3148 (N_3148,N_2912,N_2882);
or U3149 (N_3149,N_2917,N_2994);
or U3150 (N_3150,N_2835,N_2837);
nor U3151 (N_3151,N_2840,N_2852);
nand U3152 (N_3152,N_2950,N_2949);
nand U3153 (N_3153,N_2953,N_2835);
nand U3154 (N_3154,N_2976,N_2892);
and U3155 (N_3155,N_2950,N_2876);
or U3156 (N_3156,N_2885,N_2847);
nor U3157 (N_3157,N_2927,N_2940);
nor U3158 (N_3158,N_2848,N_2873);
nor U3159 (N_3159,N_2967,N_2889);
nor U3160 (N_3160,N_2806,N_2858);
or U3161 (N_3161,N_2889,N_2931);
nand U3162 (N_3162,N_2819,N_2880);
nand U3163 (N_3163,N_2992,N_2830);
nand U3164 (N_3164,N_2993,N_2836);
and U3165 (N_3165,N_2821,N_2953);
or U3166 (N_3166,N_2986,N_2895);
and U3167 (N_3167,N_2941,N_2853);
nor U3168 (N_3168,N_2866,N_2956);
nand U3169 (N_3169,N_2897,N_2894);
or U3170 (N_3170,N_2806,N_2823);
or U3171 (N_3171,N_2961,N_2809);
or U3172 (N_3172,N_2851,N_2841);
nand U3173 (N_3173,N_2832,N_2935);
or U3174 (N_3174,N_2902,N_2949);
or U3175 (N_3175,N_2838,N_2843);
nand U3176 (N_3176,N_2986,N_2964);
and U3177 (N_3177,N_2931,N_2933);
and U3178 (N_3178,N_2948,N_2924);
and U3179 (N_3179,N_2960,N_2914);
nor U3180 (N_3180,N_2920,N_2815);
and U3181 (N_3181,N_2975,N_2847);
and U3182 (N_3182,N_2978,N_2831);
nor U3183 (N_3183,N_2849,N_2958);
nand U3184 (N_3184,N_2970,N_2898);
nor U3185 (N_3185,N_2923,N_2802);
and U3186 (N_3186,N_2897,N_2963);
and U3187 (N_3187,N_2838,N_2938);
nor U3188 (N_3188,N_2901,N_2876);
or U3189 (N_3189,N_2937,N_2986);
or U3190 (N_3190,N_2955,N_2817);
nor U3191 (N_3191,N_2800,N_2916);
and U3192 (N_3192,N_2879,N_2914);
nand U3193 (N_3193,N_2845,N_2906);
nor U3194 (N_3194,N_2806,N_2931);
nor U3195 (N_3195,N_2879,N_2833);
or U3196 (N_3196,N_2935,N_2852);
nand U3197 (N_3197,N_2846,N_2996);
and U3198 (N_3198,N_2934,N_2970);
and U3199 (N_3199,N_2857,N_2900);
or U3200 (N_3200,N_3151,N_3000);
or U3201 (N_3201,N_3096,N_3043);
or U3202 (N_3202,N_3094,N_3008);
nor U3203 (N_3203,N_3017,N_3146);
or U3204 (N_3204,N_3058,N_3167);
or U3205 (N_3205,N_3108,N_3143);
or U3206 (N_3206,N_3119,N_3186);
nor U3207 (N_3207,N_3191,N_3052);
or U3208 (N_3208,N_3003,N_3135);
or U3209 (N_3209,N_3071,N_3120);
and U3210 (N_3210,N_3172,N_3041);
and U3211 (N_3211,N_3114,N_3182);
nand U3212 (N_3212,N_3034,N_3196);
nand U3213 (N_3213,N_3161,N_3020);
nor U3214 (N_3214,N_3060,N_3045);
and U3215 (N_3215,N_3183,N_3171);
nor U3216 (N_3216,N_3074,N_3103);
nor U3217 (N_3217,N_3198,N_3144);
or U3218 (N_3218,N_3177,N_3173);
nor U3219 (N_3219,N_3073,N_3072);
or U3220 (N_3220,N_3145,N_3085);
and U3221 (N_3221,N_3106,N_3004);
nand U3222 (N_3222,N_3134,N_3057);
or U3223 (N_3223,N_3112,N_3054);
and U3224 (N_3224,N_3010,N_3076);
nand U3225 (N_3225,N_3037,N_3123);
nand U3226 (N_3226,N_3166,N_3040);
and U3227 (N_3227,N_3097,N_3049);
or U3228 (N_3228,N_3086,N_3091);
nand U3229 (N_3229,N_3111,N_3067);
nor U3230 (N_3230,N_3092,N_3019);
and U3231 (N_3231,N_3031,N_3180);
or U3232 (N_3232,N_3065,N_3053);
or U3233 (N_3233,N_3062,N_3070);
or U3234 (N_3234,N_3176,N_3050);
and U3235 (N_3235,N_3026,N_3175);
and U3236 (N_3236,N_3185,N_3142);
nand U3237 (N_3237,N_3088,N_3115);
nor U3238 (N_3238,N_3007,N_3027);
nand U3239 (N_3239,N_3124,N_3153);
and U3240 (N_3240,N_3002,N_3035);
nor U3241 (N_3241,N_3001,N_3018);
or U3242 (N_3242,N_3078,N_3121);
nor U3243 (N_3243,N_3136,N_3055);
nor U3244 (N_3244,N_3098,N_3051);
or U3245 (N_3245,N_3100,N_3129);
and U3246 (N_3246,N_3046,N_3148);
nand U3247 (N_3247,N_3199,N_3133);
and U3248 (N_3248,N_3081,N_3022);
and U3249 (N_3249,N_3154,N_3168);
and U3250 (N_3250,N_3126,N_3197);
nor U3251 (N_3251,N_3080,N_3087);
nor U3252 (N_3252,N_3117,N_3156);
nor U3253 (N_3253,N_3044,N_3024);
or U3254 (N_3254,N_3130,N_3089);
nor U3255 (N_3255,N_3102,N_3016);
or U3256 (N_3256,N_3162,N_3033);
nand U3257 (N_3257,N_3083,N_3039);
nor U3258 (N_3258,N_3109,N_3132);
or U3259 (N_3259,N_3158,N_3169);
and U3260 (N_3260,N_3061,N_3042);
nand U3261 (N_3261,N_3194,N_3059);
nor U3262 (N_3262,N_3150,N_3107);
and U3263 (N_3263,N_3138,N_3118);
nor U3264 (N_3264,N_3157,N_3140);
or U3265 (N_3265,N_3164,N_3137);
nand U3266 (N_3266,N_3069,N_3063);
nand U3267 (N_3267,N_3104,N_3079);
or U3268 (N_3268,N_3192,N_3099);
nand U3269 (N_3269,N_3187,N_3110);
nand U3270 (N_3270,N_3101,N_3015);
or U3271 (N_3271,N_3011,N_3032);
or U3272 (N_3272,N_3122,N_3077);
and U3273 (N_3273,N_3149,N_3029);
or U3274 (N_3274,N_3005,N_3064);
nand U3275 (N_3275,N_3189,N_3066);
and U3276 (N_3276,N_3179,N_3093);
and U3277 (N_3277,N_3127,N_3021);
nand U3278 (N_3278,N_3181,N_3116);
or U3279 (N_3279,N_3141,N_3084);
or U3280 (N_3280,N_3025,N_3174);
or U3281 (N_3281,N_3125,N_3068);
nor U3282 (N_3282,N_3023,N_3131);
or U3283 (N_3283,N_3170,N_3013);
and U3284 (N_3284,N_3159,N_3193);
or U3285 (N_3285,N_3075,N_3152);
and U3286 (N_3286,N_3165,N_3128);
and U3287 (N_3287,N_3048,N_3184);
and U3288 (N_3288,N_3147,N_3105);
nand U3289 (N_3289,N_3082,N_3113);
nand U3290 (N_3290,N_3012,N_3056);
nor U3291 (N_3291,N_3038,N_3095);
and U3292 (N_3292,N_3014,N_3009);
or U3293 (N_3293,N_3028,N_3195);
or U3294 (N_3294,N_3155,N_3006);
nand U3295 (N_3295,N_3190,N_3047);
nand U3296 (N_3296,N_3163,N_3188);
nand U3297 (N_3297,N_3160,N_3178);
and U3298 (N_3298,N_3030,N_3036);
nor U3299 (N_3299,N_3090,N_3139);
nand U3300 (N_3300,N_3198,N_3095);
nand U3301 (N_3301,N_3021,N_3015);
or U3302 (N_3302,N_3196,N_3173);
or U3303 (N_3303,N_3021,N_3051);
nand U3304 (N_3304,N_3094,N_3152);
nor U3305 (N_3305,N_3187,N_3036);
nand U3306 (N_3306,N_3135,N_3144);
nor U3307 (N_3307,N_3143,N_3136);
nor U3308 (N_3308,N_3103,N_3071);
nand U3309 (N_3309,N_3012,N_3091);
or U3310 (N_3310,N_3161,N_3097);
nand U3311 (N_3311,N_3036,N_3163);
nor U3312 (N_3312,N_3089,N_3051);
nor U3313 (N_3313,N_3091,N_3141);
or U3314 (N_3314,N_3119,N_3160);
nand U3315 (N_3315,N_3016,N_3052);
nand U3316 (N_3316,N_3031,N_3098);
nand U3317 (N_3317,N_3177,N_3175);
nor U3318 (N_3318,N_3109,N_3036);
nor U3319 (N_3319,N_3166,N_3187);
and U3320 (N_3320,N_3030,N_3164);
and U3321 (N_3321,N_3127,N_3084);
xor U3322 (N_3322,N_3142,N_3082);
nor U3323 (N_3323,N_3134,N_3063);
or U3324 (N_3324,N_3186,N_3098);
or U3325 (N_3325,N_3147,N_3165);
nor U3326 (N_3326,N_3048,N_3180);
nor U3327 (N_3327,N_3046,N_3111);
or U3328 (N_3328,N_3083,N_3032);
or U3329 (N_3329,N_3051,N_3029);
or U3330 (N_3330,N_3150,N_3121);
and U3331 (N_3331,N_3008,N_3065);
and U3332 (N_3332,N_3101,N_3150);
and U3333 (N_3333,N_3194,N_3046);
nand U3334 (N_3334,N_3020,N_3183);
nor U3335 (N_3335,N_3119,N_3135);
nor U3336 (N_3336,N_3102,N_3127);
nor U3337 (N_3337,N_3055,N_3051);
nor U3338 (N_3338,N_3158,N_3128);
and U3339 (N_3339,N_3020,N_3104);
nor U3340 (N_3340,N_3158,N_3166);
and U3341 (N_3341,N_3062,N_3186);
or U3342 (N_3342,N_3011,N_3066);
and U3343 (N_3343,N_3005,N_3171);
nand U3344 (N_3344,N_3060,N_3127);
and U3345 (N_3345,N_3152,N_3102);
nand U3346 (N_3346,N_3089,N_3100);
or U3347 (N_3347,N_3146,N_3044);
and U3348 (N_3348,N_3149,N_3089);
nor U3349 (N_3349,N_3035,N_3055);
and U3350 (N_3350,N_3073,N_3147);
and U3351 (N_3351,N_3199,N_3155);
nor U3352 (N_3352,N_3032,N_3025);
nand U3353 (N_3353,N_3150,N_3022);
nor U3354 (N_3354,N_3009,N_3072);
or U3355 (N_3355,N_3058,N_3009);
and U3356 (N_3356,N_3002,N_3040);
and U3357 (N_3357,N_3084,N_3123);
and U3358 (N_3358,N_3170,N_3138);
nand U3359 (N_3359,N_3075,N_3136);
or U3360 (N_3360,N_3159,N_3117);
nand U3361 (N_3361,N_3153,N_3030);
nor U3362 (N_3362,N_3047,N_3154);
nor U3363 (N_3363,N_3019,N_3095);
and U3364 (N_3364,N_3016,N_3081);
nand U3365 (N_3365,N_3004,N_3005);
nand U3366 (N_3366,N_3081,N_3120);
and U3367 (N_3367,N_3043,N_3021);
nor U3368 (N_3368,N_3021,N_3040);
xnor U3369 (N_3369,N_3179,N_3002);
or U3370 (N_3370,N_3181,N_3194);
or U3371 (N_3371,N_3131,N_3183);
and U3372 (N_3372,N_3150,N_3118);
nand U3373 (N_3373,N_3017,N_3036);
nand U3374 (N_3374,N_3187,N_3169);
or U3375 (N_3375,N_3049,N_3062);
nand U3376 (N_3376,N_3055,N_3156);
nor U3377 (N_3377,N_3198,N_3191);
and U3378 (N_3378,N_3026,N_3138);
and U3379 (N_3379,N_3089,N_3142);
and U3380 (N_3380,N_3029,N_3195);
or U3381 (N_3381,N_3139,N_3103);
or U3382 (N_3382,N_3111,N_3082);
and U3383 (N_3383,N_3169,N_3049);
xor U3384 (N_3384,N_3134,N_3165);
nor U3385 (N_3385,N_3085,N_3193);
and U3386 (N_3386,N_3113,N_3142);
nand U3387 (N_3387,N_3036,N_3041);
nor U3388 (N_3388,N_3033,N_3040);
and U3389 (N_3389,N_3150,N_3141);
nand U3390 (N_3390,N_3136,N_3173);
nor U3391 (N_3391,N_3152,N_3053);
or U3392 (N_3392,N_3185,N_3131);
or U3393 (N_3393,N_3139,N_3002);
nor U3394 (N_3394,N_3103,N_3030);
or U3395 (N_3395,N_3107,N_3003);
and U3396 (N_3396,N_3155,N_3073);
or U3397 (N_3397,N_3196,N_3055);
and U3398 (N_3398,N_3002,N_3004);
and U3399 (N_3399,N_3086,N_3072);
nand U3400 (N_3400,N_3386,N_3210);
or U3401 (N_3401,N_3346,N_3306);
and U3402 (N_3402,N_3270,N_3271);
nand U3403 (N_3403,N_3266,N_3360);
nor U3404 (N_3404,N_3282,N_3285);
nand U3405 (N_3405,N_3324,N_3269);
or U3406 (N_3406,N_3305,N_3246);
nor U3407 (N_3407,N_3368,N_3329);
or U3408 (N_3408,N_3314,N_3348);
or U3409 (N_3409,N_3311,N_3223);
nor U3410 (N_3410,N_3370,N_3297);
and U3411 (N_3411,N_3365,N_3352);
and U3412 (N_3412,N_3242,N_3310);
and U3413 (N_3413,N_3273,N_3251);
or U3414 (N_3414,N_3294,N_3215);
nor U3415 (N_3415,N_3379,N_3367);
nor U3416 (N_3416,N_3250,N_3366);
and U3417 (N_3417,N_3385,N_3323);
or U3418 (N_3418,N_3369,N_3397);
nor U3419 (N_3419,N_3298,N_3286);
nand U3420 (N_3420,N_3353,N_3384);
and U3421 (N_3421,N_3300,N_3301);
or U3422 (N_3422,N_3345,N_3299);
nand U3423 (N_3423,N_3339,N_3265);
nand U3424 (N_3424,N_3238,N_3331);
xor U3425 (N_3425,N_3227,N_3380);
and U3426 (N_3426,N_3293,N_3214);
or U3427 (N_3427,N_3391,N_3207);
or U3428 (N_3428,N_3230,N_3376);
or U3429 (N_3429,N_3244,N_3392);
nand U3430 (N_3430,N_3290,N_3222);
nand U3431 (N_3431,N_3302,N_3268);
and U3432 (N_3432,N_3204,N_3337);
nor U3433 (N_3433,N_3387,N_3307);
and U3434 (N_3434,N_3228,N_3281);
and U3435 (N_3435,N_3260,N_3333);
nand U3436 (N_3436,N_3274,N_3358);
nor U3437 (N_3437,N_3364,N_3218);
or U3438 (N_3438,N_3327,N_3381);
or U3439 (N_3439,N_3389,N_3377);
nand U3440 (N_3440,N_3334,N_3320);
nand U3441 (N_3441,N_3241,N_3236);
nor U3442 (N_3442,N_3350,N_3219);
nand U3443 (N_3443,N_3295,N_3374);
or U3444 (N_3444,N_3213,N_3232);
nor U3445 (N_3445,N_3254,N_3308);
or U3446 (N_3446,N_3292,N_3205);
nand U3447 (N_3447,N_3383,N_3344);
nor U3448 (N_3448,N_3351,N_3208);
nand U3449 (N_3449,N_3328,N_3280);
and U3450 (N_3450,N_3239,N_3343);
nor U3451 (N_3451,N_3259,N_3388);
or U3452 (N_3452,N_3362,N_3378);
nor U3453 (N_3453,N_3315,N_3296);
nor U3454 (N_3454,N_3396,N_3326);
and U3455 (N_3455,N_3224,N_3288);
nand U3456 (N_3456,N_3363,N_3338);
nor U3457 (N_3457,N_3357,N_3216);
and U3458 (N_3458,N_3203,N_3336);
or U3459 (N_3459,N_3325,N_3247);
and U3460 (N_3460,N_3399,N_3304);
or U3461 (N_3461,N_3316,N_3283);
nor U3462 (N_3462,N_3211,N_3356);
or U3463 (N_3463,N_3245,N_3382);
or U3464 (N_3464,N_3291,N_3319);
nor U3465 (N_3465,N_3335,N_3221);
nand U3466 (N_3466,N_3341,N_3220);
or U3467 (N_3467,N_3375,N_3234);
and U3468 (N_3468,N_3371,N_3229);
and U3469 (N_3469,N_3309,N_3263);
or U3470 (N_3470,N_3275,N_3279);
nor U3471 (N_3471,N_3277,N_3253);
and U3472 (N_3472,N_3209,N_3258);
nor U3473 (N_3473,N_3373,N_3330);
nor U3474 (N_3474,N_3252,N_3354);
nor U3475 (N_3475,N_3217,N_3243);
or U3476 (N_3476,N_3226,N_3361);
and U3477 (N_3477,N_3332,N_3255);
nor U3478 (N_3478,N_3398,N_3390);
and U3479 (N_3479,N_3322,N_3202);
or U3480 (N_3480,N_3240,N_3342);
and U3481 (N_3481,N_3340,N_3372);
nand U3482 (N_3482,N_3237,N_3287);
or U3483 (N_3483,N_3289,N_3200);
or U3484 (N_3484,N_3212,N_3264);
nand U3485 (N_3485,N_3347,N_3231);
xor U3486 (N_3486,N_3321,N_3261);
or U3487 (N_3487,N_3349,N_3249);
or U3488 (N_3488,N_3272,N_3256);
or U3489 (N_3489,N_3267,N_3318);
xor U3490 (N_3490,N_3276,N_3233);
nand U3491 (N_3491,N_3395,N_3284);
nor U3492 (N_3492,N_3313,N_3359);
nand U3493 (N_3493,N_3257,N_3248);
nor U3494 (N_3494,N_3317,N_3235);
or U3495 (N_3495,N_3393,N_3355);
and U3496 (N_3496,N_3312,N_3225);
or U3497 (N_3497,N_3278,N_3303);
nor U3498 (N_3498,N_3201,N_3262);
and U3499 (N_3499,N_3206,N_3394);
or U3500 (N_3500,N_3207,N_3241);
or U3501 (N_3501,N_3363,N_3339);
nor U3502 (N_3502,N_3223,N_3377);
and U3503 (N_3503,N_3262,N_3210);
nor U3504 (N_3504,N_3283,N_3253);
or U3505 (N_3505,N_3299,N_3323);
nor U3506 (N_3506,N_3263,N_3367);
nor U3507 (N_3507,N_3398,N_3281);
nand U3508 (N_3508,N_3397,N_3248);
nand U3509 (N_3509,N_3372,N_3331);
and U3510 (N_3510,N_3327,N_3270);
nor U3511 (N_3511,N_3372,N_3257);
nor U3512 (N_3512,N_3226,N_3335);
or U3513 (N_3513,N_3394,N_3267);
nor U3514 (N_3514,N_3205,N_3229);
nor U3515 (N_3515,N_3218,N_3303);
nand U3516 (N_3516,N_3310,N_3337);
or U3517 (N_3517,N_3261,N_3337);
nand U3518 (N_3518,N_3377,N_3352);
nor U3519 (N_3519,N_3315,N_3397);
and U3520 (N_3520,N_3388,N_3220);
nor U3521 (N_3521,N_3235,N_3316);
or U3522 (N_3522,N_3357,N_3220);
and U3523 (N_3523,N_3278,N_3358);
nor U3524 (N_3524,N_3350,N_3392);
or U3525 (N_3525,N_3270,N_3260);
nor U3526 (N_3526,N_3294,N_3216);
or U3527 (N_3527,N_3325,N_3330);
nor U3528 (N_3528,N_3360,N_3396);
xor U3529 (N_3529,N_3346,N_3233);
and U3530 (N_3530,N_3227,N_3202);
nor U3531 (N_3531,N_3379,N_3215);
nor U3532 (N_3532,N_3390,N_3207);
nand U3533 (N_3533,N_3215,N_3392);
nor U3534 (N_3534,N_3369,N_3273);
or U3535 (N_3535,N_3278,N_3375);
nand U3536 (N_3536,N_3263,N_3316);
nand U3537 (N_3537,N_3311,N_3326);
and U3538 (N_3538,N_3205,N_3320);
nor U3539 (N_3539,N_3279,N_3246);
nand U3540 (N_3540,N_3324,N_3284);
nor U3541 (N_3541,N_3392,N_3363);
and U3542 (N_3542,N_3368,N_3290);
nor U3543 (N_3543,N_3232,N_3200);
xor U3544 (N_3544,N_3364,N_3369);
and U3545 (N_3545,N_3317,N_3333);
or U3546 (N_3546,N_3384,N_3234);
nand U3547 (N_3547,N_3394,N_3359);
nor U3548 (N_3548,N_3362,N_3224);
nor U3549 (N_3549,N_3327,N_3359);
and U3550 (N_3550,N_3373,N_3378);
nor U3551 (N_3551,N_3356,N_3226);
nand U3552 (N_3552,N_3210,N_3377);
and U3553 (N_3553,N_3387,N_3302);
nor U3554 (N_3554,N_3392,N_3245);
nor U3555 (N_3555,N_3292,N_3222);
and U3556 (N_3556,N_3240,N_3387);
nand U3557 (N_3557,N_3277,N_3302);
nor U3558 (N_3558,N_3376,N_3334);
or U3559 (N_3559,N_3322,N_3328);
or U3560 (N_3560,N_3266,N_3241);
nor U3561 (N_3561,N_3210,N_3391);
nor U3562 (N_3562,N_3394,N_3224);
nor U3563 (N_3563,N_3326,N_3386);
nand U3564 (N_3564,N_3360,N_3241);
nor U3565 (N_3565,N_3379,N_3383);
nor U3566 (N_3566,N_3295,N_3304);
and U3567 (N_3567,N_3217,N_3301);
or U3568 (N_3568,N_3364,N_3247);
nor U3569 (N_3569,N_3204,N_3381);
and U3570 (N_3570,N_3342,N_3216);
or U3571 (N_3571,N_3351,N_3366);
nand U3572 (N_3572,N_3389,N_3390);
and U3573 (N_3573,N_3263,N_3379);
or U3574 (N_3574,N_3297,N_3238);
or U3575 (N_3575,N_3275,N_3285);
and U3576 (N_3576,N_3341,N_3366);
and U3577 (N_3577,N_3361,N_3386);
or U3578 (N_3578,N_3395,N_3225);
nand U3579 (N_3579,N_3370,N_3348);
nand U3580 (N_3580,N_3397,N_3305);
nand U3581 (N_3581,N_3246,N_3247);
nand U3582 (N_3582,N_3266,N_3364);
nor U3583 (N_3583,N_3267,N_3307);
nand U3584 (N_3584,N_3243,N_3256);
and U3585 (N_3585,N_3399,N_3312);
and U3586 (N_3586,N_3247,N_3349);
or U3587 (N_3587,N_3246,N_3399);
nor U3588 (N_3588,N_3290,N_3200);
and U3589 (N_3589,N_3242,N_3230);
or U3590 (N_3590,N_3291,N_3384);
and U3591 (N_3591,N_3296,N_3215);
nor U3592 (N_3592,N_3226,N_3295);
or U3593 (N_3593,N_3254,N_3293);
and U3594 (N_3594,N_3322,N_3228);
nor U3595 (N_3595,N_3316,N_3362);
or U3596 (N_3596,N_3289,N_3309);
nor U3597 (N_3597,N_3289,N_3211);
nand U3598 (N_3598,N_3263,N_3351);
xor U3599 (N_3599,N_3388,N_3216);
nand U3600 (N_3600,N_3486,N_3557);
or U3601 (N_3601,N_3527,N_3540);
and U3602 (N_3602,N_3593,N_3442);
and U3603 (N_3603,N_3549,N_3573);
or U3604 (N_3604,N_3520,N_3546);
nand U3605 (N_3605,N_3488,N_3460);
or U3606 (N_3606,N_3476,N_3529);
nand U3607 (N_3607,N_3485,N_3499);
nand U3608 (N_3608,N_3577,N_3487);
and U3609 (N_3609,N_3462,N_3567);
nand U3610 (N_3610,N_3563,N_3532);
nor U3611 (N_3611,N_3430,N_3467);
and U3612 (N_3612,N_3425,N_3587);
nand U3613 (N_3613,N_3490,N_3531);
and U3614 (N_3614,N_3554,N_3582);
nor U3615 (N_3615,N_3451,N_3519);
and U3616 (N_3616,N_3400,N_3579);
nor U3617 (N_3617,N_3436,N_3544);
and U3618 (N_3618,N_3591,N_3433);
or U3619 (N_3619,N_3541,N_3407);
nand U3620 (N_3620,N_3457,N_3585);
or U3621 (N_3621,N_3421,N_3576);
or U3622 (N_3622,N_3470,N_3453);
and U3623 (N_3623,N_3454,N_3592);
nor U3624 (N_3624,N_3583,N_3477);
nor U3625 (N_3625,N_3510,N_3492);
nor U3626 (N_3626,N_3524,N_3501);
or U3627 (N_3627,N_3590,N_3427);
or U3628 (N_3628,N_3459,N_3533);
and U3629 (N_3629,N_3491,N_3575);
or U3630 (N_3630,N_3562,N_3447);
nand U3631 (N_3631,N_3494,N_3571);
nand U3632 (N_3632,N_3560,N_3543);
and U3633 (N_3633,N_3479,N_3414);
nand U3634 (N_3634,N_3535,N_3565);
or U3635 (N_3635,N_3599,N_3581);
nand U3636 (N_3636,N_3422,N_3511);
nor U3637 (N_3637,N_3443,N_3439);
and U3638 (N_3638,N_3555,N_3474);
nor U3639 (N_3639,N_3547,N_3572);
or U3640 (N_3640,N_3420,N_3466);
or U3641 (N_3641,N_3507,N_3437);
and U3642 (N_3642,N_3429,N_3448);
nor U3643 (N_3643,N_3584,N_3536);
nor U3644 (N_3644,N_3440,N_3548);
and U3645 (N_3645,N_3598,N_3500);
and U3646 (N_3646,N_3574,N_3446);
and U3647 (N_3647,N_3495,N_3506);
nand U3648 (N_3648,N_3449,N_3566);
nor U3649 (N_3649,N_3426,N_3435);
or U3650 (N_3650,N_3505,N_3512);
nor U3651 (N_3651,N_3596,N_3509);
and U3652 (N_3652,N_3589,N_3408);
nor U3653 (N_3653,N_3450,N_3406);
and U3654 (N_3654,N_3431,N_3412);
nor U3655 (N_3655,N_3525,N_3502);
or U3656 (N_3656,N_3539,N_3515);
and U3657 (N_3657,N_3482,N_3468);
or U3658 (N_3658,N_3418,N_3415);
nor U3659 (N_3659,N_3434,N_3461);
nor U3660 (N_3660,N_3514,N_3409);
or U3661 (N_3661,N_3538,N_3497);
and U3662 (N_3662,N_3597,N_3402);
or U3663 (N_3663,N_3458,N_3428);
nor U3664 (N_3664,N_3523,N_3516);
nand U3665 (N_3665,N_3595,N_3586);
nand U3666 (N_3666,N_3534,N_3404);
and U3667 (N_3667,N_3551,N_3465);
nand U3668 (N_3668,N_3456,N_3526);
and U3669 (N_3669,N_3556,N_3550);
nand U3670 (N_3670,N_3588,N_3521);
nand U3671 (N_3671,N_3455,N_3475);
nor U3672 (N_3672,N_3545,N_3558);
or U3673 (N_3673,N_3564,N_3405);
or U3674 (N_3674,N_3498,N_3438);
nor U3675 (N_3675,N_3444,N_3578);
or U3676 (N_3676,N_3561,N_3528);
or U3677 (N_3677,N_3594,N_3423);
nand U3678 (N_3678,N_3552,N_3481);
nor U3679 (N_3679,N_3559,N_3493);
nor U3680 (N_3680,N_3441,N_3553);
or U3681 (N_3681,N_3504,N_3463);
or U3682 (N_3682,N_3464,N_3478);
and U3683 (N_3683,N_3472,N_3508);
or U3684 (N_3684,N_3537,N_3480);
nor U3685 (N_3685,N_3469,N_3484);
nand U3686 (N_3686,N_3416,N_3522);
nand U3687 (N_3687,N_3517,N_3569);
nand U3688 (N_3688,N_3518,N_3471);
or U3689 (N_3689,N_3452,N_3413);
nand U3690 (N_3690,N_3580,N_3410);
nor U3691 (N_3691,N_3496,N_3489);
or U3692 (N_3692,N_3530,N_3568);
and U3693 (N_3693,N_3411,N_3473);
nor U3694 (N_3694,N_3503,N_3445);
and U3695 (N_3695,N_3513,N_3432);
or U3696 (N_3696,N_3542,N_3424);
nor U3697 (N_3697,N_3570,N_3483);
nand U3698 (N_3698,N_3401,N_3419);
nand U3699 (N_3699,N_3403,N_3417);
nor U3700 (N_3700,N_3591,N_3420);
nand U3701 (N_3701,N_3495,N_3564);
or U3702 (N_3702,N_3418,N_3400);
nand U3703 (N_3703,N_3431,N_3583);
and U3704 (N_3704,N_3517,N_3507);
nand U3705 (N_3705,N_3423,N_3494);
and U3706 (N_3706,N_3544,N_3419);
or U3707 (N_3707,N_3414,N_3534);
nand U3708 (N_3708,N_3448,N_3501);
nor U3709 (N_3709,N_3432,N_3536);
nand U3710 (N_3710,N_3538,N_3573);
or U3711 (N_3711,N_3552,N_3568);
nand U3712 (N_3712,N_3493,N_3515);
or U3713 (N_3713,N_3567,N_3489);
and U3714 (N_3714,N_3434,N_3432);
nor U3715 (N_3715,N_3466,N_3585);
nor U3716 (N_3716,N_3590,N_3405);
nand U3717 (N_3717,N_3462,N_3404);
or U3718 (N_3718,N_3486,N_3426);
nand U3719 (N_3719,N_3447,N_3479);
and U3720 (N_3720,N_3433,N_3462);
or U3721 (N_3721,N_3523,N_3524);
nor U3722 (N_3722,N_3437,N_3434);
or U3723 (N_3723,N_3510,N_3546);
or U3724 (N_3724,N_3511,N_3508);
nor U3725 (N_3725,N_3401,N_3540);
and U3726 (N_3726,N_3479,N_3478);
nor U3727 (N_3727,N_3505,N_3486);
or U3728 (N_3728,N_3577,N_3504);
nor U3729 (N_3729,N_3480,N_3440);
nand U3730 (N_3730,N_3447,N_3565);
nand U3731 (N_3731,N_3547,N_3455);
or U3732 (N_3732,N_3537,N_3404);
nand U3733 (N_3733,N_3469,N_3406);
nand U3734 (N_3734,N_3560,N_3501);
and U3735 (N_3735,N_3532,N_3531);
and U3736 (N_3736,N_3517,N_3473);
nor U3737 (N_3737,N_3507,N_3493);
nand U3738 (N_3738,N_3594,N_3484);
nor U3739 (N_3739,N_3466,N_3592);
nand U3740 (N_3740,N_3452,N_3465);
and U3741 (N_3741,N_3569,N_3432);
or U3742 (N_3742,N_3427,N_3494);
and U3743 (N_3743,N_3542,N_3440);
and U3744 (N_3744,N_3427,N_3472);
and U3745 (N_3745,N_3451,N_3484);
and U3746 (N_3746,N_3550,N_3537);
or U3747 (N_3747,N_3426,N_3462);
or U3748 (N_3748,N_3560,N_3485);
nor U3749 (N_3749,N_3530,N_3572);
nand U3750 (N_3750,N_3576,N_3424);
nor U3751 (N_3751,N_3435,N_3523);
or U3752 (N_3752,N_3476,N_3469);
nand U3753 (N_3753,N_3443,N_3551);
and U3754 (N_3754,N_3577,N_3583);
nand U3755 (N_3755,N_3453,N_3527);
or U3756 (N_3756,N_3530,N_3552);
nor U3757 (N_3757,N_3467,N_3444);
and U3758 (N_3758,N_3431,N_3424);
nor U3759 (N_3759,N_3591,N_3598);
nand U3760 (N_3760,N_3559,N_3553);
nand U3761 (N_3761,N_3561,N_3403);
nand U3762 (N_3762,N_3431,N_3586);
nand U3763 (N_3763,N_3471,N_3443);
or U3764 (N_3764,N_3578,N_3512);
and U3765 (N_3765,N_3414,N_3571);
and U3766 (N_3766,N_3589,N_3436);
nand U3767 (N_3767,N_3452,N_3551);
nand U3768 (N_3768,N_3573,N_3423);
nor U3769 (N_3769,N_3448,N_3544);
and U3770 (N_3770,N_3550,N_3448);
and U3771 (N_3771,N_3449,N_3510);
nand U3772 (N_3772,N_3467,N_3490);
nor U3773 (N_3773,N_3577,N_3448);
or U3774 (N_3774,N_3584,N_3447);
nand U3775 (N_3775,N_3535,N_3503);
or U3776 (N_3776,N_3559,N_3426);
and U3777 (N_3777,N_3550,N_3528);
nor U3778 (N_3778,N_3476,N_3460);
or U3779 (N_3779,N_3565,N_3457);
nor U3780 (N_3780,N_3518,N_3541);
nand U3781 (N_3781,N_3490,N_3496);
and U3782 (N_3782,N_3544,N_3481);
nand U3783 (N_3783,N_3430,N_3454);
and U3784 (N_3784,N_3558,N_3448);
and U3785 (N_3785,N_3450,N_3495);
or U3786 (N_3786,N_3599,N_3477);
nor U3787 (N_3787,N_3476,N_3583);
and U3788 (N_3788,N_3560,N_3496);
and U3789 (N_3789,N_3531,N_3581);
xor U3790 (N_3790,N_3563,N_3493);
nand U3791 (N_3791,N_3495,N_3545);
or U3792 (N_3792,N_3517,N_3480);
xnor U3793 (N_3793,N_3561,N_3405);
nand U3794 (N_3794,N_3485,N_3492);
and U3795 (N_3795,N_3562,N_3522);
and U3796 (N_3796,N_3539,N_3548);
nor U3797 (N_3797,N_3591,N_3587);
or U3798 (N_3798,N_3404,N_3416);
and U3799 (N_3799,N_3456,N_3508);
nand U3800 (N_3800,N_3605,N_3680);
and U3801 (N_3801,N_3731,N_3638);
and U3802 (N_3802,N_3723,N_3754);
nand U3803 (N_3803,N_3643,N_3603);
or U3804 (N_3804,N_3671,N_3662);
or U3805 (N_3805,N_3792,N_3768);
or U3806 (N_3806,N_3689,N_3631);
or U3807 (N_3807,N_3733,N_3746);
and U3808 (N_3808,N_3741,N_3699);
nand U3809 (N_3809,N_3628,N_3645);
and U3810 (N_3810,N_3737,N_3644);
and U3811 (N_3811,N_3647,N_3751);
nor U3812 (N_3812,N_3614,N_3727);
and U3813 (N_3813,N_3750,N_3637);
nor U3814 (N_3814,N_3778,N_3725);
nor U3815 (N_3815,N_3707,N_3782);
nand U3816 (N_3816,N_3797,N_3715);
nand U3817 (N_3817,N_3774,N_3666);
and U3818 (N_3818,N_3695,N_3613);
or U3819 (N_3819,N_3642,N_3732);
nand U3820 (N_3820,N_3606,N_3757);
and U3821 (N_3821,N_3604,N_3617);
nor U3822 (N_3822,N_3658,N_3787);
or U3823 (N_3823,N_3675,N_3688);
nor U3824 (N_3824,N_3704,N_3677);
or U3825 (N_3825,N_3611,N_3679);
xnor U3826 (N_3826,N_3667,N_3706);
nand U3827 (N_3827,N_3610,N_3678);
or U3828 (N_3828,N_3761,N_3690);
nor U3829 (N_3829,N_3655,N_3608);
and U3830 (N_3830,N_3618,N_3670);
nor U3831 (N_3831,N_3600,N_3619);
or U3832 (N_3832,N_3659,N_3789);
and U3833 (N_3833,N_3629,N_3771);
or U3834 (N_3834,N_3687,N_3626);
nor U3835 (N_3835,N_3669,N_3716);
nor U3836 (N_3836,N_3639,N_3601);
nand U3837 (N_3837,N_3770,N_3758);
and U3838 (N_3838,N_3632,N_3640);
and U3839 (N_3839,N_3747,N_3795);
nor U3840 (N_3840,N_3790,N_3705);
nand U3841 (N_3841,N_3703,N_3788);
and U3842 (N_3842,N_3739,N_3729);
nand U3843 (N_3843,N_3649,N_3785);
or U3844 (N_3844,N_3663,N_3759);
and U3845 (N_3845,N_3624,N_3708);
or U3846 (N_3846,N_3641,N_3749);
nor U3847 (N_3847,N_3625,N_3766);
nor U3848 (N_3848,N_3752,N_3775);
nor U3849 (N_3849,N_3664,N_3657);
nand U3850 (N_3850,N_3620,N_3779);
xnor U3851 (N_3851,N_3630,N_3772);
nor U3852 (N_3852,N_3681,N_3734);
or U3853 (N_3853,N_3694,N_3753);
and U3854 (N_3854,N_3794,N_3665);
nand U3855 (N_3855,N_3701,N_3661);
and U3856 (N_3856,N_3654,N_3738);
or U3857 (N_3857,N_3748,N_3698);
xnor U3858 (N_3858,N_3615,N_3602);
nor U3859 (N_3859,N_3783,N_3686);
nand U3860 (N_3860,N_3636,N_3743);
nand U3861 (N_3861,N_3769,N_3672);
nor U3862 (N_3862,N_3650,N_3653);
and U3863 (N_3863,N_3682,N_3767);
nor U3864 (N_3864,N_3710,N_3683);
and U3865 (N_3865,N_3676,N_3717);
nor U3866 (N_3866,N_3684,N_3773);
or U3867 (N_3867,N_3721,N_3740);
and U3868 (N_3868,N_3634,N_3607);
nor U3869 (N_3869,N_3712,N_3728);
nor U3870 (N_3870,N_3693,N_3616);
nor U3871 (N_3871,N_3623,N_3730);
or U3872 (N_3872,N_3756,N_3622);
nand U3873 (N_3873,N_3777,N_3755);
nor U3874 (N_3874,N_3691,N_3714);
or U3875 (N_3875,N_3744,N_3786);
nor U3876 (N_3876,N_3702,N_3799);
xnor U3877 (N_3877,N_3652,N_3621);
and U3878 (N_3878,N_3745,N_3711);
or U3879 (N_3879,N_3660,N_3763);
and U3880 (N_3880,N_3718,N_3735);
nor U3881 (N_3881,N_3720,N_3791);
nor U3882 (N_3882,N_3656,N_3724);
nand U3883 (N_3883,N_3776,N_3781);
or U3884 (N_3884,N_3742,N_3764);
nand U3885 (N_3885,N_3646,N_3793);
nand U3886 (N_3886,N_3700,N_3648);
nand U3887 (N_3887,N_3784,N_3765);
nor U3888 (N_3888,N_3713,N_3609);
or U3889 (N_3889,N_3633,N_3726);
or U3890 (N_3890,N_3673,N_3692);
nor U3891 (N_3891,N_3719,N_3780);
nand U3892 (N_3892,N_3709,N_3736);
nor U3893 (N_3893,N_3651,N_3627);
nor U3894 (N_3894,N_3796,N_3668);
nor U3895 (N_3895,N_3762,N_3722);
or U3896 (N_3896,N_3760,N_3674);
nand U3897 (N_3897,N_3685,N_3697);
nand U3898 (N_3898,N_3612,N_3635);
or U3899 (N_3899,N_3798,N_3696);
nor U3900 (N_3900,N_3679,N_3704);
nand U3901 (N_3901,N_3713,N_3651);
nor U3902 (N_3902,N_3671,N_3792);
or U3903 (N_3903,N_3625,N_3770);
nor U3904 (N_3904,N_3677,N_3694);
or U3905 (N_3905,N_3634,N_3761);
nand U3906 (N_3906,N_3647,N_3653);
nand U3907 (N_3907,N_3764,N_3690);
and U3908 (N_3908,N_3714,N_3749);
nand U3909 (N_3909,N_3651,N_3621);
nand U3910 (N_3910,N_3710,N_3711);
or U3911 (N_3911,N_3673,N_3779);
or U3912 (N_3912,N_3730,N_3796);
nor U3913 (N_3913,N_3621,N_3695);
nand U3914 (N_3914,N_3796,N_3708);
or U3915 (N_3915,N_3715,N_3693);
and U3916 (N_3916,N_3779,N_3756);
or U3917 (N_3917,N_3651,N_3780);
and U3918 (N_3918,N_3731,N_3732);
or U3919 (N_3919,N_3705,N_3708);
or U3920 (N_3920,N_3764,N_3789);
or U3921 (N_3921,N_3773,N_3675);
and U3922 (N_3922,N_3761,N_3785);
nor U3923 (N_3923,N_3795,N_3724);
or U3924 (N_3924,N_3741,N_3782);
nand U3925 (N_3925,N_3600,N_3681);
nand U3926 (N_3926,N_3742,N_3776);
xor U3927 (N_3927,N_3772,N_3750);
or U3928 (N_3928,N_3677,N_3671);
nor U3929 (N_3929,N_3736,N_3680);
nand U3930 (N_3930,N_3711,N_3744);
or U3931 (N_3931,N_3749,N_3726);
and U3932 (N_3932,N_3637,N_3793);
nor U3933 (N_3933,N_3747,N_3619);
and U3934 (N_3934,N_3712,N_3613);
nand U3935 (N_3935,N_3774,N_3618);
nand U3936 (N_3936,N_3678,N_3748);
nor U3937 (N_3937,N_3629,N_3669);
nand U3938 (N_3938,N_3799,N_3609);
and U3939 (N_3939,N_3716,N_3763);
and U3940 (N_3940,N_3772,N_3617);
nand U3941 (N_3941,N_3727,N_3666);
nor U3942 (N_3942,N_3601,N_3735);
or U3943 (N_3943,N_3769,N_3662);
nand U3944 (N_3944,N_3695,N_3759);
nor U3945 (N_3945,N_3716,N_3741);
nor U3946 (N_3946,N_3729,N_3678);
or U3947 (N_3947,N_3625,N_3767);
nor U3948 (N_3948,N_3735,N_3680);
nor U3949 (N_3949,N_3747,N_3625);
or U3950 (N_3950,N_3757,N_3782);
nand U3951 (N_3951,N_3734,N_3680);
nand U3952 (N_3952,N_3609,N_3604);
nand U3953 (N_3953,N_3771,N_3782);
and U3954 (N_3954,N_3630,N_3681);
or U3955 (N_3955,N_3727,N_3768);
and U3956 (N_3956,N_3681,N_3687);
and U3957 (N_3957,N_3680,N_3647);
or U3958 (N_3958,N_3791,N_3757);
and U3959 (N_3959,N_3751,N_3615);
or U3960 (N_3960,N_3731,N_3769);
or U3961 (N_3961,N_3662,N_3767);
nand U3962 (N_3962,N_3675,N_3626);
nor U3963 (N_3963,N_3697,N_3618);
and U3964 (N_3964,N_3688,N_3703);
nand U3965 (N_3965,N_3684,N_3644);
nand U3966 (N_3966,N_3639,N_3762);
nor U3967 (N_3967,N_3749,N_3653);
and U3968 (N_3968,N_3686,N_3687);
nand U3969 (N_3969,N_3766,N_3772);
nor U3970 (N_3970,N_3684,N_3799);
nor U3971 (N_3971,N_3766,N_3793);
or U3972 (N_3972,N_3650,N_3728);
nand U3973 (N_3973,N_3609,N_3765);
nor U3974 (N_3974,N_3734,N_3672);
nand U3975 (N_3975,N_3673,N_3714);
nor U3976 (N_3976,N_3799,N_3641);
nor U3977 (N_3977,N_3684,N_3769);
and U3978 (N_3978,N_3749,N_3615);
nor U3979 (N_3979,N_3766,N_3729);
nand U3980 (N_3980,N_3771,N_3795);
and U3981 (N_3981,N_3667,N_3679);
nor U3982 (N_3982,N_3646,N_3739);
nor U3983 (N_3983,N_3613,N_3658);
nand U3984 (N_3984,N_3706,N_3726);
nand U3985 (N_3985,N_3677,N_3623);
nor U3986 (N_3986,N_3738,N_3642);
or U3987 (N_3987,N_3797,N_3615);
and U3988 (N_3988,N_3701,N_3736);
nand U3989 (N_3989,N_3670,N_3680);
nand U3990 (N_3990,N_3748,N_3612);
and U3991 (N_3991,N_3726,N_3709);
nand U3992 (N_3992,N_3665,N_3778);
and U3993 (N_3993,N_3774,N_3689);
nor U3994 (N_3994,N_3614,N_3661);
nand U3995 (N_3995,N_3731,N_3712);
nand U3996 (N_3996,N_3753,N_3770);
nor U3997 (N_3997,N_3688,N_3604);
nor U3998 (N_3998,N_3770,N_3739);
nand U3999 (N_3999,N_3717,N_3635);
and U4000 (N_4000,N_3803,N_3950);
nor U4001 (N_4001,N_3975,N_3968);
or U4002 (N_4002,N_3934,N_3992);
nor U4003 (N_4003,N_3874,N_3863);
nand U4004 (N_4004,N_3936,N_3962);
nor U4005 (N_4005,N_3955,N_3849);
and U4006 (N_4006,N_3935,N_3822);
nor U4007 (N_4007,N_3883,N_3991);
and U4008 (N_4008,N_3836,N_3841);
and U4009 (N_4009,N_3825,N_3983);
and U4010 (N_4010,N_3909,N_3930);
and U4011 (N_4011,N_3891,N_3969);
or U4012 (N_4012,N_3818,N_3830);
nor U4013 (N_4013,N_3868,N_3855);
and U4014 (N_4014,N_3900,N_3949);
nor U4015 (N_4015,N_3915,N_3921);
or U4016 (N_4016,N_3903,N_3873);
or U4017 (N_4017,N_3925,N_3929);
nand U4018 (N_4018,N_3954,N_3808);
and U4019 (N_4019,N_3899,N_3990);
nand U4020 (N_4020,N_3882,N_3987);
nor U4021 (N_4021,N_3942,N_3923);
and U4022 (N_4022,N_3911,N_3860);
or U4023 (N_4023,N_3869,N_3848);
nor U4024 (N_4024,N_3959,N_3933);
and U4025 (N_4025,N_3846,N_3888);
and U4026 (N_4026,N_3828,N_3928);
and U4027 (N_4027,N_3813,N_3844);
nor U4028 (N_4028,N_3988,N_3858);
or U4029 (N_4029,N_3958,N_3937);
nor U4030 (N_4030,N_3811,N_3829);
or U4031 (N_4031,N_3941,N_3815);
nor U4032 (N_4032,N_3963,N_3807);
and U4033 (N_4033,N_3993,N_3995);
and U4034 (N_4034,N_3998,N_3943);
or U4035 (N_4035,N_3897,N_3814);
xor U4036 (N_4036,N_3820,N_3812);
and U4037 (N_4037,N_3932,N_3896);
or U4038 (N_4038,N_3997,N_3871);
and U4039 (N_4039,N_3839,N_3852);
xnor U4040 (N_4040,N_3905,N_3878);
or U4041 (N_4041,N_3856,N_3823);
nor U4042 (N_4042,N_3947,N_3981);
nor U4043 (N_4043,N_3977,N_3895);
nand U4044 (N_4044,N_3999,N_3908);
nand U4045 (N_4045,N_3948,N_3979);
or U4046 (N_4046,N_3970,N_3845);
nand U4047 (N_4047,N_3945,N_3837);
and U4048 (N_4048,N_3966,N_3922);
and U4049 (N_4049,N_3879,N_3831);
or U4050 (N_4050,N_3876,N_3952);
or U4051 (N_4051,N_3972,N_3916);
or U4052 (N_4052,N_3980,N_3918);
nand U4053 (N_4053,N_3989,N_3847);
nor U4054 (N_4054,N_3854,N_3939);
nand U4055 (N_4055,N_3843,N_3907);
nor U4056 (N_4056,N_3842,N_3976);
or U4057 (N_4057,N_3940,N_3971);
nor U4058 (N_4058,N_3835,N_3859);
nand U4059 (N_4059,N_3885,N_3890);
or U4060 (N_4060,N_3819,N_3985);
and U4061 (N_4061,N_3924,N_3801);
nor U4062 (N_4062,N_3964,N_3804);
or U4063 (N_4063,N_3838,N_3800);
nand U4064 (N_4064,N_3864,N_3862);
and U4065 (N_4065,N_3861,N_3827);
and U4066 (N_4066,N_3904,N_3978);
nand U4067 (N_4067,N_3994,N_3821);
and U4068 (N_4068,N_3953,N_3894);
nand U4069 (N_4069,N_3809,N_3880);
nand U4070 (N_4070,N_3938,N_3886);
nand U4071 (N_4071,N_3920,N_3957);
or U4072 (N_4072,N_3857,N_3867);
or U4073 (N_4073,N_3802,N_3996);
nand U4074 (N_4074,N_3806,N_3986);
nand U4075 (N_4075,N_3866,N_3917);
and U4076 (N_4076,N_3850,N_3875);
or U4077 (N_4077,N_3912,N_3901);
nand U4078 (N_4078,N_3982,N_3805);
or U4079 (N_4079,N_3919,N_3951);
and U4080 (N_4080,N_3810,N_3898);
nor U4081 (N_4081,N_3967,N_3865);
and U4082 (N_4082,N_3984,N_3824);
nand U4083 (N_4083,N_3817,N_3931);
or U4084 (N_4084,N_3840,N_3902);
nand U4085 (N_4085,N_3960,N_3884);
or U4086 (N_4086,N_3887,N_3973);
nand U4087 (N_4087,N_3961,N_3826);
or U4088 (N_4088,N_3834,N_3889);
nand U4089 (N_4089,N_3892,N_3926);
or U4090 (N_4090,N_3851,N_3974);
nor U4091 (N_4091,N_3914,N_3877);
and U4092 (N_4092,N_3832,N_3870);
or U4093 (N_4093,N_3833,N_3853);
nor U4094 (N_4094,N_3872,N_3906);
or U4095 (N_4095,N_3910,N_3893);
nand U4096 (N_4096,N_3956,N_3946);
or U4097 (N_4097,N_3965,N_3927);
or U4098 (N_4098,N_3913,N_3881);
and U4099 (N_4099,N_3944,N_3816);
and U4100 (N_4100,N_3934,N_3813);
nor U4101 (N_4101,N_3865,N_3954);
nand U4102 (N_4102,N_3939,N_3907);
nand U4103 (N_4103,N_3829,N_3854);
or U4104 (N_4104,N_3969,N_3879);
or U4105 (N_4105,N_3969,N_3995);
nand U4106 (N_4106,N_3891,N_3868);
and U4107 (N_4107,N_3940,N_3831);
or U4108 (N_4108,N_3999,N_3930);
nand U4109 (N_4109,N_3948,N_3841);
nand U4110 (N_4110,N_3974,N_3809);
nor U4111 (N_4111,N_3806,N_3996);
nor U4112 (N_4112,N_3906,N_3885);
and U4113 (N_4113,N_3946,N_3802);
nand U4114 (N_4114,N_3816,N_3994);
nor U4115 (N_4115,N_3800,N_3849);
or U4116 (N_4116,N_3931,N_3930);
nor U4117 (N_4117,N_3992,N_3887);
and U4118 (N_4118,N_3812,N_3867);
or U4119 (N_4119,N_3860,N_3898);
nand U4120 (N_4120,N_3869,N_3978);
and U4121 (N_4121,N_3810,N_3840);
xor U4122 (N_4122,N_3940,N_3907);
nand U4123 (N_4123,N_3891,N_3913);
and U4124 (N_4124,N_3993,N_3983);
nor U4125 (N_4125,N_3970,N_3977);
nor U4126 (N_4126,N_3866,N_3966);
and U4127 (N_4127,N_3959,N_3920);
or U4128 (N_4128,N_3807,N_3943);
and U4129 (N_4129,N_3902,N_3914);
nor U4130 (N_4130,N_3905,N_3821);
nand U4131 (N_4131,N_3855,N_3991);
or U4132 (N_4132,N_3936,N_3943);
nand U4133 (N_4133,N_3907,N_3934);
nand U4134 (N_4134,N_3945,N_3906);
or U4135 (N_4135,N_3981,N_3960);
nor U4136 (N_4136,N_3957,N_3911);
nor U4137 (N_4137,N_3917,N_3833);
and U4138 (N_4138,N_3816,N_3826);
or U4139 (N_4139,N_3902,N_3906);
and U4140 (N_4140,N_3915,N_3845);
nand U4141 (N_4141,N_3885,N_3977);
and U4142 (N_4142,N_3980,N_3920);
or U4143 (N_4143,N_3874,N_3902);
and U4144 (N_4144,N_3854,N_3967);
nor U4145 (N_4145,N_3924,N_3856);
nor U4146 (N_4146,N_3944,N_3865);
or U4147 (N_4147,N_3952,N_3813);
or U4148 (N_4148,N_3984,N_3948);
and U4149 (N_4149,N_3984,N_3992);
nor U4150 (N_4150,N_3864,N_3886);
or U4151 (N_4151,N_3858,N_3888);
nor U4152 (N_4152,N_3838,N_3945);
nor U4153 (N_4153,N_3832,N_3986);
or U4154 (N_4154,N_3862,N_3966);
and U4155 (N_4155,N_3863,N_3857);
and U4156 (N_4156,N_3818,N_3921);
or U4157 (N_4157,N_3876,N_3843);
nor U4158 (N_4158,N_3943,N_3881);
and U4159 (N_4159,N_3965,N_3918);
or U4160 (N_4160,N_3968,N_3952);
nand U4161 (N_4161,N_3842,N_3922);
or U4162 (N_4162,N_3941,N_3903);
xnor U4163 (N_4163,N_3828,N_3995);
nand U4164 (N_4164,N_3955,N_3817);
and U4165 (N_4165,N_3813,N_3953);
and U4166 (N_4166,N_3938,N_3821);
nand U4167 (N_4167,N_3916,N_3819);
nand U4168 (N_4168,N_3867,N_3984);
nor U4169 (N_4169,N_3950,N_3984);
nor U4170 (N_4170,N_3966,N_3809);
nand U4171 (N_4171,N_3824,N_3974);
nor U4172 (N_4172,N_3813,N_3812);
and U4173 (N_4173,N_3818,N_3852);
nand U4174 (N_4174,N_3975,N_3865);
or U4175 (N_4175,N_3864,N_3937);
nand U4176 (N_4176,N_3872,N_3974);
or U4177 (N_4177,N_3870,N_3876);
and U4178 (N_4178,N_3960,N_3815);
nand U4179 (N_4179,N_3840,N_3960);
nor U4180 (N_4180,N_3845,N_3923);
or U4181 (N_4181,N_3990,N_3812);
nor U4182 (N_4182,N_3832,N_3946);
and U4183 (N_4183,N_3837,N_3840);
nand U4184 (N_4184,N_3829,N_3846);
nor U4185 (N_4185,N_3982,N_3855);
nand U4186 (N_4186,N_3869,N_3847);
or U4187 (N_4187,N_3890,N_3939);
nor U4188 (N_4188,N_3890,N_3899);
and U4189 (N_4189,N_3925,N_3904);
or U4190 (N_4190,N_3979,N_3998);
and U4191 (N_4191,N_3982,N_3884);
and U4192 (N_4192,N_3863,N_3893);
or U4193 (N_4193,N_3898,N_3868);
xor U4194 (N_4194,N_3914,N_3874);
and U4195 (N_4195,N_3946,N_3888);
nor U4196 (N_4196,N_3981,N_3879);
and U4197 (N_4197,N_3977,N_3976);
or U4198 (N_4198,N_3939,N_3983);
or U4199 (N_4199,N_3896,N_3824);
nand U4200 (N_4200,N_4130,N_4142);
and U4201 (N_4201,N_4167,N_4110);
or U4202 (N_4202,N_4135,N_4092);
nand U4203 (N_4203,N_4080,N_4084);
nand U4204 (N_4204,N_4045,N_4073);
nand U4205 (N_4205,N_4151,N_4000);
nor U4206 (N_4206,N_4091,N_4197);
or U4207 (N_4207,N_4119,N_4020);
and U4208 (N_4208,N_4006,N_4191);
nand U4209 (N_4209,N_4025,N_4124);
or U4210 (N_4210,N_4164,N_4097);
nor U4211 (N_4211,N_4048,N_4143);
nand U4212 (N_4212,N_4046,N_4004);
nand U4213 (N_4213,N_4137,N_4033);
nand U4214 (N_4214,N_4035,N_4005);
nor U4215 (N_4215,N_4082,N_4052);
or U4216 (N_4216,N_4077,N_4106);
nor U4217 (N_4217,N_4144,N_4180);
nand U4218 (N_4218,N_4121,N_4136);
nand U4219 (N_4219,N_4199,N_4147);
nor U4220 (N_4220,N_4177,N_4050);
nor U4221 (N_4221,N_4002,N_4146);
and U4222 (N_4222,N_4187,N_4026);
or U4223 (N_4223,N_4161,N_4039);
or U4224 (N_4224,N_4064,N_4040);
and U4225 (N_4225,N_4126,N_4175);
or U4226 (N_4226,N_4008,N_4190);
and U4227 (N_4227,N_4015,N_4024);
nor U4228 (N_4228,N_4001,N_4032);
nand U4229 (N_4229,N_4007,N_4043);
nor U4230 (N_4230,N_4059,N_4065);
nand U4231 (N_4231,N_4113,N_4060);
nor U4232 (N_4232,N_4100,N_4163);
or U4233 (N_4233,N_4185,N_4103);
and U4234 (N_4234,N_4122,N_4150);
nand U4235 (N_4235,N_4022,N_4018);
or U4236 (N_4236,N_4049,N_4192);
nand U4237 (N_4237,N_4047,N_4034);
or U4238 (N_4238,N_4105,N_4108);
nand U4239 (N_4239,N_4062,N_4029);
or U4240 (N_4240,N_4078,N_4195);
nor U4241 (N_4241,N_4125,N_4179);
or U4242 (N_4242,N_4074,N_4037);
nand U4243 (N_4243,N_4038,N_4068);
or U4244 (N_4244,N_4087,N_4152);
and U4245 (N_4245,N_4194,N_4154);
nand U4246 (N_4246,N_4042,N_4099);
nor U4247 (N_4247,N_4069,N_4061);
nor U4248 (N_4248,N_4066,N_4117);
or U4249 (N_4249,N_4156,N_4003);
nand U4250 (N_4250,N_4085,N_4019);
or U4251 (N_4251,N_4114,N_4023);
and U4252 (N_4252,N_4071,N_4162);
and U4253 (N_4253,N_4010,N_4056);
xor U4254 (N_4254,N_4123,N_4057);
or U4255 (N_4255,N_4129,N_4182);
and U4256 (N_4256,N_4102,N_4196);
nor U4257 (N_4257,N_4021,N_4094);
or U4258 (N_4258,N_4111,N_4158);
nor U4259 (N_4259,N_4168,N_4083);
nand U4260 (N_4260,N_4149,N_4189);
or U4261 (N_4261,N_4176,N_4159);
and U4262 (N_4262,N_4198,N_4051);
or U4263 (N_4263,N_4090,N_4132);
nor U4264 (N_4264,N_4067,N_4089);
or U4265 (N_4265,N_4184,N_4101);
and U4266 (N_4266,N_4027,N_4139);
nor U4267 (N_4267,N_4169,N_4140);
nor U4268 (N_4268,N_4145,N_4112);
nor U4269 (N_4269,N_4134,N_4041);
and U4270 (N_4270,N_4014,N_4017);
nor U4271 (N_4271,N_4141,N_4173);
and U4272 (N_4272,N_4031,N_4053);
or U4273 (N_4273,N_4095,N_4098);
nor U4274 (N_4274,N_4070,N_4058);
nor U4275 (N_4275,N_4153,N_4079);
nand U4276 (N_4276,N_4171,N_4193);
nor U4277 (N_4277,N_4107,N_4076);
nor U4278 (N_4278,N_4081,N_4186);
or U4279 (N_4279,N_4012,N_4088);
nor U4280 (N_4280,N_4181,N_4166);
or U4281 (N_4281,N_4104,N_4028);
or U4282 (N_4282,N_4115,N_4157);
xor U4283 (N_4283,N_4011,N_4009);
or U4284 (N_4284,N_4160,N_4138);
nor U4285 (N_4285,N_4072,N_4096);
nor U4286 (N_4286,N_4174,N_4131);
or U4287 (N_4287,N_4127,N_4109);
and U4288 (N_4288,N_4116,N_4030);
nand U4289 (N_4289,N_4133,N_4016);
xor U4290 (N_4290,N_4120,N_4063);
nand U4291 (N_4291,N_4086,N_4148);
or U4292 (N_4292,N_4055,N_4044);
or U4293 (N_4293,N_4170,N_4178);
and U4294 (N_4294,N_4165,N_4036);
nor U4295 (N_4295,N_4013,N_4118);
or U4296 (N_4296,N_4128,N_4054);
or U4297 (N_4297,N_4075,N_4155);
nand U4298 (N_4298,N_4183,N_4172);
and U4299 (N_4299,N_4093,N_4188);
nor U4300 (N_4300,N_4018,N_4016);
nor U4301 (N_4301,N_4113,N_4165);
nor U4302 (N_4302,N_4119,N_4063);
and U4303 (N_4303,N_4033,N_4138);
or U4304 (N_4304,N_4068,N_4032);
and U4305 (N_4305,N_4019,N_4110);
nand U4306 (N_4306,N_4160,N_4134);
and U4307 (N_4307,N_4092,N_4115);
nand U4308 (N_4308,N_4123,N_4100);
or U4309 (N_4309,N_4022,N_4150);
nand U4310 (N_4310,N_4060,N_4029);
or U4311 (N_4311,N_4105,N_4137);
or U4312 (N_4312,N_4078,N_4036);
or U4313 (N_4313,N_4091,N_4093);
nor U4314 (N_4314,N_4134,N_4136);
nand U4315 (N_4315,N_4019,N_4060);
and U4316 (N_4316,N_4035,N_4127);
nor U4317 (N_4317,N_4029,N_4016);
nor U4318 (N_4318,N_4081,N_4058);
nor U4319 (N_4319,N_4015,N_4093);
nor U4320 (N_4320,N_4090,N_4043);
nor U4321 (N_4321,N_4021,N_4148);
nor U4322 (N_4322,N_4032,N_4028);
nand U4323 (N_4323,N_4036,N_4084);
nand U4324 (N_4324,N_4000,N_4043);
nand U4325 (N_4325,N_4027,N_4076);
nor U4326 (N_4326,N_4008,N_4125);
and U4327 (N_4327,N_4118,N_4185);
and U4328 (N_4328,N_4193,N_4080);
and U4329 (N_4329,N_4156,N_4084);
nand U4330 (N_4330,N_4130,N_4137);
and U4331 (N_4331,N_4029,N_4039);
nand U4332 (N_4332,N_4107,N_4003);
nand U4333 (N_4333,N_4012,N_4031);
or U4334 (N_4334,N_4032,N_4152);
or U4335 (N_4335,N_4047,N_4172);
and U4336 (N_4336,N_4152,N_4178);
nor U4337 (N_4337,N_4085,N_4182);
nand U4338 (N_4338,N_4059,N_4152);
nand U4339 (N_4339,N_4078,N_4015);
nor U4340 (N_4340,N_4022,N_4048);
nand U4341 (N_4341,N_4191,N_4118);
or U4342 (N_4342,N_4010,N_4003);
or U4343 (N_4343,N_4196,N_4147);
nor U4344 (N_4344,N_4126,N_4119);
and U4345 (N_4345,N_4053,N_4159);
nor U4346 (N_4346,N_4095,N_4051);
nor U4347 (N_4347,N_4143,N_4104);
nor U4348 (N_4348,N_4177,N_4154);
or U4349 (N_4349,N_4179,N_4050);
nand U4350 (N_4350,N_4138,N_4191);
or U4351 (N_4351,N_4184,N_4182);
and U4352 (N_4352,N_4186,N_4021);
nor U4353 (N_4353,N_4168,N_4123);
nor U4354 (N_4354,N_4110,N_4157);
nand U4355 (N_4355,N_4034,N_4100);
nor U4356 (N_4356,N_4062,N_4072);
nor U4357 (N_4357,N_4146,N_4182);
nand U4358 (N_4358,N_4133,N_4141);
nand U4359 (N_4359,N_4186,N_4076);
nand U4360 (N_4360,N_4049,N_4048);
nand U4361 (N_4361,N_4036,N_4197);
nand U4362 (N_4362,N_4158,N_4036);
or U4363 (N_4363,N_4016,N_4005);
nor U4364 (N_4364,N_4119,N_4055);
nor U4365 (N_4365,N_4192,N_4030);
nor U4366 (N_4366,N_4051,N_4171);
and U4367 (N_4367,N_4028,N_4152);
and U4368 (N_4368,N_4039,N_4088);
or U4369 (N_4369,N_4083,N_4094);
and U4370 (N_4370,N_4036,N_4096);
and U4371 (N_4371,N_4101,N_4043);
nor U4372 (N_4372,N_4103,N_4083);
nand U4373 (N_4373,N_4039,N_4142);
nand U4374 (N_4374,N_4132,N_4189);
and U4375 (N_4375,N_4178,N_4089);
and U4376 (N_4376,N_4163,N_4089);
and U4377 (N_4377,N_4083,N_4020);
nor U4378 (N_4378,N_4007,N_4143);
nand U4379 (N_4379,N_4045,N_4174);
or U4380 (N_4380,N_4165,N_4074);
nand U4381 (N_4381,N_4059,N_4184);
or U4382 (N_4382,N_4140,N_4077);
and U4383 (N_4383,N_4077,N_4195);
or U4384 (N_4384,N_4177,N_4049);
nand U4385 (N_4385,N_4014,N_4008);
nor U4386 (N_4386,N_4068,N_4077);
nand U4387 (N_4387,N_4157,N_4046);
nor U4388 (N_4388,N_4011,N_4115);
and U4389 (N_4389,N_4147,N_4110);
nand U4390 (N_4390,N_4185,N_4090);
nor U4391 (N_4391,N_4122,N_4033);
or U4392 (N_4392,N_4046,N_4006);
or U4393 (N_4393,N_4052,N_4004);
nand U4394 (N_4394,N_4143,N_4133);
xnor U4395 (N_4395,N_4061,N_4086);
nor U4396 (N_4396,N_4152,N_4089);
or U4397 (N_4397,N_4169,N_4111);
or U4398 (N_4398,N_4047,N_4073);
nand U4399 (N_4399,N_4183,N_4070);
or U4400 (N_4400,N_4294,N_4354);
nand U4401 (N_4401,N_4352,N_4245);
nand U4402 (N_4402,N_4201,N_4217);
nor U4403 (N_4403,N_4297,N_4262);
and U4404 (N_4404,N_4377,N_4225);
nor U4405 (N_4405,N_4360,N_4373);
and U4406 (N_4406,N_4205,N_4235);
or U4407 (N_4407,N_4221,N_4226);
and U4408 (N_4408,N_4241,N_4250);
or U4409 (N_4409,N_4339,N_4345);
nor U4410 (N_4410,N_4394,N_4362);
nand U4411 (N_4411,N_4359,N_4260);
nand U4412 (N_4412,N_4278,N_4223);
or U4413 (N_4413,N_4218,N_4330);
and U4414 (N_4414,N_4295,N_4308);
and U4415 (N_4415,N_4288,N_4307);
and U4416 (N_4416,N_4388,N_4399);
or U4417 (N_4417,N_4349,N_4365);
and U4418 (N_4418,N_4296,N_4385);
and U4419 (N_4419,N_4328,N_4323);
and U4420 (N_4420,N_4267,N_4375);
and U4421 (N_4421,N_4322,N_4243);
nand U4422 (N_4422,N_4222,N_4285);
nor U4423 (N_4423,N_4351,N_4206);
and U4424 (N_4424,N_4334,N_4263);
nand U4425 (N_4425,N_4341,N_4270);
nand U4426 (N_4426,N_4211,N_4287);
nand U4427 (N_4427,N_4369,N_4316);
and U4428 (N_4428,N_4311,N_4280);
and U4429 (N_4429,N_4387,N_4258);
nor U4430 (N_4430,N_4265,N_4212);
nor U4431 (N_4431,N_4396,N_4281);
nor U4432 (N_4432,N_4268,N_4273);
or U4433 (N_4433,N_4363,N_4277);
and U4434 (N_4434,N_4256,N_4283);
or U4435 (N_4435,N_4234,N_4228);
nand U4436 (N_4436,N_4350,N_4272);
nand U4437 (N_4437,N_4395,N_4233);
nand U4438 (N_4438,N_4202,N_4264);
nor U4439 (N_4439,N_4384,N_4276);
or U4440 (N_4440,N_4361,N_4368);
nor U4441 (N_4441,N_4254,N_4238);
xnor U4442 (N_4442,N_4244,N_4237);
or U4443 (N_4443,N_4380,N_4383);
or U4444 (N_4444,N_4397,N_4248);
and U4445 (N_4445,N_4242,N_4253);
nand U4446 (N_4446,N_4340,N_4329);
nand U4447 (N_4447,N_4358,N_4305);
or U4448 (N_4448,N_4210,N_4392);
nand U4449 (N_4449,N_4338,N_4292);
nand U4450 (N_4450,N_4331,N_4324);
nor U4451 (N_4451,N_4304,N_4259);
nor U4452 (N_4452,N_4357,N_4303);
nand U4453 (N_4453,N_4378,N_4333);
nor U4454 (N_4454,N_4208,N_4291);
and U4455 (N_4455,N_4261,N_4213);
nand U4456 (N_4456,N_4236,N_4367);
nand U4457 (N_4457,N_4389,N_4209);
and U4458 (N_4458,N_4372,N_4249);
nand U4459 (N_4459,N_4310,N_4309);
nor U4460 (N_4460,N_4274,N_4301);
nor U4461 (N_4461,N_4216,N_4393);
xnor U4462 (N_4462,N_4300,N_4214);
nor U4463 (N_4463,N_4381,N_4229);
nand U4464 (N_4464,N_4298,N_4227);
nor U4465 (N_4465,N_4335,N_4320);
and U4466 (N_4466,N_4220,N_4370);
and U4467 (N_4467,N_4325,N_4231);
nand U4468 (N_4468,N_4203,N_4318);
nand U4469 (N_4469,N_4290,N_4313);
nor U4470 (N_4470,N_4279,N_4302);
nor U4471 (N_4471,N_4200,N_4364);
nor U4472 (N_4472,N_4269,N_4326);
and U4473 (N_4473,N_4391,N_4284);
and U4474 (N_4474,N_4366,N_4376);
or U4475 (N_4475,N_4255,N_4275);
nor U4476 (N_4476,N_4232,N_4327);
or U4477 (N_4477,N_4299,N_4355);
or U4478 (N_4478,N_4224,N_4315);
nor U4479 (N_4479,N_4282,N_4319);
or U4480 (N_4480,N_4215,N_4371);
nor U4481 (N_4481,N_4379,N_4332);
and U4482 (N_4482,N_4247,N_4219);
or U4483 (N_4483,N_4342,N_4356);
and U4484 (N_4484,N_4252,N_4337);
or U4485 (N_4485,N_4312,N_4204);
nand U4486 (N_4486,N_4306,N_4240);
nand U4487 (N_4487,N_4382,N_4374);
or U4488 (N_4488,N_4293,N_4336);
and U4489 (N_4489,N_4346,N_4390);
or U4490 (N_4490,N_4271,N_4207);
nand U4491 (N_4491,N_4246,N_4348);
nand U4492 (N_4492,N_4344,N_4353);
nand U4493 (N_4493,N_4239,N_4321);
nand U4494 (N_4494,N_4230,N_4266);
nand U4495 (N_4495,N_4317,N_4343);
nand U4496 (N_4496,N_4347,N_4386);
nand U4497 (N_4497,N_4314,N_4286);
nand U4498 (N_4498,N_4257,N_4289);
nor U4499 (N_4499,N_4251,N_4398);
nand U4500 (N_4500,N_4292,N_4350);
xor U4501 (N_4501,N_4383,N_4258);
or U4502 (N_4502,N_4361,N_4319);
nand U4503 (N_4503,N_4261,N_4390);
and U4504 (N_4504,N_4364,N_4379);
nor U4505 (N_4505,N_4353,N_4393);
nor U4506 (N_4506,N_4361,N_4354);
and U4507 (N_4507,N_4284,N_4243);
nand U4508 (N_4508,N_4210,N_4252);
nor U4509 (N_4509,N_4261,N_4219);
or U4510 (N_4510,N_4291,N_4337);
or U4511 (N_4511,N_4283,N_4355);
nor U4512 (N_4512,N_4254,N_4242);
nor U4513 (N_4513,N_4231,N_4265);
and U4514 (N_4514,N_4282,N_4212);
and U4515 (N_4515,N_4342,N_4263);
nand U4516 (N_4516,N_4294,N_4215);
nand U4517 (N_4517,N_4278,N_4273);
nor U4518 (N_4518,N_4227,N_4331);
and U4519 (N_4519,N_4243,N_4236);
nand U4520 (N_4520,N_4217,N_4354);
or U4521 (N_4521,N_4256,N_4251);
and U4522 (N_4522,N_4235,N_4313);
or U4523 (N_4523,N_4380,N_4216);
nand U4524 (N_4524,N_4335,N_4378);
nand U4525 (N_4525,N_4359,N_4288);
and U4526 (N_4526,N_4237,N_4235);
or U4527 (N_4527,N_4251,N_4245);
nor U4528 (N_4528,N_4246,N_4264);
nand U4529 (N_4529,N_4232,N_4240);
and U4530 (N_4530,N_4379,N_4385);
nor U4531 (N_4531,N_4310,N_4220);
nand U4532 (N_4532,N_4234,N_4392);
and U4533 (N_4533,N_4329,N_4322);
nor U4534 (N_4534,N_4264,N_4382);
nor U4535 (N_4535,N_4260,N_4285);
nand U4536 (N_4536,N_4266,N_4394);
nand U4537 (N_4537,N_4341,N_4362);
nor U4538 (N_4538,N_4335,N_4227);
nor U4539 (N_4539,N_4248,N_4256);
or U4540 (N_4540,N_4349,N_4232);
and U4541 (N_4541,N_4210,N_4217);
nand U4542 (N_4542,N_4306,N_4272);
and U4543 (N_4543,N_4203,N_4396);
and U4544 (N_4544,N_4216,N_4348);
and U4545 (N_4545,N_4269,N_4300);
nor U4546 (N_4546,N_4325,N_4304);
nand U4547 (N_4547,N_4277,N_4358);
or U4548 (N_4548,N_4200,N_4222);
or U4549 (N_4549,N_4354,N_4387);
or U4550 (N_4550,N_4284,N_4214);
nor U4551 (N_4551,N_4293,N_4253);
or U4552 (N_4552,N_4222,N_4293);
nor U4553 (N_4553,N_4398,N_4270);
or U4554 (N_4554,N_4378,N_4346);
or U4555 (N_4555,N_4399,N_4378);
nor U4556 (N_4556,N_4391,N_4379);
and U4557 (N_4557,N_4239,N_4354);
nor U4558 (N_4558,N_4350,N_4391);
or U4559 (N_4559,N_4258,N_4365);
nor U4560 (N_4560,N_4301,N_4237);
or U4561 (N_4561,N_4252,N_4377);
nand U4562 (N_4562,N_4219,N_4244);
nor U4563 (N_4563,N_4306,N_4359);
nor U4564 (N_4564,N_4291,N_4284);
nand U4565 (N_4565,N_4304,N_4398);
and U4566 (N_4566,N_4373,N_4346);
nor U4567 (N_4567,N_4345,N_4313);
and U4568 (N_4568,N_4339,N_4233);
or U4569 (N_4569,N_4207,N_4256);
nand U4570 (N_4570,N_4209,N_4307);
nand U4571 (N_4571,N_4321,N_4341);
nor U4572 (N_4572,N_4233,N_4313);
and U4573 (N_4573,N_4324,N_4383);
nand U4574 (N_4574,N_4385,N_4314);
or U4575 (N_4575,N_4398,N_4246);
nand U4576 (N_4576,N_4291,N_4279);
nor U4577 (N_4577,N_4382,N_4386);
and U4578 (N_4578,N_4377,N_4357);
nand U4579 (N_4579,N_4251,N_4319);
and U4580 (N_4580,N_4234,N_4341);
or U4581 (N_4581,N_4331,N_4355);
nand U4582 (N_4582,N_4230,N_4362);
and U4583 (N_4583,N_4218,N_4372);
or U4584 (N_4584,N_4399,N_4266);
or U4585 (N_4585,N_4200,N_4321);
nor U4586 (N_4586,N_4254,N_4287);
or U4587 (N_4587,N_4307,N_4316);
nand U4588 (N_4588,N_4361,N_4268);
nor U4589 (N_4589,N_4375,N_4275);
and U4590 (N_4590,N_4313,N_4227);
and U4591 (N_4591,N_4241,N_4280);
nor U4592 (N_4592,N_4377,N_4338);
or U4593 (N_4593,N_4254,N_4207);
nand U4594 (N_4594,N_4375,N_4300);
nand U4595 (N_4595,N_4224,N_4289);
and U4596 (N_4596,N_4226,N_4219);
and U4597 (N_4597,N_4351,N_4305);
nor U4598 (N_4598,N_4312,N_4346);
or U4599 (N_4599,N_4224,N_4266);
or U4600 (N_4600,N_4446,N_4584);
and U4601 (N_4601,N_4411,N_4413);
nor U4602 (N_4602,N_4572,N_4580);
and U4603 (N_4603,N_4432,N_4594);
and U4604 (N_4604,N_4467,N_4571);
or U4605 (N_4605,N_4478,N_4473);
and U4606 (N_4606,N_4483,N_4425);
or U4607 (N_4607,N_4477,N_4490);
and U4608 (N_4608,N_4420,N_4451);
or U4609 (N_4609,N_4585,N_4564);
nor U4610 (N_4610,N_4547,N_4579);
nand U4611 (N_4611,N_4439,N_4530);
nor U4612 (N_4612,N_4575,N_4592);
and U4613 (N_4613,N_4501,N_4402);
or U4614 (N_4614,N_4559,N_4442);
nor U4615 (N_4615,N_4489,N_4441);
and U4616 (N_4616,N_4534,N_4498);
nor U4617 (N_4617,N_4505,N_4454);
or U4618 (N_4618,N_4544,N_4521);
nor U4619 (N_4619,N_4458,N_4511);
and U4620 (N_4620,N_4496,N_4428);
nand U4621 (N_4621,N_4497,N_4408);
nor U4622 (N_4622,N_4515,N_4405);
or U4623 (N_4623,N_4465,N_4485);
nand U4624 (N_4624,N_4563,N_4593);
nor U4625 (N_4625,N_4598,N_4470);
nor U4626 (N_4626,N_4416,N_4461);
nand U4627 (N_4627,N_4596,N_4565);
nor U4628 (N_4628,N_4509,N_4510);
nand U4629 (N_4629,N_4436,N_4401);
or U4630 (N_4630,N_4551,N_4576);
and U4631 (N_4631,N_4591,N_4536);
and U4632 (N_4632,N_4526,N_4537);
nand U4633 (N_4633,N_4476,N_4586);
nor U4634 (N_4634,N_4421,N_4430);
nand U4635 (N_4635,N_4403,N_4545);
or U4636 (N_4636,N_4406,N_4508);
nor U4637 (N_4637,N_4414,N_4494);
and U4638 (N_4638,N_4480,N_4456);
nand U4639 (N_4639,N_4589,N_4469);
or U4640 (N_4640,N_4459,N_4427);
nand U4641 (N_4641,N_4460,N_4455);
nand U4642 (N_4642,N_4529,N_4475);
and U4643 (N_4643,N_4434,N_4499);
and U4644 (N_4644,N_4527,N_4440);
or U4645 (N_4645,N_4502,N_4588);
and U4646 (N_4646,N_4532,N_4525);
and U4647 (N_4647,N_4518,N_4562);
or U4648 (N_4648,N_4554,N_4520);
and U4649 (N_4649,N_4541,N_4558);
nand U4650 (N_4650,N_4561,N_4472);
and U4651 (N_4651,N_4512,N_4409);
nor U4652 (N_4652,N_4404,N_4550);
xor U4653 (N_4653,N_4443,N_4597);
xnor U4654 (N_4654,N_4433,N_4552);
nor U4655 (N_4655,N_4542,N_4418);
nand U4656 (N_4656,N_4448,N_4500);
or U4657 (N_4657,N_4438,N_4531);
nand U4658 (N_4658,N_4484,N_4555);
nor U4659 (N_4659,N_4410,N_4516);
nor U4660 (N_4660,N_4517,N_4493);
and U4661 (N_4661,N_4549,N_4435);
nor U4662 (N_4662,N_4444,N_4417);
nor U4663 (N_4663,N_4587,N_4569);
nor U4664 (N_4664,N_4538,N_4577);
or U4665 (N_4665,N_4445,N_4487);
nand U4666 (N_4666,N_4415,N_4422);
and U4667 (N_4667,N_4453,N_4546);
nor U4668 (N_4668,N_4429,N_4486);
and U4669 (N_4669,N_4424,N_4447);
nor U4670 (N_4670,N_4570,N_4514);
or U4671 (N_4671,N_4513,N_4507);
nand U4672 (N_4672,N_4578,N_4407);
nor U4673 (N_4673,N_4419,N_4573);
or U4674 (N_4674,N_4582,N_4599);
nor U4675 (N_4675,N_4495,N_4426);
and U4676 (N_4676,N_4457,N_4548);
nand U4677 (N_4677,N_4412,N_4479);
and U4678 (N_4678,N_4583,N_4540);
and U4679 (N_4679,N_4503,N_4522);
or U4680 (N_4680,N_4450,N_4560);
nand U4681 (N_4681,N_4528,N_4533);
or U4682 (N_4682,N_4535,N_4581);
nand U4683 (N_4683,N_4567,N_4590);
xor U4684 (N_4684,N_4423,N_4464);
and U4685 (N_4685,N_4474,N_4491);
and U4686 (N_4686,N_4482,N_4539);
and U4687 (N_4687,N_4566,N_4466);
or U4688 (N_4688,N_4431,N_4488);
nor U4689 (N_4689,N_4468,N_4543);
or U4690 (N_4690,N_4471,N_4481);
xnor U4691 (N_4691,N_4553,N_4523);
xnor U4692 (N_4692,N_4574,N_4556);
nor U4693 (N_4693,N_4462,N_4524);
and U4694 (N_4694,N_4568,N_4492);
nand U4695 (N_4695,N_4506,N_4437);
nor U4696 (N_4696,N_4449,N_4463);
or U4697 (N_4697,N_4519,N_4504);
and U4698 (N_4698,N_4557,N_4400);
and U4699 (N_4699,N_4452,N_4595);
and U4700 (N_4700,N_4474,N_4433);
and U4701 (N_4701,N_4598,N_4506);
nand U4702 (N_4702,N_4535,N_4449);
nor U4703 (N_4703,N_4502,N_4449);
nand U4704 (N_4704,N_4524,N_4473);
and U4705 (N_4705,N_4493,N_4465);
and U4706 (N_4706,N_4581,N_4518);
and U4707 (N_4707,N_4448,N_4466);
nor U4708 (N_4708,N_4416,N_4460);
nor U4709 (N_4709,N_4454,N_4571);
and U4710 (N_4710,N_4539,N_4522);
nand U4711 (N_4711,N_4566,N_4483);
and U4712 (N_4712,N_4551,N_4410);
and U4713 (N_4713,N_4474,N_4526);
or U4714 (N_4714,N_4573,N_4556);
or U4715 (N_4715,N_4443,N_4464);
or U4716 (N_4716,N_4421,N_4582);
xor U4717 (N_4717,N_4412,N_4559);
and U4718 (N_4718,N_4504,N_4567);
or U4719 (N_4719,N_4406,N_4431);
or U4720 (N_4720,N_4467,N_4524);
nor U4721 (N_4721,N_4459,N_4575);
nand U4722 (N_4722,N_4489,N_4539);
or U4723 (N_4723,N_4546,N_4590);
nor U4724 (N_4724,N_4443,N_4412);
nand U4725 (N_4725,N_4523,N_4564);
nor U4726 (N_4726,N_4522,N_4545);
or U4727 (N_4727,N_4557,N_4413);
nor U4728 (N_4728,N_4512,N_4573);
and U4729 (N_4729,N_4497,N_4588);
or U4730 (N_4730,N_4528,N_4569);
nand U4731 (N_4731,N_4545,N_4437);
nand U4732 (N_4732,N_4423,N_4597);
nand U4733 (N_4733,N_4441,N_4453);
nand U4734 (N_4734,N_4529,N_4444);
and U4735 (N_4735,N_4504,N_4430);
nand U4736 (N_4736,N_4500,N_4564);
and U4737 (N_4737,N_4460,N_4515);
nor U4738 (N_4738,N_4429,N_4520);
and U4739 (N_4739,N_4510,N_4595);
and U4740 (N_4740,N_4429,N_4432);
or U4741 (N_4741,N_4521,N_4586);
or U4742 (N_4742,N_4526,N_4467);
nor U4743 (N_4743,N_4438,N_4471);
nor U4744 (N_4744,N_4590,N_4597);
nor U4745 (N_4745,N_4443,N_4570);
nor U4746 (N_4746,N_4553,N_4543);
or U4747 (N_4747,N_4446,N_4435);
nor U4748 (N_4748,N_4463,N_4597);
or U4749 (N_4749,N_4504,N_4568);
nor U4750 (N_4750,N_4426,N_4517);
nor U4751 (N_4751,N_4512,N_4550);
and U4752 (N_4752,N_4419,N_4592);
or U4753 (N_4753,N_4574,N_4444);
and U4754 (N_4754,N_4546,N_4541);
nor U4755 (N_4755,N_4514,N_4440);
nand U4756 (N_4756,N_4570,N_4528);
nand U4757 (N_4757,N_4595,N_4435);
nand U4758 (N_4758,N_4545,N_4484);
nand U4759 (N_4759,N_4529,N_4465);
and U4760 (N_4760,N_4490,N_4577);
and U4761 (N_4761,N_4501,N_4598);
nor U4762 (N_4762,N_4417,N_4465);
and U4763 (N_4763,N_4447,N_4557);
nor U4764 (N_4764,N_4561,N_4424);
nand U4765 (N_4765,N_4581,N_4441);
and U4766 (N_4766,N_4577,N_4582);
and U4767 (N_4767,N_4516,N_4557);
nand U4768 (N_4768,N_4410,N_4567);
nand U4769 (N_4769,N_4523,N_4417);
or U4770 (N_4770,N_4585,N_4533);
nand U4771 (N_4771,N_4516,N_4453);
nand U4772 (N_4772,N_4438,N_4500);
and U4773 (N_4773,N_4415,N_4546);
nor U4774 (N_4774,N_4415,N_4572);
and U4775 (N_4775,N_4511,N_4406);
nand U4776 (N_4776,N_4435,N_4417);
nor U4777 (N_4777,N_4438,N_4586);
nand U4778 (N_4778,N_4482,N_4556);
nor U4779 (N_4779,N_4517,N_4555);
and U4780 (N_4780,N_4541,N_4534);
and U4781 (N_4781,N_4401,N_4485);
and U4782 (N_4782,N_4492,N_4424);
nor U4783 (N_4783,N_4456,N_4530);
nor U4784 (N_4784,N_4403,N_4526);
or U4785 (N_4785,N_4421,N_4584);
and U4786 (N_4786,N_4543,N_4524);
and U4787 (N_4787,N_4465,N_4489);
nor U4788 (N_4788,N_4525,N_4443);
or U4789 (N_4789,N_4596,N_4519);
nor U4790 (N_4790,N_4597,N_4442);
or U4791 (N_4791,N_4594,N_4470);
and U4792 (N_4792,N_4418,N_4492);
or U4793 (N_4793,N_4518,N_4463);
nand U4794 (N_4794,N_4581,N_4455);
and U4795 (N_4795,N_4433,N_4443);
or U4796 (N_4796,N_4596,N_4465);
and U4797 (N_4797,N_4590,N_4471);
nor U4798 (N_4798,N_4481,N_4561);
and U4799 (N_4799,N_4436,N_4517);
and U4800 (N_4800,N_4686,N_4732);
or U4801 (N_4801,N_4753,N_4643);
nand U4802 (N_4802,N_4728,N_4706);
nor U4803 (N_4803,N_4724,N_4720);
nor U4804 (N_4804,N_4759,N_4612);
nor U4805 (N_4805,N_4701,N_4787);
and U4806 (N_4806,N_4719,N_4696);
or U4807 (N_4807,N_4667,N_4655);
and U4808 (N_4808,N_4697,N_4657);
and U4809 (N_4809,N_4650,N_4642);
or U4810 (N_4810,N_4754,N_4631);
nand U4811 (N_4811,N_4646,N_4708);
or U4812 (N_4812,N_4758,N_4752);
nand U4813 (N_4813,N_4718,N_4671);
nor U4814 (N_4814,N_4741,N_4651);
and U4815 (N_4815,N_4633,N_4620);
nor U4816 (N_4816,N_4771,N_4679);
nand U4817 (N_4817,N_4704,N_4665);
or U4818 (N_4818,N_4647,N_4702);
and U4819 (N_4819,N_4674,N_4675);
nor U4820 (N_4820,N_4769,N_4779);
and U4821 (N_4821,N_4727,N_4623);
nand U4822 (N_4822,N_4761,N_4768);
and U4823 (N_4823,N_4621,N_4681);
or U4824 (N_4824,N_4619,N_4630);
nand U4825 (N_4825,N_4694,N_4690);
nor U4826 (N_4826,N_4756,N_4793);
nor U4827 (N_4827,N_4716,N_4640);
nand U4828 (N_4828,N_4774,N_4604);
nor U4829 (N_4829,N_4711,N_4698);
or U4830 (N_4830,N_4618,N_4764);
nor U4831 (N_4831,N_4789,N_4788);
nand U4832 (N_4832,N_4603,N_4760);
nand U4833 (N_4833,N_4743,N_4726);
nor U4834 (N_4834,N_4654,N_4750);
or U4835 (N_4835,N_4742,N_4699);
nor U4836 (N_4836,N_4748,N_4637);
and U4837 (N_4837,N_4682,N_4721);
nand U4838 (N_4838,N_4649,N_4625);
nand U4839 (N_4839,N_4658,N_4795);
or U4840 (N_4840,N_4744,N_4723);
nor U4841 (N_4841,N_4712,N_4629);
and U4842 (N_4842,N_4688,N_4740);
and U4843 (N_4843,N_4783,N_4773);
nor U4844 (N_4844,N_4670,N_4660);
nand U4845 (N_4845,N_4607,N_4736);
or U4846 (N_4846,N_4772,N_4796);
nand U4847 (N_4847,N_4766,N_4669);
nand U4848 (N_4848,N_4762,N_4755);
nand U4849 (N_4849,N_4613,N_4725);
and U4850 (N_4850,N_4678,N_4608);
nor U4851 (N_4851,N_4729,N_4749);
nor U4852 (N_4852,N_4733,N_4715);
nor U4853 (N_4853,N_4745,N_4689);
or U4854 (N_4854,N_4731,N_4684);
or U4855 (N_4855,N_4661,N_4730);
and U4856 (N_4856,N_4757,N_4797);
or U4857 (N_4857,N_4794,N_4710);
nor U4858 (N_4858,N_4644,N_4705);
nand U4859 (N_4859,N_4747,N_4792);
nand U4860 (N_4860,N_4606,N_4735);
and U4861 (N_4861,N_4739,N_4641);
or U4862 (N_4862,N_4778,N_4635);
or U4863 (N_4863,N_4685,N_4663);
nor U4864 (N_4864,N_4648,N_4717);
and U4865 (N_4865,N_4653,N_4799);
nand U4866 (N_4866,N_4770,N_4692);
and U4867 (N_4867,N_4602,N_4765);
and U4868 (N_4868,N_4738,N_4628);
or U4869 (N_4869,N_4737,N_4652);
nor U4870 (N_4870,N_4777,N_4614);
nor U4871 (N_4871,N_4676,N_4751);
or U4872 (N_4872,N_4687,N_4636);
or U4873 (N_4873,N_4605,N_4713);
xnor U4874 (N_4874,N_4683,N_4609);
nand U4875 (N_4875,N_4709,N_4610);
and U4876 (N_4876,N_4722,N_4763);
or U4877 (N_4877,N_4707,N_4786);
nand U4878 (N_4878,N_4798,N_4668);
and U4879 (N_4879,N_4664,N_4677);
nand U4880 (N_4880,N_4672,N_4638);
nor U4881 (N_4881,N_4656,N_4600);
nand U4882 (N_4882,N_4617,N_4624);
nor U4883 (N_4883,N_4611,N_4680);
or U4884 (N_4884,N_4601,N_4693);
or U4885 (N_4885,N_4627,N_4734);
nor U4886 (N_4886,N_4645,N_4622);
or U4887 (N_4887,N_4691,N_4780);
and U4888 (N_4888,N_4703,N_4659);
or U4889 (N_4889,N_4695,N_4626);
nor U4890 (N_4890,N_4616,N_4639);
nor U4891 (N_4891,N_4746,N_4700);
nand U4892 (N_4892,N_4632,N_4785);
nand U4893 (N_4893,N_4784,N_4775);
or U4894 (N_4894,N_4782,N_4781);
nand U4895 (N_4895,N_4673,N_4767);
and U4896 (N_4896,N_4776,N_4634);
nor U4897 (N_4897,N_4790,N_4791);
or U4898 (N_4898,N_4615,N_4662);
or U4899 (N_4899,N_4714,N_4666);
nand U4900 (N_4900,N_4697,N_4681);
or U4901 (N_4901,N_4783,N_4629);
or U4902 (N_4902,N_4796,N_4649);
nand U4903 (N_4903,N_4657,N_4784);
xor U4904 (N_4904,N_4717,N_4683);
nor U4905 (N_4905,N_4799,N_4627);
and U4906 (N_4906,N_4747,N_4618);
nand U4907 (N_4907,N_4673,N_4628);
and U4908 (N_4908,N_4620,N_4654);
or U4909 (N_4909,N_4761,N_4659);
or U4910 (N_4910,N_4755,N_4630);
nor U4911 (N_4911,N_4641,N_4679);
and U4912 (N_4912,N_4651,N_4644);
and U4913 (N_4913,N_4603,N_4685);
nor U4914 (N_4914,N_4734,N_4762);
nor U4915 (N_4915,N_4652,N_4681);
or U4916 (N_4916,N_4696,N_4759);
nand U4917 (N_4917,N_4787,N_4637);
and U4918 (N_4918,N_4600,N_4780);
nand U4919 (N_4919,N_4637,N_4791);
and U4920 (N_4920,N_4698,N_4716);
or U4921 (N_4921,N_4724,N_4649);
and U4922 (N_4922,N_4623,N_4793);
nor U4923 (N_4923,N_4706,N_4789);
xnor U4924 (N_4924,N_4765,N_4705);
or U4925 (N_4925,N_4615,N_4783);
and U4926 (N_4926,N_4709,N_4789);
and U4927 (N_4927,N_4692,N_4745);
and U4928 (N_4928,N_4621,N_4698);
or U4929 (N_4929,N_4632,N_4647);
and U4930 (N_4930,N_4731,N_4640);
and U4931 (N_4931,N_4660,N_4772);
nor U4932 (N_4932,N_4784,N_4709);
and U4933 (N_4933,N_4644,N_4620);
nor U4934 (N_4934,N_4724,N_4725);
nor U4935 (N_4935,N_4732,N_4758);
nor U4936 (N_4936,N_4797,N_4735);
and U4937 (N_4937,N_4645,N_4665);
and U4938 (N_4938,N_4733,N_4755);
nor U4939 (N_4939,N_4698,N_4673);
nand U4940 (N_4940,N_4642,N_4683);
nand U4941 (N_4941,N_4751,N_4741);
nand U4942 (N_4942,N_4736,N_4760);
nor U4943 (N_4943,N_4785,N_4727);
nand U4944 (N_4944,N_4723,N_4674);
xor U4945 (N_4945,N_4787,N_4682);
and U4946 (N_4946,N_4671,N_4633);
nor U4947 (N_4947,N_4765,N_4661);
nor U4948 (N_4948,N_4738,N_4607);
or U4949 (N_4949,N_4649,N_4789);
nor U4950 (N_4950,N_4632,N_4662);
and U4951 (N_4951,N_4785,N_4772);
nand U4952 (N_4952,N_4628,N_4612);
nand U4953 (N_4953,N_4722,N_4732);
nand U4954 (N_4954,N_4753,N_4696);
or U4955 (N_4955,N_4613,N_4668);
nor U4956 (N_4956,N_4695,N_4689);
nand U4957 (N_4957,N_4671,N_4790);
nor U4958 (N_4958,N_4695,N_4750);
or U4959 (N_4959,N_4735,N_4682);
or U4960 (N_4960,N_4642,N_4780);
nand U4961 (N_4961,N_4748,N_4776);
or U4962 (N_4962,N_4630,N_4668);
nand U4963 (N_4963,N_4627,N_4748);
nor U4964 (N_4964,N_4767,N_4611);
and U4965 (N_4965,N_4721,N_4670);
nor U4966 (N_4966,N_4774,N_4779);
nand U4967 (N_4967,N_4656,N_4709);
and U4968 (N_4968,N_4749,N_4744);
nor U4969 (N_4969,N_4663,N_4747);
or U4970 (N_4970,N_4694,N_4641);
nor U4971 (N_4971,N_4786,N_4611);
or U4972 (N_4972,N_4698,N_4646);
or U4973 (N_4973,N_4791,N_4678);
nor U4974 (N_4974,N_4682,N_4658);
nor U4975 (N_4975,N_4757,N_4719);
nor U4976 (N_4976,N_4778,N_4623);
and U4977 (N_4977,N_4721,N_4634);
nand U4978 (N_4978,N_4767,N_4741);
nor U4979 (N_4979,N_4628,N_4761);
nor U4980 (N_4980,N_4687,N_4637);
or U4981 (N_4981,N_4693,N_4633);
nor U4982 (N_4982,N_4749,N_4684);
and U4983 (N_4983,N_4791,N_4776);
nor U4984 (N_4984,N_4673,N_4720);
nand U4985 (N_4985,N_4777,N_4690);
nor U4986 (N_4986,N_4792,N_4666);
nor U4987 (N_4987,N_4676,N_4748);
and U4988 (N_4988,N_4746,N_4727);
nand U4989 (N_4989,N_4610,N_4711);
and U4990 (N_4990,N_4794,N_4674);
or U4991 (N_4991,N_4634,N_4757);
nand U4992 (N_4992,N_4722,N_4630);
nand U4993 (N_4993,N_4695,N_4711);
and U4994 (N_4994,N_4680,N_4770);
nand U4995 (N_4995,N_4682,N_4764);
nand U4996 (N_4996,N_4620,N_4696);
nor U4997 (N_4997,N_4782,N_4702);
and U4998 (N_4998,N_4694,N_4624);
nand U4999 (N_4999,N_4741,N_4734);
nor UO_0 (O_0,N_4990,N_4999);
nand UO_1 (O_1,N_4929,N_4989);
nand UO_2 (O_2,N_4832,N_4905);
nand UO_3 (O_3,N_4970,N_4824);
and UO_4 (O_4,N_4850,N_4925);
and UO_5 (O_5,N_4831,N_4977);
or UO_6 (O_6,N_4968,N_4984);
and UO_7 (O_7,N_4888,N_4963);
and UO_8 (O_8,N_4872,N_4947);
nand UO_9 (O_9,N_4852,N_4950);
or UO_10 (O_10,N_4954,N_4897);
or UO_11 (O_11,N_4843,N_4960);
nand UO_12 (O_12,N_4800,N_4955);
nor UO_13 (O_13,N_4879,N_4933);
nor UO_14 (O_14,N_4978,N_4875);
and UO_15 (O_15,N_4874,N_4961);
and UO_16 (O_16,N_4932,N_4986);
nand UO_17 (O_17,N_4987,N_4823);
nand UO_18 (O_18,N_4869,N_4944);
and UO_19 (O_19,N_4939,N_4935);
and UO_20 (O_20,N_4991,N_4847);
nand UO_21 (O_21,N_4808,N_4949);
nand UO_22 (O_22,N_4856,N_4959);
nor UO_23 (O_23,N_4878,N_4916);
and UO_24 (O_24,N_4828,N_4833);
or UO_25 (O_25,N_4988,N_4862);
and UO_26 (O_26,N_4965,N_4851);
nand UO_27 (O_27,N_4857,N_4868);
and UO_28 (O_28,N_4973,N_4863);
or UO_29 (O_29,N_4845,N_4890);
and UO_30 (O_30,N_4972,N_4894);
nand UO_31 (O_31,N_4956,N_4880);
and UO_32 (O_32,N_4899,N_4817);
nand UO_33 (O_33,N_4957,N_4861);
or UO_34 (O_34,N_4951,N_4952);
nor UO_35 (O_35,N_4865,N_4809);
nand UO_36 (O_36,N_4853,N_4962);
or UO_37 (O_37,N_4964,N_4811);
or UO_38 (O_38,N_4901,N_4889);
nor UO_39 (O_39,N_4994,N_4837);
and UO_40 (O_40,N_4806,N_4822);
nor UO_41 (O_41,N_4941,N_4923);
or UO_42 (O_42,N_4814,N_4815);
and UO_43 (O_43,N_4945,N_4909);
or UO_44 (O_44,N_4807,N_4835);
or UO_45 (O_45,N_4915,N_4971);
and UO_46 (O_46,N_4882,N_4820);
or UO_47 (O_47,N_4854,N_4805);
or UO_48 (O_48,N_4911,N_4810);
and UO_49 (O_49,N_4934,N_4836);
and UO_50 (O_50,N_4848,N_4921);
nor UO_51 (O_51,N_4948,N_4849);
nand UO_52 (O_52,N_4887,N_4922);
or UO_53 (O_53,N_4803,N_4884);
or UO_54 (O_54,N_4981,N_4967);
and UO_55 (O_55,N_4895,N_4919);
and UO_56 (O_56,N_4844,N_4883);
nand UO_57 (O_57,N_4812,N_4896);
and UO_58 (O_58,N_4906,N_4937);
nand UO_59 (O_59,N_4886,N_4827);
and UO_60 (O_60,N_4969,N_4930);
and UO_61 (O_61,N_4859,N_4900);
or UO_62 (O_62,N_4936,N_4910);
or UO_63 (O_63,N_4855,N_4928);
and UO_64 (O_64,N_4873,N_4931);
or UO_65 (O_65,N_4892,N_4864);
nand UO_66 (O_66,N_4871,N_4943);
and UO_67 (O_67,N_4993,N_4966);
or UO_68 (O_68,N_4942,N_4913);
or UO_69 (O_69,N_4876,N_4842);
nor UO_70 (O_70,N_4924,N_4996);
nand UO_71 (O_71,N_4997,N_4983);
nor UO_72 (O_72,N_4881,N_4825);
nand UO_73 (O_73,N_4870,N_4946);
nor UO_74 (O_74,N_4885,N_4914);
nand UO_75 (O_75,N_4953,N_4877);
nor UO_76 (O_76,N_4912,N_4834);
or UO_77 (O_77,N_4907,N_4867);
nand UO_78 (O_78,N_4958,N_4938);
and UO_79 (O_79,N_4918,N_4940);
and UO_80 (O_80,N_4830,N_4813);
and UO_81 (O_81,N_4927,N_4839);
and UO_82 (O_82,N_4891,N_4908);
and UO_83 (O_83,N_4829,N_4976);
nor UO_84 (O_84,N_4926,N_4985);
or UO_85 (O_85,N_4975,N_4802);
and UO_86 (O_86,N_4821,N_4904);
nor UO_87 (O_87,N_4816,N_4818);
nor UO_88 (O_88,N_4840,N_4920);
xor UO_89 (O_89,N_4903,N_4838);
nand UO_90 (O_90,N_4804,N_4992);
and UO_91 (O_91,N_4858,N_4801);
or UO_92 (O_92,N_4866,N_4998);
nand UO_93 (O_93,N_4893,N_4846);
or UO_94 (O_94,N_4898,N_4819);
and UO_95 (O_95,N_4974,N_4980);
and UO_96 (O_96,N_4995,N_4841);
nor UO_97 (O_97,N_4917,N_4860);
and UO_98 (O_98,N_4979,N_4902);
nand UO_99 (O_99,N_4826,N_4982);
xor UO_100 (O_100,N_4989,N_4937);
and UO_101 (O_101,N_4950,N_4805);
nand UO_102 (O_102,N_4941,N_4990);
nor UO_103 (O_103,N_4879,N_4924);
xor UO_104 (O_104,N_4972,N_4815);
nand UO_105 (O_105,N_4993,N_4901);
nand UO_106 (O_106,N_4895,N_4943);
nand UO_107 (O_107,N_4965,N_4922);
and UO_108 (O_108,N_4973,N_4983);
nor UO_109 (O_109,N_4852,N_4832);
and UO_110 (O_110,N_4843,N_4942);
nand UO_111 (O_111,N_4899,N_4867);
nand UO_112 (O_112,N_4838,N_4897);
nor UO_113 (O_113,N_4815,N_4986);
or UO_114 (O_114,N_4910,N_4962);
nor UO_115 (O_115,N_4977,N_4902);
nand UO_116 (O_116,N_4971,N_4818);
or UO_117 (O_117,N_4920,N_4913);
nor UO_118 (O_118,N_4972,N_4842);
or UO_119 (O_119,N_4843,N_4883);
and UO_120 (O_120,N_4851,N_4844);
and UO_121 (O_121,N_4824,N_4821);
and UO_122 (O_122,N_4836,N_4886);
nor UO_123 (O_123,N_4934,N_4911);
nand UO_124 (O_124,N_4881,N_4927);
nor UO_125 (O_125,N_4934,N_4850);
or UO_126 (O_126,N_4876,N_4875);
nor UO_127 (O_127,N_4929,N_4982);
and UO_128 (O_128,N_4974,N_4845);
nand UO_129 (O_129,N_4820,N_4995);
or UO_130 (O_130,N_4920,N_4889);
nor UO_131 (O_131,N_4976,N_4982);
or UO_132 (O_132,N_4982,N_4951);
and UO_133 (O_133,N_4803,N_4938);
or UO_134 (O_134,N_4967,N_4934);
nand UO_135 (O_135,N_4811,N_4988);
or UO_136 (O_136,N_4859,N_4843);
and UO_137 (O_137,N_4923,N_4829);
nand UO_138 (O_138,N_4865,N_4893);
and UO_139 (O_139,N_4853,N_4887);
and UO_140 (O_140,N_4956,N_4857);
or UO_141 (O_141,N_4821,N_4831);
nand UO_142 (O_142,N_4936,N_4867);
and UO_143 (O_143,N_4978,N_4936);
nand UO_144 (O_144,N_4858,N_4978);
nor UO_145 (O_145,N_4977,N_4853);
and UO_146 (O_146,N_4852,N_4988);
nand UO_147 (O_147,N_4863,N_4897);
or UO_148 (O_148,N_4975,N_4821);
nor UO_149 (O_149,N_4994,N_4919);
and UO_150 (O_150,N_4906,N_4925);
or UO_151 (O_151,N_4915,N_4839);
or UO_152 (O_152,N_4924,N_4808);
or UO_153 (O_153,N_4934,N_4944);
nand UO_154 (O_154,N_4847,N_4904);
nand UO_155 (O_155,N_4884,N_4942);
and UO_156 (O_156,N_4848,N_4832);
and UO_157 (O_157,N_4975,N_4847);
or UO_158 (O_158,N_4859,N_4985);
and UO_159 (O_159,N_4935,N_4913);
nor UO_160 (O_160,N_4975,N_4916);
and UO_161 (O_161,N_4940,N_4997);
nor UO_162 (O_162,N_4946,N_4971);
and UO_163 (O_163,N_4865,N_4815);
xnor UO_164 (O_164,N_4968,N_4947);
or UO_165 (O_165,N_4942,N_4920);
and UO_166 (O_166,N_4815,N_4923);
and UO_167 (O_167,N_4996,N_4806);
xor UO_168 (O_168,N_4865,N_4958);
and UO_169 (O_169,N_4961,N_4829);
nand UO_170 (O_170,N_4871,N_4910);
or UO_171 (O_171,N_4938,N_4831);
and UO_172 (O_172,N_4958,N_4971);
or UO_173 (O_173,N_4936,N_4856);
nand UO_174 (O_174,N_4982,N_4925);
or UO_175 (O_175,N_4915,N_4867);
nor UO_176 (O_176,N_4821,N_4843);
nor UO_177 (O_177,N_4879,N_4869);
nand UO_178 (O_178,N_4957,N_4855);
nand UO_179 (O_179,N_4917,N_4813);
nand UO_180 (O_180,N_4957,N_4874);
or UO_181 (O_181,N_4939,N_4800);
and UO_182 (O_182,N_4995,N_4990);
nor UO_183 (O_183,N_4973,N_4803);
nor UO_184 (O_184,N_4932,N_4949);
nand UO_185 (O_185,N_4906,N_4939);
nor UO_186 (O_186,N_4856,N_4849);
and UO_187 (O_187,N_4985,N_4832);
and UO_188 (O_188,N_4870,N_4974);
nor UO_189 (O_189,N_4972,N_4995);
or UO_190 (O_190,N_4971,N_4903);
or UO_191 (O_191,N_4801,N_4931);
nand UO_192 (O_192,N_4858,N_4868);
nand UO_193 (O_193,N_4928,N_4927);
nor UO_194 (O_194,N_4827,N_4899);
nand UO_195 (O_195,N_4979,N_4923);
nor UO_196 (O_196,N_4823,N_4805);
nor UO_197 (O_197,N_4918,N_4873);
nand UO_198 (O_198,N_4877,N_4879);
nor UO_199 (O_199,N_4958,N_4905);
nand UO_200 (O_200,N_4905,N_4884);
or UO_201 (O_201,N_4857,N_4850);
or UO_202 (O_202,N_4824,N_4958);
and UO_203 (O_203,N_4801,N_4965);
or UO_204 (O_204,N_4826,N_4923);
and UO_205 (O_205,N_4901,N_4807);
nand UO_206 (O_206,N_4808,N_4822);
nor UO_207 (O_207,N_4955,N_4823);
nor UO_208 (O_208,N_4962,N_4872);
and UO_209 (O_209,N_4852,N_4823);
and UO_210 (O_210,N_4979,N_4894);
nand UO_211 (O_211,N_4980,N_4984);
or UO_212 (O_212,N_4995,N_4921);
nor UO_213 (O_213,N_4826,N_4972);
nand UO_214 (O_214,N_4888,N_4929);
nand UO_215 (O_215,N_4981,N_4835);
nor UO_216 (O_216,N_4980,N_4954);
nand UO_217 (O_217,N_4836,N_4864);
nor UO_218 (O_218,N_4871,N_4838);
nor UO_219 (O_219,N_4818,N_4848);
or UO_220 (O_220,N_4842,N_4877);
or UO_221 (O_221,N_4936,N_4816);
nand UO_222 (O_222,N_4887,N_4947);
or UO_223 (O_223,N_4814,N_4926);
nor UO_224 (O_224,N_4980,N_4852);
nor UO_225 (O_225,N_4967,N_4988);
nor UO_226 (O_226,N_4849,N_4941);
nor UO_227 (O_227,N_4917,N_4952);
or UO_228 (O_228,N_4908,N_4967);
and UO_229 (O_229,N_4968,N_4894);
nand UO_230 (O_230,N_4962,N_4865);
nor UO_231 (O_231,N_4926,N_4958);
nor UO_232 (O_232,N_4979,N_4816);
nor UO_233 (O_233,N_4939,N_4891);
and UO_234 (O_234,N_4831,N_4983);
nor UO_235 (O_235,N_4931,N_4929);
or UO_236 (O_236,N_4831,N_4953);
nand UO_237 (O_237,N_4876,N_4935);
nand UO_238 (O_238,N_4949,N_4989);
nor UO_239 (O_239,N_4974,N_4839);
or UO_240 (O_240,N_4878,N_4821);
and UO_241 (O_241,N_4856,N_4899);
nor UO_242 (O_242,N_4923,N_4894);
and UO_243 (O_243,N_4912,N_4983);
and UO_244 (O_244,N_4936,N_4863);
nor UO_245 (O_245,N_4966,N_4808);
or UO_246 (O_246,N_4885,N_4819);
nand UO_247 (O_247,N_4878,N_4982);
and UO_248 (O_248,N_4973,N_4862);
nor UO_249 (O_249,N_4840,N_4894);
nand UO_250 (O_250,N_4951,N_4975);
nor UO_251 (O_251,N_4999,N_4918);
or UO_252 (O_252,N_4944,N_4941);
or UO_253 (O_253,N_4989,N_4908);
nor UO_254 (O_254,N_4962,N_4939);
and UO_255 (O_255,N_4861,N_4953);
and UO_256 (O_256,N_4925,N_4846);
nand UO_257 (O_257,N_4907,N_4977);
or UO_258 (O_258,N_4855,N_4828);
nor UO_259 (O_259,N_4955,N_4975);
or UO_260 (O_260,N_4886,N_4847);
nor UO_261 (O_261,N_4883,N_4925);
or UO_262 (O_262,N_4938,N_4829);
and UO_263 (O_263,N_4884,N_4808);
nor UO_264 (O_264,N_4806,N_4906);
nor UO_265 (O_265,N_4990,N_4800);
nor UO_266 (O_266,N_4948,N_4854);
nand UO_267 (O_267,N_4883,N_4840);
nand UO_268 (O_268,N_4808,N_4898);
xnor UO_269 (O_269,N_4875,N_4819);
and UO_270 (O_270,N_4834,N_4902);
nand UO_271 (O_271,N_4804,N_4960);
nand UO_272 (O_272,N_4846,N_4901);
nor UO_273 (O_273,N_4923,N_4996);
and UO_274 (O_274,N_4987,N_4817);
nand UO_275 (O_275,N_4807,N_4929);
or UO_276 (O_276,N_4931,N_4995);
and UO_277 (O_277,N_4800,N_4894);
nor UO_278 (O_278,N_4988,N_4945);
or UO_279 (O_279,N_4858,N_4824);
nand UO_280 (O_280,N_4849,N_4845);
and UO_281 (O_281,N_4858,N_4990);
nor UO_282 (O_282,N_4976,N_4984);
nor UO_283 (O_283,N_4853,N_4934);
and UO_284 (O_284,N_4806,N_4927);
nor UO_285 (O_285,N_4819,N_4986);
nand UO_286 (O_286,N_4972,N_4962);
nand UO_287 (O_287,N_4840,N_4927);
nor UO_288 (O_288,N_4985,N_4842);
nand UO_289 (O_289,N_4871,N_4819);
and UO_290 (O_290,N_4875,N_4962);
and UO_291 (O_291,N_4944,N_4800);
nor UO_292 (O_292,N_4967,N_4965);
and UO_293 (O_293,N_4823,N_4962);
and UO_294 (O_294,N_4830,N_4801);
nand UO_295 (O_295,N_4955,N_4801);
nor UO_296 (O_296,N_4917,N_4857);
or UO_297 (O_297,N_4902,N_4980);
nor UO_298 (O_298,N_4804,N_4981);
nand UO_299 (O_299,N_4997,N_4896);
nor UO_300 (O_300,N_4973,N_4964);
or UO_301 (O_301,N_4934,N_4829);
nand UO_302 (O_302,N_4854,N_4937);
and UO_303 (O_303,N_4891,N_4802);
and UO_304 (O_304,N_4888,N_4863);
nor UO_305 (O_305,N_4948,N_4984);
nor UO_306 (O_306,N_4968,N_4852);
or UO_307 (O_307,N_4889,N_4855);
nor UO_308 (O_308,N_4852,N_4822);
nor UO_309 (O_309,N_4885,N_4933);
or UO_310 (O_310,N_4965,N_4802);
nor UO_311 (O_311,N_4896,N_4914);
or UO_312 (O_312,N_4960,N_4876);
or UO_313 (O_313,N_4937,N_4936);
and UO_314 (O_314,N_4890,N_4886);
nor UO_315 (O_315,N_4919,N_4923);
or UO_316 (O_316,N_4859,N_4803);
nand UO_317 (O_317,N_4903,N_4835);
nand UO_318 (O_318,N_4900,N_4994);
and UO_319 (O_319,N_4894,N_4990);
and UO_320 (O_320,N_4965,N_4815);
or UO_321 (O_321,N_4957,N_4989);
nand UO_322 (O_322,N_4875,N_4961);
and UO_323 (O_323,N_4850,N_4808);
nand UO_324 (O_324,N_4895,N_4948);
nor UO_325 (O_325,N_4992,N_4813);
and UO_326 (O_326,N_4880,N_4835);
or UO_327 (O_327,N_4869,N_4877);
or UO_328 (O_328,N_4897,N_4924);
and UO_329 (O_329,N_4943,N_4839);
nor UO_330 (O_330,N_4967,N_4963);
nor UO_331 (O_331,N_4828,N_4915);
nand UO_332 (O_332,N_4822,N_4854);
and UO_333 (O_333,N_4936,N_4853);
and UO_334 (O_334,N_4800,N_4813);
nand UO_335 (O_335,N_4803,N_4897);
nor UO_336 (O_336,N_4930,N_4810);
nor UO_337 (O_337,N_4843,N_4854);
nor UO_338 (O_338,N_4971,N_4808);
nand UO_339 (O_339,N_4827,N_4980);
or UO_340 (O_340,N_4825,N_4991);
and UO_341 (O_341,N_4856,N_4940);
nand UO_342 (O_342,N_4813,N_4863);
and UO_343 (O_343,N_4966,N_4947);
or UO_344 (O_344,N_4834,N_4959);
nor UO_345 (O_345,N_4822,N_4959);
nor UO_346 (O_346,N_4882,N_4943);
nor UO_347 (O_347,N_4929,N_4862);
or UO_348 (O_348,N_4872,N_4826);
or UO_349 (O_349,N_4805,N_4928);
nand UO_350 (O_350,N_4869,N_4953);
and UO_351 (O_351,N_4904,N_4827);
nand UO_352 (O_352,N_4810,N_4855);
nor UO_353 (O_353,N_4956,N_4800);
nor UO_354 (O_354,N_4914,N_4867);
nand UO_355 (O_355,N_4906,N_4972);
or UO_356 (O_356,N_4814,N_4973);
xor UO_357 (O_357,N_4859,N_4801);
or UO_358 (O_358,N_4831,N_4841);
and UO_359 (O_359,N_4970,N_4960);
and UO_360 (O_360,N_4969,N_4800);
nand UO_361 (O_361,N_4955,N_4867);
and UO_362 (O_362,N_4901,N_4845);
xor UO_363 (O_363,N_4908,N_4973);
nand UO_364 (O_364,N_4927,N_4923);
nand UO_365 (O_365,N_4955,N_4970);
xor UO_366 (O_366,N_4961,N_4997);
nand UO_367 (O_367,N_4926,N_4817);
nor UO_368 (O_368,N_4845,N_4807);
and UO_369 (O_369,N_4877,N_4912);
nand UO_370 (O_370,N_4860,N_4811);
nor UO_371 (O_371,N_4979,N_4831);
and UO_372 (O_372,N_4821,N_4871);
and UO_373 (O_373,N_4807,N_4993);
nor UO_374 (O_374,N_4933,N_4953);
nand UO_375 (O_375,N_4956,N_4803);
or UO_376 (O_376,N_4966,N_4973);
and UO_377 (O_377,N_4972,N_4867);
or UO_378 (O_378,N_4869,N_4921);
nor UO_379 (O_379,N_4905,N_4959);
nand UO_380 (O_380,N_4996,N_4959);
nand UO_381 (O_381,N_4987,N_4840);
or UO_382 (O_382,N_4813,N_4935);
nand UO_383 (O_383,N_4892,N_4830);
nor UO_384 (O_384,N_4833,N_4812);
nor UO_385 (O_385,N_4873,N_4976);
nor UO_386 (O_386,N_4840,N_4831);
and UO_387 (O_387,N_4851,N_4966);
nor UO_388 (O_388,N_4844,N_4815);
or UO_389 (O_389,N_4938,N_4964);
or UO_390 (O_390,N_4832,N_4934);
nand UO_391 (O_391,N_4905,N_4887);
nor UO_392 (O_392,N_4986,N_4919);
and UO_393 (O_393,N_4839,N_4841);
nand UO_394 (O_394,N_4954,N_4878);
xnor UO_395 (O_395,N_4852,N_4897);
nor UO_396 (O_396,N_4994,N_4989);
and UO_397 (O_397,N_4847,N_4990);
or UO_398 (O_398,N_4817,N_4954);
or UO_399 (O_399,N_4818,N_4933);
nand UO_400 (O_400,N_4852,N_4937);
or UO_401 (O_401,N_4838,N_4890);
nor UO_402 (O_402,N_4888,N_4893);
nand UO_403 (O_403,N_4903,N_4904);
or UO_404 (O_404,N_4982,N_4894);
or UO_405 (O_405,N_4837,N_4835);
nor UO_406 (O_406,N_4854,N_4875);
nor UO_407 (O_407,N_4812,N_4949);
nand UO_408 (O_408,N_4886,N_4998);
or UO_409 (O_409,N_4983,N_4904);
and UO_410 (O_410,N_4841,N_4881);
and UO_411 (O_411,N_4861,N_4993);
or UO_412 (O_412,N_4970,N_4863);
or UO_413 (O_413,N_4896,N_4804);
and UO_414 (O_414,N_4905,N_4909);
and UO_415 (O_415,N_4803,N_4812);
nor UO_416 (O_416,N_4826,N_4829);
nand UO_417 (O_417,N_4930,N_4865);
nand UO_418 (O_418,N_4875,N_4999);
xor UO_419 (O_419,N_4995,N_4822);
or UO_420 (O_420,N_4862,N_4946);
or UO_421 (O_421,N_4856,N_4962);
nor UO_422 (O_422,N_4941,N_4866);
or UO_423 (O_423,N_4855,N_4876);
nand UO_424 (O_424,N_4980,N_4916);
or UO_425 (O_425,N_4888,N_4961);
nand UO_426 (O_426,N_4964,N_4857);
and UO_427 (O_427,N_4918,N_4858);
and UO_428 (O_428,N_4869,N_4993);
nand UO_429 (O_429,N_4849,N_4937);
and UO_430 (O_430,N_4911,N_4891);
or UO_431 (O_431,N_4872,N_4870);
or UO_432 (O_432,N_4842,N_4830);
and UO_433 (O_433,N_4857,N_4906);
or UO_434 (O_434,N_4925,N_4820);
nor UO_435 (O_435,N_4916,N_4971);
nand UO_436 (O_436,N_4862,N_4844);
nand UO_437 (O_437,N_4980,N_4983);
or UO_438 (O_438,N_4987,N_4972);
nand UO_439 (O_439,N_4892,N_4840);
or UO_440 (O_440,N_4974,N_4981);
nand UO_441 (O_441,N_4928,N_4808);
or UO_442 (O_442,N_4914,N_4814);
and UO_443 (O_443,N_4813,N_4927);
nor UO_444 (O_444,N_4894,N_4863);
and UO_445 (O_445,N_4992,N_4927);
nand UO_446 (O_446,N_4859,N_4851);
or UO_447 (O_447,N_4918,N_4885);
nand UO_448 (O_448,N_4969,N_4935);
or UO_449 (O_449,N_4994,N_4910);
and UO_450 (O_450,N_4895,N_4813);
or UO_451 (O_451,N_4979,N_4966);
nor UO_452 (O_452,N_4856,N_4831);
and UO_453 (O_453,N_4800,N_4878);
or UO_454 (O_454,N_4841,N_4908);
or UO_455 (O_455,N_4993,N_4847);
nand UO_456 (O_456,N_4844,N_4970);
or UO_457 (O_457,N_4953,N_4976);
or UO_458 (O_458,N_4859,N_4867);
and UO_459 (O_459,N_4862,N_4848);
nor UO_460 (O_460,N_4936,N_4833);
and UO_461 (O_461,N_4944,N_4950);
or UO_462 (O_462,N_4800,N_4865);
xnor UO_463 (O_463,N_4837,N_4954);
nor UO_464 (O_464,N_4803,N_4885);
xor UO_465 (O_465,N_4850,N_4927);
nor UO_466 (O_466,N_4936,N_4824);
or UO_467 (O_467,N_4911,N_4989);
nand UO_468 (O_468,N_4924,N_4994);
nand UO_469 (O_469,N_4875,N_4842);
and UO_470 (O_470,N_4947,N_4809);
nand UO_471 (O_471,N_4827,N_4857);
or UO_472 (O_472,N_4848,N_4837);
or UO_473 (O_473,N_4971,N_4822);
or UO_474 (O_474,N_4841,N_4924);
nor UO_475 (O_475,N_4800,N_4850);
or UO_476 (O_476,N_4996,N_4984);
nand UO_477 (O_477,N_4951,N_4853);
or UO_478 (O_478,N_4972,N_4898);
xor UO_479 (O_479,N_4945,N_4940);
nor UO_480 (O_480,N_4809,N_4811);
nor UO_481 (O_481,N_4909,N_4852);
or UO_482 (O_482,N_4998,N_4873);
or UO_483 (O_483,N_4916,N_4988);
or UO_484 (O_484,N_4884,N_4844);
nand UO_485 (O_485,N_4903,N_4858);
and UO_486 (O_486,N_4883,N_4953);
or UO_487 (O_487,N_4932,N_4988);
or UO_488 (O_488,N_4831,N_4923);
nand UO_489 (O_489,N_4907,N_4932);
nor UO_490 (O_490,N_4834,N_4866);
and UO_491 (O_491,N_4863,N_4999);
nand UO_492 (O_492,N_4984,N_4919);
and UO_493 (O_493,N_4843,N_4950);
nand UO_494 (O_494,N_4884,N_4816);
and UO_495 (O_495,N_4814,N_4823);
nor UO_496 (O_496,N_4990,N_4804);
and UO_497 (O_497,N_4870,N_4941);
or UO_498 (O_498,N_4850,N_4928);
and UO_499 (O_499,N_4933,N_4911);
or UO_500 (O_500,N_4839,N_4868);
nor UO_501 (O_501,N_4841,N_4948);
nand UO_502 (O_502,N_4988,N_4834);
and UO_503 (O_503,N_4854,N_4856);
and UO_504 (O_504,N_4832,N_4884);
nor UO_505 (O_505,N_4946,N_4901);
nand UO_506 (O_506,N_4948,N_4980);
and UO_507 (O_507,N_4850,N_4881);
nand UO_508 (O_508,N_4949,N_4963);
or UO_509 (O_509,N_4886,N_4832);
or UO_510 (O_510,N_4929,N_4864);
and UO_511 (O_511,N_4905,N_4928);
nor UO_512 (O_512,N_4859,N_4915);
nand UO_513 (O_513,N_4968,N_4844);
nand UO_514 (O_514,N_4969,N_4947);
or UO_515 (O_515,N_4809,N_4817);
nand UO_516 (O_516,N_4974,N_4876);
and UO_517 (O_517,N_4847,N_4962);
and UO_518 (O_518,N_4800,N_4856);
nor UO_519 (O_519,N_4855,N_4894);
or UO_520 (O_520,N_4805,N_4842);
nand UO_521 (O_521,N_4925,N_4947);
and UO_522 (O_522,N_4934,N_4887);
nand UO_523 (O_523,N_4968,N_4979);
and UO_524 (O_524,N_4829,N_4832);
or UO_525 (O_525,N_4851,N_4835);
or UO_526 (O_526,N_4934,N_4844);
and UO_527 (O_527,N_4801,N_4883);
or UO_528 (O_528,N_4837,N_4960);
nand UO_529 (O_529,N_4834,N_4905);
or UO_530 (O_530,N_4971,N_4994);
nand UO_531 (O_531,N_4954,N_4839);
or UO_532 (O_532,N_4972,N_4805);
or UO_533 (O_533,N_4808,N_4903);
and UO_534 (O_534,N_4955,N_4905);
or UO_535 (O_535,N_4813,N_4824);
and UO_536 (O_536,N_4858,N_4841);
nor UO_537 (O_537,N_4830,N_4918);
nand UO_538 (O_538,N_4997,N_4831);
and UO_539 (O_539,N_4885,N_4837);
or UO_540 (O_540,N_4918,N_4987);
or UO_541 (O_541,N_4922,N_4836);
or UO_542 (O_542,N_4852,N_4876);
and UO_543 (O_543,N_4958,N_4833);
xor UO_544 (O_544,N_4976,N_4874);
nor UO_545 (O_545,N_4986,N_4876);
or UO_546 (O_546,N_4812,N_4843);
and UO_547 (O_547,N_4864,N_4861);
and UO_548 (O_548,N_4998,N_4893);
nand UO_549 (O_549,N_4970,N_4834);
nand UO_550 (O_550,N_4848,N_4915);
or UO_551 (O_551,N_4924,N_4914);
and UO_552 (O_552,N_4845,N_4921);
or UO_553 (O_553,N_4988,N_4933);
or UO_554 (O_554,N_4850,N_4958);
and UO_555 (O_555,N_4859,N_4884);
nand UO_556 (O_556,N_4900,N_4934);
or UO_557 (O_557,N_4951,N_4804);
nand UO_558 (O_558,N_4887,N_4910);
and UO_559 (O_559,N_4893,N_4819);
and UO_560 (O_560,N_4809,N_4837);
nor UO_561 (O_561,N_4987,N_4877);
nor UO_562 (O_562,N_4902,N_4879);
nor UO_563 (O_563,N_4923,N_4847);
or UO_564 (O_564,N_4988,N_4867);
and UO_565 (O_565,N_4833,N_4981);
and UO_566 (O_566,N_4831,N_4918);
nand UO_567 (O_567,N_4837,N_4847);
nor UO_568 (O_568,N_4818,N_4995);
and UO_569 (O_569,N_4877,N_4972);
nand UO_570 (O_570,N_4864,N_4930);
nor UO_571 (O_571,N_4964,N_4950);
and UO_572 (O_572,N_4972,N_4838);
nor UO_573 (O_573,N_4819,N_4955);
nand UO_574 (O_574,N_4918,N_4939);
and UO_575 (O_575,N_4982,N_4887);
nor UO_576 (O_576,N_4949,N_4940);
and UO_577 (O_577,N_4978,N_4948);
nand UO_578 (O_578,N_4855,N_4959);
nand UO_579 (O_579,N_4995,N_4926);
nor UO_580 (O_580,N_4991,N_4832);
or UO_581 (O_581,N_4893,N_4990);
nor UO_582 (O_582,N_4932,N_4831);
nor UO_583 (O_583,N_4956,N_4906);
nand UO_584 (O_584,N_4855,N_4905);
and UO_585 (O_585,N_4916,N_4800);
nor UO_586 (O_586,N_4914,N_4888);
nor UO_587 (O_587,N_4890,N_4999);
xor UO_588 (O_588,N_4841,N_4885);
and UO_589 (O_589,N_4909,N_4811);
nand UO_590 (O_590,N_4887,N_4921);
nor UO_591 (O_591,N_4902,N_4848);
nand UO_592 (O_592,N_4938,N_4965);
or UO_593 (O_593,N_4885,N_4804);
nand UO_594 (O_594,N_4885,N_4822);
or UO_595 (O_595,N_4865,N_4948);
nand UO_596 (O_596,N_4819,N_4815);
and UO_597 (O_597,N_4951,N_4922);
nor UO_598 (O_598,N_4949,N_4958);
nor UO_599 (O_599,N_4983,N_4929);
nor UO_600 (O_600,N_4929,N_4884);
and UO_601 (O_601,N_4862,N_4867);
and UO_602 (O_602,N_4845,N_4955);
xor UO_603 (O_603,N_4932,N_4947);
nand UO_604 (O_604,N_4916,N_4855);
and UO_605 (O_605,N_4963,N_4831);
or UO_606 (O_606,N_4927,N_4967);
and UO_607 (O_607,N_4987,N_4976);
and UO_608 (O_608,N_4994,N_4930);
xnor UO_609 (O_609,N_4932,N_4869);
nor UO_610 (O_610,N_4807,N_4921);
and UO_611 (O_611,N_4933,N_4829);
or UO_612 (O_612,N_4919,N_4937);
and UO_613 (O_613,N_4944,N_4973);
or UO_614 (O_614,N_4976,N_4868);
xor UO_615 (O_615,N_4964,N_4820);
nor UO_616 (O_616,N_4853,N_4889);
or UO_617 (O_617,N_4899,N_4911);
nor UO_618 (O_618,N_4900,N_4860);
nand UO_619 (O_619,N_4856,N_4996);
nand UO_620 (O_620,N_4842,N_4943);
nor UO_621 (O_621,N_4905,N_4946);
or UO_622 (O_622,N_4879,N_4926);
or UO_623 (O_623,N_4850,N_4975);
nand UO_624 (O_624,N_4841,N_4862);
nor UO_625 (O_625,N_4827,N_4885);
nand UO_626 (O_626,N_4817,N_4928);
nor UO_627 (O_627,N_4920,N_4875);
or UO_628 (O_628,N_4947,N_4941);
xnor UO_629 (O_629,N_4831,N_4873);
or UO_630 (O_630,N_4922,N_4821);
nor UO_631 (O_631,N_4819,N_4809);
and UO_632 (O_632,N_4834,N_4867);
or UO_633 (O_633,N_4815,N_4863);
and UO_634 (O_634,N_4893,N_4937);
or UO_635 (O_635,N_4833,N_4826);
and UO_636 (O_636,N_4940,N_4964);
nor UO_637 (O_637,N_4823,N_4862);
and UO_638 (O_638,N_4889,N_4891);
and UO_639 (O_639,N_4963,N_4974);
nand UO_640 (O_640,N_4959,N_4806);
nand UO_641 (O_641,N_4975,N_4875);
nor UO_642 (O_642,N_4809,N_4886);
nand UO_643 (O_643,N_4957,N_4845);
nor UO_644 (O_644,N_4850,N_4899);
nor UO_645 (O_645,N_4979,N_4937);
nor UO_646 (O_646,N_4994,N_4824);
nand UO_647 (O_647,N_4981,N_4875);
and UO_648 (O_648,N_4980,N_4825);
and UO_649 (O_649,N_4980,N_4949);
nand UO_650 (O_650,N_4887,N_4980);
or UO_651 (O_651,N_4982,N_4835);
and UO_652 (O_652,N_4848,N_4906);
nor UO_653 (O_653,N_4813,N_4918);
or UO_654 (O_654,N_4870,N_4807);
nand UO_655 (O_655,N_4946,N_4914);
or UO_656 (O_656,N_4800,N_4897);
and UO_657 (O_657,N_4935,N_4856);
and UO_658 (O_658,N_4941,N_4899);
nor UO_659 (O_659,N_4808,N_4887);
xor UO_660 (O_660,N_4952,N_4834);
nor UO_661 (O_661,N_4898,N_4805);
nor UO_662 (O_662,N_4839,N_4956);
nor UO_663 (O_663,N_4845,N_4884);
and UO_664 (O_664,N_4975,N_4911);
nor UO_665 (O_665,N_4842,N_4927);
or UO_666 (O_666,N_4928,N_4807);
nor UO_667 (O_667,N_4988,N_4826);
nand UO_668 (O_668,N_4801,N_4972);
nand UO_669 (O_669,N_4964,N_4890);
or UO_670 (O_670,N_4931,N_4817);
and UO_671 (O_671,N_4836,N_4850);
nand UO_672 (O_672,N_4916,N_4842);
and UO_673 (O_673,N_4803,N_4894);
nand UO_674 (O_674,N_4990,N_4888);
nor UO_675 (O_675,N_4835,N_4868);
or UO_676 (O_676,N_4920,N_4936);
and UO_677 (O_677,N_4897,N_4883);
or UO_678 (O_678,N_4928,N_4902);
nand UO_679 (O_679,N_4972,N_4904);
nand UO_680 (O_680,N_4816,N_4978);
nand UO_681 (O_681,N_4912,N_4899);
and UO_682 (O_682,N_4864,N_4903);
nand UO_683 (O_683,N_4913,N_4959);
and UO_684 (O_684,N_4875,N_4881);
or UO_685 (O_685,N_4810,N_4929);
nor UO_686 (O_686,N_4994,N_4944);
or UO_687 (O_687,N_4908,N_4862);
nor UO_688 (O_688,N_4831,N_4994);
nor UO_689 (O_689,N_4868,N_4957);
nor UO_690 (O_690,N_4860,N_4972);
or UO_691 (O_691,N_4961,N_4801);
nand UO_692 (O_692,N_4827,N_4846);
nor UO_693 (O_693,N_4923,N_4872);
or UO_694 (O_694,N_4926,N_4951);
nand UO_695 (O_695,N_4817,N_4905);
nand UO_696 (O_696,N_4900,N_4969);
or UO_697 (O_697,N_4883,N_4850);
or UO_698 (O_698,N_4860,N_4946);
nand UO_699 (O_699,N_4891,N_4999);
nand UO_700 (O_700,N_4862,N_4957);
or UO_701 (O_701,N_4881,N_4812);
or UO_702 (O_702,N_4800,N_4843);
nand UO_703 (O_703,N_4819,N_4905);
nor UO_704 (O_704,N_4909,N_4835);
nand UO_705 (O_705,N_4907,N_4949);
nand UO_706 (O_706,N_4964,N_4881);
nand UO_707 (O_707,N_4950,N_4832);
or UO_708 (O_708,N_4914,N_4949);
or UO_709 (O_709,N_4872,N_4873);
nor UO_710 (O_710,N_4999,N_4828);
and UO_711 (O_711,N_4922,N_4997);
and UO_712 (O_712,N_4925,N_4841);
and UO_713 (O_713,N_4993,N_4895);
and UO_714 (O_714,N_4993,N_4842);
nand UO_715 (O_715,N_4985,N_4911);
nor UO_716 (O_716,N_4882,N_4963);
and UO_717 (O_717,N_4857,N_4992);
nor UO_718 (O_718,N_4850,N_4816);
nor UO_719 (O_719,N_4863,N_4945);
nand UO_720 (O_720,N_4853,N_4837);
and UO_721 (O_721,N_4956,N_4882);
nor UO_722 (O_722,N_4877,N_4952);
and UO_723 (O_723,N_4956,N_4823);
and UO_724 (O_724,N_4868,N_4913);
and UO_725 (O_725,N_4964,N_4873);
nor UO_726 (O_726,N_4958,N_4927);
nand UO_727 (O_727,N_4986,N_4987);
and UO_728 (O_728,N_4808,N_4995);
nand UO_729 (O_729,N_4890,N_4892);
or UO_730 (O_730,N_4804,N_4906);
and UO_731 (O_731,N_4886,N_4891);
nand UO_732 (O_732,N_4941,N_4904);
nand UO_733 (O_733,N_4968,N_4915);
and UO_734 (O_734,N_4949,N_4926);
or UO_735 (O_735,N_4938,N_4822);
nand UO_736 (O_736,N_4873,N_4960);
nor UO_737 (O_737,N_4899,N_4848);
or UO_738 (O_738,N_4987,N_4863);
nor UO_739 (O_739,N_4822,N_4960);
nand UO_740 (O_740,N_4909,N_4898);
nor UO_741 (O_741,N_4909,N_4825);
nand UO_742 (O_742,N_4972,N_4963);
or UO_743 (O_743,N_4928,N_4853);
or UO_744 (O_744,N_4855,N_4998);
nor UO_745 (O_745,N_4986,N_4971);
or UO_746 (O_746,N_4976,N_4833);
or UO_747 (O_747,N_4938,N_4888);
nor UO_748 (O_748,N_4960,N_4890);
nor UO_749 (O_749,N_4851,N_4833);
or UO_750 (O_750,N_4818,N_4803);
nor UO_751 (O_751,N_4994,N_4933);
and UO_752 (O_752,N_4848,N_4991);
nand UO_753 (O_753,N_4956,N_4824);
and UO_754 (O_754,N_4811,N_4821);
nor UO_755 (O_755,N_4927,N_4814);
or UO_756 (O_756,N_4865,N_4872);
or UO_757 (O_757,N_4960,N_4877);
or UO_758 (O_758,N_4833,N_4840);
nand UO_759 (O_759,N_4841,N_4826);
nand UO_760 (O_760,N_4992,N_4999);
or UO_761 (O_761,N_4882,N_4847);
nor UO_762 (O_762,N_4986,N_4923);
or UO_763 (O_763,N_4941,N_4999);
nor UO_764 (O_764,N_4937,N_4986);
or UO_765 (O_765,N_4877,N_4926);
and UO_766 (O_766,N_4837,N_4880);
and UO_767 (O_767,N_4987,N_4943);
and UO_768 (O_768,N_4861,N_4808);
nor UO_769 (O_769,N_4918,N_4837);
or UO_770 (O_770,N_4838,N_4847);
nand UO_771 (O_771,N_4883,N_4914);
and UO_772 (O_772,N_4832,N_4834);
nand UO_773 (O_773,N_4986,N_4941);
and UO_774 (O_774,N_4935,N_4872);
and UO_775 (O_775,N_4876,N_4970);
nand UO_776 (O_776,N_4887,N_4825);
and UO_777 (O_777,N_4909,N_4978);
nand UO_778 (O_778,N_4893,N_4999);
nand UO_779 (O_779,N_4801,N_4935);
and UO_780 (O_780,N_4817,N_4874);
nand UO_781 (O_781,N_4936,N_4954);
nand UO_782 (O_782,N_4893,N_4896);
nand UO_783 (O_783,N_4922,N_4947);
nand UO_784 (O_784,N_4954,N_4913);
nand UO_785 (O_785,N_4978,N_4993);
nand UO_786 (O_786,N_4864,N_4990);
nand UO_787 (O_787,N_4963,N_4952);
nor UO_788 (O_788,N_4830,N_4912);
nor UO_789 (O_789,N_4874,N_4835);
nand UO_790 (O_790,N_4881,N_4968);
nor UO_791 (O_791,N_4903,N_4900);
or UO_792 (O_792,N_4997,N_4877);
nor UO_793 (O_793,N_4846,N_4912);
or UO_794 (O_794,N_4884,N_4961);
nand UO_795 (O_795,N_4883,N_4912);
or UO_796 (O_796,N_4945,N_4870);
or UO_797 (O_797,N_4976,N_4825);
nand UO_798 (O_798,N_4819,N_4987);
and UO_799 (O_799,N_4964,N_4879);
nand UO_800 (O_800,N_4827,N_4822);
and UO_801 (O_801,N_4877,N_4871);
and UO_802 (O_802,N_4878,N_4897);
and UO_803 (O_803,N_4867,N_4827);
nor UO_804 (O_804,N_4929,N_4866);
nor UO_805 (O_805,N_4824,N_4914);
or UO_806 (O_806,N_4930,N_4980);
nor UO_807 (O_807,N_4968,N_4847);
nor UO_808 (O_808,N_4863,N_4857);
nor UO_809 (O_809,N_4965,N_4837);
nand UO_810 (O_810,N_4874,N_4861);
or UO_811 (O_811,N_4820,N_4852);
and UO_812 (O_812,N_4867,N_4828);
nand UO_813 (O_813,N_4810,N_4869);
and UO_814 (O_814,N_4836,N_4894);
nand UO_815 (O_815,N_4901,N_4967);
and UO_816 (O_816,N_4935,N_4947);
nand UO_817 (O_817,N_4970,N_4940);
or UO_818 (O_818,N_4965,N_4879);
nand UO_819 (O_819,N_4828,N_4990);
and UO_820 (O_820,N_4949,N_4922);
and UO_821 (O_821,N_4899,N_4843);
nor UO_822 (O_822,N_4899,N_4864);
and UO_823 (O_823,N_4934,N_4816);
nand UO_824 (O_824,N_4848,N_4801);
or UO_825 (O_825,N_4911,N_4908);
nand UO_826 (O_826,N_4996,N_4840);
and UO_827 (O_827,N_4994,N_4850);
nor UO_828 (O_828,N_4866,N_4832);
and UO_829 (O_829,N_4896,N_4811);
or UO_830 (O_830,N_4893,N_4899);
nand UO_831 (O_831,N_4830,N_4993);
and UO_832 (O_832,N_4913,N_4892);
or UO_833 (O_833,N_4830,N_4901);
nor UO_834 (O_834,N_4941,N_4924);
or UO_835 (O_835,N_4948,N_4940);
nor UO_836 (O_836,N_4882,N_4955);
or UO_837 (O_837,N_4942,N_4890);
or UO_838 (O_838,N_4923,N_4860);
nor UO_839 (O_839,N_4811,N_4881);
nor UO_840 (O_840,N_4846,N_4878);
or UO_841 (O_841,N_4910,N_4823);
nor UO_842 (O_842,N_4862,N_4928);
nand UO_843 (O_843,N_4898,N_4923);
or UO_844 (O_844,N_4978,N_4957);
and UO_845 (O_845,N_4915,N_4817);
nand UO_846 (O_846,N_4889,N_4979);
or UO_847 (O_847,N_4968,N_4889);
nor UO_848 (O_848,N_4867,N_4872);
or UO_849 (O_849,N_4817,N_4823);
and UO_850 (O_850,N_4945,N_4865);
and UO_851 (O_851,N_4817,N_4844);
or UO_852 (O_852,N_4805,N_4932);
nor UO_853 (O_853,N_4844,N_4874);
nand UO_854 (O_854,N_4892,N_4869);
nand UO_855 (O_855,N_4827,N_4986);
or UO_856 (O_856,N_4987,N_4929);
nand UO_857 (O_857,N_4805,N_4852);
and UO_858 (O_858,N_4931,N_4820);
nor UO_859 (O_859,N_4853,N_4831);
and UO_860 (O_860,N_4870,N_4940);
and UO_861 (O_861,N_4905,N_4877);
nor UO_862 (O_862,N_4943,N_4827);
nor UO_863 (O_863,N_4879,N_4885);
and UO_864 (O_864,N_4909,N_4984);
nand UO_865 (O_865,N_4971,N_4908);
nor UO_866 (O_866,N_4855,N_4961);
or UO_867 (O_867,N_4919,N_4899);
or UO_868 (O_868,N_4915,N_4914);
and UO_869 (O_869,N_4866,N_4835);
and UO_870 (O_870,N_4965,N_4944);
nand UO_871 (O_871,N_4826,N_4843);
and UO_872 (O_872,N_4936,N_4944);
nor UO_873 (O_873,N_4910,N_4815);
or UO_874 (O_874,N_4889,N_4819);
nand UO_875 (O_875,N_4828,N_4922);
or UO_876 (O_876,N_4814,N_4829);
xnor UO_877 (O_877,N_4859,N_4861);
or UO_878 (O_878,N_4982,N_4958);
and UO_879 (O_879,N_4820,N_4956);
nor UO_880 (O_880,N_4996,N_4905);
nor UO_881 (O_881,N_4925,N_4984);
nor UO_882 (O_882,N_4997,N_4812);
and UO_883 (O_883,N_4995,N_4911);
and UO_884 (O_884,N_4891,N_4946);
nand UO_885 (O_885,N_4927,N_4861);
or UO_886 (O_886,N_4851,N_4837);
or UO_887 (O_887,N_4954,N_4951);
or UO_888 (O_888,N_4839,N_4877);
nand UO_889 (O_889,N_4880,N_4925);
nand UO_890 (O_890,N_4891,N_4873);
or UO_891 (O_891,N_4954,N_4844);
and UO_892 (O_892,N_4994,N_4880);
nor UO_893 (O_893,N_4835,N_4907);
and UO_894 (O_894,N_4892,N_4934);
nand UO_895 (O_895,N_4984,N_4961);
nand UO_896 (O_896,N_4889,N_4938);
and UO_897 (O_897,N_4807,N_4944);
or UO_898 (O_898,N_4935,N_4841);
or UO_899 (O_899,N_4891,N_4896);
nand UO_900 (O_900,N_4909,N_4942);
nand UO_901 (O_901,N_4842,N_4850);
and UO_902 (O_902,N_4996,N_4907);
or UO_903 (O_903,N_4868,N_4819);
and UO_904 (O_904,N_4915,N_4977);
or UO_905 (O_905,N_4823,N_4981);
nand UO_906 (O_906,N_4995,N_4854);
or UO_907 (O_907,N_4957,N_4843);
and UO_908 (O_908,N_4905,N_4847);
nand UO_909 (O_909,N_4831,N_4896);
nor UO_910 (O_910,N_4946,N_4879);
and UO_911 (O_911,N_4861,N_4809);
and UO_912 (O_912,N_4920,N_4891);
nand UO_913 (O_913,N_4844,N_4974);
and UO_914 (O_914,N_4920,N_4838);
and UO_915 (O_915,N_4942,N_4877);
or UO_916 (O_916,N_4916,N_4953);
nand UO_917 (O_917,N_4800,N_4980);
nor UO_918 (O_918,N_4870,N_4923);
or UO_919 (O_919,N_4893,N_4968);
nand UO_920 (O_920,N_4957,N_4838);
nor UO_921 (O_921,N_4892,N_4943);
nor UO_922 (O_922,N_4802,N_4970);
nand UO_923 (O_923,N_4954,N_4876);
nor UO_924 (O_924,N_4941,N_4926);
or UO_925 (O_925,N_4890,N_4998);
and UO_926 (O_926,N_4870,N_4954);
nor UO_927 (O_927,N_4957,N_4851);
or UO_928 (O_928,N_4802,N_4985);
nor UO_929 (O_929,N_4943,N_4804);
or UO_930 (O_930,N_4940,N_4920);
xnor UO_931 (O_931,N_4882,N_4928);
and UO_932 (O_932,N_4815,N_4971);
nand UO_933 (O_933,N_4875,N_4840);
and UO_934 (O_934,N_4876,N_4854);
or UO_935 (O_935,N_4956,N_4888);
and UO_936 (O_936,N_4838,N_4810);
xor UO_937 (O_937,N_4858,N_4810);
or UO_938 (O_938,N_4941,N_4942);
or UO_939 (O_939,N_4857,N_4998);
or UO_940 (O_940,N_4986,N_4829);
nor UO_941 (O_941,N_4934,N_4818);
or UO_942 (O_942,N_4894,N_4824);
xor UO_943 (O_943,N_4910,N_4822);
nor UO_944 (O_944,N_4904,N_4824);
and UO_945 (O_945,N_4811,N_4966);
and UO_946 (O_946,N_4921,N_4844);
or UO_947 (O_947,N_4911,N_4809);
nand UO_948 (O_948,N_4886,N_4932);
nor UO_949 (O_949,N_4845,N_4838);
or UO_950 (O_950,N_4868,N_4986);
nor UO_951 (O_951,N_4923,N_4959);
nand UO_952 (O_952,N_4844,N_4946);
nor UO_953 (O_953,N_4819,N_4839);
nor UO_954 (O_954,N_4874,N_4973);
nand UO_955 (O_955,N_4830,N_4838);
nor UO_956 (O_956,N_4933,N_4837);
nand UO_957 (O_957,N_4891,N_4904);
or UO_958 (O_958,N_4945,N_4893);
nor UO_959 (O_959,N_4930,N_4802);
nand UO_960 (O_960,N_4989,N_4900);
nor UO_961 (O_961,N_4894,N_4930);
nand UO_962 (O_962,N_4815,N_4946);
or UO_963 (O_963,N_4857,N_4845);
or UO_964 (O_964,N_4825,N_4848);
and UO_965 (O_965,N_4981,N_4836);
or UO_966 (O_966,N_4976,N_4971);
xor UO_967 (O_967,N_4879,N_4913);
nor UO_968 (O_968,N_4900,N_4890);
and UO_969 (O_969,N_4854,N_4814);
or UO_970 (O_970,N_4900,N_4875);
or UO_971 (O_971,N_4976,N_4863);
nor UO_972 (O_972,N_4961,N_4989);
or UO_973 (O_973,N_4918,N_4980);
nor UO_974 (O_974,N_4981,N_4818);
and UO_975 (O_975,N_4978,N_4853);
xnor UO_976 (O_976,N_4855,N_4915);
and UO_977 (O_977,N_4928,N_4948);
or UO_978 (O_978,N_4868,N_4941);
or UO_979 (O_979,N_4851,N_4983);
nor UO_980 (O_980,N_4998,N_4992);
nand UO_981 (O_981,N_4908,N_4880);
nor UO_982 (O_982,N_4921,N_4907);
nand UO_983 (O_983,N_4941,N_4916);
nand UO_984 (O_984,N_4942,N_4846);
nor UO_985 (O_985,N_4927,N_4873);
or UO_986 (O_986,N_4856,N_4978);
and UO_987 (O_987,N_4822,N_4884);
nand UO_988 (O_988,N_4990,N_4968);
and UO_989 (O_989,N_4907,N_4979);
nand UO_990 (O_990,N_4883,N_4812);
nand UO_991 (O_991,N_4994,N_4982);
or UO_992 (O_992,N_4897,N_4964);
or UO_993 (O_993,N_4834,N_4977);
nor UO_994 (O_994,N_4922,N_4925);
nor UO_995 (O_995,N_4932,N_4960);
nor UO_996 (O_996,N_4951,N_4809);
nand UO_997 (O_997,N_4980,N_4821);
and UO_998 (O_998,N_4907,N_4801);
or UO_999 (O_999,N_4808,N_4973);
endmodule