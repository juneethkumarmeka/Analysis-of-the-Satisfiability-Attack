module basic_750_5000_1000_25_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_680,In_280);
or U1 (N_1,In_273,In_622);
or U2 (N_2,In_604,In_488);
nor U3 (N_3,In_37,In_748);
nand U4 (N_4,In_608,In_587);
or U5 (N_5,In_29,In_218);
and U6 (N_6,In_695,In_696);
nand U7 (N_7,In_499,In_170);
nor U8 (N_8,In_89,In_114);
and U9 (N_9,In_109,In_50);
or U10 (N_10,In_708,In_405);
nor U11 (N_11,In_683,In_615);
or U12 (N_12,In_589,In_38);
nand U13 (N_13,In_585,In_27);
nor U14 (N_14,In_353,In_34);
and U15 (N_15,In_100,In_289);
and U16 (N_16,In_704,In_621);
and U17 (N_17,In_456,In_466);
nor U18 (N_18,In_199,In_327);
nor U19 (N_19,In_586,In_215);
or U20 (N_20,In_362,In_225);
and U21 (N_21,In_49,In_335);
nand U22 (N_22,In_338,In_549);
xnor U23 (N_23,In_623,In_619);
nor U24 (N_24,In_23,In_560);
nand U25 (N_25,In_40,In_687);
nor U26 (N_26,In_437,In_378);
and U27 (N_27,In_397,In_506);
nor U28 (N_28,In_87,In_337);
nand U29 (N_29,In_270,In_133);
nand U30 (N_30,In_484,In_504);
nor U31 (N_31,In_471,In_173);
or U32 (N_32,In_112,In_33);
nand U33 (N_33,In_415,In_111);
xor U34 (N_34,In_375,In_749);
nand U35 (N_35,In_366,In_737);
nand U36 (N_36,In_276,In_581);
nand U37 (N_37,In_633,In_47);
nor U38 (N_38,In_743,In_71);
and U39 (N_39,In_194,In_438);
nor U40 (N_40,In_599,In_340);
xnor U41 (N_41,In_607,In_56);
or U42 (N_42,In_285,In_107);
xor U43 (N_43,In_511,In_252);
nor U44 (N_44,In_474,In_342);
nand U45 (N_45,In_147,In_446);
and U46 (N_46,In_148,In_283);
nand U47 (N_47,In_277,In_146);
or U48 (N_48,In_52,In_205);
nand U49 (N_49,In_306,In_677);
xnor U50 (N_50,In_125,In_571);
and U51 (N_51,In_16,In_121);
and U52 (N_52,In_541,In_598);
nand U53 (N_53,In_175,In_35);
nor U54 (N_54,In_674,In_428);
or U55 (N_55,In_203,In_126);
or U56 (N_56,In_644,In_162);
xnor U57 (N_57,In_152,In_359);
nor U58 (N_58,In_729,In_236);
nand U59 (N_59,In_99,In_709);
xnor U60 (N_60,In_216,In_408);
xor U61 (N_61,In_97,In_514);
or U62 (N_62,In_63,In_554);
nor U63 (N_63,In_193,In_185);
and U64 (N_64,In_630,In_635);
nand U65 (N_65,In_544,In_217);
xor U66 (N_66,In_245,In_36);
nor U67 (N_67,In_386,In_463);
nand U68 (N_68,In_72,In_518);
nand U69 (N_69,In_640,In_527);
and U70 (N_70,In_449,In_624);
or U71 (N_71,In_235,In_284);
nor U72 (N_72,In_537,In_20);
nand U73 (N_73,In_394,In_41);
nand U74 (N_74,In_361,In_180);
nor U75 (N_75,In_450,In_320);
or U76 (N_76,In_746,In_356);
nor U77 (N_77,In_314,In_742);
xnor U78 (N_78,In_584,In_435);
nor U79 (N_79,In_357,In_32);
xnor U80 (N_80,In_461,In_86);
nand U81 (N_81,In_528,In_460);
or U82 (N_82,In_489,In_578);
xor U83 (N_83,In_740,In_226);
and U84 (N_84,In_200,In_324);
and U85 (N_85,In_564,In_613);
xor U86 (N_86,In_717,In_464);
or U87 (N_87,In_614,In_690);
nor U88 (N_88,In_303,In_331);
and U89 (N_89,In_697,In_81);
or U90 (N_90,In_64,In_715);
nand U91 (N_91,In_457,In_196);
xor U92 (N_92,In_102,In_177);
or U93 (N_93,In_51,In_719);
nand U94 (N_94,In_354,In_430);
and U95 (N_95,In_155,In_264);
and U96 (N_96,In_288,In_591);
or U97 (N_97,In_667,In_151);
and U98 (N_98,In_470,In_583);
or U99 (N_99,In_714,In_547);
xnor U100 (N_100,In_28,In_649);
and U101 (N_101,In_332,In_650);
and U102 (N_102,In_374,In_479);
nand U103 (N_103,In_171,In_57);
nand U104 (N_104,In_90,In_648);
xor U105 (N_105,In_293,In_682);
or U106 (N_106,In_487,In_25);
nand U107 (N_107,In_164,In_316);
or U108 (N_108,In_486,In_684);
nand U109 (N_109,In_31,In_116);
nor U110 (N_110,In_427,In_536);
nor U111 (N_111,In_414,In_381);
nand U112 (N_112,In_592,In_694);
nand U113 (N_113,In_319,In_496);
and U114 (N_114,In_91,In_723);
and U115 (N_115,In_647,In_253);
xor U116 (N_116,In_351,In_383);
nor U117 (N_117,In_576,In_83);
nand U118 (N_118,In_222,In_131);
and U119 (N_119,In_224,In_279);
and U120 (N_120,In_30,In_572);
xor U121 (N_121,In_389,In_521);
or U122 (N_122,In_189,In_418);
and U123 (N_123,In_401,In_7);
xnor U124 (N_124,In_720,In_664);
nand U125 (N_125,In_14,In_653);
nand U126 (N_126,In_500,In_371);
nor U127 (N_127,In_343,In_570);
xnor U128 (N_128,In_485,In_198);
nor U129 (N_129,In_73,In_142);
xnor U130 (N_130,In_78,In_92);
or U131 (N_131,In_294,In_19);
or U132 (N_132,In_601,In_478);
and U133 (N_133,In_655,In_699);
nor U134 (N_134,In_60,In_55);
nor U135 (N_135,In_533,In_241);
and U136 (N_136,In_515,In_75);
xor U137 (N_137,In_272,In_300);
and U138 (N_138,In_439,In_158);
nor U139 (N_139,In_214,In_65);
xnor U140 (N_140,In_588,In_297);
nor U141 (N_141,In_168,In_358);
nor U142 (N_142,In_46,In_594);
xnor U143 (N_143,In_365,In_445);
nor U144 (N_144,In_255,In_642);
xnor U145 (N_145,In_254,In_281);
and U146 (N_146,In_390,In_686);
xnor U147 (N_147,In_3,In_422);
nand U148 (N_148,In_665,In_535);
and U149 (N_149,In_301,In_231);
and U150 (N_150,In_261,In_669);
or U151 (N_151,In_223,In_101);
or U152 (N_152,In_550,In_219);
nor U153 (N_153,In_491,In_373);
nor U154 (N_154,In_728,In_602);
nor U155 (N_155,In_228,In_259);
or U156 (N_156,In_237,In_507);
nor U157 (N_157,In_286,In_269);
xor U158 (N_158,In_675,In_325);
nand U159 (N_159,In_256,In_447);
nand U160 (N_160,In_278,In_404);
or U161 (N_161,In_700,In_380);
nor U162 (N_162,In_569,In_423);
or U163 (N_163,In_117,In_266);
or U164 (N_164,In_207,In_258);
xnor U165 (N_165,In_128,In_676);
or U166 (N_166,In_721,In_600);
xnor U167 (N_167,In_419,In_118);
xnor U168 (N_168,In_190,In_392);
xnor U169 (N_169,In_287,In_628);
and U170 (N_170,In_307,In_367);
xnor U171 (N_171,In_476,In_744);
xnor U172 (N_172,In_302,In_211);
nor U173 (N_173,In_482,In_291);
xor U174 (N_174,In_573,In_227);
nand U175 (N_175,In_662,In_103);
nor U176 (N_176,In_609,In_716);
nor U177 (N_177,In_197,In_693);
xnor U178 (N_178,In_712,In_119);
and U179 (N_179,In_597,In_13);
and U180 (N_180,In_534,In_232);
or U181 (N_181,In_730,In_240);
nor U182 (N_182,In_339,In_520);
nand U183 (N_183,In_315,In_657);
and U184 (N_184,In_540,In_627);
xor U185 (N_185,In_641,In_341);
nand U186 (N_186,In_136,In_738);
nor U187 (N_187,In_681,In_452);
or U188 (N_188,In_326,In_495);
nand U189 (N_189,In_59,In_698);
xnor U190 (N_190,In_0,In_330);
nand U191 (N_191,In_620,In_249);
nor U192 (N_192,In_54,In_165);
nand U193 (N_193,In_74,In_559);
or U194 (N_194,In_274,In_673);
xnor U195 (N_195,In_106,In_710);
xor U196 (N_196,In_458,In_651);
or U197 (N_197,In_93,In_141);
nor U198 (N_198,In_124,In_68);
nor U199 (N_199,In_192,In_552);
nand U200 (N_200,In_483,In_234);
nor U201 (N_201,In_184,N_5);
and U202 (N_202,In_387,In_388);
and U203 (N_203,In_711,In_490);
nand U204 (N_204,In_161,In_579);
and U205 (N_205,In_725,In_603);
or U206 (N_206,N_101,N_3);
nand U207 (N_207,In_79,In_149);
xnor U208 (N_208,In_741,In_671);
xnor U209 (N_209,In_221,In_220);
nor U210 (N_210,N_64,N_116);
xnor U211 (N_211,In_181,N_148);
and U212 (N_212,In_548,N_40);
and U213 (N_213,In_260,In_120);
nor U214 (N_214,In_299,In_210);
and U215 (N_215,In_562,In_637);
and U216 (N_216,In_558,In_154);
nand U217 (N_217,In_312,N_80);
or U218 (N_218,In_113,In_317);
and U219 (N_219,In_618,N_48);
and U220 (N_220,N_182,N_98);
and U221 (N_221,N_84,In_409);
nor U222 (N_222,In_58,N_179);
xnor U223 (N_223,In_104,N_35);
nand U224 (N_224,In_436,N_88);
xnor U225 (N_225,N_121,In_88);
and U226 (N_226,In_248,N_106);
and U227 (N_227,In_167,N_128);
and U228 (N_228,In_553,N_85);
nand U229 (N_229,N_107,N_177);
nor U230 (N_230,In_233,In_542);
nor U231 (N_231,In_736,In_703);
and U232 (N_232,In_352,N_67);
or U233 (N_233,N_171,N_140);
and U234 (N_234,N_139,In_242);
nor U235 (N_235,In_308,N_104);
xnor U236 (N_236,In_243,In_138);
xor U237 (N_237,N_147,In_345);
nand U238 (N_238,N_6,N_100);
nand U239 (N_239,In_497,In_313);
and U240 (N_240,In_179,In_257);
xnor U241 (N_241,N_86,In_660);
or U242 (N_242,N_0,In_509);
or U243 (N_243,In_531,In_372);
and U244 (N_244,In_523,In_344);
xnor U245 (N_245,N_163,N_27);
or U246 (N_246,N_161,N_24);
or U247 (N_247,N_180,In_632);
nor U248 (N_248,N_105,N_2);
nor U249 (N_249,In_166,In_267);
nand U250 (N_250,In_426,N_168);
or U251 (N_251,In_605,In_183);
and U252 (N_252,In_400,In_123);
or U253 (N_253,In_455,N_47);
nand U254 (N_254,N_150,In_17);
and U255 (N_255,In_9,In_62);
or U256 (N_256,In_718,N_93);
xnor U257 (N_257,In_393,In_140);
and U258 (N_258,N_77,N_70);
or U259 (N_259,In_467,In_172);
and U260 (N_260,N_169,N_162);
or U261 (N_261,In_182,In_735);
nor U262 (N_262,N_141,N_9);
nand U263 (N_263,In_363,N_71);
nor U264 (N_264,N_191,In_453);
xor U265 (N_265,In_678,In_347);
nor U266 (N_266,N_26,N_53);
and U267 (N_267,N_103,In_472);
and U268 (N_268,N_165,In_379);
nor U269 (N_269,N_54,N_49);
nand U270 (N_270,In_658,In_85);
nand U271 (N_271,In_262,In_668);
and U272 (N_272,In_526,In_425);
and U273 (N_273,In_656,In_395);
nor U274 (N_274,In_145,In_398);
nand U275 (N_275,N_113,N_74);
nand U276 (N_276,In_512,In_80);
and U277 (N_277,In_568,N_115);
nor U278 (N_278,In_144,In_296);
xnor U279 (N_279,In_105,N_72);
and U280 (N_280,N_132,In_555);
nand U281 (N_281,In_292,In_574);
nor U282 (N_282,N_19,N_31);
and U283 (N_283,In_5,In_502);
nor U284 (N_284,N_151,N_38);
xor U285 (N_285,N_138,In_160);
xnor U286 (N_286,In_692,In_503);
nand U287 (N_287,In_413,N_90);
nand U288 (N_288,N_96,In_135);
xnor U289 (N_289,In_501,In_639);
or U290 (N_290,In_417,In_517);
nor U291 (N_291,In_465,In_593);
nand U292 (N_292,N_58,In_505);
nor U293 (N_293,N_110,In_429);
or U294 (N_294,N_146,N_89);
and U295 (N_295,N_155,In_96);
xor U296 (N_296,In_477,N_153);
nor U297 (N_297,N_25,N_59);
and U298 (N_298,In_204,In_577);
nor U299 (N_299,N_73,In_545);
nor U300 (N_300,N_112,N_44);
nand U301 (N_301,In_412,In_580);
or U302 (N_302,In_516,In_733);
and U303 (N_303,In_1,In_567);
or U304 (N_304,In_745,In_209);
or U305 (N_305,N_158,In_606);
nand U306 (N_306,In_329,In_26);
xor U307 (N_307,N_83,N_76);
and U308 (N_308,In_318,In_727);
or U309 (N_309,N_120,N_152);
nor U310 (N_310,N_56,N_29);
nor U311 (N_311,N_57,In_298);
and U312 (N_312,In_275,In_230);
xor U313 (N_313,In_462,In_66);
nor U314 (N_314,In_410,N_144);
and U315 (N_315,N_20,In_195);
nor U316 (N_316,In_238,In_188);
or U317 (N_317,In_132,N_92);
nand U318 (N_318,In_355,N_4);
and U319 (N_319,In_44,In_213);
nor U320 (N_320,In_688,In_522);
xor U321 (N_321,N_17,In_659);
or U322 (N_322,In_82,In_631);
and U323 (N_323,In_201,In_475);
and U324 (N_324,N_8,In_661);
nand U325 (N_325,In_646,In_61);
nor U326 (N_326,N_126,N_193);
and U327 (N_327,In_634,In_726);
nand U328 (N_328,In_566,In_178);
nor U329 (N_329,N_41,N_15);
nand U330 (N_330,In_176,In_724);
nand U331 (N_331,In_596,In_350);
or U332 (N_332,N_130,In_557);
nand U333 (N_333,In_529,N_87);
and U334 (N_334,In_739,N_187);
nor U335 (N_335,N_133,In_493);
and U336 (N_336,In_747,In_370);
xnor U337 (N_337,N_62,In_645);
nor U338 (N_338,In_643,In_384);
nand U339 (N_339,In_612,In_459);
nand U340 (N_340,In_229,In_510);
xnor U341 (N_341,In_638,In_2);
nand U342 (N_342,In_39,In_616);
and U343 (N_343,In_705,In_130);
xor U344 (N_344,In_186,In_702);
nor U345 (N_345,In_282,In_411);
nand U346 (N_346,In_115,In_239);
xnor U347 (N_347,In_212,In_443);
xor U348 (N_348,In_440,N_197);
and U349 (N_349,In_556,N_45);
nand U350 (N_350,N_28,N_176);
nor U351 (N_351,In_67,In_543);
nand U352 (N_352,In_336,In_304);
nor U353 (N_353,In_98,N_117);
nand U354 (N_354,N_23,In_290);
xor U355 (N_355,N_184,In_391);
xor U356 (N_356,In_346,In_108);
xnor U357 (N_357,N_192,In_402);
nor U358 (N_358,In_595,In_94);
and U359 (N_359,In_43,N_109);
xnor U360 (N_360,In_382,In_69);
nor U361 (N_361,N_118,In_268);
nor U362 (N_362,In_538,N_145);
and U363 (N_363,In_334,N_61);
xor U364 (N_364,N_170,In_208);
xor U365 (N_365,N_82,N_18);
nand U366 (N_366,In_385,In_10);
nor U367 (N_367,N_167,N_175);
nor U368 (N_368,N_1,In_448);
nand U369 (N_369,In_139,In_498);
nand U370 (N_370,In_672,In_403);
xnor U371 (N_371,N_55,In_473);
xnor U372 (N_372,N_143,N_78);
and U373 (N_373,In_406,N_99);
or U374 (N_374,In_45,N_119);
nand U375 (N_375,In_323,In_663);
nor U376 (N_376,In_582,N_186);
or U377 (N_377,N_189,In_247);
or U378 (N_378,In_734,N_42);
or U379 (N_379,In_561,N_166);
xnor U380 (N_380,In_666,In_513);
xor U381 (N_381,In_24,N_21);
and U382 (N_382,In_444,In_629);
nand U383 (N_383,In_480,In_652);
nor U384 (N_384,In_360,N_81);
and U385 (N_385,In_707,In_187);
or U386 (N_386,In_713,In_431);
xnor U387 (N_387,N_154,In_169);
or U388 (N_388,N_94,In_494);
or U389 (N_389,In_530,N_134);
xnor U390 (N_390,In_469,In_15);
or U391 (N_391,In_481,In_129);
or U392 (N_392,In_376,N_7);
nand U393 (N_393,N_185,In_468);
and U394 (N_394,N_32,In_434);
or U395 (N_395,N_135,In_636);
xor U396 (N_396,In_309,N_14);
and U397 (N_397,In_396,N_68);
and U398 (N_398,N_172,In_654);
and U399 (N_399,In_322,N_127);
xor U400 (N_400,In_202,N_164);
or U401 (N_401,In_122,N_181);
nand U402 (N_402,In_524,N_340);
nand U403 (N_403,N_223,N_380);
nor U404 (N_404,In_701,N_95);
and U405 (N_405,In_333,N_367);
and U406 (N_406,N_294,In_246);
and U407 (N_407,N_325,N_304);
nor U408 (N_408,N_312,N_249);
and U409 (N_409,In_625,In_563);
and U410 (N_410,N_216,N_260);
or U411 (N_411,In_433,In_263);
nand U412 (N_412,N_111,In_508);
and U413 (N_413,In_685,N_270);
and U414 (N_414,In_244,N_214);
nand U415 (N_415,N_224,N_244);
or U416 (N_416,N_358,N_157);
xnor U417 (N_417,N_242,N_239);
nand U418 (N_418,N_395,N_365);
nand U419 (N_419,In_610,In_565);
nand U420 (N_420,In_11,In_679);
xor U421 (N_421,In_53,In_137);
nand U422 (N_422,In_706,In_156);
nor U423 (N_423,N_259,N_11);
nand U424 (N_424,N_210,N_306);
nand U425 (N_425,N_322,N_379);
and U426 (N_426,N_376,N_334);
or U427 (N_427,N_240,N_227);
nand U428 (N_428,N_383,N_201);
or U429 (N_429,N_203,N_256);
and U430 (N_430,N_308,N_12);
and U431 (N_431,In_551,N_381);
and U432 (N_432,N_370,N_362);
nor U433 (N_433,N_198,N_225);
or U434 (N_434,N_344,N_310);
and U435 (N_435,N_237,N_302);
xnor U436 (N_436,N_389,N_220);
nor U437 (N_437,N_373,N_43);
or U438 (N_438,N_290,In_250);
xnor U439 (N_439,N_289,In_153);
and U440 (N_440,N_114,N_337);
nand U441 (N_441,N_34,In_70);
and U442 (N_442,In_6,N_399);
and U443 (N_443,N_60,N_397);
and U444 (N_444,N_282,In_617);
xor U445 (N_445,N_196,In_368);
nor U446 (N_446,N_160,N_298);
or U447 (N_447,N_124,N_262);
nand U448 (N_448,N_343,In_157);
nor U449 (N_449,N_222,In_127);
and U450 (N_450,N_13,N_374);
or U451 (N_451,N_263,N_392);
nand U452 (N_452,N_190,N_274);
and U453 (N_453,N_388,N_385);
and U454 (N_454,N_320,N_221);
nor U455 (N_455,N_291,In_143);
xnor U456 (N_456,N_37,In_525);
nand U457 (N_457,In_691,N_253);
and U458 (N_458,N_22,N_356);
and U459 (N_459,In_150,N_39);
nor U460 (N_460,N_295,N_313);
and U461 (N_461,N_238,N_178);
nand U462 (N_462,N_361,N_50);
nand U463 (N_463,N_318,In_4);
nand U464 (N_464,N_398,In_48);
nor U465 (N_465,N_267,N_333);
and U466 (N_466,N_183,N_394);
and U467 (N_467,N_314,N_357);
nand U468 (N_468,N_366,In_424);
nand U469 (N_469,N_287,N_297);
xnor U470 (N_470,In_364,N_354);
nor U471 (N_471,N_137,N_209);
xor U472 (N_472,In_575,N_315);
nor U473 (N_473,N_350,N_331);
or U474 (N_474,In_174,N_338);
or U475 (N_475,In_539,In_442);
xor U476 (N_476,N_378,N_255);
nor U477 (N_477,N_387,N_236);
and U478 (N_478,N_79,N_275);
xor U479 (N_479,In_492,N_396);
nand U480 (N_480,N_369,In_271);
nor U481 (N_481,In_369,N_125);
or U482 (N_482,N_226,N_328);
and U483 (N_483,In_251,N_352);
and U484 (N_484,In_76,N_131);
or U485 (N_485,N_329,N_332);
and U486 (N_486,In_590,In_722);
xor U487 (N_487,N_51,N_91);
or U488 (N_488,In_191,In_407);
or U489 (N_489,N_258,N_280);
nand U490 (N_490,N_254,In_611);
or U491 (N_491,In_12,N_363);
or U492 (N_492,N_123,N_271);
nor U493 (N_493,N_300,N_159);
and U494 (N_494,In_432,N_129);
nand U495 (N_495,In_265,N_377);
nor U496 (N_496,N_391,N_212);
xnor U497 (N_497,N_384,In_311);
and U498 (N_498,In_454,In_42);
nor U499 (N_499,N_327,N_273);
nand U500 (N_500,In_421,N_195);
xor U501 (N_501,N_215,In_134);
nand U502 (N_502,N_359,N_336);
xor U503 (N_503,In_546,N_233);
nand U504 (N_504,In_399,N_299);
xor U505 (N_505,N_231,In_95);
nand U506 (N_506,N_269,N_63);
xnor U507 (N_507,N_202,N_342);
and U508 (N_508,In_84,N_355);
or U509 (N_509,N_247,N_174);
nor U510 (N_510,N_208,N_206);
or U511 (N_511,N_228,N_217);
or U512 (N_512,N_309,N_321);
nand U513 (N_513,N_142,N_235);
or U514 (N_514,N_351,N_173);
or U515 (N_515,N_218,N_265);
xnor U516 (N_516,N_303,N_52);
xor U517 (N_517,N_317,In_348);
nand U518 (N_518,N_279,N_229);
and U519 (N_519,In_377,N_136);
nand U520 (N_520,N_188,N_272);
xor U521 (N_521,In_18,N_250);
nand U522 (N_522,N_278,N_33);
xnor U523 (N_523,N_30,In_110);
nand U524 (N_524,N_293,In_732);
xnor U525 (N_525,N_10,In_295);
nand U526 (N_526,N_345,N_277);
and U527 (N_527,N_211,N_346);
nand U528 (N_528,In_519,In_22);
nor U529 (N_529,N_292,N_296);
and U530 (N_530,N_353,N_268);
nand U531 (N_531,N_371,N_97);
nand U532 (N_532,In_321,N_122);
xnor U533 (N_533,N_281,N_248);
nor U534 (N_534,N_316,N_319);
nand U535 (N_535,In_349,N_16);
nand U536 (N_536,N_199,N_301);
xnor U537 (N_537,N_349,In_305);
nand U538 (N_538,In_328,N_285);
nand U539 (N_539,In_689,N_207);
nand U540 (N_540,N_108,In_159);
nand U541 (N_541,N_348,N_276);
and U542 (N_542,N_326,N_156);
nor U543 (N_543,In_206,N_284);
nand U544 (N_544,N_149,In_77);
nand U545 (N_545,N_36,N_386);
and U546 (N_546,N_264,N_382);
nand U547 (N_547,N_102,N_243);
xnor U548 (N_548,N_194,N_46);
or U549 (N_549,N_66,N_252);
nor U550 (N_550,In_670,N_245);
and U551 (N_551,N_261,N_234);
nor U552 (N_552,N_375,N_372);
xor U553 (N_553,In_626,N_368);
nand U554 (N_554,N_204,N_347);
xnor U555 (N_555,N_230,N_330);
or U556 (N_556,N_339,N_390);
xnor U557 (N_557,N_360,N_65);
nor U558 (N_558,N_283,N_205);
xnor U559 (N_559,N_286,In_21);
nor U560 (N_560,N_257,In_420);
xnor U561 (N_561,N_323,N_266);
or U562 (N_562,In_8,N_232);
nand U563 (N_563,N_393,N_219);
nor U564 (N_564,N_75,In_310);
nor U565 (N_565,In_451,N_364);
and U566 (N_566,N_324,N_288);
xnor U567 (N_567,N_305,N_251);
and U568 (N_568,N_246,N_341);
nand U569 (N_569,In_163,N_200);
or U570 (N_570,N_69,N_213);
nand U571 (N_571,N_335,In_532);
and U572 (N_572,N_241,N_307);
nand U573 (N_573,N_311,In_416);
nand U574 (N_574,In_441,In_731);
nor U575 (N_575,In_263,In_21);
nand U576 (N_576,N_277,N_260);
nor U577 (N_577,N_317,In_143);
and U578 (N_578,N_328,N_373);
or U579 (N_579,N_159,N_12);
or U580 (N_580,N_214,N_205);
xor U581 (N_581,N_372,N_124);
nor U582 (N_582,In_706,N_259);
or U583 (N_583,N_297,N_258);
and U584 (N_584,N_395,N_224);
nor U585 (N_585,In_22,N_328);
or U586 (N_586,N_36,N_380);
and U587 (N_587,N_66,N_296);
xnor U588 (N_588,In_368,N_319);
nor U589 (N_589,In_691,N_234);
and U590 (N_590,N_202,N_97);
xnor U591 (N_591,N_267,In_143);
and U592 (N_592,In_575,N_300);
xnor U593 (N_593,N_263,N_240);
xor U594 (N_594,N_256,In_625);
or U595 (N_595,N_231,N_255);
or U596 (N_596,In_348,In_420);
or U597 (N_597,N_369,In_416);
nand U598 (N_598,N_288,In_271);
nor U599 (N_599,In_95,In_6);
xnor U600 (N_600,N_415,N_407);
or U601 (N_601,N_406,N_501);
nor U602 (N_602,N_551,N_549);
or U603 (N_603,N_510,N_491);
nand U604 (N_604,N_598,N_535);
or U605 (N_605,N_433,N_420);
and U606 (N_606,N_405,N_539);
or U607 (N_607,N_479,N_476);
or U608 (N_608,N_596,N_515);
and U609 (N_609,N_497,N_526);
nand U610 (N_610,N_496,N_409);
or U611 (N_611,N_457,N_524);
nor U612 (N_612,N_593,N_584);
nand U613 (N_613,N_430,N_558);
xor U614 (N_614,N_452,N_520);
xnor U615 (N_615,N_440,N_489);
and U616 (N_616,N_421,N_464);
nor U617 (N_617,N_404,N_599);
nor U618 (N_618,N_571,N_547);
nor U619 (N_619,N_482,N_521);
and U620 (N_620,N_578,N_597);
and U621 (N_621,N_522,N_590);
xor U622 (N_622,N_460,N_592);
nand U623 (N_623,N_562,N_577);
xor U624 (N_624,N_569,N_447);
or U625 (N_625,N_438,N_534);
nand U626 (N_626,N_556,N_595);
nand U627 (N_627,N_424,N_472);
nor U628 (N_628,N_448,N_498);
and U629 (N_629,N_572,N_400);
or U630 (N_630,N_532,N_449);
xor U631 (N_631,N_467,N_579);
xnor U632 (N_632,N_517,N_588);
and U633 (N_633,N_507,N_540);
and U634 (N_634,N_566,N_475);
nor U635 (N_635,N_499,N_477);
nor U636 (N_636,N_525,N_570);
xor U637 (N_637,N_533,N_453);
and U638 (N_638,N_466,N_431);
or U639 (N_639,N_473,N_506);
xor U640 (N_640,N_469,N_586);
nor U641 (N_641,N_436,N_410);
xor U642 (N_642,N_443,N_468);
or U643 (N_643,N_495,N_518);
and U644 (N_644,N_531,N_455);
nand U645 (N_645,N_542,N_417);
and U646 (N_646,N_563,N_444);
nand U647 (N_647,N_543,N_458);
and U648 (N_648,N_544,N_509);
or U649 (N_649,N_575,N_555);
or U650 (N_650,N_594,N_454);
and U651 (N_651,N_459,N_441);
or U652 (N_652,N_439,N_402);
or U653 (N_653,N_564,N_486);
nand U654 (N_654,N_508,N_529);
nor U655 (N_655,N_528,N_483);
or U656 (N_656,N_451,N_591);
xor U657 (N_657,N_541,N_545);
nor U658 (N_658,N_492,N_435);
or U659 (N_659,N_548,N_559);
and U660 (N_660,N_413,N_502);
xnor U661 (N_661,N_546,N_401);
xnor U662 (N_662,N_581,N_462);
nor U663 (N_663,N_493,N_583);
nand U664 (N_664,N_511,N_527);
or U665 (N_665,N_536,N_429);
nor U666 (N_666,N_552,N_480);
xor U667 (N_667,N_519,N_434);
nand U668 (N_668,N_446,N_470);
and U669 (N_669,N_425,N_585);
xor U670 (N_670,N_478,N_456);
xnor U671 (N_671,N_487,N_554);
xor U672 (N_672,N_411,N_550);
nand U673 (N_673,N_505,N_538);
nor U674 (N_674,N_450,N_574);
nor U675 (N_675,N_481,N_408);
and U676 (N_676,N_553,N_490);
nand U677 (N_677,N_427,N_514);
or U678 (N_678,N_426,N_576);
and U679 (N_679,N_414,N_442);
xor U680 (N_680,N_463,N_416);
xnor U681 (N_681,N_560,N_589);
or U682 (N_682,N_465,N_488);
nor U683 (N_683,N_471,N_484);
or U684 (N_684,N_418,N_537);
and U685 (N_685,N_428,N_503);
nor U686 (N_686,N_422,N_485);
or U687 (N_687,N_504,N_587);
and U688 (N_688,N_423,N_432);
xor U689 (N_689,N_474,N_582);
nand U690 (N_690,N_419,N_403);
or U691 (N_691,N_512,N_494);
or U692 (N_692,N_437,N_513);
and U693 (N_693,N_565,N_412);
nand U694 (N_694,N_557,N_561);
nand U695 (N_695,N_530,N_567);
nor U696 (N_696,N_516,N_568);
or U697 (N_697,N_580,N_500);
nand U698 (N_698,N_573,N_461);
or U699 (N_699,N_445,N_523);
xnor U700 (N_700,N_585,N_565);
and U701 (N_701,N_591,N_491);
nor U702 (N_702,N_430,N_427);
and U703 (N_703,N_554,N_467);
nand U704 (N_704,N_454,N_488);
or U705 (N_705,N_543,N_472);
and U706 (N_706,N_411,N_438);
or U707 (N_707,N_523,N_453);
or U708 (N_708,N_563,N_595);
nor U709 (N_709,N_448,N_506);
and U710 (N_710,N_431,N_588);
nor U711 (N_711,N_505,N_543);
nand U712 (N_712,N_430,N_544);
nand U713 (N_713,N_542,N_575);
nor U714 (N_714,N_448,N_518);
nand U715 (N_715,N_582,N_440);
nor U716 (N_716,N_569,N_485);
or U717 (N_717,N_540,N_407);
and U718 (N_718,N_456,N_476);
or U719 (N_719,N_557,N_565);
nor U720 (N_720,N_527,N_487);
nand U721 (N_721,N_477,N_502);
nor U722 (N_722,N_511,N_477);
and U723 (N_723,N_442,N_435);
nor U724 (N_724,N_530,N_541);
or U725 (N_725,N_483,N_492);
or U726 (N_726,N_458,N_588);
xor U727 (N_727,N_476,N_580);
and U728 (N_728,N_577,N_434);
and U729 (N_729,N_409,N_445);
nor U730 (N_730,N_522,N_580);
and U731 (N_731,N_517,N_544);
nand U732 (N_732,N_577,N_424);
and U733 (N_733,N_597,N_598);
and U734 (N_734,N_501,N_560);
nand U735 (N_735,N_580,N_541);
and U736 (N_736,N_530,N_473);
and U737 (N_737,N_432,N_549);
or U738 (N_738,N_419,N_489);
and U739 (N_739,N_535,N_446);
and U740 (N_740,N_406,N_496);
and U741 (N_741,N_522,N_584);
nor U742 (N_742,N_495,N_410);
or U743 (N_743,N_515,N_459);
nand U744 (N_744,N_516,N_416);
nand U745 (N_745,N_548,N_525);
nor U746 (N_746,N_417,N_434);
xnor U747 (N_747,N_469,N_555);
nor U748 (N_748,N_508,N_582);
nor U749 (N_749,N_573,N_556);
nor U750 (N_750,N_554,N_413);
nor U751 (N_751,N_525,N_544);
nand U752 (N_752,N_461,N_422);
xnor U753 (N_753,N_495,N_451);
nand U754 (N_754,N_520,N_485);
nand U755 (N_755,N_482,N_483);
and U756 (N_756,N_577,N_595);
nor U757 (N_757,N_427,N_416);
or U758 (N_758,N_567,N_584);
nand U759 (N_759,N_575,N_468);
and U760 (N_760,N_458,N_462);
nand U761 (N_761,N_518,N_454);
nand U762 (N_762,N_590,N_405);
xnor U763 (N_763,N_575,N_432);
xnor U764 (N_764,N_412,N_460);
and U765 (N_765,N_570,N_420);
nor U766 (N_766,N_486,N_594);
and U767 (N_767,N_452,N_563);
and U768 (N_768,N_452,N_522);
or U769 (N_769,N_586,N_575);
nand U770 (N_770,N_569,N_521);
nand U771 (N_771,N_427,N_570);
nor U772 (N_772,N_578,N_467);
nor U773 (N_773,N_434,N_472);
nor U774 (N_774,N_538,N_580);
nor U775 (N_775,N_525,N_504);
nand U776 (N_776,N_563,N_593);
and U777 (N_777,N_578,N_542);
or U778 (N_778,N_521,N_494);
nor U779 (N_779,N_452,N_497);
nand U780 (N_780,N_400,N_482);
nor U781 (N_781,N_437,N_577);
nand U782 (N_782,N_427,N_522);
and U783 (N_783,N_581,N_505);
nor U784 (N_784,N_423,N_487);
nor U785 (N_785,N_590,N_421);
or U786 (N_786,N_528,N_527);
xnor U787 (N_787,N_458,N_492);
nand U788 (N_788,N_558,N_530);
xnor U789 (N_789,N_404,N_513);
xor U790 (N_790,N_402,N_431);
nand U791 (N_791,N_423,N_534);
or U792 (N_792,N_413,N_573);
xor U793 (N_793,N_541,N_488);
xnor U794 (N_794,N_454,N_464);
or U795 (N_795,N_526,N_433);
or U796 (N_796,N_406,N_482);
xnor U797 (N_797,N_539,N_517);
or U798 (N_798,N_566,N_511);
xnor U799 (N_799,N_529,N_408);
nor U800 (N_800,N_720,N_791);
nand U801 (N_801,N_681,N_654);
or U802 (N_802,N_788,N_607);
nor U803 (N_803,N_748,N_715);
or U804 (N_804,N_662,N_758);
xor U805 (N_805,N_650,N_760);
nand U806 (N_806,N_642,N_765);
nor U807 (N_807,N_759,N_622);
nand U808 (N_808,N_731,N_764);
nor U809 (N_809,N_610,N_721);
nand U810 (N_810,N_713,N_766);
and U811 (N_811,N_677,N_750);
and U812 (N_812,N_796,N_768);
or U813 (N_813,N_769,N_795);
or U814 (N_814,N_704,N_763);
xnor U815 (N_815,N_726,N_648);
xnor U816 (N_816,N_635,N_645);
nand U817 (N_817,N_618,N_767);
xor U818 (N_818,N_786,N_694);
and U819 (N_819,N_798,N_782);
and U820 (N_820,N_779,N_699);
xor U821 (N_821,N_789,N_696);
and U822 (N_822,N_676,N_669);
and U823 (N_823,N_776,N_611);
xnor U824 (N_824,N_605,N_714);
or U825 (N_825,N_702,N_683);
nor U826 (N_826,N_665,N_743);
nor U827 (N_827,N_753,N_738);
or U828 (N_828,N_604,N_633);
nor U829 (N_829,N_701,N_752);
and U830 (N_830,N_628,N_690);
nand U831 (N_831,N_736,N_719);
nand U832 (N_832,N_793,N_762);
or U833 (N_833,N_686,N_615);
nand U834 (N_834,N_614,N_603);
nand U835 (N_835,N_717,N_777);
or U836 (N_836,N_712,N_613);
and U837 (N_837,N_641,N_755);
nand U838 (N_838,N_653,N_689);
xor U839 (N_839,N_672,N_756);
or U840 (N_840,N_697,N_783);
and U841 (N_841,N_659,N_706);
and U842 (N_842,N_740,N_725);
nor U843 (N_843,N_797,N_707);
and U844 (N_844,N_606,N_733);
or U845 (N_845,N_727,N_638);
xnor U846 (N_846,N_774,N_711);
or U847 (N_847,N_761,N_716);
or U848 (N_848,N_637,N_739);
nand U849 (N_849,N_671,N_680);
or U850 (N_850,N_749,N_631);
nor U851 (N_851,N_770,N_724);
xnor U852 (N_852,N_656,N_600);
nand U853 (N_853,N_670,N_623);
or U854 (N_854,N_709,N_602);
xor U855 (N_855,N_688,N_754);
nand U856 (N_856,N_691,N_772);
nand U857 (N_857,N_734,N_679);
nand U858 (N_858,N_632,N_609);
and U859 (N_859,N_673,N_705);
nor U860 (N_860,N_682,N_608);
and U861 (N_861,N_601,N_771);
nand U862 (N_862,N_723,N_678);
xnor U863 (N_863,N_745,N_652);
and U864 (N_864,N_693,N_781);
nand U865 (N_865,N_646,N_773);
and U866 (N_866,N_746,N_667);
nor U867 (N_867,N_708,N_790);
and U868 (N_868,N_630,N_674);
and U869 (N_869,N_751,N_664);
nor U870 (N_870,N_675,N_744);
nor U871 (N_871,N_735,N_666);
nor U872 (N_872,N_732,N_658);
and U873 (N_873,N_616,N_794);
nor U874 (N_874,N_692,N_722);
nor U875 (N_875,N_780,N_757);
xnor U876 (N_876,N_624,N_728);
or U877 (N_877,N_643,N_737);
and U878 (N_878,N_778,N_660);
nor U879 (N_879,N_612,N_647);
nor U880 (N_880,N_661,N_620);
xnor U881 (N_881,N_639,N_747);
or U882 (N_882,N_718,N_655);
xnor U883 (N_883,N_687,N_629);
xor U884 (N_884,N_730,N_619);
or U885 (N_885,N_785,N_617);
xor U886 (N_886,N_742,N_700);
nor U887 (N_887,N_657,N_644);
nor U888 (N_888,N_626,N_710);
xor U889 (N_889,N_663,N_792);
or U890 (N_890,N_729,N_695);
and U891 (N_891,N_698,N_636);
and U892 (N_892,N_668,N_627);
xor U893 (N_893,N_775,N_799);
xor U894 (N_894,N_640,N_787);
nand U895 (N_895,N_685,N_649);
nand U896 (N_896,N_651,N_634);
xnor U897 (N_897,N_684,N_741);
nand U898 (N_898,N_703,N_625);
or U899 (N_899,N_621,N_784);
nor U900 (N_900,N_761,N_780);
xor U901 (N_901,N_663,N_741);
nor U902 (N_902,N_626,N_603);
and U903 (N_903,N_626,N_794);
xnor U904 (N_904,N_769,N_665);
and U905 (N_905,N_654,N_669);
or U906 (N_906,N_693,N_664);
nor U907 (N_907,N_760,N_644);
xor U908 (N_908,N_785,N_708);
and U909 (N_909,N_668,N_736);
xnor U910 (N_910,N_663,N_782);
xor U911 (N_911,N_632,N_725);
nand U912 (N_912,N_609,N_660);
and U913 (N_913,N_661,N_663);
xor U914 (N_914,N_624,N_672);
nand U915 (N_915,N_606,N_605);
xnor U916 (N_916,N_631,N_766);
or U917 (N_917,N_746,N_745);
and U918 (N_918,N_771,N_622);
xor U919 (N_919,N_714,N_744);
nor U920 (N_920,N_715,N_660);
xnor U921 (N_921,N_706,N_605);
and U922 (N_922,N_699,N_709);
or U923 (N_923,N_680,N_610);
nor U924 (N_924,N_610,N_702);
nand U925 (N_925,N_659,N_686);
nand U926 (N_926,N_697,N_799);
and U927 (N_927,N_744,N_793);
and U928 (N_928,N_664,N_672);
nand U929 (N_929,N_785,N_767);
and U930 (N_930,N_729,N_687);
nand U931 (N_931,N_747,N_742);
and U932 (N_932,N_713,N_748);
nand U933 (N_933,N_685,N_693);
nand U934 (N_934,N_668,N_741);
nor U935 (N_935,N_635,N_618);
nor U936 (N_936,N_662,N_672);
xor U937 (N_937,N_657,N_775);
xor U938 (N_938,N_626,N_668);
nand U939 (N_939,N_622,N_694);
nor U940 (N_940,N_627,N_793);
xor U941 (N_941,N_643,N_675);
and U942 (N_942,N_736,N_608);
nand U943 (N_943,N_695,N_640);
or U944 (N_944,N_709,N_796);
and U945 (N_945,N_674,N_776);
nand U946 (N_946,N_629,N_712);
or U947 (N_947,N_707,N_658);
and U948 (N_948,N_730,N_637);
xor U949 (N_949,N_642,N_793);
or U950 (N_950,N_607,N_752);
or U951 (N_951,N_772,N_762);
nor U952 (N_952,N_690,N_605);
nor U953 (N_953,N_724,N_692);
nor U954 (N_954,N_775,N_742);
or U955 (N_955,N_669,N_777);
nand U956 (N_956,N_751,N_743);
nor U957 (N_957,N_741,N_752);
xnor U958 (N_958,N_765,N_717);
xor U959 (N_959,N_795,N_717);
or U960 (N_960,N_768,N_757);
and U961 (N_961,N_798,N_638);
and U962 (N_962,N_759,N_704);
and U963 (N_963,N_702,N_796);
xor U964 (N_964,N_655,N_674);
and U965 (N_965,N_700,N_677);
xnor U966 (N_966,N_659,N_673);
or U967 (N_967,N_780,N_655);
nand U968 (N_968,N_754,N_791);
and U969 (N_969,N_662,N_644);
and U970 (N_970,N_762,N_605);
nand U971 (N_971,N_773,N_659);
or U972 (N_972,N_709,N_630);
nor U973 (N_973,N_772,N_734);
nor U974 (N_974,N_646,N_605);
and U975 (N_975,N_611,N_726);
and U976 (N_976,N_764,N_650);
nand U977 (N_977,N_600,N_658);
nor U978 (N_978,N_777,N_753);
xor U979 (N_979,N_745,N_658);
nand U980 (N_980,N_755,N_713);
nand U981 (N_981,N_703,N_612);
nor U982 (N_982,N_703,N_658);
nand U983 (N_983,N_766,N_625);
nor U984 (N_984,N_746,N_610);
or U985 (N_985,N_707,N_725);
nand U986 (N_986,N_649,N_784);
nand U987 (N_987,N_795,N_651);
or U988 (N_988,N_644,N_688);
or U989 (N_989,N_733,N_680);
xor U990 (N_990,N_669,N_764);
xnor U991 (N_991,N_714,N_632);
xnor U992 (N_992,N_787,N_710);
xnor U993 (N_993,N_784,N_706);
or U994 (N_994,N_683,N_708);
and U995 (N_995,N_610,N_614);
xnor U996 (N_996,N_746,N_682);
xnor U997 (N_997,N_745,N_648);
nand U998 (N_998,N_607,N_600);
nor U999 (N_999,N_745,N_637);
or U1000 (N_1000,N_896,N_920);
nand U1001 (N_1001,N_952,N_889);
nor U1002 (N_1002,N_921,N_816);
xnor U1003 (N_1003,N_843,N_954);
nand U1004 (N_1004,N_809,N_811);
nor U1005 (N_1005,N_994,N_940);
nor U1006 (N_1006,N_914,N_841);
or U1007 (N_1007,N_910,N_849);
nand U1008 (N_1008,N_856,N_851);
xnor U1009 (N_1009,N_912,N_974);
or U1010 (N_1010,N_805,N_862);
nor U1011 (N_1011,N_853,N_875);
and U1012 (N_1012,N_986,N_842);
nand U1013 (N_1013,N_987,N_931);
xnor U1014 (N_1014,N_878,N_959);
xnor U1015 (N_1015,N_953,N_876);
nor U1016 (N_1016,N_937,N_887);
and U1017 (N_1017,N_904,N_833);
nand U1018 (N_1018,N_846,N_903);
and U1019 (N_1019,N_916,N_897);
xnor U1020 (N_1020,N_882,N_957);
and U1021 (N_1021,N_939,N_832);
or U1022 (N_1022,N_871,N_941);
nand U1023 (N_1023,N_980,N_858);
nor U1024 (N_1024,N_866,N_915);
nor U1025 (N_1025,N_956,N_963);
or U1026 (N_1026,N_885,N_966);
or U1027 (N_1027,N_864,N_983);
and U1028 (N_1028,N_881,N_932);
nand U1029 (N_1029,N_852,N_961);
nor U1030 (N_1030,N_928,N_823);
nor U1031 (N_1031,N_902,N_814);
nor U1032 (N_1032,N_955,N_818);
and U1033 (N_1033,N_872,N_988);
and U1034 (N_1034,N_982,N_831);
and U1035 (N_1035,N_984,N_946);
nor U1036 (N_1036,N_883,N_913);
and U1037 (N_1037,N_822,N_861);
or U1038 (N_1038,N_929,N_948);
nor U1039 (N_1039,N_965,N_865);
xnor U1040 (N_1040,N_996,N_894);
nand U1041 (N_1041,N_830,N_892);
xor U1042 (N_1042,N_976,N_869);
or U1043 (N_1043,N_962,N_874);
nand U1044 (N_1044,N_808,N_924);
or U1045 (N_1045,N_947,N_847);
xnor U1046 (N_1046,N_825,N_879);
nand U1047 (N_1047,N_857,N_993);
and U1048 (N_1048,N_991,N_801);
nand U1049 (N_1049,N_817,N_806);
xor U1050 (N_1050,N_880,N_975);
or U1051 (N_1051,N_848,N_978);
nand U1052 (N_1052,N_938,N_829);
nor U1053 (N_1053,N_999,N_967);
xor U1054 (N_1054,N_868,N_972);
nor U1055 (N_1055,N_971,N_977);
nor U1056 (N_1056,N_908,N_828);
and U1057 (N_1057,N_803,N_951);
nand U1058 (N_1058,N_863,N_989);
and U1059 (N_1059,N_936,N_895);
nand U1060 (N_1060,N_891,N_935);
xnor U1061 (N_1061,N_819,N_901);
xor U1062 (N_1062,N_985,N_836);
or U1063 (N_1063,N_930,N_899);
nor U1064 (N_1064,N_838,N_870);
xnor U1065 (N_1065,N_859,N_997);
nor U1066 (N_1066,N_867,N_860);
xor U1067 (N_1067,N_890,N_812);
nor U1068 (N_1068,N_942,N_950);
and U1069 (N_1069,N_958,N_898);
xor U1070 (N_1070,N_844,N_960);
or U1071 (N_1071,N_906,N_893);
or U1072 (N_1072,N_839,N_979);
nand U1073 (N_1073,N_800,N_807);
nand U1074 (N_1074,N_925,N_888);
and U1075 (N_1075,N_834,N_900);
xnor U1076 (N_1076,N_877,N_922);
nand U1077 (N_1077,N_998,N_837);
xor U1078 (N_1078,N_827,N_973);
nor U1079 (N_1079,N_813,N_804);
and U1080 (N_1080,N_884,N_907);
nor U1081 (N_1081,N_826,N_926);
nand U1082 (N_1082,N_964,N_815);
and U1083 (N_1083,N_923,N_917);
nor U1084 (N_1084,N_820,N_802);
nor U1085 (N_1085,N_934,N_855);
nor U1086 (N_1086,N_810,N_919);
and U1087 (N_1087,N_824,N_949);
and U1088 (N_1088,N_944,N_943);
or U1089 (N_1089,N_909,N_927);
nand U1090 (N_1090,N_854,N_886);
or U1091 (N_1091,N_992,N_840);
or U1092 (N_1092,N_970,N_968);
and U1093 (N_1093,N_990,N_933);
xnor U1094 (N_1094,N_969,N_905);
xnor U1095 (N_1095,N_845,N_945);
nor U1096 (N_1096,N_835,N_981);
nor U1097 (N_1097,N_995,N_821);
xor U1098 (N_1098,N_850,N_873);
and U1099 (N_1099,N_918,N_911);
and U1100 (N_1100,N_976,N_941);
xnor U1101 (N_1101,N_822,N_860);
xor U1102 (N_1102,N_855,N_891);
xor U1103 (N_1103,N_819,N_891);
and U1104 (N_1104,N_893,N_942);
and U1105 (N_1105,N_856,N_881);
nor U1106 (N_1106,N_879,N_817);
nand U1107 (N_1107,N_921,N_914);
and U1108 (N_1108,N_922,N_882);
and U1109 (N_1109,N_925,N_986);
xor U1110 (N_1110,N_946,N_861);
xor U1111 (N_1111,N_810,N_997);
and U1112 (N_1112,N_920,N_831);
and U1113 (N_1113,N_829,N_995);
or U1114 (N_1114,N_999,N_912);
or U1115 (N_1115,N_978,N_961);
and U1116 (N_1116,N_995,N_924);
nand U1117 (N_1117,N_904,N_982);
nand U1118 (N_1118,N_845,N_900);
xnor U1119 (N_1119,N_961,N_933);
nand U1120 (N_1120,N_845,N_893);
and U1121 (N_1121,N_850,N_971);
or U1122 (N_1122,N_980,N_810);
xor U1123 (N_1123,N_892,N_957);
and U1124 (N_1124,N_901,N_848);
nor U1125 (N_1125,N_831,N_806);
xnor U1126 (N_1126,N_809,N_830);
nand U1127 (N_1127,N_892,N_966);
or U1128 (N_1128,N_975,N_887);
and U1129 (N_1129,N_984,N_841);
nand U1130 (N_1130,N_898,N_995);
xnor U1131 (N_1131,N_853,N_890);
xor U1132 (N_1132,N_848,N_823);
xor U1133 (N_1133,N_894,N_808);
nand U1134 (N_1134,N_884,N_903);
nand U1135 (N_1135,N_929,N_824);
or U1136 (N_1136,N_807,N_872);
xnor U1137 (N_1137,N_982,N_964);
or U1138 (N_1138,N_884,N_814);
or U1139 (N_1139,N_879,N_836);
xor U1140 (N_1140,N_894,N_814);
nor U1141 (N_1141,N_987,N_947);
nand U1142 (N_1142,N_953,N_939);
or U1143 (N_1143,N_981,N_992);
nand U1144 (N_1144,N_954,N_817);
nor U1145 (N_1145,N_871,N_959);
nand U1146 (N_1146,N_930,N_829);
or U1147 (N_1147,N_813,N_818);
and U1148 (N_1148,N_939,N_919);
and U1149 (N_1149,N_832,N_914);
nand U1150 (N_1150,N_930,N_995);
and U1151 (N_1151,N_923,N_997);
nand U1152 (N_1152,N_945,N_895);
xor U1153 (N_1153,N_912,N_929);
nor U1154 (N_1154,N_981,N_842);
or U1155 (N_1155,N_853,N_938);
nand U1156 (N_1156,N_885,N_868);
nand U1157 (N_1157,N_899,N_904);
and U1158 (N_1158,N_960,N_976);
or U1159 (N_1159,N_876,N_909);
or U1160 (N_1160,N_852,N_908);
and U1161 (N_1161,N_962,N_857);
or U1162 (N_1162,N_844,N_952);
and U1163 (N_1163,N_868,N_961);
and U1164 (N_1164,N_860,N_960);
xnor U1165 (N_1165,N_925,N_821);
and U1166 (N_1166,N_829,N_923);
or U1167 (N_1167,N_964,N_944);
xor U1168 (N_1168,N_875,N_924);
nor U1169 (N_1169,N_808,N_889);
nor U1170 (N_1170,N_827,N_993);
nand U1171 (N_1171,N_974,N_891);
nor U1172 (N_1172,N_816,N_887);
or U1173 (N_1173,N_964,N_939);
nand U1174 (N_1174,N_971,N_918);
or U1175 (N_1175,N_985,N_860);
xor U1176 (N_1176,N_965,N_989);
nor U1177 (N_1177,N_898,N_908);
nor U1178 (N_1178,N_930,N_901);
xnor U1179 (N_1179,N_868,N_870);
nor U1180 (N_1180,N_851,N_868);
nor U1181 (N_1181,N_840,N_859);
and U1182 (N_1182,N_833,N_919);
xnor U1183 (N_1183,N_802,N_953);
nor U1184 (N_1184,N_983,N_922);
nor U1185 (N_1185,N_849,N_942);
or U1186 (N_1186,N_929,N_967);
xnor U1187 (N_1187,N_828,N_935);
nor U1188 (N_1188,N_833,N_837);
or U1189 (N_1189,N_886,N_906);
nor U1190 (N_1190,N_987,N_855);
and U1191 (N_1191,N_961,N_869);
and U1192 (N_1192,N_954,N_923);
nand U1193 (N_1193,N_946,N_969);
and U1194 (N_1194,N_927,N_849);
nand U1195 (N_1195,N_803,N_808);
nand U1196 (N_1196,N_917,N_891);
and U1197 (N_1197,N_926,N_961);
nand U1198 (N_1198,N_843,N_995);
nand U1199 (N_1199,N_839,N_930);
and U1200 (N_1200,N_1062,N_1026);
xor U1201 (N_1201,N_1149,N_1098);
nand U1202 (N_1202,N_1089,N_1183);
xor U1203 (N_1203,N_1068,N_1064);
and U1204 (N_1204,N_1143,N_1069);
nand U1205 (N_1205,N_1043,N_1017);
xor U1206 (N_1206,N_1138,N_1056);
nor U1207 (N_1207,N_1193,N_1086);
nor U1208 (N_1208,N_1165,N_1030);
or U1209 (N_1209,N_1004,N_1097);
or U1210 (N_1210,N_1073,N_1019);
and U1211 (N_1211,N_1035,N_1197);
nand U1212 (N_1212,N_1101,N_1013);
or U1213 (N_1213,N_1157,N_1127);
nor U1214 (N_1214,N_1132,N_1095);
nand U1215 (N_1215,N_1119,N_1159);
and U1216 (N_1216,N_1071,N_1052);
xor U1217 (N_1217,N_1114,N_1009);
xor U1218 (N_1218,N_1074,N_1185);
nand U1219 (N_1219,N_1025,N_1146);
xnor U1220 (N_1220,N_1042,N_1198);
xnor U1221 (N_1221,N_1006,N_1135);
nor U1222 (N_1222,N_1134,N_1072);
xor U1223 (N_1223,N_1172,N_1126);
and U1224 (N_1224,N_1037,N_1090);
and U1225 (N_1225,N_1173,N_1100);
or U1226 (N_1226,N_1049,N_1021);
and U1227 (N_1227,N_1000,N_1192);
xnor U1228 (N_1228,N_1137,N_1170);
nand U1229 (N_1229,N_1094,N_1187);
xnor U1230 (N_1230,N_1080,N_1015);
nand U1231 (N_1231,N_1194,N_1048);
or U1232 (N_1232,N_1005,N_1178);
xor U1233 (N_1233,N_1024,N_1123);
nor U1234 (N_1234,N_1140,N_1020);
and U1235 (N_1235,N_1148,N_1113);
or U1236 (N_1236,N_1115,N_1151);
xnor U1237 (N_1237,N_1153,N_1182);
xor U1238 (N_1238,N_1168,N_1029);
or U1239 (N_1239,N_1108,N_1063);
xor U1240 (N_1240,N_1033,N_1003);
nand U1241 (N_1241,N_1107,N_1103);
and U1242 (N_1242,N_1083,N_1016);
and U1243 (N_1243,N_1070,N_1058);
and U1244 (N_1244,N_1184,N_1053);
xnor U1245 (N_1245,N_1039,N_1120);
or U1246 (N_1246,N_1117,N_1139);
nor U1247 (N_1247,N_1175,N_1136);
xnor U1248 (N_1248,N_1106,N_1181);
and U1249 (N_1249,N_1162,N_1038);
and U1250 (N_1250,N_1079,N_1188);
nand U1251 (N_1251,N_1023,N_1014);
xnor U1252 (N_1252,N_1160,N_1131);
and U1253 (N_1253,N_1196,N_1142);
and U1254 (N_1254,N_1018,N_1105);
or U1255 (N_1255,N_1176,N_1096);
or U1256 (N_1256,N_1189,N_1034);
and U1257 (N_1257,N_1118,N_1116);
nand U1258 (N_1258,N_1154,N_1028);
or U1259 (N_1259,N_1047,N_1166);
nor U1260 (N_1260,N_1190,N_1133);
xor U1261 (N_1261,N_1010,N_1167);
nor U1262 (N_1262,N_1044,N_1040);
nor U1263 (N_1263,N_1102,N_1060);
nor U1264 (N_1264,N_1082,N_1124);
xor U1265 (N_1265,N_1195,N_1001);
nand U1266 (N_1266,N_1059,N_1121);
xor U1267 (N_1267,N_1144,N_1085);
nor U1268 (N_1268,N_1177,N_1051);
nand U1269 (N_1269,N_1055,N_1128);
or U1270 (N_1270,N_1066,N_1174);
xor U1271 (N_1271,N_1179,N_1088);
or U1272 (N_1272,N_1156,N_1150);
xor U1273 (N_1273,N_1099,N_1031);
nor U1274 (N_1274,N_1130,N_1111);
and U1275 (N_1275,N_1067,N_1041);
xnor U1276 (N_1276,N_1022,N_1036);
or U1277 (N_1277,N_1012,N_1191);
or U1278 (N_1278,N_1161,N_1169);
and U1279 (N_1279,N_1158,N_1141);
and U1280 (N_1280,N_1045,N_1199);
and U1281 (N_1281,N_1050,N_1164);
xnor U1282 (N_1282,N_1078,N_1152);
nor U1283 (N_1283,N_1046,N_1077);
or U1284 (N_1284,N_1180,N_1007);
nor U1285 (N_1285,N_1110,N_1125);
and U1286 (N_1286,N_1054,N_1087);
nor U1287 (N_1287,N_1122,N_1084);
or U1288 (N_1288,N_1104,N_1109);
and U1289 (N_1289,N_1112,N_1008);
nand U1290 (N_1290,N_1145,N_1129);
or U1291 (N_1291,N_1065,N_1155);
or U1292 (N_1292,N_1147,N_1091);
nor U1293 (N_1293,N_1186,N_1002);
or U1294 (N_1294,N_1027,N_1092);
or U1295 (N_1295,N_1163,N_1171);
and U1296 (N_1296,N_1081,N_1011);
nand U1297 (N_1297,N_1075,N_1032);
or U1298 (N_1298,N_1061,N_1057);
nand U1299 (N_1299,N_1076,N_1093);
and U1300 (N_1300,N_1034,N_1192);
nor U1301 (N_1301,N_1141,N_1067);
or U1302 (N_1302,N_1191,N_1045);
and U1303 (N_1303,N_1162,N_1195);
xnor U1304 (N_1304,N_1198,N_1193);
nand U1305 (N_1305,N_1041,N_1092);
xnor U1306 (N_1306,N_1068,N_1028);
xnor U1307 (N_1307,N_1176,N_1005);
nand U1308 (N_1308,N_1181,N_1057);
and U1309 (N_1309,N_1138,N_1114);
nand U1310 (N_1310,N_1068,N_1199);
or U1311 (N_1311,N_1135,N_1065);
and U1312 (N_1312,N_1021,N_1131);
or U1313 (N_1313,N_1158,N_1163);
xnor U1314 (N_1314,N_1001,N_1002);
and U1315 (N_1315,N_1004,N_1016);
xnor U1316 (N_1316,N_1069,N_1071);
nor U1317 (N_1317,N_1039,N_1065);
nor U1318 (N_1318,N_1124,N_1015);
and U1319 (N_1319,N_1030,N_1031);
nand U1320 (N_1320,N_1030,N_1069);
and U1321 (N_1321,N_1035,N_1103);
or U1322 (N_1322,N_1117,N_1008);
or U1323 (N_1323,N_1052,N_1188);
and U1324 (N_1324,N_1011,N_1034);
nand U1325 (N_1325,N_1100,N_1106);
nor U1326 (N_1326,N_1193,N_1083);
nor U1327 (N_1327,N_1112,N_1127);
and U1328 (N_1328,N_1197,N_1139);
or U1329 (N_1329,N_1050,N_1184);
and U1330 (N_1330,N_1164,N_1084);
or U1331 (N_1331,N_1072,N_1199);
xor U1332 (N_1332,N_1108,N_1049);
nor U1333 (N_1333,N_1102,N_1195);
nor U1334 (N_1334,N_1008,N_1170);
nand U1335 (N_1335,N_1159,N_1151);
nor U1336 (N_1336,N_1169,N_1138);
and U1337 (N_1337,N_1125,N_1095);
and U1338 (N_1338,N_1037,N_1105);
nand U1339 (N_1339,N_1122,N_1096);
or U1340 (N_1340,N_1081,N_1198);
or U1341 (N_1341,N_1188,N_1159);
nand U1342 (N_1342,N_1026,N_1140);
or U1343 (N_1343,N_1102,N_1027);
or U1344 (N_1344,N_1000,N_1070);
and U1345 (N_1345,N_1023,N_1143);
nor U1346 (N_1346,N_1118,N_1039);
xnor U1347 (N_1347,N_1104,N_1191);
xor U1348 (N_1348,N_1164,N_1126);
and U1349 (N_1349,N_1041,N_1036);
and U1350 (N_1350,N_1003,N_1127);
and U1351 (N_1351,N_1052,N_1121);
nor U1352 (N_1352,N_1143,N_1018);
xnor U1353 (N_1353,N_1145,N_1093);
and U1354 (N_1354,N_1029,N_1078);
nor U1355 (N_1355,N_1189,N_1056);
nand U1356 (N_1356,N_1085,N_1154);
nand U1357 (N_1357,N_1175,N_1070);
nand U1358 (N_1358,N_1000,N_1037);
or U1359 (N_1359,N_1118,N_1031);
xnor U1360 (N_1360,N_1066,N_1198);
nor U1361 (N_1361,N_1199,N_1196);
or U1362 (N_1362,N_1010,N_1066);
and U1363 (N_1363,N_1112,N_1150);
nor U1364 (N_1364,N_1148,N_1014);
or U1365 (N_1365,N_1101,N_1080);
or U1366 (N_1366,N_1025,N_1117);
and U1367 (N_1367,N_1057,N_1026);
nor U1368 (N_1368,N_1015,N_1001);
nor U1369 (N_1369,N_1043,N_1127);
and U1370 (N_1370,N_1199,N_1176);
nand U1371 (N_1371,N_1034,N_1053);
nor U1372 (N_1372,N_1033,N_1058);
xor U1373 (N_1373,N_1080,N_1017);
xor U1374 (N_1374,N_1196,N_1094);
xnor U1375 (N_1375,N_1088,N_1007);
or U1376 (N_1376,N_1183,N_1035);
xor U1377 (N_1377,N_1074,N_1095);
nand U1378 (N_1378,N_1048,N_1081);
nand U1379 (N_1379,N_1035,N_1158);
or U1380 (N_1380,N_1090,N_1123);
nand U1381 (N_1381,N_1187,N_1168);
or U1382 (N_1382,N_1032,N_1098);
and U1383 (N_1383,N_1171,N_1025);
nand U1384 (N_1384,N_1127,N_1085);
or U1385 (N_1385,N_1168,N_1036);
xnor U1386 (N_1386,N_1062,N_1049);
nor U1387 (N_1387,N_1109,N_1123);
and U1388 (N_1388,N_1047,N_1071);
nand U1389 (N_1389,N_1152,N_1199);
or U1390 (N_1390,N_1094,N_1082);
nor U1391 (N_1391,N_1126,N_1051);
xor U1392 (N_1392,N_1136,N_1195);
xor U1393 (N_1393,N_1123,N_1035);
nor U1394 (N_1394,N_1010,N_1139);
nand U1395 (N_1395,N_1097,N_1167);
or U1396 (N_1396,N_1030,N_1191);
or U1397 (N_1397,N_1082,N_1149);
xnor U1398 (N_1398,N_1011,N_1019);
nor U1399 (N_1399,N_1149,N_1052);
nor U1400 (N_1400,N_1317,N_1207);
nor U1401 (N_1401,N_1287,N_1298);
xor U1402 (N_1402,N_1372,N_1235);
nor U1403 (N_1403,N_1376,N_1387);
xor U1404 (N_1404,N_1234,N_1290);
nand U1405 (N_1405,N_1327,N_1389);
nand U1406 (N_1406,N_1245,N_1229);
nand U1407 (N_1407,N_1244,N_1388);
and U1408 (N_1408,N_1300,N_1340);
and U1409 (N_1409,N_1237,N_1370);
nand U1410 (N_1410,N_1253,N_1367);
and U1411 (N_1411,N_1261,N_1307);
xor U1412 (N_1412,N_1220,N_1304);
and U1413 (N_1413,N_1267,N_1275);
nor U1414 (N_1414,N_1201,N_1284);
or U1415 (N_1415,N_1329,N_1277);
and U1416 (N_1416,N_1316,N_1319);
xnor U1417 (N_1417,N_1301,N_1215);
nor U1418 (N_1418,N_1364,N_1398);
xnor U1419 (N_1419,N_1305,N_1233);
nand U1420 (N_1420,N_1224,N_1303);
and U1421 (N_1421,N_1283,N_1213);
or U1422 (N_1422,N_1365,N_1390);
nand U1423 (N_1423,N_1369,N_1271);
or U1424 (N_1424,N_1204,N_1205);
nand U1425 (N_1425,N_1252,N_1243);
nand U1426 (N_1426,N_1339,N_1276);
and U1427 (N_1427,N_1363,N_1256);
xnor U1428 (N_1428,N_1313,N_1306);
nor U1429 (N_1429,N_1251,N_1209);
or U1430 (N_1430,N_1315,N_1236);
nand U1431 (N_1431,N_1357,N_1285);
and U1432 (N_1432,N_1248,N_1335);
nor U1433 (N_1433,N_1366,N_1362);
or U1434 (N_1434,N_1217,N_1297);
and U1435 (N_1435,N_1324,N_1318);
nor U1436 (N_1436,N_1348,N_1343);
or U1437 (N_1437,N_1383,N_1247);
or U1438 (N_1438,N_1344,N_1399);
xor U1439 (N_1439,N_1231,N_1295);
and U1440 (N_1440,N_1241,N_1240);
or U1441 (N_1441,N_1311,N_1296);
xor U1442 (N_1442,N_1395,N_1242);
or U1443 (N_1443,N_1333,N_1264);
and U1444 (N_1444,N_1352,N_1336);
and U1445 (N_1445,N_1226,N_1354);
nor U1446 (N_1446,N_1259,N_1384);
nand U1447 (N_1447,N_1223,N_1393);
and U1448 (N_1448,N_1396,N_1230);
nand U1449 (N_1449,N_1227,N_1374);
nor U1450 (N_1450,N_1214,N_1254);
and U1451 (N_1451,N_1342,N_1265);
or U1452 (N_1452,N_1282,N_1210);
nand U1453 (N_1453,N_1381,N_1239);
xnor U1454 (N_1454,N_1211,N_1375);
nand U1455 (N_1455,N_1349,N_1299);
nand U1456 (N_1456,N_1377,N_1257);
and U1457 (N_1457,N_1216,N_1255);
and U1458 (N_1458,N_1280,N_1378);
and U1459 (N_1459,N_1379,N_1302);
nor U1460 (N_1460,N_1310,N_1358);
xnor U1461 (N_1461,N_1206,N_1391);
xor U1462 (N_1462,N_1320,N_1273);
or U1463 (N_1463,N_1212,N_1222);
nor U1464 (N_1464,N_1292,N_1380);
nand U1465 (N_1465,N_1382,N_1356);
nor U1466 (N_1466,N_1328,N_1326);
xnor U1467 (N_1467,N_1373,N_1385);
nor U1468 (N_1468,N_1394,N_1269);
nor U1469 (N_1469,N_1322,N_1351);
or U1470 (N_1470,N_1294,N_1323);
nand U1471 (N_1471,N_1225,N_1359);
or U1472 (N_1472,N_1350,N_1334);
xnor U1473 (N_1473,N_1325,N_1361);
or U1474 (N_1474,N_1386,N_1321);
xor U1475 (N_1475,N_1314,N_1258);
or U1476 (N_1476,N_1203,N_1221);
nand U1477 (N_1477,N_1392,N_1368);
or U1478 (N_1478,N_1347,N_1200);
xnor U1479 (N_1479,N_1345,N_1338);
or U1480 (N_1480,N_1263,N_1272);
nor U1481 (N_1481,N_1289,N_1278);
and U1482 (N_1482,N_1341,N_1288);
nor U1483 (N_1483,N_1218,N_1228);
and U1484 (N_1484,N_1270,N_1337);
xnor U1485 (N_1485,N_1202,N_1293);
or U1486 (N_1486,N_1262,N_1397);
or U1487 (N_1487,N_1308,N_1279);
and U1488 (N_1488,N_1219,N_1232);
or U1489 (N_1489,N_1346,N_1360);
or U1490 (N_1490,N_1250,N_1249);
or U1491 (N_1491,N_1281,N_1312);
xnor U1492 (N_1492,N_1208,N_1371);
nor U1493 (N_1493,N_1268,N_1260);
nand U1494 (N_1494,N_1246,N_1286);
xor U1495 (N_1495,N_1309,N_1274);
nor U1496 (N_1496,N_1291,N_1355);
and U1497 (N_1497,N_1238,N_1330);
and U1498 (N_1498,N_1266,N_1332);
nand U1499 (N_1499,N_1331,N_1353);
or U1500 (N_1500,N_1212,N_1261);
nor U1501 (N_1501,N_1245,N_1356);
or U1502 (N_1502,N_1363,N_1264);
or U1503 (N_1503,N_1345,N_1208);
xnor U1504 (N_1504,N_1294,N_1265);
nor U1505 (N_1505,N_1366,N_1237);
xor U1506 (N_1506,N_1348,N_1290);
or U1507 (N_1507,N_1243,N_1222);
nand U1508 (N_1508,N_1373,N_1302);
and U1509 (N_1509,N_1230,N_1378);
or U1510 (N_1510,N_1360,N_1272);
and U1511 (N_1511,N_1214,N_1235);
and U1512 (N_1512,N_1289,N_1368);
and U1513 (N_1513,N_1268,N_1274);
nor U1514 (N_1514,N_1299,N_1232);
nand U1515 (N_1515,N_1375,N_1338);
or U1516 (N_1516,N_1393,N_1349);
xnor U1517 (N_1517,N_1331,N_1388);
or U1518 (N_1518,N_1318,N_1250);
xor U1519 (N_1519,N_1277,N_1227);
and U1520 (N_1520,N_1201,N_1339);
and U1521 (N_1521,N_1262,N_1309);
nor U1522 (N_1522,N_1396,N_1213);
or U1523 (N_1523,N_1263,N_1398);
and U1524 (N_1524,N_1270,N_1216);
and U1525 (N_1525,N_1205,N_1322);
xor U1526 (N_1526,N_1220,N_1309);
and U1527 (N_1527,N_1275,N_1222);
nor U1528 (N_1528,N_1225,N_1268);
nand U1529 (N_1529,N_1206,N_1255);
nor U1530 (N_1530,N_1264,N_1262);
and U1531 (N_1531,N_1210,N_1354);
and U1532 (N_1532,N_1320,N_1265);
and U1533 (N_1533,N_1383,N_1333);
xnor U1534 (N_1534,N_1347,N_1305);
nor U1535 (N_1535,N_1379,N_1342);
xor U1536 (N_1536,N_1202,N_1261);
or U1537 (N_1537,N_1399,N_1291);
or U1538 (N_1538,N_1202,N_1283);
nand U1539 (N_1539,N_1301,N_1277);
and U1540 (N_1540,N_1286,N_1267);
xnor U1541 (N_1541,N_1239,N_1304);
and U1542 (N_1542,N_1279,N_1252);
nand U1543 (N_1543,N_1312,N_1364);
and U1544 (N_1544,N_1303,N_1381);
xnor U1545 (N_1545,N_1308,N_1288);
and U1546 (N_1546,N_1386,N_1360);
and U1547 (N_1547,N_1315,N_1296);
and U1548 (N_1548,N_1368,N_1219);
and U1549 (N_1549,N_1287,N_1321);
or U1550 (N_1550,N_1293,N_1358);
nor U1551 (N_1551,N_1306,N_1297);
xor U1552 (N_1552,N_1280,N_1388);
xnor U1553 (N_1553,N_1286,N_1265);
nand U1554 (N_1554,N_1272,N_1306);
xnor U1555 (N_1555,N_1216,N_1264);
xor U1556 (N_1556,N_1344,N_1232);
xor U1557 (N_1557,N_1212,N_1335);
xnor U1558 (N_1558,N_1284,N_1356);
nor U1559 (N_1559,N_1289,N_1252);
xnor U1560 (N_1560,N_1312,N_1236);
nand U1561 (N_1561,N_1208,N_1381);
or U1562 (N_1562,N_1293,N_1324);
and U1563 (N_1563,N_1210,N_1367);
nor U1564 (N_1564,N_1323,N_1303);
nor U1565 (N_1565,N_1362,N_1381);
or U1566 (N_1566,N_1227,N_1282);
xnor U1567 (N_1567,N_1256,N_1302);
xnor U1568 (N_1568,N_1331,N_1308);
and U1569 (N_1569,N_1340,N_1235);
and U1570 (N_1570,N_1212,N_1284);
and U1571 (N_1571,N_1263,N_1380);
or U1572 (N_1572,N_1293,N_1221);
xnor U1573 (N_1573,N_1214,N_1260);
or U1574 (N_1574,N_1301,N_1212);
or U1575 (N_1575,N_1312,N_1265);
nand U1576 (N_1576,N_1391,N_1252);
xor U1577 (N_1577,N_1292,N_1363);
nor U1578 (N_1578,N_1249,N_1375);
or U1579 (N_1579,N_1277,N_1232);
nor U1580 (N_1580,N_1230,N_1206);
nor U1581 (N_1581,N_1390,N_1262);
or U1582 (N_1582,N_1284,N_1361);
nand U1583 (N_1583,N_1333,N_1399);
xnor U1584 (N_1584,N_1387,N_1314);
nand U1585 (N_1585,N_1297,N_1349);
xnor U1586 (N_1586,N_1359,N_1360);
nand U1587 (N_1587,N_1217,N_1280);
or U1588 (N_1588,N_1240,N_1297);
xor U1589 (N_1589,N_1356,N_1318);
nand U1590 (N_1590,N_1200,N_1284);
and U1591 (N_1591,N_1204,N_1312);
nand U1592 (N_1592,N_1395,N_1275);
and U1593 (N_1593,N_1244,N_1358);
and U1594 (N_1594,N_1229,N_1238);
nor U1595 (N_1595,N_1274,N_1334);
xnor U1596 (N_1596,N_1283,N_1378);
and U1597 (N_1597,N_1319,N_1209);
nand U1598 (N_1598,N_1313,N_1394);
nor U1599 (N_1599,N_1239,N_1229);
nor U1600 (N_1600,N_1433,N_1427);
nor U1601 (N_1601,N_1570,N_1406);
nor U1602 (N_1602,N_1405,N_1552);
nand U1603 (N_1603,N_1424,N_1585);
or U1604 (N_1604,N_1498,N_1574);
and U1605 (N_1605,N_1537,N_1509);
and U1606 (N_1606,N_1512,N_1468);
and U1607 (N_1607,N_1402,N_1593);
or U1608 (N_1608,N_1418,N_1588);
or U1609 (N_1609,N_1556,N_1571);
xnor U1610 (N_1610,N_1408,N_1457);
and U1611 (N_1611,N_1454,N_1489);
xor U1612 (N_1612,N_1583,N_1425);
and U1613 (N_1613,N_1526,N_1500);
nand U1614 (N_1614,N_1459,N_1482);
xor U1615 (N_1615,N_1569,N_1563);
xor U1616 (N_1616,N_1466,N_1463);
xnor U1617 (N_1617,N_1525,N_1437);
nor U1618 (N_1618,N_1524,N_1496);
and U1619 (N_1619,N_1493,N_1404);
nand U1620 (N_1620,N_1444,N_1484);
xor U1621 (N_1621,N_1415,N_1547);
xnor U1622 (N_1622,N_1590,N_1460);
xor U1623 (N_1623,N_1486,N_1565);
nor U1624 (N_1624,N_1573,N_1551);
nor U1625 (N_1625,N_1452,N_1520);
nor U1626 (N_1626,N_1548,N_1472);
nand U1627 (N_1627,N_1453,N_1411);
or U1628 (N_1628,N_1501,N_1532);
nor U1629 (N_1629,N_1555,N_1580);
nor U1630 (N_1630,N_1464,N_1592);
xnor U1631 (N_1631,N_1403,N_1518);
nor U1632 (N_1632,N_1490,N_1533);
and U1633 (N_1633,N_1455,N_1510);
nand U1634 (N_1634,N_1462,N_1440);
nor U1635 (N_1635,N_1523,N_1575);
xnor U1636 (N_1636,N_1499,N_1587);
xnor U1637 (N_1637,N_1446,N_1430);
nor U1638 (N_1638,N_1560,N_1538);
nand U1639 (N_1639,N_1449,N_1502);
xor U1640 (N_1640,N_1572,N_1550);
and U1641 (N_1641,N_1544,N_1407);
or U1642 (N_1642,N_1485,N_1535);
nand U1643 (N_1643,N_1599,N_1409);
and U1644 (N_1644,N_1469,N_1432);
xnor U1645 (N_1645,N_1400,N_1507);
and U1646 (N_1646,N_1562,N_1494);
and U1647 (N_1647,N_1594,N_1516);
and U1648 (N_1648,N_1578,N_1577);
xor U1649 (N_1649,N_1504,N_1595);
nand U1650 (N_1650,N_1428,N_1441);
nand U1651 (N_1651,N_1456,N_1439);
xor U1652 (N_1652,N_1567,N_1536);
nand U1653 (N_1653,N_1417,N_1442);
xor U1654 (N_1654,N_1519,N_1545);
or U1655 (N_1655,N_1508,N_1549);
nand U1656 (N_1656,N_1530,N_1491);
nor U1657 (N_1657,N_1438,N_1421);
xnor U1658 (N_1658,N_1445,N_1554);
xor U1659 (N_1659,N_1443,N_1434);
or U1660 (N_1660,N_1476,N_1426);
or U1661 (N_1661,N_1558,N_1447);
nor U1662 (N_1662,N_1461,N_1506);
nor U1663 (N_1663,N_1413,N_1475);
and U1664 (N_1664,N_1470,N_1521);
nor U1665 (N_1665,N_1488,N_1513);
xor U1666 (N_1666,N_1465,N_1511);
xnor U1667 (N_1667,N_1422,N_1596);
or U1668 (N_1668,N_1522,N_1477);
nand U1669 (N_1669,N_1487,N_1528);
nand U1670 (N_1670,N_1480,N_1527);
nand U1671 (N_1671,N_1497,N_1581);
and U1672 (N_1672,N_1529,N_1531);
xnor U1673 (N_1673,N_1582,N_1553);
or U1674 (N_1674,N_1479,N_1557);
and U1675 (N_1675,N_1412,N_1517);
or U1676 (N_1676,N_1410,N_1514);
nand U1677 (N_1677,N_1435,N_1414);
and U1678 (N_1678,N_1561,N_1568);
and U1679 (N_1679,N_1597,N_1564);
nand U1680 (N_1680,N_1586,N_1579);
xor U1681 (N_1681,N_1566,N_1436);
or U1682 (N_1682,N_1458,N_1419);
xor U1683 (N_1683,N_1559,N_1505);
nand U1684 (N_1684,N_1542,N_1515);
or U1685 (N_1685,N_1598,N_1429);
or U1686 (N_1686,N_1546,N_1576);
or U1687 (N_1687,N_1451,N_1481);
nor U1688 (N_1688,N_1483,N_1495);
xnor U1689 (N_1689,N_1416,N_1591);
or U1690 (N_1690,N_1420,N_1473);
xor U1691 (N_1691,N_1471,N_1584);
nor U1692 (N_1692,N_1543,N_1540);
or U1693 (N_1693,N_1503,N_1539);
nand U1694 (N_1694,N_1589,N_1401);
nand U1695 (N_1695,N_1492,N_1450);
nand U1696 (N_1696,N_1474,N_1534);
nand U1697 (N_1697,N_1448,N_1467);
xor U1698 (N_1698,N_1423,N_1541);
or U1699 (N_1699,N_1431,N_1478);
nor U1700 (N_1700,N_1471,N_1506);
nand U1701 (N_1701,N_1465,N_1568);
or U1702 (N_1702,N_1408,N_1465);
nor U1703 (N_1703,N_1488,N_1451);
nand U1704 (N_1704,N_1539,N_1498);
xor U1705 (N_1705,N_1509,N_1439);
nor U1706 (N_1706,N_1592,N_1530);
xor U1707 (N_1707,N_1425,N_1569);
and U1708 (N_1708,N_1557,N_1553);
and U1709 (N_1709,N_1470,N_1515);
and U1710 (N_1710,N_1463,N_1501);
or U1711 (N_1711,N_1455,N_1509);
xor U1712 (N_1712,N_1411,N_1565);
or U1713 (N_1713,N_1427,N_1538);
or U1714 (N_1714,N_1529,N_1535);
nand U1715 (N_1715,N_1457,N_1581);
or U1716 (N_1716,N_1419,N_1599);
nand U1717 (N_1717,N_1510,N_1438);
nor U1718 (N_1718,N_1520,N_1411);
xor U1719 (N_1719,N_1581,N_1548);
nand U1720 (N_1720,N_1555,N_1585);
or U1721 (N_1721,N_1415,N_1418);
or U1722 (N_1722,N_1546,N_1566);
and U1723 (N_1723,N_1556,N_1453);
and U1724 (N_1724,N_1517,N_1403);
or U1725 (N_1725,N_1597,N_1433);
and U1726 (N_1726,N_1491,N_1587);
and U1727 (N_1727,N_1480,N_1464);
or U1728 (N_1728,N_1559,N_1406);
nor U1729 (N_1729,N_1445,N_1517);
nor U1730 (N_1730,N_1515,N_1558);
xor U1731 (N_1731,N_1475,N_1549);
and U1732 (N_1732,N_1523,N_1424);
nand U1733 (N_1733,N_1494,N_1458);
nand U1734 (N_1734,N_1542,N_1596);
nor U1735 (N_1735,N_1499,N_1578);
nand U1736 (N_1736,N_1501,N_1479);
nor U1737 (N_1737,N_1436,N_1577);
or U1738 (N_1738,N_1470,N_1504);
xor U1739 (N_1739,N_1406,N_1586);
or U1740 (N_1740,N_1580,N_1582);
and U1741 (N_1741,N_1441,N_1419);
nor U1742 (N_1742,N_1450,N_1504);
nor U1743 (N_1743,N_1403,N_1586);
nand U1744 (N_1744,N_1542,N_1449);
or U1745 (N_1745,N_1566,N_1477);
nand U1746 (N_1746,N_1508,N_1598);
nor U1747 (N_1747,N_1455,N_1586);
and U1748 (N_1748,N_1448,N_1506);
nand U1749 (N_1749,N_1525,N_1481);
xor U1750 (N_1750,N_1483,N_1408);
xnor U1751 (N_1751,N_1410,N_1523);
nand U1752 (N_1752,N_1446,N_1580);
and U1753 (N_1753,N_1502,N_1404);
nor U1754 (N_1754,N_1462,N_1418);
and U1755 (N_1755,N_1496,N_1448);
and U1756 (N_1756,N_1443,N_1446);
nand U1757 (N_1757,N_1470,N_1401);
nand U1758 (N_1758,N_1443,N_1502);
nand U1759 (N_1759,N_1558,N_1568);
xnor U1760 (N_1760,N_1435,N_1556);
nand U1761 (N_1761,N_1457,N_1594);
and U1762 (N_1762,N_1418,N_1576);
or U1763 (N_1763,N_1517,N_1486);
nand U1764 (N_1764,N_1547,N_1439);
or U1765 (N_1765,N_1498,N_1490);
or U1766 (N_1766,N_1439,N_1562);
xnor U1767 (N_1767,N_1464,N_1472);
and U1768 (N_1768,N_1417,N_1569);
and U1769 (N_1769,N_1448,N_1525);
or U1770 (N_1770,N_1452,N_1456);
or U1771 (N_1771,N_1501,N_1459);
nand U1772 (N_1772,N_1523,N_1496);
nand U1773 (N_1773,N_1532,N_1579);
nor U1774 (N_1774,N_1439,N_1519);
xnor U1775 (N_1775,N_1570,N_1434);
nand U1776 (N_1776,N_1400,N_1499);
or U1777 (N_1777,N_1401,N_1522);
and U1778 (N_1778,N_1561,N_1570);
and U1779 (N_1779,N_1589,N_1557);
nand U1780 (N_1780,N_1522,N_1598);
or U1781 (N_1781,N_1444,N_1426);
and U1782 (N_1782,N_1529,N_1482);
nor U1783 (N_1783,N_1536,N_1455);
or U1784 (N_1784,N_1404,N_1419);
or U1785 (N_1785,N_1431,N_1493);
xor U1786 (N_1786,N_1577,N_1509);
nor U1787 (N_1787,N_1491,N_1414);
xnor U1788 (N_1788,N_1538,N_1503);
or U1789 (N_1789,N_1597,N_1418);
or U1790 (N_1790,N_1585,N_1483);
and U1791 (N_1791,N_1451,N_1534);
and U1792 (N_1792,N_1415,N_1434);
xor U1793 (N_1793,N_1404,N_1476);
or U1794 (N_1794,N_1403,N_1474);
xnor U1795 (N_1795,N_1504,N_1502);
or U1796 (N_1796,N_1590,N_1552);
and U1797 (N_1797,N_1412,N_1545);
or U1798 (N_1798,N_1598,N_1545);
nor U1799 (N_1799,N_1495,N_1526);
and U1800 (N_1800,N_1655,N_1775);
and U1801 (N_1801,N_1739,N_1717);
or U1802 (N_1802,N_1632,N_1788);
nand U1803 (N_1803,N_1610,N_1732);
nor U1804 (N_1804,N_1631,N_1797);
xnor U1805 (N_1805,N_1718,N_1609);
and U1806 (N_1806,N_1798,N_1625);
or U1807 (N_1807,N_1623,N_1629);
nor U1808 (N_1808,N_1656,N_1628);
nand U1809 (N_1809,N_1689,N_1637);
nand U1810 (N_1810,N_1690,N_1607);
and U1811 (N_1811,N_1793,N_1639);
nand U1812 (N_1812,N_1773,N_1729);
nor U1813 (N_1813,N_1749,N_1666);
or U1814 (N_1814,N_1673,N_1756);
and U1815 (N_1815,N_1702,N_1722);
or U1816 (N_1816,N_1734,N_1707);
xor U1817 (N_1817,N_1752,N_1687);
and U1818 (N_1818,N_1693,N_1737);
nor U1819 (N_1819,N_1699,N_1755);
xnor U1820 (N_1820,N_1647,N_1649);
or U1821 (N_1821,N_1781,N_1665);
nor U1822 (N_1822,N_1611,N_1696);
nand U1823 (N_1823,N_1660,N_1671);
and U1824 (N_1824,N_1748,N_1680);
or U1825 (N_1825,N_1640,N_1743);
xor U1826 (N_1826,N_1713,N_1613);
xnor U1827 (N_1827,N_1771,N_1705);
or U1828 (N_1828,N_1731,N_1643);
and U1829 (N_1829,N_1764,N_1763);
or U1830 (N_1830,N_1683,N_1723);
nand U1831 (N_1831,N_1667,N_1700);
xor U1832 (N_1832,N_1777,N_1669);
xor U1833 (N_1833,N_1653,N_1697);
xor U1834 (N_1834,N_1612,N_1642);
nor U1835 (N_1835,N_1741,N_1728);
nor U1836 (N_1836,N_1636,N_1608);
xnor U1837 (N_1837,N_1716,N_1651);
and U1838 (N_1838,N_1709,N_1603);
nor U1839 (N_1839,N_1678,N_1715);
nor U1840 (N_1840,N_1691,N_1652);
nand U1841 (N_1841,N_1768,N_1638);
and U1842 (N_1842,N_1767,N_1796);
nand U1843 (N_1843,N_1626,N_1724);
xnor U1844 (N_1844,N_1658,N_1633);
nor U1845 (N_1845,N_1659,N_1782);
nor U1846 (N_1846,N_1604,N_1661);
nor U1847 (N_1847,N_1688,N_1674);
nor U1848 (N_1848,N_1686,N_1606);
or U1849 (N_1849,N_1645,N_1621);
nand U1850 (N_1850,N_1754,N_1605);
nor U1851 (N_1851,N_1618,N_1783);
and U1852 (N_1852,N_1784,N_1654);
xor U1853 (N_1853,N_1711,N_1634);
nand U1854 (N_1854,N_1779,N_1769);
xor U1855 (N_1855,N_1663,N_1670);
or U1856 (N_1856,N_1714,N_1774);
or U1857 (N_1857,N_1772,N_1706);
nor U1858 (N_1858,N_1792,N_1751);
xnor U1859 (N_1859,N_1794,N_1615);
nand U1860 (N_1860,N_1646,N_1712);
nor U1861 (N_1861,N_1770,N_1685);
or U1862 (N_1862,N_1692,N_1760);
nor U1863 (N_1863,N_1744,N_1622);
or U1864 (N_1864,N_1630,N_1727);
nor U1865 (N_1865,N_1644,N_1684);
nand U1866 (N_1866,N_1672,N_1635);
xnor U1867 (N_1867,N_1662,N_1791);
or U1868 (N_1868,N_1627,N_1790);
and U1869 (N_1869,N_1738,N_1761);
and U1870 (N_1870,N_1740,N_1776);
nor U1871 (N_1871,N_1600,N_1720);
and U1872 (N_1872,N_1725,N_1746);
nand U1873 (N_1873,N_1616,N_1762);
xnor U1874 (N_1874,N_1668,N_1648);
nor U1875 (N_1875,N_1745,N_1602);
nor U1876 (N_1876,N_1701,N_1726);
nor U1877 (N_1877,N_1795,N_1703);
nor U1878 (N_1878,N_1758,N_1733);
xor U1879 (N_1879,N_1679,N_1614);
xor U1880 (N_1880,N_1736,N_1682);
nor U1881 (N_1881,N_1780,N_1641);
and U1882 (N_1882,N_1708,N_1742);
nor U1883 (N_1883,N_1617,N_1799);
nor U1884 (N_1884,N_1619,N_1694);
and U1885 (N_1885,N_1765,N_1657);
or U1886 (N_1886,N_1786,N_1695);
nand U1887 (N_1887,N_1624,N_1710);
and U1888 (N_1888,N_1759,N_1620);
or U1889 (N_1889,N_1730,N_1719);
nand U1890 (N_1890,N_1664,N_1721);
nand U1891 (N_1891,N_1677,N_1778);
xor U1892 (N_1892,N_1735,N_1789);
and U1893 (N_1893,N_1675,N_1757);
or U1894 (N_1894,N_1676,N_1681);
and U1895 (N_1895,N_1750,N_1698);
or U1896 (N_1896,N_1753,N_1747);
or U1897 (N_1897,N_1601,N_1704);
nor U1898 (N_1898,N_1787,N_1785);
or U1899 (N_1899,N_1766,N_1650);
nand U1900 (N_1900,N_1702,N_1706);
and U1901 (N_1901,N_1795,N_1791);
nand U1902 (N_1902,N_1773,N_1733);
and U1903 (N_1903,N_1692,N_1745);
or U1904 (N_1904,N_1615,N_1624);
xnor U1905 (N_1905,N_1678,N_1637);
or U1906 (N_1906,N_1756,N_1759);
nand U1907 (N_1907,N_1708,N_1616);
and U1908 (N_1908,N_1674,N_1686);
nand U1909 (N_1909,N_1606,N_1683);
xor U1910 (N_1910,N_1718,N_1651);
xnor U1911 (N_1911,N_1744,N_1794);
and U1912 (N_1912,N_1684,N_1671);
or U1913 (N_1913,N_1732,N_1760);
xnor U1914 (N_1914,N_1682,N_1798);
xnor U1915 (N_1915,N_1701,N_1739);
xnor U1916 (N_1916,N_1723,N_1704);
or U1917 (N_1917,N_1752,N_1639);
and U1918 (N_1918,N_1685,N_1618);
or U1919 (N_1919,N_1785,N_1690);
nand U1920 (N_1920,N_1661,N_1690);
nor U1921 (N_1921,N_1789,N_1625);
and U1922 (N_1922,N_1689,N_1797);
or U1923 (N_1923,N_1788,N_1668);
or U1924 (N_1924,N_1638,N_1796);
and U1925 (N_1925,N_1791,N_1615);
nand U1926 (N_1926,N_1602,N_1640);
xnor U1927 (N_1927,N_1791,N_1683);
nand U1928 (N_1928,N_1690,N_1796);
xor U1929 (N_1929,N_1653,N_1760);
xnor U1930 (N_1930,N_1716,N_1686);
xnor U1931 (N_1931,N_1640,N_1643);
or U1932 (N_1932,N_1724,N_1742);
nand U1933 (N_1933,N_1786,N_1657);
nor U1934 (N_1934,N_1629,N_1780);
or U1935 (N_1935,N_1601,N_1638);
or U1936 (N_1936,N_1745,N_1765);
and U1937 (N_1937,N_1625,N_1619);
or U1938 (N_1938,N_1660,N_1688);
or U1939 (N_1939,N_1613,N_1682);
and U1940 (N_1940,N_1606,N_1650);
nand U1941 (N_1941,N_1753,N_1662);
nand U1942 (N_1942,N_1781,N_1663);
and U1943 (N_1943,N_1688,N_1706);
nand U1944 (N_1944,N_1621,N_1685);
nor U1945 (N_1945,N_1685,N_1745);
or U1946 (N_1946,N_1604,N_1773);
or U1947 (N_1947,N_1637,N_1762);
xor U1948 (N_1948,N_1665,N_1727);
nor U1949 (N_1949,N_1743,N_1783);
xnor U1950 (N_1950,N_1734,N_1785);
nand U1951 (N_1951,N_1779,N_1688);
and U1952 (N_1952,N_1784,N_1742);
and U1953 (N_1953,N_1654,N_1721);
xor U1954 (N_1954,N_1799,N_1630);
nor U1955 (N_1955,N_1761,N_1785);
nand U1956 (N_1956,N_1604,N_1638);
nand U1957 (N_1957,N_1614,N_1712);
xor U1958 (N_1958,N_1615,N_1604);
nand U1959 (N_1959,N_1707,N_1690);
or U1960 (N_1960,N_1722,N_1748);
and U1961 (N_1961,N_1647,N_1674);
nor U1962 (N_1962,N_1735,N_1725);
nand U1963 (N_1963,N_1683,N_1784);
nand U1964 (N_1964,N_1774,N_1696);
nor U1965 (N_1965,N_1601,N_1784);
xor U1966 (N_1966,N_1610,N_1650);
nor U1967 (N_1967,N_1641,N_1653);
or U1968 (N_1968,N_1719,N_1633);
nand U1969 (N_1969,N_1793,N_1725);
xnor U1970 (N_1970,N_1703,N_1601);
nor U1971 (N_1971,N_1779,N_1628);
xnor U1972 (N_1972,N_1673,N_1637);
or U1973 (N_1973,N_1771,N_1765);
nand U1974 (N_1974,N_1628,N_1606);
nor U1975 (N_1975,N_1715,N_1682);
xor U1976 (N_1976,N_1770,N_1774);
xnor U1977 (N_1977,N_1789,N_1660);
nand U1978 (N_1978,N_1717,N_1612);
xor U1979 (N_1979,N_1736,N_1616);
nand U1980 (N_1980,N_1759,N_1657);
and U1981 (N_1981,N_1783,N_1698);
xor U1982 (N_1982,N_1679,N_1658);
nor U1983 (N_1983,N_1616,N_1625);
nand U1984 (N_1984,N_1641,N_1765);
nor U1985 (N_1985,N_1701,N_1757);
nand U1986 (N_1986,N_1623,N_1703);
xnor U1987 (N_1987,N_1710,N_1751);
nand U1988 (N_1988,N_1770,N_1715);
nand U1989 (N_1989,N_1671,N_1685);
nor U1990 (N_1990,N_1613,N_1731);
nor U1991 (N_1991,N_1769,N_1696);
nand U1992 (N_1992,N_1631,N_1735);
xnor U1993 (N_1993,N_1729,N_1742);
and U1994 (N_1994,N_1786,N_1773);
or U1995 (N_1995,N_1646,N_1683);
and U1996 (N_1996,N_1600,N_1780);
nand U1997 (N_1997,N_1767,N_1610);
or U1998 (N_1998,N_1704,N_1655);
or U1999 (N_1999,N_1601,N_1676);
nand U2000 (N_2000,N_1822,N_1976);
or U2001 (N_2001,N_1869,N_1849);
nor U2002 (N_2002,N_1816,N_1885);
xor U2003 (N_2003,N_1858,N_1979);
nor U2004 (N_2004,N_1827,N_1866);
nor U2005 (N_2005,N_1810,N_1940);
nor U2006 (N_2006,N_1928,N_1930);
and U2007 (N_2007,N_1814,N_1909);
xor U2008 (N_2008,N_1874,N_1917);
or U2009 (N_2009,N_1932,N_1856);
nor U2010 (N_2010,N_1853,N_1995);
or U2011 (N_2011,N_1802,N_1936);
and U2012 (N_2012,N_1915,N_1873);
xor U2013 (N_2013,N_1913,N_1844);
and U2014 (N_2014,N_1835,N_1947);
nor U2015 (N_2015,N_1967,N_1883);
xnor U2016 (N_2016,N_1875,N_1884);
nor U2017 (N_2017,N_1811,N_1889);
nand U2018 (N_2018,N_1959,N_1993);
xor U2019 (N_2019,N_1933,N_1990);
and U2020 (N_2020,N_1965,N_1862);
nor U2021 (N_2021,N_1824,N_1978);
xor U2022 (N_2022,N_1899,N_1960);
nor U2023 (N_2023,N_1901,N_1969);
nand U2024 (N_2024,N_1872,N_1946);
or U2025 (N_2025,N_1961,N_1949);
nor U2026 (N_2026,N_1837,N_1803);
xor U2027 (N_2027,N_1954,N_1914);
and U2028 (N_2028,N_1958,N_1882);
xor U2029 (N_2029,N_1985,N_1854);
xor U2030 (N_2030,N_1941,N_1881);
or U2031 (N_2031,N_1921,N_1938);
nand U2032 (N_2032,N_1834,N_1939);
xnor U2033 (N_2033,N_1868,N_1876);
or U2034 (N_2034,N_1852,N_1905);
and U2035 (N_2035,N_1898,N_1839);
and U2036 (N_2036,N_1997,N_1871);
nand U2037 (N_2037,N_1804,N_1820);
xor U2038 (N_2038,N_1998,N_1867);
xor U2039 (N_2039,N_1815,N_1886);
nand U2040 (N_2040,N_1987,N_1999);
xor U2041 (N_2041,N_1847,N_1896);
nor U2042 (N_2042,N_1972,N_1974);
or U2043 (N_2043,N_1991,N_1966);
nor U2044 (N_2044,N_1956,N_1963);
xor U2045 (N_2045,N_1924,N_1906);
nand U2046 (N_2046,N_1908,N_1840);
nor U2047 (N_2047,N_1808,N_1937);
nor U2048 (N_2048,N_1911,N_1894);
or U2049 (N_2049,N_1929,N_1904);
xor U2050 (N_2050,N_1968,N_1984);
nor U2051 (N_2051,N_1846,N_1920);
nand U2052 (N_2052,N_1948,N_1870);
nand U2053 (N_2053,N_1813,N_1848);
and U2054 (N_2054,N_1831,N_1879);
or U2055 (N_2055,N_1880,N_1892);
or U2056 (N_2056,N_1994,N_1926);
and U2057 (N_2057,N_1895,N_1925);
nand U2058 (N_2058,N_1919,N_1829);
xnor U2059 (N_2059,N_1859,N_1857);
nand U2060 (N_2060,N_1893,N_1942);
nand U2061 (N_2061,N_1845,N_1897);
nand U2062 (N_2062,N_1833,N_1817);
nand U2063 (N_2063,N_1821,N_1981);
nand U2064 (N_2064,N_1982,N_1843);
and U2065 (N_2065,N_1916,N_1934);
or U2066 (N_2066,N_1912,N_1971);
nand U2067 (N_2067,N_1953,N_1865);
and U2068 (N_2068,N_1955,N_1950);
nand U2069 (N_2069,N_1992,N_1801);
nor U2070 (N_2070,N_1855,N_1973);
and U2071 (N_2071,N_1996,N_1828);
nand U2072 (N_2072,N_1935,N_1952);
nor U2073 (N_2073,N_1864,N_1975);
xnor U2074 (N_2074,N_1951,N_1836);
xor U2075 (N_2075,N_1923,N_1826);
or U2076 (N_2076,N_1805,N_1922);
xor U2077 (N_2077,N_1860,N_1988);
or U2078 (N_2078,N_1910,N_1891);
nand U2079 (N_2079,N_1842,N_1851);
and U2080 (N_2080,N_1863,N_1903);
nand U2081 (N_2081,N_1986,N_1825);
or U2082 (N_2082,N_1861,N_1943);
and U2083 (N_2083,N_1809,N_1877);
nand U2084 (N_2084,N_1819,N_1812);
xor U2085 (N_2085,N_1878,N_1980);
or U2086 (N_2086,N_1957,N_1970);
xor U2087 (N_2087,N_1944,N_1945);
or U2088 (N_2088,N_1962,N_1807);
or U2089 (N_2089,N_1850,N_1900);
or U2090 (N_2090,N_1902,N_1907);
nand U2091 (N_2091,N_1823,N_1977);
nand U2092 (N_2092,N_1983,N_1830);
nor U2093 (N_2093,N_1918,N_1841);
and U2094 (N_2094,N_1887,N_1927);
nand U2095 (N_2095,N_1888,N_1964);
or U2096 (N_2096,N_1890,N_1989);
or U2097 (N_2097,N_1832,N_1838);
nand U2098 (N_2098,N_1818,N_1806);
nor U2099 (N_2099,N_1931,N_1800);
and U2100 (N_2100,N_1939,N_1935);
nand U2101 (N_2101,N_1918,N_1965);
or U2102 (N_2102,N_1885,N_1957);
nor U2103 (N_2103,N_1868,N_1816);
nand U2104 (N_2104,N_1884,N_1956);
xnor U2105 (N_2105,N_1874,N_1945);
and U2106 (N_2106,N_1928,N_1967);
nand U2107 (N_2107,N_1988,N_1908);
nand U2108 (N_2108,N_1953,N_1972);
xor U2109 (N_2109,N_1817,N_1977);
or U2110 (N_2110,N_1936,N_1816);
and U2111 (N_2111,N_1805,N_1863);
nand U2112 (N_2112,N_1967,N_1850);
and U2113 (N_2113,N_1999,N_1882);
nor U2114 (N_2114,N_1870,N_1802);
nor U2115 (N_2115,N_1921,N_1987);
and U2116 (N_2116,N_1857,N_1936);
xor U2117 (N_2117,N_1896,N_1975);
nor U2118 (N_2118,N_1854,N_1852);
and U2119 (N_2119,N_1824,N_1939);
nand U2120 (N_2120,N_1829,N_1880);
xnor U2121 (N_2121,N_1992,N_1962);
nand U2122 (N_2122,N_1840,N_1978);
xor U2123 (N_2123,N_1989,N_1858);
and U2124 (N_2124,N_1874,N_1864);
nand U2125 (N_2125,N_1857,N_1830);
nand U2126 (N_2126,N_1874,N_1998);
xor U2127 (N_2127,N_1826,N_1822);
nand U2128 (N_2128,N_1985,N_1809);
or U2129 (N_2129,N_1946,N_1840);
and U2130 (N_2130,N_1996,N_1820);
xnor U2131 (N_2131,N_1900,N_1946);
nand U2132 (N_2132,N_1848,N_1957);
and U2133 (N_2133,N_1939,N_1811);
or U2134 (N_2134,N_1801,N_1996);
or U2135 (N_2135,N_1825,N_1949);
or U2136 (N_2136,N_1885,N_1869);
or U2137 (N_2137,N_1921,N_1974);
or U2138 (N_2138,N_1924,N_1936);
or U2139 (N_2139,N_1826,N_1858);
and U2140 (N_2140,N_1873,N_1800);
xor U2141 (N_2141,N_1866,N_1925);
nor U2142 (N_2142,N_1944,N_1989);
xnor U2143 (N_2143,N_1966,N_1915);
nor U2144 (N_2144,N_1832,N_1812);
or U2145 (N_2145,N_1871,N_1879);
or U2146 (N_2146,N_1991,N_1981);
or U2147 (N_2147,N_1870,N_1915);
xor U2148 (N_2148,N_1926,N_1827);
nand U2149 (N_2149,N_1908,N_1817);
xnor U2150 (N_2150,N_1863,N_1849);
or U2151 (N_2151,N_1931,N_1885);
nor U2152 (N_2152,N_1852,N_1803);
nand U2153 (N_2153,N_1862,N_1804);
or U2154 (N_2154,N_1995,N_1948);
and U2155 (N_2155,N_1948,N_1807);
or U2156 (N_2156,N_1914,N_1978);
nor U2157 (N_2157,N_1905,N_1817);
nand U2158 (N_2158,N_1871,N_1850);
and U2159 (N_2159,N_1999,N_1984);
xor U2160 (N_2160,N_1932,N_1974);
nor U2161 (N_2161,N_1885,N_1887);
nor U2162 (N_2162,N_1923,N_1857);
nand U2163 (N_2163,N_1814,N_1900);
nand U2164 (N_2164,N_1956,N_1918);
or U2165 (N_2165,N_1850,N_1874);
and U2166 (N_2166,N_1938,N_1859);
or U2167 (N_2167,N_1979,N_1960);
nand U2168 (N_2168,N_1934,N_1855);
or U2169 (N_2169,N_1801,N_1973);
nand U2170 (N_2170,N_1963,N_1938);
and U2171 (N_2171,N_1970,N_1904);
or U2172 (N_2172,N_1884,N_1808);
nor U2173 (N_2173,N_1938,N_1874);
nand U2174 (N_2174,N_1920,N_1886);
or U2175 (N_2175,N_1848,N_1956);
nand U2176 (N_2176,N_1992,N_1988);
nand U2177 (N_2177,N_1953,N_1976);
or U2178 (N_2178,N_1864,N_1825);
and U2179 (N_2179,N_1864,N_1899);
xor U2180 (N_2180,N_1966,N_1963);
xnor U2181 (N_2181,N_1815,N_1904);
nor U2182 (N_2182,N_1896,N_1995);
and U2183 (N_2183,N_1885,N_1886);
or U2184 (N_2184,N_1970,N_1991);
or U2185 (N_2185,N_1870,N_1958);
nand U2186 (N_2186,N_1900,N_1821);
and U2187 (N_2187,N_1935,N_1823);
or U2188 (N_2188,N_1912,N_1870);
or U2189 (N_2189,N_1873,N_1833);
nor U2190 (N_2190,N_1949,N_1932);
nor U2191 (N_2191,N_1992,N_1848);
and U2192 (N_2192,N_1988,N_1865);
nand U2193 (N_2193,N_1928,N_1936);
nand U2194 (N_2194,N_1899,N_1923);
nor U2195 (N_2195,N_1942,N_1963);
xnor U2196 (N_2196,N_1927,N_1968);
nor U2197 (N_2197,N_1942,N_1866);
nor U2198 (N_2198,N_1948,N_1833);
and U2199 (N_2199,N_1858,N_1982);
and U2200 (N_2200,N_2081,N_2039);
and U2201 (N_2201,N_2143,N_2130);
nor U2202 (N_2202,N_2051,N_2125);
xor U2203 (N_2203,N_2028,N_2122);
xor U2204 (N_2204,N_2004,N_2072);
and U2205 (N_2205,N_2007,N_2157);
nor U2206 (N_2206,N_2060,N_2038);
or U2207 (N_2207,N_2133,N_2080);
or U2208 (N_2208,N_2054,N_2131);
or U2209 (N_2209,N_2059,N_2018);
xor U2210 (N_2210,N_2178,N_2194);
nor U2211 (N_2211,N_2156,N_2005);
xor U2212 (N_2212,N_2033,N_2154);
nor U2213 (N_2213,N_2104,N_2041);
nor U2214 (N_2214,N_2098,N_2086);
and U2215 (N_2215,N_2047,N_2074);
or U2216 (N_2216,N_2010,N_2153);
nor U2217 (N_2217,N_2083,N_2031);
and U2218 (N_2218,N_2148,N_2069);
xor U2219 (N_2219,N_2030,N_2147);
nor U2220 (N_2220,N_2094,N_2021);
nand U2221 (N_2221,N_2076,N_2052);
nor U2222 (N_2222,N_2009,N_2128);
nand U2223 (N_2223,N_2106,N_2132);
nand U2224 (N_2224,N_2110,N_2056);
and U2225 (N_2225,N_2105,N_2196);
nand U2226 (N_2226,N_2102,N_2029);
nor U2227 (N_2227,N_2096,N_2090);
nand U2228 (N_2228,N_2100,N_2070);
nand U2229 (N_2229,N_2037,N_2036);
or U2230 (N_2230,N_2119,N_2162);
and U2231 (N_2231,N_2192,N_2167);
xnor U2232 (N_2232,N_2075,N_2176);
xnor U2233 (N_2233,N_2011,N_2191);
and U2234 (N_2234,N_2186,N_2113);
nand U2235 (N_2235,N_2181,N_2164);
nor U2236 (N_2236,N_2139,N_2180);
nand U2237 (N_2237,N_2062,N_2043);
nor U2238 (N_2238,N_2170,N_2103);
nand U2239 (N_2239,N_2198,N_2182);
nand U2240 (N_2240,N_2166,N_2095);
and U2241 (N_2241,N_2050,N_2114);
xnor U2242 (N_2242,N_2129,N_2013);
or U2243 (N_2243,N_2078,N_2158);
or U2244 (N_2244,N_2024,N_2188);
and U2245 (N_2245,N_2073,N_2014);
nand U2246 (N_2246,N_2115,N_2177);
nand U2247 (N_2247,N_2197,N_2032);
nor U2248 (N_2248,N_2002,N_2116);
nand U2249 (N_2249,N_2058,N_2082);
or U2250 (N_2250,N_2123,N_2149);
and U2251 (N_2251,N_2199,N_2173);
nor U2252 (N_2252,N_2184,N_2121);
nor U2253 (N_2253,N_2023,N_2183);
or U2254 (N_2254,N_2120,N_2112);
or U2255 (N_2255,N_2019,N_2045);
nand U2256 (N_2256,N_2000,N_2034);
xnor U2257 (N_2257,N_2109,N_2111);
nand U2258 (N_2258,N_2017,N_2093);
nand U2259 (N_2259,N_2084,N_2141);
nor U2260 (N_2260,N_2053,N_2142);
nand U2261 (N_2261,N_2160,N_2063);
xor U2262 (N_2262,N_2066,N_2161);
nor U2263 (N_2263,N_2126,N_2079);
nor U2264 (N_2264,N_2134,N_2144);
nor U2265 (N_2265,N_2174,N_2049);
nand U2266 (N_2266,N_2169,N_2136);
and U2267 (N_2267,N_2065,N_2087);
xnor U2268 (N_2268,N_2108,N_2145);
and U2269 (N_2269,N_2097,N_2187);
nor U2270 (N_2270,N_2118,N_2027);
nand U2271 (N_2271,N_2155,N_2171);
or U2272 (N_2272,N_2117,N_2064);
or U2273 (N_2273,N_2168,N_2046);
xor U2274 (N_2274,N_2048,N_2175);
and U2275 (N_2275,N_2193,N_2146);
nand U2276 (N_2276,N_2159,N_2138);
or U2277 (N_2277,N_2068,N_2088);
and U2278 (N_2278,N_2185,N_2040);
and U2279 (N_2279,N_2089,N_2001);
xor U2280 (N_2280,N_2016,N_2057);
and U2281 (N_2281,N_2042,N_2091);
and U2282 (N_2282,N_2107,N_2085);
and U2283 (N_2283,N_2150,N_2151);
nor U2284 (N_2284,N_2061,N_2101);
and U2285 (N_2285,N_2124,N_2003);
or U2286 (N_2286,N_2140,N_2165);
nand U2287 (N_2287,N_2152,N_2071);
xnor U2288 (N_2288,N_2135,N_2127);
nor U2289 (N_2289,N_2179,N_2189);
nand U2290 (N_2290,N_2022,N_2015);
nand U2291 (N_2291,N_2092,N_2172);
and U2292 (N_2292,N_2035,N_2163);
nor U2293 (N_2293,N_2190,N_2012);
nand U2294 (N_2294,N_2055,N_2067);
or U2295 (N_2295,N_2025,N_2006);
or U2296 (N_2296,N_2077,N_2026);
nor U2297 (N_2297,N_2195,N_2137);
or U2298 (N_2298,N_2099,N_2044);
and U2299 (N_2299,N_2020,N_2008);
and U2300 (N_2300,N_2136,N_2038);
or U2301 (N_2301,N_2016,N_2024);
and U2302 (N_2302,N_2022,N_2162);
xor U2303 (N_2303,N_2144,N_2067);
or U2304 (N_2304,N_2069,N_2138);
nand U2305 (N_2305,N_2098,N_2023);
nand U2306 (N_2306,N_2130,N_2144);
nor U2307 (N_2307,N_2046,N_2055);
nand U2308 (N_2308,N_2013,N_2157);
xor U2309 (N_2309,N_2061,N_2051);
nor U2310 (N_2310,N_2113,N_2053);
and U2311 (N_2311,N_2074,N_2112);
nor U2312 (N_2312,N_2158,N_2159);
xor U2313 (N_2313,N_2084,N_2161);
nand U2314 (N_2314,N_2034,N_2196);
and U2315 (N_2315,N_2066,N_2199);
or U2316 (N_2316,N_2122,N_2190);
xor U2317 (N_2317,N_2029,N_2124);
and U2318 (N_2318,N_2120,N_2113);
nor U2319 (N_2319,N_2038,N_2076);
nor U2320 (N_2320,N_2120,N_2117);
nand U2321 (N_2321,N_2127,N_2050);
nand U2322 (N_2322,N_2027,N_2154);
or U2323 (N_2323,N_2167,N_2000);
or U2324 (N_2324,N_2091,N_2026);
xor U2325 (N_2325,N_2186,N_2021);
nor U2326 (N_2326,N_2176,N_2108);
xor U2327 (N_2327,N_2026,N_2037);
and U2328 (N_2328,N_2050,N_2076);
and U2329 (N_2329,N_2136,N_2148);
nand U2330 (N_2330,N_2020,N_2130);
or U2331 (N_2331,N_2063,N_2054);
xor U2332 (N_2332,N_2150,N_2029);
nor U2333 (N_2333,N_2026,N_2082);
xor U2334 (N_2334,N_2132,N_2114);
or U2335 (N_2335,N_2078,N_2118);
nand U2336 (N_2336,N_2157,N_2057);
xnor U2337 (N_2337,N_2166,N_2148);
and U2338 (N_2338,N_2081,N_2186);
or U2339 (N_2339,N_2165,N_2142);
and U2340 (N_2340,N_2053,N_2148);
xor U2341 (N_2341,N_2171,N_2092);
and U2342 (N_2342,N_2068,N_2070);
or U2343 (N_2343,N_2086,N_2114);
nor U2344 (N_2344,N_2190,N_2196);
nand U2345 (N_2345,N_2045,N_2120);
xor U2346 (N_2346,N_2187,N_2101);
nand U2347 (N_2347,N_2002,N_2139);
nor U2348 (N_2348,N_2046,N_2193);
xnor U2349 (N_2349,N_2111,N_2162);
and U2350 (N_2350,N_2046,N_2187);
or U2351 (N_2351,N_2048,N_2055);
nor U2352 (N_2352,N_2007,N_2136);
nor U2353 (N_2353,N_2102,N_2090);
and U2354 (N_2354,N_2193,N_2081);
nand U2355 (N_2355,N_2135,N_2133);
or U2356 (N_2356,N_2137,N_2119);
and U2357 (N_2357,N_2061,N_2161);
nor U2358 (N_2358,N_2111,N_2114);
nand U2359 (N_2359,N_2099,N_2019);
xnor U2360 (N_2360,N_2035,N_2106);
or U2361 (N_2361,N_2139,N_2165);
nand U2362 (N_2362,N_2041,N_2076);
or U2363 (N_2363,N_2174,N_2075);
and U2364 (N_2364,N_2111,N_2027);
nor U2365 (N_2365,N_2179,N_2169);
nand U2366 (N_2366,N_2169,N_2036);
nor U2367 (N_2367,N_2041,N_2094);
nand U2368 (N_2368,N_2158,N_2050);
xor U2369 (N_2369,N_2001,N_2189);
nand U2370 (N_2370,N_2153,N_2052);
or U2371 (N_2371,N_2074,N_2065);
and U2372 (N_2372,N_2169,N_2067);
or U2373 (N_2373,N_2060,N_2027);
nand U2374 (N_2374,N_2079,N_2071);
and U2375 (N_2375,N_2143,N_2001);
xnor U2376 (N_2376,N_2017,N_2133);
nand U2377 (N_2377,N_2154,N_2050);
nand U2378 (N_2378,N_2009,N_2045);
nor U2379 (N_2379,N_2138,N_2149);
nand U2380 (N_2380,N_2008,N_2107);
nor U2381 (N_2381,N_2009,N_2019);
nor U2382 (N_2382,N_2168,N_2035);
nor U2383 (N_2383,N_2029,N_2082);
and U2384 (N_2384,N_2018,N_2044);
nor U2385 (N_2385,N_2009,N_2054);
and U2386 (N_2386,N_2078,N_2184);
and U2387 (N_2387,N_2059,N_2016);
xor U2388 (N_2388,N_2060,N_2021);
xnor U2389 (N_2389,N_2050,N_2013);
xnor U2390 (N_2390,N_2131,N_2081);
nor U2391 (N_2391,N_2105,N_2090);
nand U2392 (N_2392,N_2186,N_2083);
nand U2393 (N_2393,N_2179,N_2093);
or U2394 (N_2394,N_2043,N_2102);
nand U2395 (N_2395,N_2139,N_2029);
nand U2396 (N_2396,N_2133,N_2139);
nor U2397 (N_2397,N_2001,N_2023);
xnor U2398 (N_2398,N_2186,N_2071);
nor U2399 (N_2399,N_2049,N_2094);
and U2400 (N_2400,N_2250,N_2251);
nand U2401 (N_2401,N_2261,N_2233);
nand U2402 (N_2402,N_2334,N_2360);
nor U2403 (N_2403,N_2339,N_2206);
xnor U2404 (N_2404,N_2220,N_2388);
or U2405 (N_2405,N_2393,N_2211);
xor U2406 (N_2406,N_2293,N_2271);
nand U2407 (N_2407,N_2291,N_2312);
or U2408 (N_2408,N_2228,N_2346);
and U2409 (N_2409,N_2231,N_2280);
or U2410 (N_2410,N_2319,N_2387);
xor U2411 (N_2411,N_2239,N_2362);
xor U2412 (N_2412,N_2345,N_2236);
nand U2413 (N_2413,N_2370,N_2243);
nor U2414 (N_2414,N_2306,N_2369);
and U2415 (N_2415,N_2318,N_2273);
nand U2416 (N_2416,N_2287,N_2321);
and U2417 (N_2417,N_2230,N_2331);
and U2418 (N_2418,N_2323,N_2315);
or U2419 (N_2419,N_2340,N_2390);
nor U2420 (N_2420,N_2295,N_2214);
or U2421 (N_2421,N_2235,N_2299);
xor U2422 (N_2422,N_2292,N_2358);
and U2423 (N_2423,N_2378,N_2309);
nand U2424 (N_2424,N_2355,N_2352);
xnor U2425 (N_2425,N_2366,N_2373);
nor U2426 (N_2426,N_2217,N_2265);
nor U2427 (N_2427,N_2353,N_2224);
and U2428 (N_2428,N_2242,N_2308);
nand U2429 (N_2429,N_2269,N_2394);
nand U2430 (N_2430,N_2263,N_2210);
nor U2431 (N_2431,N_2262,N_2286);
xor U2432 (N_2432,N_2377,N_2347);
nand U2433 (N_2433,N_2254,N_2202);
or U2434 (N_2434,N_2344,N_2332);
nor U2435 (N_2435,N_2311,N_2255);
xnor U2436 (N_2436,N_2221,N_2303);
nor U2437 (N_2437,N_2281,N_2245);
or U2438 (N_2438,N_2335,N_2320);
and U2439 (N_2439,N_2244,N_2259);
xnor U2440 (N_2440,N_2257,N_2368);
nand U2441 (N_2441,N_2359,N_2266);
xor U2442 (N_2442,N_2307,N_2237);
nor U2443 (N_2443,N_2380,N_2276);
xor U2444 (N_2444,N_2213,N_2392);
nand U2445 (N_2445,N_2324,N_2326);
or U2446 (N_2446,N_2399,N_2215);
nor U2447 (N_2447,N_2225,N_2238);
nor U2448 (N_2448,N_2289,N_2357);
xnor U2449 (N_2449,N_2252,N_2205);
xor U2450 (N_2450,N_2301,N_2374);
xor U2451 (N_2451,N_2284,N_2201);
nand U2452 (N_2452,N_2338,N_2207);
xor U2453 (N_2453,N_2283,N_2372);
nand U2454 (N_2454,N_2395,N_2288);
nor U2455 (N_2455,N_2351,N_2267);
or U2456 (N_2456,N_2212,N_2364);
or U2457 (N_2457,N_2381,N_2337);
or U2458 (N_2458,N_2277,N_2328);
xnor U2459 (N_2459,N_2229,N_2296);
nand U2460 (N_2460,N_2365,N_2297);
nand U2461 (N_2461,N_2268,N_2219);
and U2462 (N_2462,N_2272,N_2305);
nand U2463 (N_2463,N_2376,N_2253);
nand U2464 (N_2464,N_2314,N_2200);
nor U2465 (N_2465,N_2216,N_2258);
xor U2466 (N_2466,N_2264,N_2397);
xor U2467 (N_2467,N_2218,N_2384);
and U2468 (N_2468,N_2232,N_2270);
nor U2469 (N_2469,N_2350,N_2398);
and U2470 (N_2470,N_2383,N_2385);
xnor U2471 (N_2471,N_2316,N_2313);
and U2472 (N_2472,N_2391,N_2325);
nand U2473 (N_2473,N_2222,N_2367);
xor U2474 (N_2474,N_2246,N_2349);
or U2475 (N_2475,N_2223,N_2290);
or U2476 (N_2476,N_2278,N_2227);
xor U2477 (N_2477,N_2302,N_2363);
nor U2478 (N_2478,N_2285,N_2389);
or U2479 (N_2479,N_2333,N_2342);
or U2480 (N_2480,N_2375,N_2322);
or U2481 (N_2481,N_2275,N_2209);
and U2482 (N_2482,N_2327,N_2203);
xor U2483 (N_2483,N_2336,N_2329);
nor U2484 (N_2484,N_2379,N_2386);
xnor U2485 (N_2485,N_2298,N_2343);
nand U2486 (N_2486,N_2279,N_2356);
xnor U2487 (N_2487,N_2330,N_2371);
nor U2488 (N_2488,N_2396,N_2240);
xnor U2489 (N_2489,N_2354,N_2248);
xor U2490 (N_2490,N_2361,N_2204);
and U2491 (N_2491,N_2247,N_2226);
or U2492 (N_2492,N_2249,N_2348);
nor U2493 (N_2493,N_2234,N_2208);
xnor U2494 (N_2494,N_2241,N_2282);
xnor U2495 (N_2495,N_2300,N_2310);
or U2496 (N_2496,N_2260,N_2317);
and U2497 (N_2497,N_2294,N_2341);
or U2498 (N_2498,N_2256,N_2304);
xor U2499 (N_2499,N_2274,N_2382);
nand U2500 (N_2500,N_2308,N_2294);
nor U2501 (N_2501,N_2241,N_2253);
nor U2502 (N_2502,N_2312,N_2378);
nand U2503 (N_2503,N_2261,N_2307);
and U2504 (N_2504,N_2367,N_2236);
xnor U2505 (N_2505,N_2369,N_2380);
xnor U2506 (N_2506,N_2265,N_2244);
nand U2507 (N_2507,N_2301,N_2308);
xor U2508 (N_2508,N_2287,N_2248);
xor U2509 (N_2509,N_2265,N_2264);
or U2510 (N_2510,N_2366,N_2273);
and U2511 (N_2511,N_2275,N_2372);
nor U2512 (N_2512,N_2297,N_2394);
and U2513 (N_2513,N_2222,N_2373);
and U2514 (N_2514,N_2363,N_2204);
nor U2515 (N_2515,N_2239,N_2332);
or U2516 (N_2516,N_2209,N_2280);
nor U2517 (N_2517,N_2272,N_2238);
xnor U2518 (N_2518,N_2240,N_2301);
or U2519 (N_2519,N_2248,N_2276);
or U2520 (N_2520,N_2293,N_2354);
nor U2521 (N_2521,N_2237,N_2308);
or U2522 (N_2522,N_2303,N_2203);
xnor U2523 (N_2523,N_2365,N_2260);
nand U2524 (N_2524,N_2283,N_2207);
nand U2525 (N_2525,N_2264,N_2387);
nor U2526 (N_2526,N_2248,N_2289);
nand U2527 (N_2527,N_2231,N_2204);
or U2528 (N_2528,N_2203,N_2225);
or U2529 (N_2529,N_2378,N_2216);
or U2530 (N_2530,N_2295,N_2271);
and U2531 (N_2531,N_2234,N_2233);
or U2532 (N_2532,N_2366,N_2307);
or U2533 (N_2533,N_2370,N_2360);
and U2534 (N_2534,N_2392,N_2390);
nand U2535 (N_2535,N_2221,N_2275);
xor U2536 (N_2536,N_2224,N_2332);
nor U2537 (N_2537,N_2252,N_2317);
and U2538 (N_2538,N_2215,N_2355);
or U2539 (N_2539,N_2216,N_2261);
xnor U2540 (N_2540,N_2237,N_2229);
nor U2541 (N_2541,N_2380,N_2313);
nand U2542 (N_2542,N_2320,N_2227);
xnor U2543 (N_2543,N_2231,N_2379);
nor U2544 (N_2544,N_2368,N_2321);
xnor U2545 (N_2545,N_2212,N_2221);
xnor U2546 (N_2546,N_2232,N_2202);
xnor U2547 (N_2547,N_2203,N_2312);
xnor U2548 (N_2548,N_2280,N_2250);
xor U2549 (N_2549,N_2273,N_2288);
and U2550 (N_2550,N_2344,N_2351);
xor U2551 (N_2551,N_2361,N_2205);
xor U2552 (N_2552,N_2373,N_2377);
nor U2553 (N_2553,N_2289,N_2261);
nand U2554 (N_2554,N_2296,N_2253);
xor U2555 (N_2555,N_2293,N_2355);
or U2556 (N_2556,N_2299,N_2287);
and U2557 (N_2557,N_2253,N_2260);
nor U2558 (N_2558,N_2228,N_2309);
and U2559 (N_2559,N_2299,N_2246);
xor U2560 (N_2560,N_2335,N_2297);
xnor U2561 (N_2561,N_2292,N_2362);
xnor U2562 (N_2562,N_2318,N_2208);
nor U2563 (N_2563,N_2244,N_2222);
and U2564 (N_2564,N_2224,N_2295);
nand U2565 (N_2565,N_2217,N_2214);
or U2566 (N_2566,N_2275,N_2288);
and U2567 (N_2567,N_2286,N_2364);
and U2568 (N_2568,N_2261,N_2280);
xnor U2569 (N_2569,N_2332,N_2381);
or U2570 (N_2570,N_2296,N_2367);
nand U2571 (N_2571,N_2386,N_2200);
and U2572 (N_2572,N_2342,N_2247);
or U2573 (N_2573,N_2247,N_2321);
or U2574 (N_2574,N_2267,N_2278);
xor U2575 (N_2575,N_2336,N_2260);
xnor U2576 (N_2576,N_2354,N_2386);
or U2577 (N_2577,N_2311,N_2327);
or U2578 (N_2578,N_2370,N_2230);
or U2579 (N_2579,N_2237,N_2214);
nor U2580 (N_2580,N_2294,N_2366);
and U2581 (N_2581,N_2244,N_2218);
nand U2582 (N_2582,N_2263,N_2383);
xor U2583 (N_2583,N_2231,N_2221);
xnor U2584 (N_2584,N_2221,N_2373);
nand U2585 (N_2585,N_2219,N_2348);
and U2586 (N_2586,N_2319,N_2361);
and U2587 (N_2587,N_2223,N_2382);
and U2588 (N_2588,N_2286,N_2314);
nor U2589 (N_2589,N_2239,N_2371);
nor U2590 (N_2590,N_2331,N_2277);
xor U2591 (N_2591,N_2378,N_2241);
nand U2592 (N_2592,N_2214,N_2241);
and U2593 (N_2593,N_2342,N_2239);
nand U2594 (N_2594,N_2312,N_2347);
and U2595 (N_2595,N_2296,N_2256);
nor U2596 (N_2596,N_2316,N_2384);
xor U2597 (N_2597,N_2395,N_2233);
or U2598 (N_2598,N_2289,N_2377);
xnor U2599 (N_2599,N_2252,N_2320);
and U2600 (N_2600,N_2405,N_2466);
nor U2601 (N_2601,N_2421,N_2409);
or U2602 (N_2602,N_2563,N_2444);
or U2603 (N_2603,N_2413,N_2406);
and U2604 (N_2604,N_2401,N_2502);
xor U2605 (N_2605,N_2496,N_2418);
nand U2606 (N_2606,N_2528,N_2522);
nand U2607 (N_2607,N_2426,N_2585);
nor U2608 (N_2608,N_2550,N_2488);
nor U2609 (N_2609,N_2472,N_2524);
nor U2610 (N_2610,N_2478,N_2476);
nand U2611 (N_2611,N_2440,N_2541);
xnor U2612 (N_2612,N_2419,N_2568);
nor U2613 (N_2613,N_2464,N_2507);
nand U2614 (N_2614,N_2567,N_2412);
and U2615 (N_2615,N_2420,N_2498);
xor U2616 (N_2616,N_2554,N_2495);
and U2617 (N_2617,N_2519,N_2523);
nor U2618 (N_2618,N_2455,N_2587);
xor U2619 (N_2619,N_2576,N_2453);
nor U2620 (N_2620,N_2536,N_2530);
or U2621 (N_2621,N_2400,N_2517);
and U2622 (N_2622,N_2415,N_2410);
nand U2623 (N_2623,N_2459,N_2577);
xor U2624 (N_2624,N_2434,N_2544);
nand U2625 (N_2625,N_2474,N_2408);
nor U2626 (N_2626,N_2407,N_2532);
or U2627 (N_2627,N_2486,N_2548);
nor U2628 (N_2628,N_2553,N_2423);
and U2629 (N_2629,N_2460,N_2580);
and U2630 (N_2630,N_2551,N_2583);
nor U2631 (N_2631,N_2468,N_2525);
or U2632 (N_2632,N_2512,N_2475);
nor U2633 (N_2633,N_2473,N_2581);
or U2634 (N_2634,N_2471,N_2579);
nor U2635 (N_2635,N_2490,N_2540);
nor U2636 (N_2636,N_2492,N_2594);
nand U2637 (N_2637,N_2574,N_2456);
or U2638 (N_2638,N_2566,N_2561);
or U2639 (N_2639,N_2484,N_2596);
and U2640 (N_2640,N_2573,N_2485);
nor U2641 (N_2641,N_2597,N_2510);
or U2642 (N_2642,N_2452,N_2547);
xnor U2643 (N_2643,N_2569,N_2531);
and U2644 (N_2644,N_2454,N_2416);
or U2645 (N_2645,N_2521,N_2427);
nor U2646 (N_2646,N_2586,N_2590);
nor U2647 (N_2647,N_2450,N_2527);
nor U2648 (N_2648,N_2487,N_2529);
xnor U2649 (N_2649,N_2584,N_2433);
nand U2650 (N_2650,N_2598,N_2489);
xor U2651 (N_2651,N_2564,N_2500);
and U2652 (N_2652,N_2439,N_2477);
nand U2653 (N_2653,N_2565,N_2430);
nand U2654 (N_2654,N_2501,N_2417);
and U2655 (N_2655,N_2447,N_2402);
or U2656 (N_2656,N_2504,N_2497);
nor U2657 (N_2657,N_2494,N_2446);
and U2658 (N_2658,N_2438,N_2578);
nor U2659 (N_2659,N_2589,N_2506);
nor U2660 (N_2660,N_2463,N_2509);
nor U2661 (N_2661,N_2479,N_2559);
nor U2662 (N_2662,N_2537,N_2461);
xnor U2663 (N_2663,N_2552,N_2514);
nand U2664 (N_2664,N_2428,N_2595);
or U2665 (N_2665,N_2425,N_2445);
nor U2666 (N_2666,N_2414,N_2543);
nand U2667 (N_2667,N_2424,N_2526);
and U2668 (N_2668,N_2555,N_2441);
or U2669 (N_2669,N_2535,N_2451);
nor U2670 (N_2670,N_2469,N_2470);
xnor U2671 (N_2671,N_2505,N_2481);
xor U2672 (N_2672,N_2513,N_2499);
or U2673 (N_2673,N_2575,N_2465);
or U2674 (N_2674,N_2549,N_2582);
and U2675 (N_2675,N_2533,N_2449);
and U2676 (N_2676,N_2546,N_2467);
nor U2677 (N_2677,N_2592,N_2593);
and U2678 (N_2678,N_2491,N_2435);
nand U2679 (N_2679,N_2457,N_2483);
xnor U2680 (N_2680,N_2480,N_2437);
xor U2681 (N_2681,N_2557,N_2591);
xnor U2682 (N_2682,N_2508,N_2482);
and U2683 (N_2683,N_2429,N_2545);
nand U2684 (N_2684,N_2520,N_2516);
xnor U2685 (N_2685,N_2572,N_2558);
nand U2686 (N_2686,N_2432,N_2458);
nand U2687 (N_2687,N_2570,N_2443);
nand U2688 (N_2688,N_2404,N_2493);
nand U2689 (N_2689,N_2462,N_2448);
or U2690 (N_2690,N_2422,N_2556);
and U2691 (N_2691,N_2518,N_2542);
xor U2692 (N_2692,N_2562,N_2411);
xnor U2693 (N_2693,N_2442,N_2436);
nor U2694 (N_2694,N_2599,N_2538);
or U2695 (N_2695,N_2588,N_2560);
or U2696 (N_2696,N_2515,N_2511);
and U2697 (N_2697,N_2431,N_2403);
nor U2698 (N_2698,N_2534,N_2503);
nor U2699 (N_2699,N_2539,N_2571);
nand U2700 (N_2700,N_2598,N_2491);
or U2701 (N_2701,N_2506,N_2565);
and U2702 (N_2702,N_2552,N_2535);
or U2703 (N_2703,N_2406,N_2456);
xnor U2704 (N_2704,N_2547,N_2579);
xnor U2705 (N_2705,N_2554,N_2497);
or U2706 (N_2706,N_2415,N_2483);
and U2707 (N_2707,N_2474,N_2443);
and U2708 (N_2708,N_2548,N_2494);
nand U2709 (N_2709,N_2470,N_2416);
nor U2710 (N_2710,N_2454,N_2545);
and U2711 (N_2711,N_2543,N_2437);
xnor U2712 (N_2712,N_2530,N_2404);
nand U2713 (N_2713,N_2530,N_2417);
or U2714 (N_2714,N_2501,N_2484);
nor U2715 (N_2715,N_2540,N_2420);
xnor U2716 (N_2716,N_2485,N_2410);
or U2717 (N_2717,N_2580,N_2547);
and U2718 (N_2718,N_2449,N_2499);
or U2719 (N_2719,N_2589,N_2544);
xnor U2720 (N_2720,N_2570,N_2522);
xor U2721 (N_2721,N_2560,N_2477);
nor U2722 (N_2722,N_2477,N_2590);
and U2723 (N_2723,N_2550,N_2400);
nand U2724 (N_2724,N_2547,N_2482);
and U2725 (N_2725,N_2408,N_2510);
xor U2726 (N_2726,N_2533,N_2504);
nand U2727 (N_2727,N_2586,N_2462);
and U2728 (N_2728,N_2583,N_2528);
nand U2729 (N_2729,N_2574,N_2489);
xor U2730 (N_2730,N_2477,N_2531);
nor U2731 (N_2731,N_2580,N_2590);
nor U2732 (N_2732,N_2592,N_2476);
xnor U2733 (N_2733,N_2483,N_2458);
xor U2734 (N_2734,N_2430,N_2484);
xor U2735 (N_2735,N_2549,N_2483);
nor U2736 (N_2736,N_2466,N_2497);
or U2737 (N_2737,N_2477,N_2540);
nand U2738 (N_2738,N_2546,N_2569);
xnor U2739 (N_2739,N_2465,N_2454);
nand U2740 (N_2740,N_2576,N_2572);
nor U2741 (N_2741,N_2562,N_2465);
or U2742 (N_2742,N_2569,N_2520);
and U2743 (N_2743,N_2427,N_2522);
nand U2744 (N_2744,N_2528,N_2475);
xor U2745 (N_2745,N_2442,N_2421);
nor U2746 (N_2746,N_2589,N_2421);
or U2747 (N_2747,N_2570,N_2450);
or U2748 (N_2748,N_2431,N_2456);
and U2749 (N_2749,N_2554,N_2494);
and U2750 (N_2750,N_2436,N_2576);
nand U2751 (N_2751,N_2555,N_2508);
xor U2752 (N_2752,N_2589,N_2548);
xnor U2753 (N_2753,N_2433,N_2411);
xnor U2754 (N_2754,N_2410,N_2447);
or U2755 (N_2755,N_2408,N_2460);
and U2756 (N_2756,N_2405,N_2593);
xnor U2757 (N_2757,N_2595,N_2405);
and U2758 (N_2758,N_2511,N_2514);
or U2759 (N_2759,N_2458,N_2434);
or U2760 (N_2760,N_2522,N_2578);
xor U2761 (N_2761,N_2472,N_2497);
and U2762 (N_2762,N_2406,N_2513);
xnor U2763 (N_2763,N_2566,N_2492);
or U2764 (N_2764,N_2407,N_2499);
xnor U2765 (N_2765,N_2458,N_2569);
xnor U2766 (N_2766,N_2492,N_2433);
and U2767 (N_2767,N_2496,N_2461);
or U2768 (N_2768,N_2435,N_2486);
and U2769 (N_2769,N_2492,N_2508);
xor U2770 (N_2770,N_2532,N_2449);
nor U2771 (N_2771,N_2560,N_2567);
xor U2772 (N_2772,N_2400,N_2450);
nor U2773 (N_2773,N_2497,N_2450);
and U2774 (N_2774,N_2521,N_2558);
xor U2775 (N_2775,N_2407,N_2436);
nand U2776 (N_2776,N_2513,N_2485);
and U2777 (N_2777,N_2507,N_2482);
nand U2778 (N_2778,N_2453,N_2455);
xor U2779 (N_2779,N_2452,N_2469);
nand U2780 (N_2780,N_2432,N_2487);
and U2781 (N_2781,N_2440,N_2528);
nand U2782 (N_2782,N_2471,N_2415);
and U2783 (N_2783,N_2571,N_2481);
nand U2784 (N_2784,N_2493,N_2489);
and U2785 (N_2785,N_2460,N_2532);
and U2786 (N_2786,N_2428,N_2518);
and U2787 (N_2787,N_2509,N_2514);
nor U2788 (N_2788,N_2414,N_2405);
and U2789 (N_2789,N_2431,N_2556);
and U2790 (N_2790,N_2481,N_2409);
nor U2791 (N_2791,N_2490,N_2419);
or U2792 (N_2792,N_2467,N_2444);
nand U2793 (N_2793,N_2415,N_2585);
nand U2794 (N_2794,N_2492,N_2543);
nor U2795 (N_2795,N_2521,N_2414);
xor U2796 (N_2796,N_2559,N_2464);
or U2797 (N_2797,N_2458,N_2566);
or U2798 (N_2798,N_2503,N_2489);
or U2799 (N_2799,N_2562,N_2528);
or U2800 (N_2800,N_2677,N_2789);
nand U2801 (N_2801,N_2791,N_2771);
xnor U2802 (N_2802,N_2607,N_2724);
nor U2803 (N_2803,N_2657,N_2679);
xor U2804 (N_2804,N_2788,N_2762);
and U2805 (N_2805,N_2623,N_2611);
nand U2806 (N_2806,N_2695,N_2617);
or U2807 (N_2807,N_2661,N_2625);
xnor U2808 (N_2808,N_2738,N_2665);
nor U2809 (N_2809,N_2663,N_2610);
or U2810 (N_2810,N_2733,N_2747);
and U2811 (N_2811,N_2720,N_2683);
nor U2812 (N_2812,N_2775,N_2659);
and U2813 (N_2813,N_2674,N_2698);
xnor U2814 (N_2814,N_2614,N_2774);
xor U2815 (N_2815,N_2647,N_2780);
nor U2816 (N_2816,N_2670,N_2669);
xnor U2817 (N_2817,N_2776,N_2787);
nor U2818 (N_2818,N_2620,N_2742);
nand U2819 (N_2819,N_2729,N_2730);
or U2820 (N_2820,N_2628,N_2778);
nand U2821 (N_2821,N_2668,N_2633);
nand U2822 (N_2822,N_2785,N_2728);
xnor U2823 (N_2823,N_2767,N_2651);
or U2824 (N_2824,N_2686,N_2681);
or U2825 (N_2825,N_2601,N_2758);
and U2826 (N_2826,N_2676,N_2717);
and U2827 (N_2827,N_2682,N_2640);
nor U2828 (N_2828,N_2786,N_2777);
and U2829 (N_2829,N_2632,N_2693);
nor U2830 (N_2830,N_2662,N_2783);
and U2831 (N_2831,N_2752,N_2678);
nand U2832 (N_2832,N_2710,N_2731);
xor U2833 (N_2833,N_2772,N_2675);
nand U2834 (N_2834,N_2630,N_2779);
nand U2835 (N_2835,N_2646,N_2692);
and U2836 (N_2836,N_2604,N_2644);
nor U2837 (N_2837,N_2672,N_2653);
xnor U2838 (N_2838,N_2746,N_2721);
and U2839 (N_2839,N_2613,N_2685);
xnor U2840 (N_2840,N_2616,N_2741);
xnor U2841 (N_2841,N_2643,N_2799);
and U2842 (N_2842,N_2658,N_2627);
and U2843 (N_2843,N_2696,N_2726);
or U2844 (N_2844,N_2709,N_2744);
nand U2845 (N_2845,N_2602,N_2773);
xor U2846 (N_2846,N_2745,N_2603);
nor U2847 (N_2847,N_2629,N_2794);
nand U2848 (N_2848,N_2751,N_2756);
nor U2849 (N_2849,N_2792,N_2708);
nand U2850 (N_2850,N_2739,N_2723);
or U2851 (N_2851,N_2722,N_2700);
or U2852 (N_2852,N_2687,N_2734);
nand U2853 (N_2853,N_2635,N_2714);
and U2854 (N_2854,N_2768,N_2624);
xnor U2855 (N_2855,N_2621,N_2725);
nand U2856 (N_2856,N_2688,N_2732);
xnor U2857 (N_2857,N_2740,N_2600);
and U2858 (N_2858,N_2684,N_2618);
nand U2859 (N_2859,N_2605,N_2790);
xnor U2860 (N_2860,N_2638,N_2769);
nor U2861 (N_2861,N_2671,N_2718);
nand U2862 (N_2862,N_2689,N_2703);
and U2863 (N_2863,N_2736,N_2694);
or U2864 (N_2864,N_2760,N_2699);
and U2865 (N_2865,N_2716,N_2609);
nor U2866 (N_2866,N_2754,N_2798);
or U2867 (N_2867,N_2743,N_2619);
xnor U2868 (N_2868,N_2770,N_2704);
and U2869 (N_2869,N_2648,N_2713);
or U2870 (N_2870,N_2702,N_2645);
nor U2871 (N_2871,N_2622,N_2764);
and U2872 (N_2872,N_2680,N_2707);
xnor U2873 (N_2873,N_2765,N_2691);
nor U2874 (N_2874,N_2711,N_2757);
nor U2875 (N_2875,N_2615,N_2705);
and U2876 (N_2876,N_2750,N_2650);
nor U2877 (N_2877,N_2795,N_2782);
and U2878 (N_2878,N_2636,N_2749);
or U2879 (N_2879,N_2690,N_2660);
and U2880 (N_2880,N_2715,N_2639);
nor U2881 (N_2881,N_2781,N_2641);
and U2882 (N_2882,N_2656,N_2761);
xor U2883 (N_2883,N_2766,N_2637);
xnor U2884 (N_2884,N_2666,N_2608);
or U2885 (N_2885,N_2634,N_2748);
or U2886 (N_2886,N_2649,N_2753);
nand U2887 (N_2887,N_2664,N_2654);
nor U2888 (N_2888,N_2626,N_2631);
and U2889 (N_2889,N_2793,N_2667);
xor U2890 (N_2890,N_2612,N_2652);
nand U2891 (N_2891,N_2642,N_2735);
nand U2892 (N_2892,N_2759,N_2712);
nand U2893 (N_2893,N_2697,N_2606);
nor U2894 (N_2894,N_2797,N_2755);
and U2895 (N_2895,N_2737,N_2673);
xnor U2896 (N_2896,N_2784,N_2763);
or U2897 (N_2897,N_2719,N_2655);
nand U2898 (N_2898,N_2796,N_2727);
xor U2899 (N_2899,N_2701,N_2706);
xor U2900 (N_2900,N_2602,N_2640);
nand U2901 (N_2901,N_2647,N_2698);
xnor U2902 (N_2902,N_2717,N_2746);
xor U2903 (N_2903,N_2784,N_2726);
xor U2904 (N_2904,N_2625,N_2721);
and U2905 (N_2905,N_2617,N_2774);
nand U2906 (N_2906,N_2655,N_2687);
nor U2907 (N_2907,N_2667,N_2723);
xnor U2908 (N_2908,N_2784,N_2630);
and U2909 (N_2909,N_2786,N_2696);
xor U2910 (N_2910,N_2637,N_2689);
nor U2911 (N_2911,N_2751,N_2604);
nor U2912 (N_2912,N_2713,N_2716);
and U2913 (N_2913,N_2685,N_2645);
nor U2914 (N_2914,N_2732,N_2731);
or U2915 (N_2915,N_2787,N_2687);
or U2916 (N_2916,N_2785,N_2683);
nor U2917 (N_2917,N_2701,N_2638);
nand U2918 (N_2918,N_2775,N_2663);
xnor U2919 (N_2919,N_2657,N_2665);
nor U2920 (N_2920,N_2617,N_2625);
nand U2921 (N_2921,N_2608,N_2652);
nor U2922 (N_2922,N_2758,N_2740);
or U2923 (N_2923,N_2613,N_2668);
and U2924 (N_2924,N_2766,N_2703);
and U2925 (N_2925,N_2662,N_2698);
nor U2926 (N_2926,N_2792,N_2752);
and U2927 (N_2927,N_2699,N_2652);
and U2928 (N_2928,N_2632,N_2659);
and U2929 (N_2929,N_2625,N_2674);
and U2930 (N_2930,N_2719,N_2667);
and U2931 (N_2931,N_2759,N_2609);
or U2932 (N_2932,N_2741,N_2651);
xnor U2933 (N_2933,N_2600,N_2635);
nand U2934 (N_2934,N_2629,N_2736);
or U2935 (N_2935,N_2651,N_2712);
xor U2936 (N_2936,N_2612,N_2763);
and U2937 (N_2937,N_2786,N_2725);
xnor U2938 (N_2938,N_2682,N_2784);
nor U2939 (N_2939,N_2662,N_2771);
and U2940 (N_2940,N_2733,N_2639);
nand U2941 (N_2941,N_2618,N_2729);
xnor U2942 (N_2942,N_2741,N_2689);
nand U2943 (N_2943,N_2644,N_2694);
nand U2944 (N_2944,N_2702,N_2680);
or U2945 (N_2945,N_2618,N_2631);
or U2946 (N_2946,N_2745,N_2765);
and U2947 (N_2947,N_2693,N_2717);
and U2948 (N_2948,N_2675,N_2681);
or U2949 (N_2949,N_2775,N_2722);
nor U2950 (N_2950,N_2622,N_2761);
nand U2951 (N_2951,N_2661,N_2680);
xnor U2952 (N_2952,N_2785,N_2664);
xnor U2953 (N_2953,N_2768,N_2655);
or U2954 (N_2954,N_2718,N_2728);
and U2955 (N_2955,N_2656,N_2643);
nor U2956 (N_2956,N_2656,N_2630);
or U2957 (N_2957,N_2685,N_2757);
nor U2958 (N_2958,N_2695,N_2618);
or U2959 (N_2959,N_2616,N_2690);
xor U2960 (N_2960,N_2673,N_2649);
or U2961 (N_2961,N_2688,N_2726);
or U2962 (N_2962,N_2770,N_2674);
or U2963 (N_2963,N_2743,N_2721);
xor U2964 (N_2964,N_2730,N_2761);
and U2965 (N_2965,N_2713,N_2661);
or U2966 (N_2966,N_2666,N_2658);
and U2967 (N_2967,N_2632,N_2678);
or U2968 (N_2968,N_2665,N_2659);
nand U2969 (N_2969,N_2608,N_2636);
or U2970 (N_2970,N_2629,N_2642);
and U2971 (N_2971,N_2618,N_2619);
xor U2972 (N_2972,N_2719,N_2622);
nand U2973 (N_2973,N_2765,N_2768);
xnor U2974 (N_2974,N_2649,N_2708);
and U2975 (N_2975,N_2723,N_2653);
nand U2976 (N_2976,N_2791,N_2617);
and U2977 (N_2977,N_2671,N_2666);
nand U2978 (N_2978,N_2618,N_2687);
xor U2979 (N_2979,N_2741,N_2657);
nor U2980 (N_2980,N_2782,N_2691);
nor U2981 (N_2981,N_2639,N_2727);
and U2982 (N_2982,N_2774,N_2751);
xnor U2983 (N_2983,N_2776,N_2689);
nand U2984 (N_2984,N_2642,N_2790);
nor U2985 (N_2985,N_2739,N_2657);
or U2986 (N_2986,N_2748,N_2675);
and U2987 (N_2987,N_2602,N_2729);
xor U2988 (N_2988,N_2673,N_2622);
nor U2989 (N_2989,N_2625,N_2623);
nor U2990 (N_2990,N_2719,N_2787);
nand U2991 (N_2991,N_2685,N_2618);
or U2992 (N_2992,N_2620,N_2627);
and U2993 (N_2993,N_2675,N_2625);
or U2994 (N_2994,N_2637,N_2785);
nand U2995 (N_2995,N_2748,N_2693);
nand U2996 (N_2996,N_2792,N_2694);
xor U2997 (N_2997,N_2745,N_2776);
nor U2998 (N_2998,N_2640,N_2633);
nand U2999 (N_2999,N_2635,N_2606);
and U3000 (N_3000,N_2861,N_2810);
xor U3001 (N_3001,N_2899,N_2996);
nand U3002 (N_3002,N_2978,N_2868);
nor U3003 (N_3003,N_2869,N_2831);
or U3004 (N_3004,N_2801,N_2816);
or U3005 (N_3005,N_2938,N_2917);
xnor U3006 (N_3006,N_2960,N_2814);
or U3007 (N_3007,N_2942,N_2968);
and U3008 (N_3008,N_2975,N_2981);
nand U3009 (N_3009,N_2955,N_2992);
nor U3010 (N_3010,N_2957,N_2807);
and U3011 (N_3011,N_2943,N_2826);
or U3012 (N_3012,N_2974,N_2930);
nand U3013 (N_3013,N_2908,N_2856);
and U3014 (N_3014,N_2809,N_2895);
nand U3015 (N_3015,N_2844,N_2841);
or U3016 (N_3016,N_2838,N_2980);
xnor U3017 (N_3017,N_2886,N_2910);
xnor U3018 (N_3018,N_2846,N_2945);
or U3019 (N_3019,N_2865,N_2973);
nor U3020 (N_3020,N_2825,N_2836);
or U3021 (N_3021,N_2934,N_2994);
and U3022 (N_3022,N_2839,N_2958);
xor U3023 (N_3023,N_2843,N_2859);
and U3024 (N_3024,N_2935,N_2920);
nor U3025 (N_3025,N_2890,N_2904);
xor U3026 (N_3026,N_2997,N_2876);
nand U3027 (N_3027,N_2933,N_2857);
nand U3028 (N_3028,N_2882,N_2830);
and U3029 (N_3029,N_2971,N_2834);
and U3030 (N_3030,N_2940,N_2840);
or U3031 (N_3031,N_2907,N_2903);
nor U3032 (N_3032,N_2905,N_2873);
and U3033 (N_3033,N_2811,N_2969);
or U3034 (N_3034,N_2879,N_2970);
and U3035 (N_3035,N_2884,N_2953);
or U3036 (N_3036,N_2914,N_2983);
and U3037 (N_3037,N_2972,N_2928);
or U3038 (N_3038,N_2999,N_2924);
and U3039 (N_3039,N_2932,N_2912);
nor U3040 (N_3040,N_2991,N_2835);
and U3041 (N_3041,N_2875,N_2894);
or U3042 (N_3042,N_2906,N_2897);
and U3043 (N_3043,N_2853,N_2995);
nor U3044 (N_3044,N_2850,N_2989);
nor U3045 (N_3045,N_2842,N_2847);
xnor U3046 (N_3046,N_2963,N_2818);
and U3047 (N_3047,N_2959,N_2946);
nand U3048 (N_3048,N_2845,N_2949);
nand U3049 (N_3049,N_2936,N_2979);
nor U3050 (N_3050,N_2874,N_2966);
or U3051 (N_3051,N_2866,N_2800);
nor U3052 (N_3052,N_2948,N_2944);
or U3053 (N_3053,N_2923,N_2804);
xnor U3054 (N_3054,N_2821,N_2820);
xor U3055 (N_3055,N_2998,N_2878);
and U3056 (N_3056,N_2880,N_2956);
nor U3057 (N_3057,N_2922,N_2954);
nor U3058 (N_3058,N_2967,N_2976);
or U3059 (N_3059,N_2911,N_2915);
nor U3060 (N_3060,N_2984,N_2871);
nor U3061 (N_3061,N_2916,N_2863);
nand U3062 (N_3062,N_2855,N_2817);
and U3063 (N_3063,N_2877,N_2828);
and U3064 (N_3064,N_2990,N_2921);
nor U3065 (N_3065,N_2862,N_2829);
or U3066 (N_3066,N_2867,N_2926);
and U3067 (N_3067,N_2803,N_2872);
nand U3068 (N_3068,N_2909,N_2813);
nor U3069 (N_3069,N_2819,N_2883);
nor U3070 (N_3070,N_2888,N_2827);
xnor U3071 (N_3071,N_2993,N_2927);
and U3072 (N_3072,N_2902,N_2852);
and U3073 (N_3073,N_2977,N_2964);
and U3074 (N_3074,N_2824,N_2858);
or U3075 (N_3075,N_2947,N_2851);
xnor U3076 (N_3076,N_2812,N_2848);
nor U3077 (N_3077,N_2985,N_2986);
xnor U3078 (N_3078,N_2987,N_2889);
nand U3079 (N_3079,N_2887,N_2941);
xor U3080 (N_3080,N_2832,N_2962);
nand U3081 (N_3081,N_2896,N_2925);
and U3082 (N_3082,N_2881,N_2952);
and U3083 (N_3083,N_2901,N_2891);
nand U3084 (N_3084,N_2854,N_2892);
and U3085 (N_3085,N_2937,N_2805);
nand U3086 (N_3086,N_2931,N_2885);
and U3087 (N_3087,N_2893,N_2929);
xnor U3088 (N_3088,N_2919,N_2833);
or U3089 (N_3089,N_2982,N_2950);
or U3090 (N_3090,N_2864,N_2837);
nor U3091 (N_3091,N_2913,N_2806);
xnor U3092 (N_3092,N_2900,N_2802);
nand U3093 (N_3093,N_2939,N_2860);
xor U3094 (N_3094,N_2918,N_2822);
and U3095 (N_3095,N_2823,N_2988);
xor U3096 (N_3096,N_2815,N_2961);
xnor U3097 (N_3097,N_2849,N_2965);
nor U3098 (N_3098,N_2951,N_2808);
nand U3099 (N_3099,N_2898,N_2870);
xor U3100 (N_3100,N_2916,N_2947);
nor U3101 (N_3101,N_2881,N_2813);
nand U3102 (N_3102,N_2935,N_2805);
and U3103 (N_3103,N_2883,N_2886);
and U3104 (N_3104,N_2870,N_2969);
or U3105 (N_3105,N_2835,N_2866);
or U3106 (N_3106,N_2935,N_2869);
and U3107 (N_3107,N_2820,N_2846);
and U3108 (N_3108,N_2943,N_2895);
or U3109 (N_3109,N_2840,N_2813);
nand U3110 (N_3110,N_2852,N_2875);
and U3111 (N_3111,N_2992,N_2949);
or U3112 (N_3112,N_2986,N_2859);
nand U3113 (N_3113,N_2810,N_2962);
and U3114 (N_3114,N_2911,N_2879);
and U3115 (N_3115,N_2969,N_2994);
and U3116 (N_3116,N_2876,N_2808);
or U3117 (N_3117,N_2888,N_2964);
nand U3118 (N_3118,N_2852,N_2994);
nor U3119 (N_3119,N_2953,N_2864);
and U3120 (N_3120,N_2864,N_2975);
and U3121 (N_3121,N_2935,N_2913);
and U3122 (N_3122,N_2988,N_2989);
nor U3123 (N_3123,N_2926,N_2958);
or U3124 (N_3124,N_2976,N_2867);
and U3125 (N_3125,N_2838,N_2881);
nand U3126 (N_3126,N_2968,N_2950);
nand U3127 (N_3127,N_2803,N_2822);
xnor U3128 (N_3128,N_2854,N_2822);
and U3129 (N_3129,N_2809,N_2896);
xor U3130 (N_3130,N_2891,N_2957);
and U3131 (N_3131,N_2966,N_2869);
nand U3132 (N_3132,N_2896,N_2914);
xnor U3133 (N_3133,N_2876,N_2987);
xor U3134 (N_3134,N_2847,N_2907);
nand U3135 (N_3135,N_2937,N_2918);
or U3136 (N_3136,N_2944,N_2913);
nand U3137 (N_3137,N_2914,N_2927);
or U3138 (N_3138,N_2862,N_2974);
nor U3139 (N_3139,N_2992,N_2818);
nor U3140 (N_3140,N_2978,N_2835);
nor U3141 (N_3141,N_2800,N_2828);
nor U3142 (N_3142,N_2918,N_2910);
xor U3143 (N_3143,N_2849,N_2962);
nor U3144 (N_3144,N_2951,N_2823);
nand U3145 (N_3145,N_2899,N_2813);
nand U3146 (N_3146,N_2893,N_2821);
and U3147 (N_3147,N_2826,N_2824);
nor U3148 (N_3148,N_2886,N_2925);
nand U3149 (N_3149,N_2932,N_2817);
or U3150 (N_3150,N_2988,N_2844);
xor U3151 (N_3151,N_2948,N_2942);
and U3152 (N_3152,N_2832,N_2988);
and U3153 (N_3153,N_2897,N_2959);
or U3154 (N_3154,N_2861,N_2947);
or U3155 (N_3155,N_2825,N_2921);
nor U3156 (N_3156,N_2821,N_2961);
nor U3157 (N_3157,N_2979,N_2851);
nand U3158 (N_3158,N_2818,N_2803);
nand U3159 (N_3159,N_2816,N_2980);
nor U3160 (N_3160,N_2954,N_2897);
and U3161 (N_3161,N_2826,N_2896);
and U3162 (N_3162,N_2884,N_2890);
nor U3163 (N_3163,N_2979,N_2872);
and U3164 (N_3164,N_2980,N_2865);
and U3165 (N_3165,N_2905,N_2937);
or U3166 (N_3166,N_2829,N_2958);
nor U3167 (N_3167,N_2985,N_2947);
or U3168 (N_3168,N_2962,N_2879);
nor U3169 (N_3169,N_2886,N_2941);
nand U3170 (N_3170,N_2996,N_2869);
and U3171 (N_3171,N_2942,N_2892);
nor U3172 (N_3172,N_2972,N_2934);
nor U3173 (N_3173,N_2829,N_2973);
and U3174 (N_3174,N_2954,N_2943);
xor U3175 (N_3175,N_2958,N_2864);
nor U3176 (N_3176,N_2990,N_2901);
xor U3177 (N_3177,N_2944,N_2977);
nor U3178 (N_3178,N_2862,N_2910);
or U3179 (N_3179,N_2850,N_2841);
or U3180 (N_3180,N_2823,N_2961);
nand U3181 (N_3181,N_2935,N_2934);
xnor U3182 (N_3182,N_2816,N_2900);
or U3183 (N_3183,N_2803,N_2905);
or U3184 (N_3184,N_2883,N_2888);
nand U3185 (N_3185,N_2876,N_2880);
nor U3186 (N_3186,N_2961,N_2982);
nand U3187 (N_3187,N_2877,N_2963);
nor U3188 (N_3188,N_2937,N_2887);
nor U3189 (N_3189,N_2866,N_2985);
nor U3190 (N_3190,N_2856,N_2967);
nor U3191 (N_3191,N_2926,N_2861);
and U3192 (N_3192,N_2969,N_2822);
and U3193 (N_3193,N_2992,N_2896);
nand U3194 (N_3194,N_2871,N_2870);
xnor U3195 (N_3195,N_2877,N_2894);
or U3196 (N_3196,N_2818,N_2847);
and U3197 (N_3197,N_2951,N_2967);
nand U3198 (N_3198,N_2893,N_2906);
nor U3199 (N_3199,N_2841,N_2947);
or U3200 (N_3200,N_3126,N_3038);
nor U3201 (N_3201,N_3151,N_3031);
and U3202 (N_3202,N_3141,N_3192);
or U3203 (N_3203,N_3173,N_3195);
xor U3204 (N_3204,N_3129,N_3056);
nand U3205 (N_3205,N_3066,N_3013);
nor U3206 (N_3206,N_3189,N_3142);
or U3207 (N_3207,N_3080,N_3067);
or U3208 (N_3208,N_3057,N_3033);
or U3209 (N_3209,N_3042,N_3069);
or U3210 (N_3210,N_3154,N_3158);
nand U3211 (N_3211,N_3039,N_3064);
nand U3212 (N_3212,N_3132,N_3091);
nor U3213 (N_3213,N_3100,N_3007);
and U3214 (N_3214,N_3012,N_3193);
and U3215 (N_3215,N_3146,N_3155);
or U3216 (N_3216,N_3106,N_3134);
nor U3217 (N_3217,N_3183,N_3089);
or U3218 (N_3218,N_3150,N_3085);
nand U3219 (N_3219,N_3164,N_3122);
xnor U3220 (N_3220,N_3130,N_3025);
nor U3221 (N_3221,N_3112,N_3147);
and U3222 (N_3222,N_3179,N_3198);
xor U3223 (N_3223,N_3186,N_3078);
or U3224 (N_3224,N_3006,N_3019);
nor U3225 (N_3225,N_3040,N_3003);
nor U3226 (N_3226,N_3037,N_3099);
xor U3227 (N_3227,N_3167,N_3138);
xor U3228 (N_3228,N_3079,N_3088);
nor U3229 (N_3229,N_3156,N_3030);
xnor U3230 (N_3230,N_3063,N_3052);
or U3231 (N_3231,N_3087,N_3095);
or U3232 (N_3232,N_3175,N_3169);
or U3233 (N_3233,N_3086,N_3054);
and U3234 (N_3234,N_3051,N_3010);
nand U3235 (N_3235,N_3046,N_3116);
xnor U3236 (N_3236,N_3120,N_3065);
xor U3237 (N_3237,N_3090,N_3184);
xnor U3238 (N_3238,N_3117,N_3136);
xor U3239 (N_3239,N_3014,N_3199);
xnor U3240 (N_3240,N_3152,N_3143);
xor U3241 (N_3241,N_3171,N_3018);
and U3242 (N_3242,N_3190,N_3172);
and U3243 (N_3243,N_3174,N_3123);
or U3244 (N_3244,N_3165,N_3005);
nand U3245 (N_3245,N_3027,N_3118);
nor U3246 (N_3246,N_3097,N_3043);
nor U3247 (N_3247,N_3166,N_3029);
or U3248 (N_3248,N_3028,N_3177);
nor U3249 (N_3249,N_3103,N_3075);
nor U3250 (N_3250,N_3109,N_3157);
and U3251 (N_3251,N_3178,N_3124);
or U3252 (N_3252,N_3015,N_3176);
xnor U3253 (N_3253,N_3050,N_3096);
and U3254 (N_3254,N_3185,N_3004);
xor U3255 (N_3255,N_3140,N_3188);
nand U3256 (N_3256,N_3002,N_3145);
xor U3257 (N_3257,N_3016,N_3168);
nor U3258 (N_3258,N_3022,N_3160);
nand U3259 (N_3259,N_3045,N_3044);
nor U3260 (N_3260,N_3036,N_3101);
xnor U3261 (N_3261,N_3162,N_3148);
xor U3262 (N_3262,N_3094,N_3068);
nand U3263 (N_3263,N_3073,N_3113);
xor U3264 (N_3264,N_3170,N_3108);
nand U3265 (N_3265,N_3128,N_3081);
and U3266 (N_3266,N_3092,N_3009);
nand U3267 (N_3267,N_3149,N_3114);
xnor U3268 (N_3268,N_3053,N_3182);
nor U3269 (N_3269,N_3197,N_3041);
or U3270 (N_3270,N_3060,N_3180);
or U3271 (N_3271,N_3077,N_3076);
or U3272 (N_3272,N_3071,N_3061);
and U3273 (N_3273,N_3181,N_3023);
or U3274 (N_3274,N_3115,N_3049);
and U3275 (N_3275,N_3191,N_3137);
and U3276 (N_3276,N_3131,N_3159);
nor U3277 (N_3277,N_3024,N_3011);
xnor U3278 (N_3278,N_3110,N_3032);
and U3279 (N_3279,N_3194,N_3121);
nand U3280 (N_3280,N_3196,N_3058);
nor U3281 (N_3281,N_3127,N_3083);
or U3282 (N_3282,N_3084,N_3062);
xnor U3283 (N_3283,N_3098,N_3104);
nor U3284 (N_3284,N_3139,N_3070);
or U3285 (N_3285,N_3102,N_3163);
nand U3286 (N_3286,N_3008,N_3026);
or U3287 (N_3287,N_3048,N_3082);
nand U3288 (N_3288,N_3153,N_3034);
xnor U3289 (N_3289,N_3021,N_3074);
or U3290 (N_3290,N_3111,N_3105);
and U3291 (N_3291,N_3125,N_3001);
or U3292 (N_3292,N_3161,N_3135);
and U3293 (N_3293,N_3020,N_3107);
nor U3294 (N_3294,N_3017,N_3047);
or U3295 (N_3295,N_3133,N_3059);
nand U3296 (N_3296,N_3119,N_3055);
or U3297 (N_3297,N_3072,N_3144);
nand U3298 (N_3298,N_3093,N_3035);
and U3299 (N_3299,N_3187,N_3000);
nand U3300 (N_3300,N_3190,N_3123);
nand U3301 (N_3301,N_3034,N_3030);
and U3302 (N_3302,N_3017,N_3102);
nor U3303 (N_3303,N_3006,N_3004);
nor U3304 (N_3304,N_3093,N_3155);
and U3305 (N_3305,N_3089,N_3145);
nand U3306 (N_3306,N_3034,N_3101);
or U3307 (N_3307,N_3042,N_3151);
and U3308 (N_3308,N_3106,N_3089);
nor U3309 (N_3309,N_3028,N_3065);
nor U3310 (N_3310,N_3179,N_3017);
nor U3311 (N_3311,N_3007,N_3013);
nor U3312 (N_3312,N_3036,N_3198);
or U3313 (N_3313,N_3133,N_3047);
or U3314 (N_3314,N_3192,N_3041);
nand U3315 (N_3315,N_3128,N_3076);
xor U3316 (N_3316,N_3153,N_3187);
nand U3317 (N_3317,N_3103,N_3143);
nor U3318 (N_3318,N_3090,N_3003);
or U3319 (N_3319,N_3189,N_3193);
and U3320 (N_3320,N_3177,N_3088);
and U3321 (N_3321,N_3171,N_3095);
xnor U3322 (N_3322,N_3177,N_3057);
or U3323 (N_3323,N_3138,N_3122);
or U3324 (N_3324,N_3016,N_3025);
and U3325 (N_3325,N_3188,N_3019);
nand U3326 (N_3326,N_3097,N_3006);
or U3327 (N_3327,N_3179,N_3075);
nand U3328 (N_3328,N_3006,N_3101);
and U3329 (N_3329,N_3126,N_3001);
nor U3330 (N_3330,N_3197,N_3089);
or U3331 (N_3331,N_3025,N_3109);
and U3332 (N_3332,N_3114,N_3095);
nor U3333 (N_3333,N_3128,N_3172);
and U3334 (N_3334,N_3014,N_3017);
and U3335 (N_3335,N_3020,N_3110);
nand U3336 (N_3336,N_3093,N_3069);
nor U3337 (N_3337,N_3136,N_3110);
nand U3338 (N_3338,N_3177,N_3006);
or U3339 (N_3339,N_3088,N_3048);
nor U3340 (N_3340,N_3115,N_3112);
xnor U3341 (N_3341,N_3174,N_3134);
xnor U3342 (N_3342,N_3170,N_3075);
xor U3343 (N_3343,N_3096,N_3127);
or U3344 (N_3344,N_3145,N_3041);
and U3345 (N_3345,N_3173,N_3183);
and U3346 (N_3346,N_3029,N_3074);
nand U3347 (N_3347,N_3165,N_3126);
or U3348 (N_3348,N_3072,N_3170);
or U3349 (N_3349,N_3098,N_3122);
or U3350 (N_3350,N_3037,N_3101);
and U3351 (N_3351,N_3131,N_3172);
nor U3352 (N_3352,N_3138,N_3054);
nor U3353 (N_3353,N_3176,N_3110);
xor U3354 (N_3354,N_3023,N_3138);
and U3355 (N_3355,N_3177,N_3023);
xor U3356 (N_3356,N_3119,N_3052);
nand U3357 (N_3357,N_3101,N_3199);
or U3358 (N_3358,N_3186,N_3031);
nor U3359 (N_3359,N_3076,N_3172);
xor U3360 (N_3360,N_3040,N_3066);
xor U3361 (N_3361,N_3135,N_3098);
xor U3362 (N_3362,N_3174,N_3021);
nor U3363 (N_3363,N_3091,N_3006);
nand U3364 (N_3364,N_3051,N_3071);
and U3365 (N_3365,N_3028,N_3002);
nand U3366 (N_3366,N_3144,N_3130);
xor U3367 (N_3367,N_3005,N_3173);
or U3368 (N_3368,N_3121,N_3086);
and U3369 (N_3369,N_3091,N_3173);
xnor U3370 (N_3370,N_3003,N_3073);
nand U3371 (N_3371,N_3161,N_3114);
or U3372 (N_3372,N_3161,N_3068);
and U3373 (N_3373,N_3127,N_3023);
and U3374 (N_3374,N_3195,N_3066);
xor U3375 (N_3375,N_3075,N_3024);
nand U3376 (N_3376,N_3195,N_3128);
nand U3377 (N_3377,N_3142,N_3154);
xnor U3378 (N_3378,N_3025,N_3101);
or U3379 (N_3379,N_3193,N_3042);
xor U3380 (N_3380,N_3116,N_3053);
and U3381 (N_3381,N_3049,N_3136);
nor U3382 (N_3382,N_3003,N_3188);
or U3383 (N_3383,N_3074,N_3088);
xnor U3384 (N_3384,N_3172,N_3100);
or U3385 (N_3385,N_3186,N_3170);
nand U3386 (N_3386,N_3182,N_3044);
nor U3387 (N_3387,N_3150,N_3072);
xor U3388 (N_3388,N_3022,N_3066);
nor U3389 (N_3389,N_3130,N_3149);
or U3390 (N_3390,N_3079,N_3174);
or U3391 (N_3391,N_3002,N_3090);
nand U3392 (N_3392,N_3167,N_3155);
xnor U3393 (N_3393,N_3154,N_3037);
and U3394 (N_3394,N_3041,N_3049);
nor U3395 (N_3395,N_3013,N_3158);
or U3396 (N_3396,N_3002,N_3074);
nor U3397 (N_3397,N_3160,N_3044);
and U3398 (N_3398,N_3006,N_3186);
nor U3399 (N_3399,N_3111,N_3078);
and U3400 (N_3400,N_3359,N_3215);
nor U3401 (N_3401,N_3348,N_3373);
or U3402 (N_3402,N_3396,N_3315);
and U3403 (N_3403,N_3311,N_3319);
nor U3404 (N_3404,N_3216,N_3241);
or U3405 (N_3405,N_3252,N_3254);
nor U3406 (N_3406,N_3243,N_3265);
nor U3407 (N_3407,N_3251,N_3238);
and U3408 (N_3408,N_3314,N_3245);
and U3409 (N_3409,N_3271,N_3361);
xnor U3410 (N_3410,N_3240,N_3378);
and U3411 (N_3411,N_3323,N_3212);
or U3412 (N_3412,N_3304,N_3266);
and U3413 (N_3413,N_3330,N_3381);
xnor U3414 (N_3414,N_3355,N_3318);
or U3415 (N_3415,N_3325,N_3306);
or U3416 (N_3416,N_3225,N_3377);
nand U3417 (N_3417,N_3299,N_3205);
or U3418 (N_3418,N_3296,N_3365);
nor U3419 (N_3419,N_3388,N_3261);
or U3420 (N_3420,N_3263,N_3267);
or U3421 (N_3421,N_3395,N_3357);
nor U3422 (N_3422,N_3346,N_3276);
nand U3423 (N_3423,N_3344,N_3347);
nand U3424 (N_3424,N_3226,N_3356);
and U3425 (N_3425,N_3260,N_3264);
and U3426 (N_3426,N_3389,N_3201);
nor U3427 (N_3427,N_3317,N_3235);
xnor U3428 (N_3428,N_3287,N_3221);
nor U3429 (N_3429,N_3305,N_3321);
nand U3430 (N_3430,N_3393,N_3200);
nor U3431 (N_3431,N_3310,N_3326);
and U3432 (N_3432,N_3283,N_3291);
nor U3433 (N_3433,N_3229,N_3383);
and U3434 (N_3434,N_3208,N_3244);
nor U3435 (N_3435,N_3313,N_3268);
nor U3436 (N_3436,N_3248,N_3272);
and U3437 (N_3437,N_3258,N_3209);
nor U3438 (N_3438,N_3354,N_3385);
and U3439 (N_3439,N_3397,N_3239);
nor U3440 (N_3440,N_3242,N_3368);
nor U3441 (N_3441,N_3379,N_3297);
nor U3442 (N_3442,N_3340,N_3320);
and U3443 (N_3443,N_3207,N_3308);
or U3444 (N_3444,N_3222,N_3284);
xnor U3445 (N_3445,N_3275,N_3342);
nand U3446 (N_3446,N_3333,N_3211);
xnor U3447 (N_3447,N_3391,N_3329);
and U3448 (N_3448,N_3206,N_3334);
and U3449 (N_3449,N_3327,N_3390);
and U3450 (N_3450,N_3367,N_3280);
and U3451 (N_3451,N_3213,N_3210);
and U3452 (N_3452,N_3362,N_3293);
xnor U3453 (N_3453,N_3274,N_3371);
nand U3454 (N_3454,N_3302,N_3231);
nand U3455 (N_3455,N_3374,N_3233);
or U3456 (N_3456,N_3237,N_3298);
and U3457 (N_3457,N_3277,N_3380);
nand U3458 (N_3458,N_3394,N_3331);
xor U3459 (N_3459,N_3290,N_3307);
xor U3460 (N_3460,N_3382,N_3351);
or U3461 (N_3461,N_3324,N_3328);
nor U3462 (N_3462,N_3282,N_3384);
nand U3463 (N_3463,N_3341,N_3286);
xnor U3464 (N_3464,N_3303,N_3228);
nand U3465 (N_3465,N_3281,N_3218);
nor U3466 (N_3466,N_3364,N_3223);
and U3467 (N_3467,N_3269,N_3387);
nand U3468 (N_3468,N_3358,N_3295);
nor U3469 (N_3469,N_3316,N_3292);
xor U3470 (N_3470,N_3363,N_3230);
nor U3471 (N_3471,N_3337,N_3236);
nand U3472 (N_3472,N_3262,N_3339);
and U3473 (N_3473,N_3202,N_3386);
or U3474 (N_3474,N_3372,N_3256);
or U3475 (N_3475,N_3353,N_3259);
or U3476 (N_3476,N_3289,N_3336);
and U3477 (N_3477,N_3253,N_3246);
nor U3478 (N_3478,N_3214,N_3309);
xor U3479 (N_3479,N_3369,N_3370);
or U3480 (N_3480,N_3270,N_3219);
nand U3481 (N_3481,N_3345,N_3294);
or U3482 (N_3482,N_3343,N_3279);
or U3483 (N_3483,N_3232,N_3249);
and U3484 (N_3484,N_3332,N_3352);
xnor U3485 (N_3485,N_3227,N_3217);
xnor U3486 (N_3486,N_3250,N_3220);
xor U3487 (N_3487,N_3322,N_3335);
xnor U3488 (N_3488,N_3247,N_3203);
nor U3489 (N_3489,N_3399,N_3273);
and U3490 (N_3490,N_3204,N_3366);
or U3491 (N_3491,N_3350,N_3392);
and U3492 (N_3492,N_3234,N_3288);
xor U3493 (N_3493,N_3398,N_3375);
xnor U3494 (N_3494,N_3301,N_3338);
xor U3495 (N_3495,N_3360,N_3285);
and U3496 (N_3496,N_3278,N_3257);
and U3497 (N_3497,N_3376,N_3224);
nor U3498 (N_3498,N_3255,N_3300);
or U3499 (N_3499,N_3349,N_3312);
xnor U3500 (N_3500,N_3372,N_3266);
nand U3501 (N_3501,N_3292,N_3319);
and U3502 (N_3502,N_3222,N_3294);
nor U3503 (N_3503,N_3346,N_3348);
xor U3504 (N_3504,N_3220,N_3297);
nor U3505 (N_3505,N_3264,N_3388);
nand U3506 (N_3506,N_3229,N_3276);
xor U3507 (N_3507,N_3291,N_3369);
nor U3508 (N_3508,N_3295,N_3225);
nor U3509 (N_3509,N_3299,N_3262);
nand U3510 (N_3510,N_3216,N_3257);
nor U3511 (N_3511,N_3328,N_3322);
nand U3512 (N_3512,N_3286,N_3394);
and U3513 (N_3513,N_3334,N_3239);
xnor U3514 (N_3514,N_3273,N_3295);
and U3515 (N_3515,N_3349,N_3261);
xor U3516 (N_3516,N_3260,N_3238);
or U3517 (N_3517,N_3210,N_3242);
xor U3518 (N_3518,N_3327,N_3295);
and U3519 (N_3519,N_3386,N_3314);
nand U3520 (N_3520,N_3339,N_3240);
nand U3521 (N_3521,N_3373,N_3350);
and U3522 (N_3522,N_3336,N_3211);
nor U3523 (N_3523,N_3307,N_3343);
and U3524 (N_3524,N_3316,N_3252);
xor U3525 (N_3525,N_3358,N_3348);
or U3526 (N_3526,N_3259,N_3369);
nand U3527 (N_3527,N_3204,N_3300);
or U3528 (N_3528,N_3260,N_3329);
and U3529 (N_3529,N_3278,N_3288);
nor U3530 (N_3530,N_3335,N_3326);
nor U3531 (N_3531,N_3308,N_3246);
nand U3532 (N_3532,N_3268,N_3244);
xnor U3533 (N_3533,N_3376,N_3283);
nor U3534 (N_3534,N_3344,N_3398);
nor U3535 (N_3535,N_3224,N_3254);
nand U3536 (N_3536,N_3376,N_3338);
or U3537 (N_3537,N_3273,N_3250);
and U3538 (N_3538,N_3318,N_3299);
nand U3539 (N_3539,N_3294,N_3338);
and U3540 (N_3540,N_3360,N_3275);
xor U3541 (N_3541,N_3288,N_3238);
nor U3542 (N_3542,N_3396,N_3262);
xor U3543 (N_3543,N_3289,N_3250);
or U3544 (N_3544,N_3288,N_3380);
nand U3545 (N_3545,N_3339,N_3398);
nand U3546 (N_3546,N_3256,N_3216);
and U3547 (N_3547,N_3308,N_3234);
or U3548 (N_3548,N_3253,N_3283);
nand U3549 (N_3549,N_3324,N_3253);
nand U3550 (N_3550,N_3261,N_3282);
and U3551 (N_3551,N_3367,N_3335);
or U3552 (N_3552,N_3260,N_3257);
nand U3553 (N_3553,N_3382,N_3268);
nand U3554 (N_3554,N_3367,N_3260);
or U3555 (N_3555,N_3235,N_3209);
nor U3556 (N_3556,N_3385,N_3372);
nand U3557 (N_3557,N_3317,N_3205);
or U3558 (N_3558,N_3266,N_3333);
nand U3559 (N_3559,N_3278,N_3242);
nor U3560 (N_3560,N_3294,N_3307);
and U3561 (N_3561,N_3296,N_3394);
nand U3562 (N_3562,N_3267,N_3234);
or U3563 (N_3563,N_3254,N_3202);
and U3564 (N_3564,N_3231,N_3385);
or U3565 (N_3565,N_3215,N_3349);
nor U3566 (N_3566,N_3346,N_3265);
nor U3567 (N_3567,N_3230,N_3321);
nor U3568 (N_3568,N_3239,N_3336);
nor U3569 (N_3569,N_3241,N_3344);
or U3570 (N_3570,N_3291,N_3384);
nand U3571 (N_3571,N_3351,N_3315);
nand U3572 (N_3572,N_3341,N_3221);
nand U3573 (N_3573,N_3389,N_3313);
and U3574 (N_3574,N_3338,N_3235);
and U3575 (N_3575,N_3380,N_3383);
and U3576 (N_3576,N_3202,N_3209);
xnor U3577 (N_3577,N_3386,N_3200);
or U3578 (N_3578,N_3397,N_3368);
xor U3579 (N_3579,N_3397,N_3267);
nand U3580 (N_3580,N_3213,N_3250);
nand U3581 (N_3581,N_3372,N_3366);
nand U3582 (N_3582,N_3387,N_3244);
nor U3583 (N_3583,N_3213,N_3307);
nand U3584 (N_3584,N_3264,N_3238);
nor U3585 (N_3585,N_3336,N_3308);
nand U3586 (N_3586,N_3201,N_3335);
nor U3587 (N_3587,N_3323,N_3222);
nor U3588 (N_3588,N_3397,N_3395);
nand U3589 (N_3589,N_3228,N_3318);
and U3590 (N_3590,N_3296,N_3276);
xor U3591 (N_3591,N_3313,N_3211);
and U3592 (N_3592,N_3348,N_3257);
nor U3593 (N_3593,N_3378,N_3276);
nor U3594 (N_3594,N_3301,N_3361);
nor U3595 (N_3595,N_3251,N_3321);
nand U3596 (N_3596,N_3348,N_3343);
nand U3597 (N_3597,N_3311,N_3228);
or U3598 (N_3598,N_3218,N_3289);
xnor U3599 (N_3599,N_3344,N_3324);
or U3600 (N_3600,N_3490,N_3429);
and U3601 (N_3601,N_3416,N_3472);
or U3602 (N_3602,N_3526,N_3413);
nor U3603 (N_3603,N_3488,N_3451);
nor U3604 (N_3604,N_3421,N_3443);
nand U3605 (N_3605,N_3541,N_3497);
xnor U3606 (N_3606,N_3598,N_3410);
and U3607 (N_3607,N_3529,N_3583);
or U3608 (N_3608,N_3407,N_3500);
xor U3609 (N_3609,N_3570,N_3512);
nand U3610 (N_3610,N_3462,N_3491);
nand U3611 (N_3611,N_3556,N_3597);
xor U3612 (N_3612,N_3502,N_3523);
or U3613 (N_3613,N_3554,N_3439);
nor U3614 (N_3614,N_3571,N_3542);
and U3615 (N_3615,N_3474,N_3404);
nand U3616 (N_3616,N_3585,N_3485);
nand U3617 (N_3617,N_3587,N_3511);
or U3618 (N_3618,N_3543,N_3418);
and U3619 (N_3619,N_3509,N_3454);
xnor U3620 (N_3620,N_3469,N_3520);
nor U3621 (N_3621,N_3465,N_3470);
or U3622 (N_3622,N_3591,N_3463);
or U3623 (N_3623,N_3577,N_3401);
xor U3624 (N_3624,N_3422,N_3513);
nand U3625 (N_3625,N_3563,N_3524);
and U3626 (N_3626,N_3517,N_3449);
nor U3627 (N_3627,N_3546,N_3547);
xor U3628 (N_3628,N_3483,N_3433);
nor U3629 (N_3629,N_3535,N_3540);
xor U3630 (N_3630,N_3514,N_3544);
xor U3631 (N_3631,N_3414,N_3412);
nor U3632 (N_3632,N_3492,N_3521);
nor U3633 (N_3633,N_3559,N_3417);
or U3634 (N_3634,N_3549,N_3552);
nor U3635 (N_3635,N_3473,N_3420);
or U3636 (N_3636,N_3567,N_3586);
and U3637 (N_3637,N_3530,N_3450);
nand U3638 (N_3638,N_3578,N_3440);
or U3639 (N_3639,N_3402,N_3565);
nor U3640 (N_3640,N_3489,N_3484);
and U3641 (N_3641,N_3411,N_3499);
nor U3642 (N_3642,N_3548,N_3475);
or U3643 (N_3643,N_3522,N_3561);
or U3644 (N_3644,N_3564,N_3581);
and U3645 (N_3645,N_3536,N_3467);
nor U3646 (N_3646,N_3441,N_3539);
or U3647 (N_3647,N_3507,N_3452);
nand U3648 (N_3648,N_3464,N_3400);
nor U3649 (N_3649,N_3589,N_3466);
and U3650 (N_3650,N_3493,N_3506);
nand U3651 (N_3651,N_3592,N_3498);
nand U3652 (N_3652,N_3518,N_3456);
nor U3653 (N_3653,N_3432,N_3476);
nor U3654 (N_3654,N_3423,N_3480);
or U3655 (N_3655,N_3496,N_3447);
and U3656 (N_3656,N_3428,N_3445);
or U3657 (N_3657,N_3588,N_3505);
and U3658 (N_3658,N_3582,N_3482);
xnor U3659 (N_3659,N_3551,N_3495);
and U3660 (N_3660,N_3550,N_3486);
or U3661 (N_3661,N_3504,N_3458);
and U3662 (N_3662,N_3430,N_3455);
nand U3663 (N_3663,N_3487,N_3427);
nand U3664 (N_3664,N_3560,N_3408);
or U3665 (N_3665,N_3508,N_3576);
and U3666 (N_3666,N_3527,N_3442);
nand U3667 (N_3667,N_3436,N_3534);
or U3668 (N_3668,N_3579,N_3479);
nand U3669 (N_3669,N_3460,N_3446);
and U3670 (N_3670,N_3453,N_3438);
nand U3671 (N_3671,N_3537,N_3569);
nor U3672 (N_3672,N_3515,N_3405);
xor U3673 (N_3673,N_3573,N_3415);
xor U3674 (N_3674,N_3566,N_3580);
or U3675 (N_3675,N_3533,N_3575);
nand U3676 (N_3676,N_3403,N_3584);
or U3677 (N_3677,N_3477,N_3457);
xor U3678 (N_3678,N_3532,N_3431);
xnor U3679 (N_3679,N_3461,N_3459);
nand U3680 (N_3680,N_3419,N_3562);
and U3681 (N_3681,N_3545,N_3426);
nor U3682 (N_3682,N_3590,N_3444);
nand U3683 (N_3683,N_3596,N_3593);
xor U3684 (N_3684,N_3599,N_3574);
nand U3685 (N_3685,N_3531,N_3435);
xor U3686 (N_3686,N_3471,N_3406);
xnor U3687 (N_3687,N_3525,N_3557);
nand U3688 (N_3688,N_3528,N_3568);
nand U3689 (N_3689,N_3425,N_3553);
and U3690 (N_3690,N_3555,N_3519);
xor U3691 (N_3691,N_3494,N_3409);
nor U3692 (N_3692,N_3595,N_3510);
nand U3693 (N_3693,N_3468,N_3503);
or U3694 (N_3694,N_3538,N_3478);
and U3695 (N_3695,N_3434,N_3437);
xor U3696 (N_3696,N_3424,N_3501);
nor U3697 (N_3697,N_3594,N_3481);
or U3698 (N_3698,N_3572,N_3516);
and U3699 (N_3699,N_3448,N_3558);
nand U3700 (N_3700,N_3586,N_3526);
or U3701 (N_3701,N_3493,N_3426);
or U3702 (N_3702,N_3568,N_3508);
and U3703 (N_3703,N_3429,N_3451);
nor U3704 (N_3704,N_3511,N_3500);
and U3705 (N_3705,N_3578,N_3476);
nor U3706 (N_3706,N_3512,N_3591);
xnor U3707 (N_3707,N_3580,N_3560);
and U3708 (N_3708,N_3493,N_3527);
nor U3709 (N_3709,N_3540,N_3545);
nand U3710 (N_3710,N_3404,N_3421);
or U3711 (N_3711,N_3542,N_3418);
or U3712 (N_3712,N_3519,N_3503);
and U3713 (N_3713,N_3509,N_3535);
and U3714 (N_3714,N_3509,N_3578);
xor U3715 (N_3715,N_3599,N_3406);
nand U3716 (N_3716,N_3404,N_3424);
nor U3717 (N_3717,N_3523,N_3450);
or U3718 (N_3718,N_3472,N_3596);
and U3719 (N_3719,N_3423,N_3432);
xor U3720 (N_3720,N_3462,N_3496);
nand U3721 (N_3721,N_3542,N_3495);
or U3722 (N_3722,N_3426,N_3508);
nand U3723 (N_3723,N_3454,N_3535);
nor U3724 (N_3724,N_3424,N_3562);
nor U3725 (N_3725,N_3522,N_3519);
nand U3726 (N_3726,N_3522,N_3459);
xnor U3727 (N_3727,N_3501,N_3583);
or U3728 (N_3728,N_3523,N_3599);
nor U3729 (N_3729,N_3575,N_3460);
and U3730 (N_3730,N_3431,N_3429);
nor U3731 (N_3731,N_3483,N_3471);
and U3732 (N_3732,N_3438,N_3575);
or U3733 (N_3733,N_3518,N_3564);
xnor U3734 (N_3734,N_3528,N_3532);
or U3735 (N_3735,N_3564,N_3497);
xor U3736 (N_3736,N_3490,N_3463);
nand U3737 (N_3737,N_3400,N_3505);
or U3738 (N_3738,N_3599,N_3409);
xor U3739 (N_3739,N_3546,N_3591);
and U3740 (N_3740,N_3477,N_3456);
or U3741 (N_3741,N_3565,N_3574);
nand U3742 (N_3742,N_3470,N_3512);
nand U3743 (N_3743,N_3518,N_3426);
and U3744 (N_3744,N_3573,N_3435);
nand U3745 (N_3745,N_3596,N_3419);
nand U3746 (N_3746,N_3519,N_3599);
xnor U3747 (N_3747,N_3495,N_3588);
and U3748 (N_3748,N_3549,N_3514);
or U3749 (N_3749,N_3527,N_3441);
nor U3750 (N_3750,N_3455,N_3447);
nand U3751 (N_3751,N_3497,N_3490);
or U3752 (N_3752,N_3552,N_3453);
nand U3753 (N_3753,N_3446,N_3496);
nor U3754 (N_3754,N_3427,N_3555);
nor U3755 (N_3755,N_3554,N_3570);
xor U3756 (N_3756,N_3568,N_3504);
nand U3757 (N_3757,N_3596,N_3520);
and U3758 (N_3758,N_3406,N_3450);
nand U3759 (N_3759,N_3460,N_3424);
or U3760 (N_3760,N_3524,N_3442);
and U3761 (N_3761,N_3413,N_3580);
nor U3762 (N_3762,N_3528,N_3515);
xnor U3763 (N_3763,N_3497,N_3577);
or U3764 (N_3764,N_3449,N_3488);
and U3765 (N_3765,N_3519,N_3457);
nor U3766 (N_3766,N_3525,N_3406);
nor U3767 (N_3767,N_3429,N_3480);
or U3768 (N_3768,N_3454,N_3543);
and U3769 (N_3769,N_3444,N_3541);
nand U3770 (N_3770,N_3414,N_3497);
xnor U3771 (N_3771,N_3526,N_3415);
and U3772 (N_3772,N_3478,N_3497);
and U3773 (N_3773,N_3550,N_3423);
and U3774 (N_3774,N_3471,N_3411);
nand U3775 (N_3775,N_3480,N_3503);
nand U3776 (N_3776,N_3571,N_3439);
or U3777 (N_3777,N_3425,N_3437);
nor U3778 (N_3778,N_3479,N_3486);
nor U3779 (N_3779,N_3559,N_3533);
nor U3780 (N_3780,N_3445,N_3599);
xor U3781 (N_3781,N_3470,N_3472);
nand U3782 (N_3782,N_3503,N_3570);
nor U3783 (N_3783,N_3537,N_3455);
nor U3784 (N_3784,N_3420,N_3490);
and U3785 (N_3785,N_3476,N_3510);
xnor U3786 (N_3786,N_3479,N_3420);
xnor U3787 (N_3787,N_3493,N_3460);
and U3788 (N_3788,N_3498,N_3465);
nand U3789 (N_3789,N_3415,N_3447);
xnor U3790 (N_3790,N_3415,N_3568);
nor U3791 (N_3791,N_3588,N_3491);
xnor U3792 (N_3792,N_3551,N_3586);
nor U3793 (N_3793,N_3437,N_3440);
and U3794 (N_3794,N_3505,N_3413);
xnor U3795 (N_3795,N_3542,N_3589);
or U3796 (N_3796,N_3563,N_3464);
and U3797 (N_3797,N_3484,N_3403);
and U3798 (N_3798,N_3415,N_3407);
xor U3799 (N_3799,N_3416,N_3535);
xnor U3800 (N_3800,N_3629,N_3637);
or U3801 (N_3801,N_3699,N_3719);
or U3802 (N_3802,N_3673,N_3617);
nor U3803 (N_3803,N_3683,N_3635);
nand U3804 (N_3804,N_3791,N_3651);
or U3805 (N_3805,N_3650,N_3727);
xor U3806 (N_3806,N_3752,N_3711);
xnor U3807 (N_3807,N_3761,N_3609);
nand U3808 (N_3808,N_3643,N_3670);
nor U3809 (N_3809,N_3689,N_3797);
nor U3810 (N_3810,N_3615,N_3760);
and U3811 (N_3811,N_3721,N_3776);
nand U3812 (N_3812,N_3747,N_3697);
and U3813 (N_3813,N_3764,N_3724);
xnor U3814 (N_3814,N_3620,N_3785);
nand U3815 (N_3815,N_3630,N_3777);
and U3816 (N_3816,N_3744,N_3649);
or U3817 (N_3817,N_3624,N_3675);
xor U3818 (N_3818,N_3743,N_3745);
or U3819 (N_3819,N_3680,N_3723);
nand U3820 (N_3820,N_3728,N_3715);
xor U3821 (N_3821,N_3755,N_3606);
xor U3822 (N_3822,N_3634,N_3706);
nand U3823 (N_3823,N_3799,N_3687);
xnor U3824 (N_3824,N_3748,N_3774);
xor U3825 (N_3825,N_3654,N_3779);
or U3826 (N_3826,N_3773,N_3664);
nor U3827 (N_3827,N_3746,N_3766);
nand U3828 (N_3828,N_3681,N_3713);
xnor U3829 (N_3829,N_3759,N_3682);
or U3830 (N_3830,N_3717,N_3667);
or U3831 (N_3831,N_3738,N_3603);
xor U3832 (N_3832,N_3605,N_3647);
nor U3833 (N_3833,N_3663,N_3705);
nor U3834 (N_3834,N_3616,N_3787);
and U3835 (N_3835,N_3685,N_3691);
nand U3836 (N_3836,N_3636,N_3781);
nand U3837 (N_3837,N_3611,N_3739);
nor U3838 (N_3838,N_3631,N_3622);
nor U3839 (N_3839,N_3729,N_3703);
and U3840 (N_3840,N_3753,N_3621);
nand U3841 (N_3841,N_3775,N_3741);
and U3842 (N_3842,N_3619,N_3742);
nand U3843 (N_3843,N_3679,N_3704);
or U3844 (N_3844,N_3608,N_3790);
nor U3845 (N_3845,N_3757,N_3734);
or U3846 (N_3846,N_3716,N_3690);
xor U3847 (N_3847,N_3710,N_3770);
xnor U3848 (N_3848,N_3698,N_3701);
or U3849 (N_3849,N_3639,N_3794);
or U3850 (N_3850,N_3633,N_3661);
and U3851 (N_3851,N_3771,N_3686);
or U3852 (N_3852,N_3600,N_3618);
nand U3853 (N_3853,N_3731,N_3749);
nand U3854 (N_3854,N_3694,N_3660);
and U3855 (N_3855,N_3750,N_3718);
nand U3856 (N_3856,N_3767,N_3688);
or U3857 (N_3857,N_3788,N_3625);
and U3858 (N_3858,N_3638,N_3754);
and U3859 (N_3859,N_3726,N_3700);
nand U3860 (N_3860,N_3758,N_3778);
or U3861 (N_3861,N_3626,N_3662);
nand U3862 (N_3862,N_3632,N_3784);
or U3863 (N_3863,N_3659,N_3708);
and U3864 (N_3864,N_3786,N_3740);
nand U3865 (N_3865,N_3602,N_3684);
or U3866 (N_3866,N_3607,N_3737);
xnor U3867 (N_3867,N_3725,N_3614);
or U3868 (N_3868,N_3730,N_3722);
or U3869 (N_3869,N_3665,N_3628);
or U3870 (N_3870,N_3610,N_3669);
or U3871 (N_3871,N_3627,N_3656);
xor U3872 (N_3872,N_3709,N_3658);
nand U3873 (N_3873,N_3601,N_3756);
xnor U3874 (N_3874,N_3648,N_3736);
nor U3875 (N_3875,N_3652,N_3780);
nor U3876 (N_3876,N_3641,N_3733);
nor U3877 (N_3877,N_3612,N_3646);
xor U3878 (N_3878,N_3672,N_3692);
and U3879 (N_3879,N_3676,N_3604);
xnor U3880 (N_3880,N_3623,N_3678);
or U3881 (N_3881,N_3789,N_3735);
and U3882 (N_3882,N_3762,N_3671);
nor U3883 (N_3883,N_3657,N_3666);
or U3884 (N_3884,N_3640,N_3714);
and U3885 (N_3885,N_3696,N_3720);
or U3886 (N_3886,N_3693,N_3769);
or U3887 (N_3887,N_3751,N_3674);
nor U3888 (N_3888,N_3783,N_3613);
nand U3889 (N_3889,N_3677,N_3763);
nand U3890 (N_3890,N_3668,N_3798);
nand U3891 (N_3891,N_3655,N_3782);
or U3892 (N_3892,N_3707,N_3793);
nor U3893 (N_3893,N_3772,N_3768);
nor U3894 (N_3894,N_3702,N_3795);
nor U3895 (N_3895,N_3796,N_3645);
nand U3896 (N_3896,N_3695,N_3653);
or U3897 (N_3897,N_3712,N_3644);
nor U3898 (N_3898,N_3642,N_3765);
nand U3899 (N_3899,N_3732,N_3792);
nor U3900 (N_3900,N_3660,N_3632);
or U3901 (N_3901,N_3658,N_3785);
nor U3902 (N_3902,N_3724,N_3793);
nor U3903 (N_3903,N_3709,N_3619);
xor U3904 (N_3904,N_3683,N_3793);
xnor U3905 (N_3905,N_3683,N_3637);
nand U3906 (N_3906,N_3617,N_3789);
or U3907 (N_3907,N_3651,N_3649);
nand U3908 (N_3908,N_3778,N_3688);
or U3909 (N_3909,N_3744,N_3728);
and U3910 (N_3910,N_3717,N_3662);
nor U3911 (N_3911,N_3773,N_3660);
nor U3912 (N_3912,N_3712,N_3748);
nor U3913 (N_3913,N_3749,N_3771);
xor U3914 (N_3914,N_3696,N_3703);
nand U3915 (N_3915,N_3617,N_3766);
and U3916 (N_3916,N_3688,N_3677);
or U3917 (N_3917,N_3741,N_3651);
and U3918 (N_3918,N_3729,N_3661);
nor U3919 (N_3919,N_3762,N_3601);
and U3920 (N_3920,N_3636,N_3706);
and U3921 (N_3921,N_3695,N_3778);
or U3922 (N_3922,N_3737,N_3711);
and U3923 (N_3923,N_3766,N_3613);
or U3924 (N_3924,N_3682,N_3631);
nor U3925 (N_3925,N_3792,N_3779);
or U3926 (N_3926,N_3681,N_3632);
xor U3927 (N_3927,N_3799,N_3768);
nor U3928 (N_3928,N_3667,N_3666);
nand U3929 (N_3929,N_3686,N_3743);
and U3930 (N_3930,N_3661,N_3671);
and U3931 (N_3931,N_3735,N_3617);
xor U3932 (N_3932,N_3795,N_3641);
or U3933 (N_3933,N_3741,N_3725);
or U3934 (N_3934,N_3795,N_3651);
nand U3935 (N_3935,N_3710,N_3748);
and U3936 (N_3936,N_3710,N_3617);
nor U3937 (N_3937,N_3737,N_3741);
xnor U3938 (N_3938,N_3727,N_3645);
or U3939 (N_3939,N_3767,N_3618);
nand U3940 (N_3940,N_3616,N_3630);
or U3941 (N_3941,N_3622,N_3601);
and U3942 (N_3942,N_3616,N_3791);
or U3943 (N_3943,N_3684,N_3679);
and U3944 (N_3944,N_3734,N_3788);
or U3945 (N_3945,N_3629,N_3747);
nand U3946 (N_3946,N_3689,N_3749);
and U3947 (N_3947,N_3600,N_3625);
nand U3948 (N_3948,N_3728,N_3711);
or U3949 (N_3949,N_3689,N_3777);
or U3950 (N_3950,N_3793,N_3772);
xor U3951 (N_3951,N_3647,N_3662);
nor U3952 (N_3952,N_3621,N_3721);
and U3953 (N_3953,N_3609,N_3792);
and U3954 (N_3954,N_3767,N_3681);
and U3955 (N_3955,N_3659,N_3696);
or U3956 (N_3956,N_3735,N_3731);
xnor U3957 (N_3957,N_3779,N_3651);
nand U3958 (N_3958,N_3690,N_3710);
nor U3959 (N_3959,N_3709,N_3720);
nor U3960 (N_3960,N_3603,N_3628);
and U3961 (N_3961,N_3751,N_3750);
xnor U3962 (N_3962,N_3712,N_3768);
xnor U3963 (N_3963,N_3735,N_3616);
nor U3964 (N_3964,N_3727,N_3708);
and U3965 (N_3965,N_3684,N_3726);
nor U3966 (N_3966,N_3698,N_3721);
and U3967 (N_3967,N_3788,N_3658);
nor U3968 (N_3968,N_3610,N_3786);
and U3969 (N_3969,N_3676,N_3788);
nand U3970 (N_3970,N_3632,N_3728);
and U3971 (N_3971,N_3619,N_3728);
xnor U3972 (N_3972,N_3604,N_3629);
xnor U3973 (N_3973,N_3791,N_3668);
xor U3974 (N_3974,N_3602,N_3763);
or U3975 (N_3975,N_3779,N_3653);
xnor U3976 (N_3976,N_3782,N_3695);
and U3977 (N_3977,N_3696,N_3605);
nor U3978 (N_3978,N_3668,N_3600);
nor U3979 (N_3979,N_3702,N_3636);
xnor U3980 (N_3980,N_3722,N_3726);
nand U3981 (N_3981,N_3782,N_3600);
and U3982 (N_3982,N_3724,N_3648);
nand U3983 (N_3983,N_3734,N_3719);
or U3984 (N_3984,N_3652,N_3681);
xnor U3985 (N_3985,N_3760,N_3799);
nand U3986 (N_3986,N_3766,N_3688);
xnor U3987 (N_3987,N_3655,N_3673);
and U3988 (N_3988,N_3783,N_3666);
and U3989 (N_3989,N_3618,N_3672);
nor U3990 (N_3990,N_3682,N_3788);
nor U3991 (N_3991,N_3784,N_3709);
xor U3992 (N_3992,N_3739,N_3758);
or U3993 (N_3993,N_3737,N_3658);
nand U3994 (N_3994,N_3634,N_3710);
nand U3995 (N_3995,N_3659,N_3600);
and U3996 (N_3996,N_3600,N_3793);
nand U3997 (N_3997,N_3631,N_3730);
and U3998 (N_3998,N_3713,N_3709);
xor U3999 (N_3999,N_3763,N_3703);
or U4000 (N_4000,N_3859,N_3913);
or U4001 (N_4001,N_3922,N_3877);
nor U4002 (N_4002,N_3973,N_3879);
nor U4003 (N_4003,N_3992,N_3830);
nor U4004 (N_4004,N_3820,N_3962);
and U4005 (N_4005,N_3919,N_3801);
nand U4006 (N_4006,N_3905,N_3835);
and U4007 (N_4007,N_3903,N_3822);
nor U4008 (N_4008,N_3845,N_3950);
nor U4009 (N_4009,N_3897,N_3999);
or U4010 (N_4010,N_3951,N_3906);
nand U4011 (N_4011,N_3967,N_3865);
xor U4012 (N_4012,N_3867,N_3971);
or U4013 (N_4013,N_3963,N_3969);
nor U4014 (N_4014,N_3964,N_3812);
nand U4015 (N_4015,N_3948,N_3981);
nor U4016 (N_4016,N_3979,N_3895);
and U4017 (N_4017,N_3930,N_3956);
or U4018 (N_4018,N_3952,N_3954);
nor U4019 (N_4019,N_3840,N_3957);
or U4020 (N_4020,N_3890,N_3996);
xnor U4021 (N_4021,N_3838,N_3953);
and U4022 (N_4022,N_3887,N_3866);
nor U4023 (N_4023,N_3857,N_3871);
nand U4024 (N_4024,N_3975,N_3818);
and U4025 (N_4025,N_3892,N_3809);
nand U4026 (N_4026,N_3824,N_3885);
and U4027 (N_4027,N_3886,N_3873);
and U4028 (N_4028,N_3938,N_3931);
or U4029 (N_4029,N_3803,N_3862);
and U4030 (N_4030,N_3884,N_3904);
or U4031 (N_4031,N_3933,N_3861);
xnor U4032 (N_4032,N_3978,N_3937);
nand U4033 (N_4033,N_3970,N_3984);
or U4034 (N_4034,N_3907,N_3856);
nand U4035 (N_4035,N_3825,N_3831);
nor U4036 (N_4036,N_3917,N_3908);
or U4037 (N_4037,N_3961,N_3945);
nor U4038 (N_4038,N_3805,N_3814);
xor U4039 (N_4039,N_3888,N_3842);
and U4040 (N_4040,N_3853,N_3878);
nand U4041 (N_4041,N_3910,N_3921);
xnor U4042 (N_4042,N_3816,N_3974);
nand U4043 (N_4043,N_3934,N_3839);
and U4044 (N_4044,N_3960,N_3965);
nor U4045 (N_4045,N_3843,N_3935);
nor U4046 (N_4046,N_3918,N_3883);
and U4047 (N_4047,N_3943,N_3985);
and U4048 (N_4048,N_3946,N_3914);
or U4049 (N_4049,N_3989,N_3990);
and U4050 (N_4050,N_3902,N_3896);
and U4051 (N_4051,N_3939,N_3844);
nor U4052 (N_4052,N_3899,N_3958);
or U4053 (N_4053,N_3834,N_3941);
nor U4054 (N_4054,N_3864,N_3912);
xnor U4055 (N_4055,N_3852,N_3972);
nand U4056 (N_4056,N_3909,N_3993);
nor U4057 (N_4057,N_3829,N_3928);
nand U4058 (N_4058,N_3841,N_3942);
xor U4059 (N_4059,N_3959,N_3807);
or U4060 (N_4060,N_3920,N_3846);
xor U4061 (N_4061,N_3987,N_3947);
and U4062 (N_4062,N_3977,N_3940);
nor U4063 (N_4063,N_3923,N_3995);
nand U4064 (N_4064,N_3936,N_3806);
nand U4065 (N_4065,N_3968,N_3875);
nor U4066 (N_4066,N_3915,N_3929);
and U4067 (N_4067,N_3881,N_3836);
nand U4068 (N_4068,N_3924,N_3893);
nor U4069 (N_4069,N_3982,N_3813);
xor U4070 (N_4070,N_3837,N_3832);
or U4071 (N_4071,N_3870,N_3944);
and U4072 (N_4072,N_3802,N_3983);
xor U4073 (N_4073,N_3819,N_3826);
nor U4074 (N_4074,N_3815,N_3901);
and U4075 (N_4075,N_3882,N_3991);
nand U4076 (N_4076,N_3828,N_3804);
nand U4077 (N_4077,N_3849,N_3949);
or U4078 (N_4078,N_3891,N_3874);
and U4079 (N_4079,N_3955,N_3858);
nand U4080 (N_4080,N_3926,N_3817);
or U4081 (N_4081,N_3833,N_3800);
xnor U4082 (N_4082,N_3868,N_3927);
xnor U4083 (N_4083,N_3911,N_3850);
and U4084 (N_4084,N_3880,N_3916);
and U4085 (N_4085,N_3998,N_3827);
and U4086 (N_4086,N_3900,N_3848);
nor U4087 (N_4087,N_3821,N_3925);
or U4088 (N_4088,N_3863,N_3810);
nand U4089 (N_4089,N_3894,N_3811);
nor U4090 (N_4090,N_3966,N_3994);
or U4091 (N_4091,N_3860,N_3872);
nor U4092 (N_4092,N_3869,N_3876);
xor U4093 (N_4093,N_3851,N_3932);
nor U4094 (N_4094,N_3976,N_3898);
nor U4095 (N_4095,N_3823,N_3847);
or U4096 (N_4096,N_3997,N_3980);
nor U4097 (N_4097,N_3986,N_3988);
and U4098 (N_4098,N_3854,N_3808);
nand U4099 (N_4099,N_3855,N_3889);
and U4100 (N_4100,N_3997,N_3977);
nor U4101 (N_4101,N_3986,N_3892);
xnor U4102 (N_4102,N_3802,N_3962);
xnor U4103 (N_4103,N_3950,N_3857);
and U4104 (N_4104,N_3951,N_3928);
nor U4105 (N_4105,N_3916,N_3871);
xor U4106 (N_4106,N_3893,N_3949);
or U4107 (N_4107,N_3956,N_3942);
nor U4108 (N_4108,N_3973,N_3825);
nand U4109 (N_4109,N_3858,N_3938);
xnor U4110 (N_4110,N_3833,N_3831);
nand U4111 (N_4111,N_3905,N_3805);
nor U4112 (N_4112,N_3943,N_3849);
nand U4113 (N_4113,N_3885,N_3975);
xnor U4114 (N_4114,N_3883,N_3875);
xor U4115 (N_4115,N_3982,N_3920);
and U4116 (N_4116,N_3934,N_3875);
or U4117 (N_4117,N_3851,N_3923);
nor U4118 (N_4118,N_3811,N_3887);
and U4119 (N_4119,N_3963,N_3860);
and U4120 (N_4120,N_3816,N_3814);
nand U4121 (N_4121,N_3908,N_3881);
nor U4122 (N_4122,N_3874,N_3811);
xnor U4123 (N_4123,N_3899,N_3835);
nor U4124 (N_4124,N_3910,N_3824);
and U4125 (N_4125,N_3871,N_3865);
nor U4126 (N_4126,N_3999,N_3966);
nand U4127 (N_4127,N_3925,N_3820);
nand U4128 (N_4128,N_3917,N_3984);
nor U4129 (N_4129,N_3890,N_3913);
nor U4130 (N_4130,N_3922,N_3854);
and U4131 (N_4131,N_3913,N_3981);
nor U4132 (N_4132,N_3888,N_3884);
or U4133 (N_4133,N_3990,N_3911);
nor U4134 (N_4134,N_3910,N_3967);
xnor U4135 (N_4135,N_3816,N_3836);
nand U4136 (N_4136,N_3929,N_3951);
xor U4137 (N_4137,N_3804,N_3968);
xor U4138 (N_4138,N_3821,N_3943);
and U4139 (N_4139,N_3970,N_3900);
or U4140 (N_4140,N_3861,N_3810);
or U4141 (N_4141,N_3987,N_3817);
nor U4142 (N_4142,N_3998,N_3852);
and U4143 (N_4143,N_3884,N_3843);
nand U4144 (N_4144,N_3992,N_3930);
xnor U4145 (N_4145,N_3859,N_3996);
xor U4146 (N_4146,N_3815,N_3942);
xor U4147 (N_4147,N_3860,N_3804);
nor U4148 (N_4148,N_3947,N_3844);
nand U4149 (N_4149,N_3978,N_3806);
and U4150 (N_4150,N_3823,N_3813);
nand U4151 (N_4151,N_3847,N_3874);
or U4152 (N_4152,N_3909,N_3937);
nand U4153 (N_4153,N_3857,N_3891);
nor U4154 (N_4154,N_3917,N_3816);
nor U4155 (N_4155,N_3901,N_3976);
xor U4156 (N_4156,N_3866,N_3908);
xor U4157 (N_4157,N_3905,N_3910);
or U4158 (N_4158,N_3892,N_3847);
nor U4159 (N_4159,N_3962,N_3909);
or U4160 (N_4160,N_3834,N_3875);
and U4161 (N_4161,N_3919,N_3888);
nor U4162 (N_4162,N_3985,N_3850);
nor U4163 (N_4163,N_3856,N_3924);
nand U4164 (N_4164,N_3959,N_3912);
and U4165 (N_4165,N_3853,N_3818);
nor U4166 (N_4166,N_3802,N_3880);
nor U4167 (N_4167,N_3927,N_3841);
or U4168 (N_4168,N_3863,N_3957);
or U4169 (N_4169,N_3850,N_3839);
xnor U4170 (N_4170,N_3831,N_3875);
nand U4171 (N_4171,N_3922,N_3827);
and U4172 (N_4172,N_3803,N_3948);
or U4173 (N_4173,N_3881,N_3812);
nand U4174 (N_4174,N_3890,N_3993);
xnor U4175 (N_4175,N_3912,N_3898);
nand U4176 (N_4176,N_3879,N_3840);
or U4177 (N_4177,N_3822,N_3999);
xnor U4178 (N_4178,N_3994,N_3991);
or U4179 (N_4179,N_3861,N_3958);
nand U4180 (N_4180,N_3844,N_3893);
and U4181 (N_4181,N_3935,N_3870);
and U4182 (N_4182,N_3880,N_3990);
nor U4183 (N_4183,N_3819,N_3997);
xnor U4184 (N_4184,N_3895,N_3865);
and U4185 (N_4185,N_3816,N_3892);
nand U4186 (N_4186,N_3875,N_3930);
xnor U4187 (N_4187,N_3853,N_3913);
nor U4188 (N_4188,N_3947,N_3927);
and U4189 (N_4189,N_3986,N_3953);
nand U4190 (N_4190,N_3856,N_3822);
and U4191 (N_4191,N_3915,N_3873);
and U4192 (N_4192,N_3814,N_3956);
nand U4193 (N_4193,N_3869,N_3808);
nand U4194 (N_4194,N_3894,N_3807);
nor U4195 (N_4195,N_3821,N_3970);
nand U4196 (N_4196,N_3942,N_3924);
nor U4197 (N_4197,N_3819,N_3976);
nand U4198 (N_4198,N_3945,N_3939);
xor U4199 (N_4199,N_3967,N_3803);
nor U4200 (N_4200,N_4190,N_4078);
or U4201 (N_4201,N_4141,N_4108);
nand U4202 (N_4202,N_4050,N_4059);
nor U4203 (N_4203,N_4147,N_4189);
nand U4204 (N_4204,N_4086,N_4063);
nor U4205 (N_4205,N_4116,N_4162);
nor U4206 (N_4206,N_4045,N_4186);
nor U4207 (N_4207,N_4173,N_4129);
or U4208 (N_4208,N_4156,N_4058);
nor U4209 (N_4209,N_4046,N_4111);
nor U4210 (N_4210,N_4198,N_4197);
or U4211 (N_4211,N_4069,N_4168);
xor U4212 (N_4212,N_4160,N_4085);
nand U4213 (N_4213,N_4099,N_4021);
nor U4214 (N_4214,N_4145,N_4096);
nand U4215 (N_4215,N_4179,N_4133);
xor U4216 (N_4216,N_4163,N_4033);
xor U4217 (N_4217,N_4054,N_4070);
and U4218 (N_4218,N_4164,N_4126);
nand U4219 (N_4219,N_4074,N_4065);
nand U4220 (N_4220,N_4068,N_4082);
or U4221 (N_4221,N_4088,N_4150);
nand U4222 (N_4222,N_4114,N_4073);
or U4223 (N_4223,N_4007,N_4006);
and U4224 (N_4224,N_4064,N_4098);
xor U4225 (N_4225,N_4158,N_4060);
nor U4226 (N_4226,N_4191,N_4009);
and U4227 (N_4227,N_4148,N_4041);
nor U4228 (N_4228,N_4022,N_4053);
nand U4229 (N_4229,N_4003,N_4015);
nor U4230 (N_4230,N_4030,N_4130);
xor U4231 (N_4231,N_4176,N_4194);
or U4232 (N_4232,N_4062,N_4180);
xor U4233 (N_4233,N_4020,N_4127);
nor U4234 (N_4234,N_4093,N_4044);
nor U4235 (N_4235,N_4090,N_4018);
nor U4236 (N_4236,N_4101,N_4138);
and U4237 (N_4237,N_4095,N_4055);
or U4238 (N_4238,N_4137,N_4120);
xor U4239 (N_4239,N_4155,N_4036);
xnor U4240 (N_4240,N_4187,N_4121);
and U4241 (N_4241,N_4031,N_4172);
nand U4242 (N_4242,N_4113,N_4104);
xor U4243 (N_4243,N_4097,N_4136);
or U4244 (N_4244,N_4185,N_4011);
nor U4245 (N_4245,N_4174,N_4029);
nor U4246 (N_4246,N_4183,N_4013);
xnor U4247 (N_4247,N_4010,N_4028);
xor U4248 (N_4248,N_4142,N_4023);
and U4249 (N_4249,N_4083,N_4102);
nor U4250 (N_4250,N_4094,N_4056);
and U4251 (N_4251,N_4115,N_4170);
nor U4252 (N_4252,N_4135,N_4112);
xnor U4253 (N_4253,N_4152,N_4181);
xnor U4254 (N_4254,N_4140,N_4017);
nand U4255 (N_4255,N_4057,N_4146);
nor U4256 (N_4256,N_4080,N_4109);
nand U4257 (N_4257,N_4084,N_4125);
xnor U4258 (N_4258,N_4161,N_4128);
nand U4259 (N_4259,N_4134,N_4040);
xnor U4260 (N_4260,N_4014,N_4081);
nand U4261 (N_4261,N_4153,N_4066);
or U4262 (N_4262,N_4171,N_4144);
nor U4263 (N_4263,N_4032,N_4106);
nor U4264 (N_4264,N_4043,N_4092);
nand U4265 (N_4265,N_4124,N_4002);
or U4266 (N_4266,N_4024,N_4004);
xnor U4267 (N_4267,N_4117,N_4034);
and U4268 (N_4268,N_4077,N_4118);
and U4269 (N_4269,N_4061,N_4182);
xor U4270 (N_4270,N_4157,N_4119);
xnor U4271 (N_4271,N_4035,N_4166);
and U4272 (N_4272,N_4131,N_4076);
xnor U4273 (N_4273,N_4196,N_4001);
nand U4274 (N_4274,N_4178,N_4123);
and U4275 (N_4275,N_4167,N_4000);
nor U4276 (N_4276,N_4087,N_4079);
and U4277 (N_4277,N_4052,N_4100);
nor U4278 (N_4278,N_4105,N_4175);
xor U4279 (N_4279,N_4103,N_4177);
nand U4280 (N_4280,N_4195,N_4075);
xnor U4281 (N_4281,N_4047,N_4005);
nor U4282 (N_4282,N_4067,N_4139);
and U4283 (N_4283,N_4184,N_4132);
nor U4284 (N_4284,N_4192,N_4165);
nand U4285 (N_4285,N_4149,N_4169);
nor U4286 (N_4286,N_4089,N_4091);
nor U4287 (N_4287,N_4154,N_4048);
or U4288 (N_4288,N_4008,N_4037);
xnor U4289 (N_4289,N_4122,N_4107);
or U4290 (N_4290,N_4071,N_4143);
nand U4291 (N_4291,N_4193,N_4012);
and U4292 (N_4292,N_4016,N_4199);
nor U4293 (N_4293,N_4188,N_4072);
nor U4294 (N_4294,N_4026,N_4051);
xor U4295 (N_4295,N_4159,N_4027);
nor U4296 (N_4296,N_4049,N_4042);
or U4297 (N_4297,N_4025,N_4110);
or U4298 (N_4298,N_4019,N_4039);
nand U4299 (N_4299,N_4151,N_4038);
nor U4300 (N_4300,N_4092,N_4076);
xnor U4301 (N_4301,N_4160,N_4156);
and U4302 (N_4302,N_4162,N_4138);
and U4303 (N_4303,N_4034,N_4116);
or U4304 (N_4304,N_4188,N_4076);
xnor U4305 (N_4305,N_4100,N_4150);
or U4306 (N_4306,N_4133,N_4030);
or U4307 (N_4307,N_4109,N_4111);
nand U4308 (N_4308,N_4109,N_4057);
or U4309 (N_4309,N_4048,N_4042);
xor U4310 (N_4310,N_4042,N_4085);
nand U4311 (N_4311,N_4110,N_4186);
and U4312 (N_4312,N_4082,N_4189);
xor U4313 (N_4313,N_4005,N_4085);
and U4314 (N_4314,N_4018,N_4074);
and U4315 (N_4315,N_4011,N_4142);
or U4316 (N_4316,N_4167,N_4183);
and U4317 (N_4317,N_4156,N_4048);
xor U4318 (N_4318,N_4164,N_4145);
xnor U4319 (N_4319,N_4137,N_4027);
or U4320 (N_4320,N_4104,N_4169);
or U4321 (N_4321,N_4003,N_4045);
or U4322 (N_4322,N_4187,N_4196);
and U4323 (N_4323,N_4139,N_4146);
xor U4324 (N_4324,N_4101,N_4142);
or U4325 (N_4325,N_4186,N_4008);
nand U4326 (N_4326,N_4193,N_4059);
and U4327 (N_4327,N_4199,N_4050);
or U4328 (N_4328,N_4017,N_4096);
xor U4329 (N_4329,N_4013,N_4161);
nand U4330 (N_4330,N_4163,N_4023);
nor U4331 (N_4331,N_4004,N_4143);
nor U4332 (N_4332,N_4136,N_4007);
xnor U4333 (N_4333,N_4026,N_4191);
or U4334 (N_4334,N_4086,N_4002);
or U4335 (N_4335,N_4146,N_4105);
or U4336 (N_4336,N_4053,N_4089);
or U4337 (N_4337,N_4171,N_4062);
and U4338 (N_4338,N_4114,N_4116);
nor U4339 (N_4339,N_4118,N_4058);
or U4340 (N_4340,N_4138,N_4015);
nand U4341 (N_4341,N_4111,N_4105);
and U4342 (N_4342,N_4057,N_4197);
and U4343 (N_4343,N_4197,N_4032);
and U4344 (N_4344,N_4090,N_4100);
nand U4345 (N_4345,N_4183,N_4001);
nor U4346 (N_4346,N_4183,N_4094);
and U4347 (N_4347,N_4132,N_4046);
nor U4348 (N_4348,N_4095,N_4134);
xor U4349 (N_4349,N_4054,N_4183);
and U4350 (N_4350,N_4122,N_4170);
xnor U4351 (N_4351,N_4155,N_4097);
xnor U4352 (N_4352,N_4189,N_4031);
nor U4353 (N_4353,N_4034,N_4018);
and U4354 (N_4354,N_4117,N_4135);
and U4355 (N_4355,N_4128,N_4087);
or U4356 (N_4356,N_4011,N_4013);
or U4357 (N_4357,N_4168,N_4034);
nand U4358 (N_4358,N_4071,N_4029);
and U4359 (N_4359,N_4097,N_4087);
xnor U4360 (N_4360,N_4127,N_4177);
nor U4361 (N_4361,N_4063,N_4105);
xor U4362 (N_4362,N_4179,N_4067);
and U4363 (N_4363,N_4031,N_4091);
xor U4364 (N_4364,N_4197,N_4181);
nor U4365 (N_4365,N_4170,N_4001);
nor U4366 (N_4366,N_4000,N_4047);
nand U4367 (N_4367,N_4064,N_4044);
xor U4368 (N_4368,N_4010,N_4017);
or U4369 (N_4369,N_4185,N_4040);
xnor U4370 (N_4370,N_4128,N_4025);
nand U4371 (N_4371,N_4183,N_4047);
or U4372 (N_4372,N_4056,N_4059);
or U4373 (N_4373,N_4046,N_4067);
or U4374 (N_4374,N_4156,N_4001);
and U4375 (N_4375,N_4039,N_4197);
nand U4376 (N_4376,N_4128,N_4140);
or U4377 (N_4377,N_4055,N_4167);
nor U4378 (N_4378,N_4035,N_4143);
nor U4379 (N_4379,N_4141,N_4107);
or U4380 (N_4380,N_4053,N_4087);
or U4381 (N_4381,N_4140,N_4102);
nor U4382 (N_4382,N_4031,N_4013);
xor U4383 (N_4383,N_4037,N_4161);
or U4384 (N_4384,N_4033,N_4100);
xnor U4385 (N_4385,N_4067,N_4090);
nand U4386 (N_4386,N_4147,N_4116);
xnor U4387 (N_4387,N_4156,N_4060);
and U4388 (N_4388,N_4085,N_4019);
or U4389 (N_4389,N_4091,N_4129);
and U4390 (N_4390,N_4138,N_4126);
and U4391 (N_4391,N_4015,N_4051);
nand U4392 (N_4392,N_4014,N_4139);
or U4393 (N_4393,N_4182,N_4183);
or U4394 (N_4394,N_4126,N_4027);
or U4395 (N_4395,N_4014,N_4153);
or U4396 (N_4396,N_4002,N_4079);
nand U4397 (N_4397,N_4006,N_4095);
nor U4398 (N_4398,N_4191,N_4086);
and U4399 (N_4399,N_4091,N_4054);
xor U4400 (N_4400,N_4374,N_4211);
or U4401 (N_4401,N_4265,N_4391);
or U4402 (N_4402,N_4384,N_4208);
nor U4403 (N_4403,N_4318,N_4249);
nor U4404 (N_4404,N_4336,N_4282);
or U4405 (N_4405,N_4328,N_4223);
and U4406 (N_4406,N_4314,N_4321);
nand U4407 (N_4407,N_4362,N_4288);
and U4408 (N_4408,N_4242,N_4316);
and U4409 (N_4409,N_4298,N_4258);
nand U4410 (N_4410,N_4326,N_4370);
xnor U4411 (N_4411,N_4308,N_4279);
or U4412 (N_4412,N_4335,N_4226);
and U4413 (N_4413,N_4270,N_4218);
and U4414 (N_4414,N_4204,N_4262);
nand U4415 (N_4415,N_4360,N_4236);
nor U4416 (N_4416,N_4274,N_4250);
or U4417 (N_4417,N_4216,N_4319);
nor U4418 (N_4418,N_4214,N_4395);
and U4419 (N_4419,N_4387,N_4306);
nand U4420 (N_4420,N_4244,N_4296);
nor U4421 (N_4421,N_4289,N_4213);
or U4422 (N_4422,N_4348,N_4295);
xor U4423 (N_4423,N_4359,N_4327);
xnor U4424 (N_4424,N_4220,N_4245);
nor U4425 (N_4425,N_4202,N_4369);
nand U4426 (N_4426,N_4325,N_4361);
xor U4427 (N_4427,N_4247,N_4355);
nor U4428 (N_4428,N_4263,N_4379);
or U4429 (N_4429,N_4378,N_4261);
nand U4430 (N_4430,N_4290,N_4397);
or U4431 (N_4431,N_4390,N_4230);
xnor U4432 (N_4432,N_4256,N_4252);
and U4433 (N_4433,N_4219,N_4353);
and U4434 (N_4434,N_4217,N_4373);
xnor U4435 (N_4435,N_4210,N_4382);
xor U4436 (N_4436,N_4205,N_4372);
xnor U4437 (N_4437,N_4225,N_4315);
and U4438 (N_4438,N_4364,N_4313);
nand U4439 (N_4439,N_4281,N_4206);
nor U4440 (N_4440,N_4300,N_4293);
nand U4441 (N_4441,N_4255,N_4303);
nand U4442 (N_4442,N_4292,N_4273);
and U4443 (N_4443,N_4354,N_4254);
nand U4444 (N_4444,N_4341,N_4294);
nand U4445 (N_4445,N_4330,N_4302);
xor U4446 (N_4446,N_4238,N_4345);
or U4447 (N_4447,N_4367,N_4349);
or U4448 (N_4448,N_4394,N_4253);
or U4449 (N_4449,N_4232,N_4285);
or U4450 (N_4450,N_4264,N_4371);
nor U4451 (N_4451,N_4200,N_4277);
nor U4452 (N_4452,N_4333,N_4251);
nor U4453 (N_4453,N_4358,N_4332);
nand U4454 (N_4454,N_4299,N_4320);
nand U4455 (N_4455,N_4385,N_4234);
or U4456 (N_4456,N_4398,N_4203);
or U4457 (N_4457,N_4305,N_4337);
xor U4458 (N_4458,N_4393,N_4227);
xnor U4459 (N_4459,N_4368,N_4271);
and U4460 (N_4460,N_4363,N_4260);
and U4461 (N_4461,N_4346,N_4283);
nand U4462 (N_4462,N_4304,N_4381);
nor U4463 (N_4463,N_4248,N_4257);
xor U4464 (N_4464,N_4380,N_4329);
xor U4465 (N_4465,N_4356,N_4224);
nand U4466 (N_4466,N_4243,N_4259);
xnor U4467 (N_4467,N_4229,N_4311);
xnor U4468 (N_4468,N_4383,N_4352);
or U4469 (N_4469,N_4392,N_4386);
nand U4470 (N_4470,N_4399,N_4275);
nor U4471 (N_4471,N_4340,N_4344);
or U4472 (N_4472,N_4239,N_4351);
nor U4473 (N_4473,N_4267,N_4228);
nand U4474 (N_4474,N_4331,N_4241);
or U4475 (N_4475,N_4339,N_4221);
or U4476 (N_4476,N_4338,N_4286);
nor U4477 (N_4477,N_4209,N_4278);
nand U4478 (N_4478,N_4291,N_4246);
or U4479 (N_4479,N_4301,N_4317);
nand U4480 (N_4480,N_4347,N_4357);
and U4481 (N_4481,N_4376,N_4343);
or U4482 (N_4482,N_4212,N_4233);
nand U4483 (N_4483,N_4297,N_4389);
nand U4484 (N_4484,N_4268,N_4377);
nor U4485 (N_4485,N_4334,N_4235);
xnor U4486 (N_4486,N_4266,N_4240);
nand U4487 (N_4487,N_4396,N_4280);
nand U4488 (N_4488,N_4276,N_4231);
or U4489 (N_4489,N_4312,N_4342);
nor U4490 (N_4490,N_4207,N_4284);
nand U4491 (N_4491,N_4215,N_4388);
nor U4492 (N_4492,N_4324,N_4309);
or U4493 (N_4493,N_4269,N_4322);
nand U4494 (N_4494,N_4323,N_4201);
nor U4495 (N_4495,N_4222,N_4307);
nor U4496 (N_4496,N_4287,N_4272);
nor U4497 (N_4497,N_4237,N_4366);
nor U4498 (N_4498,N_4310,N_4350);
nor U4499 (N_4499,N_4375,N_4365);
or U4500 (N_4500,N_4328,N_4350);
and U4501 (N_4501,N_4211,N_4203);
or U4502 (N_4502,N_4296,N_4344);
and U4503 (N_4503,N_4375,N_4217);
and U4504 (N_4504,N_4307,N_4367);
and U4505 (N_4505,N_4238,N_4335);
nor U4506 (N_4506,N_4357,N_4281);
or U4507 (N_4507,N_4288,N_4273);
and U4508 (N_4508,N_4302,N_4212);
nor U4509 (N_4509,N_4224,N_4286);
or U4510 (N_4510,N_4271,N_4230);
xnor U4511 (N_4511,N_4205,N_4248);
xor U4512 (N_4512,N_4375,N_4379);
or U4513 (N_4513,N_4303,N_4323);
and U4514 (N_4514,N_4277,N_4341);
or U4515 (N_4515,N_4291,N_4289);
xor U4516 (N_4516,N_4261,N_4361);
nor U4517 (N_4517,N_4264,N_4388);
and U4518 (N_4518,N_4371,N_4286);
nand U4519 (N_4519,N_4291,N_4300);
or U4520 (N_4520,N_4346,N_4261);
nand U4521 (N_4521,N_4256,N_4277);
nor U4522 (N_4522,N_4206,N_4397);
nor U4523 (N_4523,N_4201,N_4298);
and U4524 (N_4524,N_4243,N_4388);
and U4525 (N_4525,N_4318,N_4342);
xor U4526 (N_4526,N_4344,N_4254);
nor U4527 (N_4527,N_4384,N_4236);
xor U4528 (N_4528,N_4261,N_4270);
nand U4529 (N_4529,N_4375,N_4351);
nor U4530 (N_4530,N_4361,N_4311);
xor U4531 (N_4531,N_4393,N_4282);
and U4532 (N_4532,N_4241,N_4380);
or U4533 (N_4533,N_4367,N_4312);
nand U4534 (N_4534,N_4280,N_4209);
xor U4535 (N_4535,N_4371,N_4334);
xnor U4536 (N_4536,N_4247,N_4263);
and U4537 (N_4537,N_4267,N_4201);
or U4538 (N_4538,N_4276,N_4241);
nor U4539 (N_4539,N_4262,N_4330);
and U4540 (N_4540,N_4275,N_4233);
xor U4541 (N_4541,N_4278,N_4358);
nand U4542 (N_4542,N_4291,N_4316);
or U4543 (N_4543,N_4201,N_4352);
nor U4544 (N_4544,N_4390,N_4329);
xnor U4545 (N_4545,N_4238,N_4296);
nor U4546 (N_4546,N_4285,N_4222);
nor U4547 (N_4547,N_4394,N_4337);
xnor U4548 (N_4548,N_4388,N_4340);
or U4549 (N_4549,N_4399,N_4264);
xnor U4550 (N_4550,N_4272,N_4214);
nor U4551 (N_4551,N_4385,N_4384);
nand U4552 (N_4552,N_4283,N_4305);
and U4553 (N_4553,N_4359,N_4207);
nor U4554 (N_4554,N_4228,N_4247);
and U4555 (N_4555,N_4278,N_4296);
and U4556 (N_4556,N_4268,N_4308);
nor U4557 (N_4557,N_4216,N_4266);
or U4558 (N_4558,N_4347,N_4372);
or U4559 (N_4559,N_4348,N_4302);
or U4560 (N_4560,N_4394,N_4307);
nor U4561 (N_4561,N_4332,N_4353);
or U4562 (N_4562,N_4337,N_4296);
nor U4563 (N_4563,N_4276,N_4224);
and U4564 (N_4564,N_4259,N_4235);
or U4565 (N_4565,N_4292,N_4385);
and U4566 (N_4566,N_4271,N_4292);
xor U4567 (N_4567,N_4379,N_4340);
and U4568 (N_4568,N_4319,N_4239);
nor U4569 (N_4569,N_4226,N_4235);
and U4570 (N_4570,N_4272,N_4308);
nand U4571 (N_4571,N_4399,N_4356);
nand U4572 (N_4572,N_4220,N_4320);
xnor U4573 (N_4573,N_4250,N_4251);
nor U4574 (N_4574,N_4345,N_4328);
or U4575 (N_4575,N_4252,N_4273);
or U4576 (N_4576,N_4313,N_4306);
and U4577 (N_4577,N_4276,N_4352);
nand U4578 (N_4578,N_4399,N_4253);
xor U4579 (N_4579,N_4372,N_4391);
and U4580 (N_4580,N_4291,N_4354);
nand U4581 (N_4581,N_4318,N_4200);
and U4582 (N_4582,N_4364,N_4352);
nand U4583 (N_4583,N_4371,N_4359);
xor U4584 (N_4584,N_4359,N_4386);
and U4585 (N_4585,N_4248,N_4246);
nor U4586 (N_4586,N_4203,N_4391);
or U4587 (N_4587,N_4321,N_4231);
xor U4588 (N_4588,N_4389,N_4300);
xor U4589 (N_4589,N_4380,N_4374);
nand U4590 (N_4590,N_4237,N_4256);
or U4591 (N_4591,N_4307,N_4219);
xor U4592 (N_4592,N_4392,N_4396);
nand U4593 (N_4593,N_4233,N_4324);
or U4594 (N_4594,N_4219,N_4291);
and U4595 (N_4595,N_4328,N_4374);
and U4596 (N_4596,N_4373,N_4261);
nand U4597 (N_4597,N_4374,N_4387);
nor U4598 (N_4598,N_4217,N_4284);
nor U4599 (N_4599,N_4260,N_4288);
xor U4600 (N_4600,N_4489,N_4574);
or U4601 (N_4601,N_4464,N_4554);
nor U4602 (N_4602,N_4434,N_4555);
nor U4603 (N_4603,N_4427,N_4479);
or U4604 (N_4604,N_4473,N_4506);
nor U4605 (N_4605,N_4496,N_4482);
or U4606 (N_4606,N_4586,N_4589);
nand U4607 (N_4607,N_4546,N_4543);
nor U4608 (N_4608,N_4519,N_4444);
and U4609 (N_4609,N_4592,N_4532);
xor U4610 (N_4610,N_4420,N_4558);
nor U4611 (N_4611,N_4469,N_4407);
xor U4612 (N_4612,N_4440,N_4557);
or U4613 (N_4613,N_4597,N_4432);
or U4614 (N_4614,N_4591,N_4425);
xnor U4615 (N_4615,N_4566,N_4581);
nor U4616 (N_4616,N_4494,N_4426);
nand U4617 (N_4617,N_4499,N_4450);
or U4618 (N_4618,N_4595,N_4477);
nand U4619 (N_4619,N_4486,N_4488);
nand U4620 (N_4620,N_4578,N_4553);
xnor U4621 (N_4621,N_4556,N_4405);
or U4622 (N_4622,N_4525,N_4562);
nand U4623 (N_4623,N_4573,N_4483);
nand U4624 (N_4624,N_4510,N_4474);
nand U4625 (N_4625,N_4548,N_4570);
xor U4626 (N_4626,N_4416,N_4435);
nand U4627 (N_4627,N_4534,N_4528);
xnor U4628 (N_4628,N_4403,N_4413);
or U4629 (N_4629,N_4536,N_4422);
nor U4630 (N_4630,N_4447,N_4448);
nand U4631 (N_4631,N_4599,N_4585);
xor U4632 (N_4632,N_4431,N_4409);
nand U4633 (N_4633,N_4421,N_4455);
nor U4634 (N_4634,N_4576,N_4560);
and U4635 (N_4635,N_4593,N_4590);
nand U4636 (N_4636,N_4502,N_4402);
xnor U4637 (N_4637,N_4584,N_4476);
nand U4638 (N_4638,N_4454,N_4484);
nand U4639 (N_4639,N_4439,N_4514);
or U4640 (N_4640,N_4485,N_4437);
nor U4641 (N_4641,N_4563,N_4516);
or U4642 (N_4642,N_4478,N_4461);
nor U4643 (N_4643,N_4547,N_4412);
nor U4644 (N_4644,N_4531,N_4527);
and U4645 (N_4645,N_4517,N_4419);
nand U4646 (N_4646,N_4433,N_4411);
xor U4647 (N_4647,N_4436,N_4513);
and U4648 (N_4648,N_4491,N_4598);
and U4649 (N_4649,N_4452,N_4508);
nor U4650 (N_4650,N_4400,N_4518);
nand U4651 (N_4651,N_4544,N_4580);
nor U4652 (N_4652,N_4569,N_4538);
and U4653 (N_4653,N_4559,N_4551);
xor U4654 (N_4654,N_4524,N_4530);
xnor U4655 (N_4655,N_4501,N_4571);
and U4656 (N_4656,N_4453,N_4442);
or U4657 (N_4657,N_4415,N_4458);
or U4658 (N_4658,N_4511,N_4568);
and U4659 (N_4659,N_4429,N_4509);
nand U4660 (N_4660,N_4404,N_4428);
xnor U4661 (N_4661,N_4583,N_4468);
or U4662 (N_4662,N_4490,N_4500);
nand U4663 (N_4663,N_4441,N_4572);
and U4664 (N_4664,N_4467,N_4503);
or U4665 (N_4665,N_4504,N_4577);
nand U4666 (N_4666,N_4423,N_4410);
and U4667 (N_4667,N_4549,N_4417);
nor U4668 (N_4668,N_4575,N_4424);
xnor U4669 (N_4669,N_4451,N_4588);
or U4670 (N_4670,N_4564,N_4462);
xnor U4671 (N_4671,N_4498,N_4545);
nor U4672 (N_4672,N_4471,N_4515);
nor U4673 (N_4673,N_4418,N_4596);
nor U4674 (N_4674,N_4443,N_4582);
xnor U4675 (N_4675,N_4408,N_4430);
nor U4676 (N_4676,N_4497,N_4487);
and U4677 (N_4677,N_4523,N_4526);
xnor U4678 (N_4678,N_4537,N_4540);
nand U4679 (N_4679,N_4512,N_4579);
xnor U4680 (N_4680,N_4495,N_4470);
nand U4681 (N_4681,N_4463,N_4438);
nor U4682 (N_4682,N_4521,N_4480);
nand U4683 (N_4683,N_4522,N_4449);
nand U4684 (N_4684,N_4481,N_4542);
or U4685 (N_4685,N_4507,N_4529);
or U4686 (N_4686,N_4552,N_4414);
and U4687 (N_4687,N_4587,N_4565);
nand U4688 (N_4688,N_4505,N_4459);
nand U4689 (N_4689,N_4533,N_4466);
xor U4690 (N_4690,N_4550,N_4535);
or U4691 (N_4691,N_4465,N_4406);
and U4692 (N_4692,N_4472,N_4520);
xnor U4693 (N_4693,N_4492,N_4460);
nand U4694 (N_4694,N_4457,N_4493);
nor U4695 (N_4695,N_4475,N_4567);
nand U4696 (N_4696,N_4594,N_4561);
nor U4697 (N_4697,N_4541,N_4539);
and U4698 (N_4698,N_4456,N_4445);
xnor U4699 (N_4699,N_4401,N_4446);
or U4700 (N_4700,N_4496,N_4469);
xor U4701 (N_4701,N_4411,N_4496);
nand U4702 (N_4702,N_4588,N_4511);
and U4703 (N_4703,N_4538,N_4590);
and U4704 (N_4704,N_4428,N_4590);
or U4705 (N_4705,N_4433,N_4408);
xor U4706 (N_4706,N_4556,N_4457);
or U4707 (N_4707,N_4554,N_4521);
and U4708 (N_4708,N_4514,N_4458);
nand U4709 (N_4709,N_4483,N_4599);
xnor U4710 (N_4710,N_4466,N_4581);
nor U4711 (N_4711,N_4538,N_4408);
nand U4712 (N_4712,N_4448,N_4464);
xor U4713 (N_4713,N_4416,N_4589);
nand U4714 (N_4714,N_4448,N_4516);
nand U4715 (N_4715,N_4454,N_4590);
nor U4716 (N_4716,N_4588,N_4416);
and U4717 (N_4717,N_4558,N_4520);
nand U4718 (N_4718,N_4574,N_4400);
or U4719 (N_4719,N_4485,N_4488);
nor U4720 (N_4720,N_4500,N_4476);
nor U4721 (N_4721,N_4443,N_4551);
nor U4722 (N_4722,N_4499,N_4528);
or U4723 (N_4723,N_4497,N_4455);
nand U4724 (N_4724,N_4512,N_4422);
xnor U4725 (N_4725,N_4563,N_4595);
and U4726 (N_4726,N_4472,N_4492);
xnor U4727 (N_4727,N_4483,N_4591);
or U4728 (N_4728,N_4431,N_4562);
nand U4729 (N_4729,N_4417,N_4444);
nor U4730 (N_4730,N_4405,N_4419);
nand U4731 (N_4731,N_4502,N_4536);
nand U4732 (N_4732,N_4538,N_4552);
xnor U4733 (N_4733,N_4489,N_4439);
xor U4734 (N_4734,N_4427,N_4499);
and U4735 (N_4735,N_4596,N_4535);
nand U4736 (N_4736,N_4493,N_4542);
nor U4737 (N_4737,N_4505,N_4482);
and U4738 (N_4738,N_4495,N_4591);
xor U4739 (N_4739,N_4452,N_4526);
xnor U4740 (N_4740,N_4471,N_4502);
xnor U4741 (N_4741,N_4450,N_4479);
nand U4742 (N_4742,N_4501,N_4550);
nor U4743 (N_4743,N_4515,N_4566);
nor U4744 (N_4744,N_4547,N_4434);
nand U4745 (N_4745,N_4570,N_4509);
nor U4746 (N_4746,N_4452,N_4541);
xor U4747 (N_4747,N_4402,N_4549);
nor U4748 (N_4748,N_4492,N_4502);
or U4749 (N_4749,N_4404,N_4438);
or U4750 (N_4750,N_4579,N_4439);
xnor U4751 (N_4751,N_4535,N_4571);
xor U4752 (N_4752,N_4431,N_4542);
nor U4753 (N_4753,N_4529,N_4409);
and U4754 (N_4754,N_4570,N_4564);
or U4755 (N_4755,N_4568,N_4587);
or U4756 (N_4756,N_4591,N_4461);
and U4757 (N_4757,N_4559,N_4478);
and U4758 (N_4758,N_4547,N_4494);
nand U4759 (N_4759,N_4413,N_4554);
or U4760 (N_4760,N_4494,N_4500);
nor U4761 (N_4761,N_4535,N_4481);
nor U4762 (N_4762,N_4487,N_4574);
or U4763 (N_4763,N_4420,N_4418);
or U4764 (N_4764,N_4440,N_4453);
and U4765 (N_4765,N_4462,N_4430);
nand U4766 (N_4766,N_4514,N_4436);
xor U4767 (N_4767,N_4473,N_4562);
and U4768 (N_4768,N_4416,N_4501);
or U4769 (N_4769,N_4499,N_4480);
xor U4770 (N_4770,N_4523,N_4486);
nand U4771 (N_4771,N_4450,N_4562);
and U4772 (N_4772,N_4516,N_4482);
xor U4773 (N_4773,N_4599,N_4403);
nor U4774 (N_4774,N_4444,N_4556);
and U4775 (N_4775,N_4476,N_4499);
nor U4776 (N_4776,N_4530,N_4550);
nor U4777 (N_4777,N_4513,N_4550);
nor U4778 (N_4778,N_4409,N_4544);
or U4779 (N_4779,N_4505,N_4598);
or U4780 (N_4780,N_4497,N_4479);
nand U4781 (N_4781,N_4574,N_4571);
nor U4782 (N_4782,N_4563,N_4517);
nor U4783 (N_4783,N_4491,N_4567);
or U4784 (N_4784,N_4543,N_4426);
nor U4785 (N_4785,N_4594,N_4510);
or U4786 (N_4786,N_4518,N_4548);
and U4787 (N_4787,N_4507,N_4535);
and U4788 (N_4788,N_4533,N_4408);
nand U4789 (N_4789,N_4468,N_4544);
xnor U4790 (N_4790,N_4499,N_4537);
xor U4791 (N_4791,N_4508,N_4433);
or U4792 (N_4792,N_4586,N_4569);
xnor U4793 (N_4793,N_4572,N_4503);
and U4794 (N_4794,N_4403,N_4470);
or U4795 (N_4795,N_4573,N_4517);
nand U4796 (N_4796,N_4431,N_4413);
nor U4797 (N_4797,N_4471,N_4404);
nor U4798 (N_4798,N_4586,N_4442);
or U4799 (N_4799,N_4574,N_4430);
and U4800 (N_4800,N_4648,N_4746);
nand U4801 (N_4801,N_4737,N_4781);
and U4802 (N_4802,N_4755,N_4756);
and U4803 (N_4803,N_4727,N_4773);
and U4804 (N_4804,N_4687,N_4743);
and U4805 (N_4805,N_4751,N_4766);
or U4806 (N_4806,N_4714,N_4679);
xnor U4807 (N_4807,N_4612,N_4702);
nor U4808 (N_4808,N_4658,N_4762);
nand U4809 (N_4809,N_4778,N_4626);
or U4810 (N_4810,N_4661,N_4749);
nor U4811 (N_4811,N_4733,N_4771);
nand U4812 (N_4812,N_4681,N_4744);
nor U4813 (N_4813,N_4631,N_4682);
or U4814 (N_4814,N_4639,N_4772);
or U4815 (N_4815,N_4685,N_4622);
nor U4816 (N_4816,N_4720,N_4660);
and U4817 (N_4817,N_4786,N_4796);
or U4818 (N_4818,N_4705,N_4767);
or U4819 (N_4819,N_4764,N_4676);
or U4820 (N_4820,N_4712,N_4719);
and U4821 (N_4821,N_4604,N_4704);
nand U4822 (N_4822,N_4613,N_4640);
or U4823 (N_4823,N_4698,N_4638);
or U4824 (N_4824,N_4793,N_4745);
nand U4825 (N_4825,N_4754,N_4721);
nand U4826 (N_4826,N_4627,N_4670);
and U4827 (N_4827,N_4699,N_4625);
and U4828 (N_4828,N_4747,N_4668);
or U4829 (N_4829,N_4601,N_4758);
nand U4830 (N_4830,N_4618,N_4689);
nand U4831 (N_4831,N_4610,N_4665);
xnor U4832 (N_4832,N_4726,N_4730);
nand U4833 (N_4833,N_4715,N_4798);
and U4834 (N_4834,N_4605,N_4652);
nand U4835 (N_4835,N_4600,N_4633);
nor U4836 (N_4836,N_4779,N_4635);
and U4837 (N_4837,N_4630,N_4710);
xnor U4838 (N_4838,N_4775,N_4619);
nor U4839 (N_4839,N_4628,N_4617);
nand U4840 (N_4840,N_4683,N_4697);
nand U4841 (N_4841,N_4717,N_4760);
nand U4842 (N_4842,N_4761,N_4782);
or U4843 (N_4843,N_4700,N_4784);
xor U4844 (N_4844,N_4653,N_4728);
nor U4845 (N_4845,N_4713,N_4656);
or U4846 (N_4846,N_4723,N_4711);
xor U4847 (N_4847,N_4606,N_4794);
or U4848 (N_4848,N_4799,N_4603);
nor U4849 (N_4849,N_4738,N_4611);
or U4850 (N_4850,N_4791,N_4787);
nor U4851 (N_4851,N_4690,N_4752);
xor U4852 (N_4852,N_4768,N_4789);
and U4853 (N_4853,N_4675,N_4680);
nand U4854 (N_4854,N_4674,N_4607);
nor U4855 (N_4855,N_4795,N_4616);
or U4856 (N_4856,N_4722,N_4739);
and U4857 (N_4857,N_4691,N_4777);
and U4858 (N_4858,N_4763,N_4792);
nor U4859 (N_4859,N_4783,N_4678);
xor U4860 (N_4860,N_4669,N_4732);
nor U4861 (N_4861,N_4731,N_4688);
or U4862 (N_4862,N_4694,N_4788);
nand U4863 (N_4863,N_4602,N_4729);
and U4864 (N_4864,N_4634,N_4757);
xor U4865 (N_4865,N_4742,N_4701);
nand U4866 (N_4866,N_4636,N_4692);
nand U4867 (N_4867,N_4624,N_4769);
xor U4868 (N_4868,N_4671,N_4696);
xnor U4869 (N_4869,N_4655,N_4666);
nor U4870 (N_4870,N_4765,N_4663);
xnor U4871 (N_4871,N_4659,N_4753);
nand U4872 (N_4872,N_4662,N_4693);
nor U4873 (N_4873,N_4632,N_4647);
and U4874 (N_4874,N_4759,N_4748);
nor U4875 (N_4875,N_4621,N_4708);
nand U4876 (N_4876,N_4620,N_4724);
or U4877 (N_4877,N_4649,N_4686);
nor U4878 (N_4878,N_4637,N_4776);
xor U4879 (N_4879,N_4750,N_4608);
xnor U4880 (N_4880,N_4695,N_4718);
xnor U4881 (N_4881,N_4734,N_4673);
and U4882 (N_4882,N_4642,N_4650);
nand U4883 (N_4883,N_4706,N_4797);
nand U4884 (N_4884,N_4770,N_4709);
nand U4885 (N_4885,N_4684,N_4667);
nor U4886 (N_4886,N_4672,N_4644);
nand U4887 (N_4887,N_4740,N_4646);
nand U4888 (N_4888,N_4657,N_4645);
and U4889 (N_4889,N_4735,N_4790);
or U4890 (N_4890,N_4716,N_4654);
or U4891 (N_4891,N_4614,N_4615);
nor U4892 (N_4892,N_4741,N_4774);
or U4893 (N_4893,N_4677,N_4651);
nand U4894 (N_4894,N_4785,N_4609);
or U4895 (N_4895,N_4643,N_4641);
or U4896 (N_4896,N_4664,N_4623);
or U4897 (N_4897,N_4736,N_4707);
xnor U4898 (N_4898,N_4703,N_4629);
xnor U4899 (N_4899,N_4780,N_4725);
xor U4900 (N_4900,N_4601,N_4792);
nor U4901 (N_4901,N_4703,N_4708);
or U4902 (N_4902,N_4708,N_4636);
nand U4903 (N_4903,N_4700,N_4660);
or U4904 (N_4904,N_4798,N_4742);
nor U4905 (N_4905,N_4647,N_4655);
nor U4906 (N_4906,N_4645,N_4697);
or U4907 (N_4907,N_4654,N_4729);
xor U4908 (N_4908,N_4797,N_4777);
nor U4909 (N_4909,N_4623,N_4715);
nor U4910 (N_4910,N_4727,N_4628);
and U4911 (N_4911,N_4745,N_4649);
and U4912 (N_4912,N_4680,N_4664);
nand U4913 (N_4913,N_4681,N_4692);
nand U4914 (N_4914,N_4738,N_4662);
or U4915 (N_4915,N_4675,N_4709);
xor U4916 (N_4916,N_4687,N_4762);
or U4917 (N_4917,N_4788,N_4733);
or U4918 (N_4918,N_4695,N_4624);
nand U4919 (N_4919,N_4693,N_4670);
nor U4920 (N_4920,N_4682,N_4788);
and U4921 (N_4921,N_4621,N_4637);
and U4922 (N_4922,N_4630,N_4786);
and U4923 (N_4923,N_4700,N_4713);
xnor U4924 (N_4924,N_4644,N_4642);
and U4925 (N_4925,N_4720,N_4798);
and U4926 (N_4926,N_4669,N_4637);
and U4927 (N_4927,N_4654,N_4617);
nand U4928 (N_4928,N_4701,N_4765);
and U4929 (N_4929,N_4712,N_4601);
and U4930 (N_4930,N_4720,N_4791);
xnor U4931 (N_4931,N_4666,N_4794);
or U4932 (N_4932,N_4721,N_4763);
xor U4933 (N_4933,N_4787,N_4651);
nand U4934 (N_4934,N_4799,N_4718);
xor U4935 (N_4935,N_4768,N_4718);
nor U4936 (N_4936,N_4661,N_4794);
nor U4937 (N_4937,N_4764,N_4710);
xnor U4938 (N_4938,N_4741,N_4763);
and U4939 (N_4939,N_4602,N_4712);
nand U4940 (N_4940,N_4696,N_4778);
and U4941 (N_4941,N_4692,N_4743);
nor U4942 (N_4942,N_4640,N_4773);
nand U4943 (N_4943,N_4771,N_4737);
nand U4944 (N_4944,N_4728,N_4787);
xor U4945 (N_4945,N_4785,N_4712);
nand U4946 (N_4946,N_4619,N_4792);
xnor U4947 (N_4947,N_4634,N_4740);
xnor U4948 (N_4948,N_4645,N_4714);
and U4949 (N_4949,N_4750,N_4688);
xnor U4950 (N_4950,N_4762,N_4689);
or U4951 (N_4951,N_4622,N_4722);
nor U4952 (N_4952,N_4667,N_4669);
nor U4953 (N_4953,N_4612,N_4728);
nand U4954 (N_4954,N_4699,N_4775);
or U4955 (N_4955,N_4709,N_4666);
nand U4956 (N_4956,N_4663,N_4653);
xor U4957 (N_4957,N_4662,N_4751);
xor U4958 (N_4958,N_4782,N_4664);
or U4959 (N_4959,N_4709,N_4700);
nor U4960 (N_4960,N_4603,N_4636);
and U4961 (N_4961,N_4696,N_4612);
or U4962 (N_4962,N_4699,N_4604);
nand U4963 (N_4963,N_4705,N_4698);
or U4964 (N_4964,N_4644,N_4772);
or U4965 (N_4965,N_4777,N_4782);
nor U4966 (N_4966,N_4674,N_4748);
or U4967 (N_4967,N_4705,N_4792);
and U4968 (N_4968,N_4653,N_4751);
or U4969 (N_4969,N_4689,N_4619);
or U4970 (N_4970,N_4786,N_4654);
nor U4971 (N_4971,N_4708,N_4603);
nand U4972 (N_4972,N_4629,N_4765);
or U4973 (N_4973,N_4786,N_4766);
nor U4974 (N_4974,N_4746,N_4702);
and U4975 (N_4975,N_4648,N_4760);
and U4976 (N_4976,N_4693,N_4779);
xnor U4977 (N_4977,N_4794,N_4639);
xnor U4978 (N_4978,N_4690,N_4654);
nor U4979 (N_4979,N_4669,N_4602);
nand U4980 (N_4980,N_4740,N_4692);
or U4981 (N_4981,N_4702,N_4656);
nor U4982 (N_4982,N_4699,N_4760);
and U4983 (N_4983,N_4627,N_4774);
and U4984 (N_4984,N_4689,N_4739);
nor U4985 (N_4985,N_4642,N_4715);
and U4986 (N_4986,N_4766,N_4677);
or U4987 (N_4987,N_4646,N_4683);
nand U4988 (N_4988,N_4724,N_4638);
nand U4989 (N_4989,N_4702,N_4642);
and U4990 (N_4990,N_4676,N_4678);
nor U4991 (N_4991,N_4797,N_4752);
xnor U4992 (N_4992,N_4746,N_4731);
or U4993 (N_4993,N_4671,N_4694);
nand U4994 (N_4994,N_4609,N_4745);
nor U4995 (N_4995,N_4659,N_4743);
xor U4996 (N_4996,N_4719,N_4691);
and U4997 (N_4997,N_4692,N_4733);
and U4998 (N_4998,N_4791,N_4696);
and U4999 (N_4999,N_4681,N_4631);
or UO_0 (O_0,N_4995,N_4884);
xor UO_1 (O_1,N_4911,N_4861);
and UO_2 (O_2,N_4946,N_4821);
nand UO_3 (O_3,N_4889,N_4899);
nand UO_4 (O_4,N_4976,N_4970);
or UO_5 (O_5,N_4834,N_4837);
xnor UO_6 (O_6,N_4886,N_4986);
nand UO_7 (O_7,N_4982,N_4871);
nand UO_8 (O_8,N_4887,N_4981);
xor UO_9 (O_9,N_4967,N_4936);
and UO_10 (O_10,N_4851,N_4902);
or UO_11 (O_11,N_4932,N_4814);
and UO_12 (O_12,N_4848,N_4804);
nand UO_13 (O_13,N_4812,N_4874);
xnor UO_14 (O_14,N_4811,N_4964);
nand UO_15 (O_15,N_4987,N_4923);
and UO_16 (O_16,N_4898,N_4957);
nor UO_17 (O_17,N_4838,N_4979);
nand UO_18 (O_18,N_4990,N_4803);
or UO_19 (O_19,N_4845,N_4829);
and UO_20 (O_20,N_4996,N_4823);
or UO_21 (O_21,N_4989,N_4901);
nor UO_22 (O_22,N_4916,N_4891);
nor UO_23 (O_23,N_4855,N_4962);
and UO_24 (O_24,N_4840,N_4894);
or UO_25 (O_25,N_4992,N_4893);
nor UO_26 (O_26,N_4802,N_4817);
xor UO_27 (O_27,N_4949,N_4921);
nand UO_28 (O_28,N_4933,N_4961);
and UO_29 (O_29,N_4863,N_4953);
or UO_30 (O_30,N_4984,N_4930);
and UO_31 (O_31,N_4879,N_4927);
or UO_32 (O_32,N_4807,N_4928);
xnor UO_33 (O_33,N_4922,N_4931);
or UO_34 (O_34,N_4881,N_4983);
xnor UO_35 (O_35,N_4943,N_4913);
nor UO_36 (O_36,N_4935,N_4882);
nor UO_37 (O_37,N_4846,N_4939);
or UO_38 (O_38,N_4998,N_4854);
or UO_39 (O_39,N_4912,N_4900);
xnor UO_40 (O_40,N_4810,N_4828);
nor UO_41 (O_41,N_4905,N_4841);
nor UO_42 (O_42,N_4826,N_4824);
xnor UO_43 (O_43,N_4868,N_4806);
and UO_44 (O_44,N_4896,N_4819);
and UO_45 (O_45,N_4864,N_4867);
xnor UO_46 (O_46,N_4842,N_4937);
or UO_47 (O_47,N_4862,N_4951);
and UO_48 (O_48,N_4839,N_4909);
nor UO_49 (O_49,N_4994,N_4917);
nand UO_50 (O_50,N_4958,N_4952);
or UO_51 (O_51,N_4903,N_4849);
xor UO_52 (O_52,N_4800,N_4869);
xnor UO_53 (O_53,N_4836,N_4968);
nor UO_54 (O_54,N_4914,N_4908);
and UO_55 (O_55,N_4866,N_4915);
nand UO_56 (O_56,N_4934,N_4942);
xor UO_57 (O_57,N_4941,N_4830);
xnor UO_58 (O_58,N_4978,N_4897);
xnor UO_59 (O_59,N_4865,N_4926);
nor UO_60 (O_60,N_4929,N_4856);
nor UO_61 (O_61,N_4973,N_4993);
xor UO_62 (O_62,N_4910,N_4954);
nand UO_63 (O_63,N_4805,N_4924);
nand UO_64 (O_64,N_4873,N_4999);
or UO_65 (O_65,N_4940,N_4835);
and UO_66 (O_66,N_4831,N_4971);
nor UO_67 (O_67,N_4966,N_4820);
or UO_68 (O_68,N_4963,N_4904);
nor UO_69 (O_69,N_4991,N_4918);
or UO_70 (O_70,N_4997,N_4880);
or UO_71 (O_71,N_4956,N_4890);
nand UO_72 (O_72,N_4825,N_4833);
or UO_73 (O_73,N_4859,N_4948);
and UO_74 (O_74,N_4920,N_4895);
or UO_75 (O_75,N_4809,N_4843);
or UO_76 (O_76,N_4870,N_4985);
nor UO_77 (O_77,N_4944,N_4950);
and UO_78 (O_78,N_4969,N_4945);
and UO_79 (O_79,N_4876,N_4816);
and UO_80 (O_80,N_4974,N_4813);
and UO_81 (O_81,N_4850,N_4885);
xnor UO_82 (O_82,N_4906,N_4844);
xor UO_83 (O_83,N_4938,N_4877);
or UO_84 (O_84,N_4965,N_4822);
nor UO_85 (O_85,N_4925,N_4827);
xor UO_86 (O_86,N_4947,N_4980);
nor UO_87 (O_87,N_4972,N_4960);
xnor UO_88 (O_88,N_4815,N_4847);
nor UO_89 (O_89,N_4858,N_4808);
nand UO_90 (O_90,N_4878,N_4801);
and UO_91 (O_91,N_4857,N_4907);
xnor UO_92 (O_92,N_4872,N_4883);
and UO_93 (O_93,N_4919,N_4832);
nand UO_94 (O_94,N_4977,N_4875);
or UO_95 (O_95,N_4818,N_4959);
nor UO_96 (O_96,N_4852,N_4892);
nand UO_97 (O_97,N_4975,N_4955);
nor UO_98 (O_98,N_4888,N_4853);
and UO_99 (O_99,N_4988,N_4860);
and UO_100 (O_100,N_4995,N_4940);
nand UO_101 (O_101,N_4829,N_4918);
xnor UO_102 (O_102,N_4957,N_4817);
xnor UO_103 (O_103,N_4964,N_4859);
xor UO_104 (O_104,N_4845,N_4938);
nor UO_105 (O_105,N_4965,N_4994);
xor UO_106 (O_106,N_4864,N_4862);
and UO_107 (O_107,N_4843,N_4867);
and UO_108 (O_108,N_4971,N_4907);
nand UO_109 (O_109,N_4963,N_4978);
xor UO_110 (O_110,N_4903,N_4982);
nand UO_111 (O_111,N_4871,N_4930);
nor UO_112 (O_112,N_4824,N_4830);
nor UO_113 (O_113,N_4854,N_4866);
or UO_114 (O_114,N_4836,N_4820);
and UO_115 (O_115,N_4926,N_4991);
nand UO_116 (O_116,N_4845,N_4924);
nand UO_117 (O_117,N_4882,N_4994);
and UO_118 (O_118,N_4879,N_4978);
nor UO_119 (O_119,N_4973,N_4927);
xnor UO_120 (O_120,N_4937,N_4851);
or UO_121 (O_121,N_4987,N_4945);
and UO_122 (O_122,N_4919,N_4856);
and UO_123 (O_123,N_4885,N_4851);
xnor UO_124 (O_124,N_4815,N_4832);
nor UO_125 (O_125,N_4839,N_4814);
xor UO_126 (O_126,N_4958,N_4830);
nand UO_127 (O_127,N_4967,N_4832);
nand UO_128 (O_128,N_4956,N_4982);
xor UO_129 (O_129,N_4965,N_4920);
nand UO_130 (O_130,N_4873,N_4866);
nand UO_131 (O_131,N_4900,N_4949);
nor UO_132 (O_132,N_4948,N_4902);
nand UO_133 (O_133,N_4848,N_4962);
and UO_134 (O_134,N_4833,N_4939);
nor UO_135 (O_135,N_4918,N_4842);
and UO_136 (O_136,N_4901,N_4927);
or UO_137 (O_137,N_4868,N_4880);
nor UO_138 (O_138,N_4826,N_4957);
nor UO_139 (O_139,N_4819,N_4823);
nor UO_140 (O_140,N_4949,N_4834);
or UO_141 (O_141,N_4847,N_4802);
nor UO_142 (O_142,N_4848,N_4919);
nand UO_143 (O_143,N_4883,N_4897);
nand UO_144 (O_144,N_4955,N_4824);
nand UO_145 (O_145,N_4918,N_4960);
xnor UO_146 (O_146,N_4941,N_4978);
nand UO_147 (O_147,N_4867,N_4859);
xor UO_148 (O_148,N_4815,N_4920);
nand UO_149 (O_149,N_4912,N_4851);
and UO_150 (O_150,N_4910,N_4908);
nor UO_151 (O_151,N_4996,N_4947);
nand UO_152 (O_152,N_4946,N_4846);
and UO_153 (O_153,N_4864,N_4977);
xnor UO_154 (O_154,N_4872,N_4951);
nand UO_155 (O_155,N_4962,N_4900);
and UO_156 (O_156,N_4870,N_4975);
or UO_157 (O_157,N_4881,N_4902);
nand UO_158 (O_158,N_4837,N_4919);
nand UO_159 (O_159,N_4858,N_4973);
nand UO_160 (O_160,N_4840,N_4841);
and UO_161 (O_161,N_4867,N_4892);
and UO_162 (O_162,N_4820,N_4931);
and UO_163 (O_163,N_4942,N_4895);
and UO_164 (O_164,N_4975,N_4978);
and UO_165 (O_165,N_4922,N_4802);
or UO_166 (O_166,N_4901,N_4823);
and UO_167 (O_167,N_4915,N_4959);
nand UO_168 (O_168,N_4866,N_4919);
or UO_169 (O_169,N_4958,N_4872);
xnor UO_170 (O_170,N_4867,N_4905);
or UO_171 (O_171,N_4835,N_4823);
nor UO_172 (O_172,N_4868,N_4896);
or UO_173 (O_173,N_4863,N_4817);
and UO_174 (O_174,N_4937,N_4896);
nor UO_175 (O_175,N_4955,N_4834);
or UO_176 (O_176,N_4901,N_4945);
or UO_177 (O_177,N_4809,N_4935);
and UO_178 (O_178,N_4846,N_4816);
and UO_179 (O_179,N_4893,N_4873);
and UO_180 (O_180,N_4961,N_4851);
nand UO_181 (O_181,N_4911,N_4892);
xnor UO_182 (O_182,N_4897,N_4986);
nand UO_183 (O_183,N_4983,N_4828);
and UO_184 (O_184,N_4866,N_4926);
xnor UO_185 (O_185,N_4927,N_4947);
xor UO_186 (O_186,N_4865,N_4811);
nor UO_187 (O_187,N_4843,N_4847);
and UO_188 (O_188,N_4841,N_4975);
xor UO_189 (O_189,N_4802,N_4929);
or UO_190 (O_190,N_4922,N_4813);
nand UO_191 (O_191,N_4887,N_4846);
nand UO_192 (O_192,N_4880,N_4952);
and UO_193 (O_193,N_4945,N_4893);
or UO_194 (O_194,N_4873,N_4969);
or UO_195 (O_195,N_4951,N_4981);
xor UO_196 (O_196,N_4868,N_4878);
and UO_197 (O_197,N_4837,N_4949);
xnor UO_198 (O_198,N_4850,N_4950);
or UO_199 (O_199,N_4866,N_4813);
nand UO_200 (O_200,N_4971,N_4810);
or UO_201 (O_201,N_4966,N_4935);
or UO_202 (O_202,N_4963,N_4821);
xor UO_203 (O_203,N_4949,N_4944);
nor UO_204 (O_204,N_4995,N_4988);
and UO_205 (O_205,N_4940,N_4985);
nand UO_206 (O_206,N_4939,N_4999);
nor UO_207 (O_207,N_4890,N_4866);
nand UO_208 (O_208,N_4812,N_4897);
xor UO_209 (O_209,N_4907,N_4982);
nand UO_210 (O_210,N_4987,N_4846);
or UO_211 (O_211,N_4983,N_4937);
xnor UO_212 (O_212,N_4822,N_4805);
xor UO_213 (O_213,N_4806,N_4894);
nand UO_214 (O_214,N_4869,N_4957);
xor UO_215 (O_215,N_4828,N_4985);
and UO_216 (O_216,N_4979,N_4822);
xnor UO_217 (O_217,N_4866,N_4845);
and UO_218 (O_218,N_4937,N_4859);
and UO_219 (O_219,N_4855,N_4868);
and UO_220 (O_220,N_4954,N_4933);
and UO_221 (O_221,N_4968,N_4808);
nand UO_222 (O_222,N_4883,N_4807);
and UO_223 (O_223,N_4855,N_4937);
nor UO_224 (O_224,N_4957,N_4814);
nand UO_225 (O_225,N_4928,N_4937);
and UO_226 (O_226,N_4943,N_4915);
nor UO_227 (O_227,N_4965,N_4866);
nor UO_228 (O_228,N_4997,N_4905);
and UO_229 (O_229,N_4956,N_4870);
or UO_230 (O_230,N_4867,N_4906);
nand UO_231 (O_231,N_4950,N_4996);
and UO_232 (O_232,N_4943,N_4887);
nand UO_233 (O_233,N_4925,N_4844);
and UO_234 (O_234,N_4827,N_4880);
nand UO_235 (O_235,N_4813,N_4937);
nor UO_236 (O_236,N_4874,N_4805);
and UO_237 (O_237,N_4909,N_4885);
and UO_238 (O_238,N_4828,N_4974);
nand UO_239 (O_239,N_4837,N_4870);
or UO_240 (O_240,N_4999,N_4877);
nand UO_241 (O_241,N_4974,N_4994);
xor UO_242 (O_242,N_4997,N_4942);
nor UO_243 (O_243,N_4828,N_4862);
or UO_244 (O_244,N_4805,N_4807);
or UO_245 (O_245,N_4993,N_4807);
and UO_246 (O_246,N_4873,N_4880);
and UO_247 (O_247,N_4901,N_4957);
nor UO_248 (O_248,N_4995,N_4857);
nor UO_249 (O_249,N_4947,N_4802);
and UO_250 (O_250,N_4974,N_4993);
nor UO_251 (O_251,N_4847,N_4804);
and UO_252 (O_252,N_4935,N_4926);
xnor UO_253 (O_253,N_4975,N_4871);
nand UO_254 (O_254,N_4926,N_4956);
xor UO_255 (O_255,N_4849,N_4831);
nor UO_256 (O_256,N_4906,N_4971);
xor UO_257 (O_257,N_4909,N_4893);
xor UO_258 (O_258,N_4855,N_4934);
nor UO_259 (O_259,N_4919,N_4807);
nor UO_260 (O_260,N_4837,N_4945);
xnor UO_261 (O_261,N_4970,N_4887);
nand UO_262 (O_262,N_4935,N_4829);
xnor UO_263 (O_263,N_4988,N_4938);
and UO_264 (O_264,N_4824,N_4920);
nor UO_265 (O_265,N_4998,N_4990);
xnor UO_266 (O_266,N_4834,N_4972);
nor UO_267 (O_267,N_4966,N_4830);
or UO_268 (O_268,N_4998,N_4841);
nor UO_269 (O_269,N_4825,N_4832);
and UO_270 (O_270,N_4804,N_4879);
and UO_271 (O_271,N_4924,N_4946);
or UO_272 (O_272,N_4965,N_4829);
or UO_273 (O_273,N_4996,N_4891);
xnor UO_274 (O_274,N_4843,N_4962);
xor UO_275 (O_275,N_4864,N_4846);
or UO_276 (O_276,N_4846,N_4882);
nand UO_277 (O_277,N_4957,N_4871);
nand UO_278 (O_278,N_4970,N_4981);
and UO_279 (O_279,N_4846,N_4940);
and UO_280 (O_280,N_4984,N_4803);
nor UO_281 (O_281,N_4813,N_4848);
or UO_282 (O_282,N_4892,N_4912);
xnor UO_283 (O_283,N_4894,N_4850);
nand UO_284 (O_284,N_4805,N_4945);
and UO_285 (O_285,N_4991,N_4892);
xor UO_286 (O_286,N_4868,N_4850);
nor UO_287 (O_287,N_4857,N_4820);
nand UO_288 (O_288,N_4979,N_4929);
nor UO_289 (O_289,N_4980,N_4935);
or UO_290 (O_290,N_4990,N_4865);
xor UO_291 (O_291,N_4852,N_4890);
or UO_292 (O_292,N_4825,N_4997);
xor UO_293 (O_293,N_4922,N_4911);
nand UO_294 (O_294,N_4910,N_4962);
and UO_295 (O_295,N_4946,N_4866);
nor UO_296 (O_296,N_4830,N_4901);
xor UO_297 (O_297,N_4963,N_4827);
xnor UO_298 (O_298,N_4805,N_4845);
nand UO_299 (O_299,N_4836,N_4800);
nand UO_300 (O_300,N_4813,N_4909);
and UO_301 (O_301,N_4844,N_4950);
nand UO_302 (O_302,N_4906,N_4967);
xor UO_303 (O_303,N_4997,N_4962);
or UO_304 (O_304,N_4842,N_4925);
and UO_305 (O_305,N_4939,N_4876);
or UO_306 (O_306,N_4811,N_4882);
and UO_307 (O_307,N_4808,N_4876);
nor UO_308 (O_308,N_4816,N_4946);
or UO_309 (O_309,N_4913,N_4890);
and UO_310 (O_310,N_4834,N_4909);
nand UO_311 (O_311,N_4900,N_4905);
and UO_312 (O_312,N_4952,N_4973);
or UO_313 (O_313,N_4979,N_4882);
nand UO_314 (O_314,N_4993,N_4866);
and UO_315 (O_315,N_4873,N_4972);
or UO_316 (O_316,N_4832,N_4941);
xor UO_317 (O_317,N_4963,N_4822);
xnor UO_318 (O_318,N_4936,N_4973);
or UO_319 (O_319,N_4943,N_4850);
or UO_320 (O_320,N_4841,N_4807);
and UO_321 (O_321,N_4972,N_4901);
nor UO_322 (O_322,N_4924,N_4838);
or UO_323 (O_323,N_4902,N_4991);
nand UO_324 (O_324,N_4923,N_4812);
nor UO_325 (O_325,N_4851,N_4978);
nand UO_326 (O_326,N_4913,N_4850);
nor UO_327 (O_327,N_4870,N_4800);
nand UO_328 (O_328,N_4909,N_4874);
xnor UO_329 (O_329,N_4949,N_4909);
and UO_330 (O_330,N_4927,N_4990);
or UO_331 (O_331,N_4951,N_4860);
nand UO_332 (O_332,N_4994,N_4827);
nor UO_333 (O_333,N_4847,N_4977);
and UO_334 (O_334,N_4988,N_4947);
or UO_335 (O_335,N_4816,N_4804);
or UO_336 (O_336,N_4860,N_4804);
xor UO_337 (O_337,N_4959,N_4999);
nor UO_338 (O_338,N_4811,N_4908);
xnor UO_339 (O_339,N_4828,N_4942);
and UO_340 (O_340,N_4808,N_4880);
or UO_341 (O_341,N_4968,N_4875);
nor UO_342 (O_342,N_4916,N_4963);
and UO_343 (O_343,N_4899,N_4932);
nand UO_344 (O_344,N_4824,N_4839);
or UO_345 (O_345,N_4885,N_4973);
or UO_346 (O_346,N_4975,N_4825);
xor UO_347 (O_347,N_4956,N_4869);
or UO_348 (O_348,N_4908,N_4820);
or UO_349 (O_349,N_4996,N_4839);
or UO_350 (O_350,N_4914,N_4980);
and UO_351 (O_351,N_4948,N_4894);
nor UO_352 (O_352,N_4979,N_4875);
nand UO_353 (O_353,N_4981,N_4832);
xnor UO_354 (O_354,N_4835,N_4876);
nand UO_355 (O_355,N_4829,N_4813);
nand UO_356 (O_356,N_4806,N_4982);
nor UO_357 (O_357,N_4830,N_4864);
and UO_358 (O_358,N_4970,N_4895);
nor UO_359 (O_359,N_4985,N_4871);
or UO_360 (O_360,N_4976,N_4972);
nor UO_361 (O_361,N_4943,N_4974);
and UO_362 (O_362,N_4964,N_4979);
and UO_363 (O_363,N_4818,N_4846);
nor UO_364 (O_364,N_4933,N_4859);
nand UO_365 (O_365,N_4890,N_4896);
and UO_366 (O_366,N_4863,N_4845);
or UO_367 (O_367,N_4983,N_4879);
or UO_368 (O_368,N_4982,N_4969);
nand UO_369 (O_369,N_4929,N_4962);
and UO_370 (O_370,N_4814,N_4802);
and UO_371 (O_371,N_4934,N_4859);
nand UO_372 (O_372,N_4821,N_4961);
and UO_373 (O_373,N_4805,N_4802);
or UO_374 (O_374,N_4902,N_4963);
nor UO_375 (O_375,N_4950,N_4909);
nor UO_376 (O_376,N_4874,N_4857);
nor UO_377 (O_377,N_4873,N_4965);
and UO_378 (O_378,N_4952,N_4886);
xor UO_379 (O_379,N_4807,N_4934);
and UO_380 (O_380,N_4976,N_4910);
and UO_381 (O_381,N_4940,N_4880);
nor UO_382 (O_382,N_4831,N_4998);
and UO_383 (O_383,N_4971,N_4801);
nor UO_384 (O_384,N_4871,N_4825);
nand UO_385 (O_385,N_4950,N_4994);
nor UO_386 (O_386,N_4853,N_4903);
xor UO_387 (O_387,N_4858,N_4910);
or UO_388 (O_388,N_4808,N_4944);
nor UO_389 (O_389,N_4900,N_4827);
or UO_390 (O_390,N_4937,N_4877);
xor UO_391 (O_391,N_4937,N_4805);
xor UO_392 (O_392,N_4808,N_4888);
or UO_393 (O_393,N_4944,N_4846);
or UO_394 (O_394,N_4909,N_4916);
xnor UO_395 (O_395,N_4818,N_4996);
nand UO_396 (O_396,N_4988,N_4851);
nand UO_397 (O_397,N_4800,N_4827);
xnor UO_398 (O_398,N_4895,N_4906);
xor UO_399 (O_399,N_4906,N_4957);
or UO_400 (O_400,N_4892,N_4812);
and UO_401 (O_401,N_4899,N_4861);
or UO_402 (O_402,N_4860,N_4898);
and UO_403 (O_403,N_4997,N_4887);
nand UO_404 (O_404,N_4941,N_4880);
nor UO_405 (O_405,N_4953,N_4873);
xnor UO_406 (O_406,N_4879,N_4972);
and UO_407 (O_407,N_4824,N_4903);
or UO_408 (O_408,N_4877,N_4837);
nor UO_409 (O_409,N_4888,N_4891);
nor UO_410 (O_410,N_4865,N_4941);
nor UO_411 (O_411,N_4941,N_4859);
xnor UO_412 (O_412,N_4925,N_4835);
and UO_413 (O_413,N_4946,N_4883);
xnor UO_414 (O_414,N_4959,N_4939);
or UO_415 (O_415,N_4977,N_4820);
or UO_416 (O_416,N_4869,N_4858);
and UO_417 (O_417,N_4858,N_4855);
nor UO_418 (O_418,N_4996,N_4857);
or UO_419 (O_419,N_4996,N_4805);
nand UO_420 (O_420,N_4935,N_4937);
nand UO_421 (O_421,N_4848,N_4937);
xnor UO_422 (O_422,N_4980,N_4901);
xor UO_423 (O_423,N_4882,N_4891);
or UO_424 (O_424,N_4970,N_4829);
or UO_425 (O_425,N_4984,N_4978);
nor UO_426 (O_426,N_4878,N_4889);
or UO_427 (O_427,N_4879,N_4962);
and UO_428 (O_428,N_4959,N_4821);
xor UO_429 (O_429,N_4919,N_4863);
and UO_430 (O_430,N_4869,N_4829);
or UO_431 (O_431,N_4835,N_4932);
and UO_432 (O_432,N_4994,N_4806);
nand UO_433 (O_433,N_4863,N_4866);
or UO_434 (O_434,N_4997,N_4957);
xor UO_435 (O_435,N_4905,N_4842);
nand UO_436 (O_436,N_4894,N_4975);
nor UO_437 (O_437,N_4931,N_4954);
or UO_438 (O_438,N_4842,N_4840);
nand UO_439 (O_439,N_4835,N_4999);
nand UO_440 (O_440,N_4882,N_4934);
nand UO_441 (O_441,N_4997,N_4981);
and UO_442 (O_442,N_4926,N_4863);
nor UO_443 (O_443,N_4849,N_4971);
xor UO_444 (O_444,N_4841,N_4960);
or UO_445 (O_445,N_4939,N_4980);
nand UO_446 (O_446,N_4977,N_4949);
nand UO_447 (O_447,N_4872,N_4977);
nand UO_448 (O_448,N_4938,N_4953);
or UO_449 (O_449,N_4994,N_4914);
or UO_450 (O_450,N_4883,N_4949);
xor UO_451 (O_451,N_4840,N_4814);
or UO_452 (O_452,N_4929,N_4967);
and UO_453 (O_453,N_4864,N_4890);
or UO_454 (O_454,N_4898,N_4997);
or UO_455 (O_455,N_4862,N_4853);
nor UO_456 (O_456,N_4853,N_4925);
nand UO_457 (O_457,N_4981,N_4826);
nor UO_458 (O_458,N_4930,N_4939);
nor UO_459 (O_459,N_4888,N_4868);
and UO_460 (O_460,N_4873,N_4979);
or UO_461 (O_461,N_4977,N_4981);
or UO_462 (O_462,N_4834,N_4950);
xor UO_463 (O_463,N_4815,N_4925);
or UO_464 (O_464,N_4804,N_4978);
xor UO_465 (O_465,N_4826,N_4972);
or UO_466 (O_466,N_4819,N_4975);
or UO_467 (O_467,N_4819,N_4828);
and UO_468 (O_468,N_4820,N_4933);
or UO_469 (O_469,N_4982,N_4924);
or UO_470 (O_470,N_4964,N_4996);
and UO_471 (O_471,N_4957,N_4887);
xor UO_472 (O_472,N_4971,N_4982);
or UO_473 (O_473,N_4992,N_4990);
nand UO_474 (O_474,N_4975,N_4812);
and UO_475 (O_475,N_4871,N_4880);
xnor UO_476 (O_476,N_4972,N_4954);
and UO_477 (O_477,N_4941,N_4814);
xor UO_478 (O_478,N_4991,N_4980);
nand UO_479 (O_479,N_4912,N_4807);
nand UO_480 (O_480,N_4885,N_4916);
xor UO_481 (O_481,N_4898,N_4830);
nor UO_482 (O_482,N_4843,N_4972);
xor UO_483 (O_483,N_4988,N_4859);
nor UO_484 (O_484,N_4846,N_4898);
xor UO_485 (O_485,N_4869,N_4983);
or UO_486 (O_486,N_4808,N_4919);
nor UO_487 (O_487,N_4828,N_4878);
nand UO_488 (O_488,N_4989,N_4859);
nor UO_489 (O_489,N_4862,N_4841);
xnor UO_490 (O_490,N_4840,N_4998);
and UO_491 (O_491,N_4942,N_4970);
xor UO_492 (O_492,N_4982,N_4823);
or UO_493 (O_493,N_4839,N_4826);
xor UO_494 (O_494,N_4859,N_4806);
or UO_495 (O_495,N_4953,N_4817);
xor UO_496 (O_496,N_4871,N_4912);
nor UO_497 (O_497,N_4801,N_4814);
xor UO_498 (O_498,N_4887,N_4903);
and UO_499 (O_499,N_4962,N_4986);
and UO_500 (O_500,N_4921,N_4835);
xnor UO_501 (O_501,N_4879,N_4905);
or UO_502 (O_502,N_4853,N_4932);
nand UO_503 (O_503,N_4846,N_4999);
nor UO_504 (O_504,N_4864,N_4857);
xnor UO_505 (O_505,N_4856,N_4975);
nor UO_506 (O_506,N_4874,N_4878);
and UO_507 (O_507,N_4908,N_4866);
and UO_508 (O_508,N_4857,N_4908);
xor UO_509 (O_509,N_4841,N_4895);
nor UO_510 (O_510,N_4849,N_4821);
nor UO_511 (O_511,N_4947,N_4839);
or UO_512 (O_512,N_4958,N_4827);
and UO_513 (O_513,N_4837,N_4942);
xnor UO_514 (O_514,N_4810,N_4916);
nor UO_515 (O_515,N_4825,N_4889);
nand UO_516 (O_516,N_4832,N_4957);
and UO_517 (O_517,N_4950,N_4885);
nand UO_518 (O_518,N_4853,N_4842);
xnor UO_519 (O_519,N_4810,N_4857);
or UO_520 (O_520,N_4981,N_4810);
or UO_521 (O_521,N_4942,N_4989);
and UO_522 (O_522,N_4827,N_4897);
nand UO_523 (O_523,N_4892,N_4833);
nand UO_524 (O_524,N_4908,N_4846);
or UO_525 (O_525,N_4831,N_4904);
and UO_526 (O_526,N_4982,N_4857);
and UO_527 (O_527,N_4816,N_4812);
nor UO_528 (O_528,N_4861,N_4933);
or UO_529 (O_529,N_4928,N_4999);
nor UO_530 (O_530,N_4906,N_4911);
nor UO_531 (O_531,N_4809,N_4997);
nand UO_532 (O_532,N_4980,N_4973);
nor UO_533 (O_533,N_4859,N_4946);
nand UO_534 (O_534,N_4989,N_4881);
and UO_535 (O_535,N_4898,N_4856);
nand UO_536 (O_536,N_4911,N_4977);
or UO_537 (O_537,N_4823,N_4879);
nor UO_538 (O_538,N_4925,N_4850);
and UO_539 (O_539,N_4948,N_4975);
nor UO_540 (O_540,N_4971,N_4924);
or UO_541 (O_541,N_4988,N_4997);
nor UO_542 (O_542,N_4924,N_4855);
or UO_543 (O_543,N_4906,N_4803);
xor UO_544 (O_544,N_4993,N_4816);
or UO_545 (O_545,N_4858,N_4975);
and UO_546 (O_546,N_4828,N_4906);
and UO_547 (O_547,N_4995,N_4898);
nand UO_548 (O_548,N_4996,N_4949);
nand UO_549 (O_549,N_4810,N_4826);
or UO_550 (O_550,N_4861,N_4922);
or UO_551 (O_551,N_4890,N_4941);
and UO_552 (O_552,N_4942,N_4871);
nor UO_553 (O_553,N_4845,N_4943);
and UO_554 (O_554,N_4916,N_4946);
or UO_555 (O_555,N_4995,N_4852);
and UO_556 (O_556,N_4890,N_4977);
or UO_557 (O_557,N_4832,N_4968);
nand UO_558 (O_558,N_4961,N_4928);
nand UO_559 (O_559,N_4826,N_4945);
xnor UO_560 (O_560,N_4832,N_4977);
nand UO_561 (O_561,N_4886,N_4978);
nand UO_562 (O_562,N_4941,N_4838);
and UO_563 (O_563,N_4864,N_4925);
xor UO_564 (O_564,N_4955,N_4948);
xnor UO_565 (O_565,N_4968,N_4920);
xor UO_566 (O_566,N_4850,N_4999);
xnor UO_567 (O_567,N_4858,N_4955);
and UO_568 (O_568,N_4859,N_4871);
or UO_569 (O_569,N_4912,N_4815);
and UO_570 (O_570,N_4908,N_4806);
or UO_571 (O_571,N_4869,N_4945);
or UO_572 (O_572,N_4822,N_4854);
or UO_573 (O_573,N_4806,N_4916);
nand UO_574 (O_574,N_4803,N_4853);
nor UO_575 (O_575,N_4928,N_4874);
and UO_576 (O_576,N_4969,N_4965);
nand UO_577 (O_577,N_4960,N_4824);
or UO_578 (O_578,N_4918,N_4911);
nand UO_579 (O_579,N_4869,N_4843);
nand UO_580 (O_580,N_4820,N_4915);
or UO_581 (O_581,N_4874,N_4975);
and UO_582 (O_582,N_4801,N_4804);
and UO_583 (O_583,N_4993,N_4834);
nand UO_584 (O_584,N_4897,N_4834);
or UO_585 (O_585,N_4958,N_4826);
nor UO_586 (O_586,N_4986,N_4807);
or UO_587 (O_587,N_4834,N_4985);
and UO_588 (O_588,N_4993,N_4831);
nor UO_589 (O_589,N_4951,N_4913);
xnor UO_590 (O_590,N_4864,N_4807);
and UO_591 (O_591,N_4873,N_4853);
nand UO_592 (O_592,N_4907,N_4859);
or UO_593 (O_593,N_4874,N_4883);
and UO_594 (O_594,N_4894,N_4922);
nor UO_595 (O_595,N_4890,N_4927);
or UO_596 (O_596,N_4850,N_4896);
nand UO_597 (O_597,N_4966,N_4898);
nor UO_598 (O_598,N_4880,N_4803);
xor UO_599 (O_599,N_4822,N_4829);
nand UO_600 (O_600,N_4887,N_4969);
xor UO_601 (O_601,N_4999,N_4946);
and UO_602 (O_602,N_4971,N_4871);
xnor UO_603 (O_603,N_4943,N_4872);
xnor UO_604 (O_604,N_4901,N_4964);
nand UO_605 (O_605,N_4889,N_4981);
or UO_606 (O_606,N_4856,N_4909);
xor UO_607 (O_607,N_4870,N_4980);
nand UO_608 (O_608,N_4850,N_4878);
or UO_609 (O_609,N_4906,N_4936);
and UO_610 (O_610,N_4862,N_4950);
xor UO_611 (O_611,N_4999,N_4987);
nor UO_612 (O_612,N_4814,N_4978);
or UO_613 (O_613,N_4866,N_4977);
and UO_614 (O_614,N_4873,N_4948);
nor UO_615 (O_615,N_4812,N_4899);
nor UO_616 (O_616,N_4825,N_4952);
nor UO_617 (O_617,N_4948,N_4881);
nand UO_618 (O_618,N_4927,N_4889);
nor UO_619 (O_619,N_4952,N_4921);
or UO_620 (O_620,N_4903,N_4947);
nand UO_621 (O_621,N_4832,N_4899);
and UO_622 (O_622,N_4947,N_4818);
xor UO_623 (O_623,N_4850,N_4869);
xor UO_624 (O_624,N_4914,N_4843);
nor UO_625 (O_625,N_4847,N_4931);
nor UO_626 (O_626,N_4887,N_4835);
and UO_627 (O_627,N_4808,N_4906);
nor UO_628 (O_628,N_4835,N_4941);
nor UO_629 (O_629,N_4908,N_4812);
or UO_630 (O_630,N_4849,N_4894);
xor UO_631 (O_631,N_4818,N_4977);
and UO_632 (O_632,N_4932,N_4868);
nor UO_633 (O_633,N_4910,N_4937);
or UO_634 (O_634,N_4958,N_4945);
or UO_635 (O_635,N_4953,N_4840);
and UO_636 (O_636,N_4845,N_4998);
nor UO_637 (O_637,N_4859,N_4848);
xnor UO_638 (O_638,N_4817,N_4962);
or UO_639 (O_639,N_4802,N_4918);
xnor UO_640 (O_640,N_4986,N_4854);
and UO_641 (O_641,N_4950,N_4816);
or UO_642 (O_642,N_4944,N_4997);
nor UO_643 (O_643,N_4970,N_4860);
or UO_644 (O_644,N_4955,N_4973);
or UO_645 (O_645,N_4870,N_4970);
nor UO_646 (O_646,N_4876,N_4994);
nand UO_647 (O_647,N_4908,N_4950);
or UO_648 (O_648,N_4981,N_4805);
and UO_649 (O_649,N_4875,N_4996);
xor UO_650 (O_650,N_4829,N_4806);
xor UO_651 (O_651,N_4847,N_4919);
xnor UO_652 (O_652,N_4957,N_4842);
or UO_653 (O_653,N_4812,N_4865);
or UO_654 (O_654,N_4947,N_4933);
nor UO_655 (O_655,N_4957,N_4928);
nand UO_656 (O_656,N_4943,N_4823);
nand UO_657 (O_657,N_4884,N_4873);
and UO_658 (O_658,N_4831,N_4910);
nand UO_659 (O_659,N_4973,N_4944);
and UO_660 (O_660,N_4921,N_4962);
nor UO_661 (O_661,N_4848,N_4918);
or UO_662 (O_662,N_4846,N_4894);
xnor UO_663 (O_663,N_4949,N_4906);
xnor UO_664 (O_664,N_4963,N_4847);
nor UO_665 (O_665,N_4802,N_4867);
nand UO_666 (O_666,N_4973,N_4910);
or UO_667 (O_667,N_4953,N_4978);
nand UO_668 (O_668,N_4810,N_4995);
xnor UO_669 (O_669,N_4963,N_4900);
or UO_670 (O_670,N_4933,N_4969);
xnor UO_671 (O_671,N_4856,N_4901);
nand UO_672 (O_672,N_4804,N_4827);
xor UO_673 (O_673,N_4882,N_4838);
nor UO_674 (O_674,N_4910,N_4872);
nand UO_675 (O_675,N_4973,N_4982);
nand UO_676 (O_676,N_4875,N_4904);
nor UO_677 (O_677,N_4987,N_4924);
xor UO_678 (O_678,N_4949,N_4879);
or UO_679 (O_679,N_4828,N_4984);
nand UO_680 (O_680,N_4804,N_4909);
xor UO_681 (O_681,N_4900,N_4923);
or UO_682 (O_682,N_4958,N_4808);
or UO_683 (O_683,N_4841,N_4843);
and UO_684 (O_684,N_4868,N_4978);
and UO_685 (O_685,N_4814,N_4982);
or UO_686 (O_686,N_4823,N_4867);
nor UO_687 (O_687,N_4985,N_4991);
or UO_688 (O_688,N_4861,N_4830);
and UO_689 (O_689,N_4967,N_4961);
xnor UO_690 (O_690,N_4926,N_4815);
xor UO_691 (O_691,N_4893,N_4864);
xor UO_692 (O_692,N_4875,N_4956);
nand UO_693 (O_693,N_4999,N_4880);
or UO_694 (O_694,N_4838,N_4828);
or UO_695 (O_695,N_4915,N_4913);
or UO_696 (O_696,N_4861,N_4904);
or UO_697 (O_697,N_4884,N_4993);
nor UO_698 (O_698,N_4907,N_4827);
or UO_699 (O_699,N_4864,N_4879);
xor UO_700 (O_700,N_4843,N_4923);
nor UO_701 (O_701,N_4874,N_4868);
and UO_702 (O_702,N_4886,N_4933);
or UO_703 (O_703,N_4837,N_4892);
xnor UO_704 (O_704,N_4939,N_4977);
nand UO_705 (O_705,N_4929,N_4904);
xnor UO_706 (O_706,N_4802,N_4860);
and UO_707 (O_707,N_4892,N_4862);
xor UO_708 (O_708,N_4976,N_4832);
xnor UO_709 (O_709,N_4975,N_4846);
xor UO_710 (O_710,N_4944,N_4886);
or UO_711 (O_711,N_4883,N_4973);
xor UO_712 (O_712,N_4934,N_4992);
nand UO_713 (O_713,N_4955,N_4906);
nand UO_714 (O_714,N_4890,N_4867);
nor UO_715 (O_715,N_4877,N_4919);
and UO_716 (O_716,N_4946,N_4815);
or UO_717 (O_717,N_4921,N_4936);
and UO_718 (O_718,N_4984,N_4820);
and UO_719 (O_719,N_4982,N_4889);
xor UO_720 (O_720,N_4847,N_4909);
or UO_721 (O_721,N_4820,N_4863);
nand UO_722 (O_722,N_4827,N_4860);
and UO_723 (O_723,N_4946,N_4902);
and UO_724 (O_724,N_4903,N_4949);
nor UO_725 (O_725,N_4940,N_4939);
xnor UO_726 (O_726,N_4806,N_4938);
xor UO_727 (O_727,N_4830,N_4836);
nor UO_728 (O_728,N_4806,N_4931);
nand UO_729 (O_729,N_4884,N_4834);
nor UO_730 (O_730,N_4821,N_4902);
and UO_731 (O_731,N_4832,N_4876);
nor UO_732 (O_732,N_4991,N_4958);
and UO_733 (O_733,N_4995,N_4985);
or UO_734 (O_734,N_4814,N_4879);
and UO_735 (O_735,N_4804,N_4865);
nand UO_736 (O_736,N_4924,N_4864);
and UO_737 (O_737,N_4976,N_4887);
nand UO_738 (O_738,N_4980,N_4894);
nor UO_739 (O_739,N_4982,N_4878);
or UO_740 (O_740,N_4951,N_4810);
nand UO_741 (O_741,N_4971,N_4932);
nand UO_742 (O_742,N_4814,N_4885);
and UO_743 (O_743,N_4869,N_4919);
nand UO_744 (O_744,N_4897,N_4874);
or UO_745 (O_745,N_4918,N_4898);
nor UO_746 (O_746,N_4836,N_4909);
nor UO_747 (O_747,N_4978,N_4912);
nor UO_748 (O_748,N_4971,N_4927);
or UO_749 (O_749,N_4982,N_4994);
nor UO_750 (O_750,N_4992,N_4836);
or UO_751 (O_751,N_4947,N_4832);
and UO_752 (O_752,N_4892,N_4893);
xnor UO_753 (O_753,N_4829,N_4886);
xnor UO_754 (O_754,N_4969,N_4994);
and UO_755 (O_755,N_4983,N_4866);
nand UO_756 (O_756,N_4951,N_4953);
xor UO_757 (O_757,N_4918,N_4966);
or UO_758 (O_758,N_4872,N_4871);
xor UO_759 (O_759,N_4907,N_4970);
xnor UO_760 (O_760,N_4872,N_4815);
and UO_761 (O_761,N_4862,N_4876);
and UO_762 (O_762,N_4834,N_4851);
nor UO_763 (O_763,N_4973,N_4960);
nand UO_764 (O_764,N_4893,N_4951);
or UO_765 (O_765,N_4836,N_4940);
nor UO_766 (O_766,N_4886,N_4879);
or UO_767 (O_767,N_4949,N_4859);
nand UO_768 (O_768,N_4860,N_4896);
xnor UO_769 (O_769,N_4991,N_4940);
xor UO_770 (O_770,N_4852,N_4915);
nand UO_771 (O_771,N_4945,N_4991);
nand UO_772 (O_772,N_4819,N_4953);
and UO_773 (O_773,N_4984,N_4931);
nand UO_774 (O_774,N_4848,N_4856);
nor UO_775 (O_775,N_4896,N_4905);
nand UO_776 (O_776,N_4918,N_4833);
nand UO_777 (O_777,N_4933,N_4846);
xnor UO_778 (O_778,N_4890,N_4938);
and UO_779 (O_779,N_4912,N_4986);
nand UO_780 (O_780,N_4985,N_4964);
or UO_781 (O_781,N_4907,N_4960);
and UO_782 (O_782,N_4957,N_4890);
and UO_783 (O_783,N_4876,N_4888);
or UO_784 (O_784,N_4956,N_4900);
nand UO_785 (O_785,N_4934,N_4878);
nor UO_786 (O_786,N_4886,N_4884);
xnor UO_787 (O_787,N_4973,N_4979);
and UO_788 (O_788,N_4844,N_4891);
or UO_789 (O_789,N_4860,N_4906);
nor UO_790 (O_790,N_4837,N_4887);
nor UO_791 (O_791,N_4802,N_4897);
xor UO_792 (O_792,N_4903,N_4921);
xnor UO_793 (O_793,N_4905,N_4814);
nand UO_794 (O_794,N_4915,N_4833);
nand UO_795 (O_795,N_4885,N_4913);
and UO_796 (O_796,N_4835,N_4962);
nor UO_797 (O_797,N_4947,N_4975);
nor UO_798 (O_798,N_4927,N_4922);
xnor UO_799 (O_799,N_4847,N_4959);
nor UO_800 (O_800,N_4860,N_4820);
and UO_801 (O_801,N_4925,N_4965);
or UO_802 (O_802,N_4864,N_4901);
xor UO_803 (O_803,N_4988,N_4952);
nor UO_804 (O_804,N_4987,N_4891);
and UO_805 (O_805,N_4951,N_4868);
nand UO_806 (O_806,N_4998,N_4957);
or UO_807 (O_807,N_4904,N_4808);
nor UO_808 (O_808,N_4903,N_4873);
xnor UO_809 (O_809,N_4801,N_4864);
nand UO_810 (O_810,N_4825,N_4996);
xor UO_811 (O_811,N_4998,N_4842);
or UO_812 (O_812,N_4850,N_4930);
or UO_813 (O_813,N_4918,N_4807);
or UO_814 (O_814,N_4953,N_4976);
nand UO_815 (O_815,N_4902,N_4880);
xor UO_816 (O_816,N_4896,N_4932);
and UO_817 (O_817,N_4920,N_4927);
nand UO_818 (O_818,N_4897,N_4830);
nor UO_819 (O_819,N_4810,N_4978);
or UO_820 (O_820,N_4808,N_4861);
nor UO_821 (O_821,N_4993,N_4830);
and UO_822 (O_822,N_4870,N_4853);
and UO_823 (O_823,N_4943,N_4820);
nor UO_824 (O_824,N_4994,N_4861);
or UO_825 (O_825,N_4941,N_4827);
nand UO_826 (O_826,N_4967,N_4838);
and UO_827 (O_827,N_4948,N_4939);
nand UO_828 (O_828,N_4936,N_4871);
or UO_829 (O_829,N_4806,N_4996);
nand UO_830 (O_830,N_4983,N_4816);
nand UO_831 (O_831,N_4823,N_4989);
nand UO_832 (O_832,N_4900,N_4883);
or UO_833 (O_833,N_4925,N_4803);
nand UO_834 (O_834,N_4825,N_4801);
xnor UO_835 (O_835,N_4848,N_4898);
and UO_836 (O_836,N_4992,N_4919);
and UO_837 (O_837,N_4990,N_4908);
or UO_838 (O_838,N_4838,N_4833);
nand UO_839 (O_839,N_4828,N_4808);
and UO_840 (O_840,N_4985,N_4906);
or UO_841 (O_841,N_4855,N_4990);
and UO_842 (O_842,N_4858,N_4842);
xnor UO_843 (O_843,N_4808,N_4800);
nor UO_844 (O_844,N_4904,N_4915);
nand UO_845 (O_845,N_4818,N_4998);
nor UO_846 (O_846,N_4899,N_4980);
nand UO_847 (O_847,N_4815,N_4854);
nand UO_848 (O_848,N_4897,N_4832);
nand UO_849 (O_849,N_4947,N_4897);
and UO_850 (O_850,N_4880,N_4844);
nor UO_851 (O_851,N_4922,N_4816);
and UO_852 (O_852,N_4959,N_4845);
and UO_853 (O_853,N_4830,N_4804);
and UO_854 (O_854,N_4885,N_4892);
and UO_855 (O_855,N_4829,N_4971);
xor UO_856 (O_856,N_4922,N_4800);
nor UO_857 (O_857,N_4866,N_4912);
xor UO_858 (O_858,N_4913,N_4879);
or UO_859 (O_859,N_4848,N_4820);
xnor UO_860 (O_860,N_4855,N_4905);
or UO_861 (O_861,N_4909,N_4942);
xnor UO_862 (O_862,N_4998,N_4966);
nand UO_863 (O_863,N_4936,N_4850);
or UO_864 (O_864,N_4920,N_4870);
and UO_865 (O_865,N_4850,N_4961);
nor UO_866 (O_866,N_4862,N_4933);
and UO_867 (O_867,N_4844,N_4971);
xnor UO_868 (O_868,N_4868,N_4952);
nor UO_869 (O_869,N_4968,N_4882);
nand UO_870 (O_870,N_4827,N_4991);
nor UO_871 (O_871,N_4927,N_4911);
nand UO_872 (O_872,N_4973,N_4852);
nand UO_873 (O_873,N_4866,N_4967);
or UO_874 (O_874,N_4976,N_4969);
or UO_875 (O_875,N_4945,N_4952);
nand UO_876 (O_876,N_4828,N_4952);
and UO_877 (O_877,N_4993,N_4984);
or UO_878 (O_878,N_4863,N_4925);
xor UO_879 (O_879,N_4843,N_4874);
and UO_880 (O_880,N_4931,N_4853);
and UO_881 (O_881,N_4813,N_4973);
nor UO_882 (O_882,N_4843,N_4820);
and UO_883 (O_883,N_4941,N_4955);
nor UO_884 (O_884,N_4935,N_4860);
xnor UO_885 (O_885,N_4996,N_4927);
nor UO_886 (O_886,N_4877,N_4852);
xnor UO_887 (O_887,N_4813,N_4830);
and UO_888 (O_888,N_4809,N_4863);
nand UO_889 (O_889,N_4911,N_4905);
or UO_890 (O_890,N_4959,N_4882);
nor UO_891 (O_891,N_4972,N_4853);
or UO_892 (O_892,N_4944,N_4801);
and UO_893 (O_893,N_4839,N_4914);
or UO_894 (O_894,N_4961,N_4818);
or UO_895 (O_895,N_4988,N_4905);
xnor UO_896 (O_896,N_4983,N_4836);
xnor UO_897 (O_897,N_4983,N_4962);
xnor UO_898 (O_898,N_4893,N_4819);
nand UO_899 (O_899,N_4958,N_4948);
xor UO_900 (O_900,N_4933,N_4981);
nor UO_901 (O_901,N_4848,N_4924);
and UO_902 (O_902,N_4884,N_4854);
xnor UO_903 (O_903,N_4969,N_4962);
and UO_904 (O_904,N_4866,N_4928);
nand UO_905 (O_905,N_4943,N_4847);
nor UO_906 (O_906,N_4853,N_4828);
nand UO_907 (O_907,N_4862,N_4920);
nand UO_908 (O_908,N_4867,N_4800);
and UO_909 (O_909,N_4967,N_4951);
nand UO_910 (O_910,N_4949,N_4951);
and UO_911 (O_911,N_4893,N_4809);
or UO_912 (O_912,N_4895,N_4905);
xnor UO_913 (O_913,N_4898,N_4908);
or UO_914 (O_914,N_4891,N_4893);
and UO_915 (O_915,N_4931,N_4880);
nand UO_916 (O_916,N_4816,N_4853);
and UO_917 (O_917,N_4952,N_4998);
nand UO_918 (O_918,N_4879,N_4808);
nor UO_919 (O_919,N_4908,N_4875);
nand UO_920 (O_920,N_4805,N_4935);
xnor UO_921 (O_921,N_4911,N_4925);
nor UO_922 (O_922,N_4808,N_4948);
xnor UO_923 (O_923,N_4867,N_4896);
nand UO_924 (O_924,N_4922,N_4848);
nand UO_925 (O_925,N_4853,N_4955);
or UO_926 (O_926,N_4820,N_4974);
and UO_927 (O_927,N_4800,N_4906);
xnor UO_928 (O_928,N_4817,N_4977);
nand UO_929 (O_929,N_4897,N_4969);
and UO_930 (O_930,N_4862,N_4867);
or UO_931 (O_931,N_4977,N_4858);
xor UO_932 (O_932,N_4911,N_4985);
nor UO_933 (O_933,N_4984,N_4829);
and UO_934 (O_934,N_4965,N_4854);
xnor UO_935 (O_935,N_4820,N_4935);
and UO_936 (O_936,N_4941,N_4886);
xor UO_937 (O_937,N_4975,N_4931);
nor UO_938 (O_938,N_4879,N_4903);
nand UO_939 (O_939,N_4916,N_4841);
nand UO_940 (O_940,N_4956,N_4897);
and UO_941 (O_941,N_4809,N_4846);
and UO_942 (O_942,N_4936,N_4982);
and UO_943 (O_943,N_4925,N_4923);
xnor UO_944 (O_944,N_4893,N_4862);
nand UO_945 (O_945,N_4992,N_4884);
xor UO_946 (O_946,N_4920,N_4988);
xnor UO_947 (O_947,N_4892,N_4954);
nor UO_948 (O_948,N_4854,N_4930);
nor UO_949 (O_949,N_4899,N_4844);
or UO_950 (O_950,N_4851,N_4943);
nor UO_951 (O_951,N_4904,N_4891);
xor UO_952 (O_952,N_4923,N_4856);
nor UO_953 (O_953,N_4901,N_4850);
or UO_954 (O_954,N_4880,N_4881);
and UO_955 (O_955,N_4858,N_4949);
nand UO_956 (O_956,N_4898,N_4936);
or UO_957 (O_957,N_4911,N_4943);
xnor UO_958 (O_958,N_4986,N_4964);
nand UO_959 (O_959,N_4905,N_4939);
and UO_960 (O_960,N_4931,N_4976);
nor UO_961 (O_961,N_4841,N_4962);
and UO_962 (O_962,N_4874,N_4844);
nand UO_963 (O_963,N_4911,N_4955);
nand UO_964 (O_964,N_4991,N_4875);
xor UO_965 (O_965,N_4999,N_4832);
or UO_966 (O_966,N_4812,N_4996);
and UO_967 (O_967,N_4939,N_4965);
nand UO_968 (O_968,N_4926,N_4940);
or UO_969 (O_969,N_4897,N_4863);
and UO_970 (O_970,N_4934,N_4838);
xor UO_971 (O_971,N_4857,N_4871);
nand UO_972 (O_972,N_4905,N_4822);
and UO_973 (O_973,N_4828,N_4930);
xor UO_974 (O_974,N_4869,N_4802);
or UO_975 (O_975,N_4825,N_4935);
or UO_976 (O_976,N_4931,N_4840);
or UO_977 (O_977,N_4979,N_4920);
nor UO_978 (O_978,N_4998,N_4930);
nor UO_979 (O_979,N_4838,N_4808);
or UO_980 (O_980,N_4937,N_4857);
or UO_981 (O_981,N_4801,N_4919);
xor UO_982 (O_982,N_4928,N_4824);
nor UO_983 (O_983,N_4913,N_4918);
nor UO_984 (O_984,N_4812,N_4878);
and UO_985 (O_985,N_4840,N_4837);
nor UO_986 (O_986,N_4929,N_4801);
or UO_987 (O_987,N_4846,N_4950);
nor UO_988 (O_988,N_4800,N_4893);
xor UO_989 (O_989,N_4882,N_4866);
and UO_990 (O_990,N_4902,N_4952);
or UO_991 (O_991,N_4815,N_4938);
and UO_992 (O_992,N_4866,N_4808);
xnor UO_993 (O_993,N_4923,N_4858);
and UO_994 (O_994,N_4877,N_4821);
nand UO_995 (O_995,N_4997,N_4934);
and UO_996 (O_996,N_4802,N_4826);
nand UO_997 (O_997,N_4915,N_4808);
or UO_998 (O_998,N_4909,N_4863);
xor UO_999 (O_999,N_4981,N_4984);
endmodule