module basic_5000_50000_5000_200_levels_10xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_2672,In_212);
or U1 (N_1,In_51,In_279);
nor U2 (N_2,In_3620,In_3203);
and U3 (N_3,In_4593,In_293);
and U4 (N_4,In_4038,In_4008);
nor U5 (N_5,In_3231,In_3247);
or U6 (N_6,In_204,In_4331);
xor U7 (N_7,In_3444,In_2218);
and U8 (N_8,In_1584,In_3398);
and U9 (N_9,In_2289,In_2582);
nand U10 (N_10,In_492,In_642);
or U11 (N_11,In_4230,In_441);
and U12 (N_12,In_1357,In_3222);
nor U13 (N_13,In_2245,In_4075);
or U14 (N_14,In_300,In_1002);
and U15 (N_15,In_4813,In_3493);
or U16 (N_16,In_4445,In_3635);
or U17 (N_17,In_2286,In_3470);
nand U18 (N_18,In_3586,In_1562);
xnor U19 (N_19,In_2013,In_2921);
and U20 (N_20,In_1711,In_4487);
xnor U21 (N_21,In_3202,In_4618);
nor U22 (N_22,In_86,In_382);
nand U23 (N_23,In_1999,In_550);
nand U24 (N_24,In_4545,In_2327);
xor U25 (N_25,In_3782,In_2901);
nand U26 (N_26,In_30,In_4617);
nor U27 (N_27,In_3916,In_3336);
xor U28 (N_28,In_1590,In_1563);
nor U29 (N_29,In_4962,In_1102);
or U30 (N_30,In_3,In_1627);
or U31 (N_31,In_237,In_2250);
nand U32 (N_32,In_2100,In_4291);
or U33 (N_33,In_3564,In_3861);
or U34 (N_34,In_3577,In_1603);
or U35 (N_35,In_3109,In_4055);
nor U36 (N_36,In_2171,In_3727);
nor U37 (N_37,In_788,In_3058);
xor U38 (N_38,In_1730,In_2898);
nor U39 (N_39,In_4227,In_3843);
xnor U40 (N_40,In_4447,In_1426);
nand U41 (N_41,In_622,In_1462);
or U42 (N_42,In_2263,In_3261);
nand U43 (N_43,In_914,In_3223);
nand U44 (N_44,In_2653,In_2925);
and U45 (N_45,In_2907,In_571);
and U46 (N_46,In_2429,In_3802);
and U47 (N_47,In_1371,In_4689);
nor U48 (N_48,In_7,In_1507);
or U49 (N_49,In_2365,In_50);
and U50 (N_50,In_2081,In_503);
nor U51 (N_51,In_4179,In_83);
xor U52 (N_52,In_4773,In_3950);
xnor U53 (N_53,In_1145,In_2937);
and U54 (N_54,In_27,In_2500);
and U55 (N_55,In_250,In_1119);
nor U56 (N_56,In_3434,In_573);
nor U57 (N_57,In_3719,In_4426);
xor U58 (N_58,In_2308,In_748);
xnor U59 (N_59,In_1609,In_1015);
nor U60 (N_60,In_1342,In_4882);
and U61 (N_61,In_2232,In_2864);
nand U62 (N_62,In_4595,In_4697);
xor U63 (N_63,In_4368,In_3491);
or U64 (N_64,In_3787,In_984);
and U65 (N_65,In_1064,In_3057);
and U66 (N_66,In_2798,In_388);
nor U67 (N_67,In_4613,In_4442);
and U68 (N_68,In_3944,In_1991);
xor U69 (N_69,In_2242,In_4135);
and U70 (N_70,In_843,In_760);
or U71 (N_71,In_4413,In_1319);
nand U72 (N_72,In_63,In_1530);
nor U73 (N_73,In_2216,In_3121);
xor U74 (N_74,In_3668,In_2778);
xnor U75 (N_75,In_2865,In_2079);
and U76 (N_76,In_4764,In_4349);
nand U77 (N_77,In_3063,In_761);
nand U78 (N_78,In_1925,In_2393);
nor U79 (N_79,In_581,In_4809);
and U80 (N_80,In_3661,In_1317);
and U81 (N_81,In_3786,In_2652);
nand U82 (N_82,In_383,In_1404);
nand U83 (N_83,In_3485,In_1818);
nand U84 (N_84,In_2987,In_4673);
and U85 (N_85,In_1679,In_3189);
or U86 (N_86,In_34,In_3242);
nor U87 (N_87,In_1252,In_1370);
and U88 (N_88,In_3171,In_2063);
nand U89 (N_89,In_810,In_498);
and U90 (N_90,In_4155,In_3215);
xnor U91 (N_91,In_494,In_781);
and U92 (N_92,In_2427,In_3753);
nand U93 (N_93,In_4925,In_3913);
and U94 (N_94,In_1196,In_4502);
nor U95 (N_95,In_158,In_3298);
and U96 (N_96,In_1114,In_3928);
and U97 (N_97,In_3911,In_2868);
nor U98 (N_98,In_828,In_3572);
and U99 (N_99,In_2515,In_3300);
nor U100 (N_100,In_1551,In_2357);
nand U101 (N_101,In_4754,In_2841);
xor U102 (N_102,In_4162,In_4282);
nand U103 (N_103,In_1694,In_2387);
and U104 (N_104,In_4558,In_1501);
and U105 (N_105,In_2311,In_1918);
or U106 (N_106,In_4831,In_2852);
and U107 (N_107,In_3854,In_768);
xor U108 (N_108,In_990,In_4889);
xor U109 (N_109,In_3914,In_95);
or U110 (N_110,In_2636,In_3721);
nor U111 (N_111,In_629,In_2295);
nand U112 (N_112,In_1546,In_3770);
xor U113 (N_113,In_812,In_4430);
nor U114 (N_114,In_2655,In_4881);
nor U115 (N_115,In_532,In_1979);
or U116 (N_116,In_873,In_2473);
nand U117 (N_117,In_1200,In_2477);
xor U118 (N_118,In_3137,In_4695);
nand U119 (N_119,In_4158,In_1366);
xor U120 (N_120,In_1350,In_242);
and U121 (N_121,In_4102,In_3013);
nor U122 (N_122,In_2993,In_2256);
nand U123 (N_123,In_970,In_2619);
nand U124 (N_124,In_3471,In_3646);
xnor U125 (N_125,In_1518,In_675);
nor U126 (N_126,In_848,In_1403);
or U127 (N_127,In_4559,In_696);
nand U128 (N_128,In_2447,In_1192);
nor U129 (N_129,In_4827,In_3036);
and U130 (N_130,In_2625,In_5);
nor U131 (N_131,In_2066,In_3847);
nor U132 (N_132,In_3001,In_2396);
or U133 (N_133,In_4816,In_2708);
nand U134 (N_134,In_3772,In_3329);
xor U135 (N_135,In_4164,In_3450);
or U136 (N_136,In_1175,In_4283);
and U137 (N_137,In_2633,In_4619);
and U138 (N_138,In_1227,In_3575);
nor U139 (N_139,In_1464,In_4190);
and U140 (N_140,In_949,In_4257);
nor U141 (N_141,In_2627,In_3025);
nor U142 (N_142,In_2826,In_180);
xnor U143 (N_143,In_4492,In_1848);
nor U144 (N_144,In_4337,In_167);
nand U145 (N_145,In_4737,In_256);
xnor U146 (N_146,In_4045,In_1491);
xnor U147 (N_147,In_2744,In_1337);
or U148 (N_148,In_4687,In_2193);
xnor U149 (N_149,In_3838,In_3937);
xnor U150 (N_150,In_897,In_4350);
nor U151 (N_151,In_678,In_4260);
and U152 (N_152,In_1374,In_2463);
and U153 (N_153,In_1224,In_2374);
or U154 (N_154,In_3659,In_138);
or U155 (N_155,In_1586,In_4078);
nand U156 (N_156,In_3554,In_4043);
nand U157 (N_157,In_3645,In_1014);
nor U158 (N_158,In_1263,In_1556);
nand U159 (N_159,In_916,In_2843);
and U160 (N_160,In_1110,In_1205);
xnor U161 (N_161,In_3412,In_1011);
nor U162 (N_162,In_3437,In_4016);
and U163 (N_163,In_3680,In_2389);
and U164 (N_164,In_3875,In_1468);
nand U165 (N_165,In_3037,In_718);
nor U166 (N_166,In_1895,In_1639);
and U167 (N_167,In_4157,In_405);
xor U168 (N_168,In_521,In_1959);
and U169 (N_169,In_4698,In_3839);
or U170 (N_170,In_4148,In_4005);
and U171 (N_171,In_1702,In_2647);
nand U172 (N_172,In_4770,In_3157);
nand U173 (N_173,In_3342,In_4551);
xnor U174 (N_174,In_1054,In_2551);
or U175 (N_175,In_906,In_1634);
or U176 (N_176,In_3846,In_4986);
or U177 (N_177,In_3938,In_2153);
nand U178 (N_178,In_393,In_2398);
xnor U179 (N_179,In_4480,In_1314);
and U180 (N_180,In_3009,In_2280);
nor U181 (N_181,In_663,In_1037);
and U182 (N_182,In_745,In_4960);
or U183 (N_183,In_556,In_88);
or U184 (N_184,In_4215,In_3168);
and U185 (N_185,In_4598,In_385);
or U186 (N_186,In_4408,In_3724);
and U187 (N_187,In_3278,In_2364);
nor U188 (N_188,In_4917,In_1157);
nor U189 (N_189,In_3284,In_4700);
nand U190 (N_190,In_1613,In_2140);
or U191 (N_191,In_4467,In_3941);
nor U192 (N_192,In_2668,In_2565);
nand U193 (N_193,In_2831,In_2739);
nand U194 (N_194,In_1475,In_2645);
xor U195 (N_195,In_926,In_4250);
nor U196 (N_196,In_2342,In_3703);
or U197 (N_197,In_3014,In_3218);
nor U198 (N_198,In_3503,In_2526);
and U199 (N_199,In_553,In_942);
nor U200 (N_200,In_4649,In_2036);
xor U201 (N_201,In_4900,In_486);
xnor U202 (N_202,In_1254,In_4824);
and U203 (N_203,In_1202,In_3663);
nor U204 (N_204,In_268,In_3385);
xnor U205 (N_205,In_484,In_2956);
xor U206 (N_206,In_196,In_766);
nand U207 (N_207,In_4767,In_3055);
xnor U208 (N_208,In_4108,In_451);
nor U209 (N_209,In_3065,In_2806);
or U210 (N_210,In_946,In_836);
nor U211 (N_211,In_1940,In_3428);
nand U212 (N_212,In_3373,In_1410);
and U213 (N_213,In_1537,In_436);
nand U214 (N_214,In_3833,In_3881);
and U215 (N_215,In_2021,In_850);
or U216 (N_216,In_1174,In_3602);
nor U217 (N_217,In_3946,In_4125);
or U218 (N_218,In_2069,In_2597);
and U219 (N_219,In_3309,In_2958);
nor U220 (N_220,In_122,In_2839);
xnor U221 (N_221,In_3762,In_1163);
nor U222 (N_222,In_587,In_3041);
xnor U223 (N_223,In_1296,In_4738);
or U224 (N_224,In_46,In_1542);
or U225 (N_225,In_2998,In_2438);
nor U226 (N_226,In_2321,In_1273);
nand U227 (N_227,In_2718,In_4952);
nor U228 (N_228,In_2492,In_1621);
or U229 (N_229,In_4828,In_4171);
and U230 (N_230,In_3106,In_1868);
or U231 (N_231,In_4264,In_2705);
or U232 (N_232,In_1872,In_2566);
nor U233 (N_233,In_2641,In_341);
xnor U234 (N_234,In_2444,In_3988);
nor U235 (N_235,In_3178,In_3143);
or U236 (N_236,In_728,In_4417);
xor U237 (N_237,In_4632,In_1599);
and U238 (N_238,In_244,In_4775);
xor U239 (N_239,In_4183,In_1792);
nand U240 (N_240,In_1664,In_2361);
or U241 (N_241,In_71,In_3174);
or U242 (N_242,In_4223,In_1655);
or U243 (N_243,In_3514,In_202);
xor U244 (N_244,In_4138,In_3478);
nor U245 (N_245,In_3370,In_1845);
or U246 (N_246,In_4959,In_1983);
nand U247 (N_247,In_2061,In_4829);
or U248 (N_248,In_634,In_218);
and U249 (N_249,In_1907,In_834);
nand U250 (N_250,In_1837,In_2423);
nand U251 (N_251,In_4518,In_1593);
nand U252 (N_252,In_4957,In_2493);
nand U253 (N_253,In_4109,In_2740);
nand U254 (N_254,In_753,In_2375);
nor U255 (N_255,In_4052,In_4888);
xnor U256 (N_256,In_2455,In_4065);
xnor U257 (N_257,In_2014,In_3985);
xnor U258 (N_258,In_882,In_2189);
nand U259 (N_259,In_3998,In_857);
xor U260 (N_260,In_2975,In_937);
xor U261 (N_261,N_241,In_183);
nand U262 (N_262,In_3751,In_1529);
xor U263 (N_263,In_1550,In_3389);
xnor U264 (N_264,In_2728,In_909);
or U265 (N_265,In_2680,In_4678);
nor U266 (N_266,In_4963,In_1216);
or U267 (N_267,In_1651,In_4652);
and U268 (N_268,In_4884,In_1522);
nor U269 (N_269,In_1813,In_854);
or U270 (N_270,In_1781,In_2884);
and U271 (N_271,In_582,In_246);
nor U272 (N_272,In_844,In_1168);
nand U273 (N_273,In_3987,In_1355);
xnor U274 (N_274,In_4378,In_3685);
nand U275 (N_275,In_4616,In_1406);
nand U276 (N_276,In_621,In_3371);
nor U277 (N_277,In_2940,In_738);
nand U278 (N_278,In_2318,In_4498);
nor U279 (N_279,In_996,In_704);
nor U280 (N_280,In_1135,In_4036);
nor U281 (N_281,In_431,In_2715);
nor U282 (N_282,N_27,In_260);
xor U283 (N_283,In_4107,In_3994);
and U284 (N_284,In_4339,In_1343);
nand U285 (N_285,In_968,In_506);
xor U286 (N_286,In_4848,In_3896);
nor U287 (N_287,In_4566,In_1053);
xor U288 (N_288,In_4721,In_400);
nand U289 (N_289,In_2032,In_1121);
nor U290 (N_290,In_731,In_3032);
or U291 (N_291,N_195,In_1714);
xnor U292 (N_292,In_780,In_2938);
nand U293 (N_293,In_3259,In_3170);
and U294 (N_294,In_3636,In_4949);
nand U295 (N_295,In_2331,In_3404);
or U296 (N_296,In_1391,In_1631);
or U297 (N_297,In_2300,In_387);
and U298 (N_298,In_4175,In_2220);
or U299 (N_299,In_2019,In_3765);
or U300 (N_300,In_343,In_3246);
nor U301 (N_301,N_64,In_2310);
or U302 (N_302,In_3324,In_4757);
and U303 (N_303,In_1800,In_4066);
nand U304 (N_304,In_1187,In_2346);
or U305 (N_305,In_4948,In_3495);
nor U306 (N_306,In_4074,In_53);
nand U307 (N_307,In_4869,N_211);
nand U308 (N_308,In_2070,In_4051);
nand U309 (N_309,In_29,N_31);
xnor U310 (N_310,In_1698,In_3255);
xnor U311 (N_311,In_3297,In_2453);
nand U312 (N_312,N_139,N_36);
and U313 (N_313,In_3360,In_1221);
nand U314 (N_314,In_786,In_2943);
nor U315 (N_315,In_3673,In_1284);
nor U316 (N_316,In_1877,In_3581);
xnor U317 (N_317,In_2134,In_1065);
xor U318 (N_318,In_1238,N_96);
xnor U319 (N_319,In_3699,In_4920);
or U320 (N_320,In_2176,In_1384);
and U321 (N_321,In_2598,In_153);
nor U322 (N_322,In_478,In_4207);
xnor U323 (N_323,In_1286,In_3547);
and U324 (N_324,In_2905,In_1043);
nor U325 (N_325,In_1452,In_2424);
xor U326 (N_326,In_1796,In_3243);
xnor U327 (N_327,In_560,In_1799);
and U328 (N_328,N_160,In_3294);
nand U329 (N_329,In_2191,In_3903);
and U330 (N_330,In_2779,In_3096);
nor U331 (N_331,In_427,In_3871);
and U332 (N_332,In_2600,In_752);
nand U333 (N_333,In_2157,In_1707);
nor U334 (N_334,In_13,In_1294);
nand U335 (N_335,In_479,In_1425);
nor U336 (N_336,In_4414,In_2351);
xor U337 (N_337,In_1438,N_16);
and U338 (N_338,In_1289,In_773);
or U339 (N_339,In_1480,In_1571);
xor U340 (N_340,In_1885,In_1873);
or U341 (N_341,In_3618,In_1675);
and U342 (N_342,In_1676,In_4340);
and U343 (N_343,In_4251,In_4063);
xnor U344 (N_344,In_2887,In_2369);
nor U345 (N_345,In_2742,In_966);
xnor U346 (N_346,In_4565,In_4760);
or U347 (N_347,In_572,In_998);
nand U348 (N_348,In_822,In_4496);
nor U349 (N_349,N_12,In_1098);
nor U350 (N_350,In_2736,In_4583);
or U351 (N_351,In_3502,In_1674);
or U352 (N_352,In_4638,In_2312);
xnor U353 (N_353,In_2121,In_956);
nor U354 (N_354,In_3965,In_4685);
xor U355 (N_355,In_1585,In_2961);
xnor U356 (N_356,In_2812,In_1018);
nor U357 (N_357,In_625,In_1010);
or U358 (N_358,In_4197,In_3926);
and U359 (N_359,N_115,In_2018);
nand U360 (N_360,In_4653,In_2785);
nand U361 (N_361,In_3353,In_3117);
and U362 (N_362,In_4573,In_4819);
xnor U363 (N_363,In_1798,In_774);
nor U364 (N_364,In_3886,In_784);
nand U365 (N_365,In_4048,In_1034);
nor U366 (N_366,In_4365,In_4533);
or U367 (N_367,In_3849,In_390);
and U368 (N_368,In_4859,In_4650);
or U369 (N_369,In_1966,In_4783);
or U370 (N_370,In_28,In_2382);
and U371 (N_371,In_1352,In_3200);
and U372 (N_372,In_4299,In_378);
nand U373 (N_373,In_1269,In_1170);
and U374 (N_374,In_1444,In_959);
nand U375 (N_375,In_4577,In_1594);
nand U376 (N_376,In_500,In_2015);
and U377 (N_377,In_3570,N_44);
and U378 (N_378,In_1884,In_2888);
nor U379 (N_379,In_1922,In_1304);
and U380 (N_380,In_1368,In_3337);
xor U381 (N_381,In_4727,In_4973);
nor U382 (N_382,In_3672,In_4720);
nand U383 (N_383,In_640,In_1880);
nand U384 (N_384,In_4733,In_1734);
nand U385 (N_385,In_1422,In_1012);
and U386 (N_386,In_4374,In_4805);
xnor U387 (N_387,In_2129,In_4424);
or U388 (N_388,N_127,In_4594);
nand U389 (N_389,In_4865,In_3081);
xor U390 (N_390,In_2159,In_3400);
and U391 (N_391,In_386,In_3533);
nand U392 (N_392,In_2319,In_3446);
nor U393 (N_393,In_1239,In_4316);
and U394 (N_394,In_3904,N_175);
or U395 (N_395,In_2264,In_3757);
and U396 (N_396,In_3214,In_2316);
or U397 (N_397,In_1000,In_3158);
or U398 (N_398,In_953,In_1649);
nor U399 (N_399,In_4853,In_487);
nor U400 (N_400,In_449,In_4206);
and U401 (N_401,In_614,In_694);
nor U402 (N_402,In_1724,In_4462);
xor U403 (N_403,In_4851,In_4576);
or U404 (N_404,In_4235,In_4429);
nand U405 (N_405,In_2635,In_1299);
or U406 (N_406,In_3474,In_908);
nor U407 (N_407,In_2725,In_938);
or U408 (N_408,In_141,In_2114);
nand U409 (N_409,In_252,In_679);
or U410 (N_410,In_3534,N_225);
and U411 (N_411,In_4076,In_3052);
nor U412 (N_412,In_1887,In_1819);
xnor U413 (N_413,In_865,In_1259);
and U414 (N_414,In_2665,In_3104);
and U415 (N_415,In_2051,In_2776);
nor U416 (N_416,In_1128,In_1757);
xor U417 (N_417,In_2807,In_3971);
nand U418 (N_418,In_409,In_2758);
xor U419 (N_419,N_238,In_1693);
nor U420 (N_420,In_3455,In_1078);
xnor U421 (N_421,In_1625,In_4675);
and U422 (N_422,In_1048,In_2353);
xnor U423 (N_423,In_1946,In_1860);
xnor U424 (N_424,In_3667,In_3520);
or U425 (N_425,In_868,In_3049);
or U426 (N_426,In_2080,In_4379);
nand U427 (N_427,In_195,In_3548);
nor U428 (N_428,In_3744,In_4627);
and U429 (N_429,N_66,In_3466);
xor U430 (N_430,In_1732,In_2596);
nor U431 (N_431,In_243,In_4802);
xnor U432 (N_432,In_4112,In_3420);
nor U433 (N_433,In_4401,In_824);
or U434 (N_434,In_448,In_2354);
nand U435 (N_435,In_803,In_4755);
nor U436 (N_436,In_1081,In_2208);
nand U437 (N_437,In_1283,In_2689);
and U438 (N_438,In_2446,In_615);
nand U439 (N_439,In_2099,In_8);
and U440 (N_440,In_4605,In_2927);
nor U441 (N_441,N_207,In_2459);
or U442 (N_442,In_3964,In_2096);
nand U443 (N_443,In_2702,In_2158);
or U444 (N_444,In_4579,In_4736);
xor U445 (N_445,In_4482,In_2194);
xor U446 (N_446,In_1909,In_3417);
nor U447 (N_447,In_688,In_1127);
nor U448 (N_448,In_720,In_1295);
nand U449 (N_449,In_567,In_2829);
nand U450 (N_450,In_3760,In_3856);
and U451 (N_451,In_460,In_2543);
and U452 (N_452,N_156,In_1620);
and U453 (N_453,In_4317,In_4243);
and U454 (N_454,In_2719,In_3167);
nor U455 (N_455,In_2646,In_3225);
and U456 (N_456,In_883,In_4792);
nor U457 (N_457,In_3567,In_2409);
xnor U458 (N_458,In_1225,In_1827);
or U459 (N_459,In_434,In_325);
nand U460 (N_460,In_3026,In_1995);
or U461 (N_461,In_3494,In_4961);
and U462 (N_462,In_3648,In_627);
or U463 (N_463,In_3745,In_3603);
or U464 (N_464,In_1681,In_2624);
nand U465 (N_465,In_2580,In_4984);
nand U466 (N_466,In_4297,In_4312);
nor U467 (N_467,In_3599,In_113);
nor U468 (N_468,In_2105,In_3459);
or U469 (N_469,In_2416,In_45);
and U470 (N_470,In_1005,In_4823);
xnor U471 (N_471,In_4694,In_1510);
nor U472 (N_472,In_4569,In_3566);
xor U473 (N_473,In_3758,In_1185);
xnor U474 (N_474,In_4057,In_160);
and U475 (N_475,In_2593,In_2913);
xnor U476 (N_476,In_1178,In_3145);
nand U477 (N_477,In_207,In_2230);
and U478 (N_478,In_3669,In_971);
xnor U479 (N_479,In_2323,In_884);
and U480 (N_480,In_2752,N_71);
nor U481 (N_481,In_3558,In_3908);
xor U482 (N_482,In_2669,In_4580);
nand U483 (N_483,In_2452,In_2881);
nand U484 (N_484,In_713,In_3867);
nor U485 (N_485,In_2714,In_1326);
and U486 (N_486,In_4095,In_4489);
and U487 (N_487,In_777,In_1142);
xor U488 (N_488,In_301,In_1743);
or U489 (N_489,In_3596,In_3688);
xor U490 (N_490,In_1623,In_3810);
xor U491 (N_491,In_1692,In_889);
or U492 (N_492,In_2980,In_1842);
nor U493 (N_493,In_1423,In_518);
and U494 (N_494,In_1046,In_2584);
and U495 (N_495,In_1672,In_3276);
nand U496 (N_496,N_26,In_1708);
nand U497 (N_497,In_4448,In_1817);
and U498 (N_498,In_3028,In_1307);
and U499 (N_499,In_878,In_468);
nand U500 (N_500,In_1323,In_3201);
nor U501 (N_501,In_3414,In_2867);
or U502 (N_502,In_307,In_1553);
xnor U503 (N_503,N_260,In_1057);
nand U504 (N_504,In_381,In_2215);
nand U505 (N_505,In_3837,In_2296);
xor U506 (N_506,N_28,In_68);
nand U507 (N_507,In_206,In_4050);
nor U508 (N_508,In_1500,N_252);
or U509 (N_509,In_2336,In_2540);
xnor U510 (N_510,In_2957,In_4987);
and U511 (N_511,In_1104,In_3084);
nand U512 (N_512,In_2879,In_4037);
xor U513 (N_513,In_4586,In_4740);
and U514 (N_514,In_796,In_4412);
nor U515 (N_515,In_4292,In_2432);
nor U516 (N_516,In_2089,In_826);
nand U517 (N_517,In_1437,In_3741);
nor U518 (N_518,In_4123,In_3069);
and U519 (N_519,In_2322,In_1742);
and U520 (N_520,In_4472,In_840);
nor U521 (N_521,In_1935,In_1165);
and U522 (N_522,N_142,In_644);
nor U523 (N_523,N_384,In_4259);
and U524 (N_524,In_89,In_711);
and U525 (N_525,In_318,In_2339);
nor U526 (N_526,In_680,In_1808);
and U527 (N_527,In_3356,In_4766);
nor U528 (N_528,In_4947,In_4130);
or U529 (N_529,In_1565,N_499);
or U530 (N_530,In_2476,N_274);
and U531 (N_531,In_3447,In_4507);
nor U532 (N_532,In_4200,In_540);
xor U533 (N_533,In_4741,In_2461);
nand U534 (N_534,In_240,In_150);
xnor U535 (N_535,In_4343,In_3194);
xor U536 (N_536,In_2797,In_2040);
or U537 (N_537,In_277,In_819);
nand U538 (N_538,In_2164,In_4041);
or U539 (N_539,In_3769,In_3187);
nand U540 (N_540,In_2192,In_4274);
or U541 (N_541,In_3866,In_3034);
nand U542 (N_542,In_3399,In_2556);
xor U543 (N_543,N_138,In_2349);
nor U544 (N_544,In_2657,In_76);
and U545 (N_545,In_2882,In_471);
nor U546 (N_546,In_4040,In_2609);
xor U547 (N_547,In_2974,In_2794);
nor U548 (N_548,In_184,In_3989);
nand U549 (N_549,In_3482,N_258);
nand U550 (N_550,In_2275,In_3522);
nand U551 (N_551,In_4601,In_4013);
or U552 (N_552,In_2620,In_4383);
and U553 (N_553,In_1466,N_168);
xor U554 (N_554,In_4071,In_4511);
nand U555 (N_555,In_3984,In_1485);
nor U556 (N_556,N_278,N_72);
or U557 (N_557,In_1099,In_536);
and U558 (N_558,In_1369,In_3864);
xnor U559 (N_559,In_2403,N_83);
and U560 (N_560,In_2787,In_3605);
nor U561 (N_561,N_154,In_4967);
nand U562 (N_562,In_4835,In_2373);
and U563 (N_563,N_346,In_159);
nand U564 (N_564,In_584,In_4003);
or U565 (N_565,In_490,In_3536);
xor U566 (N_566,In_602,In_1129);
or U567 (N_567,In_3731,In_2163);
nand U568 (N_568,In_1007,N_411);
and U569 (N_569,In_3579,In_4506);
and U570 (N_570,In_2771,In_4825);
nand U571 (N_571,In_3708,In_4212);
nor U572 (N_572,In_1067,In_1017);
and U573 (N_573,In_554,In_4072);
or U574 (N_574,In_658,In_4033);
or U575 (N_575,N_354,N_357);
nand U576 (N_576,In_2002,In_3940);
xor U577 (N_577,In_3879,In_516);
or U578 (N_578,In_4384,In_144);
nand U579 (N_579,In_2803,In_4493);
nor U580 (N_580,N_176,In_2437);
nor U581 (N_581,In_1281,In_1496);
nor U582 (N_582,In_3059,In_3876);
nor U583 (N_583,In_148,In_4198);
or U584 (N_584,In_4715,In_4642);
and U585 (N_585,In_549,In_1395);
or U586 (N_586,In_2111,In_509);
nor U587 (N_587,N_81,In_1419);
and U588 (N_588,In_1558,In_510);
xnor U589 (N_589,In_371,In_1635);
xor U590 (N_590,In_1658,In_726);
nor U591 (N_591,In_2630,In_4437);
nand U592 (N_592,In_4931,N_388);
and U593 (N_593,In_3358,In_1362);
and U594 (N_594,In_763,In_177);
and U595 (N_595,In_4988,N_420);
and U596 (N_596,In_1663,In_656);
xor U597 (N_597,In_881,In_3445);
or U598 (N_598,In_4803,N_320);
nand U599 (N_599,In_2840,In_818);
xnor U600 (N_600,In_755,In_1070);
xor U601 (N_601,In_472,In_2345);
nor U602 (N_602,In_1667,In_499);
and U603 (N_603,In_1132,In_3925);
nor U604 (N_604,In_4538,In_4271);
or U605 (N_605,In_1648,In_3710);
xnor U606 (N_606,In_4213,In_1784);
nand U607 (N_607,N_361,In_2408);
nand U608 (N_608,In_1080,In_3774);
nor U609 (N_609,In_2947,In_3626);
nor U610 (N_610,In_2536,In_1063);
xnor U611 (N_611,In_930,In_3869);
and U612 (N_612,In_2834,N_308);
xnor U613 (N_613,In_3429,In_224);
nand U614 (N_614,In_1770,N_377);
xnor U615 (N_615,N_271,In_2537);
xor U616 (N_616,In_485,In_75);
or U617 (N_617,In_4796,In_3900);
or U618 (N_618,In_2084,In_1630);
or U619 (N_619,In_172,In_3481);
nor U620 (N_620,In_2183,In_3282);
nor U621 (N_621,In_1461,In_894);
and U622 (N_622,In_4064,In_130);
and U623 (N_623,In_1829,In_1197);
nand U624 (N_624,In_4781,In_1705);
or U625 (N_625,N_439,In_1446);
xnor U626 (N_626,In_2880,In_2755);
nand U627 (N_627,In_1731,In_345);
and U628 (N_628,In_3637,In_3649);
or U629 (N_629,In_825,In_3365);
nand U630 (N_630,N_336,In_2024);
xnor U631 (N_631,N_259,In_1409);
and U632 (N_632,In_2727,N_166);
nor U633 (N_633,N_9,In_2156);
nand U634 (N_634,In_4555,In_3110);
and U635 (N_635,In_3248,In_4185);
nor U636 (N_636,N_223,In_78);
xnor U637 (N_637,N_441,In_1210);
nor U638 (N_638,In_4991,N_148);
nor U639 (N_639,In_3997,In_1079);
nand U640 (N_640,N_152,In_1270);
xnor U641 (N_641,In_2441,In_1029);
or U642 (N_642,In_3240,In_2662);
or U643 (N_643,In_430,In_2517);
nand U644 (N_644,In_1291,In_3322);
or U645 (N_645,In_4730,In_1206);
and U646 (N_646,In_1396,In_1235);
xnor U647 (N_647,In_1647,In_2285);
or U648 (N_648,In_671,In_4341);
and U649 (N_649,In_880,In_4562);
or U650 (N_650,In_4203,In_3726);
nor U651 (N_651,In_3092,In_3992);
nand U652 (N_652,In_1926,In_4936);
nand U653 (N_653,In_2272,In_4443);
nand U654 (N_654,In_4602,N_116);
xor U655 (N_655,In_2465,In_3931);
nor U656 (N_656,In_2899,In_3097);
or U657 (N_657,In_3216,In_296);
nand U658 (N_658,In_4542,In_36);
and U659 (N_659,In_1894,In_4946);
nand U660 (N_660,In_2397,In_2479);
nor U661 (N_661,In_1967,In_1882);
and U662 (N_662,In_2935,In_4663);
and U663 (N_663,In_1479,N_331);
nor U664 (N_664,In_1140,In_2908);
xor U665 (N_665,In_189,In_462);
xnor U666 (N_666,In_1313,In_3576);
nand U667 (N_667,In_4958,In_2491);
nor U668 (N_668,In_3888,In_673);
xor U669 (N_669,In_3894,In_2677);
or U670 (N_670,In_3822,In_4543);
nand U671 (N_671,In_1673,In_317);
nor U672 (N_672,In_951,In_3367);
and U673 (N_673,In_4170,In_2673);
or U674 (N_674,In_807,In_102);
nor U675 (N_675,In_569,N_269);
xnor U676 (N_676,In_4534,In_1610);
and U677 (N_677,N_433,N_430);
and U678 (N_678,In_4221,In_2559);
or U679 (N_679,In_890,In_4778);
nand U680 (N_680,In_1794,In_3219);
and U681 (N_681,In_4704,In_3066);
nand U682 (N_682,In_3484,In_1539);
xnor U683 (N_683,In_710,In_2999);
and U684 (N_684,N_287,In_1365);
nand U685 (N_685,N_57,In_4703);
nor U686 (N_686,In_2087,In_3433);
xor U687 (N_687,N_338,In_1332);
nand U688 (N_688,In_2737,In_1577);
or U689 (N_689,In_169,In_1164);
nor U690 (N_690,In_3676,In_222);
nor U691 (N_691,In_2178,N_213);
xor U692 (N_692,In_1272,In_161);
and U693 (N_693,In_4363,In_3660);
and U694 (N_694,In_3435,In_2082);
xnor U695 (N_695,In_1712,In_1058);
or U696 (N_696,In_1055,In_4745);
xor U697 (N_697,In_2044,In_1069);
xnor U698 (N_698,In_495,In_3230);
and U699 (N_699,N_179,In_637);
nor U700 (N_700,In_428,In_1756);
or U701 (N_701,In_1600,In_410);
xor U702 (N_702,In_2471,In_917);
nand U703 (N_703,N_124,In_2358);
nand U704 (N_704,In_67,In_3290);
and U705 (N_705,In_1834,N_103);
nand U706 (N_706,In_4912,In_1986);
xor U707 (N_707,In_1471,In_2546);
nor U708 (N_708,In_2801,In_3832);
nand U709 (N_709,N_6,In_1387);
or U710 (N_710,N_78,In_2978);
nand U711 (N_711,In_1632,N_315);
or U712 (N_712,In_1447,In_3785);
nand U713 (N_713,In_2616,In_4096);
xor U714 (N_714,In_830,In_3657);
or U715 (N_715,In_55,In_1020);
and U716 (N_716,In_77,In_650);
nor U717 (N_717,In_4970,In_1060);
and U718 (N_718,In_892,In_1782);
nor U719 (N_719,In_1939,In_4486);
xnor U720 (N_720,In_3627,N_145);
nor U721 (N_721,In_1300,In_941);
or U722 (N_722,In_2722,In_1234);
nand U723 (N_723,In_1305,In_324);
nor U724 (N_724,In_2788,In_1381);
and U725 (N_725,In_3192,N_305);
nand U726 (N_726,In_2735,In_1052);
and U727 (N_727,In_1169,In_4346);
nand U728 (N_728,N_212,In_4758);
and U729 (N_729,In_4608,In_2825);
nor U730 (N_730,In_2857,In_3035);
or U731 (N_731,N_489,In_1195);
nand U732 (N_732,In_1751,In_4939);
nand U733 (N_733,In_1906,In_4090);
or U734 (N_734,In_4801,In_4786);
nand U735 (N_735,N_462,In_1947);
or U736 (N_736,N_483,In_327);
or U737 (N_737,In_3806,N_1);
nand U738 (N_738,In_2610,In_1822);
nand U739 (N_739,In_1118,N_11);
xor U740 (N_740,In_1949,In_1399);
and U741 (N_741,N_349,In_719);
xor U742 (N_742,N_359,In_4893);
or U743 (N_743,In_4683,N_292);
nor U744 (N_744,In_4999,In_2288);
nand U745 (N_745,In_4073,In_3291);
and U746 (N_746,N_99,In_3801);
or U747 (N_747,In_1024,N_281);
or U748 (N_748,In_2520,In_999);
nand U749 (N_749,In_3473,In_3606);
nor U750 (N_750,N_647,In_4039);
nor U751 (N_751,In_3146,N_231);
nor U752 (N_752,In_3929,In_2505);
nor U753 (N_753,In_4428,In_2273);
nand U754 (N_754,In_851,In_3048);
nor U755 (N_755,N_664,In_4871);
nand U756 (N_756,In_3100,In_368);
or U757 (N_757,N_668,N_356);
and U758 (N_758,In_466,In_4174);
nor U759 (N_759,In_1241,In_193);
and U760 (N_760,In_2514,In_2863);
or U761 (N_761,In_859,In_3537);
or U762 (N_762,In_2701,In_3007);
and U763 (N_763,In_3130,In_1716);
nor U764 (N_764,In_2490,In_2912);
and U765 (N_765,In_3085,N_313);
and U766 (N_766,In_2130,In_2819);
or U767 (N_767,N_193,In_2823);
or U768 (N_768,In_2039,N_541);
nor U769 (N_769,In_4106,In_2222);
xnor U770 (N_770,In_4490,In_4031);
xnor U771 (N_771,N_708,In_2355);
nand U772 (N_772,In_4932,N_311);
nor U773 (N_773,In_3966,In_4478);
nand U774 (N_774,In_4640,In_1932);
xnor U775 (N_775,N_663,N_186);
xor U776 (N_776,In_3611,In_3239);
and U777 (N_777,In_3615,In_2466);
or U778 (N_778,In_3734,In_2332);
and U779 (N_779,N_690,In_157);
and U780 (N_780,In_3675,In_3004);
and U781 (N_781,In_2979,In_4916);
nor U782 (N_782,N_610,In_1434);
or U783 (N_783,In_1033,In_3803);
nor U784 (N_784,In_2720,In_4361);
nor U785 (N_785,In_4751,N_709);
and U786 (N_786,In_606,In_3504);
nor U787 (N_787,N_132,In_1087);
xor U788 (N_788,In_2916,In_4539);
nand U789 (N_789,In_1643,In_570);
nand U790 (N_790,In_4347,In_1981);
or U791 (N_791,In_1764,In_4151);
nand U792 (N_792,In_3334,In_1331);
and U793 (N_793,In_4141,N_406);
xnor U794 (N_794,In_2955,In_454);
or U795 (N_795,In_3963,In_4549);
nand U796 (N_796,In_4220,In_2306);
or U797 (N_797,In_4485,In_2939);
and U798 (N_798,In_559,N_364);
xnor U799 (N_799,In_2362,In_3761);
or U800 (N_800,In_200,In_4982);
or U801 (N_801,N_73,N_733);
nand U802 (N_802,In_3740,N_487);
xor U803 (N_803,N_234,N_108);
xnor U804 (N_804,In_2754,In_2621);
xor U805 (N_805,In_1950,In_1612);
xor U806 (N_806,In_4216,In_2757);
xnor U807 (N_807,In_2866,N_366);
xor U808 (N_808,N_369,In_4924);
xor U809 (N_809,N_502,In_2395);
nor U810 (N_810,In_3286,In_4531);
and U811 (N_811,In_4582,In_821);
nor U812 (N_812,N_23,N_184);
or U813 (N_813,In_360,In_2030);
nand U814 (N_814,In_4026,In_4267);
and U815 (N_815,In_4411,In_612);
and U816 (N_816,In_1139,In_2209);
xnor U817 (N_817,In_2716,In_2305);
or U818 (N_818,In_205,In_3283);
and U819 (N_819,In_3152,In_1061);
and U820 (N_820,In_3256,In_173);
and U821 (N_821,N_562,In_1152);
nor U822 (N_822,N_140,In_4729);
or U823 (N_823,N_350,In_2877);
nor U824 (N_824,In_993,N_70);
nor U825 (N_825,N_511,In_4460);
xnor U826 (N_826,In_3386,In_2366);
nor U827 (N_827,In_1019,In_4165);
xor U828 (N_828,In_4053,In_2713);
nor U829 (N_829,In_2560,In_4068);
and U830 (N_830,In_2724,In_4798);
or U831 (N_831,In_2350,In_1257);
nand U832 (N_832,In_3423,In_2233);
and U833 (N_833,In_2817,In_960);
and U834 (N_834,In_107,In_3573);
and U835 (N_835,In_2211,In_1576);
and U836 (N_836,In_1752,In_2093);
and U837 (N_837,In_2009,In_3775);
xor U838 (N_838,In_22,In_3511);
nor U839 (N_839,In_4604,In_1701);
or U840 (N_840,In_4160,In_2160);
and U841 (N_841,In_997,In_1973);
and U842 (N_842,In_2968,In_3427);
and U843 (N_843,In_978,In_4097);
nor U844 (N_844,N_343,In_1706);
xor U845 (N_845,In_1900,In_4011);
and U846 (N_846,In_1559,In_2541);
nor U847 (N_847,In_3968,In_2302);
or U848 (N_848,In_2141,In_4739);
or U849 (N_849,In_2914,In_3804);
or U850 (N_850,In_407,In_1901);
nor U851 (N_851,In_3460,In_827);
and U852 (N_852,In_319,In_235);
xnor U853 (N_853,In_208,In_793);
and U854 (N_854,In_4093,In_4718);
and U855 (N_855,In_4540,In_3771);
or U856 (N_856,In_4779,In_330);
and U857 (N_857,In_2428,In_577);
nand U858 (N_858,In_3251,In_648);
nand U859 (N_859,In_2151,In_3134);
xor U860 (N_860,N_679,In_4444);
nand U861 (N_861,In_1984,In_315);
nor U862 (N_862,In_1494,In_3877);
nor U863 (N_863,N_172,In_3056);
or U864 (N_864,In_4585,In_3700);
and U865 (N_865,In_725,In_3250);
xor U866 (N_866,In_3430,In_1282);
nand U867 (N_867,In_1338,In_677);
or U868 (N_868,In_3975,In_4826);
xor U869 (N_869,In_668,N_648);
or U870 (N_870,In_3812,N_494);
and U871 (N_871,In_2037,In_3150);
and U872 (N_872,In_4769,N_178);
or U873 (N_873,N_297,In_1082);
or U874 (N_874,In_4020,N_310);
nand U875 (N_875,In_1943,N_660);
or U876 (N_876,N_605,In_127);
nor U877 (N_877,In_1124,In_2562);
xnor U878 (N_878,In_2115,In_2122);
nand U879 (N_879,In_1942,In_654);
nor U880 (N_880,In_682,In_82);
xnor U881 (N_881,In_266,In_1039);
nor U882 (N_882,In_1725,N_180);
nor U883 (N_883,N_680,In_4499);
nor U884 (N_884,In_2885,N_165);
nand U885 (N_885,In_2586,N_312);
or U886 (N_886,In_1797,In_3893);
and U887 (N_887,N_558,In_3671);
nand U888 (N_888,In_1276,N_522);
nand U889 (N_889,In_3730,N_173);
nor U890 (N_890,In_3381,In_4680);
xnor U891 (N_891,N_236,In_2167);
or U892 (N_892,In_342,In_1719);
or U893 (N_893,N_201,In_534);
xor U894 (N_894,In_3308,In_4847);
or U895 (N_895,In_3815,In_281);
nand U896 (N_896,N_329,In_1483);
xor U897 (N_897,In_3264,In_1538);
nand U898 (N_898,In_2276,In_4860);
nand U899 (N_899,In_3792,In_2789);
nand U900 (N_900,N_24,In_1217);
nor U901 (N_901,In_2897,N_561);
or U902 (N_902,In_2934,In_932);
or U903 (N_903,In_358,In_4599);
xnor U904 (N_904,In_2601,In_4416);
nor U905 (N_905,In_1173,In_283);
nor U906 (N_906,In_2499,In_1346);
or U907 (N_907,In_1075,In_1427);
or U908 (N_908,In_3733,In_3390);
and U909 (N_909,In_139,In_4084);
nand U910 (N_910,In_1414,In_1761);
nor U911 (N_911,N_594,N_670);
nand U912 (N_912,N_174,In_3340);
and U913 (N_913,In_3678,In_1504);
nand U914 (N_914,In_4023,In_2451);
or U915 (N_915,In_1688,In_2038);
xnor U916 (N_916,In_3996,In_2575);
xor U917 (N_917,In_4564,In_323);
xor U918 (N_918,In_3144,In_442);
nand U919 (N_919,N_699,In_174);
xnor U920 (N_920,N_582,In_757);
nand U921 (N_921,In_659,In_4571);
and U922 (N_922,In_3518,In_3835);
nand U923 (N_923,In_1832,In_4906);
xnor U924 (N_924,In_1955,In_2544);
xnor U925 (N_925,In_2008,In_4315);
or U926 (N_926,In_3842,In_3829);
nor U927 (N_927,In_3981,N_251);
nand U928 (N_928,In_4833,In_3019);
nor U929 (N_929,In_3148,In_3945);
nand U930 (N_930,In_426,In_1814);
nor U931 (N_931,In_2555,In_3431);
xor U932 (N_932,In_4261,N_456);
nand U933 (N_933,In_1865,In_3461);
and U934 (N_934,In_4058,In_835);
nand U935 (N_935,In_638,In_3623);
or U936 (N_936,In_2254,In_108);
or U937 (N_937,In_1699,In_320);
and U938 (N_938,In_3015,In_96);
xor U939 (N_939,In_2077,In_2507);
nor U940 (N_940,In_1992,In_4748);
nand U941 (N_941,In_751,In_3458);
or U942 (N_942,In_1839,In_1146);
nand U943 (N_943,In_3749,N_613);
or U944 (N_944,In_4611,In_366);
xnor U945 (N_945,In_1598,In_403);
nor U946 (N_946,In_2623,In_3610);
nor U947 (N_947,In_4371,N_68);
and U948 (N_948,N_630,N_221);
and U949 (N_949,In_4787,In_137);
nor U950 (N_950,In_4177,In_1076);
nand U951 (N_951,In_4364,In_3113);
and U952 (N_952,In_1230,In_3018);
xor U953 (N_953,In_1105,In_2976);
xnor U954 (N_954,In_2147,In_4978);
nand U955 (N_955,N_409,In_3707);
or U956 (N_956,In_1209,In_424);
or U957 (N_957,In_1375,N_121);
nor U958 (N_958,In_2637,In_4184);
nor U959 (N_959,In_2965,In_1583);
or U960 (N_960,In_418,N_143);
and U961 (N_961,In_2301,In_4795);
or U962 (N_962,N_469,In_1666);
nor U963 (N_963,In_2161,N_379);
nand U964 (N_964,In_4918,N_158);
xnor U965 (N_965,N_644,In_1085);
and U966 (N_966,In_4782,In_4709);
nor U967 (N_967,In_2692,In_2760);
and U968 (N_968,N_543,In_3862);
and U969 (N_969,N_700,In_2368);
nor U970 (N_970,In_3970,In_601);
and U971 (N_971,In_1614,In_4375);
or U972 (N_972,In_1791,N_632);
xor U973 (N_973,In_4459,In_4516);
or U974 (N_974,In_1728,In_4857);
xor U975 (N_975,In_226,In_3778);
or U976 (N_976,In_3595,In_3364);
nor U977 (N_977,In_3885,In_2629);
and U978 (N_978,In_683,In_3221);
and U979 (N_979,N_667,In_1622);
or U980 (N_980,In_1574,In_4954);
and U981 (N_981,N_275,In_365);
or U982 (N_982,In_1616,N_245);
and U983 (N_983,In_394,In_2688);
and U984 (N_984,In_2431,In_2846);
xor U985 (N_985,In_1095,In_4289);
and U986 (N_986,In_4114,N_353);
and U987 (N_987,In_2074,In_1354);
xnor U988 (N_988,In_457,In_1911);
xor U989 (N_989,In_1534,In_4512);
nand U990 (N_990,N_224,In_286);
xor U991 (N_991,In_3613,In_4163);
xnor U992 (N_992,In_2359,In_1924);
nand U993 (N_993,In_3017,In_3631);
nor U994 (N_994,N_7,In_885);
xnor U995 (N_995,In_3529,In_1172);
and U996 (N_996,In_3275,In_4178);
and U997 (N_997,In_772,In_1858);
xor U998 (N_998,In_1148,In_4913);
xor U999 (N_999,In_2426,In_4113);
xor U1000 (N_1000,In_1424,In_1347);
xor U1001 (N_1001,In_526,In_2518);
nor U1002 (N_1002,In_1569,In_1637);
or U1003 (N_1003,In_3151,N_937);
nor U1004 (N_1004,In_1402,In_251);
xnor U1005 (N_1005,In_1032,N_268);
or U1006 (N_1006,In_1802,N_723);
nand U1007 (N_1007,In_2663,In_3452);
and U1008 (N_1008,N_290,N_546);
nor U1009 (N_1009,In_3369,In_1560);
nand U1010 (N_1010,N_237,In_1443);
xor U1011 (N_1011,In_599,In_2155);
nor U1012 (N_1012,N_633,In_1207);
xor U1013 (N_1013,In_4981,In_2802);
or U1014 (N_1014,In_2527,In_1793);
nor U1015 (N_1015,N_113,In_2001);
and U1016 (N_1016,In_647,In_3499);
or U1017 (N_1017,In_2855,In_4693);
and U1018 (N_1018,In_2751,In_2142);
nand U1019 (N_1019,In_1191,In_1769);
nand U1020 (N_1020,In_4017,N_39);
or U1021 (N_1021,In_2478,In_3752);
and U1022 (N_1022,In_2392,N_98);
and U1023 (N_1023,In_384,N_878);
nor U1024 (N_1024,N_981,In_3580);
nand U1025 (N_1025,In_2411,N_615);
nor U1026 (N_1026,In_2291,In_666);
or U1027 (N_1027,In_3746,In_1659);
nand U1028 (N_1028,N_741,N_898);
and U1029 (N_1029,N_246,N_710);
or U1030 (N_1030,In_3638,In_1807);
nand U1031 (N_1031,N_773,In_776);
and U1032 (N_1032,In_4768,In_4239);
or U1033 (N_1033,N_398,In_4747);
xor U1034 (N_1034,In_4061,In_117);
nand U1035 (N_1035,In_4336,In_1988);
or U1036 (N_1036,N_464,In_3391);
nand U1037 (N_1037,In_1360,In_311);
xnor U1038 (N_1038,In_1394,In_2587);
xnor U1039 (N_1039,In_1388,N_387);
or U1040 (N_1040,In_143,In_2848);
or U1041 (N_1041,In_1898,In_2756);
nand U1042 (N_1042,In_116,In_1975);
nor U1043 (N_1043,In_867,In_1430);
nor U1044 (N_1044,In_1158,In_3609);
nand U1045 (N_1045,In_1921,In_3711);
nand U1046 (N_1046,In_2915,In_2774);
nand U1047 (N_1047,N_716,N_592);
nor U1048 (N_1048,In_413,In_1963);
or U1049 (N_1049,In_3920,In_943);
nor U1050 (N_1050,In_4903,In_4919);
and U1051 (N_1051,In_4201,In_2188);
nand U1052 (N_1052,In_596,In_445);
or U1053 (N_1053,In_546,In_4192);
and U1054 (N_1054,In_2550,In_1177);
nand U1055 (N_1055,In_322,In_395);
or U1056 (N_1056,In_4712,In_2557);
nand U1057 (N_1057,In_1521,N_646);
nand U1058 (N_1058,In_3978,In_3321);
xor U1059 (N_1059,In_2425,In_3656);
nor U1060 (N_1060,In_3402,In_1138);
nor U1061 (N_1061,In_3220,N_659);
nor U1062 (N_1062,In_4279,In_2681);
and U1063 (N_1063,In_1852,In_111);
or U1064 (N_1064,In_70,N_61);
or U1065 (N_1065,In_4120,In_631);
xor U1066 (N_1066,In_2871,In_3375);
nor U1067 (N_1067,In_939,N_617);
or U1068 (N_1068,In_2228,In_4872);
nand U1069 (N_1069,In_2488,In_455);
nor U1070 (N_1070,In_1547,In_1776);
and U1071 (N_1071,In_3288,N_301);
and U1072 (N_1072,In_4726,In_4441);
and U1073 (N_1073,N_131,N_941);
xnor U1074 (N_1074,N_450,N_890);
xnor U1075 (N_1075,In_3023,In_49);
nand U1076 (N_1076,In_4210,N_587);
nand U1077 (N_1077,In_292,In_4193);
nor U1078 (N_1078,In_1972,N_611);
and U1079 (N_1079,In_2769,In_4578);
nand U1080 (N_1080,In_79,In_3160);
or U1081 (N_1081,In_1572,In_3982);
and U1082 (N_1082,N_62,In_4377);
nor U1083 (N_1083,In_842,In_2388);
and U1084 (N_1084,N_706,In_123);
or U1085 (N_1085,In_1844,In_4993);
and U1086 (N_1086,In_4628,In_4655);
and U1087 (N_1087,In_3229,N_362);
nand U1088 (N_1088,In_1520,In_2783);
xnor U1089 (N_1089,In_1003,In_3764);
and U1090 (N_1090,In_2282,In_1996);
or U1091 (N_1091,In_2895,In_4248);
or U1092 (N_1092,In_3136,In_4699);
xor U1093 (N_1093,N_577,In_1768);
nor U1094 (N_1094,N_92,In_4077);
or U1095 (N_1095,N_19,In_2257);
or U1096 (N_1096,In_4025,In_60);
and U1097 (N_1097,N_141,In_197);
nor U1098 (N_1098,In_4592,In_3124);
nand U1099 (N_1099,In_209,In_523);
nor U1100 (N_1100,N_977,N_316);
and U1101 (N_1101,In_1682,In_443);
nor U1102 (N_1102,In_1775,In_4134);
or U1103 (N_1103,In_6,In_4933);
nor U1104 (N_1104,In_3071,In_4994);
xor U1105 (N_1105,In_583,In_1198);
nor U1106 (N_1106,In_3589,N_378);
or U1107 (N_1107,N_365,In_4067);
xnor U1108 (N_1108,In_4668,N_846);
nor U1109 (N_1109,N_556,In_1856);
nor U1110 (N_1110,In_1535,In_4500);
and U1111 (N_1111,In_4111,In_2738);
nand U1112 (N_1112,In_3779,In_3006);
and U1113 (N_1113,In_2591,N_192);
nor U1114 (N_1114,N_203,In_4990);
and U1115 (N_1115,In_744,In_1624);
nor U1116 (N_1116,In_129,N_342);
nand U1117 (N_1117,In_2504,In_1759);
nand U1118 (N_1118,In_3409,In_4318);
and U1119 (N_1119,N_868,In_2628);
and U1120 (N_1120,N_721,In_2919);
and U1121 (N_1121,In_2954,In_841);
nand U1122 (N_1122,In_4019,In_414);
nand U1123 (N_1123,N_418,In_1457);
nor U1124 (N_1124,N_395,In_4904);
nand U1125 (N_1125,In_746,N_956);
or U1126 (N_1126,In_1137,In_2054);
and U1127 (N_1127,In_994,In_2390);
and U1128 (N_1128,In_1096,N_643);
or U1129 (N_1129,In_3462,In_2890);
and U1130 (N_1130,In_856,N_992);
and U1131 (N_1131,N_528,N_177);
or U1132 (N_1132,In_872,In_219);
or U1133 (N_1133,In_2632,N_820);
nor U1134 (N_1134,In_1745,In_3650);
nand U1135 (N_1135,In_42,In_1540);
nor U1136 (N_1136,In_3594,In_4856);
nand U1137 (N_1137,In_2932,In_1717);
xnor U1138 (N_1138,In_3129,In_3190);
xnor U1139 (N_1139,In_4977,In_1278);
nand U1140 (N_1140,In_3393,In_2820);
xor U1141 (N_1141,N_135,In_4719);
nor U1142 (N_1142,In_860,N_677);
xnor U1143 (N_1143,In_1875,In_1561);
or U1144 (N_1144,In_124,In_2317);
xor U1145 (N_1145,N_926,In_4887);
or U1146 (N_1146,In_1189,In_2405);
nor U1147 (N_1147,N_597,In_4561);
or U1148 (N_1148,In_3131,N_832);
or U1149 (N_1149,In_3154,N_497);
nor U1150 (N_1150,N_373,In_3269);
xnor U1151 (N_1151,In_3957,In_4710);
and U1152 (N_1152,In_4521,In_2892);
xor U1153 (N_1153,In_4101,In_2320);
and U1154 (N_1154,In_3543,N_300);
nand U1155 (N_1155,In_2578,N_640);
xor U1156 (N_1156,In_2661,In_3930);
nor U1157 (N_1157,In_2379,In_902);
nor U1158 (N_1158,In_110,In_4849);
or U1159 (N_1159,In_213,In_3759);
nand U1160 (N_1160,N_636,In_3331);
or U1161 (N_1161,In_3682,In_4181);
or U1162 (N_1162,In_864,N_518);
or U1163 (N_1163,In_1218,In_1262);
and U1164 (N_1164,In_693,In_3318);
nor U1165 (N_1165,In_362,N_603);
xor U1166 (N_1166,In_4245,In_239);
nor U1167 (N_1167,In_121,In_983);
and U1168 (N_1168,In_291,In_4446);
nor U1169 (N_1169,In_1861,N_533);
nand U1170 (N_1170,In_4494,In_3432);
xor U1171 (N_1171,In_838,In_4454);
or U1172 (N_1172,In_769,In_1312);
or U1173 (N_1173,In_4083,In_2858);
nand U1174 (N_1174,In_4793,In_1212);
nor U1175 (N_1175,In_1824,In_3643);
nand U1176 (N_1176,In_423,In_2509);
xnor U1177 (N_1177,In_4110,In_3089);
or U1178 (N_1178,In_1642,In_845);
nor U1179 (N_1179,In_254,In_2224);
nand U1180 (N_1180,In_3583,In_4821);
or U1181 (N_1181,In_4880,N_560);
nand U1182 (N_1182,In_957,In_1181);
or U1183 (N_1183,In_3670,N_56);
nor U1184 (N_1184,In_980,In_2007);
and U1185 (N_1185,In_4877,In_3438);
and U1186 (N_1186,N_424,N_844);
xor U1187 (N_1187,In_1321,In_1805);
nand U1188 (N_1188,In_4722,In_3197);
or U1189 (N_1189,In_3624,In_4529);
and U1190 (N_1190,In_259,N_814);
or U1191 (N_1191,In_1897,N_872);
nand U1192 (N_1192,In_1748,In_4945);
nor U1193 (N_1193,In_4362,In_4452);
xor U1194 (N_1194,N_802,In_1275);
nand U1195 (N_1195,In_3653,In_3060);
xor U1196 (N_1196,In_620,In_1958);
or U1197 (N_1197,In_1804,In_3834);
nand U1198 (N_1198,N_564,In_3359);
xnor U1199 (N_1199,In_4692,N_698);
nor U1200 (N_1200,N_589,N_410);
or U1201 (N_1201,In_2484,N_711);
xor U1202 (N_1202,N_382,In_3993);
nor U1203 (N_1203,In_4998,In_440);
and U1204 (N_1204,In_4234,In_2533);
nor U1205 (N_1205,In_4537,N_440);
and U1206 (N_1206,In_1336,In_4902);
nand U1207 (N_1207,In_1150,In_2132);
nor U1208 (N_1208,In_652,In_3574);
nor U1209 (N_1209,N_163,N_332);
nand U1210 (N_1210,In_3816,N_282);
xnor U1211 (N_1211,In_3125,In_4422);
or U1212 (N_1212,In_706,N_675);
or U1213 (N_1213,In_1122,In_3701);
nand U1214 (N_1214,N_460,N_634);
nor U1215 (N_1215,In_4173,In_1670);
and U1216 (N_1216,In_3807,In_3396);
xor U1217 (N_1217,In_476,In_1353);
xnor U1218 (N_1218,In_4839,In_4373);
nand U1219 (N_1219,In_1009,In_1720);
nor U1220 (N_1220,In_3140,In_2261);
xor U1221 (N_1221,In_1442,In_1771);
xnor U1222 (N_1222,In_1536,In_3314);
and U1223 (N_1223,In_2889,In_146);
and U1224 (N_1224,In_1525,In_1329);
nor U1225 (N_1225,In_3777,N_330);
or U1226 (N_1226,N_93,In_732);
nor U1227 (N_1227,In_4049,In_4964);
xor U1228 (N_1228,In_2950,In_3848);
nor U1229 (N_1229,N_599,N_319);
nand U1230 (N_1230,In_2945,In_1570);
xor U1231 (N_1231,N_914,In_1091);
and U1232 (N_1232,In_2225,In_2497);
xnor U1233 (N_1233,In_3031,In_2928);
nand U1234 (N_1234,N_899,In_3196);
nor U1235 (N_1235,N_567,In_4302);
and U1236 (N_1236,In_1833,In_412);
nor U1237 (N_1237,In_3237,In_1253);
or U1238 (N_1238,In_4233,In_4232);
nor U1239 (N_1239,In_2123,In_422);
or U1240 (N_1240,In_1607,In_4231);
and U1241 (N_1241,N_763,In_3874);
nand U1242 (N_1242,In_513,In_2723);
nor U1243 (N_1243,In_2445,In_2119);
nand U1244 (N_1244,In_1433,In_2849);
nand U1245 (N_1245,In_2407,N_189);
or U1246 (N_1246,N_170,N_323);
and U1247 (N_1247,N_935,In_4436);
xnor U1248 (N_1248,In_4968,In_624);
nor U1249 (N_1249,In_3561,N_815);
nor U1250 (N_1250,N_505,In_2279);
xor U1251 (N_1251,In_3686,In_4194);
and U1252 (N_1252,In_188,In_481);
and U1253 (N_1253,In_155,N_1013);
nor U1254 (N_1254,N_1136,N_1124);
nand U1255 (N_1255,In_2343,N_1112);
nor U1256 (N_1256,In_4684,In_3725);
nand U1257 (N_1257,In_3723,In_4332);
nor U1258 (N_1258,In_3343,In_3232);
xnor U1259 (N_1259,In_3496,In_742);
nand U1260 (N_1260,N_355,N_13);
xnor U1261 (N_1261,N_485,In_4189);
or U1262 (N_1262,In_734,N_333);
xor U1263 (N_1263,N_965,In_1498);
or U1264 (N_1264,In_512,In_4734);
xnor U1265 (N_1265,N_35,N_417);
and U1266 (N_1266,In_1439,In_4612);
nor U1267 (N_1267,In_801,In_1130);
nor U1268 (N_1268,In_211,In_3789);
nand U1269 (N_1269,In_2538,In_4018);
xnor U1270 (N_1270,In_1944,N_375);
or U1271 (N_1271,In_3531,N_1198);
xnor U1272 (N_1272,In_4236,In_3539);
nor U1273 (N_1273,In_3505,In_3176);
nor U1274 (N_1274,In_2292,In_2297);
nor U1275 (N_1275,N_318,In_2031);
and U1276 (N_1276,N_960,In_3330);
nor U1277 (N_1277,N_1159,N_1130);
xor U1278 (N_1278,In_2460,In_3149);
nand U1279 (N_1279,In_1683,N_787);
nand U1280 (N_1280,In_2510,In_1916);
or U1281 (N_1281,In_4464,In_2967);
and U1282 (N_1282,In_1073,In_1348);
xor U1283 (N_1283,In_2485,N_380);
or U1284 (N_1284,In_670,In_2281);
xnor U1285 (N_1285,N_606,In_4176);
nand U1286 (N_1286,In_2290,In_1866);
xor U1287 (N_1287,In_808,In_4665);
or U1288 (N_1288,In_3540,In_4471);
or U1289 (N_1289,N_737,In_3456);
nand U1290 (N_1290,N_381,N_980);
nand U1291 (N_1291,N_671,In_1790);
nor U1292 (N_1292,In_1151,In_4679);
nor U1293 (N_1293,In_4280,In_1733);
xnor U1294 (N_1294,In_3467,In_4807);
nand U1295 (N_1295,In_3662,In_4750);
or U1296 (N_1296,N_747,N_414);
or U1297 (N_1297,In_3868,In_4226);
nor U1298 (N_1298,In_4281,In_3654);
nor U1299 (N_1299,In_2120,N_182);
or U1300 (N_1300,In_651,In_2474);
and U1301 (N_1301,In_2470,In_1448);
or U1302 (N_1302,N_795,N_962);
or U1303 (N_1303,In_2614,In_2168);
nor U1304 (N_1304,In_1989,In_2144);
or U1305 (N_1305,In_285,In_2442);
nand U1306 (N_1306,In_1795,In_1801);
xnor U1307 (N_1307,In_709,In_1256);
nor U1308 (N_1308,In_4836,N_109);
and U1309 (N_1309,In_265,In_132);
and U1310 (N_1310,In_2062,In_1915);
and U1311 (N_1311,N_655,In_669);
or U1312 (N_1312,In_4218,N_337);
or U1313 (N_1313,N_530,In_785);
nand U1314 (N_1314,N_481,In_3082);
and U1315 (N_1315,In_2516,N_136);
and U1316 (N_1316,In_4789,In_1363);
nor U1317 (N_1317,N_1062,N_1220);
and U1318 (N_1318,In_771,In_255);
and U1319 (N_1319,In_3939,In_4563);
and U1320 (N_1320,N_32,In_2482);
or U1321 (N_1321,N_705,N_691);
or U1322 (N_1322,In_1392,In_3413);
and U1323 (N_1323,In_4850,In_25);
nand U1324 (N_1324,In_722,In_4322);
or U1325 (N_1325,N_125,In_112);
xnor U1326 (N_1326,In_4686,In_3689);
or U1327 (N_1327,In_1606,In_2991);
or U1328 (N_1328,N_909,In_284);
nor U1329 (N_1329,N_727,N_999);
or U1330 (N_1330,In_2695,In_1993);
or U1331 (N_1331,In_4225,N_1123);
nand U1332 (N_1332,In_1044,In_530);
and U1333 (N_1333,In_3845,In_3924);
nand U1334 (N_1334,In_3349,In_4895);
and U1335 (N_1335,In_4901,In_314);
or U1336 (N_1336,N_696,N_1025);
nand U1337 (N_1337,In_4468,In_861);
or U1338 (N_1338,N_161,N_1175);
and U1339 (N_1339,In_1089,In_4570);
and U1340 (N_1340,In_2548,In_1333);
xnor U1341 (N_1341,In_4152,In_2058);
or U1342 (N_1342,In_1578,In_4082);
and U1343 (N_1343,In_1508,In_3585);
xor U1344 (N_1344,N_1235,In_3795);
and U1345 (N_1345,In_3958,N_59);
xor U1346 (N_1346,N_749,N_923);
nand U1347 (N_1347,In_1093,In_1327);
nand U1348 (N_1348,In_1441,N_1082);
and U1349 (N_1349,In_515,In_489);
or U1350 (N_1350,In_1469,In_4997);
nor U1351 (N_1351,N_591,N_973);
or U1352 (N_1352,In_3249,In_1214);
xnor U1353 (N_1353,In_927,In_2299);
nand U1354 (N_1354,N_1133,N_880);
or U1355 (N_1355,N_1033,In_2469);
and U1356 (N_1356,In_3394,N_1214);
nor U1357 (N_1357,In_2535,In_1489);
xor U1358 (N_1358,In_3418,N_654);
nand U1359 (N_1359,In_3553,N_637);
nand U1360 (N_1360,In_3439,In_2602);
nor U1361 (N_1361,N_1150,In_3405);
or U1362 (N_1362,N_419,In_4818);
and U1363 (N_1363,N_447,N_1017);
or U1364 (N_1364,N_524,In_1432);
and U1365 (N_1365,In_4144,In_247);
xnor U1366 (N_1366,In_4118,In_3078);
nor U1367 (N_1367,N_523,In_372);
nor U1368 (N_1368,In_1913,In_4817);
xor U1369 (N_1369,In_505,In_3127);
nand U1370 (N_1370,In_547,In_563);
xor U1371 (N_1371,In_3665,In_4156);
or U1372 (N_1372,In_1687,N_239);
or U1373 (N_1373,In_3161,N_1212);
and U1374 (N_1374,In_4333,In_4290);
xor U1375 (N_1375,In_1589,In_2399);
nor U1376 (N_1376,In_4581,In_4547);
or U1377 (N_1377,In_4858,In_4762);
nor U1378 (N_1378,In_3677,In_310);
and U1379 (N_1379,In_1112,N_51);
nand U1380 (N_1380,N_247,In_1786);
or U1381 (N_1381,In_3287,N_656);
xnor U1382 (N_1382,In_3267,N_401);
and U1383 (N_1383,In_2521,In_214);
and U1384 (N_1384,N_1230,In_4453);
nand U1385 (N_1385,In_558,In_2006);
xor U1386 (N_1386,In_2330,In_1828);
or U1387 (N_1387,N_1016,N_936);
or U1388 (N_1388,N_15,N_1249);
and U1389 (N_1389,In_328,In_3694);
nand U1390 (N_1390,N_286,In_4044);
nor U1391 (N_1391,In_114,In_1449);
or U1392 (N_1392,N_254,In_3175);
nand U1393 (N_1393,N_1005,N_824);
xnor U1394 (N_1394,In_100,In_1226);
xor U1395 (N_1395,In_3245,In_4530);
nor U1396 (N_1396,N_887,In_4752);
nand U1397 (N_1397,N_46,In_866);
nor U1398 (N_1398,N_344,In_2076);
and U1399 (N_1399,In_2612,In_1825);
nor U1400 (N_1400,In_258,In_4596);
xor U1401 (N_1401,In_1677,In_1532);
or U1402 (N_1402,In_3000,In_2639);
or U1403 (N_1403,In_2549,In_2667);
nor U1404 (N_1404,In_686,In_4451);
nand U1405 (N_1405,In_3642,In_1545);
and U1406 (N_1406,In_1123,In_4415);
nor U1407 (N_1407,N_537,N_578);
nand U1408 (N_1408,In_525,N_129);
xnor U1409 (N_1409,In_367,In_2792);
xnor U1410 (N_1410,In_545,In_175);
nor U1411 (N_1411,In_3578,N_991);
or U1412 (N_1412,In_3116,N_104);
xnor U1413 (N_1413,In_359,In_4435);
or U1414 (N_1414,N_222,In_278);
xnor U1415 (N_1415,In_1240,N_507);
and U1416 (N_1416,In_135,N_805);
nand U1417 (N_1417,N_809,In_2440);
nor U1418 (N_1418,In_2435,In_3542);
or U1419 (N_1419,In_3472,In_2201);
or U1420 (N_1420,In_2821,In_1244);
nor U1421 (N_1421,In_1474,In_3159);
nand U1422 (N_1422,In_924,N_208);
nor U1423 (N_1423,In_1524,In_3794);
and U1424 (N_1424,N_590,In_2923);
or U1425 (N_1425,In_1957,In_700);
xor U1426 (N_1426,N_922,In_166);
nor U1427 (N_1427,In_3951,N_862);
or U1428 (N_1428,In_257,In_4149);
or U1429 (N_1429,N_1056,In_712);
nor U1430 (N_1430,N_1020,In_3027);
and U1431 (N_1431,In_2900,In_2990);
nor U1432 (N_1432,In_2468,N_566);
nand U1433 (N_1433,In_3102,In_3408);
nand U1434 (N_1434,N_1120,In_65);
xnor U1435 (N_1435,N_34,In_522);
and U1436 (N_1436,In_4054,In_4224);
nand U1437 (N_1437,N_952,In_2960);
xor U1438 (N_1438,N_67,In_216);
or U1439 (N_1439,In_4614,In_4972);
xnor U1440 (N_1440,In_4394,In_417);
or U1441 (N_1441,N_285,In_3647);
nand U1442 (N_1442,In_4629,In_1783);
nand U1443 (N_1443,In_2072,In_4935);
or U1444 (N_1444,In_3304,In_32);
nand U1445 (N_1445,In_31,N_1149);
nand U1446 (N_1446,In_2462,In_1222);
nand U1447 (N_1447,In_811,In_2962);
nand U1448 (N_1448,In_2711,In_3821);
and U1449 (N_1449,N_864,In_782);
nand U1450 (N_1450,In_919,In_995);
nand U1451 (N_1451,In_528,In_2056);
nand U1452 (N_1452,N_1051,In_2294);
or U1453 (N_1453,In_3122,In_604);
and U1454 (N_1454,In_4405,In_4509);
nand U1455 (N_1455,In_253,In_1985);
xnor U1456 (N_1456,In_2552,In_716);
nor U1457 (N_1457,In_4182,In_354);
and U1458 (N_1458,In_2985,In_697);
or U1459 (N_1459,In_408,In_335);
or U1460 (N_1460,In_529,In_791);
or U1461 (N_1461,N_1068,In_2433);
nand U1462 (N_1462,In_104,In_2190);
or U1463 (N_1463,N_397,In_4202);
or U1464 (N_1464,N_303,In_1960);
nand U1465 (N_1465,N_474,N_263);
and U1466 (N_1466,N_1145,In_3301);
nand U1467 (N_1467,In_1809,In_4035);
nor U1468 (N_1468,In_3191,In_4166);
nor U1469 (N_1469,In_1874,In_685);
nand U1470 (N_1470,In_2594,In_352);
nor U1471 (N_1471,In_4510,In_4524);
nor U1472 (N_1472,N_848,In_1727);
nor U1473 (N_1473,In_4119,In_1090);
nor U1474 (N_1474,In_598,In_1264);
xnor U1475 (N_1475,In_4228,N_43);
or U1476 (N_1476,In_140,N_432);
or U1477 (N_1477,N_674,In_2709);
nand U1478 (N_1478,N_835,In_3088);
and U1479 (N_1479,In_3750,N_264);
nor U1480 (N_1480,In_2203,In_3155);
xor U1481 (N_1481,In_4142,In_295);
and U1482 (N_1482,N_470,In_4985);
and U1483 (N_1483,In_4861,In_496);
and U1484 (N_1484,In_1344,In_2198);
nor U1485 (N_1485,In_2360,N_525);
nand U1486 (N_1486,In_1512,In_775);
nor U1487 (N_1487,In_2384,In_4342);
and U1488 (N_1488,N_1190,N_953);
and U1489 (N_1489,In_876,In_2786);
xor U1490 (N_1490,In_2196,In_2731);
xnor U1491 (N_1491,In_1892,In_1515);
or U1492 (N_1492,In_3717,In_3008);
or U1493 (N_1493,N_84,N_693);
or U1494 (N_1494,In_350,N_328);
xor U1495 (N_1495,N_1233,In_3295);
xor U1496 (N_1496,In_1328,N_457);
xnor U1497 (N_1497,In_3754,In_3824);
and U1498 (N_1498,In_1908,N_886);
or U1499 (N_1499,In_1459,In_1544);
nor U1500 (N_1500,In_4929,N_881);
xnor U1501 (N_1501,In_2931,In_707);
nand U1502 (N_1502,N_753,In_2869);
or U1503 (N_1503,N_720,In_4222);
or U1504 (N_1504,In_4701,In_4127);
or U1505 (N_1505,N_476,In_3234);
or U1506 (N_1506,N_449,In_2679);
nand U1507 (N_1507,In_3776,In_4890);
or U1508 (N_1508,In_3588,In_1567);
xnor U1509 (N_1509,In_4527,In_4514);
or U1510 (N_1510,In_4278,In_2581);
xnor U1511 (N_1511,In_2676,In_3272);
xnor U1512 (N_1512,In_4891,N_291);
or U1513 (N_1513,N_1268,In_1934);
xnor U1514 (N_1514,In_1183,In_483);
and U1515 (N_1515,N_422,In_2942);
nor U1516 (N_1516,In_4423,In_4723);
or U1517 (N_1517,N_944,In_3509);
nor U1518 (N_1518,In_4742,In_4140);
or U1519 (N_1519,In_4761,In_282);
nor U1520 (N_1520,In_3266,In_1777);
nand U1521 (N_1521,In_3118,N_1323);
or U1522 (N_1522,In_4147,In_2088);
nor U1523 (N_1523,In_4938,In_1298);
nand U1524 (N_1524,N_219,In_541);
or U1525 (N_1525,In_1379,In_1490);
nor U1526 (N_1526,N_1216,In_2512);
and U1527 (N_1527,In_4944,In_4136);
or U1528 (N_1528,N_1247,In_103);
nand U1529 (N_1529,In_4105,In_981);
or U1530 (N_1530,In_3416,In_1136);
or U1531 (N_1531,In_3709,In_948);
and U1532 (N_1532,In_2267,In_3967);
nor U1533 (N_1533,In_4298,N_1097);
nand U1534 (N_1534,N_681,N_1483);
or U1535 (N_1535,In_2422,In_1308);
and U1536 (N_1536,In_2929,In_1665);
or U1537 (N_1537,In_2029,N_954);
nor U1538 (N_1538,N_216,In_2117);
nor U1539 (N_1539,In_1626,In_2734);
and U1540 (N_1540,In_1248,N_454);
nand U1541 (N_1541,N_1105,N_53);
or U1542 (N_1542,In_131,In_3258);
and U1543 (N_1543,In_3253,In_4397);
and U1544 (N_1544,In_4032,In_2243);
xnor U1545 (N_1545,N_1434,In_2472);
and U1546 (N_1546,In_1435,In_1021);
and U1547 (N_1547,In_377,N_436);
or U1548 (N_1548,N_1070,N_65);
xor U1549 (N_1549,N_341,In_2969);
nand U1550 (N_1550,In_2020,N_534);
or U1551 (N_1551,N_822,N_1425);
xor U1552 (N_1552,N_1185,In_2638);
xnor U1553 (N_1553,N_661,In_62);
nor U1554 (N_1554,In_4548,N_955);
nand U1555 (N_1555,N_928,In_3441);
and U1556 (N_1556,In_190,In_535);
nand U1557 (N_1557,In_2402,In_2860);
or U1558 (N_1558,In_2994,N_1393);
and U1559 (N_1559,In_1760,In_2547);
nor U1560 (N_1560,N_1055,N_501);
nand U1561 (N_1561,N_112,In_357);
and U1562 (N_1562,In_912,N_1023);
or U1563 (N_1563,In_4132,In_263);
nand U1564 (N_1564,In_1835,In_4771);
and U1565 (N_1565,In_3453,In_517);
nand U1566 (N_1566,In_2034,In_4275);
nor U1567 (N_1567,In_3652,In_450);
and U1568 (N_1568,In_304,N_921);
xnor U1569 (N_1569,In_1463,In_3039);
nand U1570 (N_1570,N_725,In_2684);
xnor U1571 (N_1571,N_309,In_4965);
nor U1572 (N_1572,N_153,In_162);
nand U1573 (N_1573,In_4724,In_3814);
and U1574 (N_1574,N_731,In_1704);
or U1575 (N_1575,In_4457,In_3165);
nand U1576 (N_1576,In_915,In_4908);
nand U1577 (N_1577,In_4610,In_2644);
or U1578 (N_1578,N_1399,In_232);
nand U1579 (N_1579,In_2963,N_1293);
and U1580 (N_1580,N_1240,In_4263);
or U1581 (N_1581,N_114,In_16);
or U1582 (N_1582,N_1297,In_2799);
or U1583 (N_1583,N_445,In_92);
nor U1584 (N_1584,In_921,In_294);
and U1585 (N_1585,In_3608,In_9);
xor U1586 (N_1586,In_804,In_3012);
xor U1587 (N_1587,In_491,In_4246);
nand U1588 (N_1588,N_893,In_1953);
nor U1589 (N_1589,In_3559,In_2795);
and U1590 (N_1590,In_661,N_903);
nand U1591 (N_1591,In_3818,N_1410);
nor U1592 (N_1592,N_831,In_578);
nand U1593 (N_1593,N_185,In_4463);
nor U1594 (N_1594,In_1762,In_739);
nor U1595 (N_1595,N_958,In_210);
nand U1596 (N_1596,In_230,N_1357);
nand U1597 (N_1597,N_837,N_200);
or U1598 (N_1598,In_3980,In_4923);
or U1599 (N_1599,In_4355,In_2608);
xor U1600 (N_1600,N_8,N_799);
or U1601 (N_1601,In_4409,In_4763);
nand U1602 (N_1602,N_321,N_1071);
nand U1603 (N_1603,N_1304,N_713);
xor U1604 (N_1604,In_1415,In_944);
and U1605 (N_1605,In_1509,In_1133);
xnor U1606 (N_1606,N_69,In_3212);
or U1607 (N_1607,In_234,In_1592);
nor U1608 (N_1608,N_745,In_1077);
or U1609 (N_1609,In_3641,N_651);
nand U1610 (N_1610,In_1268,In_1628);
nor U1611 (N_1611,In_3535,In_1611);
and U1612 (N_1612,In_903,N_1166);
nand U1613 (N_1613,N_1010,In_1506);
xor U1614 (N_1614,In_1904,In_275);
xnor U1615 (N_1615,In_1740,N_1252);
xor U1616 (N_1616,N_702,In_3374);
and U1617 (N_1617,N_1196,In_2793);
nor U1618 (N_1618,In_4696,In_3463);
or U1619 (N_1619,In_4217,In_3198);
xnor U1620 (N_1620,In_81,N_1226);
and U1621 (N_1621,N_847,In_1739);
xor U1622 (N_1622,In_1068,In_1258);
or U1623 (N_1623,In_2589,In_1938);
nor U1624 (N_1624,In_3973,In_4915);
and U1625 (N_1625,In_2246,In_593);
or U1626 (N_1626,In_1245,N_757);
and U1627 (N_1627,In_605,In_163);
nand U1628 (N_1628,In_750,N_976);
nand U1629 (N_1629,In_608,In_832);
nand U1630 (N_1630,N_1375,In_3061);
nor U1631 (N_1631,In_4403,In_4354);
or U1632 (N_1632,In_626,In_2782);
nor U1633 (N_1633,N_1412,In_764);
nor U1634 (N_1634,N_370,In_4659);
or U1635 (N_1635,N_1494,In_4950);
xnor U1636 (N_1636,In_871,In_4229);
xor U1637 (N_1637,In_2959,In_1220);
and U1638 (N_1638,In_1758,In_2108);
nand U1639 (N_1639,N_302,In_4600);
nor U1640 (N_1640,N_423,In_1511);
nor U1641 (N_1641,In_1847,In_1936);
xor U1642 (N_1642,In_416,In_2700);
nand U1643 (N_1643,N_1334,In_4062);
nor U1644 (N_1644,N_164,N_1012);
or U1645 (N_1645,N_1054,In_459);
xnor U1646 (N_1646,In_3384,In_4022);
nand U1647 (N_1647,In_170,N_326);
and U1648 (N_1648,In_4387,In_3983);
nor U1649 (N_1649,In_1125,In_119);
nand U1650 (N_1650,In_2335,In_1930);
nand U1651 (N_1651,N_21,In_3211);
nand U1652 (N_1652,In_4356,In_1097);
and U1653 (N_1653,In_2113,In_4774);
xor U1654 (N_1654,In_2344,In_4622);
nor U1655 (N_1655,N_317,In_3265);
or U1656 (N_1656,N_455,In_2103);
and U1657 (N_1657,N_1458,In_815);
and U1658 (N_1658,In_1397,N_557);
or U1659 (N_1659,In_2780,In_334);
nand U1660 (N_1660,In_2033,N_25);
and U1661 (N_1661,In_433,In_2430);
or U1662 (N_1662,In_4790,In_3344);
xnor U1663 (N_1663,In_272,In_397);
nor U1664 (N_1664,In_411,In_1831);
nand U1665 (N_1665,In_3166,N_484);
xnor U1666 (N_1666,N_729,In_1976);
xnor U1667 (N_1667,N_1121,In_4607);
nand U1668 (N_1668,N_1452,In_3289);
xnor U1669 (N_1669,In_3728,In_4293);
and U1670 (N_1670,In_1527,In_681);
and U1671 (N_1671,N_1244,N_1360);
xor U1672 (N_1672,In_2195,In_4244);
or U1673 (N_1673,In_2697,N_1480);
and U1674 (N_1674,In_2995,In_4806);
nor U1675 (N_1675,In_976,In_4366);
xnor U1676 (N_1676,N_435,In_3697);
and U1677 (N_1677,In_3296,In_1697);
or U1678 (N_1678,In_402,In_1156);
nor U1679 (N_1679,In_3292,In_2239);
xor U1680 (N_1680,In_1265,In_2911);
or U1681 (N_1681,In_4128,N_1427);
and U1682 (N_1682,In_2670,N_500);
nor U1683 (N_1683,N_631,In_2605);
xnor U1684 (N_1684,N_1271,N_695);
nand U1685 (N_1685,In_1364,In_555);
xor U1686 (N_1686,In_723,In_2970);
nor U1687 (N_1687,N_1024,In_4410);
and U1688 (N_1688,In_3919,In_3612);
and U1689 (N_1689,N_1489,In_3696);
nand U1690 (N_1690,In_3169,In_4276);
nand U1691 (N_1691,In_2486,In_1899);
xor U1692 (N_1692,In_3094,N_495);
nor U1693 (N_1693,In_2126,N_1477);
nand U1694 (N_1694,N_155,N_776);
nand U1695 (N_1695,N_1125,In_1729);
and U1696 (N_1696,In_2133,In_446);
nand U1697 (N_1697,In_1280,In_12);
nor U1698 (N_1698,In_1204,In_4630);
or U1699 (N_1699,In_1013,In_1456);
xor U1700 (N_1700,N_451,In_3788);
nor U1701 (N_1701,In_1678,In_3185);
and U1702 (N_1702,In_4830,N_672);
xnor U1703 (N_1703,N_526,N_1100);
nor U1704 (N_1704,N_267,In_4780);
xnor U1705 (N_1705,In_3107,N_1438);
xnor U1706 (N_1706,In_2494,N_60);
or U1707 (N_1707,N_579,In_3878);
nand U1708 (N_1708,In_3030,In_1171);
nand U1709 (N_1709,N_1205,In_4969);
xor U1710 (N_1710,In_2448,N_938);
xnor U1711 (N_1711,N_77,In_126);
nand U1712 (N_1712,In_2732,N_1288);
or U1713 (N_1713,In_2617,In_2449);
and U1714 (N_1714,N_480,In_1186);
xor U1715 (N_1715,In_38,N_1144);
or U1716 (N_1716,In_4631,N_616);
and U1717 (N_1717,N_468,N_1248);
and U1718 (N_1718,N_1450,In_4731);
xnor U1719 (N_1719,N_363,In_1035);
and U1720 (N_1720,In_4301,In_551);
and U1721 (N_1721,In_2138,In_3720);
nand U1722 (N_1722,In_215,In_1929);
and U1723 (N_1723,In_4484,N_1170);
nor U1724 (N_1724,In_4284,In_1345);
xnor U1725 (N_1725,In_4844,N_586);
nor U1726 (N_1726,In_4840,In_4897);
nor U1727 (N_1727,N_1197,N_520);
and U1728 (N_1728,In_3604,In_590);
xnor U1729 (N_1729,In_26,In_4497);
or U1730 (N_1730,In_2529,In_1036);
nand U1731 (N_1731,N_1255,In_348);
and U1732 (N_1732,In_4432,In_4421);
nor U1733 (N_1733,In_3103,In_3254);
nand U1734 (N_1734,In_2712,In_3584);
nor U1735 (N_1735,In_3346,In_2675);
xnor U1736 (N_1736,In_2025,In_4269);
nor U1737 (N_1737,N_598,In_429);
and U1738 (N_1738,In_4776,N_806);
nor U1739 (N_1739,In_10,In_3235);
xor U1740 (N_1740,N_1411,In_3448);
nand U1741 (N_1741,In_635,N_1469);
nor U1742 (N_1742,In_3303,N_801);
xor U1743 (N_1743,In_879,In_2583);
nor U1744 (N_1744,In_2800,In_1115);
xor U1745 (N_1745,In_1871,In_4124);
nor U1746 (N_1746,In_552,In_2252);
nor U1747 (N_1747,N_1142,In_3546);
or U1748 (N_1748,In_1188,In_1815);
or U1749 (N_1749,In_2924,N_1415);
nand U1750 (N_1750,N_1153,In_2180);
xnor U1751 (N_1751,N_5,In_2903);
nor U1752 (N_1752,N_1234,N_1609);
nor U1753 (N_1753,In_2042,In_899);
or U1754 (N_1754,N_1484,N_1521);
xor U1755 (N_1755,In_4474,In_48);
and U1756 (N_1756,In_4277,N_498);
nand U1757 (N_1757,In_3366,In_4983);
xnor U1758 (N_1758,In_2010,In_4756);
or U1759 (N_1759,In_649,In_829);
or U1760 (N_1760,In_855,In_2404);
or U1761 (N_1761,In_3883,N_1718);
nor U1762 (N_1762,N_963,In_1523);
xor U1763 (N_1763,N_117,N_1167);
nor U1764 (N_1764,In_1445,In_1401);
xnor U1765 (N_1765,In_4028,N_1269);
or U1766 (N_1766,In_2775,N_465);
nor U1767 (N_1767,In_1274,In_1820);
nor U1768 (N_1768,In_4765,N_817);
or U1769 (N_1769,In_1229,N_669);
and U1770 (N_1770,N_1173,In_1633);
nor U1771 (N_1771,In_3781,N_1294);
or U1772 (N_1772,In_3111,In_1261);
nand U1773 (N_1773,In_2226,N_1554);
or U1774 (N_1774,N_739,N_851);
xnor U1775 (N_1775,N_740,N_856);
or U1776 (N_1776,N_473,In_749);
and U1777 (N_1777,In_2854,N_111);
or U1778 (N_1778,In_33,In_2654);
xor U1779 (N_1779,In_4894,N_1692);
xnor U1780 (N_1780,N_1497,In_1602);
or U1781 (N_1781,N_906,In_3729);
and U1782 (N_1782,N_1625,N_52);
nand U1783 (N_1783,In_4296,In_3425);
or U1784 (N_1784,In_3823,In_4253);
nand U1785 (N_1785,In_3628,In_3262);
xor U1786 (N_1786,In_1285,In_3887);
nor U1787 (N_1787,In_3515,N_120);
and U1788 (N_1788,In_4137,N_1428);
or U1789 (N_1789,N_1472,In_4677);
and U1790 (N_1790,N_1319,In_3064);
and U1791 (N_1791,In_1564,In_2185);
nor U1792 (N_1792,In_2926,In_3401);
xnor U1793 (N_1793,N_1003,In_2830);
nor U1794 (N_1794,In_715,In_4187);
xor U1795 (N_1795,In_684,N_608);
nor U1796 (N_1796,N_434,N_516);
or U1797 (N_1797,N_1731,In_1147);
nor U1798 (N_1798,In_1726,In_3310);
nand U1799 (N_1799,In_2558,N_984);
nand U1800 (N_1800,N_1606,In_4477);
or U1801 (N_1801,In_3763,In_2842);
xor U1802 (N_1802,In_231,In_3932);
xnor U1803 (N_1803,In_3475,In_3681);
and U1804 (N_1804,N_1303,In_4002);
nand U1805 (N_1805,In_4007,In_4015);
and U1806 (N_1806,In_2579,In_2997);
or U1807 (N_1807,N_1700,In_1334);
xnor U1808 (N_1808,N_785,In_1022);
xnor U1809 (N_1809,N_1470,In_1016);
nand U1810 (N_1810,In_3851,N_1401);
nor U1811 (N_1811,In_2046,In_2236);
or U1812 (N_1812,N_1556,N_760);
xnor U1813 (N_1813,In_4943,N_735);
nor U1814 (N_1814,N_818,N_581);
xor U1815 (N_1815,In_2258,N_1416);
nand U1816 (N_1816,In_895,N_839);
nor U1817 (N_1817,In_1339,N_288);
or U1818 (N_1818,N_602,In_1026);
xor U1819 (N_1819,In_1541,In_886);
and U1820 (N_1820,In_1684,In_2244);
xnor U1821 (N_1821,In_3233,In_233);
nor U1822 (N_1822,In_3780,In_3901);
and U1823 (N_1823,In_4885,In_128);
and U1824 (N_1824,N_1330,In_228);
nor U1825 (N_1825,In_4168,In_2984);
or U1826 (N_1826,In_4488,In_1721);
xor U1827 (N_1827,In_4626,In_3368);
nor U1828 (N_1828,N_1044,N_1307);
nand U1829 (N_1829,In_1040,In_3206);
nor U1830 (N_1830,N_1015,In_2145);
or U1831 (N_1831,In_3095,In_2022);
and U1832 (N_1832,N_1372,In_3227);
or U1833 (N_1833,N_1576,N_1343);
xnor U1834 (N_1834,In_4713,In_106);
and U1835 (N_1835,In_1914,In_809);
xnor U1836 (N_1836,In_3895,N_486);
and U1837 (N_1837,In_4285,In_164);
and U1838 (N_1838,In_168,In_2660);
or U1839 (N_1839,In_238,In_2946);
nand U1840 (N_1840,In_3079,N_1583);
nor U1841 (N_1841,N_756,In_4644);
or U1842 (N_1842,In_1890,In_1750);
or U1843 (N_1843,N_800,N_1311);
nand U1844 (N_1844,N_1426,N_228);
xnor U1845 (N_1845,In_1696,In_1141);
and U1846 (N_1846,In_641,In_1933);
nor U1847 (N_1847,In_2694,N_1095);
nor U1848 (N_1848,In_736,N_547);
or U1849 (N_1849,In_3990,N_621);
nand U1850 (N_1850,N_1642,In_1555);
nand U1851 (N_1851,In_1869,In_962);
nor U1852 (N_1852,N_532,In_698);
xor U1853 (N_1853,N_1061,In_3571);
nor U1854 (N_1854,In_3424,N_1256);
nor U1855 (N_1855,In_11,N_780);
and U1856 (N_1856,N_1475,N_1260);
or U1857 (N_1857,N_649,N_1388);
xor U1858 (N_1858,In_1495,In_52);
and U1859 (N_1859,In_4326,In_3935);
nand U1860 (N_1860,In_1325,N_1072);
and U1861 (N_1861,N_907,N_948);
xnor U1862 (N_1862,In_2920,N_803);
or U1863 (N_1863,In_1923,In_2480);
xnor U1864 (N_1864,In_3563,N_1174);
xor U1865 (N_1865,In_3101,In_2102);
nand U1866 (N_1866,In_4352,N_1591);
and U1867 (N_1867,N_3,N_496);
and U1868 (N_1868,In_3850,In_2143);
or U1869 (N_1869,In_2177,N_946);
xor U1870 (N_1870,In_1826,N_1328);
or U1871 (N_1871,In_61,N_752);
xnor U1872 (N_1872,In_3392,In_901);
nor U1873 (N_1873,N_600,In_1573);
nor U1874 (N_1874,In_2238,In_875);
and U1875 (N_1875,In_3397,In_2152);
and U1876 (N_1876,N_777,N_504);
nor U1877 (N_1877,In_312,In_839);
xnor U1878 (N_1878,In_1997,N_1339);
and U1879 (N_1879,In_544,In_2251);
xnor U1880 (N_1880,N_1296,N_1129);
and U1881 (N_1881,In_2419,In_1047);
and U1882 (N_1882,N_860,In_2417);
nand U1883 (N_1883,N_1523,In_2049);
and U1884 (N_1884,N_1659,In_4671);
nand U1885 (N_1885,In_4812,N_682);
nand U1886 (N_1886,N_490,N_1435);
and U1887 (N_1887,In_705,In_1722);
or U1888 (N_1888,N_1152,In_3906);
nand U1889 (N_1889,In_1340,In_4541);
and U1890 (N_1890,In_3477,In_280);
xor U1891 (N_1891,In_3695,In_3320);
or U1892 (N_1892,N_49,N_248);
or U1893 (N_1893,In_1476,In_4927);
or U1894 (N_1894,N_1608,In_44);
nand U1895 (N_1895,In_1843,N_437);
nand U1896 (N_1896,In_2401,In_1881);
and U1897 (N_1897,In_290,In_3274);
nor U1898 (N_1898,N_877,N_1308);
xnor U1899 (N_1899,In_2972,In_221);
nand U1900 (N_1900,N_1018,N_1059);
or U1901 (N_1901,In_2856,In_792);
or U1902 (N_1902,In_2217,In_1023);
xnor U1903 (N_1903,In_982,In_2227);
and U1904 (N_1904,In_3486,N_811);
and U1905 (N_1905,N_1160,In_4133);
nor U1906 (N_1906,In_1413,N_54);
nor U1907 (N_1907,N_641,N_855);
or U1908 (N_1908,In_425,In_4606);
and U1909 (N_1909,N_1614,In_2717);
xnor U1910 (N_1910,N_181,In_3440);
and U1911 (N_1911,In_1267,N_335);
nor U1912 (N_1912,In_1840,N_728);
nor U1913 (N_1913,In_2363,In_1514);
nor U1914 (N_1914,N_446,In_1579);
nand U1915 (N_1915,In_3132,In_3317);
and U1916 (N_1916,N_819,N_1109);
xnor U1917 (N_1917,In_933,N_1398);
and U1918 (N_1918,N_1716,In_2016);
nand U1919 (N_1919,In_1893,In_21);
nand U1920 (N_1920,In_2481,In_4666);
nand U1921 (N_1921,In_3070,In_3590);
nand U1922 (N_1922,In_4928,In_4344);
nand U1923 (N_1923,In_2104,N_1092);
or U1924 (N_1924,In_4772,In_2511);
xnor U1925 (N_1925,In_4940,N_1143);
or U1926 (N_1926,In_4552,In_2618);
nand U1927 (N_1927,N_1267,In_543);
or U1928 (N_1928,N_827,N_1091);
nor U1929 (N_1929,In_2065,In_2298);
nand U1930 (N_1930,In_3489,N_1199);
xor U1931 (N_1931,In_3357,In_2790);
xnor U1932 (N_1932,N_1592,In_1566);
nand U1933 (N_1933,N_1282,In_1412);
and U1934 (N_1934,In_3598,In_4648);
or U1935 (N_1935,N_1156,In_3406);
nand U1936 (N_1936,In_2765,N_1704);
nor U1937 (N_1937,N_1000,In_954);
and U1938 (N_1938,In_1902,N_1191);
and U1939 (N_1939,N_673,In_1738);
and U1940 (N_1940,N_1115,In_4956);
xnor U1941 (N_1941,In_952,In_4376);
and U1942 (N_1942,In_2531,In_4536);
and U1943 (N_1943,In_452,N_1370);
and U1944 (N_1944,In_3961,N_1571);
or U1945 (N_1945,In_2075,In_2436);
nor U1946 (N_1946,In_4219,N_250);
xnor U1947 (N_1947,In_3860,In_519);
nor U1948 (N_1948,In_2941,N_905);
or U1949 (N_1949,In_3819,In_591);
nand U1950 (N_1950,In_375,In_4458);
xnor U1951 (N_1951,In_267,In_4892);
and U1952 (N_1952,In_653,N_759);
or U1953 (N_1953,In_4087,In_435);
or U1954 (N_1954,In_646,In_3858);
or U1955 (N_1955,In_1772,N_91);
and U1956 (N_1956,N_804,N_1395);
and U1957 (N_1957,In_974,N_1735);
or U1958 (N_1958,N_1647,N_1445);
nor U1959 (N_1959,N_596,N_1285);
nand U1960 (N_1960,In_4042,N_627);
nor U1961 (N_1961,In_3827,N_102);
or U1962 (N_1962,N_904,In_2506);
and U1963 (N_1963,In_4874,In_972);
xnor U1964 (N_1964,In_85,N_293);
xor U1965 (N_1965,In_2249,N_1696);
or U1966 (N_1966,In_969,N_137);
nor U1967 (N_1967,In_1744,In_3664);
xor U1968 (N_1968,In_3898,In_2340);
xor U1969 (N_1969,In_4311,In_2383);
or U1970 (N_1970,In_1320,N_1275);
xor U1971 (N_1971,In_3053,In_3090);
nand U1972 (N_1972,N_593,N_272);
xnor U1973 (N_1973,N_1229,In_2874);
nand U1974 (N_1974,In_1318,In_4989);
nor U1975 (N_1975,N_595,In_2169);
and U1976 (N_1976,In_3715,In_3046);
and U1977 (N_1977,N_1178,N_994);
nor U1978 (N_1978,In_3279,In_2386);
and U1979 (N_1979,In_2810,In_1324);
nand U1980 (N_1980,N_1361,N_257);
nand U1981 (N_1981,N_794,N_1037);
or U1982 (N_1982,In_3476,In_533);
nand U1983 (N_1983,In_1646,N_812);
and U1984 (N_1984,N_1542,In_2035);
and U1985 (N_1985,In_4854,In_806);
or U1986 (N_1986,In_3541,In_1945);
nand U1987 (N_1987,N_1098,N_1257);
or U1988 (N_1988,In_473,In_2304);
nor U1989 (N_1989,In_1948,In_2149);
or U1990 (N_1990,In_2166,N_1047);
nand U1991 (N_1991,In_1179,N_1089);
or U1992 (N_1992,N_1368,In_2875);
and U1993 (N_1993,In_4122,In_4129);
or U1994 (N_1994,In_779,In_609);
xnor U1995 (N_1995,In_4139,In_3403);
or U1996 (N_1996,N_413,N_972);
nor U1997 (N_1997,In_4523,In_2804);
and U1998 (N_1998,In_858,In_187);
or U1999 (N_1999,In_3312,N_924);
nor U2000 (N_2000,In_3952,N_894);
nor U2001 (N_2001,In_4515,In_3181);
and U2002 (N_2002,In_636,N_294);
nand U2003 (N_2003,N_347,N_1200);
xor U2004 (N_2004,In_1519,In_2746);
nor U2005 (N_2005,In_444,In_4863);
nand U2006 (N_2006,N_930,In_84);
nor U2007 (N_2007,N_1981,In_4708);
or U2008 (N_2008,N_1768,N_371);
nor U2009 (N_2009,In_1952,In_3538);
nor U2010 (N_2010,In_1841,N_1871);
nand U2011 (N_2011,N_1683,N_1353);
xnor U2012 (N_2012,In_1703,N_214);
xor U2013 (N_2013,N_1079,In_4188);
nand U2014 (N_2014,N_1502,In_4338);
or U2015 (N_2015,In_1774,N_1921);
nor U2016 (N_2016,N_1348,N_1045);
or U2017 (N_2017,In_588,In_676);
or U2018 (N_2018,In_1619,N_551);
xnor U2019 (N_2019,In_3382,In_3305);
or U2020 (N_2020,N_1373,In_2666);
or U2021 (N_2021,In_4980,N_1495);
nand U2022 (N_2022,N_1300,N_1829);
or U2023 (N_2023,N_1823,In_3468);
nand U2024 (N_2024,In_1008,N_974);
nor U2025 (N_2025,N_997,In_2170);
xor U2026 (N_2026,In_1596,In_4951);
nand U2027 (N_2027,N_849,N_327);
or U2028 (N_2028,N_1014,In_1120);
xor U2029 (N_2029,N_895,In_2525);
or U2030 (N_2030,In_2207,In_3555);
xnor U2031 (N_2031,In_911,N_1882);
and U2032 (N_2032,N_106,N_1586);
nor U2033 (N_2033,N_1347,In_2818);
xor U2034 (N_2034,In_1645,In_4574);
and U2035 (N_2035,In_353,In_4491);
xor U2036 (N_2036,In_814,N_658);
and U2037 (N_2037,In_4021,N_1362);
nor U2038 (N_2038,In_1393,In_4400);
and U2039 (N_2039,N_1861,In_3372);
or U2040 (N_2040,N_628,In_4661);
nor U2041 (N_2041,In_1581,In_3354);
xnor U2042 (N_2042,In_2067,N_939);
xor U2043 (N_2043,N_105,In_4308);
xor U2044 (N_2044,In_537,In_2078);
nand U2045 (N_2045,N_1546,In_463);
nand U2046 (N_2046,N_1064,N_843);
or U2047 (N_2047,In_58,In_1920);
xnor U2048 (N_2048,In_2603,N_171);
xnor U2049 (N_2049,In_2097,N_298);
or U2050 (N_2050,In_4370,In_586);
nor U2051 (N_2051,In_4238,In_1126);
and U2052 (N_2052,N_1102,In_3479);
and U2053 (N_2053,N_1918,N_1537);
nor U2054 (N_2054,N_779,N_1570);
and U2055 (N_2055,N_1063,N_1407);
nand U2056 (N_2056,N_1813,In_1287);
nor U2057 (N_2057,N_134,In_2259);
and U2058 (N_2058,N_1913,N_1558);
xnor U2059 (N_2059,In_1695,In_4899);
nand U2060 (N_2060,In_351,In_1001);
xnor U2061 (N_2061,N_762,N_1374);
xor U2062 (N_2062,In_955,In_3490);
nand U2063 (N_2063,N_1409,In_2748);
and U2064 (N_2064,In_1072,N_1491);
nand U2065 (N_2065,In_3870,N_1369);
xnor U2066 (N_2066,In_3323,N_1690);
or U2067 (N_2067,In_3180,In_1830);
or U2068 (N_2068,In_453,N_549);
xnor U2069 (N_2069,In_3033,In_1686);
nor U2070 (N_2070,In_2450,N_1441);
nand U2071 (N_2071,In_2200,N_1858);
xnor U2072 (N_2072,In_4688,In_1107);
nand U2073 (N_2073,In_245,N_1127);
or U2074 (N_2074,N_461,In_3387);
nand U2075 (N_2075,In_4199,In_3332);
nand U2076 (N_2076,In_4305,In_2906);
or U2077 (N_2077,In_3051,In_4634);
nor U2078 (N_2078,In_1310,In_3351);
xor U2079 (N_2079,N_90,In_2303);
and U2080 (N_2080,N_1301,In_4303);
and U2081 (N_2081,In_2564,In_4591);
or U2082 (N_2082,N_1812,N_1408);
and U2083 (N_2083,In_2213,In_2324);
or U2084 (N_2084,N_1876,In_2329);
xnor U2085 (N_2085,In_3892,In_2599);
or U2086 (N_2086,In_1998,N_87);
xor U2087 (N_2087,In_3464,N_1057);
or U2088 (N_2088,N_1896,N_1354);
xnor U2089 (N_2089,N_1126,In_420);
xor U2090 (N_2090,In_1292,N_826);
and U2091 (N_2091,In_1418,In_1106);
xor U2092 (N_2092,N_1822,In_2649);
nand U2093 (N_2093,In_1359,In_2811);
xor U2094 (N_2094,In_2206,In_264);
nand U2095 (N_2095,In_2083,In_1962);
and U2096 (N_2096,N_1454,In_4732);
nand U2097 (N_2097,In_4572,In_2567);
nand U2098 (N_2098,N_1744,In_2000);
nand U2099 (N_2099,In_3690,N_63);
and U2100 (N_2100,In_3099,In_1531);
and U2101 (N_2101,In_493,In_2650);
and U2102 (N_2102,N_1228,In_4209);
nor U2103 (N_2103,N_1215,In_4069);
nand U2104 (N_2104,In_3328,In_1836);
nor U2105 (N_2105,In_4662,In_4479);
xnor U2106 (N_2106,N_1305,N_1747);
nor U2107 (N_2107,N_1509,In_2028);
xnor U2108 (N_2108,N_1960,In_4088);
and U2109 (N_2109,N_724,In_2325);
nand U2110 (N_2110,N_1957,In_3955);
nor U2111 (N_2111,N_438,In_4804);
or U2112 (N_2112,N_552,In_3268);
and U2113 (N_2113,In_1378,In_2726);
nor U2114 (N_2114,In_1754,In_893);
nor U2115 (N_2115,In_2951,In_3209);
or U2116 (N_2116,In_4621,In_4440);
and U2117 (N_2117,N_1119,N_1803);
and U2118 (N_2118,N_1972,In_15);
nor U2119 (N_2119,N_929,In_3768);
nand U2120 (N_2120,N_1897,N_684);
nand U2121 (N_2121,N_1880,N_488);
and U2122 (N_2122,In_332,In_1669);
or U2123 (N_2123,N_1759,N_575);
nor U2124 (N_2124,In_603,N_467);
or U2125 (N_2125,N_949,In_4169);
xnor U2126 (N_2126,In_2822,N_514);
and U2127 (N_2127,In_2766,N_1147);
and U2128 (N_2128,In_630,In_1389);
nor U2129 (N_2129,In_1116,In_2125);
nand U2130 (N_2130,N_1140,In_3045);
nand U2131 (N_2131,In_2204,In_3674);
nor U2132 (N_2132,In_2643,N_1270);
nor U2133 (N_2133,N_1463,N_1253);
or U2134 (N_2134,In_3217,In_1876);
nand U2135 (N_2135,In_597,N_229);
or U2136 (N_2136,In_690,In_1297);
or U2137 (N_2137,In_2513,In_4450);
nor U2138 (N_2138,In_4161,In_3022);
or U2139 (N_2139,N_916,N_662);
xnor U2140 (N_2140,N_1448,In_2454);
and U2141 (N_2141,In_904,In_4654);
xnor U2142 (N_2142,N_1084,N_902);
nand U2143 (N_2143,In_2524,In_3852);
xor U2144 (N_2144,In_2554,In_1303);
or U2145 (N_2145,N_386,N_1111);
nand U2146 (N_2146,In_557,In_1931);
or U2147 (N_2147,In_4667,In_2210);
and U2148 (N_2148,In_2534,N_233);
or U2149 (N_2149,In_2886,In_3236);
xor U2150 (N_2150,In_3948,In_4475);
or U2151 (N_2151,N_1549,N_925);
and U2152 (N_2152,In_2607,N_1728);
nor U2153 (N_2153,In_3156,In_2205);
nor U2154 (N_2154,N_854,In_2315);
xor U2155 (N_2155,N_1828,N_1421);
and U2156 (N_2156,N_197,N_1852);
and U2157 (N_2157,N_1588,In_3523);
and U2158 (N_2158,N_1496,In_1385);
and U2159 (N_2159,In_1051,In_1917);
or U2160 (N_2160,N_1402,In_2483);
nor U2161 (N_2161,N_1384,In_3836);
and U2162 (N_2162,N_1924,In_1467);
or U2163 (N_2163,N_869,In_2508);
nor U2164 (N_2164,N_1371,N_1671);
xnor U2165 (N_2165,N_1932,In_964);
or U2166 (N_2166,N_1557,In_1351);
nor U2167 (N_2167,In_2434,N_1589);
nand U2168 (N_2168,In_3020,In_787);
nor U2169 (N_2169,In_4348,N_396);
nor U2170 (N_2170,In_1431,In_1990);
and U2171 (N_2171,N_1385,In_2532);
or U2172 (N_2172,N_701,N_1418);
nand U2173 (N_2173,In_2611,In_2128);
nor U2174 (N_2174,In_2270,N_1765);
and U2175 (N_2175,N_1975,In_2634);
nor U2176 (N_2176,In_4056,In_1951);
and U2177 (N_2177,In_576,N_358);
nor U2178 (N_2178,N_1915,In_703);
and U2179 (N_2179,In_4465,In_4528);
nor U2180 (N_2180,In_2862,In_4995);
nand U2181 (N_2181,In_3047,In_99);
and U2182 (N_2182,In_756,In_1045);
xor U2183 (N_2183,In_2896,N_1419);
xnor U2184 (N_2184,N_527,In_2356);
or U2185 (N_2185,In_297,In_2179);
nor U2186 (N_2186,N_942,N_1529);
and U2187 (N_2187,In_69,In_2109);
nand U2188 (N_2188,N_1968,In_2813);
nor U2189 (N_2189,In_524,In_1850);
xor U2190 (N_2190,N_383,N_1207);
nand U2191 (N_2191,N_97,N_232);
or U2192 (N_2192,N_1227,N_1598);
nand U2193 (N_2193,In_2269,In_2418);
and U2194 (N_2194,In_17,N_1993);
and U2195 (N_2195,N_1043,In_274);
nand U2196 (N_2196,In_3238,In_4070);
xor U2197 (N_2197,In_2671,N_122);
nand U2198 (N_2198,In_1484,In_4389);
and U2199 (N_2199,In_963,N_1703);
xor U2200 (N_2200,N_314,In_831);
xor U2201 (N_2201,N_80,In_344);
or U2202 (N_2202,In_3995,N_901);
and U2203 (N_2203,In_2542,N_1727);
nor U2204 (N_2204,In_2495,N_1350);
xor U2205 (N_2205,In_3293,N_569);
nor U2206 (N_2206,N_167,In_3426);
xor U2207 (N_2207,N_770,In_1386);
nand U2208 (N_2208,N_1832,In_152);
or U2209 (N_2209,N_1313,In_2545);
and U2210 (N_2210,In_3183,In_2733);
or U2211 (N_2211,N_243,N_876);
and U2212 (N_2212,In_3128,N_22);
and U2213 (N_2213,N_1021,In_1215);
nor U2214 (N_2214,In_4942,N_1794);
nand U2215 (N_2215,In_74,In_340);
nand U2216 (N_2216,In_3544,In_4941);
and U2217 (N_2217,In_4404,N_1710);
and U2218 (N_2218,In_2745,In_2005);
or U2219 (N_2219,In_4728,In_4483);
or U2220 (N_2220,In_1050,In_4623);
or U2221 (N_2221,In_717,In_4089);
nor U2222 (N_2222,N_218,In_2265);
nand U2223 (N_2223,N_1908,In_1608);
nor U2224 (N_2224,In_754,N_1210);
xor U2225 (N_2225,In_1854,In_3162);
nor U2226 (N_2226,N_1287,In_3880);
and U2227 (N_2227,In_4115,In_1373);
xnor U2228 (N_2228,In_1954,In_1653);
nand U2229 (N_2229,N_1320,N_1073);
or U2230 (N_2230,N_714,N_408);
nand U2231 (N_2231,N_463,In_1582);
and U2232 (N_2232,N_1397,N_1691);
xor U2233 (N_2233,N_545,In_56);
nand U2234 (N_2234,N_508,In_2502);
nor U2235 (N_2235,N_618,In_1660);
nand U2236 (N_2236,N_1892,In_3640);
xnor U2237 (N_2237,N_1748,In_870);
and U2238 (N_2238,N_199,N_544);
xor U2239 (N_2239,In_4402,In_991);
nand U2240 (N_2240,N_1490,In_2214);
and U2241 (N_2241,In_575,In_1851);
xor U2242 (N_2242,In_1595,N_1611);
nand U2243 (N_2243,N_950,In_965);
nand U2244 (N_2244,N_403,N_1773);
and U2245 (N_2245,In_2184,In_191);
nand U2246 (N_2246,N_1618,N_1237);
xor U2247 (N_2247,In_470,In_1968);
nand U2248 (N_2248,In_4690,In_3614);
and U2249 (N_2249,In_4846,N_284);
xor U2250 (N_2250,N_2005,In_3790);
or U2251 (N_2251,In_4788,In_4749);
nand U2252 (N_2252,In_4647,N_1958);
nor U2253 (N_2253,N_761,N_1417);
nand U2254 (N_2254,N_2239,N_2124);
or U2255 (N_2255,N_1316,In_2768);
nand U2256 (N_2256,In_1803,In_1502);
nor U2257 (N_2257,In_2017,In_3629);
xnor U2258 (N_2258,N_1663,N_2215);
and U2259 (N_2259,N_1164,In_1482);
xor U2260 (N_2260,In_2767,In_1891);
and U2261 (N_2261,N_2238,N_2129);
nor U2262 (N_2262,N_2052,N_919);
or U2263 (N_2263,In_4753,In_1271);
nor U2264 (N_2264,In_3977,N_1912);
nand U2265 (N_2265,In_1176,N_1631);
nor U2266 (N_2266,N_1645,N_1966);
and U2267 (N_2267,In_2237,In_4252);
or U2268 (N_2268,N_1928,In_2150);
or U2269 (N_2269,N_1840,In_1713);
or U2270 (N_2270,N_1976,In_136);
or U2271 (N_2271,N_573,N_1927);
nor U2272 (N_2272,In_992,In_2334);
xor U2273 (N_2273,In_4808,N_987);
nor U2274 (N_2274,In_133,In_2219);
nor U2275 (N_2275,N_1706,In_241);
nand U2276 (N_2276,In_2574,In_4966);
nand U2277 (N_2277,In_4249,In_3210);
nor U2278 (N_2278,N_1904,In_3936);
and U2279 (N_2279,In_1605,In_2043);
nor U2280 (N_2280,In_4546,In_467);
or U2281 (N_2281,N_1777,In_2092);
xor U2282 (N_2282,N_1548,N_1817);
nand U2283 (N_2283,N_1685,N_993);
nor U2284 (N_2284,N_1872,N_828);
nand U2285 (N_2285,In_607,N_730);
xor U2286 (N_2286,In_3119,In_3213);
xnor U2287 (N_2287,In_4481,N_202);
nand U2288 (N_2288,N_2112,In_1288);
nand U2289 (N_2289,In_2805,N_583);
or U2290 (N_2290,N_1920,In_2615);
nand U2291 (N_2291,In_1367,N_568);
nor U2292 (N_2292,N_1306,N_1040);
xnor U2293 (N_2293,N_959,N_1517);
nand U2294 (N_2294,In_3273,N_372);
nand U2295 (N_2295,In_1629,In_3299);
xor U2296 (N_2296,N_1515,In_1591);
xor U2297 (N_2297,N_988,In_3591);
or U2298 (N_2298,N_1114,N_1610);
nand U2299 (N_2299,In_1778,In_3086);
or U2300 (N_2300,N_1286,In_1870);
nor U2301 (N_2301,In_1715,In_3516);
xor U2302 (N_2302,In_1780,In_877);
or U2303 (N_2303,N_1172,N_966);
nor U2304 (N_2304,N_945,N_1687);
nor U2305 (N_2305,N_2019,In_1038);
nand U2306 (N_2306,In_3702,N_1194);
or U2307 (N_2307,In_3915,In_198);
or U2308 (N_2308,N_1512,In_4358);
xnor U2309 (N_2309,N_2225,N_1437);
or U2310 (N_2310,In_3747,In_419);
or U2311 (N_2311,In_4335,In_4797);
or U2312 (N_2312,In_1377,In_1246);
xnor U2313 (N_2313,In_165,N_1881);
nand U2314 (N_2314,N_1188,In_370);
or U2315 (N_2315,N_1569,In_3016);
xor U2316 (N_2316,In_853,In_1691);
nor U2317 (N_2317,In_816,N_1243);
nand U2318 (N_2318,N_2139,N_1724);
or U2319 (N_2319,In_4953,N_1218);
and U2320 (N_2320,N_2121,In_589);
or U2321 (N_2321,In_4425,N_1314);
or U2322 (N_2322,N_885,N_1077);
nor U2323 (N_2323,In_4711,N_1670);
nor U2324 (N_2324,In_2278,In_23);
xnor U2325 (N_2325,In_18,N_998);
nand U2326 (N_2326,In_2827,N_1824);
nand U2327 (N_2327,N_2212,In_2563);
nand U2328 (N_2328,N_1041,N_273);
and U2329 (N_2329,In_3327,In_2498);
nor U2330 (N_2330,In_3972,N_1870);
nor U2331 (N_2331,N_10,N_1810);
nor U2332 (N_2332,In_1499,In_4272);
nor U2333 (N_2333,In_3766,N_1050);
or U2334 (N_2334,N_751,N_133);
nor U2335 (N_2335,In_2073,In_2553);
nor U2336 (N_2336,In_4320,N_2194);
and U2337 (N_2337,N_850,In_269);
xor U2338 (N_2338,N_1902,In_4691);
nor U2339 (N_2339,N_638,In_3419);
nand U2340 (N_2340,In_4399,In_3067);
nor U2341 (N_2341,In_721,N_1898);
xnor U2342 (N_2342,In_289,In_2240);
nand U2343 (N_2343,N_1520,N_2200);
or U2344 (N_2344,N_1901,N_2015);
nand U2345 (N_2345,In_4307,N_1431);
nand U2346 (N_2346,In_778,In_4047);
and U2347 (N_2347,In_339,In_1361);
or U2348 (N_2348,In_2572,N_1486);
and U2349 (N_2349,N_1158,N_722);
and U2350 (N_2350,N_2186,In_4898);
nor U2351 (N_2351,N_1453,N_910);
xnor U2352 (N_2352,In_3139,N_1617);
nor U2353 (N_2353,N_1650,N_873);
nand U2354 (N_2354,In_2983,In_4553);
and U2355 (N_2355,In_2284,In_3271);
and U2356 (N_2356,In_4154,N_1578);
or U2357 (N_2357,N_1514,In_1180);
nand U2358 (N_2358,In_4294,N_2245);
xnor U2359 (N_2359,N_1154,In_2659);
nand U2360 (N_2360,N_1878,N_2044);
and U2361 (N_2361,In_4520,In_469);
nand U2362 (N_2362,In_1193,In_3383);
or U2363 (N_2363,In_2068,In_1231);
nor U2364 (N_2364,N_100,N_703);
nor U2365 (N_2365,N_1505,N_1131);
or U2366 (N_2366,N_1499,In_849);
xnor U2367 (N_2367,In_1031,N_1786);
and U2368 (N_2368,N_340,In_2832);
nor U2369 (N_2369,N_975,In_4469);
or U2370 (N_2370,In_2981,In_4099);
or U2371 (N_2371,In_3683,In_3108);
nand U2372 (N_2372,In_4707,N_1684);
nor U2373 (N_2373,In_3072,In_2274);
or U2374 (N_2374,N_1498,In_1481);
or U2375 (N_2375,N_2195,N_1265);
xnor U2376 (N_2376,In_4449,In_2851);
nor U2377 (N_2377,In_2613,N_1356);
and U2378 (N_2378,N_1637,N_1381);
nand U2379 (N_2379,In_1092,In_1650);
or U2380 (N_2380,N_1189,In_2023);
nor U2381 (N_2381,N_2192,In_1668);
or U2382 (N_2382,In_733,In_2658);
xor U2383 (N_2383,In_3098,N_2178);
or U2384 (N_2384,N_629,N_1900);
nor U2385 (N_2385,N_565,N_95);
or U2386 (N_2386,In_1478,N_626);
nand U2387 (N_2387,In_4153,N_1930);
nand U2388 (N_2388,In_2098,N_1987);
nor U2389 (N_2389,N_744,In_687);
and U2390 (N_2390,In_4784,In_3163);
nor U2391 (N_2391,In_3793,In_3126);
xnor U2392 (N_2392,In_3705,N_1141);
or U2393 (N_2393,N_1527,N_391);
or U2394 (N_2394,In_2859,In_4014);
and U2395 (N_2395,In_3632,N_477);
nor U2396 (N_2396,N_1106,N_1626);
nor U2397 (N_2397,In_199,In_3844);
xnor U2398 (N_2398,In_1199,In_227);
nor U2399 (N_2399,In_4838,In_4461);
nor U2400 (N_2400,In_2585,In_2333);
and U2401 (N_2401,N_2202,N_503);
or U2402 (N_2402,N_493,N_1946);
xnor U2403 (N_2403,In_1211,N_1090);
nand U2404 (N_2404,In_1042,N_1661);
nor U2405 (N_2405,In_356,In_4503);
nand U2406 (N_2406,N_797,In_72);
xnor U2407 (N_2407,In_1071,In_3451);
nor U2408 (N_2408,N_2207,In_2116);
xnor U2409 (N_2409,In_3600,N_783);
nand U2410 (N_2410,N_1162,N_1639);
or U2411 (N_2411,N_283,N_466);
nor U2412 (N_2412,N_256,In_4145);
xnor U2413 (N_2413,In_2750,N_2237);
or U2414 (N_2414,N_1952,N_227);
or U2415 (N_2415,In_3361,In_3622);
and U2416 (N_2416,N_1721,N_612);
xnor U2417 (N_2417,N_1866,In_1455);
and U2418 (N_2418,N_1022,N_198);
nor U2419 (N_2419,In_1977,N_1949);
xnor U2420 (N_2420,N_2221,In_2202);
nand U2421 (N_2421,In_977,In_329);
nor U2422 (N_2422,N_1181,N_1998);
or U2423 (N_2423,N_2181,In_4001);
nand U2424 (N_2424,In_1134,In_1737);
nor U2425 (N_2425,In_692,In_363);
or U2426 (N_2426,In_2833,N_2152);
or U2427 (N_2427,In_2930,N_1058);
nor U2428 (N_2428,In_4800,N_896);
nand U2429 (N_2429,In_561,N_2054);
nor U2430 (N_2430,N_1433,In_2966);
nor U2431 (N_2431,In_305,In_3422);
xnor U2432 (N_2432,N_2185,In_3557);
nor U2433 (N_2433,In_1557,In_437);
or U2434 (N_2434,N_360,N_1679);
nand U2435 (N_2435,In_548,N_1176);
xor U2436 (N_2436,In_3738,N_404);
nor U2437 (N_2437,In_4085,N_1579);
xnor U2438 (N_2438,In_564,In_421);
nand U2439 (N_2439,N_513,N_1001);
nor U2440 (N_2440,N_858,In_337);
nand U2441 (N_2441,N_1754,In_989);
and U2442 (N_2442,In_958,N_2098);
nor U2443 (N_2443,In_3644,In_4635);
or U2444 (N_2444,N_2100,N_2189);
nor U2445 (N_2445,In_2348,N_750);
nand U2446 (N_2446,In_2489,In_1006);
xor U2447 (N_2447,In_947,In_4832);
and U2448 (N_2448,N_2136,In_3173);
or U2449 (N_2449,In_2996,In_3923);
nand U2450 (N_2450,N_1997,N_2016);
nand U2451 (N_2451,In_2870,In_379);
xor U2452 (N_2452,In_568,N_1138);
nand U2453 (N_2453,N_1733,In_4820);
nand U2454 (N_2454,In_225,N_1713);
xnor U2455 (N_2455,N_1984,In_396);
and U2456 (N_2456,N_789,N_1108);
xor U2457 (N_2457,In_1309,In_2283);
or U2458 (N_2458,In_664,N_1525);
nor U2459 (N_2459,N_778,In_4864);
nand U2460 (N_2460,In_3285,N_604);
nor U2461 (N_2461,N_1382,In_43);
and U2462 (N_2462,N_512,N_1088);
nand U2463 (N_2463,N_1298,In_898);
xor U2464 (N_2464,N_624,N_431);
nand U2465 (N_2465,In_4544,N_1712);
or U2466 (N_2466,In_618,In_3087);
nand U2467 (N_2467,In_4427,In_3687);
or U2468 (N_2468,In_4024,N_1851);
nand U2469 (N_2469,N_1468,N_304);
and U2470 (N_2470,In_4875,In_1103);
xor U2471 (N_2471,N_2063,N_1873);
or U2472 (N_2472,N_1672,In_1162);
or U2473 (N_2473,In_935,N_1667);
nand U2474 (N_2474,In_3736,In_2808);
and U2475 (N_2475,In_3633,In_1390);
nand U2476 (N_2476,N_1961,In_1710);
nor U2477 (N_2477,In_2595,In_1789);
nand U2478 (N_2478,In_2573,In_655);
or U2479 (N_2479,N_1931,In_4334);
nand U2480 (N_2480,In_1644,In_3091);
xor U2481 (N_2481,In_945,N_1128);
or U2482 (N_2482,N_2013,In_4705);
and U2483 (N_2483,In_802,In_1864);
xnor U2484 (N_2484,In_3252,N_2126);
xor U2485 (N_2485,In_248,N_1595);
and U2486 (N_2486,N_1730,N_769);
nand U2487 (N_2487,N_1254,N_1788);
and U2488 (N_2488,N_2166,N_1337);
nor U2489 (N_2489,In_1436,N_1607);
nand U2490 (N_2490,In_3560,N_2113);
xnor U2491 (N_2491,In_759,In_3193);
or U2492 (N_2492,In_3959,N_1907);
nor U2493 (N_2493,N_1801,N_1508);
nand U2494 (N_2494,N_471,In_3825);
or U2495 (N_2495,In_2948,N_1078);
nand U2496 (N_2496,In_4867,N_226);
nand U2497 (N_2497,In_2309,In_4172);
and U2498 (N_2498,In_3179,In_391);
and U2499 (N_2499,In_2241,In_4682);
nor U2500 (N_2500,In_619,N_2256);
xnor U2501 (N_2501,N_1034,N_2353);
nand U2502 (N_2502,N_2161,N_2276);
xnor U2503 (N_2503,In_376,In_1311);
and U2504 (N_2504,N_394,In_3388);
xnor U2505 (N_2505,In_4879,N_2486);
nand U2506 (N_2506,N_1835,In_4406);
xnor U2507 (N_2507,In_2385,In_4508);
and U2508 (N_2508,In_4116,N_1699);
nor U2509 (N_2509,N_1723,In_2064);
or U2510 (N_2510,In_288,N_2119);
and U2511 (N_2511,N_1292,N_509);
nor U2512 (N_2512,N_2489,N_1076);
and U2513 (N_2513,In_4532,In_4395);
nand U2514 (N_2514,In_118,N_376);
and U2515 (N_2515,N_2006,In_4150);
nand U2516 (N_2516,N_1947,In_585);
nand U2517 (N_2517,In_438,N_2039);
nor U2518 (N_2518,In_1685,In_4237);
nor U2519 (N_2519,In_2229,N_2385);
nand U2520 (N_2520,N_934,In_2777);
and U2521 (N_2521,N_1251,N_2029);
nand U2522 (N_2522,N_2193,In_3582);
xnor U2523 (N_2523,In_3002,In_1233);
nand U2524 (N_2524,In_4240,In_639);
and U2525 (N_2525,N_766,In_40);
xnor U2526 (N_2526,In_3380,In_3316);
or U2527 (N_2527,N_2069,N_428);
nand U2528 (N_2528,N_1979,In_2561);
nor U2529 (N_2529,In_2686,N_1171);
and U2530 (N_2530,N_1157,In_1440);
or U2531 (N_2531,In_2212,N_1860);
or U2532 (N_2532,N_2441,In_1383);
or U2533 (N_2533,In_4393,N_1956);
nand U2534 (N_2534,In_1779,In_3177);
and U2535 (N_2535,N_1075,In_2706);
nor U2536 (N_2536,N_2410,In_1208);
nor U2537 (N_2537,In_4265,N_1654);
nand U2538 (N_2538,N_88,N_1934);
xnor U2539 (N_2539,In_3205,N_1926);
nor U2540 (N_2540,N_2482,In_2992);
and U2541 (N_2541,N_1948,N_2252);
nand U2542 (N_2542,In_3551,In_4010);
nand U2543 (N_2543,N_1568,N_510);
and U2544 (N_2544,In_1889,N_1187);
or U2545 (N_2545,In_4658,In_2973);
or U2546 (N_2546,N_2066,In_3080);
nand U2547 (N_2547,In_4456,N_1551);
and U2548 (N_2548,In_273,In_3326);
nor U2549 (N_2549,N_1827,N_1283);
or U2550 (N_2550,N_2150,In_1144);
nand U2551 (N_2551,In_501,In_1056);
nor U2552 (N_2552,In_3755,N_1036);
or U2553 (N_2553,N_538,In_54);
or U2554 (N_2554,In_2918,N_1799);
nand U2555 (N_2555,N_2415,N_1632);
nor U2556 (N_2556,N_2023,In_404);
nor U2557 (N_2557,N_554,In_3506);
nand U2558 (N_2558,N_1977,In_1513);
nand U2559 (N_2559,N_1208,N_1864);
and U2560 (N_2560,In_2071,N_1209);
nand U2561 (N_2561,N_1344,In_4955);
and U2562 (N_2562,In_3704,N_1478);
nand U2563 (N_2563,N_1333,N_2398);
nand U2564 (N_2564,N_1795,In_3658);
xnor U2565 (N_2565,In_3601,N_1561);
nor U2566 (N_2566,In_961,N_1284);
and U2567 (N_2567,In_432,N_0);
nor U2568 (N_2568,N_957,N_2437);
xor U2569 (N_2569,N_796,In_2814);
and U2570 (N_2570,In_4501,In_1232);
xor U2571 (N_2571,In_3549,N_2363);
and U2572 (N_2572,N_1681,N_1887);
and U2573 (N_2573,N_1740,In_727);
nand U2574 (N_2574,N_2429,In_1398);
xor U2575 (N_2575,N_157,In_2953);
or U2576 (N_2576,In_456,In_1846);
and U2577 (N_2577,In_3713,N_2078);
or U2578 (N_2578,N_2315,In_1143);
xor U2579 (N_2579,In_3010,In_3207);
nand U2580 (N_2580,N_1753,N_266);
nor U2581 (N_2581,In_1549,N_1726);
xor U2582 (N_2582,N_2381,In_3857);
nand U2583 (N_2583,In_115,N_1807);
and U2584 (N_2584,In_3568,N_623);
nand U2585 (N_2585,N_2233,In_3902);
xnor U2586 (N_2586,In_3545,N_2082);
and U2587 (N_2587,N_2490,In_1812);
and U2588 (N_2588,In_3859,N_194);
nand U2589 (N_2589,In_134,In_2743);
xor U2590 (N_2590,In_2421,N_1865);
nand U2591 (N_2591,N_1184,N_2137);
or U2592 (N_2592,N_657,N_1624);
nor U2593 (N_2593,N_1845,In_1028);
nor U2594 (N_2594,N_1763,N_2142);
and U2595 (N_2595,N_2038,In_3363);
nand U2596 (N_2596,In_1587,N_1085);
nor U2597 (N_2597,In_2590,In_2047);
nor U2598 (N_2598,In_236,N_2265);
xnor U2599 (N_2599,In_3044,N_2405);
xnor U2600 (N_2600,In_950,N_2076);
and U2601 (N_2601,N_2047,In_1486);
xnor U2602 (N_2602,N_1841,In_2763);
or U2603 (N_2603,In_3507,In_3021);
nand U2604 (N_2604,N_1776,N_2107);
nand U2605 (N_2605,N_2447,In_2690);
or U2606 (N_2606,In_3840,In_789);
nor U2607 (N_2607,N_2057,In_4273);
nor U2608 (N_2608,In_4674,N_280);
xor U2609 (N_2609,N_1536,N_650);
and U2610 (N_2610,N_1299,N_774);
nor U2611 (N_2611,N_1778,In_105);
xor U2612 (N_2612,N_2288,N_1324);
xnor U2613 (N_2613,In_4321,In_1260);
nand U2614 (N_2614,In_3532,N_2449);
and U2615 (N_2615,In_4455,In_3186);
nor U2616 (N_2616,In_4351,In_120);
and U2617 (N_2617,In_689,N_1338);
nand U2618 (N_2618,N_2304,N_1746);
or U2619 (N_2619,In_4398,In_1301);
nand U2620 (N_2620,In_2683,N_94);
xnor U2621 (N_2621,In_2986,N_2406);
xnor U2622 (N_2622,N_1217,N_2401);
nand U2623 (N_2623,In_1969,In_1335);
nor U2624 (N_2624,N_492,N_1612);
nand U2625 (N_2625,N_967,In_3501);
and U2626 (N_2626,N_2278,In_507);
and U2627 (N_2627,N_1781,In_4247);
nand U2628 (N_2628,In_3483,N_1278);
nor U2629 (N_2629,N_1875,In_3910);
nand U2630 (N_2630,In_4258,N_14);
xnor U2631 (N_2631,In_1785,N_1953);
nor U2632 (N_2632,N_535,In_592);
and U2633 (N_2633,In_1470,In_4329);
nand U2634 (N_2634,N_1538,N_1942);
nor U2635 (N_2635,N_1790,N_2104);
xnor U2636 (N_2636,In_1747,N_1874);
xor U2637 (N_2637,In_4834,In_4367);
nand U2638 (N_2638,In_4822,In_2127);
nor U2639 (N_2639,N_1577,N_1139);
and U2640 (N_2640,In_4029,N_2494);
nor U2641 (N_2641,N_2071,N_2080);
xor U2642 (N_2642,N_1481,N_2481);
and U2643 (N_2643,N_2268,N_2418);
nand U2644 (N_2644,N_791,In_308);
nand U2645 (N_2645,N_1613,N_1543);
nand U2646 (N_2646,N_1844,N_402);
nand U2647 (N_2647,In_1249,N_2167);
or U2648 (N_2648,N_859,N_1093);
or U2649 (N_2649,N_1087,In_900);
and U2650 (N_2650,In_3722,N_262);
nor U2651 (N_2651,In_4921,N_1163);
or U2652 (N_2652,In_1083,N_767);
or U2653 (N_2653,N_1916,N_1664);
nor U2654 (N_2654,N_2302,In_1919);
xor U2655 (N_2655,N_1562,N_2041);
nand U2656 (N_2656,N_821,In_3712);
xor U2657 (N_2657,In_4304,N_1048);
nor U2658 (N_2658,N_2327,In_398);
or U2659 (N_2659,In_3421,In_3976);
nor U2660 (N_2660,In_229,N_2197);
nor U2661 (N_2661,In_3050,N_2109);
nor U2662 (N_2662,N_2149,In_2467);
or U2663 (N_2663,N_1518,N_453);
and U2664 (N_2664,N_601,N_584);
and U2665 (N_2665,In_2891,N_1358);
nand U2666 (N_2666,In_4525,N_808);
or U2667 (N_2667,In_3003,N_130);
or U2668 (N_2668,N_2232,N_1641);
nor U2669 (N_2669,In_3449,N_553);
or U2670 (N_2670,N_908,In_2861);
xor U2671 (N_2671,In_1526,N_536);
nand U2672 (N_2672,In_447,In_701);
nand U2673 (N_2673,In_1888,In_1084);
nand U2674 (N_2674,In_3527,N_2);
or U2675 (N_2675,N_1541,N_2366);
and U2676 (N_2676,In_3899,In_1723);
nor U2677 (N_2677,In_4180,In_346);
or U2678 (N_2678,N_2050,N_1818);
nand U2679 (N_2679,In_4431,N_1601);
xor U2680 (N_2680,N_1528,N_1488);
nor U2681 (N_2681,N_842,N_1560);
nor U2682 (N_2682,In_3909,N_1792);
xor U2683 (N_2683,N_1722,In_820);
and U2684 (N_2684,N_149,In_1429);
or U2685 (N_2685,N_2289,In_929);
or U2686 (N_2686,N_2343,N_1806);
nor U2687 (N_2687,N_101,N_1202);
or U2688 (N_2688,N_1155,N_678);
nand U2689 (N_2689,In_3339,In_2687);
nand U2690 (N_2690,In_1421,N_1400);
or U2691 (N_2691,In_4664,In_4391);
xnor U2692 (N_2692,N_2143,In_156);
nor U2693 (N_2693,N_1963,N_2022);
nand U2694 (N_2694,In_514,N_2436);
or U2695 (N_2695,In_1937,In_4522);
xnor U2696 (N_2696,In_874,N_1766);
nand U2697 (N_2697,In_800,In_925);
nand U2698 (N_2698,In_3979,In_3042);
and U2699 (N_2699,In_4625,In_3974);
nand U2700 (N_2700,N_829,In_1113);
nand U2701 (N_2701,N_768,N_1281);
xnor U2702 (N_2702,In_4971,N_947);
and U2703 (N_2703,N_2065,In_2730);
nor U2704 (N_2704,In_2443,In_1025);
and U2705 (N_2705,N_2384,N_2218);
nor U2706 (N_2706,In_2045,N_2246);
and U2707 (N_2707,N_2184,N_1405);
or U2708 (N_2708,In_4505,N_969);
and U2709 (N_2709,In_3954,N_1245);
and U2710 (N_2710,N_2070,In_1159);
nand U2711 (N_2711,N_1148,N_2450);
nand U2712 (N_2712,N_2371,In_2457);
or U2713 (N_2713,N_1327,N_1701);
nor U2714 (N_2714,In_37,N_1936);
nand U2715 (N_2715,N_1894,In_3457);
and U2716 (N_2716,In_3307,N_407);
or U2717 (N_2717,N_1785,In_1277);
nor U2718 (N_2718,In_4407,N_2479);
and U2719 (N_2719,N_1317,N_1732);
nand U2720 (N_2720,N_1204,N_1223);
or U2721 (N_2721,In_1896,N_2020);
and U2722 (N_2722,N_1839,In_1859);
xor U2723 (N_2723,In_2988,N_2175);
nor U2724 (N_2724,N_1182,N_2386);
xnor U2725 (N_2725,N_1869,In_1987);
nor U2726 (N_2726,In_321,N_1837);
nor U2727 (N_2727,In_3565,N_1026);
or U2728 (N_2728,N_1457,In_3873);
nor U2729 (N_2729,N_76,N_2469);
xnor U2730 (N_2730,N_2010,N_986);
nor U2731 (N_2731,In_1167,N_255);
and U2732 (N_2732,In_702,In_4676);
xnor U2733 (N_2733,In_4557,In_2872);
or U2734 (N_2734,N_2024,In_662);
or U2735 (N_2735,N_1506,In_4121);
nand U2736 (N_2736,N_943,N_1113);
nand U2737 (N_2737,In_2883,N_412);
nand U2738 (N_2738,In_928,N_927);
and U2739 (N_2739,In_2824,In_1049);
nand U2740 (N_2740,In_2910,In_4288);
nand U2741 (N_2741,In_4143,In_1657);
xnor U2742 (N_2742,N_642,In_4433);
xor U2743 (N_2743,N_1922,In_4357);
nor U2744 (N_2744,In_1903,N_1593);
xnor U2745 (N_2745,In_347,In_4909);
nand U2746 (N_2746,In_1066,In_4079);
nand U2747 (N_2747,In_4714,In_887);
nor U2748 (N_2748,In_1477,In_1108);
and U2749 (N_2749,N_2365,N_2427);
and U2750 (N_2750,In_3693,N_517);
xor U2751 (N_2751,N_1980,In_2112);
or U2752 (N_2752,N_1524,In_2570);
nand U2753 (N_2753,N_2130,N_1605);
nand U2754 (N_2754,In_3714,N_1566);
and U2755 (N_2755,N_1638,In_975);
or U2756 (N_2756,In_1543,N_782);
and U2757 (N_2757,In_3526,N_1151);
xor U2758 (N_2758,In_4369,N_416);
or U2759 (N_2759,In_3891,In_3969);
nor U2760 (N_2760,N_482,N_559);
nand U2761 (N_2761,N_1760,In_3379);
nor U2762 (N_2762,In_2106,N_2009);
and U2763 (N_2763,In_4590,In_4330);
xnor U2764 (N_2764,In_4873,N_1636);
and U2765 (N_2765,N_2027,N_506);
nor U2766 (N_2766,N_2646,N_2513);
nand U2767 (N_2767,N_2480,N_2446);
xor U2768 (N_2768,In_3918,N_1028);
xnor U2769 (N_2769,N_1501,N_2305);
and U2770 (N_2770,In_3350,N_2688);
nand U2771 (N_2771,N_2585,N_2543);
nor U2772 (N_2772,In_4094,In_645);
nand U2773 (N_2773,N_2348,N_918);
and U2774 (N_2774,In_3244,N_2421);
xnor U2775 (N_2775,In_4725,N_2208);
xnor U2776 (N_2776,N_2570,In_1497);
and U2777 (N_2777,In_920,In_302);
xnor U2778 (N_2778,N_2008,N_1982);
nand U2779 (N_2779,N_2257,N_2428);
nor U2780 (N_2780,N_2466,N_1146);
and U2781 (N_2781,N_2049,In_1883);
xnor U2782 (N_2782,N_2651,In_2146);
or U2783 (N_2783,N_2528,N_1995);
xor U2784 (N_2784,In_1617,In_4526);
nand U2785 (N_2785,N_2296,In_2287);
xor U2786 (N_2786,N_2467,N_2615);
and U2787 (N_2787,N_2204,N_1889);
xor U2788 (N_2788,N_183,In_4876);
nand U2789 (N_2789,In_316,N_405);
or U2790 (N_2790,N_732,In_674);
nand U2791 (N_2791,N_666,In_4086);
nor U2792 (N_2792,In_90,N_1466);
nand U2793 (N_2793,N_1531,N_793);
or U2794 (N_2794,N_1677,N_1884);
nand U2795 (N_2795,N_1599,N_1682);
or U2796 (N_2796,In_1316,In_2640);
nor U2797 (N_2797,N_2158,N_2004);
nor U2798 (N_2798,N_2502,In_4328);
nand U2799 (N_2799,In_3199,In_1);
xnor U2800 (N_2800,In_392,N_1854);
xnor U2801 (N_2801,In_97,In_4669);
or U2802 (N_2802,N_1895,In_374);
and U2803 (N_2803,In_3208,N_2477);
nand U2804 (N_2804,N_2367,N_2308);
and U2805 (N_2805,N_1535,N_1035);
and U2806 (N_2806,In_3378,In_3347);
xor U2807 (N_2807,N_2317,N_1846);
nand U2808 (N_2808,N_1888,In_1074);
nor U2809 (N_2809,N_688,N_2190);
or U2810 (N_2810,In_747,N_1378);
nor U2811 (N_2811,In_1228,N_1280);
nand U2812 (N_2812,In_3492,In_3024);
nor U2813 (N_2813,In_4706,In_3306);
or U2814 (N_2814,In_1428,N_1582);
xnor U2815 (N_2815,N_2461,N_2419);
xnor U2816 (N_2816,In_1575,N_2723);
and U2817 (N_2817,In_1638,N_1355);
or U2818 (N_2818,N_1779,In_4327);
or U2819 (N_2819,In_3986,In_186);
xor U2820 (N_2820,N_2713,N_2444);
or U2821 (N_2821,N_374,In_1161);
nand U2822 (N_2822,In_2247,N_2640);
nor U2823 (N_2823,In_3922,N_1464);
and U2824 (N_2824,In_1671,N_1290);
xor U2825 (N_2825,In_1928,In_1878);
and U2826 (N_2826,In_4735,N_1564);
nor U2827 (N_2827,In_2761,N_772);
nand U2828 (N_2828,N_1346,In_852);
and U2829 (N_2829,In_3756,In_4295);
or U2830 (N_2830,In_1552,N_1891);
and U2831 (N_2831,In_4837,In_125);
nor U2832 (N_2832,In_4660,N_345);
nand U2833 (N_2833,N_2351,N_2639);
nand U2834 (N_2834,In_616,N_1007);
or U2835 (N_2835,N_1165,N_2483);
nand U2836 (N_2836,N_1742,N_1027);
and U2837 (N_2837,In_2845,In_4554);
and U2838 (N_2838,In_4870,N_1986);
xor U2839 (N_2839,In_4300,N_1883);
xor U2840 (N_2840,In_3921,N_2209);
nor U2841 (N_2841,N_42,In_1862);
or U2842 (N_2842,N_367,N_1246);
xnor U2843 (N_2843,In_4091,N_1862);
nor U2844 (N_2844,In_538,N_2676);
nand U2845 (N_2845,In_3352,N_2705);
and U2846 (N_2846,In_1088,N_1594);
and U2847 (N_2847,In_2844,N_2262);
xor U2848 (N_2848,In_1100,In_2090);
or U2849 (N_2849,N_2283,In_2909);
xnor U2850 (N_2850,N_2045,In_3138);
nor U2851 (N_2851,N_1451,In_2410);
xnor U2852 (N_2852,In_3043,In_724);
or U2853 (N_2853,N_933,In_1912);
nand U2854 (N_2854,N_1394,N_217);
or U2855 (N_2855,In_931,In_4000);
xnor U2856 (N_2856,In_3783,N_1442);
nor U2857 (N_2857,N_1919,In_3962);
or U2858 (N_2858,In_4855,N_1719);
nand U2859 (N_2859,N_619,In_3519);
xor U2860 (N_2860,In_2648,N_41);
xnor U2861 (N_2861,N_2352,N_2567);
or U2862 (N_2862,N_2347,N_2387);
xor U2863 (N_2863,N_348,N_1830);
xnor U2864 (N_2864,N_1279,N_1500);
xor U2865 (N_2865,N_2292,In_3333);
or U2866 (N_2866,N_1603,In_1242);
and U2867 (N_2867,In_2475,N_609);
or U2868 (N_2868,N_743,N_2402);
or U2869 (N_2869,N_307,N_2569);
nand U2870 (N_2870,N_2644,In_1465);
and U2871 (N_2871,N_2631,In_380);
nor U2872 (N_2872,N_2354,N_1116);
nand U2873 (N_2873,N_867,In_3315);
and U2874 (N_2874,N_704,In_1341);
nor U2875 (N_2875,In_4386,N_2379);
or U2876 (N_2876,In_1223,In_1473);
or U2877 (N_2877,In_1487,In_1974);
xnor U2878 (N_2878,N_2583,In_1971);
nand U2879 (N_2879,In_3029,N_790);
nand U2880 (N_2880,N_2226,N_2726);
or U2881 (N_2881,N_1241,N_1273);
nor U2882 (N_2882,N_1772,N_128);
nand U2883 (N_2883,In_1251,N_1655);
and U2884 (N_2884,In_1763,N_1110);
nand U2885 (N_2885,N_871,N_1757);
nor U2886 (N_2886,N_755,N_2061);
xnor U2887 (N_2887,N_719,In_3188);
nor U2888 (N_2888,N_1329,N_1621);
nor U2889 (N_2889,N_2430,In_4126);
nand U2890 (N_2890,N_1519,In_4266);
or U2891 (N_2891,In_1601,N_1135);
nand U2892 (N_2892,N_2509,N_2620);
or U2893 (N_2893,In_3684,In_3791);
and U2894 (N_2894,N_813,In_2182);
and U2895 (N_2895,N_392,N_2689);
nand U2896 (N_2896,N_875,N_2170);
xor U2897 (N_2897,N_2719,In_2371);
xor U2898 (N_2898,N_2416,N_1060);
xor U2899 (N_2899,In_1255,In_2606);
nor U2900 (N_2900,N_1049,In_2266);
nor U2901 (N_2901,N_1029,N_2090);
or U2902 (N_2902,N_2452,N_1974);
or U2903 (N_2903,N_2321,In_2487);
or U2904 (N_2904,In_2412,In_936);
and U2905 (N_2905,N_1272,In_2828);
xor U2906 (N_2906,N_900,In_1823);
or U2907 (N_2907,N_2508,N_1890);
nand U2908 (N_2908,N_1886,In_3897);
nand U2909 (N_2909,N_816,In_4372);
nor U2910 (N_2910,In_4504,N_296);
and U2911 (N_2911,In_562,N_2389);
or U2912 (N_2912,In_2055,In_1910);
and U2913 (N_2913,N_2659,N_2128);
xor U2914 (N_2914,In_4418,N_2319);
and U2915 (N_2915,N_1413,In_3415);
nor U2916 (N_2916,In_743,In_2772);
and U2917 (N_2917,N_1032,In_579);
xnor U2918 (N_2918,In_1505,N_1652);
or U2919 (N_2919,N_1809,N_2241);
xor U2920 (N_2920,In_1838,N_2749);
and U2921 (N_2921,In_2341,N_2698);
xnor U2922 (N_2922,N_2294,N_2420);
or U2923 (N_2923,N_1848,N_645);
nand U2924 (N_2924,In_4609,N_1066);
and U2925 (N_2925,N_2518,N_1122);
nor U2926 (N_2926,In_66,In_1766);
and U2927 (N_2927,In_1376,In_1160);
or U2928 (N_2928,N_2340,In_1656);
nand U2929 (N_2929,In_149,N_1695);
xor U2930 (N_2930,In_2026,In_4996);
nor U2931 (N_2931,N_1816,In_2464);
and U2932 (N_2932,In_2691,N_1083);
and U2933 (N_2933,In_2577,N_1867);
and U2934 (N_2934,N_2298,In_2853);
xor U2935 (N_2935,In_2682,In_3934);
xnor U2936 (N_2936,N_151,N_1387);
or U2937 (N_2937,N_2242,N_215);
nor U2938 (N_2938,N_1390,N_1791);
nor U2939 (N_2939,N_1107,N_479);
nand U2940 (N_2940,N_385,N_830);
nor U2941 (N_2941,N_1749,In_1420);
nand U2942 (N_2942,N_2442,N_2099);
nor U2943 (N_2943,In_4104,N_1815);
nor U2944 (N_2944,In_306,In_3498);
or U2945 (N_2945,N_2163,N_1856);
or U2946 (N_2946,In_3808,N_2576);
nor U2947 (N_2947,In_813,N_2716);
nand U2948 (N_2948,N_2191,N_786);
or U2949 (N_2949,N_2445,In_1821);
or U2950 (N_2950,N_1465,N_2103);
nand U2951 (N_2951,In_2231,N_2733);
xor U2952 (N_2952,N_1221,N_1274);
or U2953 (N_2953,In_1460,N_2597);
or U2954 (N_2954,N_123,N_1365);
xor U2955 (N_2955,N_2350,In_331);
xnor U2956 (N_2956,In_628,N_1250);
and U2957 (N_2957,N_1042,N_2369);
nor U2958 (N_2958,N_339,N_2504);
xnor U2959 (N_2959,In_2703,N_1673);
nand U2960 (N_2960,In_3153,In_985);
nor U2961 (N_2961,In_2710,N_2656);
and U2962 (N_2962,N_2413,N_2694);
xor U2963 (N_2963,N_1439,N_2033);
xnor U2964 (N_2964,In_4814,In_3569);
and U2965 (N_2965,N_2684,In_1472);
nor U2966 (N_2966,In_3241,In_891);
nand U2967 (N_2967,N_1101,N_230);
nand U2968 (N_2968,In_2420,N_2102);
nand U2969 (N_2969,In_4785,In_2091);
or U2970 (N_2970,N_1429,N_2693);
or U2971 (N_2971,In_1568,In_623);
nor U2972 (N_2972,N_1440,N_2291);
or U2973 (N_2973,N_1277,In_480);
nand U2974 (N_2974,N_2171,N_838);
nand U2975 (N_2975,N_1796,In_1041);
and U2976 (N_2976,N_1708,In_1236);
nand U2977 (N_2977,N_50,N_1392);
xor U2978 (N_2978,In_4975,N_119);
nand U2979 (N_2979,N_352,N_2234);
nor U2980 (N_2980,In_3798,N_2703);
or U2981 (N_2981,In_4670,In_1117);
and U2982 (N_2982,In_1492,In_617);
nand U2983 (N_2983,In_271,N_2132);
nor U2984 (N_2984,In_488,N_1503);
nand U2985 (N_2985,In_439,N_883);
nor U2986 (N_2986,N_2501,N_1555);
or U2987 (N_2987,N_718,In_3510);
or U2988 (N_2988,In_39,In_3280);
or U2989 (N_2989,N_2619,N_515);
or U2990 (N_2990,N_1406,In_2933);
xnor U2991 (N_2991,In_2085,N_206);
nor U2992 (N_2992,In_3953,In_1652);
xor U2993 (N_2993,In_1030,N_1859);
nand U2994 (N_2994,In_1735,N_2637);
nand U2995 (N_2995,N_2529,N_1758);
or U2996 (N_2996,N_2361,N_1396);
xnor U2997 (N_2997,N_2692,N_240);
nand U2998 (N_2998,N_4,In_1380);
xnor U2999 (N_2999,In_338,In_3943);
xor U3000 (N_3000,N_2546,N_2512);
nor U3001 (N_3001,In_1454,In_2139);
nor U3002 (N_3002,N_1222,N_1238);
nand U3003 (N_3003,In_2094,N_879);
nand U3004 (N_3004,In_2268,In_527);
and U3005 (N_3005,N_2537,N_2145);
nor U3006 (N_3006,In_2338,N_1550);
xor U3007 (N_3007,In_3277,N_2927);
nor U3008 (N_3008,N_614,In_3634);
and U3009 (N_3009,N_1711,N_572);
and U3010 (N_3010,In_4911,In_1458);
xnor U3011 (N_3011,N_2473,N_2958);
nand U3012 (N_3012,In_4466,N_2877);
nor U3013 (N_3013,N_2710,In_1718);
or U3014 (N_3014,N_2403,N_2571);
or U3015 (N_3015,N_2287,In_3960);
xnor U3016 (N_3016,In_520,N_891);
nor U3017 (N_3017,N_2629,N_1065);
or U3018 (N_3018,N_2032,N_653);
nand U3019 (N_3019,N_1377,N_1206);
and U3020 (N_3020,N_548,In_988);
nand U3021 (N_3021,N_2380,N_2611);
nand U3022 (N_3022,In_4306,In_2391);
and U3023 (N_3023,N_1447,In_987);
or U3024 (N_3024,N_2847,N_1345);
and U3025 (N_3025,In_3907,In_3797);
and U3026 (N_3026,In_1548,N_324);
nor U3027 (N_3027,N_1352,N_1474);
and U3028 (N_3028,N_1782,N_2118);
or U3029 (N_3029,N_825,In_2835);
nand U3030 (N_3030,N_2770,N_1738);
and U3031 (N_3031,N_2220,In_633);
xnor U3032 (N_3032,N_1315,N_277);
nand U3033 (N_3033,N_2206,In_2850);
nand U3034 (N_3034,N_2541,N_920);
xor U3035 (N_3035,N_2776,In_465);
xnor U3036 (N_3036,N_2876,N_1702);
and U3037 (N_3037,N_2344,N_622);
nand U3038 (N_3038,N_1225,In_2693);
nor U3039 (N_3039,N_1363,N_2932);
nor U3040 (N_3040,N_1467,N_1767);
nor U3041 (N_3041,In_1190,N_754);
nand U3042 (N_3042,N_2423,N_758);
or U3043 (N_3043,N_1473,N_2476);
nor U3044 (N_3044,In_3799,In_154);
nor U3045 (N_3045,N_1752,N_2785);
xor U3046 (N_3046,N_18,N_1389);
nand U3047 (N_3047,N_2133,N_2840);
or U3048 (N_3048,N_1201,In_1588);
nand U3049 (N_3049,N_2563,N_1693);
or U3050 (N_3050,In_4567,N_2106);
nand U3051 (N_3051,N_892,N_1923);
nor U3052 (N_3052,In_2101,In_3882);
or U3053 (N_3053,N_2231,N_2125);
and U3054 (N_3054,N_697,In_2221);
or U3055 (N_3055,N_2712,N_2593);
xor U3056 (N_3056,N_1694,In_1746);
and U3057 (N_3057,N_2108,In_986);
xor U3058 (N_3058,N_2338,N_1266);
or U3059 (N_3059,In_2523,N_2530);
and U3060 (N_3060,N_1996,In_1517);
nand U3061 (N_3061,In_3497,N_1572);
nor U3062 (N_3062,N_2000,N_2925);
or U3063 (N_3063,N_2899,N_2805);
or U3064 (N_3064,N_2263,N_2858);
nor U3065 (N_3065,In_2964,In_1597);
and U3066 (N_3066,N_2674,N_1804);
or U3067 (N_3067,N_1074,In_1554);
xnor U3068 (N_3068,N_1341,N_529);
nor U3069 (N_3069,N_2424,In_2381);
and U3070 (N_3070,N_1762,In_3338);
or U3071 (N_3071,N_2168,In_2048);
or U3072 (N_3072,N_2173,N_2979);
and U3073 (N_3073,N_1640,N_2971);
xor U3074 (N_3074,N_2696,N_2083);
or U3075 (N_3075,In_3517,N_2536);
nand U3076 (N_3076,N_2658,In_2604);
xnor U3077 (N_3077,N_1622,N_2545);
nor U3078 (N_3078,In_594,In_2235);
nor U3079 (N_3079,In_913,N_2349);
and U3080 (N_3080,N_2154,N_2722);
or U3081 (N_3081,In_1662,N_2028);
nand U3082 (N_3082,In_1219,N_82);
or U3083 (N_3083,N_1933,In_1372);
or U3084 (N_3084,N_2687,N_2824);
nor U3085 (N_3085,N_2664,In_2764);
or U3086 (N_3086,N_1750,In_660);
nor U3087 (N_3087,In_2053,N_2259);
nor U3088 (N_3088,N_2679,N_2604);
or U3089 (N_3089,In_922,N_1322);
nand U3090 (N_3090,In_1879,In_1027);
nor U3091 (N_3091,N_2273,In_4868);
nor U3092 (N_3092,N_2542,N_1533);
and U3093 (N_3093,N_2520,N_2058);
nand U3094 (N_3094,N_2751,N_2857);
and U3095 (N_3095,In_4319,N_2572);
or U3096 (N_3096,N_2610,In_2837);
xnor U3097 (N_3097,N_1239,N_2251);
xnor U3098 (N_3098,N_694,N_1534);
nor U3099 (N_3099,In_3830,N_475);
nand U3100 (N_3100,In_2181,In_3597);
or U3101 (N_3101,N_253,N_2307);
nor U3102 (N_3102,N_836,N_2831);
nand U3103 (N_3103,In_973,N_2909);
or U3104 (N_3104,N_1649,In_303);
nor U3105 (N_3105,N_2946,N_2841);
nor U3106 (N_3106,In_3991,In_2815);
nor U3107 (N_3107,N_1761,N_2661);
or U3108 (N_3108,N_2665,N_2964);
nor U3109 (N_3109,N_1476,N_1644);
xor U3110 (N_3110,N_2750,N_683);
or U3111 (N_3111,N_1955,N_2135);
and U3112 (N_3112,In_4979,In_3817);
nand U3113 (N_3113,N_742,N_2495);
xor U3114 (N_3114,In_3093,N_1755);
and U3115 (N_3115,In_3933,N_2717);
xnor U3116 (N_3116,In_4587,In_80);
nor U3117 (N_3117,In_3651,N_2364);
or U3118 (N_3118,N_2227,In_4388);
xor U3119 (N_3119,N_2370,In_1853);
xnor U3120 (N_3120,N_2531,In_4270);
nor U3121 (N_3121,N_2724,N_427);
nor U3122 (N_3122,N_1964,In_574);
nand U3123 (N_3123,N_1391,N_845);
xor U3124 (N_3124,N_2111,N_2897);
nor U3125 (N_3125,N_2085,N_2433);
and U3126 (N_3126,N_2898,N_2155);
nand U3127 (N_3127,In_3311,N_2001);
nor U3128 (N_3128,In_3077,N_1616);
xor U3129 (N_3129,N_1745,N_798);
xnor U3130 (N_3130,N_2922,N_1232);
and U3131 (N_3131,In_1293,N_1629);
nor U3132 (N_3132,N_1367,N_2600);
and U3133 (N_3133,N_2553,N_2761);
and U3134 (N_3134,In_2904,In_2678);
nor U3135 (N_3135,In_611,N_555);
nand U3136 (N_3136,N_2704,In_3407);
nand U3137 (N_3137,N_1965,In_3377);
or U3138 (N_3138,N_1717,N_2048);
nor U3139 (N_3139,N_1516,In_531);
nand U3140 (N_3140,In_708,N_1052);
xnor U3141 (N_3141,N_2547,In_313);
xnor U3142 (N_3142,N_261,N_2632);
and U3143 (N_3143,N_833,N_2848);
nand U3144 (N_3144,In_979,In_4620);
or U3145 (N_3145,In_1302,In_1109);
nor U3146 (N_3146,In_2922,N_635);
nor U3147 (N_3147,N_1990,In_504);
nand U3148 (N_3148,N_1364,In_3607);
and U3149 (N_3149,In_1194,N_190);
xor U3150 (N_3150,N_2306,In_3038);
nand U3151 (N_3151,In_2456,N_1492);
xnor U3152 (N_3152,N_2153,N_2842);
and U3153 (N_3153,In_3112,In_3524);
nand U3154 (N_3154,In_790,N_2715);
nand U3155 (N_3155,N_2608,In_795);
or U3156 (N_3156,N_1821,N_2573);
nor U3157 (N_3157,In_2372,N_2330);
and U3158 (N_3158,In_3184,In_783);
nor U3159 (N_3159,In_3552,In_474);
nand U3160 (N_3160,N_2737,In_2059);
nor U3161 (N_3161,N_2755,In_643);
and U3162 (N_3162,N_888,In_2337);
xor U3163 (N_3163,In_2530,N_2657);
and U3164 (N_3164,In_4004,N_1081);
and U3165 (N_3165,In_2012,N_2683);
and U3166 (N_3166,N_2127,N_2885);
nand U3167 (N_3167,N_2088,N_390);
nand U3168 (N_3168,N_1219,N_2891);
nor U3169 (N_3169,N_2203,In_2759);
and U3170 (N_3170,In_665,N_2937);
nand U3171 (N_3171,N_2850,N_2667);
nand U3172 (N_3172,N_1911,N_2205);
or U3173 (N_3173,N_2968,In_464);
nand U3174 (N_3174,In_4556,N_1224);
xnor U3175 (N_3175,In_1154,N_2701);
xnor U3176 (N_3176,N_2903,N_2745);
and U3177 (N_3177,N_1756,In_3956);
xor U3178 (N_3178,N_1302,In_4794);
or U3179 (N_3179,N_1526,N_1359);
nor U3180 (N_3180,N_1627,In_1767);
and U3181 (N_3181,In_4905,In_2539);
or U3182 (N_3182,N_2247,In_2753);
and U3183 (N_3183,N_1332,N_2458);
xor U3184 (N_3184,In_1094,N_917);
nor U3185 (N_3185,In_4034,N_2412);
nor U3186 (N_3186,N_1459,N_2641);
xor U3187 (N_3187,In_1451,In_3443);
and U3188 (N_3188,In_4214,In_508);
xor U3189 (N_3189,N_2827,N_2434);
nand U3190 (N_3190,N_2948,N_425);
xnor U3191 (N_3191,N_2414,In_3737);
nand U3192 (N_3192,N_2377,N_2624);
or U3193 (N_3193,N_2883,N_2596);
and U3194 (N_3194,N_1295,In_511);
nand U3195 (N_3195,In_4743,N_2455);
nand U3196 (N_3196,N_1585,N_1511);
and U3197 (N_3197,In_502,N_1137);
nor U3198 (N_3198,N_2550,N_2852);
and U3199 (N_3199,In_2626,In_4146);
and U3200 (N_3200,N_1620,N_2313);
xor U3201 (N_3201,N_1853,N_2522);
and U3202 (N_3202,N_2628,N_58);
nor U3203 (N_3203,N_1819,In_3525);
nand U3204 (N_3204,N_1774,In_2248);
or U3205 (N_3205,N_1349,N_2356);
nor U3206 (N_3206,N_2998,N_2933);
nand U3207 (N_3207,N_1422,In_4681);
nand U3208 (N_3208,In_2664,In_482);
or U3209 (N_3209,N_1985,N_1242);
nand U3210 (N_3210,N_2548,In_270);
nor U3211 (N_3211,N_2863,In_2656);
nand U3212 (N_3212,In_399,N_990);
nor U3213 (N_3213,N_2470,N_1366);
nor U3214 (N_3214,N_2671,N_2763);
xnor U3215 (N_3215,In_3826,In_336);
nand U3216 (N_3216,In_220,In_2917);
and U3217 (N_3217,In_3692,In_3718);
xnor U3218 (N_3218,N_2491,N_2686);
nand U3219 (N_3219,In_3698,N_429);
nand U3220 (N_3220,In_477,N_1736);
nand U3221 (N_3221,N_2984,N_2822);
or U3222 (N_3222,N_2976,N_2559);
nor U3223 (N_3223,In_73,N_2782);
xnor U3224 (N_3224,In_3487,In_2197);
xnor U3225 (N_3225,In_2651,N_2036);
nand U3226 (N_3226,In_109,N_2823);
nor U3227 (N_3227,N_1646,N_2138);
xor U3228 (N_3228,N_2794,In_2971);
xnor U3229 (N_3229,In_580,N_1099);
nand U3230 (N_3230,In_3949,In_3841);
and U3231 (N_3231,In_1810,N_2952);
xnor U3232 (N_3232,N_1118,N_1482);
nor U3233 (N_3233,In_1400,In_0);
nand U3234 (N_3234,N_2147,N_1456);
nor U3235 (N_3235,In_2052,In_1533);
nor U3236 (N_3236,N_2497,N_521);
nor U3237 (N_3237,In_1788,N_2623);
xor U3238 (N_3238,In_2352,N_1193);
nand U3239 (N_3239,N_2264,N_2499);
xor U3240 (N_3240,N_685,In_3616);
nor U3241 (N_3241,N_2535,N_2920);
and U3242 (N_3242,N_1676,In_730);
xor U3243 (N_3243,N_2269,N_2328);
xor U3244 (N_3244,N_2772,N_1814);
and U3245 (N_3245,N_2889,In_2749);
or U3246 (N_3246,In_151,In_1279);
or U3247 (N_3247,In_2696,N_2861);
nand U3248 (N_3248,N_2279,N_2735);
nor U3249 (N_3249,N_146,N_2339);
nor U3250 (N_3250,N_2759,In_1604);
nand U3251 (N_3251,N_2373,N_2074);
nand U3252 (N_3252,N_2341,N_1449);
nand U3253 (N_3253,In_4030,N_1833);
nand U3254 (N_3254,N_3146,N_2120);
nand U3255 (N_3255,N_2829,N_37);
nor U3256 (N_3256,N_2918,N_726);
nor U3257 (N_3257,In_2107,N_295);
or U3258 (N_3258,In_2685,N_913);
and U3259 (N_3259,N_570,In_4205);
xor U3260 (N_3260,In_2698,In_4672);
or U3261 (N_3261,N_2270,N_1547);
or U3262 (N_3262,N_389,N_2580);
nor U3263 (N_3263,In_461,N_3047);
nand U3264 (N_3264,N_2092,N_2165);
nand U3265 (N_3265,N_2818,N_1380);
or U3266 (N_3266,In_2050,N_2837);
nor U3267 (N_3267,N_3115,N_3237);
and U3268 (N_3268,In_14,N_3148);
nor U3269 (N_3269,In_4360,In_1149);
or U3270 (N_3270,In_47,N_2105);
nand U3271 (N_3271,N_2873,N_2337);
nor U3272 (N_3272,N_2556,N_2183);
or U3273 (N_3273,N_1424,N_2101);
or U3274 (N_3274,In_3562,N_2916);
and U3275 (N_3275,In_1243,N_3181);
nor U3276 (N_3276,N_2229,In_1290);
or U3277 (N_3277,In_3890,N_3079);
or U3278 (N_3278,N_2318,N_3144);
nor U3279 (N_3279,In_2367,N_2376);
or U3280 (N_3280,N_1820,N_2779);
and U3281 (N_3281,N_840,N_1404);
nor U3282 (N_3282,N_3130,N_2346);
or U3283 (N_3283,N_2983,In_2131);
and U3284 (N_3284,N_3228,N_188);
xor U3285 (N_3285,N_3192,N_1006);
or U3286 (N_3286,N_3100,N_306);
nand U3287 (N_3287,N_3180,N_3211);
xnor U3288 (N_3288,N_2094,N_2833);
and U3289 (N_3289,N_2274,N_3176);
nor U3290 (N_3290,N_3184,N_3224);
nand U3291 (N_3291,In_2415,In_3054);
xnor U3292 (N_3292,N_2440,N_1914);
nor U3293 (N_3293,In_4392,N_2067);
nand U3294 (N_3294,In_2569,N_2516);
and U3295 (N_3295,N_2322,N_191);
nand U3296 (N_3296,In_4702,N_1935);
and U3297 (N_3297,In_1358,N_689);
nand U3298 (N_3298,In_3999,N_2478);
nor U3299 (N_3299,N_1988,N_2043);
and U3300 (N_3300,In_1062,N_3204);
nor U3301 (N_3301,In_298,In_2118);
or U3302 (N_3302,In_4777,In_4589);
or U3303 (N_3303,N_2267,N_3152);
nor U3304 (N_3304,In_1315,In_3513);
nand U3305 (N_3305,In_3512,In_3639);
nor U3306 (N_3306,In_4934,N_2552);
or U3307 (N_3307,N_1648,In_610);
nor U3308 (N_3308,N_2908,In_3465);
nand U3309 (N_3309,In_4359,N_2031);
nor U3310 (N_3310,In_4131,N_2159);
nand U3311 (N_3311,N_3210,N_2258);
and U3312 (N_3312,N_2663,N_2555);
xor U3313 (N_3313,In_3884,N_2564);
xnor U3314 (N_3314,N_3063,N_1532);
or U3315 (N_3315,N_2506,N_1046);
nor U3316 (N_3316,N_3052,N_1780);
nor U3317 (N_3317,N_2517,In_4046);
nor U3318 (N_3318,N_2662,N_3084);
xor U3319 (N_3319,N_3015,N_3246);
nor U3320 (N_3320,In_2699,N_1959);
and U3321 (N_3321,N_2977,N_1847);
xor U3322 (N_3322,In_2154,N_2718);
xnor U3323 (N_3323,N_2791,In_2571);
or U3324 (N_3324,In_276,N_3214);
nor U3325 (N_3325,N_3153,In_967);
nand U3326 (N_3326,N_3215,N_2172);
xnor U3327 (N_3327,N_235,In_4560);
or U3328 (N_3328,In_3345,N_2582);
or U3329 (N_3329,N_2769,In_3811);
nor U3330 (N_3330,N_1510,N_2975);
xor U3331 (N_3331,In_741,In_1855);
and U3332 (N_3332,N_2738,N_2096);
nand U3333 (N_3333,N_3247,N_2284);
and U3334 (N_3334,N_2093,N_2432);
nand U3335 (N_3335,N_2169,N_159);
or U3336 (N_3336,In_2187,In_657);
or U3337 (N_3337,N_3043,N_2777);
xor U3338 (N_3338,N_3112,In_2347);
xor U3339 (N_3339,N_2320,N_2893);
nand U3340 (N_3340,In_1201,N_792);
nand U3341 (N_3341,N_2116,In_4584);
xor U3342 (N_3342,N_2731,N_1770);
and U3343 (N_3343,In_1863,In_3147);
or U3344 (N_3344,N_1737,N_1031);
and U3345 (N_3345,In_2124,N_3017);
nand U3346 (N_3346,N_2994,N_3046);
nand U3347 (N_3347,N_531,N_1665);
nor U3348 (N_3348,N_242,In_3655);
or U3349 (N_3349,N_1386,N_2141);
xor U3350 (N_3350,In_918,N_2579);
nor U3351 (N_3351,N_2868,N_2768);
nor U3352 (N_3352,N_3177,N_1945);
nand U3353 (N_3353,N_1383,In_2);
nor U3354 (N_3354,N_2709,In_3228);
xor U3355 (N_3355,In_3135,N_3010);
nor U3356 (N_3356,N_3239,N_3206);
nor U3357 (N_3357,N_2362,N_2734);
nor U3358 (N_3358,N_1879,N_2599);
xor U3359 (N_3359,N_2854,N_2956);
nand U3360 (N_3360,N_1906,N_3168);
nor U3361 (N_3361,N_2014,N_1941);
xnor U3362 (N_3362,N_2164,In_4196);
nand U3363 (N_3363,N_1574,N_2222);
or U3364 (N_3364,N_940,N_3229);
nand U3365 (N_3365,In_4100,N_3134);
nor U3366 (N_3366,N_2728,In_4420);
and U3367 (N_3367,N_2935,N_2201);
or U3368 (N_3368,N_2849,N_1910);
xor U3369 (N_3369,N_1183,In_1965);
or U3370 (N_3370,In_475,N_351);
nand U3371 (N_3371,In_2260,In_3436);
xnor U3372 (N_3372,N_2303,N_1734);
xnor U3373 (N_3373,N_1940,N_2230);
nand U3374 (N_3374,In_2003,N_3162);
or U3375 (N_3375,N_2300,N_1132);
nor U3376 (N_3376,N_2562,N_2943);
or U3377 (N_3377,In_798,In_2223);
nand U3378 (N_3378,In_361,N_1030);
nand U3379 (N_3379,N_1751,In_3521);
or U3380 (N_3380,N_1342,In_2174);
xor U3381 (N_3381,N_3095,N_3066);
nor U3382 (N_3382,In_3619,N_2801);
nand U3383 (N_3383,N_3156,N_3022);
and U3384 (N_3384,N_1905,In_4117);
xor U3385 (N_3385,N_3193,In_3341);
nand U3386 (N_3386,In_261,N_3191);
xor U3387 (N_3387,N_2874,N_1403);
nor U3388 (N_3388,In_3073,N_912);
nor U3389 (N_3389,In_20,N_2393);
nor U3390 (N_3390,N_2454,In_4845);
or U3391 (N_3391,In_1749,N_3081);
and U3392 (N_3392,N_47,In_91);
or U3393 (N_3393,N_1709,N_2534);
or U3394 (N_3394,N_3099,In_1111);
nor U3395 (N_3395,N_2989,N_979);
xnor U3396 (N_3396,In_2370,N_1925);
nor U3397 (N_3397,N_2598,N_1487);
xor U3398 (N_3398,N_3026,N_2151);
nor U3399 (N_3399,N_1414,N_2685);
and U3400 (N_3400,N_2266,N_2830);
xnor U3401 (N_3401,In_4639,In_3376);
nor U3402 (N_3402,N_3080,N_40);
nor U3403 (N_3403,N_2730,N_2510);
xor U3404 (N_3404,N_2802,In_3853);
and U3405 (N_3405,N_3050,In_3706);
or U3406 (N_3406,In_309,N_187);
xnor U3407 (N_3407,N_2180,N_1544);
xor U3408 (N_3408,N_2254,In_1886);
nand U3409 (N_3409,N_2261,N_2997);
and U3410 (N_3410,In_192,In_3872);
xor U3411 (N_3411,N_2714,N_2394);
xnor U3412 (N_3412,N_2214,In_4992);
or U3413 (N_3413,N_393,N_2182);
and U3414 (N_3414,N_985,N_2326);
nand U3415 (N_3415,In_3556,N_2669);
xor U3416 (N_3416,In_2148,N_748);
or U3417 (N_3417,N_2627,N_3001);
and U3418 (N_3418,N_3141,In_4815);
nor U3419 (N_3419,In_837,In_2977);
xnor U3420 (N_3420,N_2332,N_2314);
nand U3421 (N_3421,N_3173,N_2140);
or U3422 (N_3422,N_2275,In_2622);
nor U3423 (N_3423,N_2890,In_4852);
and U3424 (N_3424,In_4811,In_1503);
nor U3425 (N_3425,N_2498,N_169);
and U3426 (N_3426,N_2765,N_2253);
or U3427 (N_3427,N_3196,N_2519);
nor U3428 (N_3428,N_2586,In_4603);
nor U3429 (N_3429,N_3109,N_1885);
xnor U3430 (N_3430,N_2280,In_2057);
nand U3431 (N_3431,N_1775,N_1011);
nand U3432 (N_3432,N_2960,In_364);
nor U3433 (N_3433,N_874,N_1615);
or U3434 (N_3434,N_1231,In_4615);
xnor U3435 (N_3435,N_3065,In_714);
and U3436 (N_3436,In_4314,N_2902);
xor U3437 (N_3437,N_2471,In_1811);
xnor U3438 (N_3438,In_3889,In_667);
nand U3439 (N_3439,N_2695,N_607);
nand U3440 (N_3440,In_4656,N_3039);
nor U3441 (N_3441,In_2439,N_3249);
and U3442 (N_3442,N_2995,N_588);
or U3443 (N_3443,N_982,N_2708);
xor U3444 (N_3444,N_1002,N_89);
or U3445 (N_3445,N_3119,N_1797);
nand U3446 (N_3446,In_797,In_4641);
nand U3447 (N_3447,N_55,N_2404);
nor U3448 (N_3448,N_2865,N_2594);
nor U3449 (N_3449,N_2699,N_1009);
and U3450 (N_3450,In_41,In_1982);
nor U3451 (N_3451,N_2248,N_1325);
xnor U3452 (N_3452,N_2634,N_2949);
nor U3453 (N_3453,In_19,In_1203);
or U3454 (N_3454,N_270,N_2792);
nor U3455 (N_3455,N_2295,N_2816);
and U3456 (N_3456,In_4006,In_1640);
nand U3457 (N_3457,N_2162,N_1336);
nand U3458 (N_3458,N_1994,N_2790);
nor U3459 (N_3459,In_2528,N_2196);
or U3460 (N_3460,In_2522,In_3133);
nand U3461 (N_3461,In_823,N_3072);
nor U3462 (N_3462,N_2638,N_1584);
or U3463 (N_3463,In_497,N_2299);
nand U3464 (N_3464,N_3171,N_1455);
xnor U3465 (N_3465,N_3183,N_2468);
nand U3466 (N_3466,In_389,N_585);
nor U3467 (N_3467,N_3202,N_2443);
or U3468 (N_3468,In_765,In_3195);
xor U3469 (N_3469,N_1038,N_279);
nand U3470 (N_3470,In_4434,N_2612);
or U3471 (N_3471,N_2787,In_194);
xor U3472 (N_3472,In_1213,N_1619);
and U3473 (N_3473,N_2938,N_2796);
nor U3474 (N_3474,N_3051,N_2496);
xor U3475 (N_3475,In_3942,N_1831);
xor U3476 (N_3476,N_79,N_1335);
and U3477 (N_3477,N_75,N_2939);
nor U3478 (N_3478,In_2095,N_2702);
xnor U3479 (N_3479,In_4575,In_3820);
xnor U3480 (N_3480,N_2635,N_1789);
xnor U3481 (N_3481,N_2720,N_3241);
nand U3482 (N_3482,In_1741,N_2591);
and U3483 (N_3483,N_2533,N_2382);
xor U3484 (N_3484,In_2989,In_2086);
and U3485 (N_3485,In_4646,N_3203);
or U3486 (N_3486,N_2653,N_2439);
nand U3487 (N_3487,N_2011,N_2965);
nor U3488 (N_3488,N_2219,In_566);
and U3489 (N_3489,N_2575,N_2042);
or U3490 (N_3490,N_38,N_426);
nor U3491 (N_3491,N_1628,N_2677);
nand U3492 (N_3492,N_3233,N_2323);
or U3493 (N_3493,N_2592,In_4810);
xnor U3494 (N_3494,In_4597,In_539);
nand U3495 (N_3495,N_2844,In_4286);
xor U3496 (N_3496,N_2211,N_472);
xnor U3497 (N_3497,In_3592,N_3082);
nand U3498 (N_3498,In_4385,In_3500);
nand U3499 (N_3499,N_2957,N_2560);
xnor U3500 (N_3500,N_118,N_3045);
xnor U3501 (N_3501,In_905,N_3410);
nor U3502 (N_3502,N_3187,N_2400);
xnor U3503 (N_3503,N_2565,N_870);
and U3504 (N_3504,N_3259,N_2391);
xnor U3505 (N_3505,N_951,In_4937);
nor U3506 (N_3506,N_2285,In_3040);
or U3507 (N_3507,N_3336,In_4883);
or U3508 (N_3508,N_2224,N_3258);
nand U3509 (N_3509,In_176,N_2859);
nand U3510 (N_3510,N_3294,N_2117);
or U3511 (N_3511,N_1739,N_1771);
or U3512 (N_3512,N_2725,N_3097);
nor U3513 (N_3513,N_3058,In_3831);
nand U3514 (N_3514,N_1444,N_781);
and U3515 (N_3515,N_2465,In_1736);
and U3516 (N_3516,N_1289,N_3208);
nor U3517 (N_3517,N_3351,N_788);
and U3518 (N_3518,N_857,N_2018);
nor U3519 (N_3519,N_3305,N_3088);
nand U3520 (N_3520,N_2647,N_2334);
nand U3521 (N_3521,N_3276,In_2004);
or U3522 (N_3522,N_2771,N_2764);
nand U3523 (N_3523,N_1929,N_3489);
and U3524 (N_3524,N_17,In_3508);
nor U3525 (N_3525,N_2507,N_2951);
xor U3526 (N_3526,N_563,N_2368);
nor U3527 (N_3527,In_3114,N_3003);
nor U3528 (N_3528,N_3310,N_2521);
xnor U3529 (N_3529,N_1686,N_2249);
nand U3530 (N_3530,In_2781,N_2838);
nor U3531 (N_3531,N_3313,N_2188);
nand U3532 (N_3532,N_2072,In_3105);
or U3533 (N_3533,In_2110,N_1134);
xnor U3534 (N_3534,N_1179,In_2307);
and U3535 (N_3535,N_2811,N_2431);
nor U3536 (N_3536,N_1826,In_1690);
nand U3537 (N_3537,In_2878,N_2293);
and U3538 (N_3538,N_3452,N_3000);
nand U3539 (N_3539,N_1575,N_3316);
or U3540 (N_3540,N_3059,N_3094);
nand U3541 (N_3541,N_2538,N_3289);
or U3542 (N_3542,N_1596,In_223);
and U3543 (N_3543,N_2985,N_3075);
xnor U3544 (N_3544,N_1104,N_889);
nand U3545 (N_3545,N_2870,In_770);
or U3546 (N_3546,N_3423,N_3449);
nor U3547 (N_3547,N_3243,N_2484);
nand U3548 (N_3548,N_3389,N_2485);
xnor U3549 (N_3549,In_3917,N_1715);
or U3550 (N_3550,N_2826,N_3149);
xnor U3551 (N_3551,N_1855,In_4310);
nand U3552 (N_3552,In_4012,N_3238);
nor U3553 (N_3553,N_2904,N_3397);
and U3554 (N_3554,N_2216,N_2892);
xnor U3555 (N_3555,In_1970,N_3290);
nand U3556 (N_3556,In_1237,N_1802);
nor U3557 (N_3557,N_2081,N_2862);
and U3558 (N_3558,N_2462,In_3410);
or U3559 (N_3559,N_2574,In_4645);
nand U3560 (N_3560,In_4470,N_3458);
nand U3561 (N_3561,N_964,N_3462);
or U3562 (N_3562,N_1310,In_3076);
nand U3563 (N_3563,In_1956,In_3395);
nor U3564 (N_3564,N_3455,N_2260);
or U3565 (N_3565,In_3716,N_110);
and U3566 (N_3566,N_3373,In_4636);
xor U3567 (N_3567,In_3454,In_4651);
or U3568 (N_3568,N_3028,N_3212);
nor U3569 (N_3569,In_4103,N_3125);
nand U3570 (N_3570,N_3465,N_3487);
xnor U3571 (N_3571,N_2030,N_1863);
nor U3572 (N_3572,N_1587,N_3275);
xnor U3573 (N_3573,In_3743,N_1553);
and U3574 (N_3574,N_989,N_3231);
xnor U3575 (N_3575,N_861,In_57);
or U3576 (N_3576,In_2406,N_1843);
and U3577 (N_3577,N_3491,In_3172);
or U3578 (N_3578,N_1836,N_2037);
and U3579 (N_3579,N_3101,N_3405);
or U3580 (N_3580,In_4910,N_2311);
or U3581 (N_3581,N_3303,N_2435);
nand U3582 (N_3582,N_3357,N_3399);
xor U3583 (N_3583,N_2808,N_3034);
or U3584 (N_3584,N_3036,N_3076);
and U3585 (N_3585,N_2179,N_1326);
nor U3586 (N_3586,N_2820,In_1059);
and U3587 (N_3587,In_3224,N_2156);
and U3588 (N_3588,N_2395,N_970);
xor U3589 (N_3589,N_1991,N_2910);
and U3590 (N_3590,In_4325,N_1471);
nand U3591 (N_3591,In_1689,In_1709);
nand U3592 (N_3592,In_2944,N_1842);
nor U3593 (N_3593,N_2040,N_3086);
xnor U3594 (N_3594,N_823,N_3472);
xnor U3595 (N_3595,N_2625,N_3478);
or U3596 (N_3596,N_3242,N_2617);
or U3597 (N_3597,In_4208,N_3262);
nor U3598 (N_3598,N_2146,N_3077);
nand U3599 (N_3599,N_1857,In_415);
xnor U3600 (N_3600,N_3053,In_1849);
nor U3601 (N_3601,N_3174,N_2487);
xnor U3602 (N_3602,N_2055,N_2630);
or U3603 (N_3603,In_1153,N_3197);
nand U3604 (N_3604,N_2980,In_373);
or U3605 (N_3605,In_1356,N_2554);
or U3606 (N_3606,N_3106,N_3333);
xor U3607 (N_3607,In_2568,In_2496);
nand U3608 (N_3608,N_2752,N_2144);
nor U3609 (N_3609,N_2084,N_2021);
or U3610 (N_3610,In_2838,In_4060);
and U3611 (N_3611,In_2876,N_3277);
or U3612 (N_3612,N_2950,N_2853);
and U3613 (N_3613,In_1857,N_2325);
or U3614 (N_3614,N_2691,In_3362);
xor U3615 (N_3615,N_3271,In_4309);
and U3616 (N_3616,In_3732,N_3159);
xnor U3617 (N_3617,In_4059,N_1264);
xnor U3618 (N_3618,N_2409,N_220);
nand U3619 (N_3619,In_2172,In_2503);
nand U3620 (N_3620,N_2392,N_1658);
or U3621 (N_3621,N_807,N_3384);
nand U3622 (N_3622,N_1195,N_3375);
or U3623 (N_3623,N_2324,N_1559);
nor U3624 (N_3624,N_3090,In_600);
or U3625 (N_3625,N_3323,In_4242);
and U3626 (N_3626,N_3042,N_3358);
nor U3627 (N_3627,In_4,N_2740);
or U3628 (N_3628,N_3155,In_171);
or U3629 (N_3629,N_2860,N_3008);
nor U3630 (N_3630,N_3103,N_1825);
and U3631 (N_3631,N_2681,N_2963);
nor U3632 (N_3632,In_4255,N_2867);
nand U3633 (N_3633,N_1604,N_2095);
xor U3634 (N_3634,N_1967,N_3438);
and U3635 (N_3635,N_1834,N_2046);
and U3636 (N_3636,N_3024,N_3304);
and U3637 (N_3637,N_1651,N_1714);
xor U3638 (N_3638,N_1086,N_2505);
nand U3639 (N_3639,N_717,N_571);
xor U3640 (N_3640,N_3466,In_1382);
or U3641 (N_3641,N_3194,N_2177);
or U3642 (N_3642,N_2992,N_3260);
or U3643 (N_3643,N_3388,N_3154);
and U3644 (N_3644,N_3439,N_289);
or U3645 (N_3645,N_3286,N_3456);
xor U3646 (N_3646,In_3260,N_2603);
or U3647 (N_3647,N_1783,N_3473);
and U3648 (N_3648,N_249,N_2930);
nand U3649 (N_3649,In_1615,N_3185);
nor U3650 (N_3650,N_2697,N_2525);
and U3651 (N_3651,In_3863,N_162);
nor U3652 (N_3652,N_3060,In_565);
or U3653 (N_3653,In_3123,N_3343);
or U3654 (N_3654,In_3488,In_2836);
nor U3655 (N_3655,N_2655,N_3443);
nor U3656 (N_3656,In_35,N_2878);
and U3657 (N_3657,N_2815,In_3281);
or U3658 (N_3658,N_1720,In_1086);
nand U3659 (N_3659,In_4438,In_3735);
nand U3660 (N_3660,N_3339,N_3481);
nor U3661 (N_3661,In_1528,N_3288);
or U3662 (N_3662,In_2186,N_3129);
and U3663 (N_3663,In_2293,In_3141);
xor U3664 (N_3664,N_1261,In_4495);
and U3665 (N_3665,N_1989,In_896);
nor U3666 (N_3666,N_1669,In_4550);
nand U3667 (N_3667,N_144,N_444);
nand U3668 (N_3668,In_869,N_3347);
nor U3669 (N_3669,N_265,N_1008);
and U3670 (N_3670,N_3298,N_3442);
nand U3671 (N_3671,N_676,N_3165);
nand U3672 (N_3672,In_888,N_2900);
xor U3673 (N_3673,N_3132,In_3630);
or U3674 (N_3674,N_519,N_1080);
or U3675 (N_3675,N_3295,In_4866);
xnor U3676 (N_3676,N_3361,N_2587);
xor U3677 (N_3677,N_1180,N_2460);
nand U3678 (N_3678,N_2235,N_2086);
xnor U3679 (N_3679,N_3023,N_2643);
or U3680 (N_3680,In_3313,In_2893);
nand U3681 (N_3681,N_2590,N_2228);
or U3682 (N_3682,N_2503,N_3314);
or U3683 (N_3683,In_2413,N_3067);
nand U3684 (N_3684,N_3226,N_2947);
and U3685 (N_3685,N_3432,N_2835);
and U3686 (N_3686,N_1602,In_1450);
nand U3687 (N_3687,In_3773,N_2907);
or U3688 (N_3688,N_442,N_2157);
and U3689 (N_3689,N_3315,In_542);
nand U3690 (N_3690,N_3352,N_2417);
and U3691 (N_3691,N_2605,N_196);
xor U3692 (N_3692,N_3369,N_2618);
and U3693 (N_3693,In_1941,N_2945);
nor U3694 (N_3694,In_4633,N_2970);
or U3695 (N_3695,N_2626,In_182);
nor U3696 (N_3696,N_983,In_4353);
nand U3697 (N_3697,N_2551,N_2561);
nor U3698 (N_3698,N_3257,In_3742);
and U3699 (N_3699,N_2812,N_2966);
or U3700 (N_3700,N_2064,N_2621);
nand U3701 (N_3701,N_3205,In_4080);
nor U3702 (N_3702,N_2660,N_3348);
nand U3703 (N_3703,N_3411,In_4204);
nand U3704 (N_3704,In_3912,In_4624);
nand U3705 (N_3705,N_2199,In_1349);
or U3706 (N_3706,In_799,N_2931);
xor U3707 (N_3707,N_1565,N_1291);
or U3708 (N_3708,N_3273,In_4914);
or U3709 (N_3709,In_3739,N_2798);
nor U3710 (N_3710,N_3128,N_3278);
and U3711 (N_3711,In_4907,N_3113);
and U3712 (N_3712,In_3011,N_3497);
nand U3713 (N_3713,In_2165,N_3428);
nand U3714 (N_3714,N_1446,In_4324);
nor U3715 (N_3715,N_2784,N_3470);
xnor U3716 (N_3716,N_2645,N_3446);
nor U3717 (N_3717,N_3062,N_3102);
xnor U3718 (N_3718,N_3448,N_1950);
nand U3719 (N_3719,In_3805,N_931);
or U3720 (N_3720,N_1567,N_3021);
nand U3721 (N_3721,In_87,In_3813);
and U3722 (N_3722,N_2756,N_2388);
nor U3723 (N_3723,In_2027,N_2760);
xnor U3724 (N_3724,N_204,N_2953);
and U3725 (N_3725,N_3302,N_448);
and U3726 (N_3726,N_3447,N_3014);
nor U3727 (N_3727,N_2834,In_3927);
xor U3728 (N_3728,N_1678,N_1805);
nand U3729 (N_3729,N_3284,N_3012);
or U3730 (N_3730,N_3403,N_3108);
or U3731 (N_3731,N_1479,In_2894);
xnor U3732 (N_3732,N_576,N_3151);
nor U3733 (N_3733,N_322,N_841);
xor U3734 (N_3734,N_3394,N_3122);
nand U3735 (N_3735,In_4191,N_2929);
nor U3736 (N_3736,N_707,N_3356);
xor U3737 (N_3737,In_98,In_2936);
and U3738 (N_3738,N_1769,N_3396);
nand U3739 (N_3739,N_3425,N_3479);
nor U3740 (N_3740,N_2309,N_1563);
xor U3741 (N_3741,N_2672,In_3800);
xor U3742 (N_3742,In_3587,N_2872);
xnor U3743 (N_3743,N_3480,N_3248);
nand U3744 (N_3744,N_2851,N_3027);
nor U3745 (N_3745,N_1675,N_3422);
nor U3746 (N_3746,N_2999,N_3325);
nand U3747 (N_3747,N_2451,N_2778);
nor U3748 (N_3748,N_2670,N_2762);
nor U3749 (N_3749,N_3379,In_4716);
nor U3750 (N_3750,In_2809,N_3556);
and U3751 (N_3751,N_3735,N_3087);
and U3752 (N_3752,N_3727,N_2871);
nand U3753 (N_3753,N_2732,N_3145);
and U3754 (N_3754,N_3157,N_3734);
and U3755 (N_3755,N_2642,In_1994);
xnor U3756 (N_3756,N_3071,N_2527);
or U3757 (N_3757,N_3686,N_3287);
nand U3758 (N_3758,N_2277,N_3454);
or U3759 (N_3759,N_2148,In_1417);
nand U3760 (N_3760,In_846,N_3605);
or U3761 (N_3761,N_33,N_2680);
and U3762 (N_3762,N_2012,N_1971);
nand U3763 (N_3763,N_2375,N_2062);
nor U3764 (N_3764,In_762,In_2704);
nor U3765 (N_3765,N_3545,In_1816);
and U3766 (N_3766,N_1662,N_3429);
xnor U3767 (N_3767,N_3093,N_2793);
or U3768 (N_3768,N_2673,N_3048);
nor U3769 (N_3769,N_3567,N_1623);
and U3770 (N_3770,N_2741,N_1067);
nor U3771 (N_3771,N_1970,N_2297);
nor U3772 (N_3772,N_1432,In_4081);
nor U3773 (N_3773,In_3480,In_4517);
and U3774 (N_3774,N_3533,N_1938);
and U3775 (N_3775,N_1485,N_2866);
xnor U3776 (N_3776,N_3660,In_1407);
xnor U3777 (N_3777,N_3704,In_1408);
xnor U3778 (N_3778,N_2606,N_2881);
and U3779 (N_3779,N_2526,In_3679);
nand U3780 (N_3780,N_2991,N_3430);
xor U3781 (N_3781,N_1838,N_1680);
nor U3782 (N_3782,N_3083,In_4842);
nand U3783 (N_3783,N_2748,N_3223);
nor U3784 (N_3784,N_3218,N_415);
and U3785 (N_3785,N_2051,In_3164);
nor U3786 (N_3786,N_3114,N_3699);
nor U3787 (N_3787,In_4791,In_4535);
xnor U3788 (N_3788,N_3120,N_3500);
or U3789 (N_3789,N_3505,N_3019);
xor U3790 (N_3790,N_2372,N_3161);
and U3791 (N_3791,N_3562,N_2986);
or U3792 (N_3792,N_2609,N_968);
nor U3793 (N_3793,N_3007,N_3091);
nor U3794 (N_3794,In_4878,N_736);
or U3795 (N_3795,In_817,N_834);
nand U3796 (N_3796,N_2589,N_400);
xor U3797 (N_3797,N_3230,N_3282);
nor U3798 (N_3798,In_333,N_3520);
nor U3799 (N_3799,N_3376,In_3226);
nand U3800 (N_3800,N_715,N_3078);
xnor U3801 (N_3801,In_1322,In_1787);
or U3802 (N_3802,N_3652,N_2747);
nand U3803 (N_3803,N_897,N_3544);
nor U3804 (N_3804,N_1660,N_3198);
nor U3805 (N_3805,N_3738,N_665);
and U3806 (N_3806,N_3691,N_3418);
nor U3807 (N_3807,In_2519,N_29);
nor U3808 (N_3808,N_775,N_3730);
xnor U3809 (N_3809,N_3427,N_652);
nor U3810 (N_3810,N_3661,N_3213);
nand U3811 (N_3811,N_3664,N_3044);
and U3812 (N_3812,In_1905,N_2774);
or U3813 (N_3813,N_3535,N_3651);
nor U3814 (N_3814,N_1039,N_3569);
nor U3815 (N_3815,N_74,N_1633);
or U3816 (N_3816,N_3319,N_2775);
xnor U3817 (N_3817,N_3521,N_1705);
xnor U3818 (N_3818,N_2888,N_2832);
or U3819 (N_3819,N_687,N_2515);
nor U3820 (N_3820,N_3004,N_3671);
nor U3821 (N_3821,N_3612,N_3269);
or U3822 (N_3822,N_1999,N_2425);
nor U3823 (N_3823,N_3370,N_3701);
xor U3824 (N_3824,N_3622,In_3809);
and U3825 (N_3825,N_3696,N_2588);
nor U3826 (N_3826,N_3641,In_2234);
or U3827 (N_3827,N_2464,N_996);
nor U3828 (N_3828,N_1811,In_3865);
nor U3829 (N_3829,N_2917,N_2514);
nor U3830 (N_3830,N_2557,N_2739);
and U3831 (N_3831,N_639,N_3437);
xnor U3832 (N_3832,N_866,In_262);
and U3833 (N_3833,N_712,N_1460);
nor U3834 (N_3834,N_2390,N_3387);
nor U3835 (N_3835,N_3195,In_2949);
nand U3836 (N_3836,N_3713,N_2941);
and U3837 (N_3837,In_737,In_3621);
nor U3838 (N_3838,N_3337,N_3634);
or U3839 (N_3839,N_3390,N_2810);
nand U3840 (N_3840,N_971,N_3345);
and U3841 (N_3841,N_3240,N_2961);
nand U3842 (N_3842,N_2884,N_2813);
nand U3843 (N_3843,N_2807,N_3225);
xnor U3844 (N_3844,N_3710,N_2915);
nand U3845 (N_3845,In_145,N_3137);
nand U3846 (N_3846,N_1978,In_3530);
nor U3847 (N_3847,N_20,N_3619);
nor U3848 (N_3848,N_3111,In_2162);
and U3849 (N_3849,N_3698,In_4717);
or U3850 (N_3850,In_4382,N_3450);
xnor U3851 (N_3851,N_2358,N_2213);
nor U3852 (N_3852,N_3434,N_3061);
or U3853 (N_3853,N_3717,N_2007);
nand U3854 (N_3854,N_3732,N_1436);
or U3855 (N_3855,In_142,In_369);
xor U3856 (N_3856,In_3855,N_3618);
nand U3857 (N_3857,N_2422,N_2901);
and U3858 (N_3858,N_3175,N_3018);
nor U3859 (N_3859,N_3724,N_1318);
nand U3860 (N_3860,N_746,N_3040);
nand U3861 (N_3861,In_3120,N_2753);
nand U3862 (N_3862,N_150,N_3057);
nand U3863 (N_3863,In_2253,In_3075);
or U3864 (N_3864,N_3117,N_2924);
xor U3865 (N_3865,N_3307,N_3502);
and U3866 (N_3866,N_2806,N_3662);
xnor U3867 (N_3867,N_3261,N_3329);
and U3868 (N_3868,N_2856,N_734);
or U3869 (N_3869,N_3451,N_3338);
or U3870 (N_3870,N_3621,N_3504);
nand U3871 (N_3871,N_1161,N_3552);
and U3872 (N_3872,N_3121,In_1961);
nand U3873 (N_3873,N_2345,N_2887);
xor U3874 (N_3874,In_3784,N_2453);
xnor U3875 (N_3875,N_2766,In_4588);
and U3876 (N_3876,N_1666,N_3715);
nor U3877 (N_3877,N_3714,In_3068);
xnor U3878 (N_3878,N_3299,N_1192);
nand U3879 (N_3879,In_1101,N_915);
nor U3880 (N_3880,N_3528,In_1411);
or U3881 (N_3881,N_3049,In_4380);
xnor U3882 (N_3882,In_695,N_2131);
or U3883 (N_3883,N_2426,N_2821);
nand U3884 (N_3884,In_4186,N_3326);
nor U3885 (N_3885,N_3516,N_2355);
xor U3886 (N_3886,N_2988,N_3359);
xor U3887 (N_3887,In_4256,N_1376);
nor U3888 (N_3888,N_3742,N_2472);
and U3889 (N_3889,N_1784,N_3311);
xor U3890 (N_3890,N_1983,N_3283);
nand U3891 (N_3891,N_3032,N_3587);
and U3892 (N_3892,In_4476,N_2906);
nor U3893 (N_3893,In_2328,N_932);
nor U3894 (N_3894,N_2803,N_3702);
and U3895 (N_3895,N_3158,In_2747);
and U3896 (N_3896,N_3728,N_3690);
xnor U3897 (N_3897,N_2244,In_3074);
xnor U3898 (N_3898,N_3708,N_3558);
or U3899 (N_3899,N_3578,In_2721);
or U3900 (N_3900,In_910,N_299);
or U3901 (N_3901,N_3474,N_3201);
nor U3902 (N_3902,N_3033,N_2652);
xor U3903 (N_3903,N_3170,N_3571);
or U3904 (N_3904,N_205,N_3586);
xor U3905 (N_3905,N_2407,N_2002);
nand U3906 (N_3906,N_3721,N_1973);
nand U3907 (N_3907,N_1581,N_3492);
nand U3908 (N_3908,N_1236,N_3332);
nor U3909 (N_3909,N_3527,In_4519);
nand U3910 (N_3910,In_3263,N_3577);
xnor U3911 (N_3911,N_3608,N_3126);
nand U3912 (N_3912,N_3256,N_2581);
and U3913 (N_3913,N_2846,N_3436);
nand U3914 (N_3914,N_2864,N_3031);
nand U3915 (N_3915,N_2240,N_2566);
or U3916 (N_3916,N_3553,In_4799);
or U3917 (N_3917,N_2800,N_1903);
nor U3918 (N_3918,N_2921,N_3002);
and U3919 (N_3919,In_3270,N_1069);
nand U3920 (N_3920,N_2091,N_3016);
xor U3921 (N_3921,N_3344,N_3607);
nand U3922 (N_3922,N_3417,N_2981);
nor U3923 (N_3923,N_3255,N_3340);
nand U3924 (N_3924,N_2301,N_3322);
or U3925 (N_3925,N_3679,N_3581);
and U3926 (N_3926,N_2378,N_3615);
nor U3927 (N_3927,In_4896,N_3613);
and U3928 (N_3928,N_458,N_3720);
nand U3929 (N_3929,N_3596,N_1259);
nor U3930 (N_3930,N_2990,N_3693);
nand U3931 (N_3931,N_3650,In_185);
xor U3932 (N_3932,In_3767,N_3677);
and U3933 (N_3933,N_3309,In_863);
xnor U3934 (N_3934,N_1909,N_2919);
or U3935 (N_3935,N_3591,N_2895);
nor U3936 (N_3936,In_287,N_3483);
and U3937 (N_3937,N_882,In_847);
nor U3938 (N_3938,In_4746,N_3280);
nand U3939 (N_3939,In_1155,In_2796);
nor U3940 (N_3940,N_2746,N_3477);
nand U3941 (N_3941,N_3665,N_3471);
nor U3942 (N_3942,In_249,N_3172);
and U3943 (N_3943,N_3593,N_452);
nor U3944 (N_3944,N_3186,N_3657);
or U3945 (N_3945,N_2290,In_355);
nand U3946 (N_3946,N_2524,N_3669);
or U3947 (N_3947,N_2839,N_2744);
nor U3948 (N_3948,N_2736,In_1184);
and U3949 (N_3949,N_2134,N_3104);
nor U3950 (N_3950,N_771,N_3731);
or U3951 (N_3951,N_1169,N_2114);
nor U3952 (N_3952,N_3496,In_4974);
and U3953 (N_3953,In_2770,N_2758);
nand U3954 (N_3954,In_1250,N_3580);
and U3955 (N_3955,N_2781,N_2089);
and U3956 (N_3956,N_334,N_3270);
nor U3957 (N_3957,N_3163,N_1674);
and U3958 (N_3958,N_3606,In_2576);
or U3959 (N_3959,N_3037,In_1964);
nand U3960 (N_3960,N_3244,N_2488);
nor U3961 (N_3961,In_4419,N_2636);
nand U3962 (N_3962,In_4195,In_2501);
xnor U3963 (N_3963,N_30,N_3566);
nor U3964 (N_3964,N_3635,N_1741);
or U3965 (N_3965,N_765,In_4241);
or U3966 (N_3966,N_3096,N_2797);
nor U3967 (N_3967,In_3182,In_3319);
nor U3968 (N_3968,N_2682,N_3743);
nand U3969 (N_3969,N_3020,N_3610);
nor U3970 (N_3970,In_4930,N_3415);
nor U3971 (N_3971,N_3611,N_3296);
xor U3972 (N_3972,N_1420,N_853);
nand U3973 (N_3973,N_2973,N_3457);
and U3974 (N_3974,N_3475,In_1453);
nand U3975 (N_3975,N_3131,N_459);
or U3976 (N_3976,N_2613,In_2199);
nor U3977 (N_3977,N_2825,N_3334);
nand U3978 (N_3978,N_1688,N_1309);
xnor U3979 (N_3979,In_4027,N_3563);
xnor U3980 (N_3980,N_3292,N_3331);
nand U3981 (N_3981,N_3565,In_3115);
xnor U3982 (N_3982,N_3510,N_3085);
and U3983 (N_3983,N_3393,N_1461);
nand U3984 (N_3984,N_2272,N_3507);
and U3985 (N_3985,In_4976,In_4211);
or U3986 (N_3986,In_3325,N_3579);
nor U3987 (N_3987,N_2954,N_3364);
xnor U3988 (N_3988,N_3543,In_2902);
nand U3989 (N_3989,N_2097,N_2767);
nand U3990 (N_3990,In_4381,N_2706);
nor U3991 (N_3991,N_3354,N_2905);
and U3992 (N_3992,N_3636,N_3274);
or U3993 (N_3993,N_3055,N_2532);
xnor U3994 (N_3994,N_3604,N_3092);
nor U3995 (N_3995,N_3599,In_3005);
or U3996 (N_3996,In_4568,N_3200);
nand U3997 (N_3997,In_203,N_1539);
and U3998 (N_3998,N_1992,N_147);
nand U3999 (N_3999,In_4759,N_3377);
nand U4000 (N_4000,N_3750,N_3005);
nor U4001 (N_4001,N_3398,N_3933);
xnor U4002 (N_4002,N_3421,N_3508);
nand U4003 (N_4003,N_3962,In_178);
xnor U4004 (N_4004,In_3748,N_3957);
or U4005 (N_4005,N_3227,N_3977);
and U4006 (N_4006,N_1462,N_3190);
nand U4007 (N_4007,In_2773,In_3796);
and U4008 (N_4008,N_2828,N_580);
or U4009 (N_4009,N_2742,N_3765);
xnor U4010 (N_4010,N_3925,N_3648);
and U4011 (N_4011,N_3630,N_3683);
nand U4012 (N_4012,N_3847,N_2649);
or U4013 (N_4013,N_3740,In_4886);
nor U4014 (N_4014,N_1504,In_4287);
nand U4015 (N_4015,N_3392,N_3167);
nand U4016 (N_4016,N_3320,N_3776);
xor U4017 (N_4017,In_1405,N_1656);
nor U4018 (N_4018,N_1103,N_3998);
and U4019 (N_4019,N_3755,N_3841);
and U4020 (N_4020,N_1379,In_1806);
and U4021 (N_4021,N_3638,In_2588);
xor U4022 (N_4022,N_3413,N_3883);
or U4023 (N_4023,N_3959,N_3547);
nor U4024 (N_4024,N_3753,N_3324);
or U4025 (N_4025,In_4922,N_2843);
xnor U4026 (N_4026,N_3188,N_3892);
and U4027 (N_4027,In_2847,N_2243);
or U4028 (N_4028,N_3842,N_978);
and U4029 (N_4029,N_3263,N_3749);
nor U4030 (N_4030,N_3729,N_1850);
xor U4031 (N_4031,N_3815,N_3990);
nand U4032 (N_4032,N_3764,N_3893);
xor U4033 (N_4033,N_3938,N_3433);
nand U4034 (N_4034,N_3381,N_3926);
or U4035 (N_4035,N_3467,N_2836);
nand U4036 (N_4036,N_3903,N_3380);
nor U4037 (N_4037,N_1540,In_64);
or U4038 (N_4038,N_2814,In_1773);
nor U4039 (N_4039,N_1276,N_3658);
xnor U4040 (N_4040,N_3453,N_2463);
and U4041 (N_4041,N_3169,N_3673);
or U4042 (N_4042,N_3906,N_3802);
nand U4043 (N_4043,In_4513,N_3251);
xnor U4044 (N_4044,N_3967,N_2540);
nor U4045 (N_4045,N_3064,N_2223);
nand U4046 (N_4046,N_3523,In_1247);
or U4047 (N_4047,In_907,N_3797);
or U4048 (N_4048,N_3530,N_1340);
xor U4049 (N_4049,N_3902,N_3546);
and U4050 (N_4050,N_3589,N_574);
xor U4051 (N_4051,N_2075,In_758);
nand U4052 (N_4052,N_3285,In_3142);
or U4053 (N_4053,N_3617,N_3886);
xor U4054 (N_4054,N_3923,In_2314);
nor U4055 (N_4055,N_961,N_3829);
nand U4056 (N_4056,N_2025,N_3639);
and U4057 (N_4057,In_2784,N_3767);
nor U4058 (N_4058,N_540,N_2707);
xor U4059 (N_4059,N_3300,N_1573);
xor U4060 (N_4060,In_767,N_3575);
and U4061 (N_4061,N_3668,N_3495);
or U4062 (N_4062,N_3625,N_2942);
and U4063 (N_4063,In_4473,N_3873);
nor U4064 (N_4064,N_3772,N_3407);
nor U4065 (N_4065,N_2982,N_3947);
nor U4066 (N_4066,N_3647,N_1698);
and U4067 (N_4067,N_3921,In_406);
and U4068 (N_4068,N_3588,N_3011);
nand U4069 (N_4069,N_1168,N_2359);
nor U4070 (N_4070,N_3537,N_3025);
or U4071 (N_4071,N_3557,N_3199);
nor U4072 (N_4072,N_1729,N_3733);
nor U4073 (N_4073,N_2880,N_2936);
nand U4074 (N_4074,N_3963,N_2668);
xor U4075 (N_4075,N_3901,N_3723);
or U4076 (N_4076,N_3089,N_3640);
or U4077 (N_4077,N_3951,N_3790);
xnor U4078 (N_4078,N_3209,N_2026);
and U4079 (N_4079,N_3862,In_4396);
or U4080 (N_4080,In_4843,N_2602);
or U4081 (N_4081,N_3424,N_443);
and U4082 (N_4082,N_3268,N_3318);
and U4083 (N_4083,N_3768,In_3355);
nor U4084 (N_4084,N_1630,In_1182);
nand U4085 (N_4085,In_3083,N_3482);
nand U4086 (N_4086,N_3924,N_2845);
and U4087 (N_4087,N_3834,N_2578);
or U4088 (N_4088,N_1798,In_2642);
nor U4089 (N_4089,N_3914,In_2400);
nor U4090 (N_4090,N_3837,N_2017);
nor U4091 (N_4091,N_3939,N_2601);
xor U4092 (N_4092,N_3609,N_3856);
nor U4093 (N_4093,N_3984,N_3695);
nand U4094 (N_4094,N_1800,In_1927);
nand U4095 (N_4095,N_3789,In_691);
nor U4096 (N_4096,N_2500,N_2060);
and U4097 (N_4097,N_3468,N_3030);
xor U4098 (N_4098,N_3513,In_4744);
or U4099 (N_4099,N_2438,In_201);
or U4100 (N_4100,N_2475,N_86);
nand U4101 (N_4101,N_2523,N_3801);
or U4102 (N_4102,In_672,N_3759);
or U4103 (N_4103,N_3852,N_3784);
nor U4104 (N_4104,N_3857,N_2690);
nor U4105 (N_4105,N_3400,N_2187);
nand U4106 (N_4106,N_3602,N_539);
nand U4107 (N_4107,N_2819,N_2217);
nand U4108 (N_4108,In_2137,N_3888);
nand U4109 (N_4109,N_3395,N_3850);
and U4110 (N_4110,N_3164,N_3631);
nand U4111 (N_4111,In_2173,N_2056);
or U4112 (N_4112,N_3568,N_3908);
xnor U4113 (N_4113,N_3839,N_3777);
nor U4114 (N_4114,N_3798,N_1937);
or U4115 (N_4115,N_3851,N_2987);
nand U4116 (N_4116,N_1430,In_147);
or U4117 (N_4117,N_3147,N_3182);
nand U4118 (N_4118,N_3816,N_3469);
nor U4119 (N_4119,N_2493,In_2376);
and U4120 (N_4120,N_2996,N_3684);
or U4121 (N_4121,N_1764,In_2175);
xor U4122 (N_4122,N_3330,N_738);
nor U4123 (N_4123,N_3682,N_2789);
nand U4124 (N_4124,N_399,N_3741);
nor U4125 (N_4125,N_810,N_3368);
nand U4126 (N_4126,In_4345,N_3920);
nor U4127 (N_4127,In_2729,N_3402);
and U4128 (N_4128,N_692,In_862);
and U4129 (N_4129,N_2934,In_4323);
or U4130 (N_4130,N_3573,In_2380);
nor U4131 (N_4131,In_3666,N_3133);
and U4132 (N_4132,N_3670,In_1266);
and U4133 (N_4133,N_2896,N_3493);
or U4134 (N_4134,N_1899,N_3105);
nand U4135 (N_4135,N_542,N_2595);
and U4136 (N_4136,N_3041,N_3614);
nor U4137 (N_4137,N_2198,N_2160);
nor U4138 (N_4138,N_3846,N_3751);
nor U4139 (N_4139,N_2281,N_3672);
xor U4140 (N_4140,In_93,N_1643);
nor U4141 (N_4141,N_2073,N_3522);
or U4142 (N_4142,N_3880,N_3559);
nand U4143 (N_4143,N_3879,N_1787);
or U4144 (N_4144,N_3006,In_2458);
or U4145 (N_4145,In_1641,N_3488);
nand U4146 (N_4146,N_3810,N_2869);
and U4147 (N_4147,N_3866,N_1262);
nand U4148 (N_4148,N_3928,N_3222);
and U4149 (N_4149,N_2622,In_2707);
nand U4150 (N_4150,N_3890,N_2255);
xnor U4151 (N_4151,N_3995,N_2122);
and U4152 (N_4152,In_595,In_1330);
xnor U4153 (N_4153,N_3595,In_794);
nand U4154 (N_4154,N_3806,N_2336);
xnor U4155 (N_4155,N_3812,N_3308);
nand U4156 (N_4156,N_3961,N_3646);
nor U4157 (N_4157,In_4009,N_3594);
nand U4158 (N_4158,N_1590,N_3899);
nand U4159 (N_4159,N_3485,N_3366);
nand U4160 (N_4160,N_3628,In_3691);
or U4161 (N_4161,N_2399,N_3799);
or U4162 (N_4162,N_2408,N_1668);
xnor U4163 (N_4163,N_1177,N_3827);
xnor U4164 (N_4164,N_2912,N_3626);
nor U4165 (N_4165,N_1635,N_3118);
xor U4166 (N_4166,N_3813,N_3922);
and U4167 (N_4167,N_3511,N_421);
or U4168 (N_4168,N_3868,N_1707);
xnor U4169 (N_4169,N_3988,In_3947);
and U4170 (N_4170,N_2795,N_1263);
nor U4171 (N_4171,In_833,N_1808);
xor U4172 (N_4172,N_3688,N_3904);
nor U4173 (N_4173,N_2312,N_2614);
nand U4174 (N_4174,N_2333,N_2068);
nor U4175 (N_4175,N_3853,N_3531);
nand U4176 (N_4176,N_3718,N_3778);
xnor U4177 (N_4177,In_3335,In_3528);
nor U4178 (N_4178,N_3712,N_3135);
or U4179 (N_4179,N_1552,N_3719);
and U4180 (N_4180,N_491,In_2631);
xnor U4181 (N_4181,N_3281,N_3459);
nor U4182 (N_4182,In_2262,N_2396);
nand U4183 (N_4183,N_2411,N_3709);
nand U4184 (N_4184,N_3795,N_3667);
nand U4185 (N_4185,N_3966,N_3532);
nor U4186 (N_4186,N_3942,N_1213);
or U4187 (N_4187,N_3907,N_2568);
or U4188 (N_4188,N_3463,In_1978);
nor U4189 (N_4189,In_1765,N_2448);
or U4190 (N_4190,In_1700,N_3216);
or U4191 (N_4191,N_3675,N_3070);
nand U4192 (N_4192,N_3506,N_2271);
nand U4193 (N_4193,N_3541,N_3142);
nor U4194 (N_4194,N_3409,N_3736);
xnor U4195 (N_4195,N_2879,In_24);
or U4196 (N_4196,In_1661,N_3518);
xor U4197 (N_4197,N_3440,N_3805);
xor U4198 (N_4198,N_3221,N_2944);
nand U4199 (N_4199,N_2374,N_3494);
nand U4200 (N_4200,N_3360,In_3550);
xor U4201 (N_4201,N_1545,N_3993);
and U4202 (N_4202,N_3054,N_2914);
nor U4203 (N_4203,N_3585,N_3824);
nor U4204 (N_4204,N_3773,N_3335);
xnor U4205 (N_4205,In_4390,N_3830);
or U4206 (N_4206,In_3617,N_3756);
nand U4207 (N_4207,N_3946,N_3919);
and U4208 (N_4208,N_3989,N_3911);
and U4209 (N_4209,In_3442,N_3844);
and U4210 (N_4210,N_3814,N_1689);
nor U4211 (N_4211,N_3252,N_3891);
or U4212 (N_4212,N_1868,N_85);
and U4213 (N_4213,N_3781,N_3327);
nand U4214 (N_4214,In_1516,N_3317);
and U4215 (N_4215,N_3321,N_3279);
nor U4216 (N_4216,N_3916,N_2757);
and U4217 (N_4217,N_1951,N_3800);
nor U4218 (N_4218,N_3143,N_1597);
nor U4219 (N_4219,N_865,N_3098);
xor U4220 (N_4220,In_2952,N_3970);
nor U4221 (N_4221,N_3978,N_3796);
nor U4222 (N_4222,N_3431,In_3905);
xnor U4223 (N_4223,N_1725,N_3774);
nand U4224 (N_4224,N_2335,N_3350);
and U4225 (N_4225,In_923,N_2397);
and U4226 (N_4226,N_3794,N_3603);
and U4227 (N_4227,N_3896,N_3992);
and U4228 (N_4228,N_2544,N_3780);
xnor U4229 (N_4229,In_4657,N_3976);
nor U4230 (N_4230,In_4268,In_2255);
and U4231 (N_4231,N_3782,N_2577);
and U4232 (N_4232,N_2329,N_3788);
xor U4233 (N_4233,N_2053,N_3766);
xor U4234 (N_4234,N_2210,N_1580);
and U4235 (N_4235,N_3189,N_2654);
xnor U4236 (N_4236,N_3499,N_3754);
nor U4237 (N_4237,N_3968,N_2459);
xor U4238 (N_4238,N_3574,N_3600);
xnor U4239 (N_4239,N_2087,In_735);
nor U4240 (N_4240,N_3725,N_3975);
and U4241 (N_4241,N_3207,N_3116);
or U4242 (N_4242,N_3854,N_3771);
or U4243 (N_4243,In_632,N_1117);
and U4244 (N_4244,N_3519,N_3624);
and U4245 (N_4245,N_3775,In_3348);
or U4246 (N_4246,N_368,N_3786);
xor U4247 (N_4247,N_1657,N_3386);
nor U4248 (N_4248,N_244,N_1939);
nor U4249 (N_4249,N_3633,In_4862);
xnor U4250 (N_4250,N_4140,N_48);
or U4251 (N_4251,N_2721,N_4224);
or U4252 (N_4252,N_2913,N_1507);
and U4253 (N_4253,N_2558,N_4197);
nand U4254 (N_4254,N_4166,N_1522);
xor U4255 (N_4255,N_3597,N_1877);
and U4256 (N_4256,N_4061,N_3785);
nor U4257 (N_4257,N_4101,N_4204);
nand U4258 (N_4258,N_4200,N_4133);
nand U4259 (N_4259,N_2678,N_3341);
nand U4260 (N_4260,N_3791,N_3666);
nand U4261 (N_4261,N_4115,N_3927);
and U4262 (N_4262,N_1203,In_4092);
and U4263 (N_4263,N_3328,N_4167);
and U4264 (N_4264,N_4036,N_3503);
and U4265 (N_4265,N_2809,N_3803);
and U4266 (N_4266,N_4218,N_2926);
nand U4267 (N_4267,N_1258,N_3997);
nand U4268 (N_4268,N_4249,N_4117);
xnor U4269 (N_4269,N_3974,In_1306);
nor U4270 (N_4270,N_4160,N_4170);
nand U4271 (N_4271,In_2135,N_3910);
xor U4272 (N_4272,N_4236,N_3509);
and U4273 (N_4273,N_3253,N_3832);
xnor U4274 (N_4274,N_3912,N_3900);
or U4275 (N_4275,N_4155,N_3845);
nand U4276 (N_4276,N_4222,N_126);
nand U4277 (N_4277,N_3752,N_1053);
nand U4278 (N_4278,N_4174,N_4048);
nor U4279 (N_4279,N_4079,N_3929);
and U4280 (N_4280,N_276,N_4137);
xor U4281 (N_4281,In_4254,N_3981);
nand U4282 (N_4282,N_995,N_3236);
nor U4283 (N_4283,In_2791,N_4087);
or U4284 (N_4284,N_3642,N_4196);
nor U4285 (N_4285,N_3865,N_4045);
and U4286 (N_4286,N_3964,N_3484);
and U4287 (N_4287,N_4211,N_4057);
nand U4288 (N_4288,N_3779,N_1917);
and U4289 (N_4289,N_3840,N_4114);
xor U4290 (N_4290,N_2457,N_3692);
xnor U4291 (N_4291,N_4156,N_4147);
or U4292 (N_4292,N_3539,N_3941);
or U4293 (N_4293,In_1493,N_3534);
or U4294 (N_4294,N_4026,N_3864);
or U4295 (N_4295,N_4084,In_1416);
nand U4296 (N_4296,N_3792,In_3302);
nand U4297 (N_4297,N_4182,N_3958);
nor U4298 (N_4298,N_3524,N_4128);
or U4299 (N_4299,N_4071,N_3654);
nor U4300 (N_4300,N_4245,N_4072);
nor U4301 (N_4301,N_4074,N_4131);
or U4302 (N_4302,N_1513,N_4073);
and U4303 (N_4303,In_181,N_4220);
xnor U4304 (N_4304,N_4232,N_3944);
xor U4305 (N_4305,N_4135,N_3123);
nand U4306 (N_4306,N_4190,N_3426);
nor U4307 (N_4307,In_934,N_4123);
nor U4308 (N_4308,N_4001,N_3885);
xor U4309 (N_4309,N_2729,In_1755);
or U4310 (N_4310,N_3859,N_3748);
nand U4311 (N_4311,N_4126,N_2788);
nand U4312 (N_4312,N_3835,N_3889);
nand U4313 (N_4313,N_4248,N_2079);
or U4314 (N_4314,N_4227,N_4215);
or U4315 (N_4315,N_3737,In_740);
nand U4316 (N_4316,In_699,N_3960);
nand U4317 (N_4317,N_4091,N_3538);
and U4318 (N_4318,N_2616,N_4025);
xnor U4319 (N_4319,N_3385,N_3464);
and U4320 (N_4320,N_3913,N_3312);
nor U4321 (N_4321,N_2700,N_1893);
nand U4322 (N_4322,N_2959,N_4125);
nor U4323 (N_4323,N_2675,In_94);
nor U4324 (N_4324,In_2136,N_4106);
nand U4325 (N_4325,N_4230,N_3408);
or U4326 (N_4326,N_4082,N_2817);
and U4327 (N_4327,N_3953,N_3564);
or U4328 (N_4328,N_4040,N_4134);
nor U4329 (N_4329,N_3965,N_2648);
nand U4330 (N_4330,In_4167,N_2978);
and U4331 (N_4331,N_4148,N_3412);
or U4332 (N_4332,N_2123,N_4104);
nand U4333 (N_4333,N_4152,N_3836);
and U4334 (N_4334,N_3445,N_4111);
xnor U4335 (N_4335,N_3996,N_4122);
or U4336 (N_4336,N_3526,N_3685);
or U4337 (N_4337,N_1351,N_2783);
nor U4338 (N_4338,N_1697,N_3029);
nor U4339 (N_4339,N_3056,N_3874);
xnor U4340 (N_4340,N_1969,N_107);
and U4341 (N_4341,N_4109,N_3987);
nand U4342 (N_4342,N_3110,In_2816);
nand U4343 (N_4343,N_4054,N_2474);
nor U4344 (N_4344,N_852,N_4011);
and U4345 (N_4345,N_3342,N_4193);
xnor U4346 (N_4346,N_4180,N_4005);
nor U4347 (N_4347,N_3219,N_3808);
nand U4348 (N_4348,N_4153,N_3536);
nand U4349 (N_4349,N_4059,N_4240);
or U4350 (N_4350,N_3700,In_805);
or U4351 (N_4351,N_4055,N_4143);
or U4352 (N_4352,N_4105,N_2882);
nor U4353 (N_4353,N_1321,N_3649);
nand U4354 (N_4354,N_3909,N_3744);
nand U4355 (N_4355,N_4103,N_3867);
xnor U4356 (N_4356,In_4313,N_3822);
and U4357 (N_4357,N_3570,N_4024);
xnor U4358 (N_4358,N_4235,In_1654);
xor U4359 (N_4359,N_4205,N_4183);
and U4360 (N_4360,N_3136,N_3038);
nor U4361 (N_4361,N_3548,N_4075);
and U4362 (N_4362,N_4163,N_3297);
nor U4363 (N_4363,N_3035,N_4029);
xnor U4364 (N_4364,N_1530,N_4186);
nor U4365 (N_4365,N_2855,N_3234);
nor U4366 (N_4366,N_863,N_3490);
nand U4367 (N_4367,N_4194,N_3404);
nand U4368 (N_4368,N_1653,N_3809);
nor U4369 (N_4369,N_3265,N_4238);
nor U4370 (N_4370,In_179,N_4002);
and U4371 (N_4371,N_3220,N_3525);
or U4372 (N_4372,N_2972,N_3572);
nor U4373 (N_4373,N_4157,N_4202);
xnor U4374 (N_4374,N_3821,N_3656);
nand U4375 (N_4375,N_3542,N_4208);
nand U4376 (N_4376,N_4107,N_3620);
nand U4377 (N_4377,N_4198,N_4199);
xor U4378 (N_4378,N_4201,N_4176);
nor U4379 (N_4379,N_3918,N_2607);
nor U4380 (N_4380,N_4165,N_325);
nand U4381 (N_4381,N_3629,N_4161);
xor U4382 (N_4382,N_3979,N_2711);
xor U4383 (N_4383,N_4228,N_4003);
nand U4384 (N_4384,N_4145,N_3306);
or U4385 (N_4385,N_3956,N_3074);
or U4386 (N_4386,N_4062,N_3378);
xor U4387 (N_4387,N_3659,N_4009);
nand U4388 (N_4388,N_4112,N_4162);
or U4389 (N_4389,N_3576,N_3875);
or U4390 (N_4390,N_3009,N_625);
xnor U4391 (N_4391,In_2982,N_3166);
and U4392 (N_4392,N_4234,N_3291);
nand U4393 (N_4393,N_620,N_3627);
nand U4394 (N_4394,N_4168,In_2377);
nand U4395 (N_4395,N_4006,N_3881);
nand U4396 (N_4396,N_3674,N_3985);
xor U4397 (N_4397,N_2034,N_3367);
nand U4398 (N_4398,N_2176,In_4159);
nand U4399 (N_4399,N_3371,N_4132);
and U4400 (N_4400,N_3760,In_2762);
xnor U4401 (N_4401,N_3355,N_3414);
and U4402 (N_4402,N_2754,N_4118);
and U4403 (N_4403,N_2928,N_2174);
xnor U4404 (N_4404,N_4090,In_2271);
or U4405 (N_4405,N_4213,N_3681);
nor U4406 (N_4406,N_2077,N_1019);
or U4407 (N_4407,N_4172,N_4022);
and U4408 (N_4408,In_940,N_4116);
xor U4409 (N_4409,In_4637,N_3818);
xor U4410 (N_4410,N_3301,N_3217);
xnor U4411 (N_4411,N_3894,N_3391);
and U4412 (N_4412,N_3264,N_2035);
xor U4413 (N_4413,N_2993,N_3872);
or U4414 (N_4414,In_2592,N_3943);
and U4415 (N_4415,N_1493,N_4093);
xor U4416 (N_4416,N_3178,N_3250);
nor U4417 (N_4417,N_4042,N_1793);
xnor U4418 (N_4418,N_3435,N_3876);
xnor U4419 (N_4419,N_2316,N_4179);
and U4420 (N_4420,N_3769,N_4181);
xor U4421 (N_4421,N_4219,N_3833);
nor U4422 (N_4422,N_209,N_4136);
xnor U4423 (N_4423,N_4092,N_4243);
nand U4424 (N_4424,N_3869,N_3884);
xnor U4425 (N_4425,N_3069,N_4019);
and U4426 (N_4426,N_4064,N_4207);
xnor U4427 (N_4427,In_299,N_4223);
xor U4428 (N_4428,N_4095,N_1634);
nor U4429 (N_4429,In_2741,N_1094);
or U4430 (N_4430,N_3758,N_3346);
nand U4431 (N_4431,N_2357,N_4108);
xor U4432 (N_4432,N_3419,N_4159);
nand U4433 (N_4433,N_4016,N_3930);
or U4434 (N_4434,N_4139,N_3757);
or U4435 (N_4435,N_3746,N_3931);
and U4436 (N_4436,N_3860,N_2633);
nand U4437 (N_4437,N_3150,N_2383);
nand U4438 (N_4438,N_3954,In_2277);
nand U4439 (N_4439,N_4051,N_4031);
xor U4440 (N_4440,N_2539,N_2780);
nand U4441 (N_4441,N_3655,N_2310);
and U4442 (N_4442,In_2873,N_3793);
nand U4443 (N_4443,N_3254,N_3416);
nor U4444 (N_4444,N_2894,N_4080);
nor U4445 (N_4445,N_2342,N_2115);
or U4446 (N_4446,N_4017,N_3982);
or U4447 (N_4447,N_4192,N_3160);
nand U4448 (N_4448,N_1944,N_3476);
xor U4449 (N_4449,N_2886,N_2282);
xor U4450 (N_4450,N_3855,N_4065);
nor U4451 (N_4451,N_2875,N_3870);
nand U4452 (N_4452,N_2584,In_1488);
or U4453 (N_4453,N_4050,N_3529);
xor U4454 (N_4454,N_4034,N_3107);
nor U4455 (N_4455,N_1331,N_2940);
xnor U4456 (N_4456,N_3554,N_4088);
or U4457 (N_4457,N_4046,N_3420);
or U4458 (N_4458,N_3980,N_3807);
and U4459 (N_4459,N_3139,N_3643);
or U4460 (N_4460,N_686,N_4102);
nor U4461 (N_4461,N_2786,N_3877);
xnor U4462 (N_4462,N_4058,N_3811);
nand U4463 (N_4463,N_3819,N_4083);
nor U4464 (N_4464,N_3637,N_3632);
nor U4465 (N_4465,N_2969,N_3898);
or U4466 (N_4466,N_4184,N_4141);
xor U4467 (N_4467,N_3897,N_3703);
and U4468 (N_4468,N_3887,In_2326);
nand U4469 (N_4469,N_3266,In_59);
and U4470 (N_4470,N_1096,N_4110);
and U4471 (N_4471,N_3592,N_3551);
or U4472 (N_4472,N_4039,N_3179);
and U4473 (N_4473,N_4041,N_2923);
nand U4474 (N_4474,N_3905,N_3940);
nand U4475 (N_4475,N_4216,N_4018);
or U4476 (N_4476,N_4043,N_2360);
xor U4477 (N_4477,N_4129,In_2394);
and U4478 (N_4478,N_4020,N_4149);
nand U4479 (N_4479,N_3444,N_2331);
xor U4480 (N_4480,N_1312,N_2110);
or U4481 (N_4481,N_1423,N_4030);
or U4482 (N_4482,N_4187,N_3950);
or U4483 (N_4483,N_2773,N_3514);
nor U4484 (N_4484,N_3711,N_4185);
xor U4485 (N_4485,N_1954,In_2414);
or U4486 (N_4486,In_3828,N_3353);
nand U4487 (N_4487,N_4067,N_3663);
xnor U4488 (N_4488,N_3235,N_4119);
xnor U4489 (N_4489,N_4098,N_884);
or U4490 (N_4490,N_4053,In_3204);
or U4491 (N_4491,N_4094,N_3863);
nand U4492 (N_4492,N_3555,In_1618);
nand U4493 (N_4493,N_2511,N_3068);
nand U4494 (N_4494,N_3293,N_4242);
xor U4495 (N_4495,N_4244,In_4841);
or U4496 (N_4496,In_1980,N_3820);
nand U4497 (N_4497,N_4028,N_3971);
xor U4498 (N_4498,N_3601,N_4233);
nor U4499 (N_4499,In_1867,N_3932);
nand U4500 (N_4500,N_4388,N_4478);
xnor U4501 (N_4501,N_3678,N_4486);
nand U4502 (N_4502,N_4399,N_4209);
xnor U4503 (N_4503,N_4327,N_3694);
xor U4504 (N_4504,N_4374,N_2911);
or U4505 (N_4505,N_3138,N_4421);
and U4506 (N_4506,N_4398,N_3550);
and U4507 (N_4507,N_764,N_4448);
and U4508 (N_4508,N_3739,N_4322);
or U4509 (N_4509,N_4390,N_3374);
and U4510 (N_4510,N_2492,In_3625);
nor U4511 (N_4511,N_4491,N_3697);
nor U4512 (N_4512,N_4063,N_4469);
and U4513 (N_4513,N_4377,N_4231);
and U4514 (N_4514,N_4412,N_4089);
and U4515 (N_4515,N_3722,N_4401);
nor U4516 (N_4516,N_4237,N_4349);
nand U4517 (N_4517,N_3838,N_4445);
nand U4518 (N_4518,In_349,N_4456);
nand U4519 (N_4519,N_3831,N_2974);
and U4520 (N_4520,In_2378,N_4403);
nor U4521 (N_4521,N_3973,N_3232);
and U4522 (N_4522,N_3861,N_4206);
xor U4523 (N_4523,N_4357,N_4396);
or U4524 (N_4524,N_4359,N_4418);
xor U4525 (N_4525,N_4226,N_4474);
or U4526 (N_4526,N_4060,N_3871);
nor U4527 (N_4527,N_4385,N_4319);
or U4528 (N_4528,N_3461,N_4253);
xor U4529 (N_4529,N_4383,N_4458);
nand U4530 (N_4530,N_4373,N_4353);
and U4531 (N_4531,N_4395,N_3512);
nand U4532 (N_4532,N_2456,N_4171);
and U4533 (N_4533,N_4262,N_3915);
or U4534 (N_4534,N_4495,N_4314);
or U4535 (N_4535,N_4044,N_4414);
nor U4536 (N_4536,N_3689,N_4434);
nand U4537 (N_4537,N_3680,In_4643);
nand U4538 (N_4538,N_4246,N_4027);
nand U4539 (N_4539,N_4037,N_3073);
or U4540 (N_4540,In_217,N_210);
and U4541 (N_4541,N_3406,N_478);
or U4542 (N_4542,N_4406,N_4177);
xor U4543 (N_4543,N_911,N_4479);
nand U4544 (N_4544,N_4451,N_4300);
xnor U4545 (N_4545,N_4013,N_3986);
nand U4546 (N_4546,N_3804,N_4407);
nor U4547 (N_4547,N_2799,N_4097);
nand U4548 (N_4548,N_4266,N_3549);
and U4549 (N_4549,N_4333,N_4250);
nor U4550 (N_4550,N_4473,N_4425);
or U4551 (N_4551,N_1004,N_4330);
nand U4552 (N_4552,In_3411,N_4254);
nor U4553 (N_4553,N_4277,N_4394);
xnor U4554 (N_4554,N_4465,N_4283);
nor U4555 (N_4555,N_4023,N_4485);
nor U4556 (N_4556,In_4439,N_3560);
or U4557 (N_4557,N_4336,N_4367);
nand U4558 (N_4558,N_4306,N_4350);
nand U4559 (N_4559,N_3762,N_4008);
and U4560 (N_4560,N_4365,N_2955);
or U4561 (N_4561,In_1131,In_3593);
and U4562 (N_4562,N_4303,N_4124);
or U4563 (N_4563,In_401,N_1186);
nor U4564 (N_4564,N_4127,N_3716);
xor U4565 (N_4565,In_2060,N_4453);
and U4566 (N_4566,N_4297,N_4411);
nand U4567 (N_4567,N_4325,N_4329);
and U4568 (N_4568,N_4012,N_3983);
and U4569 (N_4569,N_4049,N_3706);
or U4570 (N_4570,N_4292,N_4299);
nor U4571 (N_4571,N_3598,N_3972);
nand U4572 (N_4572,N_4318,N_4273);
xor U4573 (N_4573,N_4393,N_4435);
nand U4574 (N_4574,N_4429,N_4386);
nand U4575 (N_4575,N_3705,N_4158);
xnor U4576 (N_4576,N_4038,N_4466);
nor U4577 (N_4577,N_4433,N_4459);
nand U4578 (N_4578,N_4309,N_4308);
nor U4579 (N_4579,N_3584,N_4307);
xnor U4580 (N_4580,N_4130,N_4035);
nand U4581 (N_4581,N_4096,N_4263);
or U4582 (N_4582,N_4070,N_4321);
nand U4583 (N_4583,N_4264,N_4428);
xor U4584 (N_4584,N_3969,N_4276);
nor U4585 (N_4585,N_4449,N_4188);
or U4586 (N_4586,N_4069,N_4369);
or U4587 (N_4587,N_4464,N_4343);
or U4588 (N_4588,N_4261,N_4275);
nand U4589 (N_4589,N_4346,N_3401);
or U4590 (N_4590,In_3257,N_4444);
and U4591 (N_4591,In_4262,N_4270);
or U4592 (N_4592,N_3895,In_4926);
and U4593 (N_4593,N_4441,N_3937);
or U4594 (N_4594,N_2743,N_4294);
and U4595 (N_4595,N_4402,N_4381);
and U4596 (N_4596,N_4274,N_4391);
nor U4597 (N_4597,N_4310,N_4081);
nor U4598 (N_4598,N_4010,N_4400);
nand U4599 (N_4599,N_3949,N_4301);
xor U4600 (N_4600,N_4068,N_4311);
nand U4601 (N_4601,N_2003,N_4033);
or U4602 (N_4602,N_4259,N_3460);
nor U4603 (N_4603,N_4476,N_4477);
xnor U4604 (N_4604,N_4488,N_4351);
or U4605 (N_4605,N_4431,N_4326);
and U4606 (N_4606,N_3362,N_4056);
nor U4607 (N_4607,N_4487,N_4032);
or U4608 (N_4608,N_4358,N_3843);
nand U4609 (N_4609,N_1443,N_4484);
nor U4610 (N_4610,N_784,N_4047);
nand U4611 (N_4611,N_4247,N_4007);
or U4612 (N_4612,N_4257,N_4175);
and U4613 (N_4613,N_4317,N_4265);
xor U4614 (N_4614,N_3365,N_1211);
xor U4615 (N_4615,N_3770,N_3707);
xnor U4616 (N_4616,N_4370,N_3590);
xnor U4617 (N_4617,N_4452,N_4410);
or U4618 (N_4618,N_4189,N_4494);
nand U4619 (N_4619,N_2236,N_4337);
xor U4620 (N_4620,N_3828,N_1743);
or U4621 (N_4621,N_3383,N_4417);
xor U4622 (N_4622,N_2666,N_4151);
or U4623 (N_4623,N_1849,N_3561);
nand U4624 (N_4624,N_4285,N_4191);
or U4625 (N_4625,N_4366,N_4338);
nor U4626 (N_4626,N_4438,N_4471);
or U4627 (N_4627,N_3349,N_3441);
nor U4628 (N_4628,N_4450,N_4066);
nor U4629 (N_4629,N_4413,N_4015);
or U4630 (N_4630,N_1943,N_3645);
and U4631 (N_4631,N_4085,N_4457);
and U4632 (N_4632,N_4382,N_3858);
nor U4633 (N_4633,N_3013,N_4397);
nand U4634 (N_4634,N_4320,N_3761);
or U4635 (N_4635,N_4363,N_3745);
nor U4636 (N_4636,N_4424,N_4360);
or U4637 (N_4637,N_4442,N_3948);
xor U4638 (N_4638,In_1166,N_4371);
nand U4639 (N_4639,In_2313,N_1962);
xor U4640 (N_4640,N_3372,N_4077);
xor U4641 (N_4641,N_4284,N_4298);
and U4642 (N_4642,N_3826,In_4098);
nor U4643 (N_4643,N_3994,N_3726);
nand U4644 (N_4644,N_4430,N_3124);
nand U4645 (N_4645,N_4447,N_4121);
nor U4646 (N_4646,N_4362,N_4282);
nor U4647 (N_4647,N_4461,N_550);
and U4648 (N_4648,N_4304,N_4324);
or U4649 (N_4649,N_4290,N_4348);
and U4650 (N_4650,N_4169,N_4463);
nor U4651 (N_4651,N_2650,N_4021);
xnor U4652 (N_4652,N_4239,N_4267);
or U4653 (N_4653,N_4295,N_3644);
xor U4654 (N_4654,N_4462,In_1680);
nor U4655 (N_4655,N_4493,In_3062);
nand U4656 (N_4656,N_2286,N_4443);
nor U4657 (N_4657,In_1636,N_4436);
nor U4658 (N_4658,N_4214,N_4352);
nor U4659 (N_4659,In_2674,N_4302);
nand U4660 (N_4660,N_4439,N_4078);
and U4661 (N_4661,N_4296,N_4251);
nor U4662 (N_4662,N_4454,N_4258);
or U4663 (N_4663,N_4256,N_3245);
or U4664 (N_4664,N_4120,N_3849);
and U4665 (N_4665,N_3823,N_4286);
nand U4666 (N_4666,N_4271,N_4499);
or U4667 (N_4667,N_2549,N_4334);
or U4668 (N_4668,N_4347,N_4482);
nand U4669 (N_4669,N_3515,N_2804);
and U4670 (N_4670,N_4279,N_4409);
nand U4671 (N_4671,In_1753,N_4217);
nand U4672 (N_4672,N_4378,N_1600);
or U4673 (N_4673,N_4492,N_4144);
xnor U4674 (N_4674,N_4332,N_4203);
xor U4675 (N_4675,In_458,N_4323);
or U4676 (N_4676,N_2727,N_4489);
and U4677 (N_4677,N_4340,N_4212);
nor U4678 (N_4678,N_4278,N_3582);
or U4679 (N_4679,In_3469,N_4255);
or U4680 (N_4680,N_4293,In_2041);
xor U4681 (N_4681,N_4316,N_3787);
nor U4682 (N_4682,N_4345,N_4004);
nor U4683 (N_4683,N_2059,N_3917);
nand U4684 (N_4684,N_4483,N_4467);
xnor U4685 (N_4685,N_4426,N_4422);
nor U4686 (N_4686,N_4164,N_4138);
and U4687 (N_4687,N_4260,N_3501);
xnor U4688 (N_4688,N_4315,N_3653);
or U4689 (N_4689,N_3382,N_3848);
and U4690 (N_4690,N_4475,N_4014);
or U4691 (N_4691,N_3763,N_4392);
nor U4692 (N_4692,N_4113,N_4341);
or U4693 (N_4693,N_4086,N_4415);
nor U4694 (N_4694,N_4052,N_3878);
nor U4695 (N_4695,N_4287,In_1004);
and U4696 (N_4696,N_3616,N_4288);
and U4697 (N_4697,N_45,N_3999);
nand U4698 (N_4698,N_4229,In_326);
or U4699 (N_4699,N_4268,In_729);
nand U4700 (N_4700,N_4178,N_4496);
or U4701 (N_4701,N_4331,N_4384);
and U4702 (N_4702,N_4356,N_4099);
or U4703 (N_4703,N_4195,N_4375);
nor U4704 (N_4704,N_4472,N_4368);
xnor U4705 (N_4705,N_4241,N_4252);
and U4706 (N_4706,N_4339,N_2967);
xor U4707 (N_4707,N_4423,N_4416);
and U4708 (N_4708,N_4361,N_3955);
xnor U4709 (N_4709,N_3623,N_4372);
xor U4710 (N_4710,N_3945,N_4291);
xnor U4711 (N_4711,N_4379,N_4405);
nor U4712 (N_4712,N_4344,N_3747);
nor U4713 (N_4713,N_4146,N_3517);
or U4714 (N_4714,In_613,N_4408);
nand U4715 (N_4715,N_4387,N_3783);
nor U4716 (N_4716,N_4100,N_3486);
or U4717 (N_4717,N_4364,N_4305);
nor U4718 (N_4718,N_3676,N_4355);
and U4719 (N_4719,N_3272,N_4312);
nor U4720 (N_4720,N_4335,N_4432);
xnor U4721 (N_4721,N_4076,N_4419);
or U4722 (N_4722,In_2011,N_4498);
nor U4723 (N_4723,N_4150,N_4225);
nand U4724 (N_4724,N_4313,N_4154);
and U4725 (N_4725,N_4455,N_3267);
nor U4726 (N_4726,N_4497,N_3882);
and U4727 (N_4727,N_4460,N_3540);
xnor U4728 (N_4728,N_4221,N_4280);
or U4729 (N_4729,N_4210,N_4437);
nand U4730 (N_4730,N_4354,N_4490);
nand U4731 (N_4731,N_3687,N_4427);
xnor U4732 (N_4732,N_3817,N_4480);
xnor U4733 (N_4733,N_4376,N_4272);
xor U4734 (N_4734,N_3140,N_2962);
nand U4735 (N_4735,N_4380,N_4173);
and U4736 (N_4736,N_2250,N_4481);
or U4737 (N_4737,N_3363,N_4389);
xnor U4738 (N_4738,N_3583,N_4281);
nand U4739 (N_4739,N_3127,N_4440);
or U4740 (N_4740,N_4470,In_101);
nand U4741 (N_4741,N_4404,In_1580);
and U4742 (N_4742,N_3935,N_3825);
xor U4743 (N_4743,N_4142,N_4446);
xnor U4744 (N_4744,N_3936,N_4342);
or U4745 (N_4745,N_4269,N_3952);
nand U4746 (N_4746,N_4289,N_3991);
nand U4747 (N_4747,N_4000,N_3498);
nor U4748 (N_4748,N_4420,N_3934);
nor U4749 (N_4749,N_4468,N_4328);
or U4750 (N_4750,N_4532,N_4650);
and U4751 (N_4751,N_4587,N_4685);
or U4752 (N_4752,N_4656,N_4707);
or U4753 (N_4753,N_4582,N_4588);
nor U4754 (N_4754,N_4573,N_4600);
and U4755 (N_4755,N_4671,N_4636);
nor U4756 (N_4756,N_4736,N_4559);
xnor U4757 (N_4757,N_4729,N_4741);
nand U4758 (N_4758,N_4718,N_4510);
or U4759 (N_4759,N_4565,N_4611);
nor U4760 (N_4760,N_4575,N_4567);
nand U4761 (N_4761,N_4562,N_4698);
xor U4762 (N_4762,N_4603,N_4618);
and U4763 (N_4763,N_4522,N_4693);
and U4764 (N_4764,N_4642,N_4675);
nand U4765 (N_4765,N_4597,N_4748);
nand U4766 (N_4766,N_4609,N_4570);
and U4767 (N_4767,N_4605,N_4647);
xor U4768 (N_4768,N_4739,N_4552);
nand U4769 (N_4769,N_4576,N_4502);
nand U4770 (N_4770,N_4749,N_4688);
nor U4771 (N_4771,N_4527,N_4695);
nand U4772 (N_4772,N_4711,N_4547);
and U4773 (N_4773,N_4732,N_4699);
or U4774 (N_4774,N_4624,N_4670);
and U4775 (N_4775,N_4725,N_4604);
nand U4776 (N_4776,N_4726,N_4507);
nor U4777 (N_4777,N_4542,N_4579);
nor U4778 (N_4778,N_4541,N_4703);
or U4779 (N_4779,N_4723,N_4713);
nor U4780 (N_4780,N_4625,N_4684);
and U4781 (N_4781,N_4512,N_4568);
nor U4782 (N_4782,N_4683,N_4538);
nand U4783 (N_4783,N_4702,N_4606);
and U4784 (N_4784,N_4710,N_4654);
xnor U4785 (N_4785,N_4530,N_4546);
and U4786 (N_4786,N_4680,N_4630);
xnor U4787 (N_4787,N_4731,N_4730);
xnor U4788 (N_4788,N_4679,N_4746);
xor U4789 (N_4789,N_4619,N_4652);
and U4790 (N_4790,N_4577,N_4591);
and U4791 (N_4791,N_4553,N_4687);
and U4792 (N_4792,N_4715,N_4673);
nor U4793 (N_4793,N_4590,N_4586);
nor U4794 (N_4794,N_4583,N_4602);
or U4795 (N_4795,N_4712,N_4706);
and U4796 (N_4796,N_4716,N_4719);
xor U4797 (N_4797,N_4520,N_4742);
xor U4798 (N_4798,N_4528,N_4620);
nor U4799 (N_4799,N_4536,N_4662);
nand U4800 (N_4800,N_4515,N_4556);
nand U4801 (N_4801,N_4627,N_4519);
or U4802 (N_4802,N_4517,N_4596);
nor U4803 (N_4803,N_4561,N_4529);
and U4804 (N_4804,N_4724,N_4728);
or U4805 (N_4805,N_4628,N_4607);
nand U4806 (N_4806,N_4646,N_4653);
nor U4807 (N_4807,N_4555,N_4660);
and U4808 (N_4808,N_4734,N_4681);
nor U4809 (N_4809,N_4505,N_4506);
nand U4810 (N_4810,N_4655,N_4735);
or U4811 (N_4811,N_4664,N_4539);
nand U4812 (N_4812,N_4640,N_4543);
nor U4813 (N_4813,N_4659,N_4544);
xor U4814 (N_4814,N_4641,N_4523);
or U4815 (N_4815,N_4580,N_4563);
nand U4816 (N_4816,N_4593,N_4557);
nor U4817 (N_4817,N_4566,N_4548);
xnor U4818 (N_4818,N_4747,N_4701);
and U4819 (N_4819,N_4537,N_4622);
xnor U4820 (N_4820,N_4638,N_4694);
nand U4821 (N_4821,N_4521,N_4540);
or U4822 (N_4822,N_4717,N_4500);
and U4823 (N_4823,N_4599,N_4745);
and U4824 (N_4824,N_4564,N_4677);
and U4825 (N_4825,N_4631,N_4569);
xor U4826 (N_4826,N_4614,N_4740);
xnor U4827 (N_4827,N_4509,N_4669);
xor U4828 (N_4828,N_4550,N_4615);
xor U4829 (N_4829,N_4727,N_4692);
or U4830 (N_4830,N_4644,N_4594);
nand U4831 (N_4831,N_4709,N_4595);
nand U4832 (N_4832,N_4589,N_4633);
or U4833 (N_4833,N_4578,N_4672);
nor U4834 (N_4834,N_4639,N_4534);
xnor U4835 (N_4835,N_4616,N_4551);
or U4836 (N_4836,N_4738,N_4558);
nor U4837 (N_4837,N_4643,N_4686);
or U4838 (N_4838,N_4610,N_4733);
and U4839 (N_4839,N_4661,N_4572);
nor U4840 (N_4840,N_4645,N_4689);
and U4841 (N_4841,N_4598,N_4514);
nand U4842 (N_4842,N_4744,N_4533);
or U4843 (N_4843,N_4584,N_4560);
or U4844 (N_4844,N_4667,N_4508);
or U4845 (N_4845,N_4743,N_4721);
nand U4846 (N_4846,N_4714,N_4626);
nand U4847 (N_4847,N_4545,N_4549);
or U4848 (N_4848,N_4658,N_4581);
xor U4849 (N_4849,N_4666,N_4696);
and U4850 (N_4850,N_4621,N_4665);
and U4851 (N_4851,N_4649,N_4674);
and U4852 (N_4852,N_4601,N_4682);
or U4853 (N_4853,N_4676,N_4690);
and U4854 (N_4854,N_4678,N_4613);
and U4855 (N_4855,N_4574,N_4526);
xor U4856 (N_4856,N_4657,N_4511);
or U4857 (N_4857,N_4635,N_4691);
nand U4858 (N_4858,N_4525,N_4704);
and U4859 (N_4859,N_4700,N_4722);
nand U4860 (N_4860,N_4663,N_4554);
xor U4861 (N_4861,N_4535,N_4608);
and U4862 (N_4862,N_4697,N_4617);
nand U4863 (N_4863,N_4705,N_4531);
and U4864 (N_4864,N_4501,N_4737);
or U4865 (N_4865,N_4503,N_4571);
and U4866 (N_4866,N_4623,N_4637);
xor U4867 (N_4867,N_4668,N_4651);
nand U4868 (N_4868,N_4524,N_4592);
nand U4869 (N_4869,N_4516,N_4518);
or U4870 (N_4870,N_4634,N_4612);
nor U4871 (N_4871,N_4629,N_4720);
nand U4872 (N_4872,N_4708,N_4632);
nor U4873 (N_4873,N_4585,N_4504);
and U4874 (N_4874,N_4648,N_4513);
or U4875 (N_4875,N_4717,N_4525);
xnor U4876 (N_4876,N_4639,N_4527);
or U4877 (N_4877,N_4637,N_4678);
nor U4878 (N_4878,N_4719,N_4627);
xnor U4879 (N_4879,N_4516,N_4546);
xnor U4880 (N_4880,N_4749,N_4587);
or U4881 (N_4881,N_4541,N_4607);
or U4882 (N_4882,N_4628,N_4525);
or U4883 (N_4883,N_4738,N_4563);
xnor U4884 (N_4884,N_4556,N_4640);
nand U4885 (N_4885,N_4580,N_4502);
or U4886 (N_4886,N_4721,N_4735);
and U4887 (N_4887,N_4673,N_4724);
and U4888 (N_4888,N_4565,N_4636);
or U4889 (N_4889,N_4564,N_4703);
nor U4890 (N_4890,N_4749,N_4644);
and U4891 (N_4891,N_4582,N_4554);
xnor U4892 (N_4892,N_4733,N_4711);
and U4893 (N_4893,N_4713,N_4655);
xor U4894 (N_4894,N_4622,N_4550);
nor U4895 (N_4895,N_4733,N_4671);
and U4896 (N_4896,N_4625,N_4653);
and U4897 (N_4897,N_4634,N_4593);
or U4898 (N_4898,N_4502,N_4647);
xnor U4899 (N_4899,N_4604,N_4606);
or U4900 (N_4900,N_4730,N_4531);
nand U4901 (N_4901,N_4690,N_4619);
nor U4902 (N_4902,N_4738,N_4592);
nand U4903 (N_4903,N_4659,N_4534);
and U4904 (N_4904,N_4549,N_4585);
or U4905 (N_4905,N_4501,N_4635);
or U4906 (N_4906,N_4725,N_4707);
and U4907 (N_4907,N_4714,N_4682);
nor U4908 (N_4908,N_4502,N_4507);
and U4909 (N_4909,N_4506,N_4628);
nor U4910 (N_4910,N_4518,N_4687);
nand U4911 (N_4911,N_4732,N_4704);
and U4912 (N_4912,N_4646,N_4596);
nor U4913 (N_4913,N_4552,N_4668);
or U4914 (N_4914,N_4748,N_4532);
or U4915 (N_4915,N_4661,N_4604);
and U4916 (N_4916,N_4532,N_4681);
and U4917 (N_4917,N_4657,N_4519);
and U4918 (N_4918,N_4734,N_4625);
nor U4919 (N_4919,N_4568,N_4736);
xnor U4920 (N_4920,N_4579,N_4532);
nor U4921 (N_4921,N_4665,N_4664);
xnor U4922 (N_4922,N_4575,N_4626);
xnor U4923 (N_4923,N_4618,N_4714);
and U4924 (N_4924,N_4651,N_4559);
nor U4925 (N_4925,N_4724,N_4684);
and U4926 (N_4926,N_4705,N_4589);
or U4927 (N_4927,N_4748,N_4691);
and U4928 (N_4928,N_4734,N_4700);
xnor U4929 (N_4929,N_4541,N_4620);
and U4930 (N_4930,N_4624,N_4608);
and U4931 (N_4931,N_4683,N_4524);
nand U4932 (N_4932,N_4528,N_4697);
and U4933 (N_4933,N_4586,N_4625);
nand U4934 (N_4934,N_4628,N_4533);
and U4935 (N_4935,N_4695,N_4533);
or U4936 (N_4936,N_4519,N_4603);
xor U4937 (N_4937,N_4681,N_4643);
and U4938 (N_4938,N_4603,N_4671);
nand U4939 (N_4939,N_4559,N_4682);
nand U4940 (N_4940,N_4632,N_4744);
nand U4941 (N_4941,N_4725,N_4700);
and U4942 (N_4942,N_4685,N_4747);
or U4943 (N_4943,N_4692,N_4687);
or U4944 (N_4944,N_4705,N_4714);
xnor U4945 (N_4945,N_4584,N_4730);
xnor U4946 (N_4946,N_4683,N_4549);
or U4947 (N_4947,N_4647,N_4707);
xnor U4948 (N_4948,N_4677,N_4533);
nor U4949 (N_4949,N_4710,N_4628);
or U4950 (N_4950,N_4582,N_4671);
and U4951 (N_4951,N_4749,N_4697);
or U4952 (N_4952,N_4727,N_4648);
xor U4953 (N_4953,N_4630,N_4511);
or U4954 (N_4954,N_4619,N_4744);
nand U4955 (N_4955,N_4631,N_4607);
or U4956 (N_4956,N_4566,N_4603);
and U4957 (N_4957,N_4652,N_4561);
nor U4958 (N_4958,N_4586,N_4667);
nand U4959 (N_4959,N_4558,N_4742);
nor U4960 (N_4960,N_4509,N_4649);
and U4961 (N_4961,N_4688,N_4508);
or U4962 (N_4962,N_4583,N_4655);
nand U4963 (N_4963,N_4515,N_4608);
nand U4964 (N_4964,N_4539,N_4737);
xnor U4965 (N_4965,N_4590,N_4538);
nand U4966 (N_4966,N_4718,N_4505);
xnor U4967 (N_4967,N_4603,N_4571);
nor U4968 (N_4968,N_4544,N_4730);
and U4969 (N_4969,N_4550,N_4599);
and U4970 (N_4970,N_4561,N_4733);
nor U4971 (N_4971,N_4702,N_4616);
xor U4972 (N_4972,N_4531,N_4739);
xor U4973 (N_4973,N_4507,N_4543);
nand U4974 (N_4974,N_4508,N_4509);
nand U4975 (N_4975,N_4732,N_4568);
nand U4976 (N_4976,N_4532,N_4616);
and U4977 (N_4977,N_4538,N_4515);
nor U4978 (N_4978,N_4537,N_4515);
nand U4979 (N_4979,N_4570,N_4736);
nor U4980 (N_4980,N_4504,N_4573);
nand U4981 (N_4981,N_4717,N_4620);
xor U4982 (N_4982,N_4715,N_4697);
or U4983 (N_4983,N_4653,N_4575);
or U4984 (N_4984,N_4563,N_4596);
or U4985 (N_4985,N_4686,N_4566);
nor U4986 (N_4986,N_4609,N_4505);
nand U4987 (N_4987,N_4656,N_4730);
or U4988 (N_4988,N_4536,N_4654);
and U4989 (N_4989,N_4687,N_4728);
nor U4990 (N_4990,N_4625,N_4668);
or U4991 (N_4991,N_4585,N_4602);
nor U4992 (N_4992,N_4559,N_4737);
nor U4993 (N_4993,N_4591,N_4531);
nand U4994 (N_4994,N_4630,N_4654);
xor U4995 (N_4995,N_4510,N_4656);
nand U4996 (N_4996,N_4650,N_4543);
nor U4997 (N_4997,N_4676,N_4680);
xor U4998 (N_4998,N_4723,N_4748);
or U4999 (N_4999,N_4636,N_4603);
and U5000 (N_5000,N_4787,N_4774);
and U5001 (N_5001,N_4895,N_4764);
or U5002 (N_5002,N_4970,N_4797);
nand U5003 (N_5003,N_4966,N_4785);
and U5004 (N_5004,N_4838,N_4858);
nand U5005 (N_5005,N_4980,N_4904);
and U5006 (N_5006,N_4820,N_4807);
nand U5007 (N_5007,N_4965,N_4977);
and U5008 (N_5008,N_4799,N_4836);
nor U5009 (N_5009,N_4892,N_4974);
xor U5010 (N_5010,N_4953,N_4755);
and U5011 (N_5011,N_4916,N_4777);
nor U5012 (N_5012,N_4770,N_4899);
nand U5013 (N_5013,N_4998,N_4833);
nand U5014 (N_5014,N_4902,N_4789);
nor U5015 (N_5015,N_4979,N_4988);
xor U5016 (N_5016,N_4927,N_4926);
nand U5017 (N_5017,N_4929,N_4985);
nand U5018 (N_5018,N_4976,N_4760);
nor U5019 (N_5019,N_4795,N_4851);
nand U5020 (N_5020,N_4995,N_4834);
nand U5021 (N_5021,N_4862,N_4948);
nand U5022 (N_5022,N_4873,N_4781);
nor U5023 (N_5023,N_4894,N_4981);
or U5024 (N_5024,N_4863,N_4945);
xnor U5025 (N_5025,N_4861,N_4989);
nor U5026 (N_5026,N_4957,N_4925);
nor U5027 (N_5027,N_4960,N_4878);
nor U5028 (N_5028,N_4994,N_4803);
nor U5029 (N_5029,N_4859,N_4896);
or U5030 (N_5030,N_4923,N_4959);
nor U5031 (N_5031,N_4829,N_4752);
nor U5032 (N_5032,N_4792,N_4866);
xnor U5033 (N_5033,N_4919,N_4881);
nand U5034 (N_5034,N_4847,N_4898);
nor U5035 (N_5035,N_4767,N_4941);
nand U5036 (N_5036,N_4986,N_4889);
xnor U5037 (N_5037,N_4796,N_4810);
nand U5038 (N_5038,N_4947,N_4907);
xor U5039 (N_5039,N_4993,N_4814);
and U5040 (N_5040,N_4900,N_4903);
nor U5041 (N_5041,N_4938,N_4856);
nand U5042 (N_5042,N_4826,N_4992);
or U5043 (N_5043,N_4805,N_4932);
xor U5044 (N_5044,N_4958,N_4906);
nor U5045 (N_5045,N_4844,N_4751);
or U5046 (N_5046,N_4936,N_4830);
and U5047 (N_5047,N_4968,N_4909);
or U5048 (N_5048,N_4943,N_4937);
xnor U5049 (N_5049,N_4821,N_4772);
nand U5050 (N_5050,N_4759,N_4818);
or U5051 (N_5051,N_4920,N_4883);
xor U5052 (N_5052,N_4912,N_4944);
nor U5053 (N_5053,N_4806,N_4869);
nor U5054 (N_5054,N_4969,N_4956);
or U5055 (N_5055,N_4880,N_4835);
nor U5056 (N_5056,N_4877,N_4850);
and U5057 (N_5057,N_4816,N_4973);
and U5058 (N_5058,N_4779,N_4884);
nor U5059 (N_5059,N_4813,N_4815);
xor U5060 (N_5060,N_4922,N_4786);
xor U5061 (N_5061,N_4822,N_4971);
xnor U5062 (N_5062,N_4778,N_4954);
and U5063 (N_5063,N_4864,N_4918);
nor U5064 (N_5064,N_4766,N_4893);
and U5065 (N_5065,N_4921,N_4784);
nand U5066 (N_5066,N_4855,N_4933);
nand U5067 (N_5067,N_4867,N_4865);
nor U5068 (N_5068,N_4999,N_4996);
nor U5069 (N_5069,N_4931,N_4843);
and U5070 (N_5070,N_4963,N_4857);
and U5071 (N_5071,N_4972,N_4901);
nor U5072 (N_5072,N_4825,N_4769);
nor U5073 (N_5073,N_4871,N_4848);
nor U5074 (N_5074,N_4991,N_4773);
nand U5075 (N_5075,N_4845,N_4808);
xor U5076 (N_5076,N_4776,N_4950);
xor U5077 (N_5077,N_4891,N_4886);
and U5078 (N_5078,N_4750,N_4832);
and U5079 (N_5079,N_4897,N_4946);
xnor U5080 (N_5080,N_4951,N_4917);
xnor U5081 (N_5081,N_4840,N_4793);
nand U5082 (N_5082,N_4928,N_4828);
xnor U5083 (N_5083,N_4768,N_4854);
xnor U5084 (N_5084,N_4765,N_4911);
xnor U5085 (N_5085,N_4964,N_4987);
and U5086 (N_5086,N_4853,N_4924);
nor U5087 (N_5087,N_4827,N_4935);
nand U5088 (N_5088,N_4756,N_4754);
and U5089 (N_5089,N_4875,N_4775);
xnor U5090 (N_5090,N_4819,N_4961);
nor U5091 (N_5091,N_4791,N_4952);
nand U5092 (N_5092,N_4842,N_4967);
xor U5093 (N_5093,N_4790,N_4915);
nor U5094 (N_5094,N_4983,N_4801);
and U5095 (N_5095,N_4860,N_4870);
nor U5096 (N_5096,N_4890,N_4783);
or U5097 (N_5097,N_4868,N_4990);
nor U5098 (N_5098,N_4905,N_4913);
xor U5099 (N_5099,N_4975,N_4885);
nand U5100 (N_5100,N_4794,N_4800);
xnor U5101 (N_5101,N_4780,N_4802);
and U5102 (N_5102,N_4824,N_4812);
nand U5103 (N_5103,N_4852,N_4978);
or U5104 (N_5104,N_4888,N_4837);
and U5105 (N_5105,N_4798,N_4934);
nand U5106 (N_5106,N_4753,N_4879);
and U5107 (N_5107,N_4940,N_4876);
nand U5108 (N_5108,N_4949,N_4908);
nor U5109 (N_5109,N_4782,N_4839);
or U5110 (N_5110,N_4887,N_4984);
nor U5111 (N_5111,N_4942,N_4882);
and U5112 (N_5112,N_4811,N_4809);
or U5113 (N_5113,N_4788,N_4841);
xnor U5114 (N_5114,N_4849,N_4910);
xor U5115 (N_5115,N_4982,N_4817);
xor U5116 (N_5116,N_4823,N_4771);
nor U5117 (N_5117,N_4846,N_4761);
xnor U5118 (N_5118,N_4872,N_4831);
nor U5119 (N_5119,N_4762,N_4930);
or U5120 (N_5120,N_4962,N_4874);
nand U5121 (N_5121,N_4804,N_4757);
xnor U5122 (N_5122,N_4763,N_4758);
or U5123 (N_5123,N_4914,N_4939);
nor U5124 (N_5124,N_4955,N_4997);
or U5125 (N_5125,N_4858,N_4781);
and U5126 (N_5126,N_4858,N_4814);
nor U5127 (N_5127,N_4859,N_4793);
nand U5128 (N_5128,N_4950,N_4833);
or U5129 (N_5129,N_4855,N_4752);
nor U5130 (N_5130,N_4888,N_4935);
xnor U5131 (N_5131,N_4795,N_4766);
or U5132 (N_5132,N_4932,N_4793);
and U5133 (N_5133,N_4913,N_4784);
and U5134 (N_5134,N_4838,N_4964);
or U5135 (N_5135,N_4992,N_4903);
nand U5136 (N_5136,N_4824,N_4794);
xnor U5137 (N_5137,N_4788,N_4918);
xor U5138 (N_5138,N_4948,N_4873);
xnor U5139 (N_5139,N_4840,N_4894);
nor U5140 (N_5140,N_4896,N_4761);
nor U5141 (N_5141,N_4940,N_4860);
nor U5142 (N_5142,N_4817,N_4972);
nor U5143 (N_5143,N_4893,N_4865);
nor U5144 (N_5144,N_4854,N_4811);
nand U5145 (N_5145,N_4982,N_4775);
nor U5146 (N_5146,N_4890,N_4847);
and U5147 (N_5147,N_4840,N_4891);
nor U5148 (N_5148,N_4780,N_4914);
or U5149 (N_5149,N_4815,N_4865);
nor U5150 (N_5150,N_4936,N_4888);
and U5151 (N_5151,N_4955,N_4848);
nor U5152 (N_5152,N_4999,N_4922);
xnor U5153 (N_5153,N_4864,N_4839);
or U5154 (N_5154,N_4820,N_4974);
xnor U5155 (N_5155,N_4979,N_4924);
or U5156 (N_5156,N_4911,N_4845);
nand U5157 (N_5157,N_4908,N_4960);
nor U5158 (N_5158,N_4789,N_4761);
or U5159 (N_5159,N_4818,N_4955);
xor U5160 (N_5160,N_4902,N_4803);
xnor U5161 (N_5161,N_4754,N_4862);
nor U5162 (N_5162,N_4830,N_4853);
nand U5163 (N_5163,N_4827,N_4793);
and U5164 (N_5164,N_4904,N_4935);
and U5165 (N_5165,N_4879,N_4810);
or U5166 (N_5166,N_4966,N_4889);
and U5167 (N_5167,N_4940,N_4933);
xnor U5168 (N_5168,N_4864,N_4798);
nor U5169 (N_5169,N_4964,N_4968);
nor U5170 (N_5170,N_4771,N_4983);
nand U5171 (N_5171,N_4969,N_4984);
nand U5172 (N_5172,N_4875,N_4857);
nand U5173 (N_5173,N_4864,N_4847);
or U5174 (N_5174,N_4892,N_4841);
xnor U5175 (N_5175,N_4840,N_4767);
nand U5176 (N_5176,N_4869,N_4886);
nor U5177 (N_5177,N_4968,N_4820);
nand U5178 (N_5178,N_4992,N_4838);
or U5179 (N_5179,N_4984,N_4999);
nand U5180 (N_5180,N_4988,N_4881);
or U5181 (N_5181,N_4999,N_4892);
or U5182 (N_5182,N_4782,N_4965);
nor U5183 (N_5183,N_4954,N_4892);
or U5184 (N_5184,N_4881,N_4863);
or U5185 (N_5185,N_4809,N_4926);
or U5186 (N_5186,N_4837,N_4890);
and U5187 (N_5187,N_4841,N_4836);
nor U5188 (N_5188,N_4866,N_4775);
and U5189 (N_5189,N_4952,N_4958);
and U5190 (N_5190,N_4905,N_4808);
nand U5191 (N_5191,N_4781,N_4952);
or U5192 (N_5192,N_4951,N_4781);
or U5193 (N_5193,N_4796,N_4784);
nand U5194 (N_5194,N_4873,N_4893);
or U5195 (N_5195,N_4800,N_4971);
and U5196 (N_5196,N_4784,N_4898);
nor U5197 (N_5197,N_4886,N_4790);
and U5198 (N_5198,N_4808,N_4811);
nand U5199 (N_5199,N_4898,N_4930);
or U5200 (N_5200,N_4876,N_4856);
nor U5201 (N_5201,N_4955,N_4922);
nand U5202 (N_5202,N_4848,N_4984);
nand U5203 (N_5203,N_4766,N_4797);
nor U5204 (N_5204,N_4909,N_4862);
and U5205 (N_5205,N_4894,N_4956);
nor U5206 (N_5206,N_4859,N_4870);
and U5207 (N_5207,N_4823,N_4795);
and U5208 (N_5208,N_4978,N_4953);
xnor U5209 (N_5209,N_4870,N_4943);
and U5210 (N_5210,N_4939,N_4877);
nor U5211 (N_5211,N_4931,N_4796);
xnor U5212 (N_5212,N_4773,N_4835);
or U5213 (N_5213,N_4967,N_4890);
xor U5214 (N_5214,N_4951,N_4836);
xnor U5215 (N_5215,N_4999,N_4936);
and U5216 (N_5216,N_4971,N_4819);
nand U5217 (N_5217,N_4862,N_4944);
nor U5218 (N_5218,N_4951,N_4881);
nand U5219 (N_5219,N_4907,N_4814);
xnor U5220 (N_5220,N_4877,N_4827);
xor U5221 (N_5221,N_4881,N_4852);
or U5222 (N_5222,N_4852,N_4867);
or U5223 (N_5223,N_4890,N_4903);
and U5224 (N_5224,N_4954,N_4863);
or U5225 (N_5225,N_4972,N_4860);
xor U5226 (N_5226,N_4981,N_4855);
or U5227 (N_5227,N_4823,N_4987);
and U5228 (N_5228,N_4937,N_4818);
and U5229 (N_5229,N_4778,N_4823);
or U5230 (N_5230,N_4963,N_4778);
nor U5231 (N_5231,N_4793,N_4860);
nand U5232 (N_5232,N_4786,N_4995);
nor U5233 (N_5233,N_4906,N_4852);
and U5234 (N_5234,N_4916,N_4941);
or U5235 (N_5235,N_4888,N_4813);
nor U5236 (N_5236,N_4917,N_4771);
or U5237 (N_5237,N_4851,N_4773);
nor U5238 (N_5238,N_4774,N_4957);
and U5239 (N_5239,N_4760,N_4883);
nor U5240 (N_5240,N_4941,N_4794);
and U5241 (N_5241,N_4764,N_4791);
nor U5242 (N_5242,N_4770,N_4994);
and U5243 (N_5243,N_4982,N_4810);
xor U5244 (N_5244,N_4906,N_4837);
and U5245 (N_5245,N_4889,N_4996);
or U5246 (N_5246,N_4880,N_4875);
nor U5247 (N_5247,N_4809,N_4866);
xor U5248 (N_5248,N_4809,N_4977);
or U5249 (N_5249,N_4936,N_4991);
or U5250 (N_5250,N_5205,N_5066);
nor U5251 (N_5251,N_5120,N_5098);
nor U5252 (N_5252,N_5024,N_5165);
and U5253 (N_5253,N_5063,N_5065);
xnor U5254 (N_5254,N_5008,N_5203);
nor U5255 (N_5255,N_5154,N_5164);
and U5256 (N_5256,N_5147,N_5187);
xor U5257 (N_5257,N_5029,N_5102);
nand U5258 (N_5258,N_5182,N_5031);
xnor U5259 (N_5259,N_5118,N_5057);
nand U5260 (N_5260,N_5109,N_5144);
and U5261 (N_5261,N_5050,N_5124);
nand U5262 (N_5262,N_5135,N_5012);
or U5263 (N_5263,N_5219,N_5070);
nand U5264 (N_5264,N_5074,N_5143);
or U5265 (N_5265,N_5104,N_5177);
xnor U5266 (N_5266,N_5033,N_5045);
and U5267 (N_5267,N_5195,N_5239);
nand U5268 (N_5268,N_5011,N_5249);
and U5269 (N_5269,N_5137,N_5041);
and U5270 (N_5270,N_5148,N_5072);
and U5271 (N_5271,N_5035,N_5176);
nand U5272 (N_5272,N_5068,N_5229);
xor U5273 (N_5273,N_5244,N_5034);
and U5274 (N_5274,N_5183,N_5119);
and U5275 (N_5275,N_5149,N_5092);
or U5276 (N_5276,N_5071,N_5095);
nor U5277 (N_5277,N_5038,N_5077);
nor U5278 (N_5278,N_5236,N_5129);
nor U5279 (N_5279,N_5245,N_5049);
and U5280 (N_5280,N_5042,N_5016);
xor U5281 (N_5281,N_5216,N_5030);
or U5282 (N_5282,N_5196,N_5127);
nor U5283 (N_5283,N_5204,N_5214);
and U5284 (N_5284,N_5125,N_5234);
nand U5285 (N_5285,N_5039,N_5108);
or U5286 (N_5286,N_5163,N_5220);
nand U5287 (N_5287,N_5088,N_5152);
nor U5288 (N_5288,N_5105,N_5082);
nor U5289 (N_5289,N_5180,N_5169);
xnor U5290 (N_5290,N_5221,N_5084);
xnor U5291 (N_5291,N_5218,N_5213);
nor U5292 (N_5292,N_5112,N_5116);
nand U5293 (N_5293,N_5043,N_5076);
xnor U5294 (N_5294,N_5141,N_5058);
or U5295 (N_5295,N_5067,N_5191);
and U5296 (N_5296,N_5040,N_5159);
xnor U5297 (N_5297,N_5210,N_5190);
or U5298 (N_5298,N_5202,N_5054);
nand U5299 (N_5299,N_5200,N_5010);
and U5300 (N_5300,N_5060,N_5184);
and U5301 (N_5301,N_5231,N_5197);
nor U5302 (N_5302,N_5132,N_5208);
or U5303 (N_5303,N_5002,N_5091);
and U5304 (N_5304,N_5153,N_5138);
and U5305 (N_5305,N_5053,N_5003);
and U5306 (N_5306,N_5121,N_5174);
xor U5307 (N_5307,N_5128,N_5188);
nand U5308 (N_5308,N_5048,N_5171);
or U5309 (N_5309,N_5090,N_5117);
xor U5310 (N_5310,N_5009,N_5007);
nand U5311 (N_5311,N_5162,N_5115);
nor U5312 (N_5312,N_5193,N_5113);
xnor U5313 (N_5313,N_5126,N_5028);
nor U5314 (N_5314,N_5103,N_5240);
or U5315 (N_5315,N_5096,N_5093);
nor U5316 (N_5316,N_5086,N_5094);
xor U5317 (N_5317,N_5005,N_5055);
xor U5318 (N_5318,N_5061,N_5242);
or U5319 (N_5319,N_5037,N_5173);
nor U5320 (N_5320,N_5142,N_5087);
nand U5321 (N_5321,N_5111,N_5014);
nor U5322 (N_5322,N_5237,N_5106);
nor U5323 (N_5323,N_5194,N_5020);
xor U5324 (N_5324,N_5224,N_5044);
or U5325 (N_5325,N_5107,N_5207);
nor U5326 (N_5326,N_5069,N_5079);
xnor U5327 (N_5327,N_5004,N_5217);
and U5328 (N_5328,N_5223,N_5025);
nor U5329 (N_5329,N_5133,N_5136);
nand U5330 (N_5330,N_5015,N_5099);
nand U5331 (N_5331,N_5059,N_5140);
or U5332 (N_5332,N_5134,N_5046);
xnor U5333 (N_5333,N_5075,N_5243);
and U5334 (N_5334,N_5013,N_5146);
xnor U5335 (N_5335,N_5123,N_5064);
nor U5336 (N_5336,N_5238,N_5026);
or U5337 (N_5337,N_5023,N_5170);
xnor U5338 (N_5338,N_5151,N_5179);
xor U5339 (N_5339,N_5051,N_5233);
and U5340 (N_5340,N_5101,N_5022);
xnor U5341 (N_5341,N_5150,N_5032);
and U5342 (N_5342,N_5222,N_5189);
nor U5343 (N_5343,N_5167,N_5110);
and U5344 (N_5344,N_5226,N_5185);
or U5345 (N_5345,N_5211,N_5100);
nand U5346 (N_5346,N_5047,N_5078);
and U5347 (N_5347,N_5166,N_5017);
nor U5348 (N_5348,N_5081,N_5158);
nor U5349 (N_5349,N_5155,N_5232);
nor U5350 (N_5350,N_5131,N_5001);
xor U5351 (N_5351,N_5198,N_5157);
or U5352 (N_5352,N_5089,N_5192);
nor U5353 (N_5353,N_5083,N_5018);
or U5354 (N_5354,N_5228,N_5006);
nand U5355 (N_5355,N_5215,N_5085);
or U5356 (N_5356,N_5021,N_5227);
nand U5357 (N_5357,N_5073,N_5139);
nor U5358 (N_5358,N_5000,N_5186);
xor U5359 (N_5359,N_5156,N_5168);
and U5360 (N_5360,N_5161,N_5178);
xnor U5361 (N_5361,N_5114,N_5247);
and U5362 (N_5362,N_5201,N_5212);
and U5363 (N_5363,N_5062,N_5027);
or U5364 (N_5364,N_5056,N_5246);
nand U5365 (N_5365,N_5160,N_5036);
nor U5366 (N_5366,N_5241,N_5206);
xnor U5367 (N_5367,N_5172,N_5248);
xnor U5368 (N_5368,N_5019,N_5080);
or U5369 (N_5369,N_5235,N_5175);
and U5370 (N_5370,N_5225,N_5199);
and U5371 (N_5371,N_5130,N_5181);
nor U5372 (N_5372,N_5209,N_5122);
xnor U5373 (N_5373,N_5097,N_5145);
nand U5374 (N_5374,N_5052,N_5230);
or U5375 (N_5375,N_5184,N_5235);
xor U5376 (N_5376,N_5052,N_5189);
nor U5377 (N_5377,N_5036,N_5229);
nand U5378 (N_5378,N_5225,N_5080);
xnor U5379 (N_5379,N_5160,N_5107);
nor U5380 (N_5380,N_5164,N_5149);
or U5381 (N_5381,N_5179,N_5019);
nand U5382 (N_5382,N_5240,N_5050);
nand U5383 (N_5383,N_5200,N_5111);
nand U5384 (N_5384,N_5113,N_5050);
or U5385 (N_5385,N_5225,N_5147);
or U5386 (N_5386,N_5033,N_5042);
or U5387 (N_5387,N_5017,N_5149);
xor U5388 (N_5388,N_5076,N_5101);
and U5389 (N_5389,N_5021,N_5012);
nor U5390 (N_5390,N_5081,N_5163);
nand U5391 (N_5391,N_5190,N_5087);
xor U5392 (N_5392,N_5237,N_5061);
xor U5393 (N_5393,N_5127,N_5170);
and U5394 (N_5394,N_5151,N_5131);
nor U5395 (N_5395,N_5203,N_5128);
and U5396 (N_5396,N_5056,N_5182);
or U5397 (N_5397,N_5155,N_5115);
nor U5398 (N_5398,N_5161,N_5019);
xnor U5399 (N_5399,N_5133,N_5058);
nor U5400 (N_5400,N_5164,N_5165);
or U5401 (N_5401,N_5041,N_5014);
or U5402 (N_5402,N_5094,N_5164);
nand U5403 (N_5403,N_5082,N_5229);
xnor U5404 (N_5404,N_5221,N_5145);
or U5405 (N_5405,N_5204,N_5065);
xnor U5406 (N_5406,N_5212,N_5041);
or U5407 (N_5407,N_5022,N_5060);
and U5408 (N_5408,N_5003,N_5101);
or U5409 (N_5409,N_5097,N_5001);
nand U5410 (N_5410,N_5181,N_5031);
nor U5411 (N_5411,N_5050,N_5197);
and U5412 (N_5412,N_5225,N_5236);
xor U5413 (N_5413,N_5249,N_5009);
nor U5414 (N_5414,N_5136,N_5101);
nand U5415 (N_5415,N_5098,N_5130);
nor U5416 (N_5416,N_5078,N_5155);
or U5417 (N_5417,N_5053,N_5025);
xnor U5418 (N_5418,N_5048,N_5196);
or U5419 (N_5419,N_5082,N_5043);
and U5420 (N_5420,N_5120,N_5177);
or U5421 (N_5421,N_5008,N_5043);
or U5422 (N_5422,N_5022,N_5102);
nor U5423 (N_5423,N_5244,N_5082);
and U5424 (N_5424,N_5207,N_5066);
nor U5425 (N_5425,N_5141,N_5088);
xor U5426 (N_5426,N_5019,N_5143);
nor U5427 (N_5427,N_5062,N_5092);
nor U5428 (N_5428,N_5005,N_5200);
or U5429 (N_5429,N_5105,N_5121);
or U5430 (N_5430,N_5041,N_5214);
and U5431 (N_5431,N_5063,N_5070);
xnor U5432 (N_5432,N_5239,N_5064);
or U5433 (N_5433,N_5068,N_5197);
xor U5434 (N_5434,N_5005,N_5182);
nor U5435 (N_5435,N_5188,N_5156);
nand U5436 (N_5436,N_5098,N_5113);
and U5437 (N_5437,N_5125,N_5075);
nand U5438 (N_5438,N_5161,N_5226);
nand U5439 (N_5439,N_5009,N_5161);
or U5440 (N_5440,N_5201,N_5023);
xnor U5441 (N_5441,N_5012,N_5025);
or U5442 (N_5442,N_5012,N_5043);
or U5443 (N_5443,N_5019,N_5243);
xor U5444 (N_5444,N_5189,N_5011);
xnor U5445 (N_5445,N_5098,N_5239);
nor U5446 (N_5446,N_5095,N_5211);
and U5447 (N_5447,N_5160,N_5219);
or U5448 (N_5448,N_5130,N_5089);
or U5449 (N_5449,N_5184,N_5174);
and U5450 (N_5450,N_5207,N_5181);
nand U5451 (N_5451,N_5028,N_5069);
xnor U5452 (N_5452,N_5166,N_5164);
nand U5453 (N_5453,N_5104,N_5076);
nor U5454 (N_5454,N_5108,N_5102);
or U5455 (N_5455,N_5073,N_5161);
nor U5456 (N_5456,N_5196,N_5071);
or U5457 (N_5457,N_5223,N_5058);
nor U5458 (N_5458,N_5112,N_5148);
nor U5459 (N_5459,N_5007,N_5065);
and U5460 (N_5460,N_5050,N_5120);
nand U5461 (N_5461,N_5005,N_5164);
nor U5462 (N_5462,N_5139,N_5230);
nor U5463 (N_5463,N_5141,N_5122);
or U5464 (N_5464,N_5198,N_5091);
nor U5465 (N_5465,N_5109,N_5050);
nand U5466 (N_5466,N_5075,N_5111);
and U5467 (N_5467,N_5057,N_5164);
nand U5468 (N_5468,N_5158,N_5050);
nor U5469 (N_5469,N_5241,N_5233);
nor U5470 (N_5470,N_5112,N_5091);
or U5471 (N_5471,N_5131,N_5104);
nand U5472 (N_5472,N_5127,N_5084);
or U5473 (N_5473,N_5194,N_5004);
nand U5474 (N_5474,N_5238,N_5130);
nor U5475 (N_5475,N_5246,N_5177);
nand U5476 (N_5476,N_5196,N_5018);
nand U5477 (N_5477,N_5099,N_5070);
nor U5478 (N_5478,N_5041,N_5104);
nor U5479 (N_5479,N_5130,N_5204);
nor U5480 (N_5480,N_5219,N_5094);
nor U5481 (N_5481,N_5140,N_5029);
or U5482 (N_5482,N_5043,N_5173);
xor U5483 (N_5483,N_5051,N_5124);
xor U5484 (N_5484,N_5118,N_5150);
nor U5485 (N_5485,N_5037,N_5002);
xor U5486 (N_5486,N_5150,N_5123);
and U5487 (N_5487,N_5021,N_5210);
nand U5488 (N_5488,N_5159,N_5245);
nand U5489 (N_5489,N_5237,N_5143);
and U5490 (N_5490,N_5208,N_5085);
or U5491 (N_5491,N_5024,N_5199);
nor U5492 (N_5492,N_5106,N_5188);
nor U5493 (N_5493,N_5226,N_5114);
or U5494 (N_5494,N_5131,N_5164);
or U5495 (N_5495,N_5071,N_5007);
nand U5496 (N_5496,N_5141,N_5225);
or U5497 (N_5497,N_5076,N_5018);
nand U5498 (N_5498,N_5223,N_5009);
xnor U5499 (N_5499,N_5039,N_5075);
or U5500 (N_5500,N_5477,N_5324);
and U5501 (N_5501,N_5437,N_5455);
or U5502 (N_5502,N_5446,N_5436);
xnor U5503 (N_5503,N_5448,N_5475);
nand U5504 (N_5504,N_5325,N_5354);
nor U5505 (N_5505,N_5495,N_5252);
xnor U5506 (N_5506,N_5385,N_5388);
and U5507 (N_5507,N_5331,N_5463);
xor U5508 (N_5508,N_5292,N_5397);
and U5509 (N_5509,N_5360,N_5444);
and U5510 (N_5510,N_5330,N_5284);
nor U5511 (N_5511,N_5470,N_5412);
nand U5512 (N_5512,N_5425,N_5409);
nor U5513 (N_5513,N_5350,N_5415);
and U5514 (N_5514,N_5469,N_5420);
nor U5515 (N_5515,N_5458,N_5499);
xor U5516 (N_5516,N_5306,N_5307);
and U5517 (N_5517,N_5456,N_5473);
or U5518 (N_5518,N_5366,N_5402);
or U5519 (N_5519,N_5260,N_5298);
nand U5520 (N_5520,N_5275,N_5309);
and U5521 (N_5521,N_5320,N_5438);
nand U5522 (N_5522,N_5404,N_5440);
and U5523 (N_5523,N_5382,N_5291);
xor U5524 (N_5524,N_5497,N_5261);
and U5525 (N_5525,N_5459,N_5482);
nand U5526 (N_5526,N_5336,N_5422);
nand U5527 (N_5527,N_5457,N_5266);
or U5528 (N_5528,N_5483,N_5281);
nor U5529 (N_5529,N_5351,N_5341);
and U5530 (N_5530,N_5478,N_5451);
and U5531 (N_5531,N_5429,N_5370);
nor U5532 (N_5532,N_5305,N_5272);
xor U5533 (N_5533,N_5380,N_5255);
or U5534 (N_5534,N_5289,N_5340);
nor U5535 (N_5535,N_5383,N_5296);
and U5536 (N_5536,N_5399,N_5349);
nand U5537 (N_5537,N_5373,N_5405);
and U5538 (N_5538,N_5427,N_5445);
nand U5539 (N_5539,N_5271,N_5277);
xnor U5540 (N_5540,N_5267,N_5329);
xnor U5541 (N_5541,N_5335,N_5414);
nand U5542 (N_5542,N_5279,N_5356);
xnor U5543 (N_5543,N_5361,N_5268);
xor U5544 (N_5544,N_5264,N_5315);
xnor U5545 (N_5545,N_5491,N_5471);
or U5546 (N_5546,N_5359,N_5316);
or U5547 (N_5547,N_5398,N_5485);
xor U5548 (N_5548,N_5406,N_5371);
nor U5549 (N_5549,N_5490,N_5396);
xor U5550 (N_5550,N_5435,N_5318);
xor U5551 (N_5551,N_5390,N_5269);
xnor U5552 (N_5552,N_5297,N_5428);
or U5553 (N_5553,N_5375,N_5358);
xnor U5554 (N_5554,N_5481,N_5327);
and U5555 (N_5555,N_5374,N_5265);
and U5556 (N_5556,N_5465,N_5372);
or U5557 (N_5557,N_5299,N_5353);
nor U5558 (N_5558,N_5301,N_5344);
and U5559 (N_5559,N_5496,N_5466);
or U5560 (N_5560,N_5310,N_5274);
and U5561 (N_5561,N_5300,N_5401);
or U5562 (N_5562,N_5431,N_5439);
nand U5563 (N_5563,N_5312,N_5416);
nand U5564 (N_5564,N_5294,N_5408);
nor U5565 (N_5565,N_5355,N_5326);
nand U5566 (N_5566,N_5413,N_5257);
nor U5567 (N_5567,N_5258,N_5494);
or U5568 (N_5568,N_5394,N_5433);
nand U5569 (N_5569,N_5389,N_5430);
or U5570 (N_5570,N_5262,N_5313);
or U5571 (N_5571,N_5323,N_5450);
nor U5572 (N_5572,N_5407,N_5319);
nor U5573 (N_5573,N_5410,N_5311);
xnor U5574 (N_5574,N_5345,N_5282);
xnor U5575 (N_5575,N_5391,N_5449);
nor U5576 (N_5576,N_5302,N_5256);
nor U5577 (N_5577,N_5259,N_5461);
xnor U5578 (N_5578,N_5280,N_5387);
xor U5579 (N_5579,N_5286,N_5432);
xnor U5580 (N_5580,N_5308,N_5443);
and U5581 (N_5581,N_5453,N_5474);
nor U5582 (N_5582,N_5270,N_5334);
nand U5583 (N_5583,N_5348,N_5283);
nor U5584 (N_5584,N_5418,N_5488);
or U5585 (N_5585,N_5338,N_5304);
nor U5586 (N_5586,N_5369,N_5480);
xnor U5587 (N_5587,N_5314,N_5384);
and U5588 (N_5588,N_5303,N_5273);
or U5589 (N_5589,N_5454,N_5346);
nor U5590 (N_5590,N_5484,N_5364);
or U5591 (N_5591,N_5343,N_5426);
nor U5592 (N_5592,N_5288,N_5357);
xor U5593 (N_5593,N_5487,N_5476);
nor U5594 (N_5594,N_5339,N_5347);
nand U5595 (N_5595,N_5368,N_5492);
and U5596 (N_5596,N_5251,N_5276);
nor U5597 (N_5597,N_5250,N_5498);
or U5598 (N_5598,N_5419,N_5376);
and U5599 (N_5599,N_5278,N_5442);
nand U5600 (N_5600,N_5393,N_5253);
and U5601 (N_5601,N_5287,N_5333);
nand U5602 (N_5602,N_5467,N_5321);
and U5603 (N_5603,N_5293,N_5452);
xnor U5604 (N_5604,N_5460,N_5434);
nor U5605 (N_5605,N_5411,N_5365);
xor U5606 (N_5606,N_5379,N_5441);
xnor U5607 (N_5607,N_5421,N_5486);
and U5608 (N_5608,N_5337,N_5493);
nor U5609 (N_5609,N_5395,N_5479);
nor U5610 (N_5610,N_5285,N_5392);
nand U5611 (N_5611,N_5462,N_5362);
or U5612 (N_5612,N_5489,N_5447);
nand U5613 (N_5613,N_5377,N_5381);
nor U5614 (N_5614,N_5263,N_5386);
or U5615 (N_5615,N_5317,N_5328);
nor U5616 (N_5616,N_5403,N_5417);
and U5617 (N_5617,N_5472,N_5332);
nor U5618 (N_5618,N_5352,N_5290);
or U5619 (N_5619,N_5464,N_5423);
nand U5620 (N_5620,N_5378,N_5363);
xor U5621 (N_5621,N_5342,N_5400);
or U5622 (N_5622,N_5424,N_5322);
xor U5623 (N_5623,N_5295,N_5367);
nand U5624 (N_5624,N_5468,N_5254);
xor U5625 (N_5625,N_5344,N_5363);
xor U5626 (N_5626,N_5471,N_5255);
or U5627 (N_5627,N_5273,N_5492);
and U5628 (N_5628,N_5288,N_5499);
and U5629 (N_5629,N_5382,N_5498);
and U5630 (N_5630,N_5420,N_5334);
nand U5631 (N_5631,N_5449,N_5281);
and U5632 (N_5632,N_5390,N_5303);
xnor U5633 (N_5633,N_5299,N_5282);
nand U5634 (N_5634,N_5404,N_5340);
nor U5635 (N_5635,N_5467,N_5336);
or U5636 (N_5636,N_5437,N_5429);
xor U5637 (N_5637,N_5281,N_5330);
and U5638 (N_5638,N_5303,N_5350);
nand U5639 (N_5639,N_5494,N_5295);
and U5640 (N_5640,N_5298,N_5276);
or U5641 (N_5641,N_5252,N_5449);
nor U5642 (N_5642,N_5323,N_5253);
and U5643 (N_5643,N_5473,N_5396);
nand U5644 (N_5644,N_5307,N_5486);
nor U5645 (N_5645,N_5403,N_5343);
nand U5646 (N_5646,N_5305,N_5389);
and U5647 (N_5647,N_5456,N_5488);
nor U5648 (N_5648,N_5273,N_5293);
xnor U5649 (N_5649,N_5339,N_5252);
and U5650 (N_5650,N_5483,N_5379);
and U5651 (N_5651,N_5431,N_5466);
nor U5652 (N_5652,N_5303,N_5484);
nor U5653 (N_5653,N_5427,N_5323);
xor U5654 (N_5654,N_5390,N_5477);
nand U5655 (N_5655,N_5304,N_5413);
nand U5656 (N_5656,N_5353,N_5293);
xnor U5657 (N_5657,N_5471,N_5476);
nand U5658 (N_5658,N_5292,N_5375);
xor U5659 (N_5659,N_5427,N_5482);
or U5660 (N_5660,N_5411,N_5495);
xor U5661 (N_5661,N_5259,N_5429);
nor U5662 (N_5662,N_5255,N_5297);
nor U5663 (N_5663,N_5371,N_5280);
or U5664 (N_5664,N_5255,N_5450);
nor U5665 (N_5665,N_5439,N_5461);
nand U5666 (N_5666,N_5312,N_5485);
nand U5667 (N_5667,N_5352,N_5303);
nor U5668 (N_5668,N_5436,N_5275);
nand U5669 (N_5669,N_5388,N_5368);
nand U5670 (N_5670,N_5404,N_5438);
nand U5671 (N_5671,N_5407,N_5408);
and U5672 (N_5672,N_5379,N_5473);
and U5673 (N_5673,N_5299,N_5260);
or U5674 (N_5674,N_5275,N_5415);
and U5675 (N_5675,N_5382,N_5451);
nor U5676 (N_5676,N_5319,N_5451);
or U5677 (N_5677,N_5334,N_5351);
or U5678 (N_5678,N_5371,N_5384);
nand U5679 (N_5679,N_5371,N_5253);
and U5680 (N_5680,N_5415,N_5363);
xnor U5681 (N_5681,N_5415,N_5408);
and U5682 (N_5682,N_5284,N_5294);
xnor U5683 (N_5683,N_5335,N_5419);
nand U5684 (N_5684,N_5270,N_5493);
and U5685 (N_5685,N_5392,N_5425);
xnor U5686 (N_5686,N_5418,N_5378);
or U5687 (N_5687,N_5481,N_5316);
nor U5688 (N_5688,N_5336,N_5461);
and U5689 (N_5689,N_5427,N_5292);
nand U5690 (N_5690,N_5317,N_5292);
nor U5691 (N_5691,N_5467,N_5353);
nor U5692 (N_5692,N_5419,N_5308);
and U5693 (N_5693,N_5273,N_5338);
or U5694 (N_5694,N_5349,N_5494);
or U5695 (N_5695,N_5339,N_5482);
xnor U5696 (N_5696,N_5404,N_5469);
nand U5697 (N_5697,N_5445,N_5367);
and U5698 (N_5698,N_5396,N_5268);
nor U5699 (N_5699,N_5350,N_5318);
xnor U5700 (N_5700,N_5424,N_5457);
nor U5701 (N_5701,N_5392,N_5368);
and U5702 (N_5702,N_5323,N_5255);
xor U5703 (N_5703,N_5338,N_5475);
nor U5704 (N_5704,N_5428,N_5262);
xnor U5705 (N_5705,N_5486,N_5303);
nor U5706 (N_5706,N_5444,N_5338);
and U5707 (N_5707,N_5323,N_5343);
xnor U5708 (N_5708,N_5486,N_5375);
nand U5709 (N_5709,N_5347,N_5359);
nand U5710 (N_5710,N_5327,N_5316);
nand U5711 (N_5711,N_5395,N_5373);
nand U5712 (N_5712,N_5306,N_5379);
or U5713 (N_5713,N_5446,N_5465);
nand U5714 (N_5714,N_5377,N_5322);
nor U5715 (N_5715,N_5374,N_5455);
or U5716 (N_5716,N_5309,N_5260);
or U5717 (N_5717,N_5440,N_5268);
nand U5718 (N_5718,N_5253,N_5276);
nor U5719 (N_5719,N_5361,N_5313);
xnor U5720 (N_5720,N_5412,N_5293);
or U5721 (N_5721,N_5290,N_5299);
and U5722 (N_5722,N_5373,N_5379);
nand U5723 (N_5723,N_5427,N_5306);
xnor U5724 (N_5724,N_5344,N_5469);
or U5725 (N_5725,N_5298,N_5458);
and U5726 (N_5726,N_5279,N_5476);
nor U5727 (N_5727,N_5294,N_5298);
and U5728 (N_5728,N_5497,N_5278);
or U5729 (N_5729,N_5273,N_5451);
and U5730 (N_5730,N_5456,N_5326);
or U5731 (N_5731,N_5333,N_5395);
nand U5732 (N_5732,N_5377,N_5481);
or U5733 (N_5733,N_5483,N_5297);
xor U5734 (N_5734,N_5355,N_5270);
and U5735 (N_5735,N_5422,N_5475);
and U5736 (N_5736,N_5299,N_5432);
and U5737 (N_5737,N_5417,N_5311);
xor U5738 (N_5738,N_5441,N_5292);
xnor U5739 (N_5739,N_5292,N_5350);
and U5740 (N_5740,N_5357,N_5458);
nand U5741 (N_5741,N_5285,N_5327);
nor U5742 (N_5742,N_5482,N_5380);
xor U5743 (N_5743,N_5291,N_5471);
and U5744 (N_5744,N_5499,N_5349);
nor U5745 (N_5745,N_5266,N_5474);
nor U5746 (N_5746,N_5313,N_5319);
nor U5747 (N_5747,N_5379,N_5270);
nor U5748 (N_5748,N_5310,N_5497);
and U5749 (N_5749,N_5381,N_5419);
nor U5750 (N_5750,N_5614,N_5507);
nand U5751 (N_5751,N_5715,N_5730);
nand U5752 (N_5752,N_5585,N_5688);
xnor U5753 (N_5753,N_5699,N_5618);
and U5754 (N_5754,N_5616,N_5552);
and U5755 (N_5755,N_5529,N_5500);
or U5756 (N_5756,N_5728,N_5667);
xnor U5757 (N_5757,N_5632,N_5747);
nand U5758 (N_5758,N_5621,N_5726);
or U5759 (N_5759,N_5735,N_5740);
xor U5760 (N_5760,N_5707,N_5564);
and U5761 (N_5761,N_5603,N_5530);
nor U5762 (N_5762,N_5695,N_5681);
nor U5763 (N_5763,N_5521,N_5648);
xor U5764 (N_5764,N_5544,N_5703);
nor U5765 (N_5765,N_5506,N_5636);
nor U5766 (N_5766,N_5567,N_5508);
and U5767 (N_5767,N_5609,N_5556);
and U5768 (N_5768,N_5612,N_5718);
nor U5769 (N_5769,N_5732,N_5587);
nand U5770 (N_5770,N_5599,N_5663);
xor U5771 (N_5771,N_5731,N_5572);
and U5772 (N_5772,N_5687,N_5694);
and U5773 (N_5773,N_5590,N_5619);
or U5774 (N_5774,N_5719,N_5513);
nor U5775 (N_5775,N_5535,N_5576);
nand U5776 (N_5776,N_5725,N_5607);
xor U5777 (N_5777,N_5524,N_5601);
or U5778 (N_5778,N_5597,N_5611);
nand U5779 (N_5779,N_5657,N_5701);
and U5780 (N_5780,N_5720,N_5671);
or U5781 (N_5781,N_5678,N_5656);
xor U5782 (N_5782,N_5709,N_5668);
and U5783 (N_5783,N_5538,N_5693);
or U5784 (N_5784,N_5654,N_5596);
or U5785 (N_5785,N_5634,N_5515);
nor U5786 (N_5786,N_5736,N_5637);
xor U5787 (N_5787,N_5723,N_5630);
xnor U5788 (N_5788,N_5631,N_5729);
and U5789 (N_5789,N_5600,N_5662);
and U5790 (N_5790,N_5595,N_5744);
xor U5791 (N_5791,N_5531,N_5604);
or U5792 (N_5792,N_5745,N_5652);
nand U5793 (N_5793,N_5643,N_5617);
nand U5794 (N_5794,N_5738,N_5522);
xor U5795 (N_5795,N_5639,N_5545);
nand U5796 (N_5796,N_5650,N_5503);
nor U5797 (N_5797,N_5742,N_5642);
xnor U5798 (N_5798,N_5537,N_5660);
xor U5799 (N_5799,N_5582,N_5565);
or U5800 (N_5800,N_5581,N_5669);
nand U5801 (N_5801,N_5505,N_5541);
or U5802 (N_5802,N_5605,N_5633);
nor U5803 (N_5803,N_5525,N_5689);
or U5804 (N_5804,N_5584,N_5520);
and U5805 (N_5805,N_5577,N_5705);
nand U5806 (N_5806,N_5638,N_5655);
nor U5807 (N_5807,N_5504,N_5517);
nor U5808 (N_5808,N_5547,N_5511);
nor U5809 (N_5809,N_5592,N_5641);
or U5810 (N_5810,N_5615,N_5749);
or U5811 (N_5811,N_5574,N_5571);
nand U5812 (N_5812,N_5627,N_5519);
and U5813 (N_5813,N_5583,N_5536);
or U5814 (N_5814,N_5651,N_5661);
xor U5815 (N_5815,N_5665,N_5512);
xnor U5816 (N_5816,N_5549,N_5546);
nor U5817 (N_5817,N_5708,N_5640);
nand U5818 (N_5818,N_5670,N_5573);
or U5819 (N_5819,N_5673,N_5591);
nand U5820 (N_5820,N_5598,N_5684);
xnor U5821 (N_5821,N_5739,N_5575);
nand U5822 (N_5822,N_5686,N_5721);
and U5823 (N_5823,N_5653,N_5586);
or U5824 (N_5824,N_5716,N_5727);
nor U5825 (N_5825,N_5722,N_5620);
and U5826 (N_5826,N_5624,N_5626);
and U5827 (N_5827,N_5579,N_5548);
nor U5828 (N_5828,N_5613,N_5717);
xnor U5829 (N_5829,N_5691,N_5558);
nand U5830 (N_5830,N_5706,N_5683);
and U5831 (N_5831,N_5589,N_5610);
and U5832 (N_5832,N_5578,N_5623);
nor U5833 (N_5833,N_5674,N_5569);
nor U5834 (N_5834,N_5690,N_5676);
and U5835 (N_5835,N_5711,N_5542);
or U5836 (N_5836,N_5550,N_5704);
xnor U5837 (N_5837,N_5555,N_5514);
xor U5838 (N_5838,N_5509,N_5724);
nor U5839 (N_5839,N_5562,N_5635);
nand U5840 (N_5840,N_5527,N_5646);
and U5841 (N_5841,N_5734,N_5710);
xnor U5842 (N_5842,N_5680,N_5560);
nand U5843 (N_5843,N_5672,N_5528);
or U5844 (N_5844,N_5554,N_5679);
and U5845 (N_5845,N_5534,N_5602);
nand U5846 (N_5846,N_5553,N_5645);
nor U5847 (N_5847,N_5593,N_5733);
and U5848 (N_5848,N_5682,N_5563);
and U5849 (N_5849,N_5628,N_5606);
nand U5850 (N_5850,N_5659,N_5714);
nor U5851 (N_5851,N_5644,N_5737);
nor U5852 (N_5852,N_5570,N_5700);
and U5853 (N_5853,N_5746,N_5685);
nand U5854 (N_5854,N_5666,N_5518);
or U5855 (N_5855,N_5696,N_5741);
nor U5856 (N_5856,N_5539,N_5625);
nor U5857 (N_5857,N_5523,N_5677);
xnor U5858 (N_5858,N_5629,N_5551);
nor U5859 (N_5859,N_5580,N_5649);
xor U5860 (N_5860,N_5568,N_5697);
or U5861 (N_5861,N_5561,N_5540);
and U5862 (N_5862,N_5658,N_5510);
nor U5863 (N_5863,N_5526,N_5559);
and U5864 (N_5864,N_5557,N_5543);
xnor U5865 (N_5865,N_5532,N_5675);
xor U5866 (N_5866,N_5743,N_5713);
and U5867 (N_5867,N_5692,N_5501);
xor U5868 (N_5868,N_5588,N_5533);
and U5869 (N_5869,N_5702,N_5594);
xor U5870 (N_5870,N_5698,N_5748);
and U5871 (N_5871,N_5664,N_5647);
nand U5872 (N_5872,N_5712,N_5516);
and U5873 (N_5873,N_5622,N_5502);
xnor U5874 (N_5874,N_5608,N_5566);
xor U5875 (N_5875,N_5592,N_5506);
or U5876 (N_5876,N_5566,N_5518);
nand U5877 (N_5877,N_5705,N_5666);
and U5878 (N_5878,N_5535,N_5680);
or U5879 (N_5879,N_5544,N_5546);
or U5880 (N_5880,N_5621,N_5557);
or U5881 (N_5881,N_5644,N_5505);
nor U5882 (N_5882,N_5675,N_5533);
xor U5883 (N_5883,N_5602,N_5594);
or U5884 (N_5884,N_5632,N_5645);
nand U5885 (N_5885,N_5520,N_5602);
and U5886 (N_5886,N_5633,N_5662);
or U5887 (N_5887,N_5739,N_5619);
nor U5888 (N_5888,N_5628,N_5572);
xnor U5889 (N_5889,N_5697,N_5631);
or U5890 (N_5890,N_5585,N_5563);
or U5891 (N_5891,N_5534,N_5681);
or U5892 (N_5892,N_5711,N_5668);
or U5893 (N_5893,N_5663,N_5725);
nor U5894 (N_5894,N_5507,N_5657);
xor U5895 (N_5895,N_5639,N_5578);
xnor U5896 (N_5896,N_5603,N_5647);
xnor U5897 (N_5897,N_5694,N_5643);
and U5898 (N_5898,N_5743,N_5640);
or U5899 (N_5899,N_5590,N_5613);
nor U5900 (N_5900,N_5739,N_5704);
xnor U5901 (N_5901,N_5701,N_5552);
nand U5902 (N_5902,N_5686,N_5633);
or U5903 (N_5903,N_5668,N_5740);
xnor U5904 (N_5904,N_5629,N_5678);
nand U5905 (N_5905,N_5587,N_5531);
or U5906 (N_5906,N_5737,N_5514);
xor U5907 (N_5907,N_5636,N_5690);
nand U5908 (N_5908,N_5639,N_5643);
nor U5909 (N_5909,N_5677,N_5749);
nor U5910 (N_5910,N_5692,N_5657);
or U5911 (N_5911,N_5700,N_5522);
nand U5912 (N_5912,N_5673,N_5706);
nand U5913 (N_5913,N_5569,N_5646);
and U5914 (N_5914,N_5523,N_5555);
nor U5915 (N_5915,N_5579,N_5635);
and U5916 (N_5916,N_5696,N_5714);
nand U5917 (N_5917,N_5678,N_5615);
nor U5918 (N_5918,N_5599,N_5575);
and U5919 (N_5919,N_5708,N_5619);
and U5920 (N_5920,N_5666,N_5641);
xnor U5921 (N_5921,N_5624,N_5639);
xnor U5922 (N_5922,N_5520,N_5653);
nor U5923 (N_5923,N_5724,N_5744);
nand U5924 (N_5924,N_5622,N_5544);
nor U5925 (N_5925,N_5533,N_5706);
nand U5926 (N_5926,N_5685,N_5666);
or U5927 (N_5927,N_5667,N_5632);
or U5928 (N_5928,N_5545,N_5686);
nand U5929 (N_5929,N_5616,N_5670);
nor U5930 (N_5930,N_5580,N_5696);
nand U5931 (N_5931,N_5613,N_5661);
nor U5932 (N_5932,N_5696,N_5726);
and U5933 (N_5933,N_5530,N_5648);
nand U5934 (N_5934,N_5586,N_5610);
and U5935 (N_5935,N_5664,N_5726);
and U5936 (N_5936,N_5671,N_5577);
nor U5937 (N_5937,N_5719,N_5645);
xor U5938 (N_5938,N_5611,N_5701);
nand U5939 (N_5939,N_5679,N_5715);
and U5940 (N_5940,N_5709,N_5632);
or U5941 (N_5941,N_5703,N_5678);
or U5942 (N_5942,N_5672,N_5652);
or U5943 (N_5943,N_5643,N_5714);
xnor U5944 (N_5944,N_5733,N_5725);
and U5945 (N_5945,N_5546,N_5512);
or U5946 (N_5946,N_5625,N_5504);
or U5947 (N_5947,N_5622,N_5672);
or U5948 (N_5948,N_5571,N_5629);
nor U5949 (N_5949,N_5742,N_5605);
nor U5950 (N_5950,N_5587,N_5711);
and U5951 (N_5951,N_5591,N_5746);
or U5952 (N_5952,N_5689,N_5547);
xnor U5953 (N_5953,N_5725,N_5749);
and U5954 (N_5954,N_5517,N_5500);
and U5955 (N_5955,N_5601,N_5591);
xnor U5956 (N_5956,N_5541,N_5644);
nor U5957 (N_5957,N_5556,N_5551);
nand U5958 (N_5958,N_5611,N_5654);
nand U5959 (N_5959,N_5523,N_5698);
nand U5960 (N_5960,N_5502,N_5743);
nand U5961 (N_5961,N_5536,N_5696);
and U5962 (N_5962,N_5582,N_5636);
or U5963 (N_5963,N_5691,N_5686);
and U5964 (N_5964,N_5510,N_5645);
xor U5965 (N_5965,N_5544,N_5589);
and U5966 (N_5966,N_5624,N_5594);
nor U5967 (N_5967,N_5646,N_5708);
nor U5968 (N_5968,N_5581,N_5623);
nor U5969 (N_5969,N_5577,N_5746);
or U5970 (N_5970,N_5705,N_5538);
or U5971 (N_5971,N_5661,N_5708);
and U5972 (N_5972,N_5586,N_5702);
nand U5973 (N_5973,N_5574,N_5504);
nand U5974 (N_5974,N_5530,N_5643);
xor U5975 (N_5975,N_5581,N_5555);
or U5976 (N_5976,N_5610,N_5566);
nand U5977 (N_5977,N_5732,N_5550);
and U5978 (N_5978,N_5562,N_5720);
xor U5979 (N_5979,N_5595,N_5659);
nor U5980 (N_5980,N_5671,N_5688);
xor U5981 (N_5981,N_5733,N_5715);
nor U5982 (N_5982,N_5679,N_5671);
or U5983 (N_5983,N_5639,N_5667);
nand U5984 (N_5984,N_5591,N_5542);
xor U5985 (N_5985,N_5730,N_5623);
nor U5986 (N_5986,N_5648,N_5735);
xor U5987 (N_5987,N_5687,N_5519);
or U5988 (N_5988,N_5606,N_5694);
nor U5989 (N_5989,N_5611,N_5567);
or U5990 (N_5990,N_5579,N_5707);
nand U5991 (N_5991,N_5734,N_5544);
nand U5992 (N_5992,N_5727,N_5568);
nor U5993 (N_5993,N_5556,N_5670);
xnor U5994 (N_5994,N_5676,N_5710);
nand U5995 (N_5995,N_5655,N_5683);
and U5996 (N_5996,N_5711,N_5613);
xor U5997 (N_5997,N_5541,N_5593);
xnor U5998 (N_5998,N_5654,N_5674);
or U5999 (N_5999,N_5582,N_5607);
xnor U6000 (N_6000,N_5762,N_5770);
and U6001 (N_6001,N_5988,N_5951);
or U6002 (N_6002,N_5810,N_5923);
and U6003 (N_6003,N_5804,N_5925);
and U6004 (N_6004,N_5815,N_5877);
xor U6005 (N_6005,N_5936,N_5757);
nor U6006 (N_6006,N_5807,N_5843);
and U6007 (N_6007,N_5873,N_5968);
and U6008 (N_6008,N_5907,N_5962);
nor U6009 (N_6009,N_5880,N_5871);
or U6010 (N_6010,N_5940,N_5959);
nor U6011 (N_6011,N_5987,N_5817);
nand U6012 (N_6012,N_5809,N_5975);
nand U6013 (N_6013,N_5950,N_5759);
or U6014 (N_6014,N_5839,N_5855);
nand U6015 (N_6015,N_5902,N_5808);
nand U6016 (N_6016,N_5995,N_5969);
nor U6017 (N_6017,N_5751,N_5778);
and U6018 (N_6018,N_5961,N_5753);
or U6019 (N_6019,N_5763,N_5957);
nor U6020 (N_6020,N_5791,N_5793);
or U6021 (N_6021,N_5891,N_5909);
nand U6022 (N_6022,N_5890,N_5800);
and U6023 (N_6023,N_5780,N_5994);
and U6024 (N_6024,N_5901,N_5992);
xnor U6025 (N_6025,N_5822,N_5869);
nand U6026 (N_6026,N_5981,N_5999);
or U6027 (N_6027,N_5892,N_5856);
and U6028 (N_6028,N_5993,N_5973);
and U6029 (N_6029,N_5868,N_5953);
nand U6030 (N_6030,N_5980,N_5946);
or U6031 (N_6031,N_5990,N_5898);
xnor U6032 (N_6032,N_5797,N_5976);
and U6033 (N_6033,N_5792,N_5921);
or U6034 (N_6034,N_5790,N_5779);
or U6035 (N_6035,N_5964,N_5883);
and U6036 (N_6036,N_5966,N_5811);
or U6037 (N_6037,N_5849,N_5764);
and U6038 (N_6038,N_5806,N_5913);
or U6039 (N_6039,N_5750,N_5943);
nand U6040 (N_6040,N_5845,N_5754);
nor U6041 (N_6041,N_5899,N_5984);
and U6042 (N_6042,N_5823,N_5760);
xnor U6043 (N_6043,N_5982,N_5852);
xnor U6044 (N_6044,N_5840,N_5916);
and U6045 (N_6045,N_5863,N_5983);
or U6046 (N_6046,N_5894,N_5918);
nor U6047 (N_6047,N_5803,N_5910);
nor U6048 (N_6048,N_5875,N_5755);
nand U6049 (N_6049,N_5912,N_5908);
nor U6050 (N_6050,N_5911,N_5882);
and U6051 (N_6051,N_5853,N_5865);
nor U6052 (N_6052,N_5781,N_5816);
or U6053 (N_6053,N_5768,N_5947);
nor U6054 (N_6054,N_5932,N_5897);
nor U6055 (N_6055,N_5796,N_5783);
nor U6056 (N_6056,N_5854,N_5787);
xor U6057 (N_6057,N_5773,N_5917);
and U6058 (N_6058,N_5906,N_5812);
and U6059 (N_6059,N_5842,N_5813);
and U6060 (N_6060,N_5928,N_5884);
and U6061 (N_6061,N_5876,N_5851);
nand U6062 (N_6062,N_5881,N_5821);
nand U6063 (N_6063,N_5986,N_5978);
nand U6064 (N_6064,N_5989,N_5786);
nor U6065 (N_6065,N_5954,N_5777);
nor U6066 (N_6066,N_5915,N_5752);
xnor U6067 (N_6067,N_5788,N_5887);
xor U6068 (N_6068,N_5935,N_5971);
and U6069 (N_6069,N_5767,N_5970);
xor U6070 (N_6070,N_5857,N_5960);
xnor U6071 (N_6071,N_5920,N_5774);
or U6072 (N_6072,N_5998,N_5766);
or U6073 (N_6073,N_5772,N_5859);
and U6074 (N_6074,N_5952,N_5848);
xor U6075 (N_6075,N_5784,N_5941);
and U6076 (N_6076,N_5775,N_5942);
xnor U6077 (N_6077,N_5896,N_5867);
nor U6078 (N_6078,N_5991,N_5945);
nor U6079 (N_6079,N_5905,N_5900);
nor U6080 (N_6080,N_5885,N_5956);
or U6081 (N_6081,N_5832,N_5972);
and U6082 (N_6082,N_5829,N_5965);
and U6083 (N_6083,N_5818,N_5838);
nor U6084 (N_6084,N_5785,N_5835);
and U6085 (N_6085,N_5841,N_5776);
nand U6086 (N_6086,N_5765,N_5979);
xnor U6087 (N_6087,N_5931,N_5798);
or U6088 (N_6088,N_5864,N_5824);
and U6089 (N_6089,N_5756,N_5844);
or U6090 (N_6090,N_5828,N_5889);
nor U6091 (N_6091,N_5836,N_5888);
nand U6092 (N_6092,N_5985,N_5834);
nor U6093 (N_6093,N_5769,N_5866);
and U6094 (N_6094,N_5948,N_5929);
xnor U6095 (N_6095,N_5850,N_5831);
and U6096 (N_6096,N_5846,N_5893);
or U6097 (N_6097,N_5967,N_5878);
nand U6098 (N_6098,N_5919,N_5903);
nor U6099 (N_6099,N_5789,N_5833);
xnor U6100 (N_6100,N_5872,N_5944);
nand U6101 (N_6101,N_5933,N_5997);
xnor U6102 (N_6102,N_5904,N_5826);
nor U6103 (N_6103,N_5922,N_5949);
or U6104 (N_6104,N_5870,N_5820);
xnor U6105 (N_6105,N_5977,N_5958);
nand U6106 (N_6106,N_5782,N_5799);
and U6107 (N_6107,N_5926,N_5847);
and U6108 (N_6108,N_5837,N_5886);
and U6109 (N_6109,N_5879,N_5761);
or U6110 (N_6110,N_5862,N_5830);
and U6111 (N_6111,N_5802,N_5861);
nor U6112 (N_6112,N_5974,N_5814);
and U6113 (N_6113,N_5819,N_5794);
xnor U6114 (N_6114,N_5858,N_5874);
or U6115 (N_6115,N_5927,N_5795);
nand U6116 (N_6116,N_5771,N_5805);
and U6117 (N_6117,N_5939,N_5914);
nand U6118 (N_6118,N_5895,N_5934);
nand U6119 (N_6119,N_5937,N_5930);
and U6120 (N_6120,N_5801,N_5825);
and U6121 (N_6121,N_5758,N_5827);
or U6122 (N_6122,N_5996,N_5924);
nor U6123 (N_6123,N_5938,N_5955);
xor U6124 (N_6124,N_5963,N_5860);
nand U6125 (N_6125,N_5845,N_5866);
or U6126 (N_6126,N_5844,N_5787);
nand U6127 (N_6127,N_5938,N_5824);
and U6128 (N_6128,N_5806,N_5805);
and U6129 (N_6129,N_5928,N_5756);
xor U6130 (N_6130,N_5966,N_5937);
nor U6131 (N_6131,N_5974,N_5967);
xor U6132 (N_6132,N_5952,N_5836);
nand U6133 (N_6133,N_5792,N_5977);
xnor U6134 (N_6134,N_5966,N_5962);
or U6135 (N_6135,N_5779,N_5817);
or U6136 (N_6136,N_5952,N_5913);
nand U6137 (N_6137,N_5844,N_5870);
nor U6138 (N_6138,N_5914,N_5769);
xnor U6139 (N_6139,N_5936,N_5917);
and U6140 (N_6140,N_5946,N_5949);
xor U6141 (N_6141,N_5763,N_5970);
xnor U6142 (N_6142,N_5834,N_5804);
nor U6143 (N_6143,N_5854,N_5769);
nor U6144 (N_6144,N_5871,N_5836);
and U6145 (N_6145,N_5911,N_5761);
xnor U6146 (N_6146,N_5865,N_5840);
or U6147 (N_6147,N_5753,N_5769);
or U6148 (N_6148,N_5926,N_5840);
or U6149 (N_6149,N_5835,N_5884);
nand U6150 (N_6150,N_5813,N_5853);
or U6151 (N_6151,N_5795,N_5923);
xnor U6152 (N_6152,N_5802,N_5961);
and U6153 (N_6153,N_5958,N_5996);
nand U6154 (N_6154,N_5832,N_5964);
nor U6155 (N_6155,N_5896,N_5788);
and U6156 (N_6156,N_5817,N_5965);
or U6157 (N_6157,N_5901,N_5903);
and U6158 (N_6158,N_5766,N_5985);
or U6159 (N_6159,N_5892,N_5940);
nor U6160 (N_6160,N_5952,N_5865);
nor U6161 (N_6161,N_5894,N_5945);
xor U6162 (N_6162,N_5847,N_5860);
and U6163 (N_6163,N_5884,N_5967);
nor U6164 (N_6164,N_5977,N_5870);
or U6165 (N_6165,N_5872,N_5775);
or U6166 (N_6166,N_5894,N_5868);
nand U6167 (N_6167,N_5854,N_5966);
or U6168 (N_6168,N_5993,N_5807);
nand U6169 (N_6169,N_5778,N_5882);
and U6170 (N_6170,N_5869,N_5799);
nand U6171 (N_6171,N_5856,N_5916);
nor U6172 (N_6172,N_5854,N_5785);
or U6173 (N_6173,N_5798,N_5759);
and U6174 (N_6174,N_5860,N_5934);
or U6175 (N_6175,N_5796,N_5789);
nor U6176 (N_6176,N_5872,N_5849);
and U6177 (N_6177,N_5999,N_5812);
nor U6178 (N_6178,N_5932,N_5776);
or U6179 (N_6179,N_5783,N_5808);
nor U6180 (N_6180,N_5940,N_5824);
xor U6181 (N_6181,N_5914,N_5993);
nand U6182 (N_6182,N_5995,N_5790);
or U6183 (N_6183,N_5768,N_5828);
nand U6184 (N_6184,N_5981,N_5833);
or U6185 (N_6185,N_5996,N_5928);
xor U6186 (N_6186,N_5805,N_5899);
nand U6187 (N_6187,N_5902,N_5876);
nand U6188 (N_6188,N_5796,N_5996);
xor U6189 (N_6189,N_5940,N_5863);
and U6190 (N_6190,N_5941,N_5893);
nor U6191 (N_6191,N_5931,N_5854);
nand U6192 (N_6192,N_5880,N_5854);
or U6193 (N_6193,N_5865,N_5984);
and U6194 (N_6194,N_5927,N_5787);
and U6195 (N_6195,N_5839,N_5891);
nand U6196 (N_6196,N_5919,N_5949);
xor U6197 (N_6197,N_5901,N_5788);
nor U6198 (N_6198,N_5988,N_5784);
and U6199 (N_6199,N_5936,N_5895);
nor U6200 (N_6200,N_5797,N_5933);
xnor U6201 (N_6201,N_5912,N_5957);
nand U6202 (N_6202,N_5777,N_5791);
and U6203 (N_6203,N_5892,N_5889);
or U6204 (N_6204,N_5788,N_5954);
nor U6205 (N_6205,N_5754,N_5862);
nand U6206 (N_6206,N_5961,N_5807);
nand U6207 (N_6207,N_5986,N_5812);
nand U6208 (N_6208,N_5811,N_5885);
and U6209 (N_6209,N_5834,N_5976);
or U6210 (N_6210,N_5757,N_5931);
or U6211 (N_6211,N_5949,N_5942);
or U6212 (N_6212,N_5944,N_5954);
and U6213 (N_6213,N_5983,N_5890);
and U6214 (N_6214,N_5823,N_5958);
xor U6215 (N_6215,N_5912,N_5757);
nor U6216 (N_6216,N_5951,N_5917);
nor U6217 (N_6217,N_5872,N_5969);
xnor U6218 (N_6218,N_5942,N_5858);
or U6219 (N_6219,N_5848,N_5823);
xnor U6220 (N_6220,N_5867,N_5903);
and U6221 (N_6221,N_5977,N_5866);
or U6222 (N_6222,N_5920,N_5768);
and U6223 (N_6223,N_5779,N_5980);
nand U6224 (N_6224,N_5832,N_5846);
and U6225 (N_6225,N_5821,N_5786);
and U6226 (N_6226,N_5872,N_5837);
nand U6227 (N_6227,N_5909,N_5890);
xnor U6228 (N_6228,N_5893,N_5909);
nor U6229 (N_6229,N_5829,N_5969);
nor U6230 (N_6230,N_5870,N_5839);
or U6231 (N_6231,N_5768,N_5845);
xor U6232 (N_6232,N_5928,N_5948);
nand U6233 (N_6233,N_5902,N_5786);
and U6234 (N_6234,N_5970,N_5772);
nand U6235 (N_6235,N_5831,N_5773);
nor U6236 (N_6236,N_5915,N_5785);
and U6237 (N_6237,N_5762,N_5976);
xnor U6238 (N_6238,N_5810,N_5997);
nor U6239 (N_6239,N_5848,N_5772);
nand U6240 (N_6240,N_5861,N_5798);
or U6241 (N_6241,N_5863,N_5756);
xnor U6242 (N_6242,N_5785,N_5784);
nand U6243 (N_6243,N_5756,N_5826);
nor U6244 (N_6244,N_5835,N_5968);
and U6245 (N_6245,N_5932,N_5847);
xor U6246 (N_6246,N_5976,N_5904);
nand U6247 (N_6247,N_5770,N_5908);
xor U6248 (N_6248,N_5764,N_5813);
nand U6249 (N_6249,N_5823,N_5844);
xor U6250 (N_6250,N_6053,N_6163);
nor U6251 (N_6251,N_6031,N_6162);
xnor U6252 (N_6252,N_6043,N_6074);
and U6253 (N_6253,N_6206,N_6219);
or U6254 (N_6254,N_6100,N_6147);
or U6255 (N_6255,N_6094,N_6138);
nand U6256 (N_6256,N_6071,N_6129);
nor U6257 (N_6257,N_6196,N_6051);
or U6258 (N_6258,N_6080,N_6126);
nand U6259 (N_6259,N_6150,N_6159);
nor U6260 (N_6260,N_6110,N_6024);
and U6261 (N_6261,N_6056,N_6115);
or U6262 (N_6262,N_6021,N_6227);
nand U6263 (N_6263,N_6226,N_6148);
nor U6264 (N_6264,N_6231,N_6067);
nand U6265 (N_6265,N_6116,N_6038);
or U6266 (N_6266,N_6003,N_6045);
or U6267 (N_6267,N_6173,N_6143);
nor U6268 (N_6268,N_6125,N_6197);
and U6269 (N_6269,N_6236,N_6055);
xnor U6270 (N_6270,N_6247,N_6142);
xnor U6271 (N_6271,N_6086,N_6122);
nor U6272 (N_6272,N_6178,N_6083);
and U6273 (N_6273,N_6033,N_6213);
nor U6274 (N_6274,N_6018,N_6019);
xor U6275 (N_6275,N_6054,N_6068);
nand U6276 (N_6276,N_6104,N_6153);
nor U6277 (N_6277,N_6199,N_6154);
nand U6278 (N_6278,N_6225,N_6136);
and U6279 (N_6279,N_6022,N_6169);
nor U6280 (N_6280,N_6012,N_6088);
and U6281 (N_6281,N_6235,N_6208);
nand U6282 (N_6282,N_6157,N_6151);
or U6283 (N_6283,N_6065,N_6165);
and U6284 (N_6284,N_6202,N_6037);
xor U6285 (N_6285,N_6092,N_6158);
nand U6286 (N_6286,N_6076,N_6057);
and U6287 (N_6287,N_6204,N_6141);
or U6288 (N_6288,N_6059,N_6113);
xor U6289 (N_6289,N_6058,N_6174);
xnor U6290 (N_6290,N_6082,N_6127);
nand U6291 (N_6291,N_6052,N_6085);
nand U6292 (N_6292,N_6184,N_6069);
or U6293 (N_6293,N_6240,N_6249);
and U6294 (N_6294,N_6101,N_6133);
and U6295 (N_6295,N_6046,N_6242);
or U6296 (N_6296,N_6171,N_6026);
nand U6297 (N_6297,N_6090,N_6049);
or U6298 (N_6298,N_6042,N_6061);
xnor U6299 (N_6299,N_6060,N_6200);
nor U6300 (N_6300,N_6016,N_6216);
nor U6301 (N_6301,N_6041,N_6095);
nand U6302 (N_6302,N_6146,N_6077);
nor U6303 (N_6303,N_6089,N_6102);
and U6304 (N_6304,N_6161,N_6114);
nor U6305 (N_6305,N_6118,N_6180);
xor U6306 (N_6306,N_6215,N_6218);
and U6307 (N_6307,N_6036,N_6070);
nand U6308 (N_6308,N_6075,N_6185);
and U6309 (N_6309,N_6011,N_6097);
or U6310 (N_6310,N_6044,N_6006);
xnor U6311 (N_6311,N_6246,N_6010);
nand U6312 (N_6312,N_6189,N_6188);
and U6313 (N_6313,N_6047,N_6194);
and U6314 (N_6314,N_6005,N_6164);
and U6315 (N_6315,N_6079,N_6093);
and U6316 (N_6316,N_6008,N_6175);
nand U6317 (N_6317,N_6048,N_6029);
and U6318 (N_6318,N_6193,N_6190);
nand U6319 (N_6319,N_6000,N_6034);
or U6320 (N_6320,N_6028,N_6217);
or U6321 (N_6321,N_6062,N_6156);
xor U6322 (N_6322,N_6137,N_6063);
nand U6323 (N_6323,N_6119,N_6081);
xor U6324 (N_6324,N_6039,N_6002);
nand U6325 (N_6325,N_6120,N_6230);
and U6326 (N_6326,N_6210,N_6107);
and U6327 (N_6327,N_6084,N_6168);
or U6328 (N_6328,N_6066,N_6130);
xor U6329 (N_6329,N_6152,N_6099);
xnor U6330 (N_6330,N_6239,N_6186);
nand U6331 (N_6331,N_6244,N_6149);
nand U6332 (N_6332,N_6245,N_6198);
xnor U6333 (N_6333,N_6108,N_6243);
or U6334 (N_6334,N_6145,N_6030);
or U6335 (N_6335,N_6179,N_6167);
nand U6336 (N_6336,N_6203,N_6195);
or U6337 (N_6337,N_6035,N_6211);
and U6338 (N_6338,N_6223,N_6087);
and U6339 (N_6339,N_6182,N_6015);
nand U6340 (N_6340,N_6009,N_6160);
xor U6341 (N_6341,N_6064,N_6234);
nor U6342 (N_6342,N_6123,N_6014);
and U6343 (N_6343,N_6155,N_6212);
and U6344 (N_6344,N_6134,N_6032);
xor U6345 (N_6345,N_6105,N_6201);
and U6346 (N_6346,N_6109,N_6007);
xor U6347 (N_6347,N_6132,N_6103);
nor U6348 (N_6348,N_6248,N_6166);
xor U6349 (N_6349,N_6224,N_6020);
nor U6350 (N_6350,N_6228,N_6237);
and U6351 (N_6351,N_6004,N_6241);
or U6352 (N_6352,N_6222,N_6139);
and U6353 (N_6353,N_6181,N_6001);
xnor U6354 (N_6354,N_6025,N_6131);
or U6355 (N_6355,N_6128,N_6209);
nand U6356 (N_6356,N_6220,N_6124);
and U6357 (N_6357,N_6017,N_6117);
nand U6358 (N_6358,N_6238,N_6106);
nor U6359 (N_6359,N_6091,N_6187);
or U6360 (N_6360,N_6205,N_6027);
and U6361 (N_6361,N_6023,N_6191);
and U6362 (N_6362,N_6013,N_6111);
or U6363 (N_6363,N_6232,N_6073);
xnor U6364 (N_6364,N_6221,N_6192);
nor U6365 (N_6365,N_6207,N_6172);
or U6366 (N_6366,N_6098,N_6233);
or U6367 (N_6367,N_6050,N_6072);
or U6368 (N_6368,N_6078,N_6176);
xnor U6369 (N_6369,N_6140,N_6040);
nor U6370 (N_6370,N_6177,N_6135);
or U6371 (N_6371,N_6170,N_6229);
xor U6372 (N_6372,N_6144,N_6121);
nand U6373 (N_6373,N_6112,N_6096);
xnor U6374 (N_6374,N_6214,N_6183);
and U6375 (N_6375,N_6046,N_6021);
nor U6376 (N_6376,N_6134,N_6131);
or U6377 (N_6377,N_6187,N_6119);
nand U6378 (N_6378,N_6131,N_6021);
or U6379 (N_6379,N_6056,N_6055);
xnor U6380 (N_6380,N_6128,N_6078);
and U6381 (N_6381,N_6239,N_6222);
nand U6382 (N_6382,N_6014,N_6033);
xor U6383 (N_6383,N_6220,N_6048);
and U6384 (N_6384,N_6092,N_6007);
or U6385 (N_6385,N_6180,N_6187);
nand U6386 (N_6386,N_6119,N_6178);
and U6387 (N_6387,N_6138,N_6111);
nand U6388 (N_6388,N_6010,N_6134);
nor U6389 (N_6389,N_6090,N_6054);
xnor U6390 (N_6390,N_6164,N_6230);
nand U6391 (N_6391,N_6084,N_6026);
and U6392 (N_6392,N_6025,N_6220);
nor U6393 (N_6393,N_6229,N_6039);
nor U6394 (N_6394,N_6239,N_6195);
nand U6395 (N_6395,N_6097,N_6137);
xor U6396 (N_6396,N_6229,N_6038);
xor U6397 (N_6397,N_6200,N_6175);
or U6398 (N_6398,N_6118,N_6155);
nand U6399 (N_6399,N_6216,N_6178);
xor U6400 (N_6400,N_6062,N_6052);
and U6401 (N_6401,N_6114,N_6043);
or U6402 (N_6402,N_6107,N_6155);
or U6403 (N_6403,N_6107,N_6078);
and U6404 (N_6404,N_6138,N_6183);
nor U6405 (N_6405,N_6151,N_6225);
nand U6406 (N_6406,N_6024,N_6002);
nor U6407 (N_6407,N_6170,N_6091);
or U6408 (N_6408,N_6196,N_6179);
and U6409 (N_6409,N_6039,N_6067);
or U6410 (N_6410,N_6065,N_6131);
nor U6411 (N_6411,N_6066,N_6222);
nor U6412 (N_6412,N_6031,N_6082);
nand U6413 (N_6413,N_6246,N_6098);
and U6414 (N_6414,N_6118,N_6067);
and U6415 (N_6415,N_6067,N_6198);
and U6416 (N_6416,N_6110,N_6209);
xor U6417 (N_6417,N_6140,N_6183);
nand U6418 (N_6418,N_6136,N_6192);
nor U6419 (N_6419,N_6026,N_6025);
or U6420 (N_6420,N_6180,N_6221);
nor U6421 (N_6421,N_6089,N_6016);
nand U6422 (N_6422,N_6233,N_6244);
nand U6423 (N_6423,N_6105,N_6185);
nand U6424 (N_6424,N_6004,N_6006);
or U6425 (N_6425,N_6056,N_6045);
or U6426 (N_6426,N_6220,N_6024);
or U6427 (N_6427,N_6049,N_6109);
xor U6428 (N_6428,N_6002,N_6236);
xnor U6429 (N_6429,N_6014,N_6208);
or U6430 (N_6430,N_6192,N_6249);
nand U6431 (N_6431,N_6159,N_6034);
nor U6432 (N_6432,N_6120,N_6075);
and U6433 (N_6433,N_6023,N_6227);
or U6434 (N_6434,N_6217,N_6150);
and U6435 (N_6435,N_6043,N_6130);
xnor U6436 (N_6436,N_6240,N_6048);
xor U6437 (N_6437,N_6007,N_6131);
nor U6438 (N_6438,N_6015,N_6139);
nand U6439 (N_6439,N_6037,N_6106);
nor U6440 (N_6440,N_6005,N_6098);
xnor U6441 (N_6441,N_6143,N_6169);
nor U6442 (N_6442,N_6000,N_6011);
or U6443 (N_6443,N_6249,N_6071);
and U6444 (N_6444,N_6112,N_6022);
xnor U6445 (N_6445,N_6123,N_6080);
and U6446 (N_6446,N_6191,N_6154);
and U6447 (N_6447,N_6032,N_6157);
xor U6448 (N_6448,N_6154,N_6151);
or U6449 (N_6449,N_6022,N_6014);
nand U6450 (N_6450,N_6017,N_6031);
and U6451 (N_6451,N_6146,N_6092);
or U6452 (N_6452,N_6009,N_6025);
or U6453 (N_6453,N_6247,N_6216);
and U6454 (N_6454,N_6185,N_6174);
or U6455 (N_6455,N_6100,N_6066);
nor U6456 (N_6456,N_6206,N_6140);
and U6457 (N_6457,N_6144,N_6155);
and U6458 (N_6458,N_6177,N_6148);
xnor U6459 (N_6459,N_6243,N_6024);
and U6460 (N_6460,N_6096,N_6059);
or U6461 (N_6461,N_6207,N_6249);
and U6462 (N_6462,N_6192,N_6193);
nor U6463 (N_6463,N_6019,N_6233);
xor U6464 (N_6464,N_6181,N_6051);
xor U6465 (N_6465,N_6132,N_6077);
or U6466 (N_6466,N_6185,N_6144);
and U6467 (N_6467,N_6239,N_6057);
nand U6468 (N_6468,N_6236,N_6015);
and U6469 (N_6469,N_6138,N_6233);
xor U6470 (N_6470,N_6133,N_6150);
and U6471 (N_6471,N_6115,N_6052);
xnor U6472 (N_6472,N_6040,N_6030);
and U6473 (N_6473,N_6031,N_6132);
xor U6474 (N_6474,N_6235,N_6055);
nor U6475 (N_6475,N_6061,N_6203);
or U6476 (N_6476,N_6229,N_6222);
nor U6477 (N_6477,N_6020,N_6023);
and U6478 (N_6478,N_6046,N_6084);
nor U6479 (N_6479,N_6153,N_6030);
and U6480 (N_6480,N_6196,N_6195);
and U6481 (N_6481,N_6154,N_6158);
nand U6482 (N_6482,N_6205,N_6016);
or U6483 (N_6483,N_6016,N_6037);
and U6484 (N_6484,N_6132,N_6156);
xnor U6485 (N_6485,N_6005,N_6018);
and U6486 (N_6486,N_6207,N_6171);
nand U6487 (N_6487,N_6176,N_6047);
nor U6488 (N_6488,N_6229,N_6225);
and U6489 (N_6489,N_6159,N_6035);
nor U6490 (N_6490,N_6139,N_6020);
nor U6491 (N_6491,N_6238,N_6194);
xor U6492 (N_6492,N_6229,N_6000);
or U6493 (N_6493,N_6062,N_6189);
and U6494 (N_6494,N_6028,N_6116);
nor U6495 (N_6495,N_6013,N_6168);
and U6496 (N_6496,N_6197,N_6023);
nand U6497 (N_6497,N_6128,N_6225);
nand U6498 (N_6498,N_6122,N_6021);
nor U6499 (N_6499,N_6055,N_6087);
nand U6500 (N_6500,N_6263,N_6370);
xor U6501 (N_6501,N_6447,N_6381);
xnor U6502 (N_6502,N_6451,N_6482);
or U6503 (N_6503,N_6322,N_6304);
nor U6504 (N_6504,N_6262,N_6252);
xnor U6505 (N_6505,N_6391,N_6455);
or U6506 (N_6506,N_6278,N_6386);
or U6507 (N_6507,N_6303,N_6290);
nand U6508 (N_6508,N_6426,N_6399);
nor U6509 (N_6509,N_6312,N_6376);
nand U6510 (N_6510,N_6352,N_6325);
nor U6511 (N_6511,N_6483,N_6436);
xnor U6512 (N_6512,N_6354,N_6372);
nor U6513 (N_6513,N_6490,N_6333);
nor U6514 (N_6514,N_6435,N_6350);
nand U6515 (N_6515,N_6294,N_6321);
and U6516 (N_6516,N_6470,N_6261);
nand U6517 (N_6517,N_6405,N_6416);
or U6518 (N_6518,N_6411,N_6412);
or U6519 (N_6519,N_6410,N_6375);
or U6520 (N_6520,N_6438,N_6433);
nor U6521 (N_6521,N_6496,N_6434);
nand U6522 (N_6522,N_6488,N_6337);
or U6523 (N_6523,N_6346,N_6291);
xor U6524 (N_6524,N_6251,N_6268);
nand U6525 (N_6525,N_6477,N_6485);
and U6526 (N_6526,N_6383,N_6397);
and U6527 (N_6527,N_6307,N_6419);
nor U6528 (N_6528,N_6260,N_6420);
nand U6529 (N_6529,N_6439,N_6403);
nand U6530 (N_6530,N_6341,N_6393);
and U6531 (N_6531,N_6314,N_6331);
xor U6532 (N_6532,N_6301,N_6457);
nor U6533 (N_6533,N_6497,N_6306);
or U6534 (N_6534,N_6284,N_6495);
nand U6535 (N_6535,N_6428,N_6368);
xor U6536 (N_6536,N_6305,N_6308);
nor U6537 (N_6537,N_6493,N_6392);
nand U6538 (N_6538,N_6300,N_6287);
and U6539 (N_6539,N_6417,N_6257);
nand U6540 (N_6540,N_6334,N_6320);
and U6541 (N_6541,N_6258,N_6423);
nand U6542 (N_6542,N_6437,N_6414);
nor U6543 (N_6543,N_6398,N_6282);
nand U6544 (N_6544,N_6345,N_6395);
and U6545 (N_6545,N_6315,N_6358);
nor U6546 (N_6546,N_6269,N_6371);
xnor U6547 (N_6547,N_6288,N_6431);
nor U6548 (N_6548,N_6448,N_6449);
nor U6549 (N_6549,N_6336,N_6342);
nand U6550 (N_6550,N_6274,N_6265);
nand U6551 (N_6551,N_6427,N_6357);
or U6552 (N_6552,N_6463,N_6384);
or U6553 (N_6553,N_6409,N_6317);
nor U6554 (N_6554,N_6316,N_6408);
and U6555 (N_6555,N_6273,N_6299);
or U6556 (N_6556,N_6276,N_6492);
nor U6557 (N_6557,N_6464,N_6298);
or U6558 (N_6558,N_6311,N_6330);
nand U6559 (N_6559,N_6347,N_6481);
xnor U6560 (N_6560,N_6476,N_6379);
nor U6561 (N_6561,N_6474,N_6388);
xor U6562 (N_6562,N_6400,N_6326);
and U6563 (N_6563,N_6430,N_6309);
and U6564 (N_6564,N_6478,N_6327);
nor U6565 (N_6565,N_6429,N_6359);
or U6566 (N_6566,N_6259,N_6421);
xnor U6567 (N_6567,N_6343,N_6486);
or U6568 (N_6568,N_6285,N_6365);
nor U6569 (N_6569,N_6382,N_6443);
nand U6570 (N_6570,N_6461,N_6329);
or U6571 (N_6571,N_6389,N_6494);
or U6572 (N_6572,N_6289,N_6394);
xor U6573 (N_6573,N_6351,N_6456);
or U6574 (N_6574,N_6498,N_6344);
nor U6575 (N_6575,N_6479,N_6332);
nand U6576 (N_6576,N_6446,N_6418);
xor U6577 (N_6577,N_6462,N_6387);
or U6578 (N_6578,N_6441,N_6264);
nor U6579 (N_6579,N_6360,N_6292);
nand U6580 (N_6580,N_6356,N_6487);
nand U6581 (N_6581,N_6415,N_6280);
nor U6582 (N_6582,N_6362,N_6297);
nand U6583 (N_6583,N_6374,N_6489);
nand U6584 (N_6584,N_6422,N_6484);
nand U6585 (N_6585,N_6338,N_6450);
nand U6586 (N_6586,N_6302,N_6324);
and U6587 (N_6587,N_6401,N_6459);
or U6588 (N_6588,N_6369,N_6271);
nor U6589 (N_6589,N_6293,N_6458);
nand U6590 (N_6590,N_6339,N_6283);
xor U6591 (N_6591,N_6465,N_6404);
and U6592 (N_6592,N_6250,N_6442);
xor U6593 (N_6593,N_6385,N_6367);
nand U6594 (N_6594,N_6266,N_6452);
and U6595 (N_6595,N_6254,N_6406);
or U6596 (N_6596,N_6281,N_6468);
nor U6597 (N_6597,N_6445,N_6253);
and U6598 (N_6598,N_6255,N_6440);
xnor U6599 (N_6599,N_6335,N_6475);
nor U6600 (N_6600,N_6467,N_6364);
xor U6601 (N_6601,N_6349,N_6270);
or U6602 (N_6602,N_6363,N_6396);
nor U6603 (N_6603,N_6340,N_6377);
xnor U6604 (N_6604,N_6402,N_6256);
nor U6605 (N_6605,N_6366,N_6296);
and U6606 (N_6606,N_6361,N_6318);
nor U6607 (N_6607,N_6380,N_6453);
nand U6608 (N_6608,N_6425,N_6286);
or U6609 (N_6609,N_6319,N_6373);
xor U6610 (N_6610,N_6499,N_6471);
nand U6611 (N_6611,N_6444,N_6413);
xor U6612 (N_6612,N_6491,N_6275);
nand U6613 (N_6613,N_6454,N_6355);
nand U6614 (N_6614,N_6432,N_6480);
or U6615 (N_6615,N_6469,N_6323);
or U6616 (N_6616,N_6279,N_6472);
nor U6617 (N_6617,N_6378,N_6277);
or U6618 (N_6618,N_6295,N_6348);
or U6619 (N_6619,N_6407,N_6460);
and U6620 (N_6620,N_6466,N_6353);
nor U6621 (N_6621,N_6272,N_6267);
nor U6622 (N_6622,N_6473,N_6424);
or U6623 (N_6623,N_6313,N_6390);
nor U6624 (N_6624,N_6310,N_6328);
and U6625 (N_6625,N_6486,N_6481);
nand U6626 (N_6626,N_6473,N_6458);
and U6627 (N_6627,N_6413,N_6479);
nor U6628 (N_6628,N_6286,N_6389);
nor U6629 (N_6629,N_6313,N_6463);
nand U6630 (N_6630,N_6434,N_6466);
xor U6631 (N_6631,N_6433,N_6474);
xor U6632 (N_6632,N_6367,N_6387);
or U6633 (N_6633,N_6453,N_6277);
xnor U6634 (N_6634,N_6354,N_6297);
nand U6635 (N_6635,N_6265,N_6268);
nor U6636 (N_6636,N_6398,N_6469);
and U6637 (N_6637,N_6487,N_6490);
nor U6638 (N_6638,N_6497,N_6398);
nand U6639 (N_6639,N_6330,N_6407);
nor U6640 (N_6640,N_6276,N_6325);
xnor U6641 (N_6641,N_6388,N_6493);
xnor U6642 (N_6642,N_6438,N_6277);
and U6643 (N_6643,N_6347,N_6259);
nand U6644 (N_6644,N_6431,N_6333);
nor U6645 (N_6645,N_6372,N_6373);
or U6646 (N_6646,N_6298,N_6321);
nor U6647 (N_6647,N_6332,N_6461);
or U6648 (N_6648,N_6278,N_6415);
or U6649 (N_6649,N_6273,N_6349);
xor U6650 (N_6650,N_6433,N_6402);
nor U6651 (N_6651,N_6488,N_6412);
nor U6652 (N_6652,N_6331,N_6440);
nor U6653 (N_6653,N_6286,N_6300);
xor U6654 (N_6654,N_6342,N_6362);
nand U6655 (N_6655,N_6261,N_6491);
nor U6656 (N_6656,N_6406,N_6381);
or U6657 (N_6657,N_6329,N_6410);
nor U6658 (N_6658,N_6257,N_6382);
nand U6659 (N_6659,N_6496,N_6354);
and U6660 (N_6660,N_6455,N_6403);
or U6661 (N_6661,N_6322,N_6456);
xor U6662 (N_6662,N_6353,N_6269);
nor U6663 (N_6663,N_6380,N_6494);
nand U6664 (N_6664,N_6365,N_6254);
and U6665 (N_6665,N_6483,N_6293);
and U6666 (N_6666,N_6461,N_6306);
and U6667 (N_6667,N_6383,N_6407);
xor U6668 (N_6668,N_6492,N_6437);
nor U6669 (N_6669,N_6498,N_6444);
or U6670 (N_6670,N_6450,N_6329);
nand U6671 (N_6671,N_6265,N_6465);
nor U6672 (N_6672,N_6432,N_6406);
or U6673 (N_6673,N_6438,N_6453);
nand U6674 (N_6674,N_6439,N_6471);
xor U6675 (N_6675,N_6281,N_6487);
or U6676 (N_6676,N_6288,N_6270);
nor U6677 (N_6677,N_6364,N_6366);
nor U6678 (N_6678,N_6320,N_6453);
xnor U6679 (N_6679,N_6384,N_6316);
nor U6680 (N_6680,N_6484,N_6266);
xor U6681 (N_6681,N_6417,N_6395);
and U6682 (N_6682,N_6328,N_6255);
or U6683 (N_6683,N_6328,N_6394);
nor U6684 (N_6684,N_6322,N_6348);
nor U6685 (N_6685,N_6461,N_6454);
and U6686 (N_6686,N_6431,N_6342);
or U6687 (N_6687,N_6362,N_6366);
and U6688 (N_6688,N_6397,N_6437);
or U6689 (N_6689,N_6276,N_6485);
nor U6690 (N_6690,N_6280,N_6392);
nand U6691 (N_6691,N_6377,N_6417);
nor U6692 (N_6692,N_6312,N_6445);
xnor U6693 (N_6693,N_6267,N_6370);
nor U6694 (N_6694,N_6477,N_6306);
nor U6695 (N_6695,N_6336,N_6394);
nor U6696 (N_6696,N_6391,N_6305);
and U6697 (N_6697,N_6467,N_6355);
xor U6698 (N_6698,N_6436,N_6484);
nor U6699 (N_6699,N_6446,N_6460);
and U6700 (N_6700,N_6362,N_6311);
xnor U6701 (N_6701,N_6291,N_6494);
nand U6702 (N_6702,N_6438,N_6478);
xnor U6703 (N_6703,N_6264,N_6299);
nor U6704 (N_6704,N_6394,N_6389);
and U6705 (N_6705,N_6498,N_6362);
xor U6706 (N_6706,N_6438,N_6397);
or U6707 (N_6707,N_6410,N_6318);
or U6708 (N_6708,N_6356,N_6373);
nor U6709 (N_6709,N_6342,N_6386);
or U6710 (N_6710,N_6386,N_6429);
nor U6711 (N_6711,N_6279,N_6487);
nand U6712 (N_6712,N_6399,N_6383);
or U6713 (N_6713,N_6257,N_6250);
nor U6714 (N_6714,N_6434,N_6287);
nor U6715 (N_6715,N_6318,N_6425);
nand U6716 (N_6716,N_6486,N_6254);
nand U6717 (N_6717,N_6359,N_6304);
nand U6718 (N_6718,N_6350,N_6287);
nor U6719 (N_6719,N_6404,N_6396);
or U6720 (N_6720,N_6376,N_6475);
and U6721 (N_6721,N_6287,N_6362);
nor U6722 (N_6722,N_6266,N_6258);
nor U6723 (N_6723,N_6474,N_6451);
or U6724 (N_6724,N_6496,N_6350);
and U6725 (N_6725,N_6468,N_6483);
xnor U6726 (N_6726,N_6425,N_6309);
xor U6727 (N_6727,N_6281,N_6306);
nand U6728 (N_6728,N_6396,N_6408);
nand U6729 (N_6729,N_6366,N_6352);
or U6730 (N_6730,N_6430,N_6366);
nand U6731 (N_6731,N_6300,N_6275);
xnor U6732 (N_6732,N_6348,N_6471);
or U6733 (N_6733,N_6363,N_6372);
or U6734 (N_6734,N_6329,N_6387);
nand U6735 (N_6735,N_6498,N_6347);
xnor U6736 (N_6736,N_6378,N_6381);
xor U6737 (N_6737,N_6365,N_6460);
and U6738 (N_6738,N_6438,N_6269);
nor U6739 (N_6739,N_6499,N_6446);
and U6740 (N_6740,N_6305,N_6358);
nor U6741 (N_6741,N_6452,N_6374);
xor U6742 (N_6742,N_6260,N_6321);
or U6743 (N_6743,N_6335,N_6431);
or U6744 (N_6744,N_6481,N_6356);
nor U6745 (N_6745,N_6261,N_6493);
nor U6746 (N_6746,N_6498,N_6267);
nand U6747 (N_6747,N_6400,N_6366);
nand U6748 (N_6748,N_6470,N_6387);
and U6749 (N_6749,N_6426,N_6299);
xnor U6750 (N_6750,N_6695,N_6561);
nand U6751 (N_6751,N_6585,N_6517);
xnor U6752 (N_6752,N_6655,N_6646);
or U6753 (N_6753,N_6719,N_6625);
and U6754 (N_6754,N_6748,N_6729);
nor U6755 (N_6755,N_6605,N_6688);
and U6756 (N_6756,N_6707,N_6575);
nor U6757 (N_6757,N_6736,N_6545);
nor U6758 (N_6758,N_6713,N_6705);
and U6759 (N_6759,N_6535,N_6744);
or U6760 (N_6760,N_6697,N_6685);
xnor U6761 (N_6761,N_6555,N_6657);
nand U6762 (N_6762,N_6531,N_6518);
nor U6763 (N_6763,N_6570,N_6659);
and U6764 (N_6764,N_6673,N_6572);
nor U6765 (N_6765,N_6714,N_6591);
nor U6766 (N_6766,N_6709,N_6542);
nand U6767 (N_6767,N_6633,N_6541);
and U6768 (N_6768,N_6666,N_6717);
xor U6769 (N_6769,N_6619,N_6601);
xnor U6770 (N_6770,N_6512,N_6574);
nand U6771 (N_6771,N_6608,N_6690);
xor U6772 (N_6772,N_6500,N_6505);
or U6773 (N_6773,N_6703,N_6735);
xor U6774 (N_6774,N_6711,N_6521);
and U6775 (N_6775,N_6581,N_6653);
nand U6776 (N_6776,N_6642,N_6661);
nand U6777 (N_6777,N_6527,N_6746);
or U6778 (N_6778,N_6507,N_6632);
and U6779 (N_6779,N_6595,N_6638);
nand U6780 (N_6780,N_6648,N_6700);
xnor U6781 (N_6781,N_6715,N_6547);
or U6782 (N_6782,N_6662,N_6613);
or U6783 (N_6783,N_6647,N_6565);
nor U6784 (N_6784,N_6698,N_6568);
or U6785 (N_6785,N_6566,N_6723);
xnor U6786 (N_6786,N_6731,N_6628);
nor U6787 (N_6787,N_6706,N_6664);
nor U6788 (N_6788,N_6600,N_6597);
nor U6789 (N_6789,N_6520,N_6615);
nor U6790 (N_6790,N_6617,N_6501);
nor U6791 (N_6791,N_6559,N_6506);
nor U6792 (N_6792,N_6534,N_6645);
nand U6793 (N_6793,N_6641,N_6553);
and U6794 (N_6794,N_6623,N_6519);
nor U6795 (N_6795,N_6684,N_6543);
or U6796 (N_6796,N_6699,N_6636);
and U6797 (N_6797,N_6676,N_6660);
nand U6798 (N_6798,N_6528,N_6590);
or U6799 (N_6799,N_6728,N_6532);
and U6800 (N_6800,N_6670,N_6672);
and U6801 (N_6801,N_6589,N_6571);
nor U6802 (N_6802,N_6671,N_6607);
xnor U6803 (N_6803,N_6624,N_6549);
xnor U6804 (N_6804,N_6739,N_6708);
nor U6805 (N_6805,N_6540,N_6742);
nor U6806 (N_6806,N_6712,N_6745);
and U6807 (N_6807,N_6665,N_6663);
xnor U6808 (N_6808,N_6612,N_6669);
or U6809 (N_6809,N_6720,N_6567);
nor U6810 (N_6810,N_6503,N_6586);
nand U6811 (N_6811,N_6515,N_6588);
xnor U6812 (N_6812,N_6630,N_6569);
xor U6813 (N_6813,N_6654,N_6573);
nand U6814 (N_6814,N_6677,N_6580);
xnor U6815 (N_6815,N_6522,N_6526);
nor U6816 (N_6816,N_6725,N_6734);
nor U6817 (N_6817,N_6609,N_6579);
and U6818 (N_6818,N_6726,N_6694);
xnor U6819 (N_6819,N_6656,N_6738);
or U6820 (N_6820,N_6516,N_6626);
nor U6821 (N_6821,N_6651,N_6618);
xor U6822 (N_6822,N_6554,N_6675);
nor U6823 (N_6823,N_6737,N_6548);
nor U6824 (N_6824,N_6639,N_6552);
or U6825 (N_6825,N_6678,N_6640);
nand U6826 (N_6826,N_6538,N_6686);
xnor U6827 (N_6827,N_6604,N_6718);
or U6828 (N_6828,N_6693,N_6616);
nor U6829 (N_6829,N_6602,N_6667);
and U6830 (N_6830,N_6603,N_6594);
nor U6831 (N_6831,N_6740,N_6556);
xnor U6832 (N_6832,N_6682,N_6701);
or U6833 (N_6833,N_6610,N_6696);
nor U6834 (N_6834,N_6599,N_6587);
xor U6835 (N_6835,N_6546,N_6502);
or U6836 (N_6836,N_6577,N_6523);
or U6837 (N_6837,N_6509,N_6564);
nand U6838 (N_6838,N_6674,N_6691);
xnor U6839 (N_6839,N_6514,N_6747);
and U6840 (N_6840,N_6544,N_6652);
xnor U6841 (N_6841,N_6710,N_6578);
nand U6842 (N_6842,N_6598,N_6724);
nand U6843 (N_6843,N_6689,N_6687);
nand U6844 (N_6844,N_6637,N_6635);
nor U6845 (N_6845,N_6649,N_6644);
xor U6846 (N_6846,N_6537,N_6621);
nor U6847 (N_6847,N_6508,N_6563);
nor U6848 (N_6848,N_6692,N_6683);
nor U6849 (N_6849,N_6627,N_6614);
nor U6850 (N_6850,N_6530,N_6557);
or U6851 (N_6851,N_6582,N_6643);
and U6852 (N_6852,N_6593,N_6727);
or U6853 (N_6853,N_6504,N_6562);
nand U6854 (N_6854,N_6510,N_6679);
nor U6855 (N_6855,N_6732,N_6629);
and U6856 (N_6856,N_6611,N_6536);
or U6857 (N_6857,N_6533,N_6733);
nor U6858 (N_6858,N_6511,N_6584);
nand U6859 (N_6859,N_6539,N_6631);
and U6860 (N_6860,N_6622,N_6560);
xor U6861 (N_6861,N_6716,N_6524);
nor U6862 (N_6862,N_6722,N_6741);
and U6863 (N_6863,N_6583,N_6596);
xor U6864 (N_6864,N_6668,N_6704);
and U6865 (N_6865,N_6730,N_6749);
nor U6866 (N_6866,N_6658,N_6606);
xor U6867 (N_6867,N_6576,N_6702);
or U6868 (N_6868,N_6558,N_6550);
xnor U6869 (N_6869,N_6680,N_6513);
and U6870 (N_6870,N_6551,N_6634);
or U6871 (N_6871,N_6529,N_6650);
xor U6872 (N_6872,N_6620,N_6592);
nand U6873 (N_6873,N_6743,N_6525);
or U6874 (N_6874,N_6681,N_6721);
nor U6875 (N_6875,N_6574,N_6677);
or U6876 (N_6876,N_6712,N_6539);
nor U6877 (N_6877,N_6613,N_6621);
or U6878 (N_6878,N_6638,N_6521);
or U6879 (N_6879,N_6607,N_6538);
and U6880 (N_6880,N_6540,N_6537);
and U6881 (N_6881,N_6518,N_6719);
nand U6882 (N_6882,N_6636,N_6719);
and U6883 (N_6883,N_6608,N_6504);
xnor U6884 (N_6884,N_6589,N_6715);
or U6885 (N_6885,N_6506,N_6741);
nand U6886 (N_6886,N_6748,N_6689);
and U6887 (N_6887,N_6700,N_6671);
nor U6888 (N_6888,N_6607,N_6699);
xnor U6889 (N_6889,N_6664,N_6707);
nand U6890 (N_6890,N_6643,N_6725);
nand U6891 (N_6891,N_6537,N_6620);
nor U6892 (N_6892,N_6681,N_6691);
and U6893 (N_6893,N_6508,N_6542);
nor U6894 (N_6894,N_6736,N_6547);
nand U6895 (N_6895,N_6636,N_6681);
nand U6896 (N_6896,N_6645,N_6683);
xnor U6897 (N_6897,N_6604,N_6723);
nor U6898 (N_6898,N_6542,N_6546);
nand U6899 (N_6899,N_6543,N_6707);
nand U6900 (N_6900,N_6720,N_6736);
xnor U6901 (N_6901,N_6687,N_6605);
or U6902 (N_6902,N_6734,N_6748);
nand U6903 (N_6903,N_6540,N_6524);
and U6904 (N_6904,N_6601,N_6720);
nor U6905 (N_6905,N_6642,N_6676);
and U6906 (N_6906,N_6633,N_6718);
nand U6907 (N_6907,N_6592,N_6588);
or U6908 (N_6908,N_6671,N_6677);
xnor U6909 (N_6909,N_6549,N_6663);
or U6910 (N_6910,N_6573,N_6561);
xor U6911 (N_6911,N_6600,N_6591);
or U6912 (N_6912,N_6684,N_6747);
nor U6913 (N_6913,N_6542,N_6600);
and U6914 (N_6914,N_6645,N_6548);
xor U6915 (N_6915,N_6688,N_6571);
nand U6916 (N_6916,N_6686,N_6682);
xnor U6917 (N_6917,N_6744,N_6696);
or U6918 (N_6918,N_6733,N_6537);
and U6919 (N_6919,N_6587,N_6736);
nand U6920 (N_6920,N_6631,N_6509);
nor U6921 (N_6921,N_6511,N_6670);
nor U6922 (N_6922,N_6584,N_6615);
or U6923 (N_6923,N_6662,N_6624);
nor U6924 (N_6924,N_6584,N_6696);
and U6925 (N_6925,N_6691,N_6569);
and U6926 (N_6926,N_6698,N_6641);
xnor U6927 (N_6927,N_6539,N_6541);
or U6928 (N_6928,N_6590,N_6613);
nor U6929 (N_6929,N_6682,N_6522);
nor U6930 (N_6930,N_6681,N_6642);
nand U6931 (N_6931,N_6558,N_6712);
nor U6932 (N_6932,N_6548,N_6516);
and U6933 (N_6933,N_6706,N_6729);
and U6934 (N_6934,N_6630,N_6521);
or U6935 (N_6935,N_6686,N_6550);
or U6936 (N_6936,N_6546,N_6715);
nand U6937 (N_6937,N_6643,N_6695);
nor U6938 (N_6938,N_6711,N_6683);
nor U6939 (N_6939,N_6616,N_6546);
nor U6940 (N_6940,N_6629,N_6549);
nand U6941 (N_6941,N_6713,N_6691);
nor U6942 (N_6942,N_6614,N_6671);
nand U6943 (N_6943,N_6516,N_6708);
xor U6944 (N_6944,N_6619,N_6535);
and U6945 (N_6945,N_6647,N_6626);
nand U6946 (N_6946,N_6635,N_6517);
nor U6947 (N_6947,N_6625,N_6528);
nand U6948 (N_6948,N_6547,N_6545);
xor U6949 (N_6949,N_6558,N_6715);
nor U6950 (N_6950,N_6646,N_6706);
nor U6951 (N_6951,N_6616,N_6539);
xnor U6952 (N_6952,N_6516,N_6563);
or U6953 (N_6953,N_6631,N_6533);
xnor U6954 (N_6954,N_6649,N_6704);
and U6955 (N_6955,N_6563,N_6733);
and U6956 (N_6956,N_6740,N_6560);
xor U6957 (N_6957,N_6637,N_6712);
nor U6958 (N_6958,N_6746,N_6545);
and U6959 (N_6959,N_6504,N_6551);
or U6960 (N_6960,N_6664,N_6527);
xnor U6961 (N_6961,N_6651,N_6611);
or U6962 (N_6962,N_6698,N_6519);
nand U6963 (N_6963,N_6696,N_6602);
xor U6964 (N_6964,N_6614,N_6692);
xnor U6965 (N_6965,N_6570,N_6683);
nand U6966 (N_6966,N_6603,N_6591);
nor U6967 (N_6967,N_6687,N_6584);
xor U6968 (N_6968,N_6646,N_6630);
nand U6969 (N_6969,N_6662,N_6502);
nand U6970 (N_6970,N_6554,N_6701);
and U6971 (N_6971,N_6660,N_6515);
nor U6972 (N_6972,N_6500,N_6601);
xor U6973 (N_6973,N_6747,N_6695);
nor U6974 (N_6974,N_6644,N_6739);
nor U6975 (N_6975,N_6619,N_6729);
nor U6976 (N_6976,N_6711,N_6579);
or U6977 (N_6977,N_6534,N_6559);
or U6978 (N_6978,N_6532,N_6669);
and U6979 (N_6979,N_6735,N_6564);
xnor U6980 (N_6980,N_6667,N_6689);
nand U6981 (N_6981,N_6667,N_6576);
nand U6982 (N_6982,N_6569,N_6562);
and U6983 (N_6983,N_6727,N_6723);
nand U6984 (N_6984,N_6694,N_6680);
nand U6985 (N_6985,N_6674,N_6710);
or U6986 (N_6986,N_6585,N_6666);
nor U6987 (N_6987,N_6648,N_6581);
or U6988 (N_6988,N_6701,N_6737);
and U6989 (N_6989,N_6731,N_6504);
or U6990 (N_6990,N_6607,N_6657);
and U6991 (N_6991,N_6652,N_6513);
xor U6992 (N_6992,N_6546,N_6631);
nor U6993 (N_6993,N_6673,N_6589);
or U6994 (N_6994,N_6715,N_6651);
or U6995 (N_6995,N_6647,N_6538);
and U6996 (N_6996,N_6535,N_6730);
or U6997 (N_6997,N_6659,N_6745);
nor U6998 (N_6998,N_6749,N_6698);
xor U6999 (N_6999,N_6723,N_6583);
xor U7000 (N_7000,N_6788,N_6843);
or U7001 (N_7001,N_6923,N_6922);
or U7002 (N_7002,N_6967,N_6789);
or U7003 (N_7003,N_6831,N_6960);
nor U7004 (N_7004,N_6840,N_6759);
or U7005 (N_7005,N_6862,N_6750);
and U7006 (N_7006,N_6914,N_6863);
nor U7007 (N_7007,N_6926,N_6776);
and U7008 (N_7008,N_6835,N_6774);
nor U7009 (N_7009,N_6818,N_6753);
and U7010 (N_7010,N_6954,N_6891);
nor U7011 (N_7011,N_6983,N_6907);
and U7012 (N_7012,N_6956,N_6844);
xnor U7013 (N_7013,N_6885,N_6880);
nor U7014 (N_7014,N_6911,N_6815);
and U7015 (N_7015,N_6790,N_6764);
nor U7016 (N_7016,N_6782,N_6942);
nand U7017 (N_7017,N_6795,N_6808);
nor U7018 (N_7018,N_6821,N_6864);
and U7019 (N_7019,N_6847,N_6872);
and U7020 (N_7020,N_6806,N_6996);
nor U7021 (N_7021,N_6785,N_6921);
nand U7022 (N_7022,N_6991,N_6841);
and U7023 (N_7023,N_6909,N_6895);
nand U7024 (N_7024,N_6781,N_6974);
or U7025 (N_7025,N_6910,N_6933);
or U7026 (N_7026,N_6934,N_6984);
xnor U7027 (N_7027,N_6856,N_6842);
nor U7028 (N_7028,N_6780,N_6938);
and U7029 (N_7029,N_6888,N_6770);
xnor U7030 (N_7030,N_6925,N_6980);
nor U7031 (N_7031,N_6825,N_6928);
xnor U7032 (N_7032,N_6773,N_6837);
or U7033 (N_7033,N_6758,N_6771);
xnor U7034 (N_7034,N_6828,N_6929);
xnor U7035 (N_7035,N_6882,N_6939);
nor U7036 (N_7036,N_6869,N_6777);
xnor U7037 (N_7037,N_6876,N_6999);
nand U7038 (N_7038,N_6778,N_6755);
or U7039 (N_7039,N_6879,N_6810);
nor U7040 (N_7040,N_6978,N_6903);
nand U7041 (N_7041,N_6887,N_6754);
nor U7042 (N_7042,N_6838,N_6951);
and U7043 (N_7043,N_6853,N_6800);
and U7044 (N_7044,N_6832,N_6982);
or U7045 (N_7045,N_6963,N_6860);
xor U7046 (N_7046,N_6819,N_6913);
or U7047 (N_7047,N_6994,N_6964);
or U7048 (N_7048,N_6944,N_6852);
nor U7049 (N_7049,N_6851,N_6868);
or U7050 (N_7050,N_6937,N_6861);
xnor U7051 (N_7051,N_6897,N_6908);
nor U7052 (N_7052,N_6905,N_6798);
nor U7053 (N_7053,N_6989,N_6892);
or U7054 (N_7054,N_6799,N_6873);
or U7055 (N_7055,N_6902,N_6784);
and U7056 (N_7056,N_6826,N_6816);
nor U7057 (N_7057,N_6920,N_6945);
or U7058 (N_7058,N_6998,N_6855);
or U7059 (N_7059,N_6932,N_6814);
or U7060 (N_7060,N_6765,N_6881);
xor U7061 (N_7061,N_6783,N_6760);
nor U7062 (N_7062,N_6890,N_6950);
nand U7063 (N_7063,N_6805,N_6820);
and U7064 (N_7064,N_6769,N_6969);
and U7065 (N_7065,N_6936,N_6796);
or U7066 (N_7066,N_6977,N_6916);
and U7067 (N_7067,N_6973,N_6833);
or U7068 (N_7068,N_6930,N_6846);
nand U7069 (N_7069,N_6987,N_6889);
xnor U7070 (N_7070,N_6807,N_6988);
xnor U7071 (N_7071,N_6767,N_6952);
and U7072 (N_7072,N_6912,N_6919);
xnor U7073 (N_7073,N_6918,N_6893);
nand U7074 (N_7074,N_6775,N_6940);
nor U7075 (N_7075,N_6866,N_6813);
nand U7076 (N_7076,N_6839,N_6875);
nand U7077 (N_7077,N_6986,N_6965);
nor U7078 (N_7078,N_6896,N_6797);
or U7079 (N_7079,N_6894,N_6823);
and U7080 (N_7080,N_6924,N_6792);
or U7081 (N_7081,N_6824,N_6957);
or U7082 (N_7082,N_6871,N_6948);
or U7083 (N_7083,N_6791,N_6786);
xnor U7084 (N_7084,N_6793,N_6975);
or U7085 (N_7085,N_6985,N_6867);
nand U7086 (N_7086,N_6762,N_6993);
nand U7087 (N_7087,N_6884,N_6834);
nor U7088 (N_7088,N_6886,N_6966);
and U7089 (N_7089,N_6757,N_6899);
or U7090 (N_7090,N_6979,N_6848);
xor U7091 (N_7091,N_6865,N_6915);
nor U7092 (N_7092,N_6959,N_6751);
or U7093 (N_7093,N_6990,N_6845);
or U7094 (N_7094,N_6811,N_6803);
and U7095 (N_7095,N_6830,N_6752);
or U7096 (N_7096,N_6953,N_6904);
nor U7097 (N_7097,N_6766,N_6857);
or U7098 (N_7098,N_6874,N_6970);
nor U7099 (N_7099,N_6961,N_6772);
nand U7100 (N_7100,N_6756,N_6877);
and U7101 (N_7101,N_6958,N_6946);
nor U7102 (N_7102,N_6955,N_6854);
and U7103 (N_7103,N_6878,N_6836);
xor U7104 (N_7104,N_6822,N_6883);
nor U7105 (N_7105,N_6801,N_6906);
nor U7106 (N_7106,N_6850,N_6763);
nor U7107 (N_7107,N_6794,N_6971);
xnor U7108 (N_7108,N_6898,N_6809);
and U7109 (N_7109,N_6817,N_6997);
or U7110 (N_7110,N_6768,N_6787);
nand U7111 (N_7111,N_6931,N_6976);
nand U7112 (N_7112,N_6779,N_6859);
nand U7113 (N_7113,N_6812,N_6949);
nand U7114 (N_7114,N_6804,N_6935);
or U7115 (N_7115,N_6992,N_6858);
and U7116 (N_7116,N_6849,N_6927);
or U7117 (N_7117,N_6962,N_6870);
nor U7118 (N_7118,N_6761,N_6900);
nand U7119 (N_7119,N_6901,N_6981);
nor U7120 (N_7120,N_6827,N_6941);
xnor U7121 (N_7121,N_6943,N_6995);
nor U7122 (N_7122,N_6968,N_6802);
and U7123 (N_7123,N_6829,N_6947);
nor U7124 (N_7124,N_6917,N_6972);
xor U7125 (N_7125,N_6899,N_6859);
or U7126 (N_7126,N_6906,N_6763);
xnor U7127 (N_7127,N_6950,N_6753);
nand U7128 (N_7128,N_6866,N_6912);
xor U7129 (N_7129,N_6928,N_6920);
nor U7130 (N_7130,N_6777,N_6970);
and U7131 (N_7131,N_6867,N_6913);
or U7132 (N_7132,N_6827,N_6814);
and U7133 (N_7133,N_6912,N_6807);
nand U7134 (N_7134,N_6980,N_6899);
or U7135 (N_7135,N_6789,N_6940);
xor U7136 (N_7136,N_6838,N_6979);
or U7137 (N_7137,N_6959,N_6831);
and U7138 (N_7138,N_6780,N_6817);
or U7139 (N_7139,N_6779,N_6783);
or U7140 (N_7140,N_6862,N_6788);
nand U7141 (N_7141,N_6869,N_6852);
xor U7142 (N_7142,N_6942,N_6764);
nand U7143 (N_7143,N_6830,N_6829);
nand U7144 (N_7144,N_6993,N_6957);
or U7145 (N_7145,N_6983,N_6935);
and U7146 (N_7146,N_6834,N_6829);
or U7147 (N_7147,N_6822,N_6754);
nor U7148 (N_7148,N_6940,N_6929);
or U7149 (N_7149,N_6915,N_6899);
xnor U7150 (N_7150,N_6953,N_6861);
nor U7151 (N_7151,N_6865,N_6802);
and U7152 (N_7152,N_6971,N_6991);
xnor U7153 (N_7153,N_6943,N_6949);
nand U7154 (N_7154,N_6894,N_6790);
or U7155 (N_7155,N_6896,N_6970);
nor U7156 (N_7156,N_6982,N_6787);
nor U7157 (N_7157,N_6949,N_6868);
and U7158 (N_7158,N_6892,N_6809);
xor U7159 (N_7159,N_6998,N_6911);
or U7160 (N_7160,N_6818,N_6946);
nand U7161 (N_7161,N_6900,N_6910);
xnor U7162 (N_7162,N_6892,N_6812);
or U7163 (N_7163,N_6813,N_6918);
xor U7164 (N_7164,N_6787,N_6990);
and U7165 (N_7165,N_6786,N_6819);
or U7166 (N_7166,N_6844,N_6996);
xnor U7167 (N_7167,N_6962,N_6904);
xor U7168 (N_7168,N_6794,N_6843);
nor U7169 (N_7169,N_6792,N_6892);
or U7170 (N_7170,N_6860,N_6965);
xor U7171 (N_7171,N_6751,N_6937);
nand U7172 (N_7172,N_6949,N_6921);
nor U7173 (N_7173,N_6922,N_6979);
and U7174 (N_7174,N_6859,N_6870);
and U7175 (N_7175,N_6926,N_6855);
nand U7176 (N_7176,N_6794,N_6819);
and U7177 (N_7177,N_6957,N_6932);
or U7178 (N_7178,N_6926,N_6961);
nor U7179 (N_7179,N_6919,N_6965);
or U7180 (N_7180,N_6959,N_6950);
nand U7181 (N_7181,N_6912,N_6924);
nor U7182 (N_7182,N_6793,N_6993);
nor U7183 (N_7183,N_6939,N_6824);
nor U7184 (N_7184,N_6944,N_6763);
xnor U7185 (N_7185,N_6872,N_6946);
xor U7186 (N_7186,N_6887,N_6904);
xor U7187 (N_7187,N_6779,N_6751);
or U7188 (N_7188,N_6796,N_6986);
or U7189 (N_7189,N_6875,N_6758);
xor U7190 (N_7190,N_6827,N_6996);
nor U7191 (N_7191,N_6873,N_6852);
xor U7192 (N_7192,N_6833,N_6831);
or U7193 (N_7193,N_6804,N_6752);
xnor U7194 (N_7194,N_6855,N_6774);
or U7195 (N_7195,N_6755,N_6926);
xor U7196 (N_7196,N_6918,N_6902);
and U7197 (N_7197,N_6894,N_6827);
nand U7198 (N_7198,N_6825,N_6855);
or U7199 (N_7199,N_6893,N_6921);
nand U7200 (N_7200,N_6969,N_6814);
nand U7201 (N_7201,N_6993,N_6998);
xnor U7202 (N_7202,N_6945,N_6896);
or U7203 (N_7203,N_6851,N_6943);
nor U7204 (N_7204,N_6773,N_6792);
nor U7205 (N_7205,N_6821,N_6867);
nor U7206 (N_7206,N_6750,N_6804);
nand U7207 (N_7207,N_6842,N_6798);
nand U7208 (N_7208,N_6794,N_6967);
and U7209 (N_7209,N_6958,N_6778);
or U7210 (N_7210,N_6766,N_6868);
xnor U7211 (N_7211,N_6973,N_6975);
or U7212 (N_7212,N_6799,N_6946);
and U7213 (N_7213,N_6941,N_6818);
nand U7214 (N_7214,N_6753,N_6768);
xnor U7215 (N_7215,N_6828,N_6820);
and U7216 (N_7216,N_6937,N_6931);
xor U7217 (N_7217,N_6800,N_6767);
xor U7218 (N_7218,N_6787,N_6909);
nor U7219 (N_7219,N_6757,N_6995);
nor U7220 (N_7220,N_6753,N_6851);
nor U7221 (N_7221,N_6824,N_6843);
or U7222 (N_7222,N_6886,N_6982);
and U7223 (N_7223,N_6991,N_6903);
or U7224 (N_7224,N_6805,N_6877);
and U7225 (N_7225,N_6851,N_6957);
xor U7226 (N_7226,N_6764,N_6850);
nor U7227 (N_7227,N_6872,N_6949);
nand U7228 (N_7228,N_6972,N_6924);
nor U7229 (N_7229,N_6895,N_6788);
xnor U7230 (N_7230,N_6984,N_6975);
xnor U7231 (N_7231,N_6911,N_6964);
nand U7232 (N_7232,N_6791,N_6919);
nand U7233 (N_7233,N_6772,N_6766);
nand U7234 (N_7234,N_6936,N_6964);
xor U7235 (N_7235,N_6904,N_6804);
nor U7236 (N_7236,N_6990,N_6905);
or U7237 (N_7237,N_6820,N_6800);
xor U7238 (N_7238,N_6797,N_6814);
nand U7239 (N_7239,N_6805,N_6908);
nor U7240 (N_7240,N_6986,N_6904);
and U7241 (N_7241,N_6952,N_6804);
nor U7242 (N_7242,N_6880,N_6779);
nand U7243 (N_7243,N_6793,N_6949);
xor U7244 (N_7244,N_6768,N_6832);
or U7245 (N_7245,N_6779,N_6887);
or U7246 (N_7246,N_6845,N_6851);
and U7247 (N_7247,N_6865,N_6929);
and U7248 (N_7248,N_6948,N_6927);
or U7249 (N_7249,N_6824,N_6938);
and U7250 (N_7250,N_7084,N_7038);
nand U7251 (N_7251,N_7207,N_7163);
xor U7252 (N_7252,N_7074,N_7123);
xor U7253 (N_7253,N_7202,N_7173);
nand U7254 (N_7254,N_7245,N_7151);
nand U7255 (N_7255,N_7119,N_7107);
and U7256 (N_7256,N_7118,N_7227);
xor U7257 (N_7257,N_7137,N_7078);
or U7258 (N_7258,N_7181,N_7114);
or U7259 (N_7259,N_7154,N_7192);
and U7260 (N_7260,N_7050,N_7172);
nand U7261 (N_7261,N_7153,N_7235);
xor U7262 (N_7262,N_7016,N_7180);
nor U7263 (N_7263,N_7193,N_7035);
or U7264 (N_7264,N_7179,N_7079);
nand U7265 (N_7265,N_7185,N_7054);
nand U7266 (N_7266,N_7162,N_7186);
or U7267 (N_7267,N_7044,N_7146);
and U7268 (N_7268,N_7222,N_7024);
and U7269 (N_7269,N_7093,N_7112);
xnor U7270 (N_7270,N_7003,N_7128);
and U7271 (N_7271,N_7135,N_7108);
and U7272 (N_7272,N_7213,N_7238);
xnor U7273 (N_7273,N_7249,N_7141);
nor U7274 (N_7274,N_7040,N_7053);
nor U7275 (N_7275,N_7198,N_7150);
xor U7276 (N_7276,N_7183,N_7066);
nor U7277 (N_7277,N_7064,N_7023);
or U7278 (N_7278,N_7058,N_7100);
and U7279 (N_7279,N_7011,N_7063);
or U7280 (N_7280,N_7020,N_7158);
nor U7281 (N_7281,N_7019,N_7212);
xnor U7282 (N_7282,N_7095,N_7129);
nand U7283 (N_7283,N_7091,N_7139);
nor U7284 (N_7284,N_7077,N_7232);
and U7285 (N_7285,N_7005,N_7029);
xnor U7286 (N_7286,N_7176,N_7226);
nor U7287 (N_7287,N_7140,N_7057);
or U7288 (N_7288,N_7004,N_7059);
nand U7289 (N_7289,N_7026,N_7142);
and U7290 (N_7290,N_7228,N_7089);
and U7291 (N_7291,N_7027,N_7189);
xor U7292 (N_7292,N_7086,N_7065);
or U7293 (N_7293,N_7076,N_7002);
xor U7294 (N_7294,N_7133,N_7229);
or U7295 (N_7295,N_7081,N_7082);
nand U7296 (N_7296,N_7170,N_7097);
xor U7297 (N_7297,N_7138,N_7014);
nand U7298 (N_7298,N_7007,N_7056);
or U7299 (N_7299,N_7070,N_7116);
or U7300 (N_7300,N_7010,N_7204);
nand U7301 (N_7301,N_7188,N_7117);
nand U7302 (N_7302,N_7194,N_7001);
nor U7303 (N_7303,N_7225,N_7203);
nand U7304 (N_7304,N_7178,N_7083);
or U7305 (N_7305,N_7006,N_7144);
or U7306 (N_7306,N_7092,N_7239);
nor U7307 (N_7307,N_7122,N_7028);
nand U7308 (N_7308,N_7008,N_7115);
and U7309 (N_7309,N_7124,N_7175);
and U7310 (N_7310,N_7171,N_7214);
nand U7311 (N_7311,N_7113,N_7051);
nand U7312 (N_7312,N_7085,N_7021);
nand U7313 (N_7313,N_7145,N_7223);
xor U7314 (N_7314,N_7132,N_7103);
nand U7315 (N_7315,N_7167,N_7060);
and U7316 (N_7316,N_7017,N_7034);
nor U7317 (N_7317,N_7219,N_7080);
or U7318 (N_7318,N_7187,N_7217);
xnor U7319 (N_7319,N_7009,N_7184);
nor U7320 (N_7320,N_7220,N_7088);
nor U7321 (N_7321,N_7157,N_7068);
nor U7322 (N_7322,N_7037,N_7196);
xor U7323 (N_7323,N_7061,N_7071);
and U7324 (N_7324,N_7248,N_7216);
xnor U7325 (N_7325,N_7218,N_7096);
or U7326 (N_7326,N_7165,N_7106);
and U7327 (N_7327,N_7148,N_7247);
or U7328 (N_7328,N_7211,N_7205);
xnor U7329 (N_7329,N_7242,N_7200);
and U7330 (N_7330,N_7075,N_7221);
nand U7331 (N_7331,N_7134,N_7210);
or U7332 (N_7332,N_7043,N_7025);
nand U7333 (N_7333,N_7120,N_7099);
xor U7334 (N_7334,N_7131,N_7030);
xor U7335 (N_7335,N_7126,N_7166);
nand U7336 (N_7336,N_7049,N_7177);
xnor U7337 (N_7337,N_7109,N_7195);
nand U7338 (N_7338,N_7110,N_7127);
nor U7339 (N_7339,N_7168,N_7036);
nor U7340 (N_7340,N_7236,N_7241);
and U7341 (N_7341,N_7201,N_7234);
xnor U7342 (N_7342,N_7243,N_7143);
xnor U7343 (N_7343,N_7244,N_7069);
nor U7344 (N_7344,N_7206,N_7094);
or U7345 (N_7345,N_7160,N_7164);
nand U7346 (N_7346,N_7208,N_7155);
xor U7347 (N_7347,N_7111,N_7047);
nor U7348 (N_7348,N_7015,N_7182);
or U7349 (N_7349,N_7240,N_7224);
nor U7350 (N_7350,N_7121,N_7055);
xor U7351 (N_7351,N_7136,N_7159);
xor U7352 (N_7352,N_7147,N_7161);
and U7353 (N_7353,N_7042,N_7215);
nor U7354 (N_7354,N_7237,N_7018);
xnor U7355 (N_7355,N_7101,N_7169);
or U7356 (N_7356,N_7073,N_7199);
xor U7357 (N_7357,N_7104,N_7067);
or U7358 (N_7358,N_7087,N_7039);
nor U7359 (N_7359,N_7022,N_7046);
or U7360 (N_7360,N_7152,N_7102);
nor U7361 (N_7361,N_7130,N_7045);
xor U7362 (N_7362,N_7032,N_7149);
nand U7363 (N_7363,N_7062,N_7125);
nor U7364 (N_7364,N_7246,N_7230);
nor U7365 (N_7365,N_7052,N_7090);
or U7366 (N_7366,N_7041,N_7209);
and U7367 (N_7367,N_7105,N_7031);
or U7368 (N_7368,N_7174,N_7190);
nand U7369 (N_7369,N_7013,N_7012);
and U7370 (N_7370,N_7048,N_7098);
and U7371 (N_7371,N_7231,N_7000);
xnor U7372 (N_7372,N_7233,N_7191);
xnor U7373 (N_7373,N_7072,N_7033);
or U7374 (N_7374,N_7156,N_7197);
nand U7375 (N_7375,N_7155,N_7174);
xnor U7376 (N_7376,N_7040,N_7132);
and U7377 (N_7377,N_7148,N_7149);
or U7378 (N_7378,N_7018,N_7005);
or U7379 (N_7379,N_7130,N_7136);
nand U7380 (N_7380,N_7028,N_7121);
nand U7381 (N_7381,N_7119,N_7071);
xor U7382 (N_7382,N_7225,N_7074);
xor U7383 (N_7383,N_7106,N_7207);
and U7384 (N_7384,N_7105,N_7074);
nor U7385 (N_7385,N_7152,N_7096);
xor U7386 (N_7386,N_7205,N_7133);
and U7387 (N_7387,N_7184,N_7156);
nand U7388 (N_7388,N_7069,N_7233);
nor U7389 (N_7389,N_7024,N_7118);
nand U7390 (N_7390,N_7017,N_7180);
nand U7391 (N_7391,N_7076,N_7022);
nor U7392 (N_7392,N_7119,N_7040);
or U7393 (N_7393,N_7022,N_7243);
xor U7394 (N_7394,N_7147,N_7171);
and U7395 (N_7395,N_7077,N_7240);
nor U7396 (N_7396,N_7031,N_7160);
or U7397 (N_7397,N_7204,N_7008);
and U7398 (N_7398,N_7092,N_7199);
nand U7399 (N_7399,N_7090,N_7168);
nand U7400 (N_7400,N_7086,N_7120);
nor U7401 (N_7401,N_7047,N_7248);
nand U7402 (N_7402,N_7109,N_7062);
nor U7403 (N_7403,N_7125,N_7180);
or U7404 (N_7404,N_7238,N_7015);
or U7405 (N_7405,N_7089,N_7097);
or U7406 (N_7406,N_7033,N_7180);
and U7407 (N_7407,N_7044,N_7213);
nand U7408 (N_7408,N_7027,N_7012);
and U7409 (N_7409,N_7211,N_7104);
xor U7410 (N_7410,N_7174,N_7160);
and U7411 (N_7411,N_7249,N_7092);
and U7412 (N_7412,N_7148,N_7033);
xor U7413 (N_7413,N_7236,N_7207);
and U7414 (N_7414,N_7241,N_7036);
or U7415 (N_7415,N_7168,N_7094);
xnor U7416 (N_7416,N_7200,N_7100);
nand U7417 (N_7417,N_7134,N_7176);
nand U7418 (N_7418,N_7057,N_7160);
xor U7419 (N_7419,N_7145,N_7103);
and U7420 (N_7420,N_7009,N_7117);
and U7421 (N_7421,N_7223,N_7073);
nand U7422 (N_7422,N_7020,N_7188);
and U7423 (N_7423,N_7019,N_7046);
or U7424 (N_7424,N_7087,N_7029);
and U7425 (N_7425,N_7204,N_7048);
xnor U7426 (N_7426,N_7229,N_7193);
and U7427 (N_7427,N_7205,N_7142);
or U7428 (N_7428,N_7069,N_7143);
nand U7429 (N_7429,N_7228,N_7005);
nor U7430 (N_7430,N_7143,N_7124);
xnor U7431 (N_7431,N_7237,N_7219);
nor U7432 (N_7432,N_7240,N_7081);
nand U7433 (N_7433,N_7160,N_7077);
nand U7434 (N_7434,N_7171,N_7003);
or U7435 (N_7435,N_7074,N_7066);
or U7436 (N_7436,N_7237,N_7132);
xor U7437 (N_7437,N_7042,N_7037);
or U7438 (N_7438,N_7219,N_7184);
nand U7439 (N_7439,N_7046,N_7010);
nand U7440 (N_7440,N_7149,N_7240);
or U7441 (N_7441,N_7083,N_7229);
nand U7442 (N_7442,N_7207,N_7063);
and U7443 (N_7443,N_7056,N_7130);
or U7444 (N_7444,N_7178,N_7110);
nor U7445 (N_7445,N_7032,N_7193);
nand U7446 (N_7446,N_7032,N_7046);
nand U7447 (N_7447,N_7170,N_7054);
nand U7448 (N_7448,N_7029,N_7047);
nand U7449 (N_7449,N_7169,N_7153);
nand U7450 (N_7450,N_7109,N_7005);
nand U7451 (N_7451,N_7074,N_7056);
nor U7452 (N_7452,N_7077,N_7204);
nand U7453 (N_7453,N_7085,N_7116);
nand U7454 (N_7454,N_7156,N_7057);
and U7455 (N_7455,N_7249,N_7061);
and U7456 (N_7456,N_7187,N_7000);
xnor U7457 (N_7457,N_7001,N_7095);
or U7458 (N_7458,N_7160,N_7154);
nand U7459 (N_7459,N_7022,N_7084);
or U7460 (N_7460,N_7105,N_7111);
or U7461 (N_7461,N_7008,N_7026);
or U7462 (N_7462,N_7061,N_7161);
nor U7463 (N_7463,N_7185,N_7247);
nand U7464 (N_7464,N_7042,N_7176);
and U7465 (N_7465,N_7092,N_7161);
xor U7466 (N_7466,N_7104,N_7037);
xor U7467 (N_7467,N_7030,N_7139);
and U7468 (N_7468,N_7151,N_7038);
nor U7469 (N_7469,N_7092,N_7019);
xnor U7470 (N_7470,N_7008,N_7144);
nor U7471 (N_7471,N_7176,N_7135);
nor U7472 (N_7472,N_7163,N_7085);
nor U7473 (N_7473,N_7118,N_7110);
xor U7474 (N_7474,N_7001,N_7152);
or U7475 (N_7475,N_7151,N_7007);
and U7476 (N_7476,N_7006,N_7032);
nand U7477 (N_7477,N_7229,N_7111);
nand U7478 (N_7478,N_7093,N_7215);
or U7479 (N_7479,N_7132,N_7187);
nor U7480 (N_7480,N_7191,N_7133);
nor U7481 (N_7481,N_7045,N_7142);
nor U7482 (N_7482,N_7002,N_7088);
and U7483 (N_7483,N_7134,N_7048);
xnor U7484 (N_7484,N_7157,N_7055);
or U7485 (N_7485,N_7008,N_7138);
or U7486 (N_7486,N_7153,N_7057);
and U7487 (N_7487,N_7022,N_7211);
xnor U7488 (N_7488,N_7002,N_7139);
or U7489 (N_7489,N_7046,N_7083);
nand U7490 (N_7490,N_7173,N_7075);
nor U7491 (N_7491,N_7180,N_7151);
or U7492 (N_7492,N_7247,N_7110);
and U7493 (N_7493,N_7009,N_7212);
or U7494 (N_7494,N_7217,N_7059);
or U7495 (N_7495,N_7044,N_7131);
or U7496 (N_7496,N_7064,N_7183);
and U7497 (N_7497,N_7132,N_7182);
and U7498 (N_7498,N_7002,N_7170);
or U7499 (N_7499,N_7050,N_7007);
or U7500 (N_7500,N_7431,N_7258);
xor U7501 (N_7501,N_7458,N_7349);
nand U7502 (N_7502,N_7407,N_7370);
nor U7503 (N_7503,N_7390,N_7279);
and U7504 (N_7504,N_7317,N_7393);
nor U7505 (N_7505,N_7283,N_7311);
nand U7506 (N_7506,N_7425,N_7356);
and U7507 (N_7507,N_7380,N_7268);
nor U7508 (N_7508,N_7413,N_7281);
nand U7509 (N_7509,N_7453,N_7432);
nand U7510 (N_7510,N_7310,N_7426);
nor U7511 (N_7511,N_7337,N_7411);
or U7512 (N_7512,N_7470,N_7299);
nor U7513 (N_7513,N_7335,N_7468);
or U7514 (N_7514,N_7290,N_7395);
nand U7515 (N_7515,N_7351,N_7348);
or U7516 (N_7516,N_7401,N_7314);
nand U7517 (N_7517,N_7376,N_7260);
and U7518 (N_7518,N_7442,N_7371);
or U7519 (N_7519,N_7386,N_7391);
nand U7520 (N_7520,N_7343,N_7353);
or U7521 (N_7521,N_7369,N_7332);
nand U7522 (N_7522,N_7344,N_7355);
nand U7523 (N_7523,N_7402,N_7307);
xnor U7524 (N_7524,N_7272,N_7338);
nand U7525 (N_7525,N_7493,N_7253);
xor U7526 (N_7526,N_7447,N_7488);
or U7527 (N_7527,N_7275,N_7398);
xor U7528 (N_7528,N_7481,N_7499);
xor U7529 (N_7529,N_7263,N_7477);
and U7530 (N_7530,N_7375,N_7464);
xnor U7531 (N_7531,N_7387,N_7416);
nand U7532 (N_7532,N_7368,N_7408);
or U7533 (N_7533,N_7342,N_7373);
or U7534 (N_7534,N_7300,N_7352);
nor U7535 (N_7535,N_7435,N_7383);
xor U7536 (N_7536,N_7329,N_7446);
or U7537 (N_7537,N_7269,N_7291);
nor U7538 (N_7538,N_7489,N_7271);
nor U7539 (N_7539,N_7436,N_7366);
nor U7540 (N_7540,N_7438,N_7457);
or U7541 (N_7541,N_7400,N_7328);
nand U7542 (N_7542,N_7490,N_7430);
or U7543 (N_7543,N_7264,N_7327);
or U7544 (N_7544,N_7434,N_7360);
xnor U7545 (N_7545,N_7282,N_7418);
nand U7546 (N_7546,N_7350,N_7469);
xor U7547 (N_7547,N_7479,N_7448);
xnor U7548 (N_7548,N_7363,N_7423);
or U7549 (N_7549,N_7491,N_7262);
nand U7550 (N_7550,N_7267,N_7306);
nand U7551 (N_7551,N_7285,N_7340);
and U7552 (N_7552,N_7276,N_7318);
and U7553 (N_7553,N_7452,N_7486);
xnor U7554 (N_7554,N_7384,N_7320);
nand U7555 (N_7555,N_7498,N_7444);
nand U7556 (N_7556,N_7424,N_7456);
or U7557 (N_7557,N_7339,N_7256);
xor U7558 (N_7558,N_7265,N_7455);
nor U7559 (N_7559,N_7428,N_7445);
nor U7560 (N_7560,N_7403,N_7379);
or U7561 (N_7561,N_7295,N_7478);
xor U7562 (N_7562,N_7462,N_7302);
or U7563 (N_7563,N_7345,N_7280);
and U7564 (N_7564,N_7412,N_7266);
and U7565 (N_7565,N_7333,N_7474);
nand U7566 (N_7566,N_7374,N_7392);
and U7567 (N_7567,N_7463,N_7313);
xnor U7568 (N_7568,N_7404,N_7450);
xor U7569 (N_7569,N_7449,N_7485);
or U7570 (N_7570,N_7270,N_7305);
nor U7571 (N_7571,N_7396,N_7322);
and U7572 (N_7572,N_7304,N_7293);
or U7573 (N_7573,N_7461,N_7324);
nand U7574 (N_7574,N_7378,N_7473);
nand U7575 (N_7575,N_7466,N_7251);
xor U7576 (N_7576,N_7397,N_7347);
xor U7577 (N_7577,N_7429,N_7296);
and U7578 (N_7578,N_7406,N_7254);
nand U7579 (N_7579,N_7292,N_7284);
and U7580 (N_7580,N_7382,N_7274);
and U7581 (N_7581,N_7409,N_7309);
or U7582 (N_7582,N_7472,N_7417);
and U7583 (N_7583,N_7331,N_7308);
and U7584 (N_7584,N_7443,N_7261);
nand U7585 (N_7585,N_7287,N_7312);
and U7586 (N_7586,N_7377,N_7467);
xor U7587 (N_7587,N_7250,N_7336);
xnor U7588 (N_7588,N_7494,N_7364);
or U7589 (N_7589,N_7297,N_7437);
and U7590 (N_7590,N_7289,N_7451);
and U7591 (N_7591,N_7294,N_7439);
nand U7592 (N_7592,N_7259,N_7475);
nor U7593 (N_7593,N_7471,N_7358);
nor U7594 (N_7594,N_7422,N_7419);
xnor U7595 (N_7595,N_7394,N_7277);
nor U7596 (N_7596,N_7341,N_7326);
nand U7597 (N_7597,N_7359,N_7315);
nand U7598 (N_7598,N_7414,N_7459);
nor U7599 (N_7599,N_7303,N_7420);
or U7600 (N_7600,N_7362,N_7483);
xnor U7601 (N_7601,N_7288,N_7286);
xnor U7602 (N_7602,N_7357,N_7484);
or U7603 (N_7603,N_7487,N_7316);
xnor U7604 (N_7604,N_7415,N_7454);
xnor U7605 (N_7605,N_7273,N_7440);
nor U7606 (N_7606,N_7323,N_7257);
nand U7607 (N_7607,N_7346,N_7255);
nand U7608 (N_7608,N_7399,N_7252);
and U7609 (N_7609,N_7405,N_7492);
xor U7610 (N_7610,N_7385,N_7465);
xnor U7611 (N_7611,N_7278,N_7319);
xnor U7612 (N_7612,N_7460,N_7497);
xnor U7613 (N_7613,N_7321,N_7330);
and U7614 (N_7614,N_7372,N_7476);
or U7615 (N_7615,N_7361,N_7389);
nand U7616 (N_7616,N_7325,N_7433);
and U7617 (N_7617,N_7298,N_7334);
or U7618 (N_7618,N_7482,N_7495);
xor U7619 (N_7619,N_7441,N_7410);
and U7620 (N_7620,N_7354,N_7421);
xnor U7621 (N_7621,N_7381,N_7496);
nand U7622 (N_7622,N_7388,N_7365);
nor U7623 (N_7623,N_7480,N_7301);
and U7624 (N_7624,N_7367,N_7427);
and U7625 (N_7625,N_7450,N_7277);
and U7626 (N_7626,N_7344,N_7376);
or U7627 (N_7627,N_7418,N_7343);
nand U7628 (N_7628,N_7412,N_7407);
nor U7629 (N_7629,N_7308,N_7432);
nor U7630 (N_7630,N_7429,N_7322);
nand U7631 (N_7631,N_7457,N_7323);
nand U7632 (N_7632,N_7251,N_7477);
and U7633 (N_7633,N_7418,N_7469);
nand U7634 (N_7634,N_7263,N_7305);
nand U7635 (N_7635,N_7373,N_7320);
and U7636 (N_7636,N_7284,N_7405);
or U7637 (N_7637,N_7270,N_7384);
nand U7638 (N_7638,N_7407,N_7319);
xor U7639 (N_7639,N_7325,N_7336);
nand U7640 (N_7640,N_7482,N_7337);
or U7641 (N_7641,N_7421,N_7411);
nor U7642 (N_7642,N_7359,N_7320);
or U7643 (N_7643,N_7379,N_7328);
nand U7644 (N_7644,N_7384,N_7390);
nor U7645 (N_7645,N_7495,N_7443);
or U7646 (N_7646,N_7297,N_7387);
xnor U7647 (N_7647,N_7496,N_7472);
nand U7648 (N_7648,N_7374,N_7347);
or U7649 (N_7649,N_7254,N_7373);
xnor U7650 (N_7650,N_7483,N_7337);
and U7651 (N_7651,N_7414,N_7499);
nand U7652 (N_7652,N_7258,N_7482);
xor U7653 (N_7653,N_7497,N_7472);
nand U7654 (N_7654,N_7496,N_7351);
nor U7655 (N_7655,N_7322,N_7413);
nand U7656 (N_7656,N_7449,N_7311);
and U7657 (N_7657,N_7314,N_7339);
xnor U7658 (N_7658,N_7376,N_7412);
nor U7659 (N_7659,N_7437,N_7471);
and U7660 (N_7660,N_7320,N_7489);
nand U7661 (N_7661,N_7390,N_7395);
nor U7662 (N_7662,N_7289,N_7434);
nor U7663 (N_7663,N_7409,N_7322);
nor U7664 (N_7664,N_7259,N_7478);
xor U7665 (N_7665,N_7286,N_7347);
nand U7666 (N_7666,N_7439,N_7462);
nand U7667 (N_7667,N_7494,N_7490);
and U7668 (N_7668,N_7426,N_7429);
xor U7669 (N_7669,N_7382,N_7337);
or U7670 (N_7670,N_7399,N_7327);
nand U7671 (N_7671,N_7313,N_7394);
nand U7672 (N_7672,N_7421,N_7446);
nor U7673 (N_7673,N_7486,N_7298);
or U7674 (N_7674,N_7271,N_7461);
and U7675 (N_7675,N_7454,N_7335);
nand U7676 (N_7676,N_7263,N_7255);
nor U7677 (N_7677,N_7368,N_7426);
nand U7678 (N_7678,N_7397,N_7269);
or U7679 (N_7679,N_7363,N_7481);
xor U7680 (N_7680,N_7436,N_7303);
or U7681 (N_7681,N_7251,N_7475);
and U7682 (N_7682,N_7339,N_7453);
nand U7683 (N_7683,N_7273,N_7316);
nor U7684 (N_7684,N_7458,N_7449);
nand U7685 (N_7685,N_7375,N_7277);
xnor U7686 (N_7686,N_7444,N_7310);
xor U7687 (N_7687,N_7367,N_7381);
and U7688 (N_7688,N_7403,N_7338);
and U7689 (N_7689,N_7417,N_7388);
nor U7690 (N_7690,N_7256,N_7475);
nor U7691 (N_7691,N_7472,N_7430);
xnor U7692 (N_7692,N_7499,N_7403);
nand U7693 (N_7693,N_7250,N_7408);
and U7694 (N_7694,N_7257,N_7348);
xor U7695 (N_7695,N_7481,N_7389);
nor U7696 (N_7696,N_7379,N_7458);
nand U7697 (N_7697,N_7386,N_7452);
and U7698 (N_7698,N_7413,N_7457);
nor U7699 (N_7699,N_7432,N_7429);
or U7700 (N_7700,N_7273,N_7402);
or U7701 (N_7701,N_7382,N_7280);
and U7702 (N_7702,N_7291,N_7448);
nand U7703 (N_7703,N_7271,N_7263);
or U7704 (N_7704,N_7446,N_7341);
xnor U7705 (N_7705,N_7386,N_7308);
and U7706 (N_7706,N_7251,N_7420);
nor U7707 (N_7707,N_7491,N_7480);
and U7708 (N_7708,N_7382,N_7342);
and U7709 (N_7709,N_7348,N_7475);
and U7710 (N_7710,N_7333,N_7273);
nor U7711 (N_7711,N_7355,N_7307);
and U7712 (N_7712,N_7420,N_7264);
or U7713 (N_7713,N_7261,N_7334);
nand U7714 (N_7714,N_7357,N_7315);
xor U7715 (N_7715,N_7310,N_7278);
and U7716 (N_7716,N_7365,N_7459);
nand U7717 (N_7717,N_7490,N_7352);
and U7718 (N_7718,N_7301,N_7442);
or U7719 (N_7719,N_7405,N_7288);
or U7720 (N_7720,N_7499,N_7259);
or U7721 (N_7721,N_7402,N_7299);
xor U7722 (N_7722,N_7490,N_7332);
and U7723 (N_7723,N_7465,N_7376);
nand U7724 (N_7724,N_7276,N_7254);
or U7725 (N_7725,N_7397,N_7494);
and U7726 (N_7726,N_7263,N_7330);
or U7727 (N_7727,N_7325,N_7467);
xor U7728 (N_7728,N_7456,N_7316);
nor U7729 (N_7729,N_7383,N_7398);
and U7730 (N_7730,N_7494,N_7475);
and U7731 (N_7731,N_7304,N_7272);
xnor U7732 (N_7732,N_7421,N_7489);
xnor U7733 (N_7733,N_7261,N_7390);
nand U7734 (N_7734,N_7301,N_7364);
and U7735 (N_7735,N_7449,N_7351);
and U7736 (N_7736,N_7319,N_7496);
or U7737 (N_7737,N_7337,N_7364);
nor U7738 (N_7738,N_7407,N_7362);
xor U7739 (N_7739,N_7450,N_7339);
nor U7740 (N_7740,N_7306,N_7419);
and U7741 (N_7741,N_7309,N_7362);
xnor U7742 (N_7742,N_7475,N_7311);
nand U7743 (N_7743,N_7324,N_7265);
and U7744 (N_7744,N_7330,N_7311);
or U7745 (N_7745,N_7316,N_7414);
and U7746 (N_7746,N_7342,N_7453);
nand U7747 (N_7747,N_7352,N_7445);
or U7748 (N_7748,N_7258,N_7430);
and U7749 (N_7749,N_7354,N_7458);
xnor U7750 (N_7750,N_7668,N_7638);
nand U7751 (N_7751,N_7653,N_7604);
and U7752 (N_7752,N_7745,N_7671);
and U7753 (N_7753,N_7590,N_7682);
xnor U7754 (N_7754,N_7571,N_7633);
nand U7755 (N_7755,N_7624,N_7570);
nand U7756 (N_7756,N_7530,N_7563);
xor U7757 (N_7757,N_7714,N_7693);
xor U7758 (N_7758,N_7615,N_7596);
nand U7759 (N_7759,N_7729,N_7584);
and U7760 (N_7760,N_7709,N_7674);
xnor U7761 (N_7761,N_7538,N_7575);
or U7762 (N_7762,N_7737,N_7514);
xor U7763 (N_7763,N_7646,N_7690);
or U7764 (N_7764,N_7577,N_7702);
and U7765 (N_7765,N_7661,N_7708);
nor U7766 (N_7766,N_7659,N_7566);
nand U7767 (N_7767,N_7618,N_7545);
nor U7768 (N_7768,N_7552,N_7664);
nand U7769 (N_7769,N_7516,N_7723);
nand U7770 (N_7770,N_7724,N_7645);
nand U7771 (N_7771,N_7573,N_7713);
or U7772 (N_7772,N_7539,N_7603);
or U7773 (N_7773,N_7707,N_7512);
nor U7774 (N_7774,N_7543,N_7678);
nand U7775 (N_7775,N_7533,N_7697);
or U7776 (N_7776,N_7675,N_7601);
or U7777 (N_7777,N_7625,N_7511);
xor U7778 (N_7778,N_7680,N_7711);
xnor U7779 (N_7779,N_7598,N_7647);
and U7780 (N_7780,N_7715,N_7666);
nand U7781 (N_7781,N_7613,N_7597);
nand U7782 (N_7782,N_7560,N_7704);
or U7783 (N_7783,N_7576,N_7643);
nand U7784 (N_7784,N_7607,N_7502);
or U7785 (N_7785,N_7578,N_7529);
nor U7786 (N_7786,N_7510,N_7665);
xor U7787 (N_7787,N_7669,N_7734);
xor U7788 (N_7788,N_7691,N_7574);
nor U7789 (N_7789,N_7507,N_7522);
nand U7790 (N_7790,N_7684,N_7585);
nor U7791 (N_7791,N_7655,N_7687);
xnor U7792 (N_7792,N_7670,N_7717);
and U7793 (N_7793,N_7733,N_7619);
or U7794 (N_7794,N_7605,N_7629);
nor U7795 (N_7795,N_7739,N_7599);
and U7796 (N_7796,N_7548,N_7551);
xnor U7797 (N_7797,N_7520,N_7531);
nor U7798 (N_7798,N_7586,N_7589);
xor U7799 (N_7799,N_7528,N_7663);
nand U7800 (N_7800,N_7611,N_7628);
and U7801 (N_7801,N_7747,N_7626);
and U7802 (N_7802,N_7698,N_7549);
nand U7803 (N_7803,N_7642,N_7662);
nand U7804 (N_7804,N_7641,N_7537);
nand U7805 (N_7805,N_7622,N_7705);
and U7806 (N_7806,N_7741,N_7583);
nand U7807 (N_7807,N_7716,N_7559);
or U7808 (N_7808,N_7746,N_7656);
xnor U7809 (N_7809,N_7620,N_7710);
or U7810 (N_7810,N_7644,N_7561);
xor U7811 (N_7811,N_7683,N_7534);
xor U7812 (N_7812,N_7701,N_7685);
and U7813 (N_7813,N_7621,N_7558);
and U7814 (N_7814,N_7593,N_7676);
and U7815 (N_7815,N_7692,N_7677);
nor U7816 (N_7816,N_7540,N_7544);
xor U7817 (N_7817,N_7667,N_7634);
nand U7818 (N_7818,N_7550,N_7536);
xor U7819 (N_7819,N_7648,N_7719);
and U7820 (N_7820,N_7727,N_7695);
nor U7821 (N_7821,N_7735,N_7616);
and U7822 (N_7822,N_7562,N_7681);
and U7823 (N_7823,N_7654,N_7588);
nor U7824 (N_7824,N_7527,N_7553);
xnor U7825 (N_7825,N_7700,N_7532);
or U7826 (N_7826,N_7631,N_7632);
xor U7827 (N_7827,N_7658,N_7696);
or U7828 (N_7828,N_7580,N_7595);
nor U7829 (N_7829,N_7689,N_7627);
nand U7830 (N_7830,N_7743,N_7657);
nor U7831 (N_7831,N_7703,N_7509);
nor U7832 (N_7832,N_7694,N_7554);
nand U7833 (N_7833,N_7649,N_7592);
xnor U7834 (N_7834,N_7606,N_7521);
nand U7835 (N_7835,N_7660,N_7567);
xor U7836 (N_7836,N_7636,N_7672);
xnor U7837 (N_7837,N_7718,N_7722);
nand U7838 (N_7838,N_7579,N_7503);
nand U7839 (N_7839,N_7526,N_7736);
xnor U7840 (N_7840,N_7508,N_7635);
nand U7841 (N_7841,N_7639,N_7673);
and U7842 (N_7842,N_7744,N_7731);
nor U7843 (N_7843,N_7608,N_7651);
nor U7844 (N_7844,N_7738,N_7581);
nor U7845 (N_7845,N_7504,N_7517);
and U7846 (N_7846,N_7557,N_7501);
nor U7847 (N_7847,N_7712,N_7609);
xor U7848 (N_7848,N_7728,N_7612);
or U7849 (N_7849,N_7568,N_7515);
xnor U7850 (N_7850,N_7600,N_7519);
or U7851 (N_7851,N_7518,N_7748);
nor U7852 (N_7852,N_7555,N_7740);
xor U7853 (N_7853,N_7594,N_7686);
nor U7854 (N_7854,N_7602,N_7524);
xnor U7855 (N_7855,N_7556,N_7564);
nor U7856 (N_7856,N_7706,N_7505);
nor U7857 (N_7857,N_7725,N_7742);
nand U7858 (N_7858,N_7587,N_7525);
or U7859 (N_7859,N_7640,N_7688);
and U7860 (N_7860,N_7650,N_7617);
nor U7861 (N_7861,N_7535,N_7726);
nor U7862 (N_7862,N_7721,N_7591);
nor U7863 (N_7863,N_7732,N_7523);
xnor U7864 (N_7864,N_7749,N_7630);
nor U7865 (N_7865,N_7614,N_7699);
and U7866 (N_7866,N_7547,N_7546);
nor U7867 (N_7867,N_7679,N_7582);
nor U7868 (N_7868,N_7637,N_7506);
nor U7869 (N_7869,N_7513,N_7541);
nor U7870 (N_7870,N_7610,N_7730);
nor U7871 (N_7871,N_7542,N_7565);
and U7872 (N_7872,N_7500,N_7652);
nor U7873 (N_7873,N_7720,N_7569);
nor U7874 (N_7874,N_7623,N_7572);
and U7875 (N_7875,N_7719,N_7536);
nor U7876 (N_7876,N_7641,N_7613);
or U7877 (N_7877,N_7590,N_7568);
and U7878 (N_7878,N_7650,N_7571);
and U7879 (N_7879,N_7624,N_7733);
and U7880 (N_7880,N_7621,N_7716);
nand U7881 (N_7881,N_7587,N_7536);
xor U7882 (N_7882,N_7501,N_7697);
or U7883 (N_7883,N_7642,N_7617);
nand U7884 (N_7884,N_7732,N_7621);
nand U7885 (N_7885,N_7677,N_7691);
xor U7886 (N_7886,N_7627,N_7613);
or U7887 (N_7887,N_7683,N_7749);
and U7888 (N_7888,N_7537,N_7505);
or U7889 (N_7889,N_7665,N_7629);
and U7890 (N_7890,N_7661,N_7572);
nand U7891 (N_7891,N_7734,N_7708);
xor U7892 (N_7892,N_7565,N_7549);
xnor U7893 (N_7893,N_7640,N_7636);
and U7894 (N_7894,N_7508,N_7523);
nor U7895 (N_7895,N_7624,N_7668);
and U7896 (N_7896,N_7571,N_7720);
or U7897 (N_7897,N_7546,N_7617);
xnor U7898 (N_7898,N_7503,N_7632);
xnor U7899 (N_7899,N_7712,N_7711);
nand U7900 (N_7900,N_7681,N_7585);
xnor U7901 (N_7901,N_7661,N_7696);
nand U7902 (N_7902,N_7645,N_7569);
or U7903 (N_7903,N_7519,N_7652);
nor U7904 (N_7904,N_7516,N_7738);
and U7905 (N_7905,N_7599,N_7681);
nand U7906 (N_7906,N_7552,N_7733);
and U7907 (N_7907,N_7657,N_7683);
and U7908 (N_7908,N_7604,N_7681);
xor U7909 (N_7909,N_7521,N_7693);
and U7910 (N_7910,N_7611,N_7526);
xnor U7911 (N_7911,N_7552,N_7641);
or U7912 (N_7912,N_7628,N_7631);
nand U7913 (N_7913,N_7572,N_7543);
and U7914 (N_7914,N_7530,N_7515);
or U7915 (N_7915,N_7527,N_7572);
and U7916 (N_7916,N_7655,N_7595);
xor U7917 (N_7917,N_7717,N_7671);
and U7918 (N_7918,N_7524,N_7668);
and U7919 (N_7919,N_7669,N_7598);
nand U7920 (N_7920,N_7640,N_7520);
nor U7921 (N_7921,N_7519,N_7511);
and U7922 (N_7922,N_7512,N_7554);
and U7923 (N_7923,N_7587,N_7531);
xor U7924 (N_7924,N_7720,N_7738);
nand U7925 (N_7925,N_7726,N_7677);
xnor U7926 (N_7926,N_7746,N_7504);
nor U7927 (N_7927,N_7675,N_7740);
xor U7928 (N_7928,N_7626,N_7736);
or U7929 (N_7929,N_7657,N_7677);
nor U7930 (N_7930,N_7505,N_7715);
nor U7931 (N_7931,N_7545,N_7549);
xnor U7932 (N_7932,N_7618,N_7562);
xor U7933 (N_7933,N_7735,N_7731);
or U7934 (N_7934,N_7582,N_7638);
or U7935 (N_7935,N_7729,N_7549);
nor U7936 (N_7936,N_7603,N_7637);
nand U7937 (N_7937,N_7539,N_7708);
and U7938 (N_7938,N_7725,N_7674);
nor U7939 (N_7939,N_7639,N_7637);
nand U7940 (N_7940,N_7587,N_7533);
nand U7941 (N_7941,N_7733,N_7725);
or U7942 (N_7942,N_7602,N_7696);
or U7943 (N_7943,N_7681,N_7655);
nor U7944 (N_7944,N_7603,N_7560);
or U7945 (N_7945,N_7618,N_7517);
xor U7946 (N_7946,N_7539,N_7611);
nand U7947 (N_7947,N_7586,N_7692);
nor U7948 (N_7948,N_7626,N_7593);
xor U7949 (N_7949,N_7722,N_7709);
xor U7950 (N_7950,N_7506,N_7527);
nand U7951 (N_7951,N_7606,N_7628);
and U7952 (N_7952,N_7616,N_7530);
or U7953 (N_7953,N_7645,N_7524);
nand U7954 (N_7954,N_7637,N_7711);
xnor U7955 (N_7955,N_7672,N_7736);
or U7956 (N_7956,N_7629,N_7630);
xor U7957 (N_7957,N_7574,N_7593);
nand U7958 (N_7958,N_7555,N_7560);
nor U7959 (N_7959,N_7610,N_7546);
xnor U7960 (N_7960,N_7615,N_7695);
nor U7961 (N_7961,N_7735,N_7673);
and U7962 (N_7962,N_7679,N_7504);
and U7963 (N_7963,N_7675,N_7606);
or U7964 (N_7964,N_7737,N_7511);
nor U7965 (N_7965,N_7657,N_7553);
or U7966 (N_7966,N_7503,N_7606);
nor U7967 (N_7967,N_7669,N_7621);
or U7968 (N_7968,N_7655,N_7677);
and U7969 (N_7969,N_7661,N_7640);
or U7970 (N_7970,N_7600,N_7545);
nor U7971 (N_7971,N_7709,N_7622);
nand U7972 (N_7972,N_7655,N_7599);
xnor U7973 (N_7973,N_7672,N_7537);
and U7974 (N_7974,N_7520,N_7576);
nor U7975 (N_7975,N_7583,N_7512);
and U7976 (N_7976,N_7525,N_7576);
xnor U7977 (N_7977,N_7507,N_7540);
or U7978 (N_7978,N_7621,N_7685);
and U7979 (N_7979,N_7700,N_7637);
or U7980 (N_7980,N_7690,N_7549);
and U7981 (N_7981,N_7634,N_7646);
nand U7982 (N_7982,N_7704,N_7613);
xor U7983 (N_7983,N_7693,N_7568);
and U7984 (N_7984,N_7532,N_7606);
nor U7985 (N_7985,N_7605,N_7708);
and U7986 (N_7986,N_7591,N_7580);
xor U7987 (N_7987,N_7684,N_7540);
or U7988 (N_7988,N_7744,N_7723);
nor U7989 (N_7989,N_7690,N_7746);
nor U7990 (N_7990,N_7525,N_7636);
or U7991 (N_7991,N_7615,N_7733);
nor U7992 (N_7992,N_7516,N_7663);
xnor U7993 (N_7993,N_7679,N_7659);
and U7994 (N_7994,N_7618,N_7715);
and U7995 (N_7995,N_7691,N_7737);
xor U7996 (N_7996,N_7575,N_7623);
and U7997 (N_7997,N_7571,N_7676);
or U7998 (N_7998,N_7632,N_7639);
xnor U7999 (N_7999,N_7555,N_7520);
xnor U8000 (N_8000,N_7884,N_7869);
nand U8001 (N_8001,N_7906,N_7927);
xnor U8002 (N_8002,N_7892,N_7820);
nor U8003 (N_8003,N_7982,N_7834);
nor U8004 (N_8004,N_7940,N_7826);
and U8005 (N_8005,N_7770,N_7885);
xor U8006 (N_8006,N_7909,N_7833);
or U8007 (N_8007,N_7903,N_7784);
nand U8008 (N_8008,N_7808,N_7935);
or U8009 (N_8009,N_7998,N_7866);
or U8010 (N_8010,N_7835,N_7943);
xor U8011 (N_8011,N_7783,N_7968);
nor U8012 (N_8012,N_7865,N_7750);
nor U8013 (N_8013,N_7953,N_7924);
nor U8014 (N_8014,N_7776,N_7999);
nor U8015 (N_8015,N_7842,N_7972);
or U8016 (N_8016,N_7923,N_7961);
and U8017 (N_8017,N_7901,N_7821);
xnor U8018 (N_8018,N_7837,N_7775);
nor U8019 (N_8019,N_7828,N_7771);
xor U8020 (N_8020,N_7929,N_7868);
nor U8021 (N_8021,N_7899,N_7755);
or U8022 (N_8022,N_7862,N_7894);
or U8023 (N_8023,N_7763,N_7993);
or U8024 (N_8024,N_7988,N_7867);
and U8025 (N_8025,N_7874,N_7839);
xor U8026 (N_8026,N_7814,N_7823);
and U8027 (N_8027,N_7804,N_7945);
or U8028 (N_8028,N_7829,N_7857);
xor U8029 (N_8029,N_7764,N_7794);
xnor U8030 (N_8030,N_7791,N_7864);
nor U8031 (N_8031,N_7856,N_7926);
or U8032 (N_8032,N_7948,N_7802);
xor U8033 (N_8033,N_7956,N_7778);
and U8034 (N_8034,N_7836,N_7878);
nand U8035 (N_8035,N_7855,N_7819);
nand U8036 (N_8036,N_7942,N_7800);
nor U8037 (N_8037,N_7782,N_7922);
or U8038 (N_8038,N_7936,N_7805);
xor U8039 (N_8039,N_7958,N_7777);
nor U8040 (N_8040,N_7832,N_7824);
or U8041 (N_8041,N_7877,N_7807);
xor U8042 (N_8042,N_7902,N_7853);
nand U8043 (N_8043,N_7930,N_7838);
or U8044 (N_8044,N_7786,N_7761);
nor U8045 (N_8045,N_7919,N_7847);
and U8046 (N_8046,N_7983,N_7974);
nor U8047 (N_8047,N_7986,N_7887);
or U8048 (N_8048,N_7787,N_7947);
xnor U8049 (N_8049,N_7789,N_7995);
nor U8050 (N_8050,N_7852,N_7818);
xor U8051 (N_8051,N_7825,N_7910);
nor U8052 (N_8052,N_7960,N_7872);
or U8053 (N_8053,N_7871,N_7753);
and U8054 (N_8054,N_7812,N_7848);
or U8055 (N_8055,N_7756,N_7827);
or U8056 (N_8056,N_7859,N_7883);
nand U8057 (N_8057,N_7815,N_7937);
nand U8058 (N_8058,N_7831,N_7767);
xor U8059 (N_8059,N_7946,N_7944);
and U8060 (N_8060,N_7758,N_7914);
nor U8061 (N_8061,N_7788,N_7760);
nand U8062 (N_8062,N_7966,N_7898);
and U8063 (N_8063,N_7939,N_7907);
or U8064 (N_8064,N_7978,N_7762);
xnor U8065 (N_8065,N_7766,N_7931);
xor U8066 (N_8066,N_7759,N_7880);
xor U8067 (N_8067,N_7964,N_7941);
nand U8068 (N_8068,N_7895,N_7987);
nor U8069 (N_8069,N_7854,N_7769);
or U8070 (N_8070,N_7757,N_7792);
nor U8071 (N_8071,N_7979,N_7888);
nor U8072 (N_8072,N_7840,N_7845);
xor U8073 (N_8073,N_7793,N_7809);
nand U8074 (N_8074,N_7882,N_7990);
and U8075 (N_8075,N_7900,N_7773);
nor U8076 (N_8076,N_7918,N_7870);
nand U8077 (N_8077,N_7886,N_7967);
or U8078 (N_8078,N_7774,N_7846);
or U8079 (N_8079,N_7992,N_7861);
and U8080 (N_8080,N_7781,N_7973);
or U8081 (N_8081,N_7904,N_7772);
nand U8082 (N_8082,N_7822,N_7799);
and U8083 (N_8083,N_7932,N_7908);
or U8084 (N_8084,N_7976,N_7949);
nor U8085 (N_8085,N_7984,N_7905);
xnor U8086 (N_8086,N_7765,N_7754);
and U8087 (N_8087,N_7876,N_7938);
or U8088 (N_8088,N_7963,N_7893);
xnor U8089 (N_8089,N_7801,N_7841);
nand U8090 (N_8090,N_7994,N_7981);
nor U8091 (N_8091,N_7969,N_7913);
xor U8092 (N_8092,N_7752,N_7875);
xnor U8093 (N_8093,N_7790,N_7957);
and U8094 (N_8094,N_7915,N_7965);
or U8095 (N_8095,N_7795,N_7817);
xor U8096 (N_8096,N_7985,N_7851);
nor U8097 (N_8097,N_7879,N_7934);
and U8098 (N_8098,N_7813,N_7850);
xor U8099 (N_8099,N_7844,N_7933);
and U8100 (N_8100,N_7810,N_7811);
or U8101 (N_8101,N_7977,N_7971);
or U8102 (N_8102,N_7950,N_7989);
nand U8103 (N_8103,N_7768,N_7996);
or U8104 (N_8104,N_7816,N_7975);
nor U8105 (N_8105,N_7916,N_7779);
nor U8106 (N_8106,N_7997,N_7803);
nand U8107 (N_8107,N_7925,N_7912);
nor U8108 (N_8108,N_7920,N_7928);
or U8109 (N_8109,N_7921,N_7860);
or U8110 (N_8110,N_7785,N_7889);
nor U8111 (N_8111,N_7991,N_7891);
nand U8112 (N_8112,N_7780,N_7896);
nand U8113 (N_8113,N_7751,N_7980);
or U8114 (N_8114,N_7951,N_7873);
or U8115 (N_8115,N_7806,N_7952);
nand U8116 (N_8116,N_7970,N_7830);
or U8117 (N_8117,N_7911,N_7863);
or U8118 (N_8118,N_7881,N_7843);
nand U8119 (N_8119,N_7849,N_7959);
xnor U8120 (N_8120,N_7890,N_7796);
or U8121 (N_8121,N_7858,N_7917);
and U8122 (N_8122,N_7955,N_7797);
nor U8123 (N_8123,N_7962,N_7798);
nor U8124 (N_8124,N_7897,N_7954);
xor U8125 (N_8125,N_7778,N_7864);
and U8126 (N_8126,N_7900,N_7858);
or U8127 (N_8127,N_7766,N_7923);
or U8128 (N_8128,N_7950,N_7893);
xnor U8129 (N_8129,N_7869,N_7909);
xnor U8130 (N_8130,N_7975,N_7830);
xnor U8131 (N_8131,N_7923,N_7904);
nand U8132 (N_8132,N_7869,N_7949);
or U8133 (N_8133,N_7995,N_7827);
xnor U8134 (N_8134,N_7880,N_7936);
or U8135 (N_8135,N_7948,N_7882);
nor U8136 (N_8136,N_7908,N_7897);
xor U8137 (N_8137,N_7902,N_7966);
nor U8138 (N_8138,N_7934,N_7913);
nor U8139 (N_8139,N_7773,N_7958);
or U8140 (N_8140,N_7811,N_7921);
or U8141 (N_8141,N_7764,N_7901);
nor U8142 (N_8142,N_7879,N_7980);
nand U8143 (N_8143,N_7913,N_7928);
nor U8144 (N_8144,N_7897,N_7764);
and U8145 (N_8145,N_7967,N_7806);
or U8146 (N_8146,N_7851,N_7899);
or U8147 (N_8147,N_7999,N_7859);
xnor U8148 (N_8148,N_7869,N_7854);
or U8149 (N_8149,N_7842,N_7829);
or U8150 (N_8150,N_7952,N_7914);
and U8151 (N_8151,N_7957,N_7857);
nand U8152 (N_8152,N_7832,N_7826);
and U8153 (N_8153,N_7955,N_7916);
and U8154 (N_8154,N_7889,N_7971);
nand U8155 (N_8155,N_7847,N_7771);
and U8156 (N_8156,N_7793,N_7831);
and U8157 (N_8157,N_7860,N_7875);
and U8158 (N_8158,N_7906,N_7751);
nor U8159 (N_8159,N_7934,N_7892);
nor U8160 (N_8160,N_7806,N_7790);
nor U8161 (N_8161,N_7856,N_7915);
nor U8162 (N_8162,N_7858,N_7874);
nand U8163 (N_8163,N_7772,N_7821);
nand U8164 (N_8164,N_7926,N_7763);
xnor U8165 (N_8165,N_7837,N_7984);
or U8166 (N_8166,N_7961,N_7939);
nor U8167 (N_8167,N_7851,N_7951);
nor U8168 (N_8168,N_7986,N_7928);
nor U8169 (N_8169,N_7833,N_7871);
xnor U8170 (N_8170,N_7926,N_7914);
nor U8171 (N_8171,N_7948,N_7763);
or U8172 (N_8172,N_7970,N_7802);
or U8173 (N_8173,N_7982,N_7778);
nor U8174 (N_8174,N_7910,N_7904);
nor U8175 (N_8175,N_7796,N_7955);
or U8176 (N_8176,N_7960,N_7940);
nand U8177 (N_8177,N_7872,N_7911);
nor U8178 (N_8178,N_7930,N_7807);
xnor U8179 (N_8179,N_7815,N_7956);
nand U8180 (N_8180,N_7908,N_7759);
or U8181 (N_8181,N_7894,N_7831);
nand U8182 (N_8182,N_7855,N_7829);
xnor U8183 (N_8183,N_7861,N_7796);
nor U8184 (N_8184,N_7973,N_7942);
or U8185 (N_8185,N_7963,N_7793);
and U8186 (N_8186,N_7871,N_7928);
nor U8187 (N_8187,N_7914,N_7821);
and U8188 (N_8188,N_7768,N_7928);
xnor U8189 (N_8189,N_7911,N_7993);
nand U8190 (N_8190,N_7786,N_7952);
nand U8191 (N_8191,N_7922,N_7910);
and U8192 (N_8192,N_7822,N_7971);
nor U8193 (N_8193,N_7789,N_7772);
nor U8194 (N_8194,N_7861,N_7957);
or U8195 (N_8195,N_7901,N_7878);
nand U8196 (N_8196,N_7781,N_7986);
and U8197 (N_8197,N_7996,N_7759);
and U8198 (N_8198,N_7806,N_7785);
and U8199 (N_8199,N_7859,N_7761);
and U8200 (N_8200,N_7960,N_7964);
and U8201 (N_8201,N_7880,N_7997);
and U8202 (N_8202,N_7951,N_7781);
nor U8203 (N_8203,N_7784,N_7890);
and U8204 (N_8204,N_7887,N_7978);
or U8205 (N_8205,N_7836,N_7904);
or U8206 (N_8206,N_7878,N_7876);
and U8207 (N_8207,N_7799,N_7857);
xnor U8208 (N_8208,N_7829,N_7971);
nor U8209 (N_8209,N_7900,N_7791);
nor U8210 (N_8210,N_7984,N_7763);
nor U8211 (N_8211,N_7805,N_7782);
nand U8212 (N_8212,N_7897,N_7936);
and U8213 (N_8213,N_7910,N_7756);
xnor U8214 (N_8214,N_7940,N_7859);
and U8215 (N_8215,N_7943,N_7760);
and U8216 (N_8216,N_7926,N_7866);
xor U8217 (N_8217,N_7983,N_7864);
or U8218 (N_8218,N_7854,N_7860);
or U8219 (N_8219,N_7963,N_7980);
nor U8220 (N_8220,N_7921,N_7898);
nand U8221 (N_8221,N_7997,N_7780);
nand U8222 (N_8222,N_7801,N_7810);
nand U8223 (N_8223,N_7993,N_7794);
nand U8224 (N_8224,N_7939,N_7947);
xnor U8225 (N_8225,N_7886,N_7840);
nor U8226 (N_8226,N_7865,N_7891);
or U8227 (N_8227,N_7762,N_7992);
xor U8228 (N_8228,N_7976,N_7924);
and U8229 (N_8229,N_7871,N_7801);
nand U8230 (N_8230,N_7843,N_7913);
nand U8231 (N_8231,N_7775,N_7777);
nor U8232 (N_8232,N_7966,N_7844);
nor U8233 (N_8233,N_7975,N_7787);
or U8234 (N_8234,N_7903,N_7763);
and U8235 (N_8235,N_7787,N_7846);
and U8236 (N_8236,N_7750,N_7913);
xnor U8237 (N_8237,N_7908,N_7771);
nand U8238 (N_8238,N_7895,N_7841);
nand U8239 (N_8239,N_7863,N_7774);
nand U8240 (N_8240,N_7822,N_7910);
or U8241 (N_8241,N_7876,N_7754);
and U8242 (N_8242,N_7969,N_7880);
nor U8243 (N_8243,N_7880,N_7830);
or U8244 (N_8244,N_7757,N_7875);
nor U8245 (N_8245,N_7918,N_7828);
xor U8246 (N_8246,N_7907,N_7777);
xor U8247 (N_8247,N_7843,N_7902);
nand U8248 (N_8248,N_7964,N_7764);
nor U8249 (N_8249,N_7842,N_7780);
nor U8250 (N_8250,N_8062,N_8073);
nor U8251 (N_8251,N_8232,N_8015);
nor U8252 (N_8252,N_8112,N_8025);
or U8253 (N_8253,N_8128,N_8008);
or U8254 (N_8254,N_8225,N_8198);
nor U8255 (N_8255,N_8194,N_8144);
nand U8256 (N_8256,N_8040,N_8204);
nand U8257 (N_8257,N_8108,N_8099);
and U8258 (N_8258,N_8067,N_8104);
or U8259 (N_8259,N_8130,N_8024);
nand U8260 (N_8260,N_8029,N_8012);
xnor U8261 (N_8261,N_8120,N_8164);
xnor U8262 (N_8262,N_8131,N_8246);
and U8263 (N_8263,N_8205,N_8145);
xnor U8264 (N_8264,N_8081,N_8002);
nand U8265 (N_8265,N_8054,N_8213);
xnor U8266 (N_8266,N_8179,N_8058);
and U8267 (N_8267,N_8001,N_8110);
nor U8268 (N_8268,N_8178,N_8132);
or U8269 (N_8269,N_8052,N_8079);
and U8270 (N_8270,N_8028,N_8239);
nor U8271 (N_8271,N_8244,N_8191);
xor U8272 (N_8272,N_8103,N_8173);
and U8273 (N_8273,N_8048,N_8053);
or U8274 (N_8274,N_8060,N_8165);
and U8275 (N_8275,N_8220,N_8169);
or U8276 (N_8276,N_8193,N_8206);
or U8277 (N_8277,N_8139,N_8214);
xor U8278 (N_8278,N_8095,N_8227);
or U8279 (N_8279,N_8037,N_8223);
or U8280 (N_8280,N_8107,N_8159);
and U8281 (N_8281,N_8155,N_8197);
nor U8282 (N_8282,N_8007,N_8189);
and U8283 (N_8283,N_8069,N_8170);
nand U8284 (N_8284,N_8013,N_8055);
nand U8285 (N_8285,N_8188,N_8044);
or U8286 (N_8286,N_8071,N_8074);
and U8287 (N_8287,N_8219,N_8038);
or U8288 (N_8288,N_8195,N_8090);
xor U8289 (N_8289,N_8160,N_8226);
or U8290 (N_8290,N_8249,N_8163);
nand U8291 (N_8291,N_8100,N_8118);
xnor U8292 (N_8292,N_8143,N_8003);
nand U8293 (N_8293,N_8089,N_8136);
nor U8294 (N_8294,N_8199,N_8083);
nand U8295 (N_8295,N_8150,N_8004);
xnor U8296 (N_8296,N_8210,N_8190);
nor U8297 (N_8297,N_8183,N_8092);
xor U8298 (N_8298,N_8181,N_8233);
and U8299 (N_8299,N_8010,N_8063);
xor U8300 (N_8300,N_8031,N_8148);
nor U8301 (N_8301,N_8072,N_8192);
and U8302 (N_8302,N_8149,N_8114);
or U8303 (N_8303,N_8140,N_8006);
or U8304 (N_8304,N_8151,N_8243);
and U8305 (N_8305,N_8236,N_8093);
nand U8306 (N_8306,N_8098,N_8000);
nor U8307 (N_8307,N_8124,N_8125);
nand U8308 (N_8308,N_8018,N_8147);
or U8309 (N_8309,N_8047,N_8202);
xnor U8310 (N_8310,N_8126,N_8096);
and U8311 (N_8311,N_8056,N_8157);
and U8312 (N_8312,N_8156,N_8014);
or U8313 (N_8313,N_8033,N_8230);
xor U8314 (N_8314,N_8011,N_8215);
or U8315 (N_8315,N_8138,N_8167);
nor U8316 (N_8316,N_8184,N_8051);
nand U8317 (N_8317,N_8080,N_8211);
nand U8318 (N_8318,N_8091,N_8087);
xor U8319 (N_8319,N_8041,N_8050);
or U8320 (N_8320,N_8088,N_8201);
and U8321 (N_8321,N_8222,N_8224);
xnor U8322 (N_8322,N_8158,N_8036);
nand U8323 (N_8323,N_8027,N_8123);
nor U8324 (N_8324,N_8049,N_8039);
or U8325 (N_8325,N_8186,N_8129);
xor U8326 (N_8326,N_8086,N_8177);
nor U8327 (N_8327,N_8133,N_8046);
nor U8328 (N_8328,N_8117,N_8111);
nand U8329 (N_8329,N_8161,N_8017);
or U8330 (N_8330,N_8097,N_8042);
and U8331 (N_8331,N_8078,N_8187);
xor U8332 (N_8332,N_8005,N_8141);
xor U8333 (N_8333,N_8105,N_8020);
nand U8334 (N_8334,N_8035,N_8221);
or U8335 (N_8335,N_8016,N_8043);
nand U8336 (N_8336,N_8142,N_8009);
nor U8337 (N_8337,N_8061,N_8106);
and U8338 (N_8338,N_8030,N_8241);
and U8339 (N_8339,N_8085,N_8162);
and U8340 (N_8340,N_8127,N_8166);
nor U8341 (N_8341,N_8076,N_8176);
xnor U8342 (N_8342,N_8135,N_8152);
nand U8343 (N_8343,N_8084,N_8153);
and U8344 (N_8344,N_8137,N_8168);
xnor U8345 (N_8345,N_8175,N_8229);
nor U8346 (N_8346,N_8200,N_8216);
nand U8347 (N_8347,N_8245,N_8077);
nor U8348 (N_8348,N_8231,N_8154);
xnor U8349 (N_8349,N_8174,N_8057);
and U8350 (N_8350,N_8208,N_8237);
nor U8351 (N_8351,N_8109,N_8116);
nand U8352 (N_8352,N_8068,N_8026);
nand U8353 (N_8353,N_8066,N_8121);
and U8354 (N_8354,N_8242,N_8235);
and U8355 (N_8355,N_8115,N_8022);
xor U8356 (N_8356,N_8146,N_8059);
or U8357 (N_8357,N_8238,N_8034);
nand U8358 (N_8358,N_8172,N_8212);
nor U8359 (N_8359,N_8021,N_8171);
nor U8360 (N_8360,N_8064,N_8228);
or U8361 (N_8361,N_8185,N_8102);
xnor U8362 (N_8362,N_8180,N_8248);
or U8363 (N_8363,N_8203,N_8075);
xnor U8364 (N_8364,N_8209,N_8234);
or U8365 (N_8365,N_8134,N_8019);
xor U8366 (N_8366,N_8032,N_8101);
nor U8367 (N_8367,N_8113,N_8247);
or U8368 (N_8368,N_8182,N_8196);
or U8369 (N_8369,N_8240,N_8082);
nor U8370 (N_8370,N_8122,N_8094);
and U8371 (N_8371,N_8119,N_8045);
or U8372 (N_8372,N_8207,N_8065);
nand U8373 (N_8373,N_8070,N_8023);
nand U8374 (N_8374,N_8218,N_8217);
nor U8375 (N_8375,N_8093,N_8231);
nand U8376 (N_8376,N_8176,N_8077);
nand U8377 (N_8377,N_8233,N_8170);
or U8378 (N_8378,N_8141,N_8154);
nor U8379 (N_8379,N_8153,N_8108);
nor U8380 (N_8380,N_8127,N_8110);
or U8381 (N_8381,N_8026,N_8086);
nor U8382 (N_8382,N_8106,N_8033);
xor U8383 (N_8383,N_8234,N_8238);
nand U8384 (N_8384,N_8093,N_8006);
and U8385 (N_8385,N_8179,N_8184);
nand U8386 (N_8386,N_8119,N_8065);
nor U8387 (N_8387,N_8100,N_8007);
nor U8388 (N_8388,N_8024,N_8017);
xor U8389 (N_8389,N_8239,N_8223);
nor U8390 (N_8390,N_8080,N_8221);
or U8391 (N_8391,N_8009,N_8228);
or U8392 (N_8392,N_8166,N_8237);
or U8393 (N_8393,N_8045,N_8204);
and U8394 (N_8394,N_8139,N_8187);
or U8395 (N_8395,N_8077,N_8199);
and U8396 (N_8396,N_8032,N_8044);
or U8397 (N_8397,N_8114,N_8235);
and U8398 (N_8398,N_8235,N_8045);
and U8399 (N_8399,N_8222,N_8022);
and U8400 (N_8400,N_8215,N_8026);
xor U8401 (N_8401,N_8121,N_8015);
xor U8402 (N_8402,N_8143,N_8108);
and U8403 (N_8403,N_8052,N_8043);
xor U8404 (N_8404,N_8199,N_8025);
or U8405 (N_8405,N_8097,N_8199);
xor U8406 (N_8406,N_8142,N_8051);
xor U8407 (N_8407,N_8169,N_8226);
xor U8408 (N_8408,N_8035,N_8069);
or U8409 (N_8409,N_8052,N_8180);
nand U8410 (N_8410,N_8228,N_8080);
nor U8411 (N_8411,N_8046,N_8080);
and U8412 (N_8412,N_8210,N_8128);
xnor U8413 (N_8413,N_8051,N_8054);
xor U8414 (N_8414,N_8109,N_8095);
nor U8415 (N_8415,N_8141,N_8008);
nand U8416 (N_8416,N_8194,N_8021);
or U8417 (N_8417,N_8102,N_8249);
or U8418 (N_8418,N_8155,N_8093);
or U8419 (N_8419,N_8057,N_8126);
and U8420 (N_8420,N_8092,N_8189);
xor U8421 (N_8421,N_8028,N_8031);
nor U8422 (N_8422,N_8106,N_8035);
or U8423 (N_8423,N_8161,N_8053);
xnor U8424 (N_8424,N_8051,N_8165);
nor U8425 (N_8425,N_8142,N_8130);
nor U8426 (N_8426,N_8155,N_8070);
nor U8427 (N_8427,N_8024,N_8179);
and U8428 (N_8428,N_8114,N_8098);
nor U8429 (N_8429,N_8198,N_8234);
nand U8430 (N_8430,N_8054,N_8108);
or U8431 (N_8431,N_8202,N_8025);
xnor U8432 (N_8432,N_8082,N_8015);
or U8433 (N_8433,N_8228,N_8103);
or U8434 (N_8434,N_8085,N_8053);
xor U8435 (N_8435,N_8192,N_8165);
nand U8436 (N_8436,N_8114,N_8060);
or U8437 (N_8437,N_8079,N_8049);
nor U8438 (N_8438,N_8089,N_8162);
and U8439 (N_8439,N_8042,N_8071);
nor U8440 (N_8440,N_8079,N_8016);
nor U8441 (N_8441,N_8239,N_8065);
nand U8442 (N_8442,N_8203,N_8164);
nand U8443 (N_8443,N_8194,N_8009);
and U8444 (N_8444,N_8147,N_8061);
nor U8445 (N_8445,N_8196,N_8088);
or U8446 (N_8446,N_8075,N_8150);
or U8447 (N_8447,N_8107,N_8152);
nand U8448 (N_8448,N_8087,N_8078);
or U8449 (N_8449,N_8110,N_8169);
and U8450 (N_8450,N_8196,N_8133);
or U8451 (N_8451,N_8158,N_8127);
xnor U8452 (N_8452,N_8163,N_8115);
or U8453 (N_8453,N_8065,N_8125);
xor U8454 (N_8454,N_8094,N_8222);
nor U8455 (N_8455,N_8216,N_8014);
and U8456 (N_8456,N_8124,N_8205);
xor U8457 (N_8457,N_8150,N_8129);
nand U8458 (N_8458,N_8239,N_8182);
xor U8459 (N_8459,N_8082,N_8017);
nor U8460 (N_8460,N_8186,N_8246);
or U8461 (N_8461,N_8040,N_8008);
and U8462 (N_8462,N_8032,N_8201);
nor U8463 (N_8463,N_8040,N_8037);
and U8464 (N_8464,N_8161,N_8216);
nand U8465 (N_8465,N_8091,N_8072);
and U8466 (N_8466,N_8117,N_8070);
nor U8467 (N_8467,N_8062,N_8026);
or U8468 (N_8468,N_8036,N_8153);
or U8469 (N_8469,N_8161,N_8126);
nor U8470 (N_8470,N_8028,N_8114);
and U8471 (N_8471,N_8141,N_8114);
and U8472 (N_8472,N_8164,N_8214);
xor U8473 (N_8473,N_8130,N_8085);
and U8474 (N_8474,N_8029,N_8101);
nor U8475 (N_8475,N_8143,N_8220);
and U8476 (N_8476,N_8220,N_8115);
and U8477 (N_8477,N_8110,N_8174);
and U8478 (N_8478,N_8204,N_8113);
nand U8479 (N_8479,N_8086,N_8232);
and U8480 (N_8480,N_8102,N_8218);
and U8481 (N_8481,N_8024,N_8140);
xnor U8482 (N_8482,N_8150,N_8013);
nor U8483 (N_8483,N_8021,N_8103);
and U8484 (N_8484,N_8177,N_8040);
nand U8485 (N_8485,N_8224,N_8082);
nor U8486 (N_8486,N_8151,N_8070);
nand U8487 (N_8487,N_8117,N_8214);
nor U8488 (N_8488,N_8215,N_8078);
xor U8489 (N_8489,N_8100,N_8019);
xor U8490 (N_8490,N_8243,N_8205);
or U8491 (N_8491,N_8076,N_8017);
or U8492 (N_8492,N_8078,N_8086);
or U8493 (N_8493,N_8099,N_8075);
and U8494 (N_8494,N_8221,N_8046);
xor U8495 (N_8495,N_8154,N_8171);
and U8496 (N_8496,N_8194,N_8089);
nor U8497 (N_8497,N_8169,N_8076);
and U8498 (N_8498,N_8137,N_8238);
xnor U8499 (N_8499,N_8117,N_8165);
nor U8500 (N_8500,N_8360,N_8385);
and U8501 (N_8501,N_8449,N_8402);
xor U8502 (N_8502,N_8321,N_8326);
xnor U8503 (N_8503,N_8362,N_8301);
xnor U8504 (N_8504,N_8394,N_8332);
nor U8505 (N_8505,N_8294,N_8405);
xnor U8506 (N_8506,N_8461,N_8298);
or U8507 (N_8507,N_8491,N_8345);
or U8508 (N_8508,N_8328,N_8463);
xor U8509 (N_8509,N_8384,N_8273);
nand U8510 (N_8510,N_8444,N_8348);
nand U8511 (N_8511,N_8254,N_8356);
nand U8512 (N_8512,N_8459,N_8325);
xor U8513 (N_8513,N_8413,N_8256);
nand U8514 (N_8514,N_8472,N_8350);
xor U8515 (N_8515,N_8478,N_8494);
nand U8516 (N_8516,N_8462,N_8331);
nand U8517 (N_8517,N_8337,N_8399);
xor U8518 (N_8518,N_8436,N_8252);
and U8519 (N_8519,N_8406,N_8264);
xnor U8520 (N_8520,N_8314,N_8260);
and U8521 (N_8521,N_8338,N_8336);
nor U8522 (N_8522,N_8471,N_8346);
nand U8523 (N_8523,N_8438,N_8349);
nor U8524 (N_8524,N_8368,N_8299);
nor U8525 (N_8525,N_8372,N_8410);
and U8526 (N_8526,N_8343,N_8416);
xor U8527 (N_8527,N_8361,N_8261);
or U8528 (N_8528,N_8378,N_8493);
xor U8529 (N_8529,N_8464,N_8443);
or U8530 (N_8530,N_8308,N_8289);
or U8531 (N_8531,N_8445,N_8412);
or U8532 (N_8532,N_8292,N_8353);
or U8533 (N_8533,N_8421,N_8380);
or U8534 (N_8534,N_8482,N_8339);
nand U8535 (N_8535,N_8423,N_8420);
nor U8536 (N_8536,N_8363,N_8408);
nand U8537 (N_8537,N_8312,N_8481);
xnor U8538 (N_8538,N_8295,N_8496);
xnor U8539 (N_8539,N_8430,N_8287);
xnor U8540 (N_8540,N_8492,N_8296);
and U8541 (N_8541,N_8476,N_8270);
xnor U8542 (N_8542,N_8383,N_8415);
or U8543 (N_8543,N_8456,N_8452);
xnor U8544 (N_8544,N_8305,N_8279);
or U8545 (N_8545,N_8390,N_8479);
nand U8546 (N_8546,N_8297,N_8475);
nand U8547 (N_8547,N_8274,N_8442);
and U8548 (N_8548,N_8495,N_8311);
nand U8549 (N_8549,N_8457,N_8377);
nand U8550 (N_8550,N_8453,N_8403);
nor U8551 (N_8551,N_8364,N_8355);
and U8552 (N_8552,N_8327,N_8469);
nand U8553 (N_8553,N_8392,N_8285);
xnor U8554 (N_8554,N_8320,N_8448);
or U8555 (N_8555,N_8439,N_8302);
or U8556 (N_8556,N_8466,N_8291);
nand U8557 (N_8557,N_8286,N_8359);
and U8558 (N_8558,N_8450,N_8486);
nand U8559 (N_8559,N_8396,N_8354);
xor U8560 (N_8560,N_8388,N_8400);
nor U8561 (N_8561,N_8446,N_8266);
xor U8562 (N_8562,N_8426,N_8447);
nor U8563 (N_8563,N_8318,N_8488);
xnor U8564 (N_8564,N_8283,N_8365);
or U8565 (N_8565,N_8409,N_8440);
nand U8566 (N_8566,N_8467,N_8379);
or U8567 (N_8567,N_8358,N_8300);
xnor U8568 (N_8568,N_8451,N_8454);
and U8569 (N_8569,N_8341,N_8330);
nor U8570 (N_8570,N_8422,N_8322);
xnor U8571 (N_8571,N_8333,N_8324);
and U8572 (N_8572,N_8376,N_8309);
nor U8573 (N_8573,N_8382,N_8428);
and U8574 (N_8574,N_8271,N_8265);
nor U8575 (N_8575,N_8329,N_8489);
nand U8576 (N_8576,N_8276,N_8281);
xor U8577 (N_8577,N_8480,N_8437);
nand U8578 (N_8578,N_8497,N_8395);
nand U8579 (N_8579,N_8347,N_8498);
and U8580 (N_8580,N_8373,N_8460);
or U8581 (N_8581,N_8398,N_8389);
nand U8582 (N_8582,N_8257,N_8351);
xnor U8583 (N_8583,N_8342,N_8458);
nor U8584 (N_8584,N_8468,N_8307);
or U8585 (N_8585,N_8272,N_8313);
nand U8586 (N_8586,N_8386,N_8404);
and U8587 (N_8587,N_8401,N_8269);
xor U8588 (N_8588,N_8310,N_8490);
nand U8589 (N_8589,N_8319,N_8431);
or U8590 (N_8590,N_8427,N_8369);
nand U8591 (N_8591,N_8419,N_8414);
or U8592 (N_8592,N_8417,N_8288);
nor U8593 (N_8593,N_8280,N_8259);
nor U8594 (N_8594,N_8268,N_8391);
and U8595 (N_8595,N_8253,N_8293);
and U8596 (N_8596,N_8334,N_8316);
nor U8597 (N_8597,N_8397,N_8323);
and U8598 (N_8598,N_8474,N_8434);
or U8599 (N_8599,N_8424,N_8425);
and U8600 (N_8600,N_8317,N_8262);
nand U8601 (N_8601,N_8277,N_8435);
nor U8602 (N_8602,N_8375,N_8411);
or U8603 (N_8603,N_8470,N_8433);
and U8604 (N_8604,N_8275,N_8315);
or U8605 (N_8605,N_8374,N_8499);
and U8606 (N_8606,N_8366,N_8473);
or U8607 (N_8607,N_8352,N_8418);
nand U8608 (N_8608,N_8306,N_8267);
or U8609 (N_8609,N_8255,N_8370);
xnor U8610 (N_8610,N_8485,N_8304);
and U8611 (N_8611,N_8441,N_8429);
nor U8612 (N_8612,N_8371,N_8357);
nand U8613 (N_8613,N_8455,N_8290);
nand U8614 (N_8614,N_8483,N_8465);
xnor U8615 (N_8615,N_8258,N_8278);
or U8616 (N_8616,N_8335,N_8387);
xor U8617 (N_8617,N_8303,N_8393);
xnor U8618 (N_8618,N_8250,N_8487);
xnor U8619 (N_8619,N_8263,N_8407);
or U8620 (N_8620,N_8251,N_8282);
and U8621 (N_8621,N_8432,N_8367);
xnor U8622 (N_8622,N_8381,N_8477);
and U8623 (N_8623,N_8484,N_8340);
and U8624 (N_8624,N_8284,N_8344);
or U8625 (N_8625,N_8306,N_8259);
nor U8626 (N_8626,N_8283,N_8466);
or U8627 (N_8627,N_8313,N_8387);
xnor U8628 (N_8628,N_8432,N_8252);
or U8629 (N_8629,N_8370,N_8346);
nor U8630 (N_8630,N_8378,N_8435);
and U8631 (N_8631,N_8407,N_8279);
nor U8632 (N_8632,N_8454,N_8289);
nand U8633 (N_8633,N_8393,N_8440);
nor U8634 (N_8634,N_8426,N_8440);
nand U8635 (N_8635,N_8377,N_8379);
xor U8636 (N_8636,N_8493,N_8363);
nand U8637 (N_8637,N_8449,N_8255);
nor U8638 (N_8638,N_8378,N_8310);
or U8639 (N_8639,N_8404,N_8349);
and U8640 (N_8640,N_8465,N_8459);
xnor U8641 (N_8641,N_8290,N_8339);
nor U8642 (N_8642,N_8462,N_8300);
and U8643 (N_8643,N_8324,N_8488);
nand U8644 (N_8644,N_8275,N_8443);
or U8645 (N_8645,N_8376,N_8477);
xnor U8646 (N_8646,N_8487,N_8357);
or U8647 (N_8647,N_8454,N_8401);
xor U8648 (N_8648,N_8276,N_8407);
nor U8649 (N_8649,N_8269,N_8256);
or U8650 (N_8650,N_8362,N_8259);
nand U8651 (N_8651,N_8367,N_8279);
and U8652 (N_8652,N_8442,N_8429);
nor U8653 (N_8653,N_8321,N_8376);
or U8654 (N_8654,N_8391,N_8387);
and U8655 (N_8655,N_8295,N_8492);
nand U8656 (N_8656,N_8293,N_8305);
nand U8657 (N_8657,N_8396,N_8475);
nor U8658 (N_8658,N_8366,N_8257);
or U8659 (N_8659,N_8459,N_8332);
nor U8660 (N_8660,N_8358,N_8307);
or U8661 (N_8661,N_8492,N_8345);
and U8662 (N_8662,N_8392,N_8456);
and U8663 (N_8663,N_8336,N_8269);
xor U8664 (N_8664,N_8442,N_8365);
or U8665 (N_8665,N_8349,N_8292);
xnor U8666 (N_8666,N_8417,N_8407);
nor U8667 (N_8667,N_8460,N_8402);
nand U8668 (N_8668,N_8345,N_8320);
nor U8669 (N_8669,N_8279,N_8276);
or U8670 (N_8670,N_8325,N_8394);
or U8671 (N_8671,N_8314,N_8369);
xnor U8672 (N_8672,N_8492,N_8437);
and U8673 (N_8673,N_8361,N_8255);
and U8674 (N_8674,N_8382,N_8316);
nor U8675 (N_8675,N_8337,N_8253);
xnor U8676 (N_8676,N_8469,N_8366);
xor U8677 (N_8677,N_8407,N_8300);
and U8678 (N_8678,N_8377,N_8272);
nand U8679 (N_8679,N_8415,N_8303);
or U8680 (N_8680,N_8448,N_8410);
or U8681 (N_8681,N_8356,N_8469);
xnor U8682 (N_8682,N_8348,N_8470);
nor U8683 (N_8683,N_8480,N_8442);
nand U8684 (N_8684,N_8356,N_8302);
xnor U8685 (N_8685,N_8323,N_8257);
nand U8686 (N_8686,N_8291,N_8290);
xor U8687 (N_8687,N_8360,N_8368);
or U8688 (N_8688,N_8308,N_8269);
nand U8689 (N_8689,N_8424,N_8303);
xnor U8690 (N_8690,N_8435,N_8434);
nand U8691 (N_8691,N_8306,N_8370);
nor U8692 (N_8692,N_8310,N_8495);
or U8693 (N_8693,N_8304,N_8298);
and U8694 (N_8694,N_8335,N_8309);
and U8695 (N_8695,N_8443,N_8408);
and U8696 (N_8696,N_8410,N_8346);
or U8697 (N_8697,N_8455,N_8413);
or U8698 (N_8698,N_8441,N_8397);
and U8699 (N_8699,N_8293,N_8480);
nor U8700 (N_8700,N_8293,N_8342);
nor U8701 (N_8701,N_8497,N_8483);
nor U8702 (N_8702,N_8260,N_8390);
xor U8703 (N_8703,N_8399,N_8288);
xor U8704 (N_8704,N_8291,N_8266);
or U8705 (N_8705,N_8333,N_8366);
nor U8706 (N_8706,N_8439,N_8404);
nand U8707 (N_8707,N_8421,N_8462);
nor U8708 (N_8708,N_8290,N_8481);
and U8709 (N_8709,N_8306,N_8356);
or U8710 (N_8710,N_8420,N_8276);
and U8711 (N_8711,N_8310,N_8439);
nor U8712 (N_8712,N_8431,N_8292);
nor U8713 (N_8713,N_8394,N_8381);
xnor U8714 (N_8714,N_8460,N_8325);
nand U8715 (N_8715,N_8415,N_8282);
xor U8716 (N_8716,N_8280,N_8427);
nor U8717 (N_8717,N_8399,N_8274);
xor U8718 (N_8718,N_8294,N_8478);
nand U8719 (N_8719,N_8438,N_8496);
or U8720 (N_8720,N_8277,N_8427);
xnor U8721 (N_8721,N_8472,N_8260);
nand U8722 (N_8722,N_8373,N_8389);
nand U8723 (N_8723,N_8298,N_8381);
nand U8724 (N_8724,N_8495,N_8397);
nand U8725 (N_8725,N_8337,N_8305);
nor U8726 (N_8726,N_8480,N_8441);
or U8727 (N_8727,N_8392,N_8376);
xnor U8728 (N_8728,N_8469,N_8442);
or U8729 (N_8729,N_8364,N_8379);
xor U8730 (N_8730,N_8297,N_8446);
or U8731 (N_8731,N_8428,N_8467);
or U8732 (N_8732,N_8424,N_8263);
xor U8733 (N_8733,N_8409,N_8333);
and U8734 (N_8734,N_8251,N_8329);
nor U8735 (N_8735,N_8468,N_8332);
or U8736 (N_8736,N_8298,N_8435);
and U8737 (N_8737,N_8470,N_8356);
nor U8738 (N_8738,N_8310,N_8484);
or U8739 (N_8739,N_8340,N_8317);
nor U8740 (N_8740,N_8258,N_8292);
or U8741 (N_8741,N_8337,N_8405);
xnor U8742 (N_8742,N_8393,N_8402);
nor U8743 (N_8743,N_8393,N_8493);
and U8744 (N_8744,N_8310,N_8321);
or U8745 (N_8745,N_8406,N_8380);
or U8746 (N_8746,N_8273,N_8318);
and U8747 (N_8747,N_8293,N_8366);
xor U8748 (N_8748,N_8344,N_8387);
or U8749 (N_8749,N_8435,N_8255);
nand U8750 (N_8750,N_8513,N_8690);
xor U8751 (N_8751,N_8747,N_8652);
xnor U8752 (N_8752,N_8705,N_8736);
xor U8753 (N_8753,N_8745,N_8589);
nor U8754 (N_8754,N_8593,N_8707);
and U8755 (N_8755,N_8710,N_8730);
xnor U8756 (N_8756,N_8700,N_8640);
or U8757 (N_8757,N_8732,N_8653);
nand U8758 (N_8758,N_8679,N_8644);
xor U8759 (N_8759,N_8697,N_8534);
or U8760 (N_8760,N_8614,N_8667);
xnor U8761 (N_8761,N_8686,N_8568);
and U8762 (N_8762,N_8727,N_8664);
or U8763 (N_8763,N_8567,N_8709);
nand U8764 (N_8764,N_8740,N_8669);
or U8765 (N_8765,N_8529,N_8523);
or U8766 (N_8766,N_8511,N_8562);
nor U8767 (N_8767,N_8655,N_8502);
and U8768 (N_8768,N_8704,N_8546);
xor U8769 (N_8769,N_8588,N_8540);
nand U8770 (N_8770,N_8711,N_8629);
nor U8771 (N_8771,N_8739,N_8583);
nand U8772 (N_8772,N_8702,N_8620);
nand U8773 (N_8773,N_8592,N_8717);
xor U8774 (N_8774,N_8603,N_8721);
and U8775 (N_8775,N_8578,N_8550);
and U8776 (N_8776,N_8555,N_8618);
and U8777 (N_8777,N_8698,N_8662);
and U8778 (N_8778,N_8744,N_8691);
xor U8779 (N_8779,N_8526,N_8577);
nand U8780 (N_8780,N_8570,N_8575);
or U8781 (N_8781,N_8569,N_8521);
and U8782 (N_8782,N_8684,N_8648);
xor U8783 (N_8783,N_8672,N_8678);
nand U8784 (N_8784,N_8579,N_8547);
or U8785 (N_8785,N_8501,N_8587);
nand U8786 (N_8786,N_8719,N_8688);
xor U8787 (N_8787,N_8656,N_8509);
and U8788 (N_8788,N_8551,N_8675);
nand U8789 (N_8789,N_8673,N_8558);
and U8790 (N_8790,N_8639,N_8731);
and U8791 (N_8791,N_8599,N_8528);
and U8792 (N_8792,N_8632,N_8602);
nor U8793 (N_8793,N_8508,N_8622);
nor U8794 (N_8794,N_8556,N_8514);
xor U8795 (N_8795,N_8597,N_8681);
and U8796 (N_8796,N_8663,N_8591);
xnor U8797 (N_8797,N_8713,N_8659);
nand U8798 (N_8798,N_8576,N_8723);
xor U8799 (N_8799,N_8604,N_8641);
nor U8800 (N_8800,N_8515,N_8613);
or U8801 (N_8801,N_8738,N_8630);
or U8802 (N_8802,N_8586,N_8584);
or U8803 (N_8803,N_8694,N_8560);
or U8804 (N_8804,N_8537,N_8522);
nor U8805 (N_8805,N_8545,N_8674);
nor U8806 (N_8806,N_8532,N_8635);
nand U8807 (N_8807,N_8541,N_8531);
nor U8808 (N_8808,N_8668,N_8600);
and U8809 (N_8809,N_8565,N_8572);
nor U8810 (N_8810,N_8611,N_8580);
xor U8811 (N_8811,N_8714,N_8696);
xnor U8812 (N_8812,N_8566,N_8615);
xnor U8813 (N_8813,N_8748,N_8728);
and U8814 (N_8814,N_8634,N_8536);
or U8815 (N_8815,N_8631,N_8559);
or U8816 (N_8816,N_8517,N_8512);
and U8817 (N_8817,N_8654,N_8637);
xnor U8818 (N_8818,N_8716,N_8595);
xor U8819 (N_8819,N_8676,N_8538);
or U8820 (N_8820,N_8544,N_8743);
nor U8821 (N_8821,N_8677,N_8670);
and U8822 (N_8822,N_8666,N_8724);
or U8823 (N_8823,N_8510,N_8612);
nor U8824 (N_8824,N_8548,N_8506);
nand U8825 (N_8825,N_8553,N_8734);
or U8826 (N_8826,N_8628,N_8720);
xor U8827 (N_8827,N_8695,N_8527);
or U8828 (N_8828,N_8657,N_8557);
nor U8829 (N_8829,N_8725,N_8516);
or U8830 (N_8830,N_8623,N_8687);
nand U8831 (N_8831,N_8683,N_8590);
and U8832 (N_8832,N_8539,N_8530);
nand U8833 (N_8833,N_8616,N_8682);
and U8834 (N_8834,N_8507,N_8564);
nand U8835 (N_8835,N_8708,N_8519);
nor U8836 (N_8836,N_8689,N_8729);
nand U8837 (N_8837,N_8524,N_8625);
xnor U8838 (N_8838,N_8504,N_8535);
and U8839 (N_8839,N_8582,N_8661);
nor U8840 (N_8840,N_8699,N_8505);
xor U8841 (N_8841,N_8571,N_8706);
or U8842 (N_8842,N_8715,N_8607);
nor U8843 (N_8843,N_8642,N_8518);
nor U8844 (N_8844,N_8601,N_8650);
and U8845 (N_8845,N_8573,N_8645);
nor U8846 (N_8846,N_8692,N_8543);
nand U8847 (N_8847,N_8722,N_8606);
nand U8848 (N_8848,N_8621,N_8742);
xor U8849 (N_8849,N_8718,N_8549);
nand U8850 (N_8850,N_8626,N_8643);
and U8851 (N_8851,N_8520,N_8680);
nand U8852 (N_8852,N_8561,N_8671);
and U8853 (N_8853,N_8685,N_8609);
xor U8854 (N_8854,N_8660,N_8610);
xor U8855 (N_8855,N_8533,N_8605);
or U8856 (N_8856,N_8633,N_8574);
nor U8857 (N_8857,N_8649,N_8735);
nor U8858 (N_8858,N_8500,N_8585);
nor U8859 (N_8859,N_8608,N_8598);
xnor U8860 (N_8860,N_8503,N_8624);
xor U8861 (N_8861,N_8703,N_8581);
or U8862 (N_8862,N_8701,N_8665);
and U8863 (N_8863,N_8647,N_8726);
or U8864 (N_8864,N_8737,N_8693);
xor U8865 (N_8865,N_8525,N_8636);
nor U8866 (N_8866,N_8746,N_8658);
and U8867 (N_8867,N_8651,N_8712);
nor U8868 (N_8868,N_8619,N_8749);
nor U8869 (N_8869,N_8596,N_8627);
nor U8870 (N_8870,N_8552,N_8594);
or U8871 (N_8871,N_8733,N_8563);
xnor U8872 (N_8872,N_8617,N_8638);
nand U8873 (N_8873,N_8542,N_8646);
nand U8874 (N_8874,N_8741,N_8554);
or U8875 (N_8875,N_8638,N_8592);
xor U8876 (N_8876,N_8683,N_8687);
xnor U8877 (N_8877,N_8581,N_8620);
or U8878 (N_8878,N_8641,N_8723);
xnor U8879 (N_8879,N_8672,N_8656);
or U8880 (N_8880,N_8688,N_8643);
xor U8881 (N_8881,N_8577,N_8597);
and U8882 (N_8882,N_8664,N_8554);
xor U8883 (N_8883,N_8531,N_8617);
nor U8884 (N_8884,N_8696,N_8576);
nor U8885 (N_8885,N_8531,N_8685);
or U8886 (N_8886,N_8586,N_8724);
or U8887 (N_8887,N_8572,N_8631);
xor U8888 (N_8888,N_8657,N_8588);
or U8889 (N_8889,N_8647,N_8696);
nand U8890 (N_8890,N_8686,N_8564);
and U8891 (N_8891,N_8736,N_8717);
or U8892 (N_8892,N_8718,N_8672);
or U8893 (N_8893,N_8629,N_8597);
nand U8894 (N_8894,N_8594,N_8705);
nor U8895 (N_8895,N_8735,N_8696);
xor U8896 (N_8896,N_8749,N_8679);
nor U8897 (N_8897,N_8546,N_8717);
or U8898 (N_8898,N_8502,N_8543);
xnor U8899 (N_8899,N_8707,N_8566);
xor U8900 (N_8900,N_8724,N_8509);
or U8901 (N_8901,N_8729,N_8512);
nand U8902 (N_8902,N_8577,N_8520);
nor U8903 (N_8903,N_8603,N_8543);
or U8904 (N_8904,N_8506,N_8553);
nor U8905 (N_8905,N_8505,N_8691);
nor U8906 (N_8906,N_8579,N_8723);
nor U8907 (N_8907,N_8706,N_8575);
xor U8908 (N_8908,N_8541,N_8529);
or U8909 (N_8909,N_8688,N_8730);
and U8910 (N_8910,N_8583,N_8514);
xor U8911 (N_8911,N_8597,N_8640);
and U8912 (N_8912,N_8703,N_8616);
or U8913 (N_8913,N_8697,N_8547);
nand U8914 (N_8914,N_8737,N_8504);
nor U8915 (N_8915,N_8545,N_8608);
or U8916 (N_8916,N_8629,N_8634);
nor U8917 (N_8917,N_8638,N_8606);
or U8918 (N_8918,N_8697,N_8500);
nand U8919 (N_8919,N_8524,N_8554);
or U8920 (N_8920,N_8660,N_8661);
nand U8921 (N_8921,N_8547,N_8575);
xnor U8922 (N_8922,N_8626,N_8637);
and U8923 (N_8923,N_8648,N_8608);
nor U8924 (N_8924,N_8735,N_8684);
xor U8925 (N_8925,N_8714,N_8740);
xnor U8926 (N_8926,N_8747,N_8717);
nor U8927 (N_8927,N_8647,N_8515);
xnor U8928 (N_8928,N_8648,N_8626);
xnor U8929 (N_8929,N_8607,N_8672);
nand U8930 (N_8930,N_8605,N_8738);
or U8931 (N_8931,N_8687,N_8560);
nor U8932 (N_8932,N_8662,N_8588);
or U8933 (N_8933,N_8720,N_8581);
nor U8934 (N_8934,N_8723,N_8730);
and U8935 (N_8935,N_8698,N_8609);
nor U8936 (N_8936,N_8513,N_8523);
and U8937 (N_8937,N_8644,N_8607);
nor U8938 (N_8938,N_8658,N_8630);
nand U8939 (N_8939,N_8661,N_8668);
xor U8940 (N_8940,N_8689,N_8570);
or U8941 (N_8941,N_8744,N_8683);
nand U8942 (N_8942,N_8705,N_8517);
and U8943 (N_8943,N_8613,N_8697);
nor U8944 (N_8944,N_8556,N_8518);
or U8945 (N_8945,N_8616,N_8731);
nand U8946 (N_8946,N_8639,N_8699);
nor U8947 (N_8947,N_8740,N_8666);
nand U8948 (N_8948,N_8684,N_8617);
or U8949 (N_8949,N_8695,N_8621);
or U8950 (N_8950,N_8599,N_8552);
nand U8951 (N_8951,N_8595,N_8685);
and U8952 (N_8952,N_8560,N_8518);
nand U8953 (N_8953,N_8658,N_8745);
nor U8954 (N_8954,N_8582,N_8747);
nor U8955 (N_8955,N_8601,N_8684);
nand U8956 (N_8956,N_8725,N_8662);
nand U8957 (N_8957,N_8688,N_8531);
nor U8958 (N_8958,N_8601,N_8624);
nor U8959 (N_8959,N_8601,N_8527);
and U8960 (N_8960,N_8508,N_8724);
and U8961 (N_8961,N_8703,N_8643);
xnor U8962 (N_8962,N_8638,N_8698);
nor U8963 (N_8963,N_8676,N_8520);
nor U8964 (N_8964,N_8635,N_8529);
or U8965 (N_8965,N_8607,N_8562);
nor U8966 (N_8966,N_8526,N_8504);
and U8967 (N_8967,N_8620,N_8624);
xnor U8968 (N_8968,N_8628,N_8588);
nor U8969 (N_8969,N_8703,N_8558);
or U8970 (N_8970,N_8702,N_8670);
nor U8971 (N_8971,N_8595,N_8648);
xor U8972 (N_8972,N_8661,N_8596);
nor U8973 (N_8973,N_8565,N_8735);
or U8974 (N_8974,N_8746,N_8617);
or U8975 (N_8975,N_8702,N_8585);
or U8976 (N_8976,N_8740,N_8578);
nor U8977 (N_8977,N_8613,N_8647);
or U8978 (N_8978,N_8706,N_8638);
xor U8979 (N_8979,N_8545,N_8502);
xor U8980 (N_8980,N_8719,N_8610);
nor U8981 (N_8981,N_8646,N_8706);
or U8982 (N_8982,N_8706,N_8727);
nand U8983 (N_8983,N_8589,N_8708);
nor U8984 (N_8984,N_8545,N_8676);
xor U8985 (N_8985,N_8504,N_8638);
or U8986 (N_8986,N_8593,N_8601);
xor U8987 (N_8987,N_8744,N_8507);
nand U8988 (N_8988,N_8748,N_8623);
nand U8989 (N_8989,N_8713,N_8641);
and U8990 (N_8990,N_8682,N_8518);
and U8991 (N_8991,N_8647,N_8510);
or U8992 (N_8992,N_8638,N_8508);
nand U8993 (N_8993,N_8566,N_8726);
xnor U8994 (N_8994,N_8588,N_8716);
xor U8995 (N_8995,N_8584,N_8747);
or U8996 (N_8996,N_8646,N_8654);
nor U8997 (N_8997,N_8670,N_8664);
and U8998 (N_8998,N_8513,N_8706);
nand U8999 (N_8999,N_8663,N_8644);
or U9000 (N_9000,N_8847,N_8802);
nand U9001 (N_9001,N_8954,N_8834);
and U9002 (N_9002,N_8965,N_8853);
or U9003 (N_9003,N_8875,N_8793);
nor U9004 (N_9004,N_8771,N_8915);
xnor U9005 (N_9005,N_8973,N_8968);
nor U9006 (N_9006,N_8930,N_8785);
nor U9007 (N_9007,N_8983,N_8960);
nand U9008 (N_9008,N_8891,N_8987);
nand U9009 (N_9009,N_8843,N_8974);
and U9010 (N_9010,N_8905,N_8901);
nor U9011 (N_9011,N_8964,N_8938);
and U9012 (N_9012,N_8775,N_8856);
and U9013 (N_9013,N_8889,N_8912);
and U9014 (N_9014,N_8830,N_8997);
and U9015 (N_9015,N_8962,N_8819);
nand U9016 (N_9016,N_8970,N_8870);
nor U9017 (N_9017,N_8943,N_8831);
nand U9018 (N_9018,N_8898,N_8772);
and U9019 (N_9019,N_8893,N_8907);
xnor U9020 (N_9020,N_8984,N_8874);
nand U9021 (N_9021,N_8778,N_8883);
nor U9022 (N_9022,N_8777,N_8823);
and U9023 (N_9023,N_8877,N_8995);
nor U9024 (N_9024,N_8825,N_8882);
and U9025 (N_9025,N_8763,N_8795);
or U9026 (N_9026,N_8986,N_8949);
nor U9027 (N_9027,N_8985,N_8854);
and U9028 (N_9028,N_8947,N_8791);
and U9029 (N_9029,N_8939,N_8850);
nor U9030 (N_9030,N_8897,N_8837);
or U9031 (N_9031,N_8796,N_8921);
and U9032 (N_9032,N_8942,N_8910);
nand U9033 (N_9033,N_8774,N_8993);
nand U9034 (N_9034,N_8754,N_8919);
nor U9035 (N_9035,N_8767,N_8818);
nand U9036 (N_9036,N_8923,N_8955);
or U9037 (N_9037,N_8876,N_8781);
and U9038 (N_9038,N_8779,N_8925);
nor U9039 (N_9039,N_8751,N_8809);
or U9040 (N_9040,N_8769,N_8892);
or U9041 (N_9041,N_8959,N_8896);
xnor U9042 (N_9042,N_8935,N_8895);
and U9043 (N_9043,N_8977,N_8851);
xor U9044 (N_9044,N_8773,N_8886);
or U9045 (N_9045,N_8758,N_8998);
or U9046 (N_9046,N_8827,N_8918);
or U9047 (N_9047,N_8826,N_8953);
xor U9048 (N_9048,N_8860,N_8928);
nand U9049 (N_9049,N_8884,N_8755);
or U9050 (N_9050,N_8979,N_8858);
and U9051 (N_9051,N_8946,N_8931);
and U9052 (N_9052,N_8994,N_8840);
nor U9053 (N_9053,N_8967,N_8963);
or U9054 (N_9054,N_8804,N_8828);
xor U9055 (N_9055,N_8845,N_8881);
xor U9056 (N_9056,N_8760,N_8934);
nor U9057 (N_9057,N_8917,N_8792);
or U9058 (N_9058,N_8878,N_8806);
nor U9059 (N_9059,N_8813,N_8757);
nand U9060 (N_9060,N_8936,N_8866);
and U9061 (N_9061,N_8846,N_8820);
or U9062 (N_9062,N_8812,N_8871);
nor U9063 (N_9063,N_8805,N_8975);
and U9064 (N_9064,N_8879,N_8855);
or U9065 (N_9065,N_8768,N_8982);
xor U9066 (N_9066,N_8865,N_8815);
and U9067 (N_9067,N_8864,N_8981);
and U9068 (N_9068,N_8969,N_8770);
nor U9069 (N_9069,N_8794,N_8797);
nor U9070 (N_9070,N_8839,N_8788);
nand U9071 (N_9071,N_8937,N_8750);
or U9072 (N_9072,N_8824,N_8990);
nor U9073 (N_9073,N_8902,N_8782);
nor U9074 (N_9074,N_8872,N_8933);
nand U9075 (N_9075,N_8958,N_8838);
nor U9076 (N_9076,N_8842,N_8894);
nand U9077 (N_9077,N_8800,N_8857);
xor U9078 (N_9078,N_8822,N_8926);
or U9079 (N_9079,N_8863,N_8980);
and U9080 (N_9080,N_8861,N_8811);
nor U9081 (N_9081,N_8786,N_8888);
nor U9082 (N_9082,N_8887,N_8948);
or U9083 (N_9083,N_8833,N_8885);
and U9084 (N_9084,N_8932,N_8852);
or U9085 (N_9085,N_8988,N_8961);
xnor U9086 (N_9086,N_8869,N_8835);
xnor U9087 (N_9087,N_8801,N_8868);
xor U9088 (N_9088,N_8780,N_8904);
nor U9089 (N_9089,N_8950,N_8927);
or U9090 (N_9090,N_8762,N_8849);
and U9091 (N_9091,N_8944,N_8752);
and U9092 (N_9092,N_8844,N_8765);
and U9093 (N_9093,N_8829,N_8821);
xor U9094 (N_9094,N_8787,N_8924);
or U9095 (N_9095,N_8940,N_8817);
and U9096 (N_9096,N_8756,N_8810);
or U9097 (N_9097,N_8900,N_8914);
nand U9098 (N_9098,N_8976,N_8761);
and U9099 (N_9099,N_8764,N_8799);
nand U9100 (N_9100,N_8798,N_8841);
and U9101 (N_9101,N_8899,N_8978);
and U9102 (N_9102,N_8903,N_8913);
or U9103 (N_9103,N_8957,N_8929);
xor U9104 (N_9104,N_8951,N_8808);
and U9105 (N_9105,N_8991,N_8920);
nand U9106 (N_9106,N_8908,N_8790);
or U9107 (N_9107,N_8945,N_8783);
nor U9108 (N_9108,N_8996,N_8922);
nor U9109 (N_9109,N_8789,N_8972);
nor U9110 (N_9110,N_8911,N_8916);
or U9111 (N_9111,N_8862,N_8941);
xnor U9112 (N_9112,N_8999,N_8816);
or U9113 (N_9113,N_8759,N_8952);
and U9114 (N_9114,N_8956,N_8992);
xor U9115 (N_9115,N_8890,N_8966);
nand U9116 (N_9116,N_8803,N_8859);
xnor U9117 (N_9117,N_8873,N_8807);
xor U9118 (N_9118,N_8906,N_8814);
nand U9119 (N_9119,N_8880,N_8909);
and U9120 (N_9120,N_8867,N_8784);
nand U9121 (N_9121,N_8776,N_8989);
xnor U9122 (N_9122,N_8848,N_8766);
and U9123 (N_9123,N_8832,N_8971);
and U9124 (N_9124,N_8836,N_8753);
and U9125 (N_9125,N_8806,N_8901);
xor U9126 (N_9126,N_8787,N_8897);
nand U9127 (N_9127,N_8959,N_8979);
and U9128 (N_9128,N_8758,N_8978);
nor U9129 (N_9129,N_8786,N_8764);
or U9130 (N_9130,N_8819,N_8873);
nor U9131 (N_9131,N_8971,N_8755);
and U9132 (N_9132,N_8808,N_8969);
and U9133 (N_9133,N_8973,N_8945);
or U9134 (N_9134,N_8755,N_8973);
or U9135 (N_9135,N_8878,N_8750);
and U9136 (N_9136,N_8978,N_8822);
nor U9137 (N_9137,N_8867,N_8760);
xnor U9138 (N_9138,N_8761,N_8857);
xor U9139 (N_9139,N_8916,N_8807);
nand U9140 (N_9140,N_8853,N_8905);
nor U9141 (N_9141,N_8874,N_8755);
and U9142 (N_9142,N_8824,N_8953);
and U9143 (N_9143,N_8995,N_8813);
nand U9144 (N_9144,N_8775,N_8787);
and U9145 (N_9145,N_8785,N_8766);
xor U9146 (N_9146,N_8935,N_8894);
nand U9147 (N_9147,N_8864,N_8855);
nand U9148 (N_9148,N_8981,N_8831);
and U9149 (N_9149,N_8765,N_8909);
xnor U9150 (N_9150,N_8756,N_8778);
or U9151 (N_9151,N_8924,N_8930);
nand U9152 (N_9152,N_8910,N_8999);
nand U9153 (N_9153,N_8937,N_8864);
or U9154 (N_9154,N_8924,N_8935);
xor U9155 (N_9155,N_8977,N_8996);
or U9156 (N_9156,N_8853,N_8921);
and U9157 (N_9157,N_8792,N_8979);
nor U9158 (N_9158,N_8973,N_8799);
and U9159 (N_9159,N_8868,N_8782);
xor U9160 (N_9160,N_8810,N_8782);
or U9161 (N_9161,N_8955,N_8933);
xor U9162 (N_9162,N_8975,N_8983);
or U9163 (N_9163,N_8864,N_8963);
or U9164 (N_9164,N_8979,N_8908);
nor U9165 (N_9165,N_8891,N_8992);
nand U9166 (N_9166,N_8834,N_8927);
or U9167 (N_9167,N_8790,N_8894);
nor U9168 (N_9168,N_8753,N_8835);
nor U9169 (N_9169,N_8832,N_8788);
or U9170 (N_9170,N_8826,N_8878);
and U9171 (N_9171,N_8877,N_8778);
xnor U9172 (N_9172,N_8927,N_8929);
or U9173 (N_9173,N_8823,N_8963);
xnor U9174 (N_9174,N_8903,N_8926);
or U9175 (N_9175,N_8860,N_8932);
or U9176 (N_9176,N_8768,N_8844);
nand U9177 (N_9177,N_8797,N_8783);
or U9178 (N_9178,N_8976,N_8878);
xor U9179 (N_9179,N_8874,N_8930);
nand U9180 (N_9180,N_8962,N_8973);
and U9181 (N_9181,N_8808,N_8829);
nor U9182 (N_9182,N_8811,N_8762);
xnor U9183 (N_9183,N_8880,N_8977);
or U9184 (N_9184,N_8937,N_8885);
nand U9185 (N_9185,N_8882,N_8897);
nor U9186 (N_9186,N_8823,N_8788);
or U9187 (N_9187,N_8939,N_8979);
and U9188 (N_9188,N_8839,N_8980);
xor U9189 (N_9189,N_8828,N_8914);
nand U9190 (N_9190,N_8791,N_8800);
and U9191 (N_9191,N_8997,N_8752);
and U9192 (N_9192,N_8799,N_8993);
nor U9193 (N_9193,N_8931,N_8815);
nand U9194 (N_9194,N_8901,N_8888);
or U9195 (N_9195,N_8756,N_8889);
nand U9196 (N_9196,N_8858,N_8943);
nand U9197 (N_9197,N_8894,N_8819);
or U9198 (N_9198,N_8912,N_8820);
xor U9199 (N_9199,N_8895,N_8944);
nand U9200 (N_9200,N_8768,N_8801);
and U9201 (N_9201,N_8964,N_8791);
nor U9202 (N_9202,N_8897,N_8871);
nand U9203 (N_9203,N_8773,N_8813);
xor U9204 (N_9204,N_8919,N_8767);
nor U9205 (N_9205,N_8753,N_8814);
nand U9206 (N_9206,N_8803,N_8996);
or U9207 (N_9207,N_8900,N_8858);
and U9208 (N_9208,N_8877,N_8774);
xor U9209 (N_9209,N_8965,N_8913);
xor U9210 (N_9210,N_8765,N_8774);
nor U9211 (N_9211,N_8772,N_8982);
or U9212 (N_9212,N_8833,N_8878);
and U9213 (N_9213,N_8757,N_8782);
nor U9214 (N_9214,N_8939,N_8883);
or U9215 (N_9215,N_8885,N_8774);
nand U9216 (N_9216,N_8828,N_8968);
xor U9217 (N_9217,N_8911,N_8981);
or U9218 (N_9218,N_8861,N_8900);
and U9219 (N_9219,N_8794,N_8839);
nand U9220 (N_9220,N_8842,N_8935);
nand U9221 (N_9221,N_8864,N_8858);
nand U9222 (N_9222,N_8763,N_8773);
xor U9223 (N_9223,N_8983,N_8864);
or U9224 (N_9224,N_8839,N_8989);
or U9225 (N_9225,N_8834,N_8889);
xnor U9226 (N_9226,N_8998,N_8971);
nand U9227 (N_9227,N_8881,N_8888);
or U9228 (N_9228,N_8922,N_8890);
and U9229 (N_9229,N_8980,N_8995);
nor U9230 (N_9230,N_8810,N_8830);
or U9231 (N_9231,N_8903,N_8810);
xnor U9232 (N_9232,N_8811,N_8947);
or U9233 (N_9233,N_8899,N_8785);
nand U9234 (N_9234,N_8797,N_8780);
nand U9235 (N_9235,N_8836,N_8977);
nor U9236 (N_9236,N_8838,N_8928);
and U9237 (N_9237,N_8776,N_8782);
or U9238 (N_9238,N_8980,N_8785);
or U9239 (N_9239,N_8835,N_8867);
or U9240 (N_9240,N_8919,N_8903);
and U9241 (N_9241,N_8820,N_8825);
nor U9242 (N_9242,N_8808,N_8897);
or U9243 (N_9243,N_8874,N_8851);
or U9244 (N_9244,N_8854,N_8831);
nand U9245 (N_9245,N_8859,N_8829);
or U9246 (N_9246,N_8752,N_8921);
or U9247 (N_9247,N_8986,N_8811);
xnor U9248 (N_9248,N_8779,N_8817);
or U9249 (N_9249,N_8823,N_8822);
or U9250 (N_9250,N_9170,N_9196);
xnor U9251 (N_9251,N_9031,N_9222);
xnor U9252 (N_9252,N_9158,N_9015);
nand U9253 (N_9253,N_9018,N_9039);
and U9254 (N_9254,N_9085,N_9001);
or U9255 (N_9255,N_9019,N_9144);
nand U9256 (N_9256,N_9043,N_9160);
nor U9257 (N_9257,N_9166,N_9204);
nor U9258 (N_9258,N_9137,N_9040);
and U9259 (N_9259,N_9184,N_9125);
or U9260 (N_9260,N_9134,N_9096);
or U9261 (N_9261,N_9094,N_9182);
nand U9262 (N_9262,N_9050,N_9017);
or U9263 (N_9263,N_9044,N_9091);
and U9264 (N_9264,N_9092,N_9037);
and U9265 (N_9265,N_9119,N_9097);
nor U9266 (N_9266,N_9235,N_9230);
nor U9267 (N_9267,N_9150,N_9034);
or U9268 (N_9268,N_9200,N_9122);
nand U9269 (N_9269,N_9082,N_9047);
and U9270 (N_9270,N_9058,N_9205);
or U9271 (N_9271,N_9198,N_9120);
and U9272 (N_9272,N_9143,N_9231);
or U9273 (N_9273,N_9070,N_9048);
nand U9274 (N_9274,N_9192,N_9236);
nand U9275 (N_9275,N_9074,N_9221);
xor U9276 (N_9276,N_9126,N_9080);
or U9277 (N_9277,N_9101,N_9249);
xor U9278 (N_9278,N_9114,N_9121);
nor U9279 (N_9279,N_9178,N_9171);
nand U9280 (N_9280,N_9027,N_9087);
xor U9281 (N_9281,N_9008,N_9075);
xor U9282 (N_9282,N_9029,N_9242);
nor U9283 (N_9283,N_9138,N_9244);
nand U9284 (N_9284,N_9148,N_9006);
or U9285 (N_9285,N_9105,N_9156);
or U9286 (N_9286,N_9099,N_9209);
xor U9287 (N_9287,N_9115,N_9110);
or U9288 (N_9288,N_9055,N_9163);
and U9289 (N_9289,N_9045,N_9218);
and U9290 (N_9290,N_9116,N_9090);
xnor U9291 (N_9291,N_9141,N_9046);
or U9292 (N_9292,N_9217,N_9003);
nor U9293 (N_9293,N_9234,N_9162);
or U9294 (N_9294,N_9147,N_9062);
xor U9295 (N_9295,N_9100,N_9157);
or U9296 (N_9296,N_9164,N_9129);
nand U9297 (N_9297,N_9131,N_9084);
and U9298 (N_9298,N_9028,N_9191);
or U9299 (N_9299,N_9103,N_9064);
or U9300 (N_9300,N_9183,N_9011);
nor U9301 (N_9301,N_9022,N_9118);
nand U9302 (N_9302,N_9241,N_9245);
nand U9303 (N_9303,N_9127,N_9023);
nand U9304 (N_9304,N_9168,N_9053);
or U9305 (N_9305,N_9177,N_9024);
or U9306 (N_9306,N_9026,N_9123);
or U9307 (N_9307,N_9223,N_9102);
nor U9308 (N_9308,N_9214,N_9220);
or U9309 (N_9309,N_9237,N_9173);
or U9310 (N_9310,N_9061,N_9007);
nand U9311 (N_9311,N_9154,N_9069);
xor U9312 (N_9312,N_9239,N_9169);
or U9313 (N_9313,N_9195,N_9113);
or U9314 (N_9314,N_9212,N_9213);
nand U9315 (N_9315,N_9051,N_9077);
nor U9316 (N_9316,N_9189,N_9229);
nor U9317 (N_9317,N_9215,N_9057);
nand U9318 (N_9318,N_9207,N_9188);
and U9319 (N_9319,N_9179,N_9104);
xor U9320 (N_9320,N_9032,N_9202);
or U9321 (N_9321,N_9232,N_9086);
nand U9322 (N_9322,N_9038,N_9009);
and U9323 (N_9323,N_9130,N_9112);
xnor U9324 (N_9324,N_9238,N_9224);
and U9325 (N_9325,N_9056,N_9049);
xnor U9326 (N_9326,N_9228,N_9194);
xnor U9327 (N_9327,N_9054,N_9206);
or U9328 (N_9328,N_9247,N_9145);
xor U9329 (N_9329,N_9211,N_9066);
and U9330 (N_9330,N_9016,N_9203);
or U9331 (N_9331,N_9185,N_9072);
xor U9332 (N_9332,N_9216,N_9065);
xor U9333 (N_9333,N_9167,N_9181);
or U9334 (N_9334,N_9165,N_9079);
nor U9335 (N_9335,N_9042,N_9176);
nand U9336 (N_9336,N_9071,N_9190);
and U9337 (N_9337,N_9159,N_9010);
or U9338 (N_9338,N_9005,N_9109);
xor U9339 (N_9339,N_9219,N_9227);
nor U9340 (N_9340,N_9243,N_9152);
and U9341 (N_9341,N_9076,N_9108);
nand U9342 (N_9342,N_9012,N_9174);
nor U9343 (N_9343,N_9248,N_9067);
and U9344 (N_9344,N_9240,N_9161);
or U9345 (N_9345,N_9201,N_9002);
nand U9346 (N_9346,N_9095,N_9059);
and U9347 (N_9347,N_9175,N_9199);
xnor U9348 (N_9348,N_9153,N_9060);
nand U9349 (N_9349,N_9149,N_9081);
nand U9350 (N_9350,N_9025,N_9117);
and U9351 (N_9351,N_9226,N_9004);
nor U9352 (N_9352,N_9132,N_9106);
xor U9353 (N_9353,N_9030,N_9172);
and U9354 (N_9354,N_9068,N_9187);
and U9355 (N_9355,N_9225,N_9020);
nor U9356 (N_9356,N_9246,N_9111);
nand U9357 (N_9357,N_9136,N_9107);
nand U9358 (N_9358,N_9036,N_9193);
nor U9359 (N_9359,N_9208,N_9089);
or U9360 (N_9360,N_9197,N_9098);
nand U9361 (N_9361,N_9133,N_9033);
or U9362 (N_9362,N_9041,N_9063);
or U9363 (N_9363,N_9088,N_9233);
nand U9364 (N_9364,N_9035,N_9140);
xor U9365 (N_9365,N_9155,N_9210);
nor U9366 (N_9366,N_9021,N_9073);
nand U9367 (N_9367,N_9083,N_9124);
nor U9368 (N_9368,N_9146,N_9093);
and U9369 (N_9369,N_9052,N_9151);
xor U9370 (N_9370,N_9186,N_9014);
xor U9371 (N_9371,N_9139,N_9142);
or U9372 (N_9372,N_9013,N_9078);
xor U9373 (N_9373,N_9180,N_9128);
nor U9374 (N_9374,N_9000,N_9135);
or U9375 (N_9375,N_9084,N_9170);
and U9376 (N_9376,N_9069,N_9164);
and U9377 (N_9377,N_9242,N_9236);
xnor U9378 (N_9378,N_9077,N_9049);
or U9379 (N_9379,N_9065,N_9037);
nor U9380 (N_9380,N_9102,N_9110);
nand U9381 (N_9381,N_9168,N_9209);
xnor U9382 (N_9382,N_9162,N_9136);
or U9383 (N_9383,N_9232,N_9016);
nor U9384 (N_9384,N_9235,N_9075);
xnor U9385 (N_9385,N_9018,N_9074);
and U9386 (N_9386,N_9209,N_9016);
nor U9387 (N_9387,N_9009,N_9163);
nand U9388 (N_9388,N_9176,N_9185);
and U9389 (N_9389,N_9191,N_9235);
or U9390 (N_9390,N_9050,N_9002);
nand U9391 (N_9391,N_9009,N_9172);
and U9392 (N_9392,N_9024,N_9028);
or U9393 (N_9393,N_9066,N_9111);
nor U9394 (N_9394,N_9011,N_9058);
or U9395 (N_9395,N_9078,N_9217);
and U9396 (N_9396,N_9236,N_9025);
and U9397 (N_9397,N_9242,N_9207);
nand U9398 (N_9398,N_9145,N_9109);
nand U9399 (N_9399,N_9027,N_9193);
or U9400 (N_9400,N_9003,N_9063);
or U9401 (N_9401,N_9185,N_9218);
nor U9402 (N_9402,N_9233,N_9061);
xor U9403 (N_9403,N_9111,N_9171);
or U9404 (N_9404,N_9124,N_9135);
nor U9405 (N_9405,N_9004,N_9224);
xor U9406 (N_9406,N_9199,N_9159);
xor U9407 (N_9407,N_9085,N_9159);
or U9408 (N_9408,N_9092,N_9229);
nand U9409 (N_9409,N_9113,N_9031);
nor U9410 (N_9410,N_9053,N_9214);
nor U9411 (N_9411,N_9182,N_9095);
nor U9412 (N_9412,N_9204,N_9188);
nand U9413 (N_9413,N_9021,N_9207);
nand U9414 (N_9414,N_9033,N_9170);
or U9415 (N_9415,N_9162,N_9202);
xor U9416 (N_9416,N_9212,N_9064);
and U9417 (N_9417,N_9166,N_9163);
nor U9418 (N_9418,N_9031,N_9139);
xnor U9419 (N_9419,N_9158,N_9020);
or U9420 (N_9420,N_9116,N_9086);
nand U9421 (N_9421,N_9075,N_9126);
nand U9422 (N_9422,N_9180,N_9117);
or U9423 (N_9423,N_9026,N_9025);
and U9424 (N_9424,N_9232,N_9052);
nand U9425 (N_9425,N_9123,N_9223);
and U9426 (N_9426,N_9059,N_9214);
and U9427 (N_9427,N_9122,N_9248);
nand U9428 (N_9428,N_9026,N_9115);
and U9429 (N_9429,N_9092,N_9038);
and U9430 (N_9430,N_9113,N_9027);
nand U9431 (N_9431,N_9189,N_9116);
xor U9432 (N_9432,N_9199,N_9036);
and U9433 (N_9433,N_9214,N_9175);
nor U9434 (N_9434,N_9184,N_9154);
xnor U9435 (N_9435,N_9215,N_9123);
and U9436 (N_9436,N_9124,N_9085);
nor U9437 (N_9437,N_9139,N_9120);
or U9438 (N_9438,N_9112,N_9183);
nor U9439 (N_9439,N_9017,N_9171);
nor U9440 (N_9440,N_9117,N_9054);
xor U9441 (N_9441,N_9228,N_9068);
xnor U9442 (N_9442,N_9156,N_9044);
xor U9443 (N_9443,N_9246,N_9107);
and U9444 (N_9444,N_9141,N_9200);
and U9445 (N_9445,N_9012,N_9184);
and U9446 (N_9446,N_9129,N_9029);
nand U9447 (N_9447,N_9177,N_9176);
nand U9448 (N_9448,N_9244,N_9046);
nand U9449 (N_9449,N_9030,N_9113);
or U9450 (N_9450,N_9147,N_9171);
or U9451 (N_9451,N_9181,N_9093);
nand U9452 (N_9452,N_9211,N_9229);
xnor U9453 (N_9453,N_9231,N_9211);
and U9454 (N_9454,N_9246,N_9233);
and U9455 (N_9455,N_9143,N_9243);
nand U9456 (N_9456,N_9092,N_9128);
or U9457 (N_9457,N_9159,N_9140);
nor U9458 (N_9458,N_9005,N_9170);
xor U9459 (N_9459,N_9055,N_9048);
nand U9460 (N_9460,N_9157,N_9237);
or U9461 (N_9461,N_9058,N_9121);
nand U9462 (N_9462,N_9046,N_9067);
and U9463 (N_9463,N_9065,N_9218);
nor U9464 (N_9464,N_9185,N_9206);
nand U9465 (N_9465,N_9233,N_9142);
nand U9466 (N_9466,N_9070,N_9024);
or U9467 (N_9467,N_9203,N_9119);
nand U9468 (N_9468,N_9090,N_9160);
xor U9469 (N_9469,N_9119,N_9102);
or U9470 (N_9470,N_9209,N_9132);
xnor U9471 (N_9471,N_9139,N_9215);
and U9472 (N_9472,N_9068,N_9061);
and U9473 (N_9473,N_9062,N_9069);
nand U9474 (N_9474,N_9195,N_9090);
nand U9475 (N_9475,N_9226,N_9214);
xor U9476 (N_9476,N_9069,N_9099);
and U9477 (N_9477,N_9184,N_9131);
nor U9478 (N_9478,N_9121,N_9247);
nor U9479 (N_9479,N_9146,N_9111);
nor U9480 (N_9480,N_9220,N_9014);
nor U9481 (N_9481,N_9176,N_9207);
nor U9482 (N_9482,N_9182,N_9121);
and U9483 (N_9483,N_9068,N_9159);
or U9484 (N_9484,N_9189,N_9222);
nor U9485 (N_9485,N_9044,N_9025);
nand U9486 (N_9486,N_9036,N_9234);
xnor U9487 (N_9487,N_9152,N_9001);
nand U9488 (N_9488,N_9174,N_9178);
nor U9489 (N_9489,N_9078,N_9091);
or U9490 (N_9490,N_9075,N_9205);
xor U9491 (N_9491,N_9007,N_9198);
nand U9492 (N_9492,N_9195,N_9057);
and U9493 (N_9493,N_9148,N_9052);
or U9494 (N_9494,N_9037,N_9157);
and U9495 (N_9495,N_9075,N_9111);
nor U9496 (N_9496,N_9129,N_9175);
and U9497 (N_9497,N_9084,N_9087);
nor U9498 (N_9498,N_9171,N_9133);
or U9499 (N_9499,N_9039,N_9031);
xnor U9500 (N_9500,N_9345,N_9270);
and U9501 (N_9501,N_9303,N_9454);
and U9502 (N_9502,N_9399,N_9479);
nand U9503 (N_9503,N_9483,N_9265);
nor U9504 (N_9504,N_9255,N_9261);
nor U9505 (N_9505,N_9367,N_9374);
or U9506 (N_9506,N_9298,N_9259);
xor U9507 (N_9507,N_9474,N_9254);
and U9508 (N_9508,N_9480,N_9438);
xnor U9509 (N_9509,N_9494,N_9421);
nor U9510 (N_9510,N_9384,N_9497);
nor U9511 (N_9511,N_9320,N_9415);
nand U9512 (N_9512,N_9444,N_9408);
or U9513 (N_9513,N_9347,N_9266);
nand U9514 (N_9514,N_9364,N_9301);
nand U9515 (N_9515,N_9429,N_9436);
nor U9516 (N_9516,N_9348,N_9441);
xor U9517 (N_9517,N_9491,N_9323);
xor U9518 (N_9518,N_9263,N_9462);
nor U9519 (N_9519,N_9431,N_9471);
or U9520 (N_9520,N_9440,N_9368);
or U9521 (N_9521,N_9433,N_9309);
xnor U9522 (N_9522,N_9279,N_9393);
nand U9523 (N_9523,N_9434,N_9290);
nand U9524 (N_9524,N_9286,N_9412);
and U9525 (N_9525,N_9416,N_9472);
nor U9526 (N_9526,N_9363,N_9486);
or U9527 (N_9527,N_9450,N_9285);
and U9528 (N_9528,N_9407,N_9280);
nand U9529 (N_9529,N_9372,N_9319);
nand U9530 (N_9530,N_9366,N_9253);
and U9531 (N_9531,N_9338,N_9273);
xor U9532 (N_9532,N_9465,N_9397);
and U9533 (N_9533,N_9312,N_9452);
xnor U9534 (N_9534,N_9250,N_9358);
and U9535 (N_9535,N_9275,N_9466);
xnor U9536 (N_9536,N_9470,N_9410);
and U9537 (N_9537,N_9477,N_9317);
xnor U9538 (N_9538,N_9356,N_9475);
nor U9539 (N_9539,N_9389,N_9446);
xor U9540 (N_9540,N_9262,N_9404);
nor U9541 (N_9541,N_9335,N_9354);
xor U9542 (N_9542,N_9401,N_9463);
nor U9543 (N_9543,N_9272,N_9449);
and U9544 (N_9544,N_9409,N_9380);
or U9545 (N_9545,N_9336,N_9304);
or U9546 (N_9546,N_9274,N_9297);
xor U9547 (N_9547,N_9496,N_9385);
and U9548 (N_9548,N_9375,N_9379);
xor U9549 (N_9549,N_9315,N_9333);
or U9550 (N_9550,N_9451,N_9457);
and U9551 (N_9551,N_9425,N_9476);
nand U9552 (N_9552,N_9313,N_9321);
nor U9553 (N_9553,N_9469,N_9365);
xnor U9554 (N_9554,N_9428,N_9377);
and U9555 (N_9555,N_9382,N_9324);
xor U9556 (N_9556,N_9299,N_9437);
or U9557 (N_9557,N_9349,N_9422);
nand U9558 (N_9558,N_9392,N_9305);
nand U9559 (N_9559,N_9258,N_9406);
xnor U9560 (N_9560,N_9281,N_9455);
xnor U9561 (N_9561,N_9340,N_9291);
xnor U9562 (N_9562,N_9473,N_9398);
or U9563 (N_9563,N_9344,N_9443);
nor U9564 (N_9564,N_9493,N_9460);
or U9565 (N_9565,N_9268,N_9316);
or U9566 (N_9566,N_9322,N_9489);
nor U9567 (N_9567,N_9332,N_9307);
nand U9568 (N_9568,N_9485,N_9487);
nand U9569 (N_9569,N_9418,N_9314);
nand U9570 (N_9570,N_9464,N_9405);
and U9571 (N_9571,N_9411,N_9490);
nand U9572 (N_9572,N_9271,N_9417);
nor U9573 (N_9573,N_9400,N_9388);
nor U9574 (N_9574,N_9495,N_9282);
nor U9575 (N_9575,N_9251,N_9287);
nor U9576 (N_9576,N_9445,N_9370);
and U9577 (N_9577,N_9387,N_9269);
xor U9578 (N_9578,N_9278,N_9378);
or U9579 (N_9579,N_9360,N_9391);
nand U9580 (N_9580,N_9403,N_9423);
nor U9581 (N_9581,N_9390,N_9355);
nand U9582 (N_9582,N_9318,N_9337);
xnor U9583 (N_9583,N_9294,N_9256);
nor U9584 (N_9584,N_9330,N_9328);
nand U9585 (N_9585,N_9383,N_9461);
and U9586 (N_9586,N_9308,N_9492);
or U9587 (N_9587,N_9342,N_9419);
nand U9588 (N_9588,N_9373,N_9499);
and U9589 (N_9589,N_9376,N_9257);
nand U9590 (N_9590,N_9442,N_9300);
xor U9591 (N_9591,N_9468,N_9459);
xnor U9592 (N_9592,N_9414,N_9252);
nand U9593 (N_9593,N_9334,N_9456);
and U9594 (N_9594,N_9260,N_9293);
and U9595 (N_9595,N_9283,N_9427);
and U9596 (N_9596,N_9331,N_9447);
and U9597 (N_9597,N_9351,N_9352);
or U9598 (N_9598,N_9264,N_9326);
or U9599 (N_9599,N_9306,N_9341);
nor U9600 (N_9600,N_9369,N_9498);
xnor U9601 (N_9601,N_9329,N_9413);
or U9602 (N_9602,N_9426,N_9357);
xor U9603 (N_9603,N_9295,N_9458);
xor U9604 (N_9604,N_9267,N_9396);
nand U9605 (N_9605,N_9310,N_9386);
nand U9606 (N_9606,N_9350,N_9484);
or U9607 (N_9607,N_9395,N_9481);
xor U9608 (N_9608,N_9353,N_9424);
or U9609 (N_9609,N_9311,N_9394);
xor U9610 (N_9610,N_9402,N_9362);
or U9611 (N_9611,N_9288,N_9346);
xnor U9612 (N_9612,N_9361,N_9371);
or U9613 (N_9613,N_9478,N_9339);
xor U9614 (N_9614,N_9277,N_9292);
nand U9615 (N_9615,N_9359,N_9488);
and U9616 (N_9616,N_9432,N_9482);
nor U9617 (N_9617,N_9439,N_9420);
nand U9618 (N_9618,N_9284,N_9289);
xnor U9619 (N_9619,N_9343,N_9327);
nand U9620 (N_9620,N_9430,N_9467);
xor U9621 (N_9621,N_9296,N_9453);
or U9622 (N_9622,N_9381,N_9276);
and U9623 (N_9623,N_9448,N_9435);
xor U9624 (N_9624,N_9325,N_9302);
nand U9625 (N_9625,N_9426,N_9486);
xnor U9626 (N_9626,N_9396,N_9476);
or U9627 (N_9627,N_9370,N_9399);
or U9628 (N_9628,N_9425,N_9407);
nor U9629 (N_9629,N_9452,N_9420);
nand U9630 (N_9630,N_9408,N_9485);
xnor U9631 (N_9631,N_9369,N_9253);
or U9632 (N_9632,N_9398,N_9444);
xnor U9633 (N_9633,N_9476,N_9366);
or U9634 (N_9634,N_9387,N_9345);
or U9635 (N_9635,N_9486,N_9447);
xnor U9636 (N_9636,N_9454,N_9387);
or U9637 (N_9637,N_9367,N_9396);
xor U9638 (N_9638,N_9393,N_9350);
or U9639 (N_9639,N_9485,N_9302);
xnor U9640 (N_9640,N_9461,N_9430);
or U9641 (N_9641,N_9282,N_9477);
nor U9642 (N_9642,N_9373,N_9407);
or U9643 (N_9643,N_9319,N_9442);
and U9644 (N_9644,N_9275,N_9351);
xor U9645 (N_9645,N_9381,N_9416);
nand U9646 (N_9646,N_9281,N_9442);
xnor U9647 (N_9647,N_9434,N_9424);
and U9648 (N_9648,N_9383,N_9394);
and U9649 (N_9649,N_9409,N_9318);
and U9650 (N_9650,N_9356,N_9259);
xnor U9651 (N_9651,N_9382,N_9415);
nor U9652 (N_9652,N_9400,N_9480);
nor U9653 (N_9653,N_9443,N_9375);
or U9654 (N_9654,N_9415,N_9326);
nor U9655 (N_9655,N_9454,N_9419);
nand U9656 (N_9656,N_9321,N_9256);
or U9657 (N_9657,N_9445,N_9383);
nand U9658 (N_9658,N_9417,N_9337);
nor U9659 (N_9659,N_9361,N_9384);
and U9660 (N_9660,N_9497,N_9383);
or U9661 (N_9661,N_9478,N_9360);
nand U9662 (N_9662,N_9491,N_9392);
nor U9663 (N_9663,N_9493,N_9339);
and U9664 (N_9664,N_9286,N_9444);
and U9665 (N_9665,N_9319,N_9475);
or U9666 (N_9666,N_9428,N_9487);
nor U9667 (N_9667,N_9409,N_9466);
nor U9668 (N_9668,N_9348,N_9256);
xnor U9669 (N_9669,N_9419,N_9464);
and U9670 (N_9670,N_9424,N_9278);
nor U9671 (N_9671,N_9354,N_9382);
nor U9672 (N_9672,N_9268,N_9314);
and U9673 (N_9673,N_9312,N_9320);
and U9674 (N_9674,N_9388,N_9311);
or U9675 (N_9675,N_9444,N_9381);
xnor U9676 (N_9676,N_9434,N_9464);
nand U9677 (N_9677,N_9378,N_9450);
nor U9678 (N_9678,N_9460,N_9468);
and U9679 (N_9679,N_9419,N_9335);
nand U9680 (N_9680,N_9279,N_9432);
or U9681 (N_9681,N_9461,N_9443);
and U9682 (N_9682,N_9490,N_9363);
xnor U9683 (N_9683,N_9367,N_9448);
nand U9684 (N_9684,N_9341,N_9318);
or U9685 (N_9685,N_9476,N_9395);
nand U9686 (N_9686,N_9347,N_9470);
xnor U9687 (N_9687,N_9408,N_9262);
or U9688 (N_9688,N_9368,N_9302);
nor U9689 (N_9689,N_9477,N_9273);
xnor U9690 (N_9690,N_9470,N_9408);
and U9691 (N_9691,N_9409,N_9306);
nand U9692 (N_9692,N_9397,N_9278);
or U9693 (N_9693,N_9337,N_9328);
nor U9694 (N_9694,N_9303,N_9397);
nand U9695 (N_9695,N_9427,N_9396);
nand U9696 (N_9696,N_9339,N_9467);
xnor U9697 (N_9697,N_9321,N_9450);
xnor U9698 (N_9698,N_9404,N_9366);
nor U9699 (N_9699,N_9290,N_9314);
or U9700 (N_9700,N_9365,N_9386);
nor U9701 (N_9701,N_9401,N_9428);
xnor U9702 (N_9702,N_9466,N_9480);
or U9703 (N_9703,N_9453,N_9264);
or U9704 (N_9704,N_9330,N_9460);
and U9705 (N_9705,N_9497,N_9343);
or U9706 (N_9706,N_9320,N_9477);
nor U9707 (N_9707,N_9469,N_9260);
or U9708 (N_9708,N_9476,N_9481);
or U9709 (N_9709,N_9273,N_9332);
nand U9710 (N_9710,N_9468,N_9329);
nand U9711 (N_9711,N_9394,N_9320);
or U9712 (N_9712,N_9416,N_9276);
nand U9713 (N_9713,N_9343,N_9486);
nand U9714 (N_9714,N_9423,N_9492);
and U9715 (N_9715,N_9414,N_9493);
and U9716 (N_9716,N_9468,N_9390);
xnor U9717 (N_9717,N_9306,N_9326);
nor U9718 (N_9718,N_9268,N_9356);
and U9719 (N_9719,N_9293,N_9488);
nand U9720 (N_9720,N_9452,N_9270);
nor U9721 (N_9721,N_9289,N_9472);
xnor U9722 (N_9722,N_9262,N_9255);
xor U9723 (N_9723,N_9303,N_9471);
nand U9724 (N_9724,N_9349,N_9418);
and U9725 (N_9725,N_9377,N_9287);
xor U9726 (N_9726,N_9295,N_9454);
nand U9727 (N_9727,N_9367,N_9277);
nand U9728 (N_9728,N_9344,N_9334);
xor U9729 (N_9729,N_9258,N_9481);
nand U9730 (N_9730,N_9376,N_9472);
nor U9731 (N_9731,N_9421,N_9322);
nand U9732 (N_9732,N_9437,N_9492);
xor U9733 (N_9733,N_9364,N_9350);
xor U9734 (N_9734,N_9385,N_9257);
xor U9735 (N_9735,N_9403,N_9287);
or U9736 (N_9736,N_9272,N_9311);
nor U9737 (N_9737,N_9283,N_9465);
xor U9738 (N_9738,N_9370,N_9379);
nand U9739 (N_9739,N_9389,N_9349);
nor U9740 (N_9740,N_9497,N_9310);
nor U9741 (N_9741,N_9313,N_9496);
nor U9742 (N_9742,N_9492,N_9341);
nor U9743 (N_9743,N_9439,N_9494);
or U9744 (N_9744,N_9466,N_9472);
or U9745 (N_9745,N_9484,N_9417);
or U9746 (N_9746,N_9331,N_9424);
or U9747 (N_9747,N_9389,N_9442);
or U9748 (N_9748,N_9303,N_9264);
xnor U9749 (N_9749,N_9296,N_9488);
xnor U9750 (N_9750,N_9557,N_9663);
and U9751 (N_9751,N_9556,N_9514);
and U9752 (N_9752,N_9725,N_9694);
nor U9753 (N_9753,N_9649,N_9540);
xnor U9754 (N_9754,N_9526,N_9722);
xnor U9755 (N_9755,N_9544,N_9515);
xor U9756 (N_9756,N_9594,N_9703);
xor U9757 (N_9757,N_9569,N_9706);
xor U9758 (N_9758,N_9713,N_9584);
xnor U9759 (N_9759,N_9736,N_9677);
or U9760 (N_9760,N_9599,N_9721);
and U9761 (N_9761,N_9534,N_9665);
or U9762 (N_9762,N_9545,N_9678);
nand U9763 (N_9763,N_9620,N_9605);
and U9764 (N_9764,N_9589,N_9704);
xor U9765 (N_9765,N_9598,N_9558);
and U9766 (N_9766,N_9525,N_9710);
nand U9767 (N_9767,N_9614,N_9524);
or U9768 (N_9768,N_9565,N_9746);
nor U9769 (N_9769,N_9607,N_9550);
xnor U9770 (N_9770,N_9689,N_9730);
nand U9771 (N_9771,N_9538,N_9692);
nand U9772 (N_9772,N_9747,N_9674);
nor U9773 (N_9773,N_9502,N_9669);
and U9774 (N_9774,N_9517,N_9571);
and U9775 (N_9775,N_9521,N_9657);
nor U9776 (N_9776,N_9593,N_9727);
or U9777 (N_9777,N_9734,N_9530);
nor U9778 (N_9778,N_9523,N_9716);
nand U9779 (N_9779,N_9611,N_9509);
nand U9780 (N_9780,N_9744,N_9682);
and U9781 (N_9781,N_9615,N_9673);
nand U9782 (N_9782,N_9576,N_9539);
xor U9783 (N_9783,N_9741,N_9648);
xor U9784 (N_9784,N_9554,N_9723);
or U9785 (N_9785,N_9552,N_9695);
nand U9786 (N_9786,N_9645,N_9728);
and U9787 (N_9787,N_9715,N_9564);
and U9788 (N_9788,N_9653,N_9572);
nand U9789 (N_9789,N_9619,N_9661);
xor U9790 (N_9790,N_9548,N_9560);
nand U9791 (N_9791,N_9688,N_9547);
nor U9792 (N_9792,N_9628,N_9519);
nand U9793 (N_9793,N_9513,N_9623);
or U9794 (N_9794,N_9506,N_9726);
or U9795 (N_9795,N_9701,N_9585);
and U9796 (N_9796,N_9510,N_9529);
nor U9797 (N_9797,N_9604,N_9575);
nand U9798 (N_9798,N_9672,N_9697);
nand U9799 (N_9799,N_9738,N_9633);
nor U9800 (N_9800,N_9651,N_9566);
nor U9801 (N_9801,N_9596,N_9543);
and U9802 (N_9802,N_9501,N_9700);
nand U9803 (N_9803,N_9608,N_9711);
xor U9804 (N_9804,N_9606,N_9717);
xnor U9805 (N_9805,N_9659,N_9743);
or U9806 (N_9806,N_9505,N_9642);
xnor U9807 (N_9807,N_9570,N_9581);
nand U9808 (N_9808,N_9504,N_9537);
or U9809 (N_9809,N_9640,N_9650);
or U9810 (N_9810,N_9693,N_9641);
and U9811 (N_9811,N_9612,N_9508);
nor U9812 (N_9812,N_9527,N_9626);
and U9813 (N_9813,N_9709,N_9740);
or U9814 (N_9814,N_9680,N_9691);
nor U9815 (N_9815,N_9532,N_9749);
and U9816 (N_9816,N_9559,N_9549);
xor U9817 (N_9817,N_9512,N_9616);
or U9818 (N_9818,N_9745,N_9541);
nor U9819 (N_9819,N_9568,N_9562);
or U9820 (N_9820,N_9702,N_9622);
xor U9821 (N_9821,N_9625,N_9518);
and U9822 (N_9822,N_9528,N_9500);
nor U9823 (N_9823,N_9655,N_9507);
xnor U9824 (N_9824,N_9601,N_9664);
nor U9825 (N_9825,N_9555,N_9573);
and U9826 (N_9826,N_9613,N_9712);
nor U9827 (N_9827,N_9577,N_9643);
and U9828 (N_9828,N_9646,N_9578);
nand U9829 (N_9829,N_9729,N_9631);
nor U9830 (N_9830,N_9684,N_9748);
and U9831 (N_9831,N_9551,N_9536);
xnor U9832 (N_9832,N_9739,N_9676);
nor U9833 (N_9833,N_9635,N_9671);
xor U9834 (N_9834,N_9681,N_9636);
nand U9835 (N_9835,N_9658,N_9662);
xnor U9836 (N_9836,N_9731,N_9685);
nand U9837 (N_9837,N_9590,N_9667);
nor U9838 (N_9838,N_9602,N_9629);
or U9839 (N_9839,N_9574,N_9600);
and U9840 (N_9840,N_9511,N_9597);
and U9841 (N_9841,N_9652,N_9719);
and U9842 (N_9842,N_9666,N_9621);
nor U9843 (N_9843,N_9546,N_9732);
or U9844 (N_9844,N_9624,N_9724);
and U9845 (N_9845,N_9656,N_9698);
nand U9846 (N_9846,N_9542,N_9668);
and U9847 (N_9847,N_9690,N_9603);
and U9848 (N_9848,N_9720,N_9634);
nor U9849 (N_9849,N_9583,N_9683);
and U9850 (N_9850,N_9718,N_9535);
or U9851 (N_9851,N_9660,N_9610);
and U9852 (N_9852,N_9707,N_9735);
xor U9853 (N_9853,N_9531,N_9579);
xnor U9854 (N_9854,N_9654,N_9737);
and U9855 (N_9855,N_9609,N_9586);
or U9856 (N_9856,N_9638,N_9533);
nand U9857 (N_9857,N_9675,N_9503);
or U9858 (N_9858,N_9617,N_9670);
nor U9859 (N_9859,N_9563,N_9618);
xor U9860 (N_9860,N_9522,N_9630);
or U9861 (N_9861,N_9647,N_9637);
or U9862 (N_9862,N_9582,N_9580);
nand U9863 (N_9863,N_9699,N_9742);
nor U9864 (N_9864,N_9567,N_9686);
or U9865 (N_9865,N_9520,N_9714);
or U9866 (N_9866,N_9516,N_9696);
nand U9867 (N_9867,N_9592,N_9587);
and U9868 (N_9868,N_9708,N_9588);
nor U9869 (N_9869,N_9644,N_9595);
and U9870 (N_9870,N_9705,N_9553);
nor U9871 (N_9871,N_9639,N_9627);
and U9872 (N_9872,N_9687,N_9591);
nand U9873 (N_9873,N_9733,N_9561);
and U9874 (N_9874,N_9632,N_9679);
xor U9875 (N_9875,N_9697,N_9623);
nand U9876 (N_9876,N_9571,N_9710);
nor U9877 (N_9877,N_9706,N_9511);
xor U9878 (N_9878,N_9541,N_9585);
nor U9879 (N_9879,N_9688,N_9502);
xnor U9880 (N_9880,N_9605,N_9526);
nand U9881 (N_9881,N_9541,N_9740);
or U9882 (N_9882,N_9706,N_9748);
nand U9883 (N_9883,N_9610,N_9671);
nor U9884 (N_9884,N_9637,N_9700);
or U9885 (N_9885,N_9514,N_9541);
nand U9886 (N_9886,N_9740,N_9508);
nand U9887 (N_9887,N_9587,N_9718);
and U9888 (N_9888,N_9701,N_9678);
nand U9889 (N_9889,N_9629,N_9639);
and U9890 (N_9890,N_9606,N_9654);
nor U9891 (N_9891,N_9540,N_9589);
xnor U9892 (N_9892,N_9514,N_9668);
and U9893 (N_9893,N_9679,N_9524);
nand U9894 (N_9894,N_9500,N_9575);
or U9895 (N_9895,N_9507,N_9563);
or U9896 (N_9896,N_9636,N_9569);
xor U9897 (N_9897,N_9666,N_9734);
nand U9898 (N_9898,N_9612,N_9509);
nor U9899 (N_9899,N_9571,N_9544);
and U9900 (N_9900,N_9632,N_9582);
and U9901 (N_9901,N_9666,N_9722);
or U9902 (N_9902,N_9638,N_9612);
or U9903 (N_9903,N_9603,N_9545);
nor U9904 (N_9904,N_9627,N_9606);
or U9905 (N_9905,N_9706,N_9679);
and U9906 (N_9906,N_9699,N_9679);
and U9907 (N_9907,N_9742,N_9599);
xor U9908 (N_9908,N_9741,N_9581);
nor U9909 (N_9909,N_9693,N_9618);
nand U9910 (N_9910,N_9740,N_9548);
xor U9911 (N_9911,N_9682,N_9733);
or U9912 (N_9912,N_9534,N_9529);
and U9913 (N_9913,N_9702,N_9618);
nand U9914 (N_9914,N_9588,N_9602);
or U9915 (N_9915,N_9643,N_9532);
and U9916 (N_9916,N_9522,N_9729);
nor U9917 (N_9917,N_9628,N_9696);
nand U9918 (N_9918,N_9733,N_9635);
nor U9919 (N_9919,N_9664,N_9551);
xnor U9920 (N_9920,N_9601,N_9597);
nand U9921 (N_9921,N_9689,N_9741);
and U9922 (N_9922,N_9617,N_9539);
xor U9923 (N_9923,N_9641,N_9568);
and U9924 (N_9924,N_9723,N_9523);
nand U9925 (N_9925,N_9715,N_9747);
and U9926 (N_9926,N_9582,N_9570);
xor U9927 (N_9927,N_9649,N_9622);
or U9928 (N_9928,N_9634,N_9581);
and U9929 (N_9929,N_9598,N_9507);
xnor U9930 (N_9930,N_9637,N_9612);
and U9931 (N_9931,N_9703,N_9536);
xor U9932 (N_9932,N_9715,N_9675);
nor U9933 (N_9933,N_9601,N_9534);
nand U9934 (N_9934,N_9662,N_9532);
nand U9935 (N_9935,N_9542,N_9739);
and U9936 (N_9936,N_9701,N_9723);
nor U9937 (N_9937,N_9733,N_9662);
and U9938 (N_9938,N_9553,N_9684);
xor U9939 (N_9939,N_9516,N_9593);
and U9940 (N_9940,N_9675,N_9701);
xor U9941 (N_9941,N_9570,N_9511);
nand U9942 (N_9942,N_9582,N_9593);
nor U9943 (N_9943,N_9591,N_9637);
xnor U9944 (N_9944,N_9729,N_9500);
xnor U9945 (N_9945,N_9658,N_9714);
xor U9946 (N_9946,N_9669,N_9608);
and U9947 (N_9947,N_9514,N_9553);
or U9948 (N_9948,N_9706,N_9613);
nand U9949 (N_9949,N_9507,N_9649);
nor U9950 (N_9950,N_9626,N_9545);
nor U9951 (N_9951,N_9686,N_9723);
nor U9952 (N_9952,N_9607,N_9615);
xor U9953 (N_9953,N_9534,N_9500);
nor U9954 (N_9954,N_9662,N_9551);
or U9955 (N_9955,N_9725,N_9562);
or U9956 (N_9956,N_9646,N_9527);
xnor U9957 (N_9957,N_9587,N_9507);
or U9958 (N_9958,N_9607,N_9595);
nor U9959 (N_9959,N_9526,N_9556);
and U9960 (N_9960,N_9533,N_9582);
and U9961 (N_9961,N_9526,N_9508);
nor U9962 (N_9962,N_9639,N_9608);
or U9963 (N_9963,N_9567,N_9500);
and U9964 (N_9964,N_9571,N_9699);
xnor U9965 (N_9965,N_9727,N_9541);
nand U9966 (N_9966,N_9510,N_9597);
nor U9967 (N_9967,N_9666,N_9612);
nor U9968 (N_9968,N_9584,N_9556);
xnor U9969 (N_9969,N_9565,N_9581);
and U9970 (N_9970,N_9630,N_9504);
xnor U9971 (N_9971,N_9717,N_9646);
nand U9972 (N_9972,N_9550,N_9533);
xor U9973 (N_9973,N_9716,N_9505);
xnor U9974 (N_9974,N_9553,N_9725);
or U9975 (N_9975,N_9665,N_9609);
or U9976 (N_9976,N_9733,N_9584);
nor U9977 (N_9977,N_9701,N_9550);
xnor U9978 (N_9978,N_9640,N_9700);
nand U9979 (N_9979,N_9721,N_9580);
and U9980 (N_9980,N_9584,N_9633);
or U9981 (N_9981,N_9535,N_9509);
or U9982 (N_9982,N_9583,N_9511);
nand U9983 (N_9983,N_9530,N_9670);
xnor U9984 (N_9984,N_9562,N_9746);
nor U9985 (N_9985,N_9719,N_9642);
xnor U9986 (N_9986,N_9637,N_9508);
or U9987 (N_9987,N_9654,N_9599);
nand U9988 (N_9988,N_9583,N_9634);
and U9989 (N_9989,N_9664,N_9518);
nand U9990 (N_9990,N_9683,N_9559);
nor U9991 (N_9991,N_9637,N_9692);
xnor U9992 (N_9992,N_9632,N_9700);
nand U9993 (N_9993,N_9674,N_9648);
xnor U9994 (N_9994,N_9736,N_9618);
or U9995 (N_9995,N_9556,N_9621);
nand U9996 (N_9996,N_9700,N_9517);
or U9997 (N_9997,N_9747,N_9698);
nand U9998 (N_9998,N_9698,N_9524);
nand U9999 (N_9999,N_9567,N_9653);
or U10000 (N_10000,N_9794,N_9950);
and U10001 (N_10001,N_9901,N_9852);
nor U10002 (N_10002,N_9966,N_9894);
nor U10003 (N_10003,N_9898,N_9890);
and U10004 (N_10004,N_9913,N_9795);
and U10005 (N_10005,N_9833,N_9844);
nand U10006 (N_10006,N_9881,N_9955);
nor U10007 (N_10007,N_9767,N_9836);
or U10008 (N_10008,N_9939,N_9991);
nor U10009 (N_10009,N_9778,N_9785);
xnor U10010 (N_10010,N_9758,N_9906);
nand U10011 (N_10011,N_9809,N_9921);
and U10012 (N_10012,N_9801,N_9864);
or U10013 (N_10013,N_9851,N_9806);
nand U10014 (N_10014,N_9958,N_9755);
or U10015 (N_10015,N_9764,N_9793);
or U10016 (N_10016,N_9997,N_9896);
nor U10017 (N_10017,N_9872,N_9902);
nor U10018 (N_10018,N_9891,N_9775);
or U10019 (N_10019,N_9944,N_9818);
or U10020 (N_10020,N_9976,N_9859);
or U10021 (N_10021,N_9879,N_9756);
nand U10022 (N_10022,N_9998,N_9798);
or U10023 (N_10023,N_9931,N_9771);
nor U10024 (N_10024,N_9762,N_9834);
xnor U10025 (N_10025,N_9912,N_9935);
or U10026 (N_10026,N_9880,N_9781);
or U10027 (N_10027,N_9923,N_9845);
or U10028 (N_10028,N_9970,N_9920);
nor U10029 (N_10029,N_9811,N_9900);
xor U10030 (N_10030,N_9968,N_9768);
nor U10031 (N_10031,N_9849,N_9910);
nor U10032 (N_10032,N_9788,N_9804);
and U10033 (N_10033,N_9817,N_9808);
nand U10034 (N_10034,N_9927,N_9919);
and U10035 (N_10035,N_9951,N_9870);
xor U10036 (N_10036,N_9986,N_9909);
xor U10037 (N_10037,N_9994,N_9942);
or U10038 (N_10038,N_9992,N_9996);
and U10039 (N_10039,N_9974,N_9869);
or U10040 (N_10040,N_9751,N_9792);
nor U10041 (N_10041,N_9757,N_9763);
nand U10042 (N_10042,N_9791,N_9874);
xor U10043 (N_10043,N_9984,N_9774);
nand U10044 (N_10044,N_9819,N_9895);
and U10045 (N_10045,N_9789,N_9948);
nor U10046 (N_10046,N_9828,N_9832);
nand U10047 (N_10047,N_9882,N_9892);
or U10048 (N_10048,N_9903,N_9853);
or U10049 (N_10049,N_9776,N_9982);
nor U10050 (N_10050,N_9868,N_9945);
or U10051 (N_10051,N_9954,N_9761);
and U10052 (N_10052,N_9752,N_9972);
nand U10053 (N_10053,N_9887,N_9889);
nand U10054 (N_10054,N_9928,N_9765);
or U10055 (N_10055,N_9782,N_9835);
or U10056 (N_10056,N_9941,N_9797);
or U10057 (N_10057,N_9799,N_9911);
and U10058 (N_10058,N_9871,N_9964);
and U10059 (N_10059,N_9899,N_9924);
and U10060 (N_10060,N_9875,N_9916);
nor U10061 (N_10061,N_9783,N_9884);
and U10062 (N_10062,N_9957,N_9814);
nand U10063 (N_10063,N_9883,N_9938);
xnor U10064 (N_10064,N_9960,N_9946);
and U10065 (N_10065,N_9971,N_9780);
xnor U10066 (N_10066,N_9842,N_9815);
nor U10067 (N_10067,N_9926,N_9840);
and U10068 (N_10068,N_9772,N_9934);
or U10069 (N_10069,N_9933,N_9973);
nor U10070 (N_10070,N_9850,N_9787);
or U10071 (N_10071,N_9800,N_9848);
xor U10072 (N_10072,N_9753,N_9965);
nor U10073 (N_10073,N_9918,N_9861);
or U10074 (N_10074,N_9867,N_9925);
nor U10075 (N_10075,N_9857,N_9963);
nor U10076 (N_10076,N_9988,N_9786);
and U10077 (N_10077,N_9952,N_9784);
and U10078 (N_10078,N_9810,N_9812);
or U10079 (N_10079,N_9846,N_9929);
or U10080 (N_10080,N_9807,N_9978);
xor U10081 (N_10081,N_9820,N_9908);
nor U10082 (N_10082,N_9805,N_9979);
or U10083 (N_10083,N_9914,N_9995);
and U10084 (N_10084,N_9754,N_9823);
nor U10085 (N_10085,N_9888,N_9987);
and U10086 (N_10086,N_9940,N_9837);
xnor U10087 (N_10087,N_9897,N_9821);
or U10088 (N_10088,N_9862,N_9905);
and U10089 (N_10089,N_9930,N_9766);
xnor U10090 (N_10090,N_9779,N_9824);
nand U10091 (N_10091,N_9777,N_9981);
nand U10092 (N_10092,N_9983,N_9773);
or U10093 (N_10093,N_9949,N_9885);
or U10094 (N_10094,N_9796,N_9989);
or U10095 (N_10095,N_9838,N_9839);
xnor U10096 (N_10096,N_9854,N_9993);
or U10097 (N_10097,N_9877,N_9863);
and U10098 (N_10098,N_9865,N_9825);
nand U10099 (N_10099,N_9943,N_9855);
xor U10100 (N_10100,N_9790,N_9967);
xor U10101 (N_10101,N_9760,N_9830);
and U10102 (N_10102,N_9962,N_9816);
nand U10103 (N_10103,N_9917,N_9866);
nand U10104 (N_10104,N_9841,N_9750);
xor U10105 (N_10105,N_9907,N_9769);
xor U10106 (N_10106,N_9827,N_9936);
nand U10107 (N_10107,N_9904,N_9975);
nor U10108 (N_10108,N_9915,N_9980);
nor U10109 (N_10109,N_9826,N_9937);
nand U10110 (N_10110,N_9873,N_9860);
or U10111 (N_10111,N_9831,N_9803);
or U10112 (N_10112,N_9893,N_9956);
nor U10113 (N_10113,N_9922,N_9843);
and U10114 (N_10114,N_9959,N_9886);
or U10115 (N_10115,N_9822,N_9858);
nor U10116 (N_10116,N_9802,N_9999);
xor U10117 (N_10117,N_9759,N_9829);
xnor U10118 (N_10118,N_9770,N_9876);
and U10119 (N_10119,N_9856,N_9947);
and U10120 (N_10120,N_9985,N_9969);
nand U10121 (N_10121,N_9932,N_9961);
nand U10122 (N_10122,N_9953,N_9990);
xnor U10123 (N_10123,N_9847,N_9977);
and U10124 (N_10124,N_9878,N_9813);
or U10125 (N_10125,N_9846,N_9967);
and U10126 (N_10126,N_9952,N_9839);
nand U10127 (N_10127,N_9979,N_9797);
and U10128 (N_10128,N_9967,N_9944);
nand U10129 (N_10129,N_9868,N_9849);
nor U10130 (N_10130,N_9882,N_9788);
and U10131 (N_10131,N_9884,N_9919);
xor U10132 (N_10132,N_9856,N_9939);
xor U10133 (N_10133,N_9831,N_9977);
or U10134 (N_10134,N_9791,N_9913);
nor U10135 (N_10135,N_9967,N_9762);
or U10136 (N_10136,N_9820,N_9759);
nand U10137 (N_10137,N_9924,N_9812);
nor U10138 (N_10138,N_9820,N_9860);
and U10139 (N_10139,N_9940,N_9810);
nor U10140 (N_10140,N_9928,N_9815);
nand U10141 (N_10141,N_9931,N_9945);
xnor U10142 (N_10142,N_9870,N_9982);
and U10143 (N_10143,N_9792,N_9856);
xor U10144 (N_10144,N_9865,N_9971);
nor U10145 (N_10145,N_9798,N_9930);
xnor U10146 (N_10146,N_9855,N_9822);
xnor U10147 (N_10147,N_9916,N_9884);
xnor U10148 (N_10148,N_9937,N_9750);
and U10149 (N_10149,N_9798,N_9821);
nor U10150 (N_10150,N_9868,N_9795);
nor U10151 (N_10151,N_9811,N_9823);
nor U10152 (N_10152,N_9923,N_9926);
and U10153 (N_10153,N_9789,N_9803);
nand U10154 (N_10154,N_9963,N_9988);
or U10155 (N_10155,N_9819,N_9944);
xor U10156 (N_10156,N_9813,N_9962);
xor U10157 (N_10157,N_9921,N_9879);
nand U10158 (N_10158,N_9875,N_9812);
or U10159 (N_10159,N_9967,N_9764);
nor U10160 (N_10160,N_9750,N_9971);
xnor U10161 (N_10161,N_9778,N_9887);
and U10162 (N_10162,N_9807,N_9815);
or U10163 (N_10163,N_9964,N_9947);
and U10164 (N_10164,N_9761,N_9805);
xor U10165 (N_10165,N_9954,N_9856);
xnor U10166 (N_10166,N_9802,N_9918);
nand U10167 (N_10167,N_9844,N_9892);
or U10168 (N_10168,N_9828,N_9895);
and U10169 (N_10169,N_9862,N_9915);
nand U10170 (N_10170,N_9796,N_9836);
or U10171 (N_10171,N_9770,N_9825);
nor U10172 (N_10172,N_9861,N_9931);
and U10173 (N_10173,N_9884,N_9973);
nor U10174 (N_10174,N_9804,N_9922);
nor U10175 (N_10175,N_9913,N_9773);
nor U10176 (N_10176,N_9956,N_9909);
nor U10177 (N_10177,N_9783,N_9955);
xor U10178 (N_10178,N_9901,N_9853);
and U10179 (N_10179,N_9964,N_9765);
xnor U10180 (N_10180,N_9781,N_9877);
nor U10181 (N_10181,N_9992,N_9755);
or U10182 (N_10182,N_9782,N_9999);
nor U10183 (N_10183,N_9940,N_9770);
or U10184 (N_10184,N_9907,N_9775);
and U10185 (N_10185,N_9930,N_9882);
nand U10186 (N_10186,N_9828,N_9868);
xnor U10187 (N_10187,N_9779,N_9992);
and U10188 (N_10188,N_9977,N_9818);
and U10189 (N_10189,N_9973,N_9866);
or U10190 (N_10190,N_9941,N_9950);
nand U10191 (N_10191,N_9953,N_9938);
and U10192 (N_10192,N_9792,N_9805);
or U10193 (N_10193,N_9922,N_9818);
and U10194 (N_10194,N_9871,N_9806);
nor U10195 (N_10195,N_9999,N_9832);
nor U10196 (N_10196,N_9843,N_9996);
xnor U10197 (N_10197,N_9970,N_9932);
nand U10198 (N_10198,N_9902,N_9893);
and U10199 (N_10199,N_9853,N_9876);
nand U10200 (N_10200,N_9884,N_9983);
xnor U10201 (N_10201,N_9939,N_9914);
and U10202 (N_10202,N_9964,N_9934);
nand U10203 (N_10203,N_9804,N_9840);
xor U10204 (N_10204,N_9810,N_9826);
xor U10205 (N_10205,N_9940,N_9806);
nand U10206 (N_10206,N_9773,N_9803);
and U10207 (N_10207,N_9843,N_9944);
nand U10208 (N_10208,N_9830,N_9828);
or U10209 (N_10209,N_9750,N_9952);
and U10210 (N_10210,N_9750,N_9759);
and U10211 (N_10211,N_9998,N_9781);
nand U10212 (N_10212,N_9907,N_9874);
nor U10213 (N_10213,N_9756,N_9787);
and U10214 (N_10214,N_9876,N_9960);
or U10215 (N_10215,N_9960,N_9797);
nor U10216 (N_10216,N_9925,N_9857);
nor U10217 (N_10217,N_9988,N_9999);
nor U10218 (N_10218,N_9852,N_9845);
and U10219 (N_10219,N_9868,N_9853);
and U10220 (N_10220,N_9851,N_9786);
xnor U10221 (N_10221,N_9856,N_9974);
nand U10222 (N_10222,N_9983,N_9826);
xnor U10223 (N_10223,N_9949,N_9919);
and U10224 (N_10224,N_9846,N_9860);
or U10225 (N_10225,N_9933,N_9802);
nand U10226 (N_10226,N_9838,N_9951);
and U10227 (N_10227,N_9998,N_9945);
nor U10228 (N_10228,N_9759,N_9913);
and U10229 (N_10229,N_9821,N_9962);
nor U10230 (N_10230,N_9919,N_9908);
xnor U10231 (N_10231,N_9817,N_9965);
and U10232 (N_10232,N_9977,N_9920);
and U10233 (N_10233,N_9758,N_9936);
and U10234 (N_10234,N_9832,N_9757);
nor U10235 (N_10235,N_9752,N_9784);
nor U10236 (N_10236,N_9861,N_9954);
and U10237 (N_10237,N_9870,N_9877);
xnor U10238 (N_10238,N_9780,N_9787);
nand U10239 (N_10239,N_9762,N_9879);
nor U10240 (N_10240,N_9941,N_9765);
and U10241 (N_10241,N_9828,N_9887);
and U10242 (N_10242,N_9833,N_9798);
nor U10243 (N_10243,N_9876,N_9785);
or U10244 (N_10244,N_9774,N_9754);
nor U10245 (N_10245,N_9773,N_9844);
nand U10246 (N_10246,N_9975,N_9796);
xor U10247 (N_10247,N_9986,N_9914);
nor U10248 (N_10248,N_9826,N_9807);
or U10249 (N_10249,N_9892,N_9782);
xor U10250 (N_10250,N_10222,N_10226);
nor U10251 (N_10251,N_10164,N_10017);
nand U10252 (N_10252,N_10086,N_10154);
xnor U10253 (N_10253,N_10053,N_10241);
and U10254 (N_10254,N_10166,N_10149);
or U10255 (N_10255,N_10189,N_10143);
nand U10256 (N_10256,N_10106,N_10192);
nand U10257 (N_10257,N_10119,N_10141);
nor U10258 (N_10258,N_10081,N_10209);
nand U10259 (N_10259,N_10133,N_10180);
and U10260 (N_10260,N_10032,N_10153);
and U10261 (N_10261,N_10083,N_10142);
nand U10262 (N_10262,N_10107,N_10056);
xor U10263 (N_10263,N_10093,N_10128);
xnor U10264 (N_10264,N_10167,N_10203);
and U10265 (N_10265,N_10240,N_10194);
and U10266 (N_10266,N_10113,N_10054);
or U10267 (N_10267,N_10176,N_10048);
nor U10268 (N_10268,N_10188,N_10012);
and U10269 (N_10269,N_10109,N_10156);
nor U10270 (N_10270,N_10218,N_10144);
or U10271 (N_10271,N_10233,N_10137);
and U10272 (N_10272,N_10232,N_10059);
nor U10273 (N_10273,N_10094,N_10158);
nand U10274 (N_10274,N_10000,N_10047);
xor U10275 (N_10275,N_10098,N_10221);
xor U10276 (N_10276,N_10183,N_10079);
and U10277 (N_10277,N_10147,N_10216);
and U10278 (N_10278,N_10114,N_10042);
or U10279 (N_10279,N_10127,N_10063);
nor U10280 (N_10280,N_10076,N_10135);
and U10281 (N_10281,N_10099,N_10084);
nor U10282 (N_10282,N_10088,N_10118);
xor U10283 (N_10283,N_10043,N_10219);
nand U10284 (N_10284,N_10136,N_10239);
xnor U10285 (N_10285,N_10037,N_10130);
xor U10286 (N_10286,N_10125,N_10033);
nor U10287 (N_10287,N_10004,N_10195);
xnor U10288 (N_10288,N_10208,N_10184);
xor U10289 (N_10289,N_10001,N_10103);
or U10290 (N_10290,N_10065,N_10161);
or U10291 (N_10291,N_10248,N_10139);
or U10292 (N_10292,N_10020,N_10191);
xnor U10293 (N_10293,N_10117,N_10181);
nand U10294 (N_10294,N_10066,N_10148);
nor U10295 (N_10295,N_10186,N_10247);
or U10296 (N_10296,N_10110,N_10177);
or U10297 (N_10297,N_10105,N_10089);
and U10298 (N_10298,N_10249,N_10046);
nand U10299 (N_10299,N_10215,N_10067);
nand U10300 (N_10300,N_10040,N_10104);
xnor U10301 (N_10301,N_10039,N_10034);
nor U10302 (N_10302,N_10058,N_10070);
nor U10303 (N_10303,N_10224,N_10207);
nor U10304 (N_10304,N_10078,N_10024);
nand U10305 (N_10305,N_10011,N_10129);
nand U10306 (N_10306,N_10073,N_10102);
or U10307 (N_10307,N_10175,N_10008);
nor U10308 (N_10308,N_10100,N_10185);
and U10309 (N_10309,N_10213,N_10199);
nor U10310 (N_10310,N_10197,N_10202);
nand U10311 (N_10311,N_10036,N_10045);
and U10312 (N_10312,N_10155,N_10075);
nor U10313 (N_10313,N_10243,N_10055);
xnor U10314 (N_10314,N_10172,N_10237);
nand U10315 (N_10315,N_10205,N_10082);
xor U10316 (N_10316,N_10227,N_10007);
and U10317 (N_10317,N_10171,N_10235);
or U10318 (N_10318,N_10121,N_10112);
and U10319 (N_10319,N_10193,N_10234);
and U10320 (N_10320,N_10062,N_10090);
xnor U10321 (N_10321,N_10223,N_10101);
nand U10322 (N_10322,N_10246,N_10145);
or U10323 (N_10323,N_10072,N_10002);
xor U10324 (N_10324,N_10157,N_10214);
nand U10325 (N_10325,N_10092,N_10087);
and U10326 (N_10326,N_10010,N_10115);
xnor U10327 (N_10327,N_10051,N_10152);
and U10328 (N_10328,N_10169,N_10026);
or U10329 (N_10329,N_10061,N_10028);
or U10330 (N_10330,N_10069,N_10220);
nand U10331 (N_10331,N_10231,N_10242);
xor U10332 (N_10332,N_10206,N_10014);
or U10333 (N_10333,N_10116,N_10052);
and U10334 (N_10334,N_10124,N_10151);
and U10335 (N_10335,N_10132,N_10173);
nor U10336 (N_10336,N_10022,N_10038);
or U10337 (N_10337,N_10163,N_10120);
and U10338 (N_10338,N_10210,N_10013);
nor U10339 (N_10339,N_10174,N_10170);
and U10340 (N_10340,N_10126,N_10050);
and U10341 (N_10341,N_10035,N_10068);
xnor U10342 (N_10342,N_10091,N_10016);
nand U10343 (N_10343,N_10230,N_10044);
nor U10344 (N_10344,N_10168,N_10018);
nand U10345 (N_10345,N_10080,N_10030);
and U10346 (N_10346,N_10077,N_10182);
nand U10347 (N_10347,N_10111,N_10200);
nor U10348 (N_10348,N_10160,N_10029);
xor U10349 (N_10349,N_10123,N_10229);
nand U10350 (N_10350,N_10064,N_10005);
nor U10351 (N_10351,N_10041,N_10108);
xnor U10352 (N_10352,N_10134,N_10178);
xnor U10353 (N_10353,N_10196,N_10131);
and U10354 (N_10354,N_10228,N_10057);
nor U10355 (N_10355,N_10003,N_10165);
nand U10356 (N_10356,N_10244,N_10198);
xnor U10357 (N_10357,N_10074,N_10138);
nand U10358 (N_10358,N_10236,N_10015);
and U10359 (N_10359,N_10217,N_10122);
or U10360 (N_10360,N_10025,N_10140);
nand U10361 (N_10361,N_10006,N_10211);
and U10362 (N_10362,N_10023,N_10071);
nor U10363 (N_10363,N_10225,N_10238);
or U10364 (N_10364,N_10204,N_10019);
nand U10365 (N_10365,N_10097,N_10021);
xor U10366 (N_10366,N_10162,N_10159);
and U10367 (N_10367,N_10031,N_10179);
and U10368 (N_10368,N_10095,N_10060);
nand U10369 (N_10369,N_10190,N_10085);
xnor U10370 (N_10370,N_10245,N_10096);
and U10371 (N_10371,N_10150,N_10049);
xnor U10372 (N_10372,N_10146,N_10201);
xor U10373 (N_10373,N_10027,N_10187);
nor U10374 (N_10374,N_10009,N_10212);
or U10375 (N_10375,N_10226,N_10012);
and U10376 (N_10376,N_10124,N_10104);
and U10377 (N_10377,N_10181,N_10209);
or U10378 (N_10378,N_10224,N_10099);
nand U10379 (N_10379,N_10149,N_10063);
and U10380 (N_10380,N_10126,N_10180);
nand U10381 (N_10381,N_10080,N_10134);
or U10382 (N_10382,N_10145,N_10157);
and U10383 (N_10383,N_10051,N_10068);
or U10384 (N_10384,N_10245,N_10117);
nand U10385 (N_10385,N_10123,N_10067);
and U10386 (N_10386,N_10148,N_10132);
nand U10387 (N_10387,N_10074,N_10112);
nand U10388 (N_10388,N_10107,N_10063);
or U10389 (N_10389,N_10137,N_10033);
nand U10390 (N_10390,N_10178,N_10014);
or U10391 (N_10391,N_10182,N_10196);
nand U10392 (N_10392,N_10201,N_10094);
nor U10393 (N_10393,N_10118,N_10205);
xor U10394 (N_10394,N_10006,N_10199);
or U10395 (N_10395,N_10223,N_10111);
and U10396 (N_10396,N_10183,N_10022);
and U10397 (N_10397,N_10214,N_10040);
xor U10398 (N_10398,N_10151,N_10044);
or U10399 (N_10399,N_10059,N_10192);
xnor U10400 (N_10400,N_10064,N_10054);
and U10401 (N_10401,N_10053,N_10140);
nand U10402 (N_10402,N_10191,N_10091);
or U10403 (N_10403,N_10237,N_10028);
nand U10404 (N_10404,N_10094,N_10146);
and U10405 (N_10405,N_10195,N_10167);
xor U10406 (N_10406,N_10195,N_10217);
nor U10407 (N_10407,N_10160,N_10193);
and U10408 (N_10408,N_10104,N_10157);
and U10409 (N_10409,N_10095,N_10106);
nor U10410 (N_10410,N_10160,N_10139);
xor U10411 (N_10411,N_10002,N_10082);
xnor U10412 (N_10412,N_10125,N_10120);
and U10413 (N_10413,N_10018,N_10215);
nand U10414 (N_10414,N_10161,N_10018);
or U10415 (N_10415,N_10112,N_10100);
or U10416 (N_10416,N_10073,N_10157);
nor U10417 (N_10417,N_10199,N_10122);
and U10418 (N_10418,N_10124,N_10176);
xor U10419 (N_10419,N_10234,N_10238);
nand U10420 (N_10420,N_10143,N_10000);
or U10421 (N_10421,N_10150,N_10223);
xor U10422 (N_10422,N_10017,N_10061);
xnor U10423 (N_10423,N_10186,N_10066);
and U10424 (N_10424,N_10092,N_10134);
nor U10425 (N_10425,N_10180,N_10084);
xnor U10426 (N_10426,N_10224,N_10102);
and U10427 (N_10427,N_10128,N_10221);
nand U10428 (N_10428,N_10208,N_10175);
or U10429 (N_10429,N_10115,N_10210);
and U10430 (N_10430,N_10203,N_10107);
or U10431 (N_10431,N_10078,N_10089);
xor U10432 (N_10432,N_10048,N_10244);
or U10433 (N_10433,N_10079,N_10142);
xnor U10434 (N_10434,N_10034,N_10075);
and U10435 (N_10435,N_10041,N_10007);
or U10436 (N_10436,N_10149,N_10244);
xor U10437 (N_10437,N_10165,N_10184);
nor U10438 (N_10438,N_10035,N_10061);
nor U10439 (N_10439,N_10012,N_10076);
nor U10440 (N_10440,N_10249,N_10040);
and U10441 (N_10441,N_10128,N_10225);
or U10442 (N_10442,N_10076,N_10037);
or U10443 (N_10443,N_10244,N_10061);
or U10444 (N_10444,N_10210,N_10042);
and U10445 (N_10445,N_10094,N_10005);
and U10446 (N_10446,N_10074,N_10011);
or U10447 (N_10447,N_10054,N_10089);
xnor U10448 (N_10448,N_10113,N_10053);
nor U10449 (N_10449,N_10046,N_10223);
nand U10450 (N_10450,N_10181,N_10104);
or U10451 (N_10451,N_10165,N_10042);
nor U10452 (N_10452,N_10206,N_10130);
nand U10453 (N_10453,N_10053,N_10038);
or U10454 (N_10454,N_10093,N_10013);
nor U10455 (N_10455,N_10072,N_10119);
or U10456 (N_10456,N_10241,N_10088);
xor U10457 (N_10457,N_10008,N_10113);
and U10458 (N_10458,N_10149,N_10075);
nand U10459 (N_10459,N_10196,N_10233);
nand U10460 (N_10460,N_10101,N_10043);
nor U10461 (N_10461,N_10246,N_10071);
nor U10462 (N_10462,N_10005,N_10241);
nor U10463 (N_10463,N_10049,N_10126);
nor U10464 (N_10464,N_10100,N_10237);
xnor U10465 (N_10465,N_10191,N_10134);
xor U10466 (N_10466,N_10190,N_10106);
nand U10467 (N_10467,N_10033,N_10087);
nor U10468 (N_10468,N_10104,N_10176);
nand U10469 (N_10469,N_10136,N_10226);
xnor U10470 (N_10470,N_10245,N_10063);
or U10471 (N_10471,N_10004,N_10106);
xnor U10472 (N_10472,N_10117,N_10111);
and U10473 (N_10473,N_10014,N_10029);
xnor U10474 (N_10474,N_10024,N_10073);
and U10475 (N_10475,N_10122,N_10187);
nand U10476 (N_10476,N_10154,N_10068);
nand U10477 (N_10477,N_10246,N_10167);
or U10478 (N_10478,N_10013,N_10031);
nor U10479 (N_10479,N_10002,N_10058);
and U10480 (N_10480,N_10214,N_10218);
xnor U10481 (N_10481,N_10213,N_10215);
xor U10482 (N_10482,N_10112,N_10129);
nand U10483 (N_10483,N_10002,N_10118);
and U10484 (N_10484,N_10151,N_10003);
nor U10485 (N_10485,N_10079,N_10096);
and U10486 (N_10486,N_10166,N_10089);
nand U10487 (N_10487,N_10152,N_10002);
nor U10488 (N_10488,N_10092,N_10039);
or U10489 (N_10489,N_10196,N_10163);
xor U10490 (N_10490,N_10091,N_10212);
nand U10491 (N_10491,N_10071,N_10136);
or U10492 (N_10492,N_10230,N_10185);
xnor U10493 (N_10493,N_10070,N_10193);
nand U10494 (N_10494,N_10185,N_10152);
nor U10495 (N_10495,N_10066,N_10010);
nor U10496 (N_10496,N_10190,N_10126);
and U10497 (N_10497,N_10220,N_10244);
nor U10498 (N_10498,N_10228,N_10046);
nand U10499 (N_10499,N_10073,N_10000);
and U10500 (N_10500,N_10426,N_10450);
xnor U10501 (N_10501,N_10431,N_10447);
nand U10502 (N_10502,N_10365,N_10466);
nand U10503 (N_10503,N_10262,N_10328);
xnor U10504 (N_10504,N_10399,N_10290);
nor U10505 (N_10505,N_10321,N_10422);
nor U10506 (N_10506,N_10438,N_10303);
nor U10507 (N_10507,N_10344,N_10346);
and U10508 (N_10508,N_10332,N_10440);
or U10509 (N_10509,N_10498,N_10402);
or U10510 (N_10510,N_10458,N_10434);
and U10511 (N_10511,N_10260,N_10288);
nor U10512 (N_10512,N_10298,N_10472);
xor U10513 (N_10513,N_10490,N_10370);
or U10514 (N_10514,N_10377,N_10347);
or U10515 (N_10515,N_10295,N_10306);
and U10516 (N_10516,N_10488,N_10289);
xnor U10517 (N_10517,N_10425,N_10356);
nor U10518 (N_10518,N_10384,N_10334);
and U10519 (N_10519,N_10461,N_10291);
and U10520 (N_10520,N_10474,N_10368);
and U10521 (N_10521,N_10300,N_10312);
and U10522 (N_10522,N_10435,N_10318);
or U10523 (N_10523,N_10266,N_10371);
nand U10524 (N_10524,N_10385,N_10330);
nand U10525 (N_10525,N_10470,N_10489);
nor U10526 (N_10526,N_10427,N_10279);
or U10527 (N_10527,N_10468,N_10310);
nand U10528 (N_10528,N_10320,N_10374);
nor U10529 (N_10529,N_10309,N_10479);
and U10530 (N_10530,N_10454,N_10452);
or U10531 (N_10531,N_10381,N_10397);
or U10532 (N_10532,N_10456,N_10405);
or U10533 (N_10533,N_10305,N_10403);
nand U10534 (N_10534,N_10378,N_10409);
nor U10535 (N_10535,N_10299,N_10419);
xor U10536 (N_10536,N_10350,N_10449);
xnor U10537 (N_10537,N_10386,N_10296);
nand U10538 (N_10538,N_10392,N_10315);
xor U10539 (N_10539,N_10317,N_10388);
or U10540 (N_10540,N_10373,N_10398);
xnor U10541 (N_10541,N_10428,N_10429);
nor U10542 (N_10542,N_10311,N_10257);
nand U10543 (N_10543,N_10277,N_10275);
and U10544 (N_10544,N_10407,N_10437);
nand U10545 (N_10545,N_10343,N_10307);
nor U10546 (N_10546,N_10406,N_10351);
nand U10547 (N_10547,N_10464,N_10459);
or U10548 (N_10548,N_10421,N_10465);
and U10549 (N_10549,N_10499,N_10482);
xnor U10550 (N_10550,N_10359,N_10462);
xnor U10551 (N_10551,N_10367,N_10369);
or U10552 (N_10552,N_10380,N_10379);
and U10553 (N_10553,N_10261,N_10448);
nor U10554 (N_10554,N_10401,N_10339);
xor U10555 (N_10555,N_10491,N_10252);
nor U10556 (N_10556,N_10280,N_10360);
or U10557 (N_10557,N_10256,N_10338);
and U10558 (N_10558,N_10362,N_10304);
nand U10559 (N_10559,N_10467,N_10441);
nand U10560 (N_10560,N_10336,N_10395);
xnor U10561 (N_10561,N_10412,N_10404);
or U10562 (N_10562,N_10476,N_10492);
and U10563 (N_10563,N_10469,N_10308);
xor U10564 (N_10564,N_10258,N_10436);
and U10565 (N_10565,N_10259,N_10278);
nand U10566 (N_10566,N_10294,N_10324);
and U10567 (N_10567,N_10282,N_10375);
nand U10568 (N_10568,N_10335,N_10313);
and U10569 (N_10569,N_10292,N_10478);
or U10570 (N_10570,N_10433,N_10293);
nand U10571 (N_10571,N_10445,N_10460);
nor U10572 (N_10572,N_10322,N_10430);
and U10573 (N_10573,N_10485,N_10391);
nor U10574 (N_10574,N_10363,N_10451);
nand U10575 (N_10575,N_10495,N_10389);
nand U10576 (N_10576,N_10416,N_10487);
or U10577 (N_10577,N_10250,N_10477);
and U10578 (N_10578,N_10393,N_10382);
xnor U10579 (N_10579,N_10268,N_10301);
xor U10580 (N_10580,N_10355,N_10314);
nand U10581 (N_10581,N_10481,N_10453);
xor U10582 (N_10582,N_10414,N_10471);
nand U10583 (N_10583,N_10273,N_10319);
and U10584 (N_10584,N_10341,N_10475);
nand U10585 (N_10585,N_10486,N_10424);
nand U10586 (N_10586,N_10331,N_10326);
nor U10587 (N_10587,N_10327,N_10394);
nand U10588 (N_10588,N_10265,N_10372);
and U10589 (N_10589,N_10333,N_10408);
or U10590 (N_10590,N_10276,N_10444);
nand U10591 (N_10591,N_10457,N_10254);
nand U10592 (N_10592,N_10493,N_10480);
nor U10593 (N_10593,N_10302,N_10271);
or U10594 (N_10594,N_10410,N_10274);
nand U10595 (N_10595,N_10270,N_10496);
xor U10596 (N_10596,N_10361,N_10264);
and U10597 (N_10597,N_10323,N_10400);
nand U10598 (N_10598,N_10442,N_10272);
nand U10599 (N_10599,N_10348,N_10396);
nand U10600 (N_10600,N_10483,N_10285);
and U10601 (N_10601,N_10325,N_10286);
nor U10602 (N_10602,N_10358,N_10439);
or U10603 (N_10603,N_10352,N_10364);
or U10604 (N_10604,N_10337,N_10316);
or U10605 (N_10605,N_10253,N_10463);
and U10606 (N_10606,N_10484,N_10411);
nor U10607 (N_10607,N_10383,N_10283);
nor U10608 (N_10608,N_10415,N_10345);
nor U10609 (N_10609,N_10267,N_10284);
nand U10610 (N_10610,N_10473,N_10418);
and U10611 (N_10611,N_10376,N_10281);
or U10612 (N_10612,N_10297,N_10354);
nor U10613 (N_10613,N_10494,N_10329);
or U10614 (N_10614,N_10357,N_10349);
nand U10615 (N_10615,N_10417,N_10353);
nand U10616 (N_10616,N_10269,N_10287);
or U10617 (N_10617,N_10446,N_10366);
xnor U10618 (N_10618,N_10390,N_10342);
and U10619 (N_10619,N_10432,N_10455);
xor U10620 (N_10620,N_10255,N_10443);
and U10621 (N_10621,N_10420,N_10413);
nor U10622 (N_10622,N_10497,N_10251);
xor U10623 (N_10623,N_10263,N_10387);
and U10624 (N_10624,N_10340,N_10423);
xnor U10625 (N_10625,N_10261,N_10449);
or U10626 (N_10626,N_10425,N_10434);
nor U10627 (N_10627,N_10414,N_10439);
and U10628 (N_10628,N_10361,N_10458);
and U10629 (N_10629,N_10351,N_10362);
and U10630 (N_10630,N_10435,N_10411);
nand U10631 (N_10631,N_10282,N_10437);
and U10632 (N_10632,N_10272,N_10449);
and U10633 (N_10633,N_10455,N_10381);
xor U10634 (N_10634,N_10488,N_10401);
and U10635 (N_10635,N_10338,N_10499);
xnor U10636 (N_10636,N_10496,N_10356);
or U10637 (N_10637,N_10382,N_10298);
xor U10638 (N_10638,N_10402,N_10473);
nand U10639 (N_10639,N_10278,N_10495);
xor U10640 (N_10640,N_10489,N_10354);
and U10641 (N_10641,N_10364,N_10466);
nand U10642 (N_10642,N_10499,N_10350);
nand U10643 (N_10643,N_10348,N_10378);
or U10644 (N_10644,N_10483,N_10451);
nor U10645 (N_10645,N_10345,N_10306);
and U10646 (N_10646,N_10381,N_10456);
xor U10647 (N_10647,N_10488,N_10287);
and U10648 (N_10648,N_10334,N_10439);
and U10649 (N_10649,N_10478,N_10332);
xnor U10650 (N_10650,N_10499,N_10374);
xnor U10651 (N_10651,N_10333,N_10354);
or U10652 (N_10652,N_10432,N_10440);
nand U10653 (N_10653,N_10336,N_10475);
nor U10654 (N_10654,N_10472,N_10441);
nand U10655 (N_10655,N_10481,N_10383);
or U10656 (N_10656,N_10291,N_10337);
xor U10657 (N_10657,N_10400,N_10301);
or U10658 (N_10658,N_10456,N_10436);
or U10659 (N_10659,N_10460,N_10287);
nand U10660 (N_10660,N_10262,N_10253);
xnor U10661 (N_10661,N_10444,N_10294);
nand U10662 (N_10662,N_10352,N_10446);
and U10663 (N_10663,N_10420,N_10333);
xnor U10664 (N_10664,N_10499,N_10298);
or U10665 (N_10665,N_10494,N_10437);
xor U10666 (N_10666,N_10312,N_10381);
xnor U10667 (N_10667,N_10388,N_10343);
nand U10668 (N_10668,N_10349,N_10447);
nor U10669 (N_10669,N_10300,N_10496);
or U10670 (N_10670,N_10408,N_10374);
xor U10671 (N_10671,N_10499,N_10489);
nor U10672 (N_10672,N_10347,N_10399);
xnor U10673 (N_10673,N_10303,N_10475);
nand U10674 (N_10674,N_10258,N_10289);
or U10675 (N_10675,N_10288,N_10397);
and U10676 (N_10676,N_10259,N_10489);
and U10677 (N_10677,N_10419,N_10307);
xor U10678 (N_10678,N_10445,N_10344);
or U10679 (N_10679,N_10367,N_10325);
or U10680 (N_10680,N_10313,N_10265);
or U10681 (N_10681,N_10496,N_10322);
or U10682 (N_10682,N_10440,N_10363);
nor U10683 (N_10683,N_10471,N_10386);
or U10684 (N_10684,N_10309,N_10353);
xnor U10685 (N_10685,N_10448,N_10339);
nor U10686 (N_10686,N_10338,N_10468);
nand U10687 (N_10687,N_10274,N_10451);
xor U10688 (N_10688,N_10477,N_10258);
xnor U10689 (N_10689,N_10453,N_10257);
nor U10690 (N_10690,N_10299,N_10288);
and U10691 (N_10691,N_10364,N_10323);
or U10692 (N_10692,N_10482,N_10328);
xor U10693 (N_10693,N_10475,N_10356);
or U10694 (N_10694,N_10329,N_10300);
nand U10695 (N_10695,N_10287,N_10274);
and U10696 (N_10696,N_10447,N_10380);
xnor U10697 (N_10697,N_10435,N_10497);
xnor U10698 (N_10698,N_10263,N_10357);
or U10699 (N_10699,N_10345,N_10389);
or U10700 (N_10700,N_10390,N_10495);
nor U10701 (N_10701,N_10456,N_10260);
nor U10702 (N_10702,N_10448,N_10421);
and U10703 (N_10703,N_10405,N_10320);
nor U10704 (N_10704,N_10403,N_10350);
or U10705 (N_10705,N_10429,N_10414);
xor U10706 (N_10706,N_10268,N_10278);
nor U10707 (N_10707,N_10449,N_10376);
or U10708 (N_10708,N_10394,N_10348);
and U10709 (N_10709,N_10277,N_10445);
and U10710 (N_10710,N_10292,N_10498);
and U10711 (N_10711,N_10267,N_10277);
and U10712 (N_10712,N_10434,N_10415);
nand U10713 (N_10713,N_10481,N_10325);
nor U10714 (N_10714,N_10357,N_10432);
nor U10715 (N_10715,N_10400,N_10330);
xnor U10716 (N_10716,N_10488,N_10458);
and U10717 (N_10717,N_10359,N_10302);
nand U10718 (N_10718,N_10397,N_10455);
nand U10719 (N_10719,N_10359,N_10380);
nor U10720 (N_10720,N_10416,N_10301);
and U10721 (N_10721,N_10408,N_10460);
or U10722 (N_10722,N_10460,N_10315);
and U10723 (N_10723,N_10423,N_10474);
and U10724 (N_10724,N_10497,N_10493);
and U10725 (N_10725,N_10496,N_10308);
nor U10726 (N_10726,N_10398,N_10463);
nor U10727 (N_10727,N_10291,N_10301);
or U10728 (N_10728,N_10424,N_10440);
or U10729 (N_10729,N_10291,N_10310);
nand U10730 (N_10730,N_10252,N_10448);
or U10731 (N_10731,N_10415,N_10382);
or U10732 (N_10732,N_10365,N_10356);
or U10733 (N_10733,N_10446,N_10472);
xnor U10734 (N_10734,N_10350,N_10345);
and U10735 (N_10735,N_10440,N_10262);
nand U10736 (N_10736,N_10498,N_10275);
nand U10737 (N_10737,N_10250,N_10251);
and U10738 (N_10738,N_10251,N_10441);
nand U10739 (N_10739,N_10467,N_10290);
nand U10740 (N_10740,N_10480,N_10426);
or U10741 (N_10741,N_10390,N_10432);
and U10742 (N_10742,N_10440,N_10386);
xnor U10743 (N_10743,N_10293,N_10398);
xnor U10744 (N_10744,N_10383,N_10387);
or U10745 (N_10745,N_10309,N_10255);
or U10746 (N_10746,N_10297,N_10258);
or U10747 (N_10747,N_10487,N_10387);
nand U10748 (N_10748,N_10350,N_10312);
and U10749 (N_10749,N_10463,N_10357);
nand U10750 (N_10750,N_10504,N_10697);
or U10751 (N_10751,N_10728,N_10628);
or U10752 (N_10752,N_10602,N_10539);
nor U10753 (N_10753,N_10501,N_10599);
xnor U10754 (N_10754,N_10631,N_10634);
or U10755 (N_10755,N_10689,N_10642);
nor U10756 (N_10756,N_10654,N_10584);
nand U10757 (N_10757,N_10702,N_10572);
nand U10758 (N_10758,N_10625,N_10554);
xnor U10759 (N_10759,N_10540,N_10607);
xor U10760 (N_10760,N_10712,N_10664);
or U10761 (N_10761,N_10617,N_10551);
and U10762 (N_10762,N_10666,N_10698);
nor U10763 (N_10763,N_10612,N_10546);
or U10764 (N_10764,N_10542,N_10692);
xor U10765 (N_10765,N_10544,N_10734);
xor U10766 (N_10766,N_10635,N_10578);
or U10767 (N_10767,N_10737,N_10574);
xor U10768 (N_10768,N_10717,N_10512);
xnor U10769 (N_10769,N_10685,N_10577);
xnor U10770 (N_10770,N_10722,N_10726);
nor U10771 (N_10771,N_10743,N_10543);
or U10772 (N_10772,N_10626,N_10509);
xnor U10773 (N_10773,N_10600,N_10529);
nor U10774 (N_10774,N_10526,N_10581);
xnor U10775 (N_10775,N_10733,N_10708);
or U10776 (N_10776,N_10649,N_10710);
or U10777 (N_10777,N_10629,N_10606);
xor U10778 (N_10778,N_10669,N_10648);
nor U10779 (N_10779,N_10541,N_10621);
or U10780 (N_10780,N_10729,N_10559);
and U10781 (N_10781,N_10638,N_10618);
xor U10782 (N_10782,N_10736,N_10695);
or U10783 (N_10783,N_10675,N_10706);
or U10784 (N_10784,N_10604,N_10705);
nand U10785 (N_10785,N_10627,N_10598);
nor U10786 (N_10786,N_10550,N_10522);
nor U10787 (N_10787,N_10592,N_10566);
nor U10788 (N_10788,N_10715,N_10514);
nor U10789 (N_10789,N_10713,N_10594);
or U10790 (N_10790,N_10677,N_10730);
and U10791 (N_10791,N_10748,N_10718);
xor U10792 (N_10792,N_10740,N_10601);
nand U10793 (N_10793,N_10747,N_10580);
xor U10794 (N_10794,N_10533,N_10537);
nor U10795 (N_10795,N_10739,N_10508);
xnor U10796 (N_10796,N_10548,N_10534);
or U10797 (N_10797,N_10745,N_10667);
nor U10798 (N_10798,N_10549,N_10741);
or U10799 (N_10799,N_10615,N_10707);
and U10800 (N_10800,N_10573,N_10700);
and U10801 (N_10801,N_10703,N_10721);
or U10802 (N_10802,N_10585,N_10555);
and U10803 (N_10803,N_10630,N_10590);
nor U10804 (N_10804,N_10576,N_10672);
xor U10805 (N_10805,N_10693,N_10701);
or U10806 (N_10806,N_10620,N_10738);
nor U10807 (N_10807,N_10662,N_10680);
xnor U10808 (N_10808,N_10524,N_10595);
and U10809 (N_10809,N_10742,N_10608);
and U10810 (N_10810,N_10647,N_10510);
xnor U10811 (N_10811,N_10731,N_10732);
xor U10812 (N_10812,N_10659,N_10694);
nand U10813 (N_10813,N_10605,N_10530);
nand U10814 (N_10814,N_10587,N_10516);
or U10815 (N_10815,N_10583,N_10586);
nand U10816 (N_10816,N_10614,N_10749);
nor U10817 (N_10817,N_10547,N_10643);
nand U10818 (N_10818,N_10517,N_10513);
or U10819 (N_10819,N_10560,N_10663);
nor U10820 (N_10820,N_10670,N_10593);
nor U10821 (N_10821,N_10678,N_10660);
nand U10822 (N_10822,N_10727,N_10565);
or U10823 (N_10823,N_10639,N_10535);
nor U10824 (N_10824,N_10686,N_10563);
nand U10825 (N_10825,N_10538,N_10506);
xnor U10826 (N_10826,N_10556,N_10633);
or U10827 (N_10827,N_10714,N_10724);
or U10828 (N_10828,N_10582,N_10519);
and U10829 (N_10829,N_10716,N_10658);
or U10830 (N_10830,N_10553,N_10589);
xnor U10831 (N_10831,N_10661,N_10562);
nand U10832 (N_10832,N_10699,N_10637);
or U10833 (N_10833,N_10668,N_10507);
nor U10834 (N_10834,N_10719,N_10656);
nand U10835 (N_10835,N_10561,N_10611);
or U10836 (N_10836,N_10684,N_10655);
or U10837 (N_10837,N_10521,N_10644);
xnor U10838 (N_10838,N_10735,N_10588);
and U10839 (N_10839,N_10690,N_10709);
nor U10840 (N_10840,N_10579,N_10632);
and U10841 (N_10841,N_10500,N_10591);
and U10842 (N_10842,N_10568,N_10681);
nor U10843 (N_10843,N_10746,N_10570);
and U10844 (N_10844,N_10723,N_10528);
nand U10845 (N_10845,N_10711,N_10624);
nand U10846 (N_10846,N_10503,N_10515);
or U10847 (N_10847,N_10518,N_10502);
xor U10848 (N_10848,N_10575,N_10683);
nand U10849 (N_10849,N_10596,N_10523);
or U10850 (N_10850,N_10652,N_10720);
and U10851 (N_10851,N_10671,N_10623);
or U10852 (N_10852,N_10650,N_10532);
xnor U10853 (N_10853,N_10619,N_10511);
or U10854 (N_10854,N_10609,N_10674);
nor U10855 (N_10855,N_10622,N_10653);
and U10856 (N_10856,N_10545,N_10744);
nand U10857 (N_10857,N_10641,N_10657);
xnor U10858 (N_10858,N_10691,N_10531);
and U10859 (N_10859,N_10687,N_10571);
or U10860 (N_10860,N_10688,N_10536);
xor U10861 (N_10861,N_10505,N_10567);
xor U10862 (N_10862,N_10676,N_10564);
xor U10863 (N_10863,N_10558,N_10597);
or U10864 (N_10864,N_10640,N_10557);
nor U10865 (N_10865,N_10616,N_10520);
and U10866 (N_10866,N_10696,N_10613);
nand U10867 (N_10867,N_10651,N_10569);
and U10868 (N_10868,N_10725,N_10525);
and U10869 (N_10869,N_10603,N_10704);
or U10870 (N_10870,N_10610,N_10552);
xnor U10871 (N_10871,N_10679,N_10636);
and U10872 (N_10872,N_10527,N_10673);
nor U10873 (N_10873,N_10665,N_10645);
xor U10874 (N_10874,N_10682,N_10646);
nand U10875 (N_10875,N_10617,N_10586);
nand U10876 (N_10876,N_10732,N_10717);
xor U10877 (N_10877,N_10741,N_10714);
nor U10878 (N_10878,N_10556,N_10667);
and U10879 (N_10879,N_10556,N_10612);
nor U10880 (N_10880,N_10620,N_10517);
or U10881 (N_10881,N_10721,N_10511);
and U10882 (N_10882,N_10635,N_10630);
nor U10883 (N_10883,N_10709,N_10576);
and U10884 (N_10884,N_10535,N_10548);
nand U10885 (N_10885,N_10625,N_10645);
nand U10886 (N_10886,N_10528,N_10692);
or U10887 (N_10887,N_10548,N_10609);
nand U10888 (N_10888,N_10715,N_10659);
or U10889 (N_10889,N_10723,N_10735);
nor U10890 (N_10890,N_10702,N_10531);
nor U10891 (N_10891,N_10503,N_10552);
and U10892 (N_10892,N_10701,N_10691);
nor U10893 (N_10893,N_10515,N_10723);
or U10894 (N_10894,N_10650,N_10641);
or U10895 (N_10895,N_10736,N_10653);
and U10896 (N_10896,N_10717,N_10510);
or U10897 (N_10897,N_10583,N_10596);
xor U10898 (N_10898,N_10671,N_10515);
or U10899 (N_10899,N_10631,N_10690);
or U10900 (N_10900,N_10641,N_10597);
xor U10901 (N_10901,N_10684,N_10660);
nand U10902 (N_10902,N_10626,N_10573);
or U10903 (N_10903,N_10668,N_10678);
or U10904 (N_10904,N_10613,N_10560);
or U10905 (N_10905,N_10622,N_10566);
nor U10906 (N_10906,N_10634,N_10655);
and U10907 (N_10907,N_10731,N_10532);
nor U10908 (N_10908,N_10633,N_10581);
and U10909 (N_10909,N_10586,N_10710);
xnor U10910 (N_10910,N_10586,N_10562);
nor U10911 (N_10911,N_10743,N_10701);
xor U10912 (N_10912,N_10602,N_10720);
xor U10913 (N_10913,N_10744,N_10723);
nor U10914 (N_10914,N_10707,N_10703);
nor U10915 (N_10915,N_10518,N_10739);
and U10916 (N_10916,N_10705,N_10718);
nor U10917 (N_10917,N_10611,N_10656);
nor U10918 (N_10918,N_10593,N_10546);
xor U10919 (N_10919,N_10549,N_10684);
nor U10920 (N_10920,N_10693,N_10593);
xnor U10921 (N_10921,N_10533,N_10582);
xor U10922 (N_10922,N_10526,N_10559);
nor U10923 (N_10923,N_10705,N_10628);
or U10924 (N_10924,N_10505,N_10609);
nor U10925 (N_10925,N_10532,N_10571);
xor U10926 (N_10926,N_10521,N_10571);
or U10927 (N_10927,N_10551,N_10595);
xnor U10928 (N_10928,N_10610,N_10710);
nand U10929 (N_10929,N_10686,N_10706);
and U10930 (N_10930,N_10565,N_10657);
nand U10931 (N_10931,N_10681,N_10558);
nand U10932 (N_10932,N_10721,N_10672);
nor U10933 (N_10933,N_10612,N_10620);
and U10934 (N_10934,N_10686,N_10722);
nor U10935 (N_10935,N_10702,N_10541);
nand U10936 (N_10936,N_10648,N_10710);
nand U10937 (N_10937,N_10561,N_10709);
or U10938 (N_10938,N_10697,N_10612);
nand U10939 (N_10939,N_10673,N_10587);
xor U10940 (N_10940,N_10709,N_10611);
nor U10941 (N_10941,N_10721,N_10586);
and U10942 (N_10942,N_10735,N_10620);
nor U10943 (N_10943,N_10731,N_10706);
or U10944 (N_10944,N_10662,N_10539);
or U10945 (N_10945,N_10507,N_10666);
nand U10946 (N_10946,N_10508,N_10534);
or U10947 (N_10947,N_10522,N_10727);
nand U10948 (N_10948,N_10633,N_10666);
or U10949 (N_10949,N_10678,N_10587);
or U10950 (N_10950,N_10673,N_10632);
nand U10951 (N_10951,N_10559,N_10642);
or U10952 (N_10952,N_10590,N_10639);
and U10953 (N_10953,N_10533,N_10612);
xor U10954 (N_10954,N_10513,N_10610);
nand U10955 (N_10955,N_10740,N_10575);
or U10956 (N_10956,N_10653,N_10724);
and U10957 (N_10957,N_10531,N_10646);
and U10958 (N_10958,N_10745,N_10580);
xnor U10959 (N_10959,N_10586,N_10559);
xor U10960 (N_10960,N_10609,N_10561);
xor U10961 (N_10961,N_10734,N_10549);
nor U10962 (N_10962,N_10632,N_10669);
nor U10963 (N_10963,N_10515,N_10726);
xor U10964 (N_10964,N_10619,N_10691);
nand U10965 (N_10965,N_10545,N_10644);
xor U10966 (N_10966,N_10554,N_10748);
and U10967 (N_10967,N_10606,N_10664);
xor U10968 (N_10968,N_10570,N_10644);
xnor U10969 (N_10969,N_10688,N_10593);
xor U10970 (N_10970,N_10527,N_10604);
and U10971 (N_10971,N_10737,N_10638);
nand U10972 (N_10972,N_10669,N_10549);
or U10973 (N_10973,N_10670,N_10548);
or U10974 (N_10974,N_10662,N_10623);
and U10975 (N_10975,N_10664,N_10513);
and U10976 (N_10976,N_10576,N_10511);
nor U10977 (N_10977,N_10615,N_10739);
and U10978 (N_10978,N_10639,N_10602);
xnor U10979 (N_10979,N_10537,N_10712);
xnor U10980 (N_10980,N_10620,N_10596);
xor U10981 (N_10981,N_10630,N_10656);
xnor U10982 (N_10982,N_10564,N_10608);
xnor U10983 (N_10983,N_10717,N_10589);
or U10984 (N_10984,N_10503,N_10660);
xnor U10985 (N_10985,N_10594,N_10602);
or U10986 (N_10986,N_10516,N_10517);
xnor U10987 (N_10987,N_10582,N_10604);
and U10988 (N_10988,N_10614,N_10696);
and U10989 (N_10989,N_10666,N_10598);
nor U10990 (N_10990,N_10550,N_10638);
nand U10991 (N_10991,N_10664,N_10624);
nor U10992 (N_10992,N_10631,N_10680);
or U10993 (N_10993,N_10736,N_10518);
nand U10994 (N_10994,N_10608,N_10646);
xor U10995 (N_10995,N_10690,N_10648);
nand U10996 (N_10996,N_10508,N_10695);
nand U10997 (N_10997,N_10696,N_10718);
or U10998 (N_10998,N_10638,N_10747);
or U10999 (N_10999,N_10519,N_10532);
or U11000 (N_11000,N_10942,N_10946);
and U11001 (N_11001,N_10768,N_10827);
or U11002 (N_11002,N_10852,N_10780);
and U11003 (N_11003,N_10868,N_10947);
and U11004 (N_11004,N_10990,N_10941);
nor U11005 (N_11005,N_10895,N_10904);
and U11006 (N_11006,N_10937,N_10853);
or U11007 (N_11007,N_10881,N_10988);
nor U11008 (N_11008,N_10960,N_10916);
and U11009 (N_11009,N_10884,N_10846);
or U11010 (N_11010,N_10981,N_10834);
or U11011 (N_11011,N_10831,N_10836);
xor U11012 (N_11012,N_10973,N_10896);
or U11013 (N_11013,N_10980,N_10806);
xnor U11014 (N_11014,N_10793,N_10871);
xnor U11015 (N_11015,N_10890,N_10903);
nor U11016 (N_11016,N_10933,N_10765);
or U11017 (N_11017,N_10804,N_10756);
nor U11018 (N_11018,N_10979,N_10835);
nor U11019 (N_11019,N_10959,N_10877);
or U11020 (N_11020,N_10923,N_10940);
and U11021 (N_11021,N_10864,N_10921);
xor U11022 (N_11022,N_10821,N_10826);
or U11023 (N_11023,N_10924,N_10810);
nor U11024 (N_11024,N_10757,N_10931);
xnor U11025 (N_11025,N_10816,N_10987);
nand U11026 (N_11026,N_10887,N_10996);
or U11027 (N_11027,N_10982,N_10754);
nor U11028 (N_11028,N_10859,N_10976);
or U11029 (N_11029,N_10812,N_10944);
nand U11030 (N_11030,N_10967,N_10808);
nor U11031 (N_11031,N_10770,N_10983);
xnor U11032 (N_11032,N_10753,N_10932);
or U11033 (N_11033,N_10855,N_10811);
xor U11034 (N_11034,N_10898,N_10902);
xnor U11035 (N_11035,N_10954,N_10917);
nor U11036 (N_11036,N_10766,N_10784);
nor U11037 (N_11037,N_10888,N_10750);
xor U11038 (N_11038,N_10799,N_10909);
and U11039 (N_11039,N_10789,N_10935);
nor U11040 (N_11040,N_10761,N_10854);
nand U11041 (N_11041,N_10752,N_10999);
and U11042 (N_11042,N_10841,N_10934);
xnor U11043 (N_11043,N_10781,N_10797);
and U11044 (N_11044,N_10995,N_10880);
nand U11045 (N_11045,N_10928,N_10778);
or U11046 (N_11046,N_10885,N_10872);
nor U11047 (N_11047,N_10971,N_10782);
xnor U11048 (N_11048,N_10956,N_10849);
or U11049 (N_11049,N_10882,N_10813);
xor U11050 (N_11050,N_10913,N_10867);
or U11051 (N_11051,N_10860,N_10794);
xor U11052 (N_11052,N_10767,N_10838);
xor U11053 (N_11053,N_10843,N_10978);
nor U11054 (N_11054,N_10861,N_10958);
or U11055 (N_11055,N_10769,N_10939);
xnor U11056 (N_11056,N_10815,N_10985);
or U11057 (N_11057,N_10863,N_10875);
or U11058 (N_11058,N_10791,N_10788);
and U11059 (N_11059,N_10907,N_10927);
or U11060 (N_11060,N_10828,N_10972);
and U11061 (N_11061,N_10930,N_10787);
nand U11062 (N_11062,N_10856,N_10886);
nor U11063 (N_11063,N_10974,N_10866);
nand U11064 (N_11064,N_10825,N_10848);
or U11065 (N_11065,N_10989,N_10986);
or U11066 (N_11066,N_10805,N_10845);
or U11067 (N_11067,N_10879,N_10893);
nand U11068 (N_11068,N_10858,N_10950);
xor U11069 (N_11069,N_10851,N_10953);
nor U11070 (N_11070,N_10798,N_10912);
nor U11071 (N_11071,N_10817,N_10964);
xnor U11072 (N_11072,N_10922,N_10993);
and U11073 (N_11073,N_10992,N_10862);
nand U11074 (N_11074,N_10844,N_10897);
xnor U11075 (N_11075,N_10955,N_10809);
or U11076 (N_11076,N_10832,N_10785);
xor U11077 (N_11077,N_10759,N_10820);
xor U11078 (N_11078,N_10777,N_10926);
and U11079 (N_11079,N_10760,N_10751);
nand U11080 (N_11080,N_10968,N_10965);
or U11081 (N_11081,N_10833,N_10929);
and U11082 (N_11082,N_10943,N_10900);
xnor U11083 (N_11083,N_10911,N_10906);
or U11084 (N_11084,N_10850,N_10915);
or U11085 (N_11085,N_10957,N_10969);
and U11086 (N_11086,N_10814,N_10774);
or U11087 (N_11087,N_10918,N_10842);
nor U11088 (N_11088,N_10763,N_10899);
nor U11089 (N_11089,N_10962,N_10819);
nor U11090 (N_11090,N_10966,N_10920);
and U11091 (N_11091,N_10889,N_10914);
nand U11092 (N_11092,N_10783,N_10792);
and U11093 (N_11093,N_10870,N_10865);
and U11094 (N_11094,N_10840,N_10824);
nand U11095 (N_11095,N_10764,N_10755);
xnor U11096 (N_11096,N_10894,N_10790);
and U11097 (N_11097,N_10977,N_10818);
and U11098 (N_11098,N_10803,N_10901);
xor U11099 (N_11099,N_10876,N_10796);
or U11100 (N_11100,N_10823,N_10994);
xor U11101 (N_11101,N_10771,N_10847);
xor U11102 (N_11102,N_10873,N_10800);
nor U11103 (N_11103,N_10822,N_10998);
or U11104 (N_11104,N_10891,N_10807);
nor U11105 (N_11105,N_10991,N_10963);
nand U11106 (N_11106,N_10801,N_10795);
nand U11107 (N_11107,N_10949,N_10773);
nand U11108 (N_11108,N_10908,N_10758);
and U11109 (N_11109,N_10874,N_10910);
nand U11110 (N_11110,N_10772,N_10883);
nor U11111 (N_11111,N_10776,N_10857);
and U11112 (N_11112,N_10892,N_10829);
xor U11113 (N_11113,N_10997,N_10802);
nor U11114 (N_11114,N_10779,N_10925);
xor U11115 (N_11115,N_10948,N_10919);
nor U11116 (N_11116,N_10830,N_10786);
xnor U11117 (N_11117,N_10951,N_10975);
and U11118 (N_11118,N_10952,N_10878);
nor U11119 (N_11119,N_10837,N_10938);
nor U11120 (N_11120,N_10945,N_10762);
nand U11121 (N_11121,N_10869,N_10961);
nand U11122 (N_11122,N_10839,N_10984);
nand U11123 (N_11123,N_10936,N_10905);
and U11124 (N_11124,N_10970,N_10775);
or U11125 (N_11125,N_10885,N_10980);
or U11126 (N_11126,N_10799,N_10763);
xor U11127 (N_11127,N_10773,N_10964);
nand U11128 (N_11128,N_10910,N_10881);
nor U11129 (N_11129,N_10883,N_10868);
nand U11130 (N_11130,N_10792,N_10891);
nor U11131 (N_11131,N_10800,N_10850);
and U11132 (N_11132,N_10812,N_10829);
nor U11133 (N_11133,N_10980,N_10825);
and U11134 (N_11134,N_10918,N_10929);
xor U11135 (N_11135,N_10886,N_10774);
and U11136 (N_11136,N_10888,N_10936);
nand U11137 (N_11137,N_10753,N_10965);
nor U11138 (N_11138,N_10819,N_10888);
nand U11139 (N_11139,N_10961,N_10807);
or U11140 (N_11140,N_10990,N_10800);
nand U11141 (N_11141,N_10882,N_10993);
or U11142 (N_11142,N_10935,N_10973);
nand U11143 (N_11143,N_10796,N_10916);
or U11144 (N_11144,N_10823,N_10877);
and U11145 (N_11145,N_10980,N_10762);
or U11146 (N_11146,N_10811,N_10875);
nand U11147 (N_11147,N_10762,N_10960);
nor U11148 (N_11148,N_10769,N_10998);
nor U11149 (N_11149,N_10877,N_10866);
or U11150 (N_11150,N_10861,N_10977);
xnor U11151 (N_11151,N_10782,N_10816);
or U11152 (N_11152,N_10772,N_10964);
nor U11153 (N_11153,N_10781,N_10846);
or U11154 (N_11154,N_10919,N_10841);
nand U11155 (N_11155,N_10882,N_10857);
nor U11156 (N_11156,N_10840,N_10936);
xor U11157 (N_11157,N_10940,N_10786);
nor U11158 (N_11158,N_10824,N_10750);
nor U11159 (N_11159,N_10912,N_10868);
nand U11160 (N_11160,N_10855,N_10899);
and U11161 (N_11161,N_10851,N_10861);
and U11162 (N_11162,N_10943,N_10926);
or U11163 (N_11163,N_10774,N_10785);
or U11164 (N_11164,N_10932,N_10861);
or U11165 (N_11165,N_10767,N_10995);
nor U11166 (N_11166,N_10916,N_10785);
and U11167 (N_11167,N_10760,N_10985);
and U11168 (N_11168,N_10761,N_10928);
or U11169 (N_11169,N_10775,N_10824);
and U11170 (N_11170,N_10809,N_10950);
xnor U11171 (N_11171,N_10981,N_10773);
xnor U11172 (N_11172,N_10770,N_10939);
and U11173 (N_11173,N_10814,N_10776);
nand U11174 (N_11174,N_10835,N_10977);
or U11175 (N_11175,N_10831,N_10923);
or U11176 (N_11176,N_10990,N_10950);
nand U11177 (N_11177,N_10993,N_10802);
nor U11178 (N_11178,N_10834,N_10835);
xor U11179 (N_11179,N_10783,N_10788);
or U11180 (N_11180,N_10906,N_10756);
nor U11181 (N_11181,N_10787,N_10896);
and U11182 (N_11182,N_10942,N_10787);
xnor U11183 (N_11183,N_10990,N_10852);
or U11184 (N_11184,N_10815,N_10897);
or U11185 (N_11185,N_10796,N_10944);
or U11186 (N_11186,N_10955,N_10784);
nand U11187 (N_11187,N_10920,N_10814);
or U11188 (N_11188,N_10817,N_10871);
and U11189 (N_11189,N_10823,N_10872);
or U11190 (N_11190,N_10755,N_10908);
xor U11191 (N_11191,N_10761,N_10877);
nand U11192 (N_11192,N_10989,N_10809);
and U11193 (N_11193,N_10760,N_10990);
or U11194 (N_11194,N_10933,N_10923);
nand U11195 (N_11195,N_10906,N_10904);
and U11196 (N_11196,N_10789,N_10940);
xor U11197 (N_11197,N_10766,N_10951);
nor U11198 (N_11198,N_10955,N_10993);
nand U11199 (N_11199,N_10850,N_10950);
and U11200 (N_11200,N_10898,N_10807);
xnor U11201 (N_11201,N_10939,N_10857);
or U11202 (N_11202,N_10943,N_10859);
and U11203 (N_11203,N_10810,N_10769);
nand U11204 (N_11204,N_10998,N_10823);
xor U11205 (N_11205,N_10829,N_10925);
or U11206 (N_11206,N_10765,N_10795);
nor U11207 (N_11207,N_10750,N_10794);
xor U11208 (N_11208,N_10915,N_10874);
xnor U11209 (N_11209,N_10907,N_10842);
nand U11210 (N_11210,N_10779,N_10931);
or U11211 (N_11211,N_10888,N_10950);
or U11212 (N_11212,N_10984,N_10825);
xnor U11213 (N_11213,N_10764,N_10991);
nor U11214 (N_11214,N_10959,N_10937);
or U11215 (N_11215,N_10985,N_10887);
or U11216 (N_11216,N_10927,N_10974);
xnor U11217 (N_11217,N_10933,N_10914);
or U11218 (N_11218,N_10986,N_10870);
and U11219 (N_11219,N_10903,N_10796);
nor U11220 (N_11220,N_10960,N_10814);
and U11221 (N_11221,N_10788,N_10953);
nor U11222 (N_11222,N_10756,N_10947);
or U11223 (N_11223,N_10970,N_10972);
or U11224 (N_11224,N_10826,N_10916);
nand U11225 (N_11225,N_10910,N_10820);
or U11226 (N_11226,N_10893,N_10777);
nor U11227 (N_11227,N_10768,N_10835);
nand U11228 (N_11228,N_10972,N_10946);
nor U11229 (N_11229,N_10777,N_10829);
or U11230 (N_11230,N_10796,N_10931);
nand U11231 (N_11231,N_10915,N_10952);
xnor U11232 (N_11232,N_10840,N_10857);
nor U11233 (N_11233,N_10908,N_10991);
nand U11234 (N_11234,N_10753,N_10755);
or U11235 (N_11235,N_10835,N_10869);
xor U11236 (N_11236,N_10987,N_10819);
nor U11237 (N_11237,N_10759,N_10752);
or U11238 (N_11238,N_10901,N_10755);
xnor U11239 (N_11239,N_10976,N_10879);
or U11240 (N_11240,N_10808,N_10984);
and U11241 (N_11241,N_10995,N_10997);
or U11242 (N_11242,N_10941,N_10908);
or U11243 (N_11243,N_10961,N_10906);
nor U11244 (N_11244,N_10754,N_10854);
and U11245 (N_11245,N_10888,N_10893);
or U11246 (N_11246,N_10995,N_10898);
nor U11247 (N_11247,N_10965,N_10809);
or U11248 (N_11248,N_10758,N_10811);
and U11249 (N_11249,N_10918,N_10778);
or U11250 (N_11250,N_11167,N_11139);
and U11251 (N_11251,N_11000,N_11217);
and U11252 (N_11252,N_11148,N_11146);
nand U11253 (N_11253,N_11232,N_11051);
xor U11254 (N_11254,N_11174,N_11060);
and U11255 (N_11255,N_11027,N_11058);
xor U11256 (N_11256,N_11114,N_11048);
and U11257 (N_11257,N_11189,N_11046);
or U11258 (N_11258,N_11013,N_11176);
xnor U11259 (N_11259,N_11211,N_11108);
and U11260 (N_11260,N_11069,N_11201);
or U11261 (N_11261,N_11221,N_11079);
nor U11262 (N_11262,N_11083,N_11208);
xnor U11263 (N_11263,N_11132,N_11244);
nand U11264 (N_11264,N_11119,N_11166);
xor U11265 (N_11265,N_11142,N_11056);
xor U11266 (N_11266,N_11003,N_11161);
and U11267 (N_11267,N_11168,N_11126);
or U11268 (N_11268,N_11188,N_11033);
xor U11269 (N_11269,N_11065,N_11054);
or U11270 (N_11270,N_11059,N_11089);
and U11271 (N_11271,N_11042,N_11052);
or U11272 (N_11272,N_11047,N_11169);
nand U11273 (N_11273,N_11122,N_11175);
and U11274 (N_11274,N_11105,N_11164);
xor U11275 (N_11275,N_11072,N_11030);
xor U11276 (N_11276,N_11112,N_11036);
nand U11277 (N_11277,N_11149,N_11032);
xnor U11278 (N_11278,N_11055,N_11016);
nor U11279 (N_11279,N_11117,N_11045);
and U11280 (N_11280,N_11192,N_11124);
nand U11281 (N_11281,N_11015,N_11239);
and U11282 (N_11282,N_11064,N_11219);
xor U11283 (N_11283,N_11110,N_11062);
or U11284 (N_11284,N_11107,N_11007);
and U11285 (N_11285,N_11120,N_11031);
and U11286 (N_11286,N_11057,N_11134);
nor U11287 (N_11287,N_11247,N_11226);
and U11288 (N_11288,N_11180,N_11145);
or U11289 (N_11289,N_11076,N_11214);
nor U11290 (N_11290,N_11231,N_11215);
or U11291 (N_11291,N_11116,N_11075);
or U11292 (N_11292,N_11184,N_11002);
nor U11293 (N_11293,N_11179,N_11008);
xor U11294 (N_11294,N_11028,N_11049);
and U11295 (N_11295,N_11135,N_11094);
nand U11296 (N_11296,N_11044,N_11001);
or U11297 (N_11297,N_11121,N_11177);
and U11298 (N_11298,N_11216,N_11086);
or U11299 (N_11299,N_11014,N_11193);
nor U11300 (N_11300,N_11202,N_11106);
or U11301 (N_11301,N_11235,N_11037);
nand U11302 (N_11302,N_11066,N_11020);
and U11303 (N_11303,N_11093,N_11229);
nor U11304 (N_11304,N_11197,N_11204);
and U11305 (N_11305,N_11171,N_11095);
and U11306 (N_11306,N_11200,N_11141);
xnor U11307 (N_11307,N_11178,N_11207);
or U11308 (N_11308,N_11103,N_11158);
or U11309 (N_11309,N_11022,N_11102);
nor U11310 (N_11310,N_11063,N_11248);
or U11311 (N_11311,N_11067,N_11078);
nand U11312 (N_11312,N_11163,N_11115);
xor U11313 (N_11313,N_11034,N_11024);
or U11314 (N_11314,N_11236,N_11196);
nor U11315 (N_11315,N_11187,N_11153);
and U11316 (N_11316,N_11010,N_11109);
nor U11317 (N_11317,N_11021,N_11203);
or U11318 (N_11318,N_11156,N_11005);
xor U11319 (N_11319,N_11151,N_11233);
xnor U11320 (N_11320,N_11137,N_11157);
and U11321 (N_11321,N_11144,N_11138);
and U11322 (N_11322,N_11006,N_11209);
and U11323 (N_11323,N_11077,N_11129);
or U11324 (N_11324,N_11099,N_11084);
xor U11325 (N_11325,N_11080,N_11071);
or U11326 (N_11326,N_11050,N_11182);
or U11327 (N_11327,N_11041,N_11053);
nor U11328 (N_11328,N_11087,N_11023);
xor U11329 (N_11329,N_11123,N_11131);
nand U11330 (N_11330,N_11068,N_11186);
or U11331 (N_11331,N_11025,N_11029);
xor U11332 (N_11332,N_11194,N_11206);
nor U11333 (N_11333,N_11073,N_11183);
or U11334 (N_11334,N_11098,N_11043);
nand U11335 (N_11335,N_11088,N_11212);
and U11336 (N_11336,N_11074,N_11162);
xor U11337 (N_11337,N_11018,N_11118);
xnor U11338 (N_11338,N_11092,N_11213);
nand U11339 (N_11339,N_11227,N_11150);
and U11340 (N_11340,N_11155,N_11017);
nand U11341 (N_11341,N_11038,N_11011);
nand U11342 (N_11342,N_11154,N_11085);
and U11343 (N_11343,N_11185,N_11104);
xor U11344 (N_11344,N_11147,N_11181);
and U11345 (N_11345,N_11224,N_11097);
nand U11346 (N_11346,N_11160,N_11225);
nand U11347 (N_11347,N_11090,N_11143);
xnor U11348 (N_11348,N_11242,N_11195);
and U11349 (N_11349,N_11061,N_11082);
nor U11350 (N_11350,N_11228,N_11240);
and U11351 (N_11351,N_11249,N_11100);
nor U11352 (N_11352,N_11040,N_11190);
nand U11353 (N_11353,N_11127,N_11245);
or U11354 (N_11354,N_11230,N_11113);
xnor U11355 (N_11355,N_11136,N_11101);
nand U11356 (N_11356,N_11091,N_11125);
nor U11357 (N_11357,N_11004,N_11243);
xor U11358 (N_11358,N_11218,N_11246);
nand U11359 (N_11359,N_11170,N_11191);
nor U11360 (N_11360,N_11019,N_11241);
xor U11361 (N_11361,N_11070,N_11130);
nor U11362 (N_11362,N_11128,N_11159);
nand U11363 (N_11363,N_11234,N_11220);
and U11364 (N_11364,N_11165,N_11223);
and U11365 (N_11365,N_11140,N_11238);
or U11366 (N_11366,N_11173,N_11012);
nand U11367 (N_11367,N_11210,N_11009);
nand U11368 (N_11368,N_11133,N_11035);
xnor U11369 (N_11369,N_11237,N_11096);
xor U11370 (N_11370,N_11152,N_11199);
xnor U11371 (N_11371,N_11198,N_11111);
or U11372 (N_11372,N_11205,N_11026);
and U11373 (N_11373,N_11081,N_11222);
nand U11374 (N_11374,N_11172,N_11039);
nand U11375 (N_11375,N_11190,N_11158);
xor U11376 (N_11376,N_11148,N_11163);
nand U11377 (N_11377,N_11069,N_11098);
and U11378 (N_11378,N_11145,N_11129);
xnor U11379 (N_11379,N_11093,N_11014);
and U11380 (N_11380,N_11194,N_11107);
or U11381 (N_11381,N_11010,N_11009);
nand U11382 (N_11382,N_11078,N_11089);
and U11383 (N_11383,N_11038,N_11124);
nor U11384 (N_11384,N_11201,N_11131);
nor U11385 (N_11385,N_11141,N_11005);
nand U11386 (N_11386,N_11058,N_11100);
xor U11387 (N_11387,N_11237,N_11022);
nand U11388 (N_11388,N_11092,N_11240);
nand U11389 (N_11389,N_11001,N_11024);
nand U11390 (N_11390,N_11160,N_11039);
or U11391 (N_11391,N_11182,N_11088);
or U11392 (N_11392,N_11057,N_11016);
nor U11393 (N_11393,N_11076,N_11021);
nor U11394 (N_11394,N_11085,N_11163);
and U11395 (N_11395,N_11247,N_11095);
and U11396 (N_11396,N_11000,N_11221);
nor U11397 (N_11397,N_11160,N_11074);
nor U11398 (N_11398,N_11032,N_11137);
nor U11399 (N_11399,N_11120,N_11023);
nand U11400 (N_11400,N_11071,N_11135);
nand U11401 (N_11401,N_11032,N_11127);
nor U11402 (N_11402,N_11232,N_11175);
nor U11403 (N_11403,N_11226,N_11049);
nor U11404 (N_11404,N_11180,N_11132);
or U11405 (N_11405,N_11238,N_11212);
xnor U11406 (N_11406,N_11148,N_11239);
or U11407 (N_11407,N_11122,N_11041);
or U11408 (N_11408,N_11234,N_11227);
nor U11409 (N_11409,N_11078,N_11071);
nor U11410 (N_11410,N_11092,N_11218);
or U11411 (N_11411,N_11013,N_11181);
or U11412 (N_11412,N_11186,N_11076);
and U11413 (N_11413,N_11217,N_11078);
xor U11414 (N_11414,N_11052,N_11018);
nor U11415 (N_11415,N_11131,N_11152);
and U11416 (N_11416,N_11107,N_11146);
and U11417 (N_11417,N_11020,N_11098);
nand U11418 (N_11418,N_11113,N_11234);
nor U11419 (N_11419,N_11052,N_11032);
and U11420 (N_11420,N_11115,N_11087);
nand U11421 (N_11421,N_11100,N_11007);
and U11422 (N_11422,N_11017,N_11138);
xnor U11423 (N_11423,N_11076,N_11179);
nand U11424 (N_11424,N_11101,N_11147);
xnor U11425 (N_11425,N_11162,N_11032);
nor U11426 (N_11426,N_11219,N_11203);
nor U11427 (N_11427,N_11026,N_11032);
xor U11428 (N_11428,N_11104,N_11140);
xor U11429 (N_11429,N_11240,N_11149);
xnor U11430 (N_11430,N_11109,N_11097);
nand U11431 (N_11431,N_11197,N_11051);
nand U11432 (N_11432,N_11021,N_11039);
or U11433 (N_11433,N_11135,N_11055);
nor U11434 (N_11434,N_11112,N_11209);
or U11435 (N_11435,N_11094,N_11031);
nor U11436 (N_11436,N_11232,N_11186);
xnor U11437 (N_11437,N_11155,N_11047);
nand U11438 (N_11438,N_11028,N_11033);
and U11439 (N_11439,N_11047,N_11133);
nor U11440 (N_11440,N_11178,N_11008);
or U11441 (N_11441,N_11168,N_11099);
nor U11442 (N_11442,N_11056,N_11097);
and U11443 (N_11443,N_11128,N_11160);
nand U11444 (N_11444,N_11114,N_11113);
nor U11445 (N_11445,N_11056,N_11245);
and U11446 (N_11446,N_11065,N_11023);
and U11447 (N_11447,N_11046,N_11224);
or U11448 (N_11448,N_11091,N_11079);
nor U11449 (N_11449,N_11110,N_11109);
or U11450 (N_11450,N_11238,N_11153);
or U11451 (N_11451,N_11034,N_11196);
nor U11452 (N_11452,N_11126,N_11133);
nand U11453 (N_11453,N_11240,N_11106);
and U11454 (N_11454,N_11076,N_11174);
and U11455 (N_11455,N_11050,N_11078);
and U11456 (N_11456,N_11094,N_11211);
xnor U11457 (N_11457,N_11056,N_11062);
nor U11458 (N_11458,N_11179,N_11032);
or U11459 (N_11459,N_11063,N_11037);
xor U11460 (N_11460,N_11064,N_11216);
xnor U11461 (N_11461,N_11132,N_11025);
and U11462 (N_11462,N_11160,N_11211);
nand U11463 (N_11463,N_11215,N_11225);
or U11464 (N_11464,N_11038,N_11018);
or U11465 (N_11465,N_11221,N_11219);
nor U11466 (N_11466,N_11125,N_11012);
and U11467 (N_11467,N_11042,N_11015);
nor U11468 (N_11468,N_11095,N_11063);
or U11469 (N_11469,N_11171,N_11087);
nand U11470 (N_11470,N_11102,N_11062);
or U11471 (N_11471,N_11181,N_11227);
xor U11472 (N_11472,N_11213,N_11102);
or U11473 (N_11473,N_11146,N_11061);
xor U11474 (N_11474,N_11212,N_11103);
or U11475 (N_11475,N_11075,N_11036);
nand U11476 (N_11476,N_11078,N_11142);
or U11477 (N_11477,N_11027,N_11223);
and U11478 (N_11478,N_11039,N_11108);
nor U11479 (N_11479,N_11104,N_11009);
nand U11480 (N_11480,N_11200,N_11225);
nor U11481 (N_11481,N_11151,N_11091);
and U11482 (N_11482,N_11074,N_11034);
nand U11483 (N_11483,N_11039,N_11229);
or U11484 (N_11484,N_11115,N_11099);
nand U11485 (N_11485,N_11138,N_11241);
or U11486 (N_11486,N_11028,N_11048);
and U11487 (N_11487,N_11221,N_11120);
xnor U11488 (N_11488,N_11089,N_11093);
and U11489 (N_11489,N_11035,N_11159);
xnor U11490 (N_11490,N_11064,N_11108);
nor U11491 (N_11491,N_11181,N_11162);
nor U11492 (N_11492,N_11008,N_11074);
and U11493 (N_11493,N_11200,N_11042);
xor U11494 (N_11494,N_11167,N_11086);
and U11495 (N_11495,N_11159,N_11218);
nor U11496 (N_11496,N_11086,N_11144);
and U11497 (N_11497,N_11195,N_11058);
or U11498 (N_11498,N_11158,N_11159);
nand U11499 (N_11499,N_11042,N_11095);
nand U11500 (N_11500,N_11348,N_11275);
or U11501 (N_11501,N_11381,N_11466);
xor U11502 (N_11502,N_11333,N_11449);
nand U11503 (N_11503,N_11486,N_11416);
or U11504 (N_11504,N_11483,N_11346);
nand U11505 (N_11505,N_11308,N_11272);
xnor U11506 (N_11506,N_11292,N_11489);
and U11507 (N_11507,N_11335,N_11443);
nor U11508 (N_11508,N_11389,N_11339);
and U11509 (N_11509,N_11465,N_11378);
nor U11510 (N_11510,N_11278,N_11329);
xnor U11511 (N_11511,N_11277,N_11344);
or U11512 (N_11512,N_11418,N_11334);
nor U11513 (N_11513,N_11349,N_11434);
xor U11514 (N_11514,N_11487,N_11287);
nor U11515 (N_11515,N_11386,N_11340);
and U11516 (N_11516,N_11498,N_11251);
nor U11517 (N_11517,N_11447,N_11379);
nand U11518 (N_11518,N_11424,N_11408);
and U11519 (N_11519,N_11281,N_11490);
and U11520 (N_11520,N_11365,N_11468);
xnor U11521 (N_11521,N_11440,N_11317);
xor U11522 (N_11522,N_11455,N_11467);
or U11523 (N_11523,N_11315,N_11338);
or U11524 (N_11524,N_11250,N_11375);
nand U11525 (N_11525,N_11450,N_11398);
and U11526 (N_11526,N_11491,N_11351);
xnor U11527 (N_11527,N_11318,N_11458);
nand U11528 (N_11528,N_11353,N_11327);
or U11529 (N_11529,N_11256,N_11369);
nor U11530 (N_11530,N_11380,N_11401);
nor U11531 (N_11531,N_11331,N_11328);
and U11532 (N_11532,N_11284,N_11493);
or U11533 (N_11533,N_11395,N_11305);
xnor U11534 (N_11534,N_11463,N_11321);
xor U11535 (N_11535,N_11410,N_11392);
nand U11536 (N_11536,N_11480,N_11319);
nand U11537 (N_11537,N_11306,N_11293);
or U11538 (N_11538,N_11442,N_11454);
and U11539 (N_11539,N_11422,N_11453);
nand U11540 (N_11540,N_11355,N_11415);
and U11541 (N_11541,N_11430,N_11368);
nand U11542 (N_11542,N_11373,N_11457);
nor U11543 (N_11543,N_11377,N_11296);
xor U11544 (N_11544,N_11356,N_11370);
nor U11545 (N_11545,N_11324,N_11421);
nand U11546 (N_11546,N_11396,N_11297);
xor U11547 (N_11547,N_11484,N_11332);
xnor U11548 (N_11548,N_11499,N_11316);
nand U11549 (N_11549,N_11413,N_11258);
nand U11550 (N_11550,N_11361,N_11304);
and U11551 (N_11551,N_11270,N_11298);
xor U11552 (N_11552,N_11451,N_11268);
or U11553 (N_11553,N_11432,N_11291);
xnor U11554 (N_11554,N_11265,N_11269);
nand U11555 (N_11555,N_11439,N_11337);
and U11556 (N_11556,N_11260,N_11302);
nor U11557 (N_11557,N_11364,N_11400);
and U11558 (N_11558,N_11267,N_11407);
nor U11559 (N_11559,N_11448,N_11322);
and U11560 (N_11560,N_11411,N_11429);
or U11561 (N_11561,N_11336,N_11300);
or U11562 (N_11562,N_11350,N_11409);
and U11563 (N_11563,N_11437,N_11475);
or U11564 (N_11564,N_11478,N_11299);
xor U11565 (N_11565,N_11419,N_11253);
xor U11566 (N_11566,N_11394,N_11459);
xnor U11567 (N_11567,N_11441,N_11280);
xor U11568 (N_11568,N_11320,N_11362);
nand U11569 (N_11569,N_11472,N_11399);
and U11570 (N_11570,N_11384,N_11360);
and U11571 (N_11571,N_11326,N_11303);
nand U11572 (N_11572,N_11295,N_11406);
nand U11573 (N_11573,N_11446,N_11387);
nand U11574 (N_11574,N_11325,N_11397);
nor U11575 (N_11575,N_11374,N_11464);
nand U11576 (N_11576,N_11435,N_11366);
and U11577 (N_11577,N_11420,N_11426);
nor U11578 (N_11578,N_11460,N_11404);
or U11579 (N_11579,N_11433,N_11470);
and U11580 (N_11580,N_11485,N_11496);
nand U11581 (N_11581,N_11388,N_11462);
nand U11582 (N_11582,N_11301,N_11390);
and U11583 (N_11583,N_11417,N_11261);
nor U11584 (N_11584,N_11482,N_11310);
or U11585 (N_11585,N_11431,N_11456);
nor U11586 (N_11586,N_11282,N_11307);
nor U11587 (N_11587,N_11289,N_11341);
and U11588 (N_11588,N_11345,N_11283);
nand U11589 (N_11589,N_11405,N_11288);
or U11590 (N_11590,N_11403,N_11358);
xnor U11591 (N_11591,N_11481,N_11436);
and U11592 (N_11592,N_11343,N_11425);
and U11593 (N_11593,N_11402,N_11438);
xor U11594 (N_11594,N_11371,N_11495);
and U11595 (N_11595,N_11257,N_11330);
and U11596 (N_11596,N_11444,N_11255);
or U11597 (N_11597,N_11263,N_11294);
xnor U11598 (N_11598,N_11279,N_11259);
nor U11599 (N_11599,N_11271,N_11385);
xor U11600 (N_11600,N_11492,N_11376);
and U11601 (N_11601,N_11423,N_11382);
or U11602 (N_11602,N_11311,N_11363);
and U11603 (N_11603,N_11347,N_11393);
or U11604 (N_11604,N_11276,N_11383);
and U11605 (N_11605,N_11479,N_11262);
xor U11606 (N_11606,N_11274,N_11473);
xor U11607 (N_11607,N_11372,N_11254);
or U11608 (N_11608,N_11497,N_11477);
nor U11609 (N_11609,N_11412,N_11252);
xor U11610 (N_11610,N_11494,N_11266);
nand U11611 (N_11611,N_11273,N_11312);
nor U11612 (N_11612,N_11476,N_11428);
nand U11613 (N_11613,N_11352,N_11314);
nor U11614 (N_11614,N_11452,N_11471);
nor U11615 (N_11615,N_11342,N_11359);
xor U11616 (N_11616,N_11286,N_11488);
xnor U11617 (N_11617,N_11469,N_11285);
nor U11618 (N_11618,N_11264,N_11461);
nor U11619 (N_11619,N_11367,N_11474);
nand U11620 (N_11620,N_11357,N_11414);
or U11621 (N_11621,N_11309,N_11427);
nand U11622 (N_11622,N_11290,N_11354);
or U11623 (N_11623,N_11445,N_11391);
nand U11624 (N_11624,N_11323,N_11313);
or U11625 (N_11625,N_11416,N_11465);
and U11626 (N_11626,N_11399,N_11285);
nor U11627 (N_11627,N_11334,N_11490);
and U11628 (N_11628,N_11319,N_11317);
or U11629 (N_11629,N_11449,N_11276);
xnor U11630 (N_11630,N_11467,N_11359);
xor U11631 (N_11631,N_11363,N_11489);
nor U11632 (N_11632,N_11311,N_11373);
or U11633 (N_11633,N_11283,N_11335);
nand U11634 (N_11634,N_11484,N_11480);
or U11635 (N_11635,N_11338,N_11368);
xor U11636 (N_11636,N_11455,N_11400);
xnor U11637 (N_11637,N_11490,N_11276);
and U11638 (N_11638,N_11428,N_11319);
nand U11639 (N_11639,N_11499,N_11274);
and U11640 (N_11640,N_11340,N_11276);
xor U11641 (N_11641,N_11466,N_11268);
nor U11642 (N_11642,N_11481,N_11268);
or U11643 (N_11643,N_11379,N_11334);
nor U11644 (N_11644,N_11368,N_11351);
or U11645 (N_11645,N_11471,N_11415);
or U11646 (N_11646,N_11323,N_11264);
nor U11647 (N_11647,N_11419,N_11482);
or U11648 (N_11648,N_11312,N_11275);
nand U11649 (N_11649,N_11476,N_11336);
or U11650 (N_11650,N_11416,N_11463);
nand U11651 (N_11651,N_11265,N_11302);
nor U11652 (N_11652,N_11354,N_11305);
xnor U11653 (N_11653,N_11283,N_11479);
xor U11654 (N_11654,N_11315,N_11363);
nor U11655 (N_11655,N_11435,N_11313);
nor U11656 (N_11656,N_11325,N_11459);
nand U11657 (N_11657,N_11411,N_11267);
nand U11658 (N_11658,N_11262,N_11433);
and U11659 (N_11659,N_11292,N_11444);
xor U11660 (N_11660,N_11424,N_11379);
xor U11661 (N_11661,N_11383,N_11412);
and U11662 (N_11662,N_11446,N_11452);
or U11663 (N_11663,N_11303,N_11345);
or U11664 (N_11664,N_11445,N_11250);
nand U11665 (N_11665,N_11349,N_11407);
nand U11666 (N_11666,N_11321,N_11442);
and U11667 (N_11667,N_11424,N_11291);
or U11668 (N_11668,N_11360,N_11300);
nand U11669 (N_11669,N_11466,N_11471);
xor U11670 (N_11670,N_11451,N_11475);
xnor U11671 (N_11671,N_11277,N_11283);
xor U11672 (N_11672,N_11409,N_11259);
nand U11673 (N_11673,N_11332,N_11373);
or U11674 (N_11674,N_11369,N_11429);
nor U11675 (N_11675,N_11499,N_11317);
xor U11676 (N_11676,N_11251,N_11291);
xnor U11677 (N_11677,N_11273,N_11306);
and U11678 (N_11678,N_11337,N_11418);
xnor U11679 (N_11679,N_11471,N_11495);
nor U11680 (N_11680,N_11294,N_11362);
nand U11681 (N_11681,N_11433,N_11420);
or U11682 (N_11682,N_11265,N_11435);
or U11683 (N_11683,N_11388,N_11313);
nand U11684 (N_11684,N_11375,N_11261);
and U11685 (N_11685,N_11471,N_11467);
xor U11686 (N_11686,N_11463,N_11397);
nand U11687 (N_11687,N_11415,N_11329);
nand U11688 (N_11688,N_11324,N_11484);
nor U11689 (N_11689,N_11356,N_11352);
nand U11690 (N_11690,N_11352,N_11427);
nand U11691 (N_11691,N_11486,N_11301);
xor U11692 (N_11692,N_11451,N_11258);
nand U11693 (N_11693,N_11253,N_11481);
nor U11694 (N_11694,N_11267,N_11250);
or U11695 (N_11695,N_11461,N_11415);
and U11696 (N_11696,N_11367,N_11487);
xnor U11697 (N_11697,N_11457,N_11278);
nand U11698 (N_11698,N_11318,N_11321);
nand U11699 (N_11699,N_11383,N_11258);
xnor U11700 (N_11700,N_11378,N_11304);
and U11701 (N_11701,N_11420,N_11348);
or U11702 (N_11702,N_11283,N_11395);
nand U11703 (N_11703,N_11357,N_11376);
nand U11704 (N_11704,N_11265,N_11489);
and U11705 (N_11705,N_11444,N_11378);
xnor U11706 (N_11706,N_11280,N_11422);
xnor U11707 (N_11707,N_11289,N_11482);
xor U11708 (N_11708,N_11499,N_11416);
nand U11709 (N_11709,N_11329,N_11268);
xnor U11710 (N_11710,N_11413,N_11312);
xnor U11711 (N_11711,N_11411,N_11399);
or U11712 (N_11712,N_11340,N_11320);
or U11713 (N_11713,N_11396,N_11279);
nor U11714 (N_11714,N_11416,N_11433);
xor U11715 (N_11715,N_11342,N_11486);
nor U11716 (N_11716,N_11368,N_11342);
or U11717 (N_11717,N_11371,N_11265);
and U11718 (N_11718,N_11295,N_11491);
nand U11719 (N_11719,N_11435,N_11434);
and U11720 (N_11720,N_11354,N_11395);
nor U11721 (N_11721,N_11496,N_11418);
xor U11722 (N_11722,N_11333,N_11372);
nor U11723 (N_11723,N_11468,N_11406);
xor U11724 (N_11724,N_11444,N_11302);
and U11725 (N_11725,N_11252,N_11337);
or U11726 (N_11726,N_11283,N_11387);
nor U11727 (N_11727,N_11480,N_11323);
and U11728 (N_11728,N_11428,N_11316);
nand U11729 (N_11729,N_11260,N_11399);
nor U11730 (N_11730,N_11296,N_11488);
nor U11731 (N_11731,N_11446,N_11279);
or U11732 (N_11732,N_11470,N_11292);
or U11733 (N_11733,N_11281,N_11406);
and U11734 (N_11734,N_11287,N_11302);
nand U11735 (N_11735,N_11389,N_11365);
or U11736 (N_11736,N_11483,N_11369);
or U11737 (N_11737,N_11407,N_11343);
nor U11738 (N_11738,N_11373,N_11297);
and U11739 (N_11739,N_11323,N_11491);
and U11740 (N_11740,N_11327,N_11261);
xnor U11741 (N_11741,N_11441,N_11495);
and U11742 (N_11742,N_11345,N_11362);
or U11743 (N_11743,N_11368,N_11253);
xnor U11744 (N_11744,N_11364,N_11375);
xnor U11745 (N_11745,N_11329,N_11385);
and U11746 (N_11746,N_11347,N_11289);
and U11747 (N_11747,N_11492,N_11403);
nand U11748 (N_11748,N_11457,N_11368);
and U11749 (N_11749,N_11403,N_11459);
and U11750 (N_11750,N_11615,N_11690);
nand U11751 (N_11751,N_11712,N_11705);
nor U11752 (N_11752,N_11646,N_11566);
or U11753 (N_11753,N_11735,N_11510);
nor U11754 (N_11754,N_11626,N_11533);
xor U11755 (N_11755,N_11663,N_11513);
nand U11756 (N_11756,N_11664,N_11744);
xor U11757 (N_11757,N_11639,N_11674);
nand U11758 (N_11758,N_11700,N_11512);
or U11759 (N_11759,N_11545,N_11643);
or U11760 (N_11760,N_11551,N_11514);
and U11761 (N_11761,N_11586,N_11628);
xnor U11762 (N_11762,N_11677,N_11549);
and U11763 (N_11763,N_11501,N_11678);
nand U11764 (N_11764,N_11613,N_11717);
or U11765 (N_11765,N_11647,N_11618);
and U11766 (N_11766,N_11668,N_11652);
xnor U11767 (N_11767,N_11509,N_11522);
nand U11768 (N_11768,N_11547,N_11746);
nand U11769 (N_11769,N_11593,N_11588);
or U11770 (N_11770,N_11644,N_11711);
nand U11771 (N_11771,N_11623,N_11536);
nand U11772 (N_11772,N_11607,N_11595);
nor U11773 (N_11773,N_11511,N_11737);
nand U11774 (N_11774,N_11503,N_11584);
nor U11775 (N_11775,N_11714,N_11600);
nand U11776 (N_11776,N_11506,N_11552);
or U11777 (N_11777,N_11715,N_11686);
nand U11778 (N_11778,N_11599,N_11624);
or U11779 (N_11779,N_11697,N_11520);
xnor U11780 (N_11780,N_11631,N_11548);
nor U11781 (N_11781,N_11537,N_11743);
nand U11782 (N_11782,N_11614,N_11728);
xor U11783 (N_11783,N_11634,N_11702);
and U11784 (N_11784,N_11565,N_11666);
or U11785 (N_11785,N_11562,N_11608);
or U11786 (N_11786,N_11541,N_11538);
xnor U11787 (N_11787,N_11683,N_11687);
nor U11788 (N_11788,N_11721,N_11703);
nor U11789 (N_11789,N_11649,N_11658);
or U11790 (N_11790,N_11741,N_11730);
xor U11791 (N_11791,N_11692,N_11617);
or U11792 (N_11792,N_11578,N_11740);
or U11793 (N_11793,N_11570,N_11580);
and U11794 (N_11794,N_11502,N_11603);
nor U11795 (N_11795,N_11555,N_11528);
nor U11796 (N_11796,N_11519,N_11560);
nand U11797 (N_11797,N_11637,N_11553);
or U11798 (N_11798,N_11694,N_11561);
nor U11799 (N_11799,N_11656,N_11747);
nor U11800 (N_11800,N_11530,N_11726);
or U11801 (N_11801,N_11587,N_11689);
xnor U11802 (N_11802,N_11698,N_11675);
nor U11803 (N_11803,N_11535,N_11736);
xor U11804 (N_11804,N_11558,N_11591);
and U11805 (N_11805,N_11660,N_11679);
nand U11806 (N_11806,N_11575,N_11665);
or U11807 (N_11807,N_11708,N_11699);
nand U11808 (N_11808,N_11713,N_11738);
and U11809 (N_11809,N_11590,N_11636);
or U11810 (N_11810,N_11707,N_11706);
nand U11811 (N_11811,N_11655,N_11567);
nand U11812 (N_11812,N_11685,N_11640);
nand U11813 (N_11813,N_11724,N_11622);
xor U11814 (N_11814,N_11582,N_11568);
nand U11815 (N_11815,N_11517,N_11629);
xnor U11816 (N_11816,N_11554,N_11709);
nor U11817 (N_11817,N_11596,N_11598);
nor U11818 (N_11818,N_11657,N_11592);
and U11819 (N_11819,N_11748,N_11589);
xnor U11820 (N_11820,N_11659,N_11563);
and U11821 (N_11821,N_11653,N_11627);
xnor U11822 (N_11822,N_11544,N_11516);
and U11823 (N_11823,N_11635,N_11564);
xor U11824 (N_11824,N_11667,N_11524);
xnor U11825 (N_11825,N_11621,N_11662);
or U11826 (N_11826,N_11576,N_11572);
and U11827 (N_11827,N_11556,N_11543);
nor U11828 (N_11828,N_11739,N_11727);
nand U11829 (N_11829,N_11557,N_11612);
nand U11830 (N_11830,N_11693,N_11725);
nor U11831 (N_11831,N_11710,N_11569);
xor U11832 (N_11832,N_11508,N_11645);
nor U11833 (N_11833,N_11505,N_11515);
xnor U11834 (N_11834,N_11648,N_11527);
or U11835 (N_11835,N_11749,N_11731);
and U11836 (N_11836,N_11732,N_11550);
nand U11837 (N_11837,N_11585,N_11688);
and U11838 (N_11838,N_11681,N_11734);
and U11839 (N_11839,N_11542,N_11573);
or U11840 (N_11840,N_11540,N_11610);
and U11841 (N_11841,N_11641,N_11500);
nor U11842 (N_11842,N_11745,N_11716);
nand U11843 (N_11843,N_11650,N_11531);
nand U11844 (N_11844,N_11718,N_11597);
nand U11845 (N_11845,N_11526,N_11701);
and U11846 (N_11846,N_11534,N_11671);
nand U11847 (N_11847,N_11720,N_11642);
and U11848 (N_11848,N_11611,N_11594);
nor U11849 (N_11849,N_11729,N_11722);
or U11850 (N_11850,N_11619,N_11521);
nand U11851 (N_11851,N_11633,N_11577);
or U11852 (N_11852,N_11601,N_11684);
and U11853 (N_11853,N_11625,N_11507);
or U11854 (N_11854,N_11695,N_11680);
nand U11855 (N_11855,N_11574,N_11525);
or U11856 (N_11856,N_11673,N_11696);
nor U11857 (N_11857,N_11704,N_11632);
nand U11858 (N_11858,N_11654,N_11532);
and U11859 (N_11859,N_11602,N_11606);
nand U11860 (N_11860,N_11669,N_11638);
nand U11861 (N_11861,N_11742,N_11539);
nand U11862 (N_11862,N_11723,N_11719);
nand U11863 (N_11863,N_11546,N_11518);
nor U11864 (N_11864,N_11609,N_11583);
nand U11865 (N_11865,N_11616,N_11571);
nor U11866 (N_11866,N_11672,N_11676);
xor U11867 (N_11867,N_11559,N_11579);
nand U11868 (N_11868,N_11504,N_11523);
or U11869 (N_11869,N_11529,N_11630);
nand U11870 (N_11870,N_11604,N_11691);
xor U11871 (N_11871,N_11581,N_11661);
xnor U11872 (N_11872,N_11682,N_11620);
and U11873 (N_11873,N_11651,N_11733);
nor U11874 (N_11874,N_11670,N_11605);
and U11875 (N_11875,N_11607,N_11551);
or U11876 (N_11876,N_11554,N_11608);
nor U11877 (N_11877,N_11512,N_11534);
xor U11878 (N_11878,N_11541,N_11748);
or U11879 (N_11879,N_11653,N_11709);
or U11880 (N_11880,N_11663,N_11530);
nor U11881 (N_11881,N_11672,N_11502);
nand U11882 (N_11882,N_11579,N_11725);
and U11883 (N_11883,N_11689,N_11687);
and U11884 (N_11884,N_11648,N_11617);
nand U11885 (N_11885,N_11583,N_11606);
nand U11886 (N_11886,N_11511,N_11717);
xor U11887 (N_11887,N_11505,N_11702);
or U11888 (N_11888,N_11668,N_11715);
xor U11889 (N_11889,N_11502,N_11732);
or U11890 (N_11890,N_11643,N_11517);
nor U11891 (N_11891,N_11585,N_11621);
and U11892 (N_11892,N_11679,N_11553);
xor U11893 (N_11893,N_11558,N_11519);
or U11894 (N_11894,N_11682,N_11556);
and U11895 (N_11895,N_11546,N_11587);
or U11896 (N_11896,N_11711,N_11547);
xnor U11897 (N_11897,N_11743,N_11519);
or U11898 (N_11898,N_11644,N_11720);
or U11899 (N_11899,N_11687,N_11616);
or U11900 (N_11900,N_11585,N_11579);
or U11901 (N_11901,N_11549,N_11520);
nand U11902 (N_11902,N_11721,N_11667);
xor U11903 (N_11903,N_11629,N_11656);
and U11904 (N_11904,N_11648,N_11646);
and U11905 (N_11905,N_11628,N_11528);
nand U11906 (N_11906,N_11620,N_11580);
or U11907 (N_11907,N_11520,N_11546);
xor U11908 (N_11908,N_11695,N_11511);
and U11909 (N_11909,N_11582,N_11643);
or U11910 (N_11910,N_11555,N_11684);
nor U11911 (N_11911,N_11534,N_11714);
nor U11912 (N_11912,N_11683,N_11645);
xor U11913 (N_11913,N_11698,N_11578);
xor U11914 (N_11914,N_11684,N_11682);
and U11915 (N_11915,N_11544,N_11644);
xnor U11916 (N_11916,N_11731,N_11593);
xor U11917 (N_11917,N_11612,N_11651);
or U11918 (N_11918,N_11569,N_11512);
nor U11919 (N_11919,N_11596,N_11535);
or U11920 (N_11920,N_11691,N_11618);
nor U11921 (N_11921,N_11614,N_11678);
nor U11922 (N_11922,N_11695,N_11738);
and U11923 (N_11923,N_11559,N_11561);
and U11924 (N_11924,N_11501,N_11648);
nor U11925 (N_11925,N_11597,N_11673);
xor U11926 (N_11926,N_11573,N_11535);
or U11927 (N_11927,N_11523,N_11633);
and U11928 (N_11928,N_11517,N_11505);
xor U11929 (N_11929,N_11511,N_11608);
xnor U11930 (N_11930,N_11646,N_11537);
and U11931 (N_11931,N_11718,N_11685);
and U11932 (N_11932,N_11701,N_11624);
or U11933 (N_11933,N_11749,N_11534);
nand U11934 (N_11934,N_11698,N_11519);
xor U11935 (N_11935,N_11718,N_11651);
or U11936 (N_11936,N_11566,N_11737);
nand U11937 (N_11937,N_11591,N_11530);
nand U11938 (N_11938,N_11699,N_11507);
nor U11939 (N_11939,N_11595,N_11739);
and U11940 (N_11940,N_11524,N_11539);
nor U11941 (N_11941,N_11527,N_11532);
xnor U11942 (N_11942,N_11529,N_11728);
or U11943 (N_11943,N_11632,N_11579);
xnor U11944 (N_11944,N_11647,N_11708);
nor U11945 (N_11945,N_11535,N_11695);
xnor U11946 (N_11946,N_11636,N_11697);
nand U11947 (N_11947,N_11749,N_11662);
xor U11948 (N_11948,N_11655,N_11738);
and U11949 (N_11949,N_11646,N_11685);
or U11950 (N_11950,N_11558,N_11536);
nand U11951 (N_11951,N_11579,N_11634);
and U11952 (N_11952,N_11594,N_11736);
nand U11953 (N_11953,N_11557,N_11642);
nor U11954 (N_11954,N_11500,N_11656);
xor U11955 (N_11955,N_11675,N_11637);
nand U11956 (N_11956,N_11663,N_11684);
and U11957 (N_11957,N_11585,N_11690);
or U11958 (N_11958,N_11626,N_11741);
xnor U11959 (N_11959,N_11523,N_11565);
nor U11960 (N_11960,N_11523,N_11667);
or U11961 (N_11961,N_11573,N_11730);
nand U11962 (N_11962,N_11693,N_11644);
nor U11963 (N_11963,N_11708,N_11651);
nand U11964 (N_11964,N_11500,N_11662);
or U11965 (N_11965,N_11504,N_11627);
xor U11966 (N_11966,N_11744,N_11597);
nor U11967 (N_11967,N_11729,N_11600);
nor U11968 (N_11968,N_11638,N_11673);
or U11969 (N_11969,N_11601,N_11612);
and U11970 (N_11970,N_11733,N_11597);
and U11971 (N_11971,N_11544,N_11558);
xor U11972 (N_11972,N_11692,N_11540);
nand U11973 (N_11973,N_11676,N_11549);
and U11974 (N_11974,N_11731,N_11528);
and U11975 (N_11975,N_11536,N_11504);
xnor U11976 (N_11976,N_11593,N_11607);
or U11977 (N_11977,N_11590,N_11509);
and U11978 (N_11978,N_11731,N_11618);
nand U11979 (N_11979,N_11681,N_11665);
xor U11980 (N_11980,N_11602,N_11615);
xor U11981 (N_11981,N_11535,N_11657);
or U11982 (N_11982,N_11591,N_11571);
xnor U11983 (N_11983,N_11723,N_11704);
and U11984 (N_11984,N_11548,N_11643);
and U11985 (N_11985,N_11504,N_11650);
xor U11986 (N_11986,N_11710,N_11668);
xnor U11987 (N_11987,N_11741,N_11617);
nor U11988 (N_11988,N_11683,N_11543);
or U11989 (N_11989,N_11620,N_11652);
or U11990 (N_11990,N_11722,N_11737);
and U11991 (N_11991,N_11580,N_11689);
xor U11992 (N_11992,N_11625,N_11527);
nor U11993 (N_11993,N_11543,N_11569);
or U11994 (N_11994,N_11737,N_11654);
xnor U11995 (N_11995,N_11605,N_11558);
and U11996 (N_11996,N_11617,N_11698);
or U11997 (N_11997,N_11562,N_11538);
nand U11998 (N_11998,N_11695,N_11503);
and U11999 (N_11999,N_11506,N_11694);
or U12000 (N_12000,N_11847,N_11761);
nor U12001 (N_12001,N_11953,N_11956);
and U12002 (N_12002,N_11998,N_11981);
and U12003 (N_12003,N_11987,N_11789);
nor U12004 (N_12004,N_11876,N_11990);
nand U12005 (N_12005,N_11913,N_11862);
nor U12006 (N_12006,N_11817,N_11877);
or U12007 (N_12007,N_11858,N_11982);
nand U12008 (N_12008,N_11965,N_11851);
xnor U12009 (N_12009,N_11841,N_11833);
nand U12010 (N_12010,N_11750,N_11773);
and U12011 (N_12011,N_11929,N_11782);
nand U12012 (N_12012,N_11934,N_11852);
xor U12013 (N_12013,N_11922,N_11801);
nor U12014 (N_12014,N_11888,N_11836);
nor U12015 (N_12015,N_11863,N_11914);
nor U12016 (N_12016,N_11924,N_11798);
or U12017 (N_12017,N_11912,N_11793);
nand U12018 (N_12018,N_11873,N_11860);
nor U12019 (N_12019,N_11875,N_11963);
or U12020 (N_12020,N_11766,N_11949);
and U12021 (N_12021,N_11986,N_11769);
nand U12022 (N_12022,N_11947,N_11822);
or U12023 (N_12023,N_11920,N_11780);
xor U12024 (N_12024,N_11972,N_11848);
nor U12025 (N_12025,N_11967,N_11814);
xor U12026 (N_12026,N_11906,N_11865);
xor U12027 (N_12027,N_11760,N_11805);
nand U12028 (N_12028,N_11806,N_11752);
or U12029 (N_12029,N_11754,N_11838);
nand U12030 (N_12030,N_11980,N_11784);
xor U12031 (N_12031,N_11893,N_11923);
and U12032 (N_12032,N_11942,N_11795);
nor U12033 (N_12033,N_11830,N_11854);
xor U12034 (N_12034,N_11903,N_11753);
xnor U12035 (N_12035,N_11900,N_11962);
nor U12036 (N_12036,N_11964,N_11783);
nand U12037 (N_12037,N_11757,N_11787);
nor U12038 (N_12038,N_11966,N_11910);
or U12039 (N_12039,N_11970,N_11855);
and U12040 (N_12040,N_11997,N_11959);
nor U12041 (N_12041,N_11845,N_11861);
xor U12042 (N_12042,N_11995,N_11973);
and U12043 (N_12043,N_11826,N_11844);
nand U12044 (N_12044,N_11974,N_11908);
or U12045 (N_12045,N_11880,N_11926);
and U12046 (N_12046,N_11802,N_11821);
xor U12047 (N_12047,N_11763,N_11792);
nor U12048 (N_12048,N_11955,N_11808);
or U12049 (N_12049,N_11899,N_11776);
and U12050 (N_12050,N_11897,N_11759);
xnor U12051 (N_12051,N_11879,N_11800);
nor U12052 (N_12052,N_11771,N_11764);
and U12053 (N_12053,N_11796,N_11874);
xnor U12054 (N_12054,N_11777,N_11939);
and U12055 (N_12055,N_11991,N_11868);
and U12056 (N_12056,N_11872,N_11916);
nor U12057 (N_12057,N_11818,N_11775);
xor U12058 (N_12058,N_11992,N_11976);
nand U12059 (N_12059,N_11938,N_11917);
and U12060 (N_12060,N_11930,N_11803);
nor U12061 (N_12061,N_11896,N_11919);
nand U12062 (N_12062,N_11932,N_11807);
nor U12063 (N_12063,N_11898,N_11905);
and U12064 (N_12064,N_11755,N_11827);
nor U12065 (N_12065,N_11902,N_11958);
and U12066 (N_12066,N_11770,N_11767);
xor U12067 (N_12067,N_11975,N_11849);
xor U12068 (N_12068,N_11884,N_11797);
nand U12069 (N_12069,N_11989,N_11889);
xor U12070 (N_12070,N_11940,N_11894);
or U12071 (N_12071,N_11936,N_11892);
xor U12072 (N_12072,N_11960,N_11819);
nand U12073 (N_12073,N_11927,N_11882);
xnor U12074 (N_12074,N_11948,N_11881);
nor U12075 (N_12075,N_11768,N_11774);
or U12076 (N_12076,N_11837,N_11824);
nand U12077 (N_12077,N_11918,N_11957);
xnor U12078 (N_12078,N_11832,N_11895);
or U12079 (N_12079,N_11961,N_11941);
nor U12080 (N_12080,N_11809,N_11968);
xnor U12081 (N_12081,N_11867,N_11781);
nor U12082 (N_12082,N_11788,N_11984);
and U12083 (N_12083,N_11871,N_11977);
and U12084 (N_12084,N_11857,N_11866);
nor U12085 (N_12085,N_11811,N_11887);
and U12086 (N_12086,N_11791,N_11785);
and U12087 (N_12087,N_11907,N_11951);
nor U12088 (N_12088,N_11999,N_11799);
or U12089 (N_12089,N_11765,N_11815);
nor U12090 (N_12090,N_11762,N_11885);
xnor U12091 (N_12091,N_11911,N_11794);
nand U12092 (N_12092,N_11790,N_11846);
or U12093 (N_12093,N_11952,N_11856);
nor U12094 (N_12094,N_11779,N_11834);
nor U12095 (N_12095,N_11820,N_11823);
and U12096 (N_12096,N_11946,N_11979);
and U12097 (N_12097,N_11925,N_11825);
nand U12098 (N_12098,N_11945,N_11869);
nand U12099 (N_12099,N_11835,N_11843);
nand U12100 (N_12100,N_11950,N_11890);
or U12101 (N_12101,N_11853,N_11883);
nand U12102 (N_12102,N_11909,N_11993);
nand U12103 (N_12103,N_11772,N_11928);
nor U12104 (N_12104,N_11969,N_11921);
xnor U12105 (N_12105,N_11971,N_11756);
or U12106 (N_12106,N_11812,N_11778);
or U12107 (N_12107,N_11994,N_11850);
or U12108 (N_12108,N_11816,N_11840);
or U12109 (N_12109,N_11937,N_11751);
xor U12110 (N_12110,N_11985,N_11901);
nand U12111 (N_12111,N_11933,N_11842);
or U12112 (N_12112,N_11859,N_11996);
xor U12113 (N_12113,N_11891,N_11904);
nand U12114 (N_12114,N_11988,N_11831);
and U12115 (N_12115,N_11886,N_11978);
and U12116 (N_12116,N_11804,N_11931);
xnor U12117 (N_12117,N_11839,N_11943);
or U12118 (N_12118,N_11878,N_11758);
nand U12119 (N_12119,N_11954,N_11915);
xor U12120 (N_12120,N_11935,N_11944);
and U12121 (N_12121,N_11810,N_11983);
xnor U12122 (N_12122,N_11870,N_11829);
nor U12123 (N_12123,N_11828,N_11813);
nor U12124 (N_12124,N_11786,N_11864);
xnor U12125 (N_12125,N_11915,N_11994);
xor U12126 (N_12126,N_11957,N_11960);
or U12127 (N_12127,N_11865,N_11891);
nand U12128 (N_12128,N_11921,N_11794);
nand U12129 (N_12129,N_11823,N_11972);
xnor U12130 (N_12130,N_11956,N_11762);
nand U12131 (N_12131,N_11757,N_11854);
xnor U12132 (N_12132,N_11906,N_11864);
nor U12133 (N_12133,N_11927,N_11801);
and U12134 (N_12134,N_11914,N_11894);
and U12135 (N_12135,N_11913,N_11849);
or U12136 (N_12136,N_11980,N_11879);
nand U12137 (N_12137,N_11877,N_11968);
and U12138 (N_12138,N_11940,N_11980);
xor U12139 (N_12139,N_11880,N_11965);
nor U12140 (N_12140,N_11900,N_11792);
nand U12141 (N_12141,N_11810,N_11976);
or U12142 (N_12142,N_11773,N_11797);
xor U12143 (N_12143,N_11774,N_11916);
xor U12144 (N_12144,N_11782,N_11966);
xor U12145 (N_12145,N_11861,N_11968);
or U12146 (N_12146,N_11910,N_11919);
and U12147 (N_12147,N_11815,N_11981);
nor U12148 (N_12148,N_11792,N_11868);
nor U12149 (N_12149,N_11804,N_11872);
xnor U12150 (N_12150,N_11978,N_11959);
nor U12151 (N_12151,N_11807,N_11893);
nor U12152 (N_12152,N_11851,N_11761);
and U12153 (N_12153,N_11899,N_11897);
xnor U12154 (N_12154,N_11951,N_11886);
and U12155 (N_12155,N_11989,N_11801);
nor U12156 (N_12156,N_11997,N_11866);
nor U12157 (N_12157,N_11805,N_11986);
nand U12158 (N_12158,N_11841,N_11922);
xor U12159 (N_12159,N_11809,N_11890);
nand U12160 (N_12160,N_11775,N_11945);
or U12161 (N_12161,N_11798,N_11774);
nor U12162 (N_12162,N_11868,N_11922);
or U12163 (N_12163,N_11812,N_11860);
nor U12164 (N_12164,N_11904,N_11765);
xnor U12165 (N_12165,N_11995,N_11982);
and U12166 (N_12166,N_11787,N_11999);
nor U12167 (N_12167,N_11958,N_11926);
and U12168 (N_12168,N_11793,N_11992);
xor U12169 (N_12169,N_11954,N_11875);
xnor U12170 (N_12170,N_11966,N_11758);
nor U12171 (N_12171,N_11862,N_11978);
xnor U12172 (N_12172,N_11935,N_11753);
and U12173 (N_12173,N_11897,N_11758);
and U12174 (N_12174,N_11801,N_11880);
and U12175 (N_12175,N_11808,N_11851);
nand U12176 (N_12176,N_11870,N_11838);
nand U12177 (N_12177,N_11799,N_11755);
nor U12178 (N_12178,N_11782,N_11794);
and U12179 (N_12179,N_11962,N_11866);
xnor U12180 (N_12180,N_11934,N_11770);
and U12181 (N_12181,N_11805,N_11919);
or U12182 (N_12182,N_11796,N_11957);
nand U12183 (N_12183,N_11983,N_11825);
or U12184 (N_12184,N_11794,N_11753);
xnor U12185 (N_12185,N_11906,N_11924);
nor U12186 (N_12186,N_11958,N_11791);
xor U12187 (N_12187,N_11950,N_11977);
xor U12188 (N_12188,N_11818,N_11927);
or U12189 (N_12189,N_11972,N_11800);
or U12190 (N_12190,N_11902,N_11778);
xor U12191 (N_12191,N_11825,N_11984);
xnor U12192 (N_12192,N_11884,N_11885);
xnor U12193 (N_12193,N_11832,N_11889);
or U12194 (N_12194,N_11800,N_11837);
xor U12195 (N_12195,N_11923,N_11796);
xnor U12196 (N_12196,N_11919,N_11901);
xor U12197 (N_12197,N_11923,N_11808);
and U12198 (N_12198,N_11768,N_11834);
and U12199 (N_12199,N_11833,N_11788);
nand U12200 (N_12200,N_11912,N_11957);
xor U12201 (N_12201,N_11896,N_11892);
nor U12202 (N_12202,N_11874,N_11895);
or U12203 (N_12203,N_11765,N_11906);
nand U12204 (N_12204,N_11896,N_11978);
nor U12205 (N_12205,N_11909,N_11887);
or U12206 (N_12206,N_11849,N_11955);
and U12207 (N_12207,N_11914,N_11772);
and U12208 (N_12208,N_11779,N_11809);
or U12209 (N_12209,N_11979,N_11858);
or U12210 (N_12210,N_11933,N_11820);
or U12211 (N_12211,N_11914,N_11816);
xnor U12212 (N_12212,N_11897,N_11753);
or U12213 (N_12213,N_11857,N_11913);
or U12214 (N_12214,N_11943,N_11818);
or U12215 (N_12215,N_11872,N_11968);
or U12216 (N_12216,N_11931,N_11881);
nand U12217 (N_12217,N_11964,N_11903);
or U12218 (N_12218,N_11881,N_11833);
or U12219 (N_12219,N_11957,N_11819);
and U12220 (N_12220,N_11969,N_11811);
or U12221 (N_12221,N_11990,N_11900);
or U12222 (N_12222,N_11892,N_11930);
xor U12223 (N_12223,N_11954,N_11777);
or U12224 (N_12224,N_11865,N_11800);
and U12225 (N_12225,N_11780,N_11772);
xnor U12226 (N_12226,N_11920,N_11873);
and U12227 (N_12227,N_11811,N_11801);
or U12228 (N_12228,N_11977,N_11899);
nor U12229 (N_12229,N_11982,N_11822);
nor U12230 (N_12230,N_11898,N_11941);
xnor U12231 (N_12231,N_11983,N_11901);
nor U12232 (N_12232,N_11965,N_11767);
nand U12233 (N_12233,N_11844,N_11994);
or U12234 (N_12234,N_11973,N_11833);
xnor U12235 (N_12235,N_11910,N_11965);
xor U12236 (N_12236,N_11848,N_11844);
nand U12237 (N_12237,N_11925,N_11969);
or U12238 (N_12238,N_11810,N_11804);
nor U12239 (N_12239,N_11875,N_11863);
nor U12240 (N_12240,N_11810,N_11799);
and U12241 (N_12241,N_11946,N_11940);
and U12242 (N_12242,N_11859,N_11884);
xnor U12243 (N_12243,N_11844,N_11997);
nand U12244 (N_12244,N_11839,N_11878);
xor U12245 (N_12245,N_11898,N_11809);
nand U12246 (N_12246,N_11888,N_11983);
nand U12247 (N_12247,N_11794,N_11919);
or U12248 (N_12248,N_11767,N_11893);
or U12249 (N_12249,N_11871,N_11862);
nor U12250 (N_12250,N_12204,N_12197);
or U12251 (N_12251,N_12013,N_12120);
or U12252 (N_12252,N_12226,N_12163);
and U12253 (N_12253,N_12168,N_12187);
or U12254 (N_12254,N_12244,N_12135);
or U12255 (N_12255,N_12094,N_12172);
nand U12256 (N_12256,N_12085,N_12096);
nand U12257 (N_12257,N_12084,N_12223);
xor U12258 (N_12258,N_12051,N_12021);
xor U12259 (N_12259,N_12067,N_12224);
and U12260 (N_12260,N_12151,N_12031);
nand U12261 (N_12261,N_12140,N_12235);
nor U12262 (N_12262,N_12158,N_12178);
xor U12263 (N_12263,N_12141,N_12248);
or U12264 (N_12264,N_12008,N_12028);
nand U12265 (N_12265,N_12077,N_12220);
nand U12266 (N_12266,N_12167,N_12227);
xnor U12267 (N_12267,N_12184,N_12225);
and U12268 (N_12268,N_12059,N_12114);
or U12269 (N_12269,N_12162,N_12170);
nand U12270 (N_12270,N_12132,N_12033);
nand U12271 (N_12271,N_12069,N_12211);
nor U12272 (N_12272,N_12221,N_12207);
nor U12273 (N_12273,N_12046,N_12029);
xor U12274 (N_12274,N_12236,N_12053);
nor U12275 (N_12275,N_12019,N_12144);
and U12276 (N_12276,N_12200,N_12115);
or U12277 (N_12277,N_12125,N_12009);
and U12278 (N_12278,N_12149,N_12217);
xor U12279 (N_12279,N_12075,N_12093);
nand U12280 (N_12280,N_12107,N_12025);
xor U12281 (N_12281,N_12157,N_12102);
or U12282 (N_12282,N_12123,N_12188);
nor U12283 (N_12283,N_12012,N_12035);
xnor U12284 (N_12284,N_12130,N_12193);
or U12285 (N_12285,N_12048,N_12159);
nand U12286 (N_12286,N_12185,N_12002);
nor U12287 (N_12287,N_12044,N_12148);
or U12288 (N_12288,N_12216,N_12212);
xnor U12289 (N_12289,N_12209,N_12198);
nand U12290 (N_12290,N_12128,N_12082);
or U12291 (N_12291,N_12108,N_12218);
nand U12292 (N_12292,N_12106,N_12234);
xnor U12293 (N_12293,N_12228,N_12214);
or U12294 (N_12294,N_12119,N_12232);
xnor U12295 (N_12295,N_12181,N_12003);
nor U12296 (N_12296,N_12074,N_12047);
nand U12297 (N_12297,N_12192,N_12055);
nor U12298 (N_12298,N_12071,N_12063);
nor U12299 (N_12299,N_12186,N_12166);
or U12300 (N_12300,N_12231,N_12097);
nor U12301 (N_12301,N_12081,N_12073);
xor U12302 (N_12302,N_12177,N_12110);
and U12303 (N_12303,N_12049,N_12099);
xnor U12304 (N_12304,N_12026,N_12092);
and U12305 (N_12305,N_12023,N_12233);
nand U12306 (N_12306,N_12241,N_12183);
and U12307 (N_12307,N_12210,N_12062);
nor U12308 (N_12308,N_12165,N_12057);
nor U12309 (N_12309,N_12152,N_12202);
or U12310 (N_12310,N_12190,N_12040);
and U12311 (N_12311,N_12004,N_12061);
xor U12312 (N_12312,N_12189,N_12169);
nand U12313 (N_12313,N_12038,N_12127);
nor U12314 (N_12314,N_12180,N_12112);
or U12315 (N_12315,N_12247,N_12032);
xnor U12316 (N_12316,N_12111,N_12215);
nor U12317 (N_12317,N_12179,N_12142);
and U12318 (N_12318,N_12042,N_12175);
nand U12319 (N_12319,N_12124,N_12100);
nor U12320 (N_12320,N_12027,N_12230);
nand U12321 (N_12321,N_12079,N_12060);
nand U12322 (N_12322,N_12146,N_12139);
or U12323 (N_12323,N_12199,N_12000);
or U12324 (N_12324,N_12229,N_12072);
or U12325 (N_12325,N_12137,N_12249);
nor U12326 (N_12326,N_12155,N_12246);
xnor U12327 (N_12327,N_12015,N_12087);
xnor U12328 (N_12328,N_12037,N_12182);
nor U12329 (N_12329,N_12153,N_12070);
nand U12330 (N_12330,N_12150,N_12054);
nand U12331 (N_12331,N_12131,N_12006);
and U12332 (N_12332,N_12173,N_12203);
or U12333 (N_12333,N_12143,N_12147);
or U12334 (N_12334,N_12208,N_12016);
nor U12335 (N_12335,N_12089,N_12036);
or U12336 (N_12336,N_12104,N_12076);
and U12337 (N_12337,N_12091,N_12161);
and U12338 (N_12338,N_12043,N_12064);
nor U12339 (N_12339,N_12039,N_12121);
xor U12340 (N_12340,N_12138,N_12205);
nor U12341 (N_12341,N_12238,N_12239);
nor U12342 (N_12342,N_12219,N_12007);
or U12343 (N_12343,N_12014,N_12237);
and U12344 (N_12344,N_12206,N_12171);
nor U12345 (N_12345,N_12136,N_12129);
xor U12346 (N_12346,N_12196,N_12242);
and U12347 (N_12347,N_12164,N_12117);
and U12348 (N_12348,N_12020,N_12160);
xor U12349 (N_12349,N_12001,N_12095);
and U12350 (N_12350,N_12105,N_12066);
and U12351 (N_12351,N_12056,N_12113);
nand U12352 (N_12352,N_12011,N_12195);
nor U12353 (N_12353,N_12068,N_12080);
nor U12354 (N_12354,N_12116,N_12240);
nand U12355 (N_12355,N_12194,N_12034);
and U12356 (N_12356,N_12213,N_12017);
and U12357 (N_12357,N_12058,N_12078);
and U12358 (N_12358,N_12145,N_12101);
or U12359 (N_12359,N_12134,N_12098);
xnor U12360 (N_12360,N_12090,N_12022);
and U12361 (N_12361,N_12030,N_12118);
or U12362 (N_12362,N_12050,N_12018);
nor U12363 (N_12363,N_12010,N_12103);
nand U12364 (N_12364,N_12052,N_12176);
or U12365 (N_12365,N_12041,N_12245);
nand U12366 (N_12366,N_12154,N_12086);
xor U12367 (N_12367,N_12156,N_12191);
and U12368 (N_12368,N_12122,N_12045);
and U12369 (N_12369,N_12243,N_12083);
nor U12370 (N_12370,N_12126,N_12088);
xor U12371 (N_12371,N_12065,N_12222);
and U12372 (N_12372,N_12005,N_12133);
or U12373 (N_12373,N_12024,N_12174);
nand U12374 (N_12374,N_12109,N_12201);
or U12375 (N_12375,N_12152,N_12080);
nand U12376 (N_12376,N_12210,N_12130);
and U12377 (N_12377,N_12127,N_12094);
nand U12378 (N_12378,N_12210,N_12224);
xnor U12379 (N_12379,N_12078,N_12212);
or U12380 (N_12380,N_12105,N_12212);
and U12381 (N_12381,N_12028,N_12062);
nor U12382 (N_12382,N_12039,N_12129);
nor U12383 (N_12383,N_12134,N_12056);
xor U12384 (N_12384,N_12155,N_12044);
nor U12385 (N_12385,N_12172,N_12114);
and U12386 (N_12386,N_12240,N_12101);
or U12387 (N_12387,N_12067,N_12063);
and U12388 (N_12388,N_12150,N_12026);
or U12389 (N_12389,N_12110,N_12167);
xor U12390 (N_12390,N_12228,N_12021);
nand U12391 (N_12391,N_12063,N_12210);
xor U12392 (N_12392,N_12123,N_12162);
nor U12393 (N_12393,N_12127,N_12138);
nand U12394 (N_12394,N_12097,N_12249);
xor U12395 (N_12395,N_12082,N_12142);
nand U12396 (N_12396,N_12007,N_12128);
nor U12397 (N_12397,N_12075,N_12229);
and U12398 (N_12398,N_12196,N_12118);
and U12399 (N_12399,N_12148,N_12198);
and U12400 (N_12400,N_12089,N_12124);
nor U12401 (N_12401,N_12203,N_12192);
or U12402 (N_12402,N_12154,N_12071);
and U12403 (N_12403,N_12228,N_12042);
or U12404 (N_12404,N_12134,N_12086);
nand U12405 (N_12405,N_12068,N_12210);
nor U12406 (N_12406,N_12047,N_12065);
and U12407 (N_12407,N_12247,N_12010);
xnor U12408 (N_12408,N_12177,N_12031);
xnor U12409 (N_12409,N_12040,N_12136);
nor U12410 (N_12410,N_12191,N_12053);
xor U12411 (N_12411,N_12050,N_12210);
nor U12412 (N_12412,N_12114,N_12159);
or U12413 (N_12413,N_12231,N_12169);
nor U12414 (N_12414,N_12130,N_12028);
or U12415 (N_12415,N_12111,N_12244);
xor U12416 (N_12416,N_12087,N_12101);
nand U12417 (N_12417,N_12126,N_12098);
and U12418 (N_12418,N_12245,N_12235);
nor U12419 (N_12419,N_12091,N_12198);
and U12420 (N_12420,N_12173,N_12196);
xnor U12421 (N_12421,N_12216,N_12061);
nor U12422 (N_12422,N_12045,N_12148);
or U12423 (N_12423,N_12249,N_12188);
xnor U12424 (N_12424,N_12189,N_12136);
xnor U12425 (N_12425,N_12176,N_12040);
and U12426 (N_12426,N_12011,N_12057);
nor U12427 (N_12427,N_12093,N_12158);
nand U12428 (N_12428,N_12025,N_12133);
nand U12429 (N_12429,N_12116,N_12179);
nor U12430 (N_12430,N_12061,N_12223);
xor U12431 (N_12431,N_12040,N_12006);
or U12432 (N_12432,N_12048,N_12216);
or U12433 (N_12433,N_12209,N_12007);
and U12434 (N_12434,N_12237,N_12229);
xnor U12435 (N_12435,N_12022,N_12072);
and U12436 (N_12436,N_12082,N_12163);
nand U12437 (N_12437,N_12066,N_12043);
nand U12438 (N_12438,N_12056,N_12227);
xnor U12439 (N_12439,N_12125,N_12101);
or U12440 (N_12440,N_12154,N_12135);
nand U12441 (N_12441,N_12164,N_12174);
nor U12442 (N_12442,N_12034,N_12098);
nor U12443 (N_12443,N_12210,N_12074);
and U12444 (N_12444,N_12054,N_12122);
or U12445 (N_12445,N_12215,N_12084);
and U12446 (N_12446,N_12176,N_12216);
or U12447 (N_12447,N_12021,N_12060);
xor U12448 (N_12448,N_12049,N_12144);
and U12449 (N_12449,N_12046,N_12021);
or U12450 (N_12450,N_12213,N_12119);
or U12451 (N_12451,N_12063,N_12196);
nand U12452 (N_12452,N_12245,N_12097);
xnor U12453 (N_12453,N_12010,N_12162);
nor U12454 (N_12454,N_12103,N_12248);
or U12455 (N_12455,N_12219,N_12122);
nand U12456 (N_12456,N_12226,N_12113);
or U12457 (N_12457,N_12103,N_12007);
or U12458 (N_12458,N_12175,N_12092);
and U12459 (N_12459,N_12044,N_12019);
xor U12460 (N_12460,N_12180,N_12145);
nand U12461 (N_12461,N_12118,N_12032);
and U12462 (N_12462,N_12142,N_12024);
nand U12463 (N_12463,N_12006,N_12226);
xor U12464 (N_12464,N_12215,N_12016);
xor U12465 (N_12465,N_12107,N_12056);
xnor U12466 (N_12466,N_12166,N_12113);
and U12467 (N_12467,N_12205,N_12211);
nor U12468 (N_12468,N_12054,N_12056);
xnor U12469 (N_12469,N_12013,N_12011);
or U12470 (N_12470,N_12069,N_12233);
xor U12471 (N_12471,N_12220,N_12164);
or U12472 (N_12472,N_12131,N_12070);
nor U12473 (N_12473,N_12153,N_12158);
and U12474 (N_12474,N_12032,N_12012);
or U12475 (N_12475,N_12086,N_12183);
xor U12476 (N_12476,N_12020,N_12134);
xnor U12477 (N_12477,N_12228,N_12070);
nor U12478 (N_12478,N_12214,N_12149);
nand U12479 (N_12479,N_12059,N_12219);
or U12480 (N_12480,N_12224,N_12243);
xor U12481 (N_12481,N_12162,N_12226);
and U12482 (N_12482,N_12155,N_12238);
and U12483 (N_12483,N_12243,N_12245);
nor U12484 (N_12484,N_12247,N_12113);
nand U12485 (N_12485,N_12134,N_12213);
or U12486 (N_12486,N_12113,N_12180);
and U12487 (N_12487,N_12086,N_12054);
nand U12488 (N_12488,N_12204,N_12062);
nand U12489 (N_12489,N_12040,N_12003);
nor U12490 (N_12490,N_12061,N_12243);
or U12491 (N_12491,N_12213,N_12107);
or U12492 (N_12492,N_12040,N_12242);
and U12493 (N_12493,N_12165,N_12111);
and U12494 (N_12494,N_12072,N_12236);
xnor U12495 (N_12495,N_12130,N_12138);
and U12496 (N_12496,N_12112,N_12096);
nor U12497 (N_12497,N_12175,N_12061);
nor U12498 (N_12498,N_12178,N_12113);
nand U12499 (N_12499,N_12019,N_12081);
and U12500 (N_12500,N_12399,N_12278);
xor U12501 (N_12501,N_12280,N_12462);
xnor U12502 (N_12502,N_12251,N_12290);
nor U12503 (N_12503,N_12275,N_12409);
and U12504 (N_12504,N_12434,N_12433);
and U12505 (N_12505,N_12259,N_12452);
and U12506 (N_12506,N_12358,N_12250);
nor U12507 (N_12507,N_12343,N_12422);
nand U12508 (N_12508,N_12256,N_12401);
nor U12509 (N_12509,N_12306,N_12309);
and U12510 (N_12510,N_12467,N_12387);
and U12511 (N_12511,N_12463,N_12483);
or U12512 (N_12512,N_12430,N_12362);
and U12513 (N_12513,N_12271,N_12455);
nand U12514 (N_12514,N_12487,N_12464);
xnor U12515 (N_12515,N_12421,N_12360);
nor U12516 (N_12516,N_12308,N_12266);
or U12517 (N_12517,N_12338,N_12393);
xnor U12518 (N_12518,N_12375,N_12313);
nand U12519 (N_12519,N_12441,N_12370);
xnor U12520 (N_12520,N_12404,N_12437);
or U12521 (N_12521,N_12276,N_12283);
nor U12522 (N_12522,N_12475,N_12453);
or U12523 (N_12523,N_12357,N_12383);
or U12524 (N_12524,N_12270,N_12395);
or U12525 (N_12525,N_12344,N_12374);
xnor U12526 (N_12526,N_12417,N_12407);
or U12527 (N_12527,N_12296,N_12496);
or U12528 (N_12528,N_12291,N_12398);
nand U12529 (N_12529,N_12397,N_12316);
nand U12530 (N_12530,N_12332,N_12350);
nand U12531 (N_12531,N_12364,N_12402);
xnor U12532 (N_12532,N_12440,N_12341);
and U12533 (N_12533,N_12326,N_12389);
nand U12534 (N_12534,N_12460,N_12448);
or U12535 (N_12535,N_12435,N_12381);
xnor U12536 (N_12536,N_12348,N_12449);
nand U12537 (N_12537,N_12254,N_12314);
nor U12538 (N_12538,N_12493,N_12289);
nand U12539 (N_12539,N_12287,N_12272);
or U12540 (N_12540,N_12408,N_12465);
nand U12541 (N_12541,N_12301,N_12263);
or U12542 (N_12542,N_12253,N_12450);
xnor U12543 (N_12543,N_12292,N_12367);
or U12544 (N_12544,N_12330,N_12443);
xnor U12545 (N_12545,N_12425,N_12413);
or U12546 (N_12546,N_12429,N_12473);
nor U12547 (N_12547,N_12428,N_12390);
nand U12548 (N_12548,N_12325,N_12469);
or U12549 (N_12549,N_12391,N_12486);
or U12550 (N_12550,N_12252,N_12356);
or U12551 (N_12551,N_12300,N_12319);
nor U12552 (N_12552,N_12318,N_12281);
nand U12553 (N_12553,N_12466,N_12478);
or U12554 (N_12554,N_12470,N_12352);
or U12555 (N_12555,N_12376,N_12497);
xnor U12556 (N_12556,N_12371,N_12378);
nand U12557 (N_12557,N_12414,N_12335);
or U12558 (N_12558,N_12365,N_12373);
nand U12559 (N_12559,N_12302,N_12489);
nor U12560 (N_12560,N_12457,N_12471);
nor U12561 (N_12561,N_12264,N_12386);
or U12562 (N_12562,N_12284,N_12353);
or U12563 (N_12563,N_12479,N_12297);
xor U12564 (N_12564,N_12322,N_12285);
nand U12565 (N_12565,N_12416,N_12418);
nor U12566 (N_12566,N_12419,N_12310);
nor U12567 (N_12567,N_12495,N_12260);
xor U12568 (N_12568,N_12359,N_12288);
or U12569 (N_12569,N_12472,N_12342);
xor U12570 (N_12570,N_12477,N_12315);
xnor U12571 (N_12571,N_12476,N_12431);
xnor U12572 (N_12572,N_12262,N_12294);
xnor U12573 (N_12573,N_12355,N_12311);
and U12574 (N_12574,N_12442,N_12267);
xor U12575 (N_12575,N_12377,N_12324);
xnor U12576 (N_12576,N_12480,N_12411);
nand U12577 (N_12577,N_12494,N_12406);
and U12578 (N_12578,N_12459,N_12400);
nand U12579 (N_12579,N_12456,N_12410);
nand U12580 (N_12580,N_12403,N_12312);
nand U12581 (N_12581,N_12498,N_12305);
or U12582 (N_12582,N_12299,N_12423);
nand U12583 (N_12583,N_12307,N_12458);
xor U12584 (N_12584,N_12394,N_12327);
or U12585 (N_12585,N_12303,N_12396);
or U12586 (N_12586,N_12384,N_12277);
nand U12587 (N_12587,N_12369,N_12388);
nor U12588 (N_12588,N_12321,N_12337);
xor U12589 (N_12589,N_12485,N_12499);
and U12590 (N_12590,N_12392,N_12257);
and U12591 (N_12591,N_12363,N_12481);
nand U12592 (N_12592,N_12368,N_12329);
and U12593 (N_12593,N_12286,N_12405);
or U12594 (N_12594,N_12491,N_12454);
nand U12595 (N_12595,N_12345,N_12444);
or U12596 (N_12596,N_12474,N_12468);
and U12597 (N_12597,N_12339,N_12451);
xnor U12598 (N_12598,N_12255,N_12320);
nand U12599 (N_12599,N_12261,N_12492);
or U12600 (N_12600,N_12354,N_12482);
nor U12601 (N_12601,N_12379,N_12427);
and U12602 (N_12602,N_12446,N_12426);
and U12603 (N_12603,N_12382,N_12298);
nand U12604 (N_12604,N_12484,N_12268);
or U12605 (N_12605,N_12323,N_12265);
xnor U12606 (N_12606,N_12385,N_12304);
and U12607 (N_12607,N_12274,N_12488);
and U12608 (N_12608,N_12445,N_12420);
nor U12609 (N_12609,N_12351,N_12415);
or U12610 (N_12610,N_12447,N_12372);
nor U12611 (N_12611,N_12424,N_12412);
xnor U12612 (N_12612,N_12438,N_12461);
or U12613 (N_12613,N_12346,N_12490);
or U12614 (N_12614,N_12340,N_12282);
nor U12615 (N_12615,N_12269,N_12347);
nand U12616 (N_12616,N_12336,N_12331);
or U12617 (N_12617,N_12432,N_12349);
xnor U12618 (N_12618,N_12436,N_12295);
nand U12619 (N_12619,N_12439,N_12333);
and U12620 (N_12620,N_12273,N_12293);
or U12621 (N_12621,N_12366,N_12334);
nand U12622 (N_12622,N_12328,N_12317);
nor U12623 (N_12623,N_12361,N_12279);
nor U12624 (N_12624,N_12380,N_12258);
nand U12625 (N_12625,N_12266,N_12317);
xor U12626 (N_12626,N_12341,N_12301);
nor U12627 (N_12627,N_12419,N_12332);
or U12628 (N_12628,N_12484,N_12443);
nand U12629 (N_12629,N_12306,N_12330);
xor U12630 (N_12630,N_12405,N_12285);
nand U12631 (N_12631,N_12338,N_12459);
or U12632 (N_12632,N_12479,N_12366);
and U12633 (N_12633,N_12490,N_12348);
nand U12634 (N_12634,N_12359,N_12463);
nand U12635 (N_12635,N_12308,N_12450);
xor U12636 (N_12636,N_12442,N_12414);
xnor U12637 (N_12637,N_12361,N_12300);
nand U12638 (N_12638,N_12267,N_12482);
nand U12639 (N_12639,N_12314,N_12256);
nor U12640 (N_12640,N_12364,N_12254);
nand U12641 (N_12641,N_12431,N_12389);
or U12642 (N_12642,N_12428,N_12256);
and U12643 (N_12643,N_12465,N_12258);
xor U12644 (N_12644,N_12482,N_12320);
and U12645 (N_12645,N_12272,N_12349);
or U12646 (N_12646,N_12484,N_12409);
and U12647 (N_12647,N_12417,N_12456);
and U12648 (N_12648,N_12270,N_12314);
or U12649 (N_12649,N_12398,N_12371);
and U12650 (N_12650,N_12266,N_12397);
nand U12651 (N_12651,N_12250,N_12252);
nand U12652 (N_12652,N_12450,N_12478);
and U12653 (N_12653,N_12486,N_12442);
and U12654 (N_12654,N_12322,N_12271);
nor U12655 (N_12655,N_12368,N_12360);
or U12656 (N_12656,N_12353,N_12319);
nor U12657 (N_12657,N_12400,N_12270);
nor U12658 (N_12658,N_12279,N_12402);
or U12659 (N_12659,N_12328,N_12255);
and U12660 (N_12660,N_12303,N_12362);
nor U12661 (N_12661,N_12400,N_12258);
nand U12662 (N_12662,N_12253,N_12290);
nor U12663 (N_12663,N_12297,N_12326);
nand U12664 (N_12664,N_12363,N_12253);
nand U12665 (N_12665,N_12341,N_12319);
nand U12666 (N_12666,N_12253,N_12312);
or U12667 (N_12667,N_12414,N_12260);
nand U12668 (N_12668,N_12263,N_12336);
xnor U12669 (N_12669,N_12377,N_12250);
or U12670 (N_12670,N_12256,N_12307);
or U12671 (N_12671,N_12306,N_12357);
nor U12672 (N_12672,N_12452,N_12368);
xnor U12673 (N_12673,N_12434,N_12361);
nor U12674 (N_12674,N_12484,N_12335);
nor U12675 (N_12675,N_12266,N_12477);
nor U12676 (N_12676,N_12449,N_12306);
nor U12677 (N_12677,N_12486,N_12453);
xor U12678 (N_12678,N_12372,N_12353);
xor U12679 (N_12679,N_12268,N_12410);
nor U12680 (N_12680,N_12272,N_12487);
nand U12681 (N_12681,N_12460,N_12279);
and U12682 (N_12682,N_12434,N_12270);
nand U12683 (N_12683,N_12269,N_12426);
nor U12684 (N_12684,N_12258,N_12278);
or U12685 (N_12685,N_12419,N_12270);
and U12686 (N_12686,N_12418,N_12348);
and U12687 (N_12687,N_12459,N_12499);
and U12688 (N_12688,N_12256,N_12298);
and U12689 (N_12689,N_12475,N_12442);
and U12690 (N_12690,N_12427,N_12465);
nand U12691 (N_12691,N_12397,N_12306);
or U12692 (N_12692,N_12269,N_12255);
nand U12693 (N_12693,N_12340,N_12435);
or U12694 (N_12694,N_12336,N_12412);
nor U12695 (N_12695,N_12461,N_12433);
or U12696 (N_12696,N_12340,N_12305);
nand U12697 (N_12697,N_12298,N_12424);
and U12698 (N_12698,N_12317,N_12420);
or U12699 (N_12699,N_12314,N_12271);
or U12700 (N_12700,N_12481,N_12304);
nor U12701 (N_12701,N_12436,N_12410);
nand U12702 (N_12702,N_12261,N_12461);
and U12703 (N_12703,N_12468,N_12252);
or U12704 (N_12704,N_12280,N_12265);
or U12705 (N_12705,N_12441,N_12296);
nand U12706 (N_12706,N_12251,N_12459);
nand U12707 (N_12707,N_12266,N_12346);
and U12708 (N_12708,N_12449,N_12327);
nand U12709 (N_12709,N_12309,N_12478);
xnor U12710 (N_12710,N_12453,N_12315);
nor U12711 (N_12711,N_12381,N_12253);
nor U12712 (N_12712,N_12267,N_12263);
nand U12713 (N_12713,N_12499,N_12318);
nand U12714 (N_12714,N_12351,N_12314);
nand U12715 (N_12715,N_12328,N_12487);
xor U12716 (N_12716,N_12291,N_12324);
nor U12717 (N_12717,N_12479,N_12262);
and U12718 (N_12718,N_12434,N_12374);
xor U12719 (N_12719,N_12312,N_12359);
nor U12720 (N_12720,N_12286,N_12498);
and U12721 (N_12721,N_12256,N_12294);
nor U12722 (N_12722,N_12283,N_12402);
nand U12723 (N_12723,N_12274,N_12471);
nand U12724 (N_12724,N_12259,N_12481);
nand U12725 (N_12725,N_12367,N_12460);
nand U12726 (N_12726,N_12285,N_12471);
or U12727 (N_12727,N_12305,N_12259);
xor U12728 (N_12728,N_12428,N_12300);
and U12729 (N_12729,N_12413,N_12428);
xnor U12730 (N_12730,N_12357,N_12270);
or U12731 (N_12731,N_12467,N_12319);
xor U12732 (N_12732,N_12499,N_12497);
and U12733 (N_12733,N_12440,N_12360);
or U12734 (N_12734,N_12395,N_12356);
nand U12735 (N_12735,N_12344,N_12323);
xor U12736 (N_12736,N_12438,N_12373);
xor U12737 (N_12737,N_12274,N_12363);
nand U12738 (N_12738,N_12440,N_12395);
or U12739 (N_12739,N_12261,N_12472);
nand U12740 (N_12740,N_12494,N_12420);
xor U12741 (N_12741,N_12462,N_12422);
and U12742 (N_12742,N_12261,N_12358);
xor U12743 (N_12743,N_12304,N_12324);
xnor U12744 (N_12744,N_12478,N_12285);
or U12745 (N_12745,N_12345,N_12361);
or U12746 (N_12746,N_12302,N_12319);
nor U12747 (N_12747,N_12475,N_12250);
nor U12748 (N_12748,N_12330,N_12394);
nor U12749 (N_12749,N_12312,N_12362);
xnor U12750 (N_12750,N_12726,N_12740);
xor U12751 (N_12751,N_12677,N_12539);
xor U12752 (N_12752,N_12631,N_12619);
nor U12753 (N_12753,N_12625,N_12581);
nand U12754 (N_12754,N_12690,N_12506);
or U12755 (N_12755,N_12664,N_12525);
nor U12756 (N_12756,N_12578,N_12545);
and U12757 (N_12757,N_12637,N_12629);
or U12758 (N_12758,N_12662,N_12630);
and U12759 (N_12759,N_12691,N_12661);
nor U12760 (N_12760,N_12674,N_12727);
and U12761 (N_12761,N_12703,N_12533);
nand U12762 (N_12762,N_12715,N_12663);
or U12763 (N_12763,N_12608,N_12747);
nand U12764 (N_12764,N_12504,N_12688);
or U12765 (N_12765,N_12573,N_12659);
or U12766 (N_12766,N_12503,N_12521);
nand U12767 (N_12767,N_12745,N_12732);
xnor U12768 (N_12768,N_12712,N_12556);
nor U12769 (N_12769,N_12591,N_12707);
or U12770 (N_12770,N_12683,N_12656);
nand U12771 (N_12771,N_12620,N_12570);
nor U12772 (N_12772,N_12604,N_12667);
xor U12773 (N_12773,N_12612,N_12529);
xnor U12774 (N_12774,N_12731,N_12669);
nand U12775 (N_12775,N_12537,N_12508);
nand U12776 (N_12776,N_12526,N_12580);
xor U12777 (N_12777,N_12623,N_12511);
nand U12778 (N_12778,N_12559,N_12644);
nand U12779 (N_12779,N_12603,N_12694);
nand U12780 (N_12780,N_12602,N_12743);
nand U12781 (N_12781,N_12558,N_12507);
nor U12782 (N_12782,N_12592,N_12706);
nor U12783 (N_12783,N_12704,N_12519);
or U12784 (N_12784,N_12647,N_12567);
xor U12785 (N_12785,N_12596,N_12512);
xnor U12786 (N_12786,N_12650,N_12717);
nor U12787 (N_12787,N_12571,N_12676);
nor U12788 (N_12788,N_12530,N_12642);
and U12789 (N_12789,N_12682,N_12628);
nand U12790 (N_12790,N_12657,N_12517);
nor U12791 (N_12791,N_12601,N_12611);
nor U12792 (N_12792,N_12749,N_12689);
and U12793 (N_12793,N_12586,N_12505);
or U12794 (N_12794,N_12531,N_12609);
nand U12795 (N_12795,N_12710,N_12624);
xnor U12796 (N_12796,N_12699,N_12648);
and U12797 (N_12797,N_12641,N_12728);
nand U12798 (N_12798,N_12742,N_12554);
xor U12799 (N_12799,N_12720,N_12543);
nand U12800 (N_12800,N_12651,N_12665);
nor U12801 (N_12801,N_12522,N_12686);
nand U12802 (N_12802,N_12627,N_12606);
nor U12803 (N_12803,N_12585,N_12709);
xor U12804 (N_12804,N_12638,N_12536);
or U12805 (N_12805,N_12698,N_12719);
xnor U12806 (N_12806,N_12621,N_12566);
or U12807 (N_12807,N_12741,N_12739);
and U12808 (N_12808,N_12716,N_12675);
and U12809 (N_12809,N_12584,N_12744);
and U12810 (N_12810,N_12668,N_12520);
nor U12811 (N_12811,N_12523,N_12542);
xor U12812 (N_12812,N_12714,N_12713);
nand U12813 (N_12813,N_12516,N_12518);
nand U12814 (N_12814,N_12605,N_12695);
nand U12815 (N_12815,N_12550,N_12737);
nand U12816 (N_12816,N_12509,N_12618);
xnor U12817 (N_12817,N_12733,N_12575);
xnor U12818 (N_12818,N_12538,N_12721);
nor U12819 (N_12819,N_12736,N_12671);
and U12820 (N_12820,N_12600,N_12649);
nand U12821 (N_12821,N_12622,N_12730);
xor U12822 (N_12822,N_12687,N_12541);
and U12823 (N_12823,N_12583,N_12515);
or U12824 (N_12824,N_12660,N_12557);
and U12825 (N_12825,N_12594,N_12501);
nor U12826 (N_12826,N_12685,N_12589);
nand U12827 (N_12827,N_12684,N_12551);
nand U12828 (N_12828,N_12574,N_12572);
or U12829 (N_12829,N_12590,N_12632);
xor U12830 (N_12830,N_12547,N_12577);
nand U12831 (N_12831,N_12673,N_12722);
xor U12832 (N_12832,N_12681,N_12534);
nor U12833 (N_12833,N_12639,N_12718);
or U12834 (N_12834,N_12635,N_12500);
nor U12835 (N_12835,N_12646,N_12535);
nor U12836 (N_12836,N_12640,N_12555);
nand U12837 (N_12837,N_12653,N_12527);
or U12838 (N_12838,N_12725,N_12702);
nor U12839 (N_12839,N_12560,N_12565);
and U12840 (N_12840,N_12697,N_12552);
nor U12841 (N_12841,N_12748,N_12636);
and U12842 (N_12842,N_12546,N_12613);
nor U12843 (N_12843,N_12633,N_12588);
or U12844 (N_12844,N_12658,N_12510);
and U12845 (N_12845,N_12502,N_12666);
nand U12846 (N_12846,N_12734,N_12672);
xnor U12847 (N_12847,N_12654,N_12729);
nor U12848 (N_12848,N_12617,N_12549);
nand U12849 (N_12849,N_12652,N_12569);
xor U12850 (N_12850,N_12607,N_12599);
nor U12851 (N_12851,N_12724,N_12576);
nand U12852 (N_12852,N_12655,N_12705);
or U12853 (N_12853,N_12670,N_12579);
or U12854 (N_12854,N_12564,N_12582);
nor U12855 (N_12855,N_12616,N_12692);
nand U12856 (N_12856,N_12696,N_12643);
nand U12857 (N_12857,N_12598,N_12568);
nand U12858 (N_12858,N_12679,N_12738);
xor U12859 (N_12859,N_12597,N_12561);
or U12860 (N_12860,N_12544,N_12513);
and U12861 (N_12861,N_12700,N_12626);
nor U12862 (N_12862,N_12587,N_12563);
and U12863 (N_12863,N_12524,N_12701);
or U12864 (N_12864,N_12532,N_12678);
xnor U12865 (N_12865,N_12593,N_12514);
or U12866 (N_12866,N_12735,N_12553);
and U12867 (N_12867,N_12711,N_12548);
nand U12868 (N_12868,N_12708,N_12680);
and U12869 (N_12869,N_12562,N_12614);
nand U12870 (N_12870,N_12746,N_12693);
and U12871 (N_12871,N_12645,N_12540);
nor U12872 (N_12872,N_12595,N_12723);
and U12873 (N_12873,N_12610,N_12634);
xor U12874 (N_12874,N_12528,N_12615);
nand U12875 (N_12875,N_12690,N_12535);
nand U12876 (N_12876,N_12556,N_12678);
or U12877 (N_12877,N_12513,N_12593);
nand U12878 (N_12878,N_12571,N_12595);
and U12879 (N_12879,N_12692,N_12707);
or U12880 (N_12880,N_12596,N_12725);
xnor U12881 (N_12881,N_12532,N_12534);
nand U12882 (N_12882,N_12513,N_12549);
nor U12883 (N_12883,N_12705,N_12665);
xnor U12884 (N_12884,N_12721,N_12572);
nor U12885 (N_12885,N_12601,N_12518);
nand U12886 (N_12886,N_12690,N_12548);
nor U12887 (N_12887,N_12516,N_12550);
nand U12888 (N_12888,N_12562,N_12743);
nand U12889 (N_12889,N_12603,N_12725);
nand U12890 (N_12890,N_12709,N_12602);
xnor U12891 (N_12891,N_12571,N_12714);
and U12892 (N_12892,N_12664,N_12523);
xnor U12893 (N_12893,N_12712,N_12562);
and U12894 (N_12894,N_12733,N_12696);
nor U12895 (N_12895,N_12717,N_12613);
nand U12896 (N_12896,N_12548,N_12502);
and U12897 (N_12897,N_12684,N_12695);
nand U12898 (N_12898,N_12723,N_12577);
nor U12899 (N_12899,N_12740,N_12556);
nor U12900 (N_12900,N_12683,N_12544);
and U12901 (N_12901,N_12698,N_12662);
nand U12902 (N_12902,N_12514,N_12512);
and U12903 (N_12903,N_12624,N_12731);
or U12904 (N_12904,N_12572,N_12691);
nand U12905 (N_12905,N_12520,N_12649);
nor U12906 (N_12906,N_12695,N_12715);
xor U12907 (N_12907,N_12589,N_12630);
and U12908 (N_12908,N_12563,N_12556);
and U12909 (N_12909,N_12639,N_12745);
xnor U12910 (N_12910,N_12536,N_12706);
nand U12911 (N_12911,N_12583,N_12508);
nand U12912 (N_12912,N_12505,N_12654);
nand U12913 (N_12913,N_12576,N_12547);
nand U12914 (N_12914,N_12522,N_12693);
or U12915 (N_12915,N_12731,N_12724);
nand U12916 (N_12916,N_12706,N_12728);
or U12917 (N_12917,N_12644,N_12504);
and U12918 (N_12918,N_12746,N_12606);
or U12919 (N_12919,N_12652,N_12720);
nand U12920 (N_12920,N_12597,N_12639);
or U12921 (N_12921,N_12671,N_12707);
nand U12922 (N_12922,N_12685,N_12545);
xor U12923 (N_12923,N_12579,N_12644);
nand U12924 (N_12924,N_12578,N_12690);
nor U12925 (N_12925,N_12658,N_12573);
and U12926 (N_12926,N_12593,N_12628);
or U12927 (N_12927,N_12530,N_12511);
and U12928 (N_12928,N_12621,N_12500);
nor U12929 (N_12929,N_12651,N_12739);
nand U12930 (N_12930,N_12541,N_12730);
xnor U12931 (N_12931,N_12631,N_12713);
xor U12932 (N_12932,N_12619,N_12654);
and U12933 (N_12933,N_12699,N_12641);
nor U12934 (N_12934,N_12643,N_12713);
or U12935 (N_12935,N_12532,N_12709);
and U12936 (N_12936,N_12702,N_12528);
xor U12937 (N_12937,N_12704,N_12623);
xor U12938 (N_12938,N_12749,N_12732);
nand U12939 (N_12939,N_12737,N_12527);
and U12940 (N_12940,N_12707,N_12680);
nor U12941 (N_12941,N_12734,N_12589);
xnor U12942 (N_12942,N_12533,N_12623);
nor U12943 (N_12943,N_12553,N_12507);
and U12944 (N_12944,N_12654,N_12522);
xor U12945 (N_12945,N_12739,N_12748);
nand U12946 (N_12946,N_12551,N_12530);
nor U12947 (N_12947,N_12661,N_12617);
nand U12948 (N_12948,N_12644,N_12556);
nor U12949 (N_12949,N_12616,N_12596);
nor U12950 (N_12950,N_12577,N_12575);
or U12951 (N_12951,N_12744,N_12619);
nor U12952 (N_12952,N_12517,N_12649);
or U12953 (N_12953,N_12657,N_12574);
and U12954 (N_12954,N_12634,N_12722);
or U12955 (N_12955,N_12699,N_12620);
nand U12956 (N_12956,N_12655,N_12716);
and U12957 (N_12957,N_12749,N_12535);
nand U12958 (N_12958,N_12697,N_12549);
and U12959 (N_12959,N_12535,N_12632);
xnor U12960 (N_12960,N_12657,N_12572);
xor U12961 (N_12961,N_12705,N_12664);
or U12962 (N_12962,N_12506,N_12724);
xnor U12963 (N_12963,N_12710,N_12652);
xor U12964 (N_12964,N_12549,N_12715);
nand U12965 (N_12965,N_12528,N_12566);
nor U12966 (N_12966,N_12698,N_12583);
nor U12967 (N_12967,N_12622,N_12664);
nand U12968 (N_12968,N_12677,N_12524);
and U12969 (N_12969,N_12549,N_12726);
or U12970 (N_12970,N_12737,N_12698);
xor U12971 (N_12971,N_12550,N_12621);
nor U12972 (N_12972,N_12740,N_12572);
and U12973 (N_12973,N_12618,N_12506);
nand U12974 (N_12974,N_12619,N_12590);
xor U12975 (N_12975,N_12707,N_12704);
nand U12976 (N_12976,N_12533,N_12592);
or U12977 (N_12977,N_12566,N_12707);
xnor U12978 (N_12978,N_12716,N_12587);
or U12979 (N_12979,N_12643,N_12624);
or U12980 (N_12980,N_12684,N_12584);
xor U12981 (N_12981,N_12600,N_12516);
xnor U12982 (N_12982,N_12644,N_12695);
and U12983 (N_12983,N_12707,N_12551);
nor U12984 (N_12984,N_12709,N_12679);
or U12985 (N_12985,N_12610,N_12524);
nand U12986 (N_12986,N_12665,N_12523);
and U12987 (N_12987,N_12550,N_12691);
xor U12988 (N_12988,N_12623,N_12660);
or U12989 (N_12989,N_12665,N_12728);
and U12990 (N_12990,N_12624,N_12693);
and U12991 (N_12991,N_12529,N_12731);
nor U12992 (N_12992,N_12572,N_12532);
xnor U12993 (N_12993,N_12696,N_12600);
nand U12994 (N_12994,N_12692,N_12634);
nand U12995 (N_12995,N_12690,N_12531);
nand U12996 (N_12996,N_12736,N_12625);
xnor U12997 (N_12997,N_12682,N_12654);
or U12998 (N_12998,N_12660,N_12741);
nor U12999 (N_12999,N_12515,N_12518);
and U13000 (N_13000,N_12899,N_12767);
and U13001 (N_13001,N_12944,N_12960);
or U13002 (N_13002,N_12969,N_12973);
nor U13003 (N_13003,N_12917,N_12820);
xnor U13004 (N_13004,N_12979,N_12827);
nor U13005 (N_13005,N_12896,N_12774);
or U13006 (N_13006,N_12753,N_12766);
nor U13007 (N_13007,N_12872,N_12994);
and U13008 (N_13008,N_12888,N_12811);
and U13009 (N_13009,N_12808,N_12787);
or U13010 (N_13010,N_12963,N_12762);
nand U13011 (N_13011,N_12794,N_12932);
or U13012 (N_13012,N_12921,N_12952);
and U13013 (N_13013,N_12895,N_12892);
xor U13014 (N_13014,N_12912,N_12800);
and U13015 (N_13015,N_12783,N_12976);
and U13016 (N_13016,N_12769,N_12931);
nor U13017 (N_13017,N_12824,N_12990);
nor U13018 (N_13018,N_12862,N_12847);
xor U13019 (N_13019,N_12771,N_12941);
nand U13020 (N_13020,N_12873,N_12844);
nand U13021 (N_13021,N_12937,N_12821);
or U13022 (N_13022,N_12949,N_12750);
xnor U13023 (N_13023,N_12829,N_12825);
and U13024 (N_13024,N_12974,N_12793);
nand U13025 (N_13025,N_12876,N_12792);
or U13026 (N_13026,N_12845,N_12954);
nand U13027 (N_13027,N_12951,N_12871);
nand U13028 (N_13028,N_12853,N_12843);
nor U13029 (N_13029,N_12883,N_12848);
or U13030 (N_13030,N_12810,N_12865);
xnor U13031 (N_13031,N_12964,N_12867);
xor U13032 (N_13032,N_12923,N_12763);
xor U13033 (N_13033,N_12910,N_12849);
or U13034 (N_13034,N_12889,N_12989);
nor U13035 (N_13035,N_12885,N_12779);
and U13036 (N_13036,N_12880,N_12982);
and U13037 (N_13037,N_12893,N_12809);
nand U13038 (N_13038,N_12773,N_12958);
xnor U13039 (N_13039,N_12785,N_12799);
xor U13040 (N_13040,N_12760,N_12993);
xnor U13041 (N_13041,N_12992,N_12863);
nand U13042 (N_13042,N_12938,N_12985);
or U13043 (N_13043,N_12836,N_12978);
nand U13044 (N_13044,N_12852,N_12860);
and U13045 (N_13045,N_12838,N_12898);
or U13046 (N_13046,N_12846,N_12831);
xnor U13047 (N_13047,N_12916,N_12984);
and U13048 (N_13048,N_12789,N_12906);
and U13049 (N_13049,N_12981,N_12959);
nand U13050 (N_13050,N_12987,N_12828);
xor U13051 (N_13051,N_12911,N_12859);
and U13052 (N_13052,N_12814,N_12834);
nor U13053 (N_13053,N_12784,N_12822);
nand U13054 (N_13054,N_12928,N_12902);
nor U13055 (N_13055,N_12761,N_12936);
and U13056 (N_13056,N_12925,N_12919);
and U13057 (N_13057,N_12839,N_12926);
and U13058 (N_13058,N_12920,N_12890);
nor U13059 (N_13059,N_12886,N_12971);
nor U13060 (N_13060,N_12980,N_12939);
and U13061 (N_13061,N_12857,N_12874);
or U13062 (N_13062,N_12927,N_12875);
and U13063 (N_13063,N_12772,N_12877);
or U13064 (N_13064,N_12754,N_12805);
nand U13065 (N_13065,N_12757,N_12837);
xor U13066 (N_13066,N_12826,N_12751);
nor U13067 (N_13067,N_12943,N_12804);
or U13068 (N_13068,N_12861,N_12780);
nand U13069 (N_13069,N_12934,N_12997);
and U13070 (N_13070,N_12786,N_12796);
xnor U13071 (N_13071,N_12864,N_12965);
nor U13072 (N_13072,N_12866,N_12819);
xnor U13073 (N_13073,N_12942,N_12768);
nand U13074 (N_13074,N_12777,N_12882);
nand U13075 (N_13075,N_12798,N_12855);
or U13076 (N_13076,N_12781,N_12770);
nand U13077 (N_13077,N_12972,N_12991);
nand U13078 (N_13078,N_12986,N_12961);
and U13079 (N_13079,N_12817,N_12795);
nand U13080 (N_13080,N_12891,N_12908);
nand U13081 (N_13081,N_12816,N_12806);
nor U13082 (N_13082,N_12948,N_12881);
nand U13083 (N_13083,N_12775,N_12957);
or U13084 (N_13084,N_12778,N_12975);
xor U13085 (N_13085,N_12758,N_12842);
or U13086 (N_13086,N_12776,N_12884);
and U13087 (N_13087,N_12933,N_12915);
and U13088 (N_13088,N_12901,N_12790);
xnor U13089 (N_13089,N_12955,N_12956);
xnor U13090 (N_13090,N_12924,N_12946);
nor U13091 (N_13091,N_12900,N_12870);
xor U13092 (N_13092,N_12947,N_12835);
xnor U13093 (N_13093,N_12935,N_12998);
or U13094 (N_13094,N_12950,N_12940);
xor U13095 (N_13095,N_12996,N_12995);
or U13096 (N_13096,N_12851,N_12929);
xnor U13097 (N_13097,N_12759,N_12967);
xor U13098 (N_13098,N_12802,N_12755);
nor U13099 (N_13099,N_12858,N_12977);
nand U13100 (N_13100,N_12887,N_12752);
or U13101 (N_13101,N_12803,N_12823);
or U13102 (N_13102,N_12815,N_12854);
nor U13103 (N_13103,N_12764,N_12812);
and U13104 (N_13104,N_12894,N_12782);
and U13105 (N_13105,N_12807,N_12930);
nand U13106 (N_13106,N_12879,N_12797);
and U13107 (N_13107,N_12832,N_12869);
nor U13108 (N_13108,N_12756,N_12968);
and U13109 (N_13109,N_12918,N_12909);
nor U13110 (N_13110,N_12818,N_12914);
xor U13111 (N_13111,N_12856,N_12813);
nand U13112 (N_13112,N_12788,N_12907);
nand U13113 (N_13113,N_12988,N_12765);
nor U13114 (N_13114,N_12962,N_12966);
and U13115 (N_13115,N_12801,N_12913);
or U13116 (N_13116,N_12904,N_12833);
xor U13117 (N_13117,N_12878,N_12953);
nand U13118 (N_13118,N_12897,N_12840);
xor U13119 (N_13119,N_12999,N_12905);
nand U13120 (N_13120,N_12945,N_12850);
and U13121 (N_13121,N_12841,N_12970);
or U13122 (N_13122,N_12922,N_12868);
nor U13123 (N_13123,N_12791,N_12830);
and U13124 (N_13124,N_12983,N_12903);
and U13125 (N_13125,N_12808,N_12962);
and U13126 (N_13126,N_12881,N_12951);
or U13127 (N_13127,N_12780,N_12868);
nand U13128 (N_13128,N_12896,N_12824);
or U13129 (N_13129,N_12928,N_12967);
or U13130 (N_13130,N_12907,N_12789);
nor U13131 (N_13131,N_12969,N_12788);
nor U13132 (N_13132,N_12912,N_12949);
nand U13133 (N_13133,N_12986,N_12935);
xnor U13134 (N_13134,N_12930,N_12983);
and U13135 (N_13135,N_12795,N_12890);
nand U13136 (N_13136,N_12983,N_12954);
or U13137 (N_13137,N_12891,N_12775);
nand U13138 (N_13138,N_12761,N_12948);
and U13139 (N_13139,N_12940,N_12848);
nand U13140 (N_13140,N_12776,N_12790);
xor U13141 (N_13141,N_12789,N_12786);
nor U13142 (N_13142,N_12951,N_12872);
and U13143 (N_13143,N_12774,N_12825);
nor U13144 (N_13144,N_12824,N_12817);
xor U13145 (N_13145,N_12810,N_12921);
nand U13146 (N_13146,N_12854,N_12802);
or U13147 (N_13147,N_12907,N_12945);
xor U13148 (N_13148,N_12782,N_12937);
nand U13149 (N_13149,N_12894,N_12827);
or U13150 (N_13150,N_12801,N_12881);
nand U13151 (N_13151,N_12767,N_12788);
xnor U13152 (N_13152,N_12912,N_12838);
xnor U13153 (N_13153,N_12988,N_12933);
or U13154 (N_13154,N_12772,N_12848);
nand U13155 (N_13155,N_12762,N_12996);
or U13156 (N_13156,N_12909,N_12766);
and U13157 (N_13157,N_12831,N_12823);
or U13158 (N_13158,N_12795,N_12841);
and U13159 (N_13159,N_12976,N_12789);
and U13160 (N_13160,N_12909,N_12959);
and U13161 (N_13161,N_12817,N_12894);
nand U13162 (N_13162,N_12754,N_12993);
and U13163 (N_13163,N_12824,N_12889);
or U13164 (N_13164,N_12889,N_12941);
nor U13165 (N_13165,N_12810,N_12766);
xnor U13166 (N_13166,N_12904,N_12886);
and U13167 (N_13167,N_12990,N_12883);
xnor U13168 (N_13168,N_12972,N_12911);
xnor U13169 (N_13169,N_12985,N_12767);
and U13170 (N_13170,N_12822,N_12880);
and U13171 (N_13171,N_12753,N_12992);
xor U13172 (N_13172,N_12985,N_12826);
or U13173 (N_13173,N_12871,N_12961);
or U13174 (N_13174,N_12859,N_12980);
or U13175 (N_13175,N_12976,N_12843);
nand U13176 (N_13176,N_12974,N_12924);
and U13177 (N_13177,N_12981,N_12926);
xor U13178 (N_13178,N_12819,N_12844);
or U13179 (N_13179,N_12988,N_12795);
nand U13180 (N_13180,N_12840,N_12760);
nor U13181 (N_13181,N_12953,N_12814);
xor U13182 (N_13182,N_12970,N_12792);
nor U13183 (N_13183,N_12995,N_12959);
nor U13184 (N_13184,N_12897,N_12958);
or U13185 (N_13185,N_12937,N_12867);
xnor U13186 (N_13186,N_12934,N_12974);
xnor U13187 (N_13187,N_12820,N_12756);
and U13188 (N_13188,N_12790,N_12802);
nand U13189 (N_13189,N_12863,N_12970);
or U13190 (N_13190,N_12965,N_12973);
nor U13191 (N_13191,N_12904,N_12841);
nor U13192 (N_13192,N_12973,N_12832);
or U13193 (N_13193,N_12936,N_12871);
and U13194 (N_13194,N_12755,N_12768);
and U13195 (N_13195,N_12908,N_12816);
xnor U13196 (N_13196,N_12878,N_12916);
and U13197 (N_13197,N_12782,N_12870);
nand U13198 (N_13198,N_12884,N_12995);
or U13199 (N_13199,N_12893,N_12890);
nor U13200 (N_13200,N_12873,N_12758);
nor U13201 (N_13201,N_12850,N_12950);
xnor U13202 (N_13202,N_12985,N_12817);
nand U13203 (N_13203,N_12761,N_12885);
and U13204 (N_13204,N_12857,N_12933);
xor U13205 (N_13205,N_12823,N_12903);
and U13206 (N_13206,N_12831,N_12849);
nand U13207 (N_13207,N_12767,N_12902);
nor U13208 (N_13208,N_12987,N_12827);
and U13209 (N_13209,N_12990,N_12874);
xnor U13210 (N_13210,N_12996,N_12932);
or U13211 (N_13211,N_12779,N_12911);
xor U13212 (N_13212,N_12989,N_12829);
nor U13213 (N_13213,N_12892,N_12761);
and U13214 (N_13214,N_12797,N_12989);
nand U13215 (N_13215,N_12962,N_12852);
xnor U13216 (N_13216,N_12981,N_12826);
xor U13217 (N_13217,N_12834,N_12843);
or U13218 (N_13218,N_12794,N_12956);
nand U13219 (N_13219,N_12860,N_12936);
xor U13220 (N_13220,N_12871,N_12790);
and U13221 (N_13221,N_12916,N_12816);
xnor U13222 (N_13222,N_12814,N_12973);
xor U13223 (N_13223,N_12988,N_12846);
xor U13224 (N_13224,N_12995,N_12781);
nand U13225 (N_13225,N_12945,N_12957);
or U13226 (N_13226,N_12984,N_12850);
or U13227 (N_13227,N_12777,N_12773);
and U13228 (N_13228,N_12765,N_12904);
xor U13229 (N_13229,N_12784,N_12802);
xnor U13230 (N_13230,N_12780,N_12750);
nor U13231 (N_13231,N_12845,N_12873);
or U13232 (N_13232,N_12928,N_12942);
nor U13233 (N_13233,N_12850,N_12915);
and U13234 (N_13234,N_12995,N_12811);
xnor U13235 (N_13235,N_12761,N_12845);
nor U13236 (N_13236,N_12818,N_12752);
nand U13237 (N_13237,N_12923,N_12838);
nor U13238 (N_13238,N_12855,N_12891);
and U13239 (N_13239,N_12851,N_12996);
xnor U13240 (N_13240,N_12946,N_12846);
xnor U13241 (N_13241,N_12870,N_12924);
and U13242 (N_13242,N_12952,N_12898);
and U13243 (N_13243,N_12833,N_12758);
and U13244 (N_13244,N_12985,N_12928);
nor U13245 (N_13245,N_12820,N_12751);
xnor U13246 (N_13246,N_12980,N_12763);
and U13247 (N_13247,N_12892,N_12987);
and U13248 (N_13248,N_12805,N_12794);
xnor U13249 (N_13249,N_12938,N_12829);
and U13250 (N_13250,N_13127,N_13015);
or U13251 (N_13251,N_13000,N_13007);
and U13252 (N_13252,N_13196,N_13123);
nor U13253 (N_13253,N_13245,N_13072);
nand U13254 (N_13254,N_13162,N_13030);
and U13255 (N_13255,N_13068,N_13141);
nor U13256 (N_13256,N_13097,N_13192);
and U13257 (N_13257,N_13101,N_13046);
and U13258 (N_13258,N_13045,N_13213);
nor U13259 (N_13259,N_13246,N_13109);
xnor U13260 (N_13260,N_13049,N_13048);
nand U13261 (N_13261,N_13009,N_13057);
and U13262 (N_13262,N_13023,N_13063);
xor U13263 (N_13263,N_13047,N_13020);
or U13264 (N_13264,N_13170,N_13155);
nor U13265 (N_13265,N_13175,N_13178);
xnor U13266 (N_13266,N_13035,N_13111);
and U13267 (N_13267,N_13104,N_13247);
nor U13268 (N_13268,N_13147,N_13157);
and U13269 (N_13269,N_13086,N_13113);
xor U13270 (N_13270,N_13146,N_13185);
nand U13271 (N_13271,N_13103,N_13166);
and U13272 (N_13272,N_13164,N_13210);
xnor U13273 (N_13273,N_13143,N_13168);
nor U13274 (N_13274,N_13225,N_13087);
or U13275 (N_13275,N_13114,N_13126);
or U13276 (N_13276,N_13004,N_13177);
or U13277 (N_13277,N_13074,N_13226);
and U13278 (N_13278,N_13021,N_13052);
nand U13279 (N_13279,N_13037,N_13218);
nand U13280 (N_13280,N_13050,N_13120);
nor U13281 (N_13281,N_13236,N_13172);
xnor U13282 (N_13282,N_13038,N_13212);
xor U13283 (N_13283,N_13179,N_13040);
nor U13284 (N_13284,N_13209,N_13075);
nand U13285 (N_13285,N_13190,N_13200);
nand U13286 (N_13286,N_13204,N_13081);
or U13287 (N_13287,N_13221,N_13159);
xor U13288 (N_13288,N_13151,N_13026);
and U13289 (N_13289,N_13059,N_13202);
xor U13290 (N_13290,N_13248,N_13090);
or U13291 (N_13291,N_13088,N_13025);
or U13292 (N_13292,N_13224,N_13003);
nand U13293 (N_13293,N_13148,N_13056);
and U13294 (N_13294,N_13098,N_13060);
nor U13295 (N_13295,N_13118,N_13034);
nand U13296 (N_13296,N_13085,N_13082);
and U13297 (N_13297,N_13054,N_13238);
or U13298 (N_13298,N_13154,N_13217);
and U13299 (N_13299,N_13091,N_13241);
xnor U13300 (N_13300,N_13207,N_13029);
nor U13301 (N_13301,N_13051,N_13061);
nor U13302 (N_13302,N_13231,N_13152);
or U13303 (N_13303,N_13189,N_13138);
xnor U13304 (N_13304,N_13070,N_13084);
xor U13305 (N_13305,N_13187,N_13032);
and U13306 (N_13306,N_13211,N_13073);
nor U13307 (N_13307,N_13095,N_13058);
or U13308 (N_13308,N_13115,N_13121);
xnor U13309 (N_13309,N_13077,N_13130);
and U13310 (N_13310,N_13180,N_13197);
or U13311 (N_13311,N_13112,N_13235);
and U13312 (N_13312,N_13001,N_13229);
or U13313 (N_13313,N_13156,N_13124);
xnor U13314 (N_13314,N_13027,N_13243);
xnor U13315 (N_13315,N_13198,N_13216);
nand U13316 (N_13316,N_13160,N_13233);
nor U13317 (N_13317,N_13105,N_13071);
nand U13318 (N_13318,N_13214,N_13008);
and U13319 (N_13319,N_13065,N_13167);
and U13320 (N_13320,N_13080,N_13145);
and U13321 (N_13321,N_13223,N_13099);
and U13322 (N_13322,N_13219,N_13036);
or U13323 (N_13323,N_13244,N_13092);
nor U13324 (N_13324,N_13079,N_13017);
or U13325 (N_13325,N_13139,N_13110);
nor U13326 (N_13326,N_13066,N_13067);
nor U13327 (N_13327,N_13194,N_13031);
xnor U13328 (N_13328,N_13011,N_13016);
or U13329 (N_13329,N_13150,N_13106);
and U13330 (N_13330,N_13227,N_13002);
or U13331 (N_13331,N_13078,N_13005);
nor U13332 (N_13332,N_13128,N_13117);
nand U13333 (N_13333,N_13094,N_13135);
and U13334 (N_13334,N_13239,N_13134);
nand U13335 (N_13335,N_13100,N_13222);
or U13336 (N_13336,N_13028,N_13228);
nand U13337 (N_13337,N_13206,N_13195);
or U13338 (N_13338,N_13230,N_13184);
xor U13339 (N_13339,N_13220,N_13234);
or U13340 (N_13340,N_13215,N_13116);
xnor U13341 (N_13341,N_13242,N_13186);
or U13342 (N_13342,N_13171,N_13125);
nor U13343 (N_13343,N_13208,N_13169);
and U13344 (N_13344,N_13193,N_13142);
nor U13345 (N_13345,N_13153,N_13108);
and U13346 (N_13346,N_13022,N_13044);
or U13347 (N_13347,N_13181,N_13237);
and U13348 (N_13348,N_13102,N_13201);
and U13349 (N_13349,N_13119,N_13174);
nand U13350 (N_13350,N_13137,N_13240);
nand U13351 (N_13351,N_13024,N_13182);
or U13352 (N_13352,N_13191,N_13203);
and U13353 (N_13353,N_13232,N_13033);
nor U13354 (N_13354,N_13129,N_13062);
nand U13355 (N_13355,N_13053,N_13183);
nor U13356 (N_13356,N_13133,N_13122);
xor U13357 (N_13357,N_13014,N_13149);
nor U13358 (N_13358,N_13136,N_13188);
and U13359 (N_13359,N_13093,N_13043);
nand U13360 (N_13360,N_13205,N_13089);
and U13361 (N_13361,N_13165,N_13096);
or U13362 (N_13362,N_13163,N_13083);
xor U13363 (N_13363,N_13041,N_13144);
nor U13364 (N_13364,N_13076,N_13176);
or U13365 (N_13365,N_13131,N_13132);
xor U13366 (N_13366,N_13249,N_13006);
or U13367 (N_13367,N_13019,N_13012);
xnor U13368 (N_13368,N_13107,N_13039);
or U13369 (N_13369,N_13010,N_13161);
and U13370 (N_13370,N_13173,N_13140);
xor U13371 (N_13371,N_13013,N_13042);
nor U13372 (N_13372,N_13158,N_13064);
and U13373 (N_13373,N_13018,N_13069);
and U13374 (N_13374,N_13055,N_13199);
nand U13375 (N_13375,N_13006,N_13152);
nor U13376 (N_13376,N_13015,N_13249);
xor U13377 (N_13377,N_13164,N_13056);
or U13378 (N_13378,N_13108,N_13086);
nor U13379 (N_13379,N_13100,N_13174);
nand U13380 (N_13380,N_13249,N_13101);
nor U13381 (N_13381,N_13213,N_13218);
and U13382 (N_13382,N_13216,N_13142);
nand U13383 (N_13383,N_13166,N_13101);
and U13384 (N_13384,N_13109,N_13214);
nor U13385 (N_13385,N_13221,N_13220);
nor U13386 (N_13386,N_13159,N_13128);
nand U13387 (N_13387,N_13097,N_13128);
xnor U13388 (N_13388,N_13143,N_13228);
or U13389 (N_13389,N_13132,N_13207);
nand U13390 (N_13390,N_13222,N_13018);
xor U13391 (N_13391,N_13047,N_13220);
nor U13392 (N_13392,N_13024,N_13071);
or U13393 (N_13393,N_13021,N_13039);
xor U13394 (N_13394,N_13204,N_13031);
xnor U13395 (N_13395,N_13170,N_13166);
or U13396 (N_13396,N_13038,N_13143);
nor U13397 (N_13397,N_13228,N_13201);
or U13398 (N_13398,N_13081,N_13134);
nor U13399 (N_13399,N_13042,N_13186);
or U13400 (N_13400,N_13203,N_13132);
xnor U13401 (N_13401,N_13193,N_13188);
nand U13402 (N_13402,N_13208,N_13111);
or U13403 (N_13403,N_13084,N_13247);
nand U13404 (N_13404,N_13173,N_13003);
or U13405 (N_13405,N_13169,N_13073);
nor U13406 (N_13406,N_13163,N_13146);
nor U13407 (N_13407,N_13099,N_13207);
nor U13408 (N_13408,N_13012,N_13000);
or U13409 (N_13409,N_13214,N_13077);
and U13410 (N_13410,N_13205,N_13122);
nor U13411 (N_13411,N_13202,N_13053);
or U13412 (N_13412,N_13141,N_13043);
nor U13413 (N_13413,N_13138,N_13225);
or U13414 (N_13414,N_13151,N_13238);
nand U13415 (N_13415,N_13238,N_13227);
or U13416 (N_13416,N_13005,N_13019);
nor U13417 (N_13417,N_13001,N_13236);
or U13418 (N_13418,N_13027,N_13128);
nor U13419 (N_13419,N_13232,N_13212);
nor U13420 (N_13420,N_13136,N_13038);
nand U13421 (N_13421,N_13026,N_13073);
and U13422 (N_13422,N_13023,N_13083);
nor U13423 (N_13423,N_13062,N_13221);
nor U13424 (N_13424,N_13218,N_13025);
nand U13425 (N_13425,N_13174,N_13086);
nor U13426 (N_13426,N_13236,N_13202);
or U13427 (N_13427,N_13083,N_13116);
and U13428 (N_13428,N_13193,N_13246);
or U13429 (N_13429,N_13244,N_13032);
or U13430 (N_13430,N_13105,N_13197);
or U13431 (N_13431,N_13010,N_13231);
or U13432 (N_13432,N_13057,N_13092);
or U13433 (N_13433,N_13110,N_13032);
or U13434 (N_13434,N_13057,N_13190);
xnor U13435 (N_13435,N_13066,N_13233);
nor U13436 (N_13436,N_13116,N_13204);
xor U13437 (N_13437,N_13123,N_13148);
or U13438 (N_13438,N_13104,N_13059);
nor U13439 (N_13439,N_13216,N_13015);
xnor U13440 (N_13440,N_13082,N_13152);
xor U13441 (N_13441,N_13037,N_13072);
nor U13442 (N_13442,N_13089,N_13109);
nand U13443 (N_13443,N_13141,N_13087);
nand U13444 (N_13444,N_13032,N_13106);
nor U13445 (N_13445,N_13022,N_13133);
and U13446 (N_13446,N_13036,N_13162);
nor U13447 (N_13447,N_13235,N_13073);
or U13448 (N_13448,N_13051,N_13214);
or U13449 (N_13449,N_13225,N_13240);
or U13450 (N_13450,N_13070,N_13111);
nand U13451 (N_13451,N_13013,N_13066);
nand U13452 (N_13452,N_13058,N_13024);
nand U13453 (N_13453,N_13228,N_13029);
or U13454 (N_13454,N_13004,N_13022);
nor U13455 (N_13455,N_13163,N_13110);
xnor U13456 (N_13456,N_13069,N_13151);
and U13457 (N_13457,N_13127,N_13156);
and U13458 (N_13458,N_13185,N_13246);
nand U13459 (N_13459,N_13189,N_13210);
nor U13460 (N_13460,N_13029,N_13023);
xor U13461 (N_13461,N_13079,N_13032);
and U13462 (N_13462,N_13206,N_13003);
nand U13463 (N_13463,N_13138,N_13200);
nor U13464 (N_13464,N_13143,N_13151);
or U13465 (N_13465,N_13050,N_13037);
or U13466 (N_13466,N_13066,N_13080);
and U13467 (N_13467,N_13018,N_13148);
xnor U13468 (N_13468,N_13205,N_13078);
nand U13469 (N_13469,N_13225,N_13019);
nand U13470 (N_13470,N_13119,N_13193);
and U13471 (N_13471,N_13015,N_13245);
or U13472 (N_13472,N_13187,N_13107);
or U13473 (N_13473,N_13039,N_13106);
or U13474 (N_13474,N_13208,N_13237);
and U13475 (N_13475,N_13224,N_13228);
or U13476 (N_13476,N_13167,N_13021);
and U13477 (N_13477,N_13110,N_13042);
and U13478 (N_13478,N_13219,N_13189);
and U13479 (N_13479,N_13179,N_13132);
and U13480 (N_13480,N_13100,N_13159);
or U13481 (N_13481,N_13016,N_13208);
xor U13482 (N_13482,N_13059,N_13097);
or U13483 (N_13483,N_13104,N_13204);
and U13484 (N_13484,N_13077,N_13026);
xor U13485 (N_13485,N_13208,N_13198);
or U13486 (N_13486,N_13210,N_13198);
and U13487 (N_13487,N_13197,N_13044);
nor U13488 (N_13488,N_13127,N_13231);
nor U13489 (N_13489,N_13192,N_13090);
or U13490 (N_13490,N_13069,N_13114);
xor U13491 (N_13491,N_13174,N_13149);
and U13492 (N_13492,N_13162,N_13091);
or U13493 (N_13493,N_13179,N_13199);
nand U13494 (N_13494,N_13006,N_13085);
or U13495 (N_13495,N_13189,N_13103);
nand U13496 (N_13496,N_13027,N_13083);
and U13497 (N_13497,N_13142,N_13153);
xnor U13498 (N_13498,N_13071,N_13097);
nor U13499 (N_13499,N_13134,N_13005);
xnor U13500 (N_13500,N_13396,N_13306);
nand U13501 (N_13501,N_13361,N_13337);
or U13502 (N_13502,N_13491,N_13354);
nor U13503 (N_13503,N_13283,N_13429);
nand U13504 (N_13504,N_13428,N_13277);
xnor U13505 (N_13505,N_13390,N_13316);
xor U13506 (N_13506,N_13297,N_13320);
xnor U13507 (N_13507,N_13397,N_13372);
nand U13508 (N_13508,N_13353,N_13492);
and U13509 (N_13509,N_13444,N_13462);
nor U13510 (N_13510,N_13410,N_13252);
xor U13511 (N_13511,N_13255,N_13323);
nand U13512 (N_13512,N_13286,N_13383);
xnor U13513 (N_13513,N_13424,N_13394);
or U13514 (N_13514,N_13425,N_13478);
xor U13515 (N_13515,N_13261,N_13395);
nor U13516 (N_13516,N_13370,N_13452);
and U13517 (N_13517,N_13262,N_13284);
nor U13518 (N_13518,N_13307,N_13263);
xnor U13519 (N_13519,N_13343,N_13391);
and U13520 (N_13520,N_13359,N_13419);
or U13521 (N_13521,N_13449,N_13331);
xnor U13522 (N_13522,N_13380,N_13399);
and U13523 (N_13523,N_13374,N_13371);
xnor U13524 (N_13524,N_13467,N_13430);
or U13525 (N_13525,N_13426,N_13456);
nor U13526 (N_13526,N_13292,N_13474);
nand U13527 (N_13527,N_13421,N_13363);
nor U13528 (N_13528,N_13433,N_13404);
xnor U13529 (N_13529,N_13260,N_13466);
or U13530 (N_13530,N_13345,N_13258);
and U13531 (N_13531,N_13443,N_13402);
or U13532 (N_13532,N_13480,N_13392);
xor U13533 (N_13533,N_13493,N_13386);
xnor U13534 (N_13534,N_13308,N_13324);
nor U13535 (N_13535,N_13264,N_13287);
and U13536 (N_13536,N_13436,N_13275);
or U13537 (N_13537,N_13470,N_13440);
and U13538 (N_13538,N_13267,N_13319);
nand U13539 (N_13539,N_13398,N_13407);
and U13540 (N_13540,N_13486,N_13327);
nand U13541 (N_13541,N_13375,N_13273);
nor U13542 (N_13542,N_13259,N_13439);
nand U13543 (N_13543,N_13411,N_13322);
or U13544 (N_13544,N_13301,N_13459);
or U13545 (N_13545,N_13473,N_13373);
nor U13546 (N_13546,N_13333,N_13329);
and U13547 (N_13547,N_13342,N_13355);
xor U13548 (N_13548,N_13257,N_13278);
nand U13549 (N_13549,N_13290,N_13321);
xnor U13550 (N_13550,N_13457,N_13418);
nor U13551 (N_13551,N_13420,N_13289);
and U13552 (N_13552,N_13282,N_13483);
nand U13553 (N_13553,N_13281,N_13296);
nor U13554 (N_13554,N_13406,N_13305);
nor U13555 (N_13555,N_13347,N_13250);
nand U13556 (N_13556,N_13340,N_13310);
and U13557 (N_13557,N_13285,N_13268);
nand U13558 (N_13558,N_13415,N_13294);
or U13559 (N_13559,N_13379,N_13302);
xor U13560 (N_13560,N_13385,N_13271);
nor U13561 (N_13561,N_13405,N_13460);
and U13562 (N_13562,N_13485,N_13311);
nor U13563 (N_13563,N_13299,N_13477);
or U13564 (N_13564,N_13272,N_13269);
nor U13565 (N_13565,N_13481,N_13414);
and U13566 (N_13566,N_13368,N_13352);
nand U13567 (N_13567,N_13441,N_13387);
nand U13568 (N_13568,N_13495,N_13427);
xor U13569 (N_13569,N_13463,N_13408);
or U13570 (N_13570,N_13348,N_13498);
xor U13571 (N_13571,N_13434,N_13300);
xnor U13572 (N_13572,N_13499,N_13376);
or U13573 (N_13573,N_13446,N_13482);
xnor U13574 (N_13574,N_13304,N_13265);
xnor U13575 (N_13575,N_13490,N_13280);
and U13576 (N_13576,N_13295,N_13403);
nor U13577 (N_13577,N_13458,N_13339);
xnor U13578 (N_13578,N_13369,N_13266);
or U13579 (N_13579,N_13346,N_13438);
nand U13580 (N_13580,N_13251,N_13479);
nor U13581 (N_13581,N_13488,N_13309);
and U13582 (N_13582,N_13365,N_13489);
nand U13583 (N_13583,N_13344,N_13471);
xor U13584 (N_13584,N_13432,N_13437);
and U13585 (N_13585,N_13475,N_13461);
and U13586 (N_13586,N_13313,N_13253);
nand U13587 (N_13587,N_13377,N_13445);
or U13588 (N_13588,N_13312,N_13468);
xnor U13589 (N_13589,N_13412,N_13279);
nor U13590 (N_13590,N_13315,N_13356);
nand U13591 (N_13591,N_13447,N_13350);
or U13592 (N_13592,N_13448,N_13497);
nand U13593 (N_13593,N_13317,N_13256);
or U13594 (N_13594,N_13384,N_13274);
and U13595 (N_13595,N_13455,N_13453);
nand U13596 (N_13596,N_13476,N_13341);
nand U13597 (N_13597,N_13435,N_13417);
nand U13598 (N_13598,N_13298,N_13442);
and U13599 (N_13599,N_13484,N_13325);
or U13600 (N_13600,N_13338,N_13293);
and U13601 (N_13601,N_13328,N_13332);
or U13602 (N_13602,N_13364,N_13270);
and U13603 (N_13603,N_13276,N_13303);
and U13604 (N_13604,N_13381,N_13351);
xnor U13605 (N_13605,N_13422,N_13413);
nand U13606 (N_13606,N_13423,N_13291);
nand U13607 (N_13607,N_13472,N_13431);
nor U13608 (N_13608,N_13378,N_13454);
nor U13609 (N_13609,N_13366,N_13335);
or U13610 (N_13610,N_13393,N_13416);
and U13611 (N_13611,N_13465,N_13357);
or U13612 (N_13612,N_13349,N_13288);
nand U13613 (N_13613,N_13469,N_13334);
xnor U13614 (N_13614,N_13336,N_13464);
or U13615 (N_13615,N_13367,N_13451);
or U13616 (N_13616,N_13314,N_13326);
nand U13617 (N_13617,N_13496,N_13400);
xnor U13618 (N_13618,N_13450,N_13494);
nand U13619 (N_13619,N_13389,N_13318);
or U13620 (N_13620,N_13360,N_13388);
and U13621 (N_13621,N_13358,N_13254);
or U13622 (N_13622,N_13330,N_13487);
and U13623 (N_13623,N_13409,N_13382);
nor U13624 (N_13624,N_13401,N_13362);
and U13625 (N_13625,N_13359,N_13353);
xor U13626 (N_13626,N_13315,N_13461);
or U13627 (N_13627,N_13439,N_13268);
nand U13628 (N_13628,N_13269,N_13404);
nand U13629 (N_13629,N_13347,N_13294);
or U13630 (N_13630,N_13336,N_13356);
and U13631 (N_13631,N_13296,N_13275);
and U13632 (N_13632,N_13425,N_13484);
and U13633 (N_13633,N_13320,N_13318);
or U13634 (N_13634,N_13436,N_13366);
nand U13635 (N_13635,N_13345,N_13396);
nand U13636 (N_13636,N_13392,N_13431);
nor U13637 (N_13637,N_13436,N_13359);
xnor U13638 (N_13638,N_13259,N_13452);
nand U13639 (N_13639,N_13352,N_13311);
nor U13640 (N_13640,N_13473,N_13322);
and U13641 (N_13641,N_13492,N_13493);
or U13642 (N_13642,N_13481,N_13408);
and U13643 (N_13643,N_13281,N_13341);
nand U13644 (N_13644,N_13496,N_13265);
nand U13645 (N_13645,N_13253,N_13319);
nor U13646 (N_13646,N_13444,N_13376);
xnor U13647 (N_13647,N_13288,N_13443);
or U13648 (N_13648,N_13374,N_13268);
xnor U13649 (N_13649,N_13464,N_13393);
nand U13650 (N_13650,N_13499,N_13440);
or U13651 (N_13651,N_13380,N_13261);
and U13652 (N_13652,N_13398,N_13406);
xnor U13653 (N_13653,N_13318,N_13280);
or U13654 (N_13654,N_13378,N_13325);
xor U13655 (N_13655,N_13373,N_13310);
nand U13656 (N_13656,N_13497,N_13418);
nand U13657 (N_13657,N_13345,N_13428);
and U13658 (N_13658,N_13286,N_13334);
xor U13659 (N_13659,N_13287,N_13464);
xnor U13660 (N_13660,N_13420,N_13460);
nand U13661 (N_13661,N_13269,N_13344);
xnor U13662 (N_13662,N_13456,N_13431);
nor U13663 (N_13663,N_13276,N_13389);
xnor U13664 (N_13664,N_13418,N_13486);
nor U13665 (N_13665,N_13363,N_13366);
xor U13666 (N_13666,N_13432,N_13448);
nor U13667 (N_13667,N_13499,N_13404);
and U13668 (N_13668,N_13281,N_13485);
and U13669 (N_13669,N_13491,N_13456);
nand U13670 (N_13670,N_13372,N_13444);
or U13671 (N_13671,N_13338,N_13350);
or U13672 (N_13672,N_13326,N_13373);
and U13673 (N_13673,N_13329,N_13421);
nand U13674 (N_13674,N_13434,N_13448);
nor U13675 (N_13675,N_13266,N_13413);
nand U13676 (N_13676,N_13321,N_13372);
and U13677 (N_13677,N_13310,N_13261);
xnor U13678 (N_13678,N_13296,N_13361);
or U13679 (N_13679,N_13480,N_13488);
nand U13680 (N_13680,N_13491,N_13274);
xnor U13681 (N_13681,N_13305,N_13457);
and U13682 (N_13682,N_13394,N_13294);
nand U13683 (N_13683,N_13255,N_13410);
nor U13684 (N_13684,N_13480,N_13404);
and U13685 (N_13685,N_13427,N_13270);
or U13686 (N_13686,N_13387,N_13358);
xnor U13687 (N_13687,N_13321,N_13320);
nand U13688 (N_13688,N_13426,N_13292);
or U13689 (N_13689,N_13461,N_13259);
xor U13690 (N_13690,N_13360,N_13410);
or U13691 (N_13691,N_13492,N_13337);
nor U13692 (N_13692,N_13282,N_13313);
or U13693 (N_13693,N_13417,N_13328);
xnor U13694 (N_13694,N_13402,N_13484);
or U13695 (N_13695,N_13265,N_13488);
or U13696 (N_13696,N_13307,N_13414);
xor U13697 (N_13697,N_13371,N_13385);
xor U13698 (N_13698,N_13271,N_13342);
nand U13699 (N_13699,N_13290,N_13365);
and U13700 (N_13700,N_13376,N_13358);
and U13701 (N_13701,N_13327,N_13406);
nand U13702 (N_13702,N_13440,N_13253);
xor U13703 (N_13703,N_13490,N_13299);
nand U13704 (N_13704,N_13498,N_13480);
nand U13705 (N_13705,N_13286,N_13325);
and U13706 (N_13706,N_13266,N_13330);
or U13707 (N_13707,N_13360,N_13496);
nand U13708 (N_13708,N_13268,N_13391);
or U13709 (N_13709,N_13317,N_13390);
nand U13710 (N_13710,N_13494,N_13417);
and U13711 (N_13711,N_13384,N_13441);
or U13712 (N_13712,N_13467,N_13421);
or U13713 (N_13713,N_13331,N_13301);
and U13714 (N_13714,N_13480,N_13368);
nor U13715 (N_13715,N_13409,N_13430);
xnor U13716 (N_13716,N_13406,N_13291);
xnor U13717 (N_13717,N_13370,N_13330);
or U13718 (N_13718,N_13380,N_13492);
or U13719 (N_13719,N_13458,N_13449);
xnor U13720 (N_13720,N_13292,N_13304);
or U13721 (N_13721,N_13487,N_13306);
nand U13722 (N_13722,N_13491,N_13359);
nand U13723 (N_13723,N_13497,N_13433);
nand U13724 (N_13724,N_13492,N_13261);
and U13725 (N_13725,N_13314,N_13472);
nor U13726 (N_13726,N_13325,N_13275);
xnor U13727 (N_13727,N_13400,N_13264);
nor U13728 (N_13728,N_13427,N_13284);
nor U13729 (N_13729,N_13421,N_13480);
nor U13730 (N_13730,N_13347,N_13422);
nand U13731 (N_13731,N_13497,N_13446);
and U13732 (N_13732,N_13480,N_13315);
xnor U13733 (N_13733,N_13281,N_13278);
nor U13734 (N_13734,N_13298,N_13425);
and U13735 (N_13735,N_13281,N_13471);
nor U13736 (N_13736,N_13265,N_13277);
nand U13737 (N_13737,N_13389,N_13373);
or U13738 (N_13738,N_13346,N_13256);
nand U13739 (N_13739,N_13460,N_13471);
nand U13740 (N_13740,N_13287,N_13331);
nor U13741 (N_13741,N_13413,N_13339);
nor U13742 (N_13742,N_13427,N_13438);
nand U13743 (N_13743,N_13469,N_13478);
nor U13744 (N_13744,N_13490,N_13312);
and U13745 (N_13745,N_13334,N_13456);
and U13746 (N_13746,N_13494,N_13352);
and U13747 (N_13747,N_13483,N_13485);
xor U13748 (N_13748,N_13334,N_13268);
or U13749 (N_13749,N_13276,N_13488);
nor U13750 (N_13750,N_13637,N_13703);
xnor U13751 (N_13751,N_13610,N_13615);
and U13752 (N_13752,N_13706,N_13577);
xnor U13753 (N_13753,N_13551,N_13733);
xnor U13754 (N_13754,N_13604,N_13679);
nor U13755 (N_13755,N_13509,N_13609);
nand U13756 (N_13756,N_13727,N_13522);
nor U13757 (N_13757,N_13695,N_13670);
xor U13758 (N_13758,N_13647,N_13666);
nor U13759 (N_13759,N_13598,N_13606);
and U13760 (N_13760,N_13541,N_13576);
nand U13761 (N_13761,N_13511,N_13704);
or U13762 (N_13762,N_13619,N_13537);
nor U13763 (N_13763,N_13588,N_13543);
nand U13764 (N_13764,N_13585,N_13746);
or U13765 (N_13765,N_13716,N_13651);
nand U13766 (N_13766,N_13687,N_13594);
nor U13767 (N_13767,N_13641,N_13663);
or U13768 (N_13768,N_13745,N_13611);
xor U13769 (N_13769,N_13653,N_13701);
nor U13770 (N_13770,N_13558,N_13623);
xor U13771 (N_13771,N_13530,N_13724);
nor U13772 (N_13772,N_13532,N_13742);
or U13773 (N_13773,N_13692,N_13673);
nor U13774 (N_13774,N_13529,N_13738);
nand U13775 (N_13775,N_13633,N_13593);
xor U13776 (N_13776,N_13741,N_13731);
and U13777 (N_13777,N_13707,N_13563);
and U13778 (N_13778,N_13675,N_13603);
nor U13779 (N_13779,N_13646,N_13693);
xor U13780 (N_13780,N_13586,N_13559);
xor U13781 (N_13781,N_13721,N_13565);
or U13782 (N_13782,N_13574,N_13717);
xnor U13783 (N_13783,N_13722,N_13730);
and U13784 (N_13784,N_13699,N_13566);
xor U13785 (N_13785,N_13664,N_13591);
nor U13786 (N_13786,N_13632,N_13728);
or U13787 (N_13787,N_13694,N_13729);
nor U13788 (N_13788,N_13640,N_13749);
nor U13789 (N_13789,N_13688,N_13554);
or U13790 (N_13790,N_13630,N_13639);
nor U13791 (N_13791,N_13700,N_13674);
nor U13792 (N_13792,N_13726,N_13601);
or U13793 (N_13793,N_13711,N_13582);
nor U13794 (N_13794,N_13581,N_13518);
nor U13795 (N_13795,N_13605,N_13523);
nand U13796 (N_13796,N_13564,N_13549);
xor U13797 (N_13797,N_13526,N_13502);
nor U13798 (N_13798,N_13571,N_13506);
or U13799 (N_13799,N_13712,N_13578);
or U13800 (N_13800,N_13686,N_13548);
nand U13801 (N_13801,N_13744,N_13710);
nand U13802 (N_13802,N_13597,N_13608);
and U13803 (N_13803,N_13570,N_13685);
nand U13804 (N_13804,N_13595,N_13552);
xnor U13805 (N_13805,N_13535,N_13650);
nor U13806 (N_13806,N_13725,N_13555);
and U13807 (N_13807,N_13705,N_13544);
and U13808 (N_13808,N_13508,N_13553);
nand U13809 (N_13809,N_13550,N_13561);
or U13810 (N_13810,N_13635,N_13513);
and U13811 (N_13811,N_13525,N_13714);
and U13812 (N_13812,N_13625,N_13678);
and U13813 (N_13813,N_13634,N_13648);
nand U13814 (N_13814,N_13584,N_13540);
nor U13815 (N_13815,N_13660,N_13533);
or U13816 (N_13816,N_13702,N_13649);
nor U13817 (N_13817,N_13708,N_13512);
and U13818 (N_13818,N_13628,N_13521);
or U13819 (N_13819,N_13528,N_13546);
and U13820 (N_13820,N_13723,N_13697);
or U13821 (N_13821,N_13562,N_13596);
nand U13822 (N_13822,N_13643,N_13573);
nor U13823 (N_13823,N_13560,N_13602);
nand U13824 (N_13824,N_13691,N_13698);
nand U13825 (N_13825,N_13547,N_13531);
nand U13826 (N_13826,N_13516,N_13556);
nand U13827 (N_13827,N_13665,N_13621);
nand U13828 (N_13828,N_13503,N_13589);
nand U13829 (N_13829,N_13654,N_13618);
nand U13830 (N_13830,N_13667,N_13568);
nand U13831 (N_13831,N_13590,N_13668);
nor U13832 (N_13832,N_13662,N_13500);
or U13833 (N_13833,N_13682,N_13583);
nor U13834 (N_13834,N_13510,N_13737);
xor U13835 (N_13835,N_13626,N_13627);
and U13836 (N_13836,N_13507,N_13683);
and U13837 (N_13837,N_13739,N_13669);
nor U13838 (N_13838,N_13504,N_13684);
nand U13839 (N_13839,N_13579,N_13636);
nor U13840 (N_13840,N_13672,N_13617);
xnor U13841 (N_13841,N_13542,N_13534);
xor U13842 (N_13842,N_13689,N_13677);
and U13843 (N_13843,N_13680,N_13718);
nand U13844 (N_13844,N_13713,N_13557);
xnor U13845 (N_13845,N_13600,N_13690);
nor U13846 (N_13846,N_13519,N_13538);
or U13847 (N_13847,N_13743,N_13539);
nor U13848 (N_13848,N_13658,N_13748);
or U13849 (N_13849,N_13616,N_13715);
nor U13850 (N_13850,N_13736,N_13676);
nor U13851 (N_13851,N_13657,N_13614);
or U13852 (N_13852,N_13652,N_13545);
xnor U13853 (N_13853,N_13638,N_13747);
nand U13854 (N_13854,N_13514,N_13536);
nand U13855 (N_13855,N_13524,N_13661);
xnor U13856 (N_13856,N_13645,N_13505);
and U13857 (N_13857,N_13709,N_13515);
nor U13858 (N_13858,N_13671,N_13732);
xnor U13859 (N_13859,N_13575,N_13740);
nor U13860 (N_13860,N_13719,N_13612);
nand U13861 (N_13861,N_13607,N_13642);
nand U13862 (N_13862,N_13517,N_13720);
and U13863 (N_13863,N_13655,N_13599);
and U13864 (N_13864,N_13569,N_13620);
nand U13865 (N_13865,N_13735,N_13624);
xor U13866 (N_13866,N_13631,N_13572);
xnor U13867 (N_13867,N_13629,N_13592);
or U13868 (N_13868,N_13567,N_13622);
nand U13869 (N_13869,N_13501,N_13659);
or U13870 (N_13870,N_13587,N_13656);
xor U13871 (N_13871,N_13644,N_13734);
and U13872 (N_13872,N_13696,N_13613);
xor U13873 (N_13873,N_13527,N_13580);
nor U13874 (N_13874,N_13681,N_13520);
xor U13875 (N_13875,N_13500,N_13692);
or U13876 (N_13876,N_13504,N_13542);
nand U13877 (N_13877,N_13568,N_13606);
and U13878 (N_13878,N_13720,N_13644);
or U13879 (N_13879,N_13684,N_13679);
nor U13880 (N_13880,N_13739,N_13746);
nor U13881 (N_13881,N_13564,N_13606);
xnor U13882 (N_13882,N_13661,N_13508);
xnor U13883 (N_13883,N_13707,N_13743);
and U13884 (N_13884,N_13672,N_13596);
or U13885 (N_13885,N_13635,N_13666);
nand U13886 (N_13886,N_13639,N_13570);
and U13887 (N_13887,N_13662,N_13717);
and U13888 (N_13888,N_13679,N_13579);
nor U13889 (N_13889,N_13523,N_13610);
nor U13890 (N_13890,N_13595,N_13556);
xnor U13891 (N_13891,N_13533,N_13575);
and U13892 (N_13892,N_13586,N_13725);
and U13893 (N_13893,N_13543,N_13558);
and U13894 (N_13894,N_13596,N_13607);
and U13895 (N_13895,N_13621,N_13673);
xnor U13896 (N_13896,N_13620,N_13554);
or U13897 (N_13897,N_13744,N_13529);
nand U13898 (N_13898,N_13642,N_13654);
or U13899 (N_13899,N_13542,N_13722);
xor U13900 (N_13900,N_13641,N_13592);
or U13901 (N_13901,N_13536,N_13616);
nor U13902 (N_13902,N_13713,N_13626);
nand U13903 (N_13903,N_13664,N_13528);
and U13904 (N_13904,N_13595,N_13667);
or U13905 (N_13905,N_13732,N_13647);
or U13906 (N_13906,N_13619,N_13704);
xor U13907 (N_13907,N_13661,N_13505);
nor U13908 (N_13908,N_13736,N_13567);
nand U13909 (N_13909,N_13704,N_13596);
nand U13910 (N_13910,N_13660,N_13560);
or U13911 (N_13911,N_13565,N_13584);
nand U13912 (N_13912,N_13560,N_13699);
or U13913 (N_13913,N_13682,N_13610);
nor U13914 (N_13914,N_13720,N_13687);
nor U13915 (N_13915,N_13558,N_13740);
and U13916 (N_13916,N_13534,N_13518);
nand U13917 (N_13917,N_13655,N_13583);
or U13918 (N_13918,N_13583,N_13745);
nor U13919 (N_13919,N_13652,N_13529);
nand U13920 (N_13920,N_13718,N_13692);
xor U13921 (N_13921,N_13710,N_13529);
xor U13922 (N_13922,N_13631,N_13563);
xor U13923 (N_13923,N_13515,N_13749);
nand U13924 (N_13924,N_13529,N_13503);
or U13925 (N_13925,N_13603,N_13502);
xnor U13926 (N_13926,N_13650,N_13640);
or U13927 (N_13927,N_13728,N_13667);
nand U13928 (N_13928,N_13564,N_13643);
or U13929 (N_13929,N_13645,N_13533);
xor U13930 (N_13930,N_13740,N_13570);
and U13931 (N_13931,N_13626,N_13526);
xor U13932 (N_13932,N_13748,N_13703);
xnor U13933 (N_13933,N_13678,N_13528);
or U13934 (N_13934,N_13740,N_13700);
nor U13935 (N_13935,N_13639,N_13541);
xor U13936 (N_13936,N_13675,N_13561);
and U13937 (N_13937,N_13733,N_13657);
or U13938 (N_13938,N_13594,N_13667);
or U13939 (N_13939,N_13692,N_13506);
nand U13940 (N_13940,N_13603,N_13548);
xor U13941 (N_13941,N_13704,N_13573);
or U13942 (N_13942,N_13671,N_13692);
nand U13943 (N_13943,N_13553,N_13627);
xor U13944 (N_13944,N_13546,N_13694);
nand U13945 (N_13945,N_13598,N_13705);
nand U13946 (N_13946,N_13740,N_13685);
or U13947 (N_13947,N_13620,N_13678);
or U13948 (N_13948,N_13607,N_13694);
xor U13949 (N_13949,N_13733,N_13692);
or U13950 (N_13950,N_13511,N_13633);
and U13951 (N_13951,N_13505,N_13647);
nand U13952 (N_13952,N_13508,N_13720);
xnor U13953 (N_13953,N_13546,N_13630);
nand U13954 (N_13954,N_13741,N_13508);
xor U13955 (N_13955,N_13606,N_13726);
xnor U13956 (N_13956,N_13664,N_13524);
and U13957 (N_13957,N_13680,N_13738);
or U13958 (N_13958,N_13668,N_13661);
or U13959 (N_13959,N_13641,N_13652);
nand U13960 (N_13960,N_13607,N_13743);
nor U13961 (N_13961,N_13520,N_13643);
nor U13962 (N_13962,N_13737,N_13607);
nand U13963 (N_13963,N_13608,N_13574);
and U13964 (N_13964,N_13566,N_13697);
xnor U13965 (N_13965,N_13553,N_13532);
or U13966 (N_13966,N_13699,N_13545);
xnor U13967 (N_13967,N_13602,N_13732);
and U13968 (N_13968,N_13564,N_13657);
nand U13969 (N_13969,N_13609,N_13604);
nand U13970 (N_13970,N_13694,N_13613);
nor U13971 (N_13971,N_13720,N_13662);
xnor U13972 (N_13972,N_13623,N_13533);
nor U13973 (N_13973,N_13655,N_13642);
xnor U13974 (N_13974,N_13618,N_13615);
and U13975 (N_13975,N_13552,N_13624);
nor U13976 (N_13976,N_13701,N_13690);
or U13977 (N_13977,N_13683,N_13642);
nand U13978 (N_13978,N_13730,N_13729);
and U13979 (N_13979,N_13535,N_13586);
or U13980 (N_13980,N_13725,N_13611);
xnor U13981 (N_13981,N_13674,N_13713);
and U13982 (N_13982,N_13631,N_13657);
nor U13983 (N_13983,N_13628,N_13526);
nor U13984 (N_13984,N_13641,N_13518);
and U13985 (N_13985,N_13576,N_13703);
nor U13986 (N_13986,N_13713,N_13711);
nand U13987 (N_13987,N_13653,N_13715);
nor U13988 (N_13988,N_13539,N_13739);
or U13989 (N_13989,N_13535,N_13537);
nor U13990 (N_13990,N_13570,N_13563);
xor U13991 (N_13991,N_13602,N_13703);
xor U13992 (N_13992,N_13634,N_13652);
xor U13993 (N_13993,N_13746,N_13725);
and U13994 (N_13994,N_13509,N_13570);
nor U13995 (N_13995,N_13613,N_13610);
xor U13996 (N_13996,N_13702,N_13621);
xnor U13997 (N_13997,N_13600,N_13630);
or U13998 (N_13998,N_13699,N_13703);
nor U13999 (N_13999,N_13681,N_13608);
nand U14000 (N_14000,N_13868,N_13807);
xor U14001 (N_14001,N_13859,N_13922);
xor U14002 (N_14002,N_13801,N_13840);
nand U14003 (N_14003,N_13758,N_13972);
xnor U14004 (N_14004,N_13926,N_13969);
or U14005 (N_14005,N_13763,N_13844);
nor U14006 (N_14006,N_13915,N_13809);
and U14007 (N_14007,N_13776,N_13950);
and U14008 (N_14008,N_13970,N_13762);
nor U14009 (N_14009,N_13949,N_13906);
nor U14010 (N_14010,N_13799,N_13914);
and U14011 (N_14011,N_13803,N_13933);
nor U14012 (N_14012,N_13897,N_13887);
and U14013 (N_14013,N_13790,N_13753);
xor U14014 (N_14014,N_13827,N_13927);
xor U14015 (N_14015,N_13759,N_13813);
nor U14016 (N_14016,N_13957,N_13929);
xnor U14017 (N_14017,N_13854,N_13769);
nand U14018 (N_14018,N_13958,N_13888);
xor U14019 (N_14019,N_13898,N_13931);
xnor U14020 (N_14020,N_13856,N_13984);
nor U14021 (N_14021,N_13766,N_13891);
or U14022 (N_14022,N_13913,N_13923);
xor U14023 (N_14023,N_13981,N_13797);
xnor U14024 (N_14024,N_13953,N_13967);
xor U14025 (N_14025,N_13858,N_13987);
or U14026 (N_14026,N_13983,N_13902);
nand U14027 (N_14027,N_13794,N_13848);
or U14028 (N_14028,N_13781,N_13966);
or U14029 (N_14029,N_13889,N_13946);
and U14030 (N_14030,N_13814,N_13826);
nand U14031 (N_14031,N_13876,N_13863);
nor U14032 (N_14032,N_13764,N_13788);
or U14033 (N_14033,N_13767,N_13978);
xnor U14034 (N_14034,N_13985,N_13991);
and U14035 (N_14035,N_13935,N_13824);
nand U14036 (N_14036,N_13785,N_13941);
or U14037 (N_14037,N_13928,N_13884);
xnor U14038 (N_14038,N_13752,N_13895);
nor U14039 (N_14039,N_13943,N_13837);
or U14040 (N_14040,N_13880,N_13832);
nand U14041 (N_14041,N_13921,N_13833);
nand U14042 (N_14042,N_13800,N_13999);
xnor U14043 (N_14043,N_13937,N_13839);
or U14044 (N_14044,N_13924,N_13835);
nor U14045 (N_14045,N_13910,N_13894);
nor U14046 (N_14046,N_13772,N_13783);
and U14047 (N_14047,N_13851,N_13770);
xnor U14048 (N_14048,N_13874,N_13979);
nand U14049 (N_14049,N_13892,N_13820);
or U14050 (N_14050,N_13817,N_13920);
nand U14051 (N_14051,N_13789,N_13756);
or U14052 (N_14052,N_13919,N_13871);
xor U14053 (N_14053,N_13791,N_13883);
and U14054 (N_14054,N_13954,N_13836);
xor U14055 (N_14055,N_13805,N_13911);
and U14056 (N_14056,N_13806,N_13912);
nand U14057 (N_14057,N_13901,N_13878);
nor U14058 (N_14058,N_13852,N_13964);
xnor U14059 (N_14059,N_13899,N_13900);
nor U14060 (N_14060,N_13793,N_13940);
xor U14061 (N_14061,N_13822,N_13877);
or U14062 (N_14062,N_13786,N_13962);
nand U14063 (N_14063,N_13829,N_13952);
and U14064 (N_14064,N_13778,N_13821);
or U14065 (N_14065,N_13944,N_13872);
and U14066 (N_14066,N_13968,N_13959);
and U14067 (N_14067,N_13867,N_13860);
and U14068 (N_14068,N_13986,N_13751);
nor U14069 (N_14069,N_13916,N_13975);
nand U14070 (N_14070,N_13761,N_13825);
or U14071 (N_14071,N_13828,N_13875);
nand U14072 (N_14072,N_13938,N_13903);
and U14073 (N_14073,N_13965,N_13784);
and U14074 (N_14074,N_13768,N_13909);
xor U14075 (N_14075,N_13792,N_13947);
nand U14076 (N_14076,N_13974,N_13896);
nand U14077 (N_14077,N_13930,N_13990);
and U14078 (N_14078,N_13780,N_13841);
or U14079 (N_14079,N_13750,N_13849);
or U14080 (N_14080,N_13996,N_13823);
nand U14081 (N_14081,N_13936,N_13818);
and U14082 (N_14082,N_13886,N_13870);
nor U14083 (N_14083,N_13760,N_13810);
xnor U14084 (N_14084,N_13908,N_13798);
or U14085 (N_14085,N_13948,N_13771);
or U14086 (N_14086,N_13997,N_13779);
nor U14087 (N_14087,N_13942,N_13834);
nor U14088 (N_14088,N_13838,N_13774);
or U14089 (N_14089,N_13861,N_13918);
nor U14090 (N_14090,N_13879,N_13773);
nor U14091 (N_14091,N_13869,N_13796);
nor U14092 (N_14092,N_13865,N_13843);
nand U14093 (N_14093,N_13932,N_13995);
xor U14094 (N_14094,N_13956,N_13804);
nand U14095 (N_14095,N_13775,N_13846);
and U14096 (N_14096,N_13815,N_13993);
or U14097 (N_14097,N_13988,N_13917);
xnor U14098 (N_14098,N_13830,N_13939);
or U14099 (N_14099,N_13971,N_13857);
xnor U14100 (N_14100,N_13982,N_13808);
nand U14101 (N_14101,N_13998,N_13755);
or U14102 (N_14102,N_13905,N_13882);
and U14103 (N_14103,N_13955,N_13989);
or U14104 (N_14104,N_13864,N_13754);
nand U14105 (N_14105,N_13994,N_13976);
nand U14106 (N_14106,N_13925,N_13812);
nand U14107 (N_14107,N_13777,N_13757);
nand U14108 (N_14108,N_13963,N_13873);
nor U14109 (N_14109,N_13890,N_13885);
and U14110 (N_14110,N_13816,N_13904);
or U14111 (N_14111,N_13893,N_13951);
and U14112 (N_14112,N_13855,N_13819);
xnor U14113 (N_14113,N_13845,N_13853);
and U14114 (N_14114,N_13977,N_13934);
and U14115 (N_14115,N_13842,N_13765);
xnor U14116 (N_14116,N_13787,N_13850);
nand U14117 (N_14117,N_13811,N_13831);
nor U14118 (N_14118,N_13782,N_13973);
or U14119 (N_14119,N_13960,N_13992);
xor U14120 (N_14120,N_13945,N_13907);
nand U14121 (N_14121,N_13980,N_13802);
xnor U14122 (N_14122,N_13847,N_13961);
xor U14123 (N_14123,N_13881,N_13866);
nand U14124 (N_14124,N_13862,N_13795);
or U14125 (N_14125,N_13831,N_13903);
xnor U14126 (N_14126,N_13977,N_13892);
nand U14127 (N_14127,N_13785,N_13827);
nand U14128 (N_14128,N_13920,N_13846);
or U14129 (N_14129,N_13923,N_13892);
nor U14130 (N_14130,N_13889,N_13787);
nand U14131 (N_14131,N_13820,N_13948);
nor U14132 (N_14132,N_13798,N_13841);
nand U14133 (N_14133,N_13800,N_13766);
nor U14134 (N_14134,N_13763,N_13911);
and U14135 (N_14135,N_13766,N_13996);
nor U14136 (N_14136,N_13822,N_13750);
or U14137 (N_14137,N_13967,N_13932);
or U14138 (N_14138,N_13808,N_13793);
nand U14139 (N_14139,N_13824,N_13786);
nor U14140 (N_14140,N_13796,N_13931);
nand U14141 (N_14141,N_13804,N_13814);
nand U14142 (N_14142,N_13928,N_13797);
xor U14143 (N_14143,N_13849,N_13947);
or U14144 (N_14144,N_13937,N_13908);
or U14145 (N_14145,N_13876,N_13870);
nor U14146 (N_14146,N_13750,N_13924);
and U14147 (N_14147,N_13969,N_13849);
nor U14148 (N_14148,N_13799,N_13788);
and U14149 (N_14149,N_13886,N_13998);
nor U14150 (N_14150,N_13760,N_13880);
or U14151 (N_14151,N_13921,N_13999);
and U14152 (N_14152,N_13931,N_13831);
xor U14153 (N_14153,N_13965,N_13797);
nand U14154 (N_14154,N_13932,N_13779);
nor U14155 (N_14155,N_13841,N_13815);
and U14156 (N_14156,N_13885,N_13844);
and U14157 (N_14157,N_13928,N_13756);
xor U14158 (N_14158,N_13974,N_13919);
xnor U14159 (N_14159,N_13871,N_13781);
nor U14160 (N_14160,N_13753,N_13883);
or U14161 (N_14161,N_13880,N_13771);
or U14162 (N_14162,N_13995,N_13917);
xnor U14163 (N_14163,N_13885,N_13773);
xor U14164 (N_14164,N_13863,N_13921);
nor U14165 (N_14165,N_13790,N_13766);
or U14166 (N_14166,N_13942,N_13881);
or U14167 (N_14167,N_13841,N_13994);
xnor U14168 (N_14168,N_13858,N_13807);
nor U14169 (N_14169,N_13991,N_13983);
and U14170 (N_14170,N_13915,N_13922);
and U14171 (N_14171,N_13951,N_13770);
and U14172 (N_14172,N_13995,N_13941);
and U14173 (N_14173,N_13789,N_13936);
nor U14174 (N_14174,N_13998,N_13941);
or U14175 (N_14175,N_13978,N_13934);
xor U14176 (N_14176,N_13784,N_13942);
nand U14177 (N_14177,N_13770,N_13850);
nor U14178 (N_14178,N_13993,N_13805);
xnor U14179 (N_14179,N_13888,N_13901);
nor U14180 (N_14180,N_13833,N_13882);
and U14181 (N_14181,N_13978,N_13931);
or U14182 (N_14182,N_13950,N_13960);
nand U14183 (N_14183,N_13842,N_13965);
nor U14184 (N_14184,N_13857,N_13988);
xnor U14185 (N_14185,N_13773,N_13915);
and U14186 (N_14186,N_13976,N_13958);
or U14187 (N_14187,N_13798,N_13889);
nor U14188 (N_14188,N_13804,N_13869);
and U14189 (N_14189,N_13916,N_13827);
nand U14190 (N_14190,N_13996,N_13976);
and U14191 (N_14191,N_13796,N_13842);
xor U14192 (N_14192,N_13995,N_13982);
or U14193 (N_14193,N_13789,N_13888);
and U14194 (N_14194,N_13780,N_13942);
nand U14195 (N_14195,N_13767,N_13789);
or U14196 (N_14196,N_13933,N_13978);
or U14197 (N_14197,N_13940,N_13908);
and U14198 (N_14198,N_13987,N_13760);
or U14199 (N_14199,N_13980,N_13818);
and U14200 (N_14200,N_13910,N_13858);
nor U14201 (N_14201,N_13972,N_13960);
or U14202 (N_14202,N_13843,N_13787);
or U14203 (N_14203,N_13933,N_13863);
xnor U14204 (N_14204,N_13820,N_13805);
and U14205 (N_14205,N_13828,N_13787);
nor U14206 (N_14206,N_13820,N_13946);
and U14207 (N_14207,N_13828,N_13919);
nor U14208 (N_14208,N_13853,N_13913);
nand U14209 (N_14209,N_13929,N_13887);
xnor U14210 (N_14210,N_13999,N_13946);
and U14211 (N_14211,N_13755,N_13754);
or U14212 (N_14212,N_13854,N_13819);
nand U14213 (N_14213,N_13777,N_13911);
nand U14214 (N_14214,N_13865,N_13935);
xnor U14215 (N_14215,N_13800,N_13864);
nor U14216 (N_14216,N_13907,N_13964);
xnor U14217 (N_14217,N_13764,N_13889);
xnor U14218 (N_14218,N_13883,N_13937);
nor U14219 (N_14219,N_13990,N_13790);
or U14220 (N_14220,N_13766,N_13889);
xor U14221 (N_14221,N_13767,N_13794);
nand U14222 (N_14222,N_13981,N_13928);
and U14223 (N_14223,N_13820,N_13798);
nand U14224 (N_14224,N_13774,N_13784);
xnor U14225 (N_14225,N_13902,N_13823);
nand U14226 (N_14226,N_13882,N_13792);
or U14227 (N_14227,N_13858,N_13941);
nand U14228 (N_14228,N_13812,N_13824);
and U14229 (N_14229,N_13932,N_13805);
or U14230 (N_14230,N_13906,N_13757);
or U14231 (N_14231,N_13792,N_13899);
or U14232 (N_14232,N_13937,N_13804);
or U14233 (N_14233,N_13788,N_13933);
nor U14234 (N_14234,N_13763,N_13987);
or U14235 (N_14235,N_13924,N_13988);
xor U14236 (N_14236,N_13806,N_13775);
nor U14237 (N_14237,N_13905,N_13990);
nand U14238 (N_14238,N_13967,N_13827);
or U14239 (N_14239,N_13861,N_13769);
or U14240 (N_14240,N_13792,N_13773);
or U14241 (N_14241,N_13847,N_13802);
and U14242 (N_14242,N_13900,N_13864);
nor U14243 (N_14243,N_13863,N_13908);
nand U14244 (N_14244,N_13843,N_13992);
or U14245 (N_14245,N_13884,N_13943);
or U14246 (N_14246,N_13770,N_13864);
and U14247 (N_14247,N_13800,N_13885);
nor U14248 (N_14248,N_13784,N_13931);
xnor U14249 (N_14249,N_13948,N_13893);
or U14250 (N_14250,N_14050,N_14140);
nand U14251 (N_14251,N_14039,N_14189);
or U14252 (N_14252,N_14207,N_14054);
nor U14253 (N_14253,N_14209,N_14215);
or U14254 (N_14254,N_14094,N_14174);
or U14255 (N_14255,N_14161,N_14180);
nand U14256 (N_14256,N_14240,N_14100);
xor U14257 (N_14257,N_14076,N_14157);
nor U14258 (N_14258,N_14142,N_14176);
xor U14259 (N_14259,N_14072,N_14159);
xor U14260 (N_14260,N_14018,N_14058);
nand U14261 (N_14261,N_14109,N_14113);
and U14262 (N_14262,N_14214,N_14037);
xor U14263 (N_14263,N_14235,N_14181);
nand U14264 (N_14264,N_14167,N_14231);
and U14265 (N_14265,N_14194,N_14036);
xor U14266 (N_14266,N_14229,N_14073);
or U14267 (N_14267,N_14020,N_14226);
xor U14268 (N_14268,N_14186,N_14218);
nand U14269 (N_14269,N_14243,N_14144);
nor U14270 (N_14270,N_14038,N_14211);
xnor U14271 (N_14271,N_14079,N_14178);
xnor U14272 (N_14272,N_14024,N_14051);
or U14273 (N_14273,N_14217,N_14083);
or U14274 (N_14274,N_14033,N_14241);
nand U14275 (N_14275,N_14119,N_14198);
or U14276 (N_14276,N_14108,N_14136);
and U14277 (N_14277,N_14089,N_14114);
and U14278 (N_14278,N_14222,N_14173);
or U14279 (N_14279,N_14216,N_14213);
xor U14280 (N_14280,N_14009,N_14154);
xor U14281 (N_14281,N_14202,N_14201);
nand U14282 (N_14282,N_14004,N_14148);
nand U14283 (N_14283,N_14099,N_14117);
and U14284 (N_14284,N_14078,N_14152);
xor U14285 (N_14285,N_14046,N_14234);
and U14286 (N_14286,N_14184,N_14044);
or U14287 (N_14287,N_14171,N_14014);
nand U14288 (N_14288,N_14121,N_14160);
xnor U14289 (N_14289,N_14238,N_14177);
or U14290 (N_14290,N_14026,N_14191);
and U14291 (N_14291,N_14056,N_14230);
xnor U14292 (N_14292,N_14132,N_14233);
and U14293 (N_14293,N_14182,N_14065);
or U14294 (N_14294,N_14059,N_14248);
and U14295 (N_14295,N_14002,N_14013);
nor U14296 (N_14296,N_14029,N_14031);
xor U14297 (N_14297,N_14011,N_14122);
and U14298 (N_14298,N_14197,N_14224);
nand U14299 (N_14299,N_14175,N_14082);
nor U14300 (N_14300,N_14055,N_14049);
xnor U14301 (N_14301,N_14162,N_14067);
and U14302 (N_14302,N_14156,N_14118);
and U14303 (N_14303,N_14110,N_14149);
nor U14304 (N_14304,N_14115,N_14012);
nor U14305 (N_14305,N_14168,N_14090);
xor U14306 (N_14306,N_14153,N_14185);
nand U14307 (N_14307,N_14223,N_14120);
xnor U14308 (N_14308,N_14021,N_14138);
or U14309 (N_14309,N_14084,N_14096);
and U14310 (N_14310,N_14028,N_14208);
nor U14311 (N_14311,N_14183,N_14069);
and U14312 (N_14312,N_14077,N_14145);
nand U14313 (N_14313,N_14066,N_14068);
xnor U14314 (N_14314,N_14212,N_14027);
nor U14315 (N_14315,N_14095,N_14228);
nor U14316 (N_14316,N_14111,N_14131);
xnor U14317 (N_14317,N_14040,N_14003);
nor U14318 (N_14318,N_14200,N_14133);
and U14319 (N_14319,N_14116,N_14048);
nand U14320 (N_14320,N_14199,N_14219);
and U14321 (N_14321,N_14101,N_14242);
and U14322 (N_14322,N_14166,N_14093);
nand U14323 (N_14323,N_14220,N_14203);
and U14324 (N_14324,N_14045,N_14103);
nand U14325 (N_14325,N_14022,N_14104);
nor U14326 (N_14326,N_14081,N_14080);
or U14327 (N_14327,N_14071,N_14225);
and U14328 (N_14328,N_14025,N_14000);
or U14329 (N_14329,N_14102,N_14106);
xor U14330 (N_14330,N_14232,N_14179);
nor U14331 (N_14331,N_14005,N_14057);
nor U14332 (N_14332,N_14210,N_14052);
nor U14333 (N_14333,N_14170,N_14006);
or U14334 (N_14334,N_14008,N_14196);
xor U14335 (N_14335,N_14035,N_14147);
nand U14336 (N_14336,N_14123,N_14017);
or U14337 (N_14337,N_14129,N_14062);
nand U14338 (N_14338,N_14074,N_14127);
xor U14339 (N_14339,N_14139,N_14098);
or U14340 (N_14340,N_14164,N_14016);
nand U14341 (N_14341,N_14187,N_14150);
nand U14342 (N_14342,N_14092,N_14195);
nor U14343 (N_14343,N_14030,N_14125);
or U14344 (N_14344,N_14128,N_14091);
and U14345 (N_14345,N_14247,N_14236);
or U14346 (N_14346,N_14239,N_14060);
nand U14347 (N_14347,N_14158,N_14227);
nand U14348 (N_14348,N_14015,N_14032);
nand U14349 (N_14349,N_14134,N_14019);
xnor U14350 (N_14350,N_14075,N_14192);
or U14351 (N_14351,N_14193,N_14135);
xor U14352 (N_14352,N_14107,N_14126);
xor U14353 (N_14353,N_14188,N_14001);
or U14354 (N_14354,N_14137,N_14086);
or U14355 (N_14355,N_14061,N_14023);
or U14356 (N_14356,N_14143,N_14070);
xnor U14357 (N_14357,N_14249,N_14007);
xor U14358 (N_14358,N_14053,N_14043);
or U14359 (N_14359,N_14105,N_14087);
xnor U14360 (N_14360,N_14172,N_14112);
nand U14361 (N_14361,N_14041,N_14010);
nand U14362 (N_14362,N_14246,N_14190);
nor U14363 (N_14363,N_14245,N_14130);
or U14364 (N_14364,N_14042,N_14047);
nor U14365 (N_14365,N_14237,N_14155);
nor U14366 (N_14366,N_14085,N_14063);
or U14367 (N_14367,N_14206,N_14124);
nor U14368 (N_14368,N_14064,N_14169);
and U14369 (N_14369,N_14204,N_14205);
nor U14370 (N_14370,N_14221,N_14163);
or U14371 (N_14371,N_14088,N_14146);
nand U14372 (N_14372,N_14244,N_14034);
or U14373 (N_14373,N_14151,N_14141);
nor U14374 (N_14374,N_14165,N_14097);
nor U14375 (N_14375,N_14249,N_14248);
xor U14376 (N_14376,N_14017,N_14063);
xnor U14377 (N_14377,N_14217,N_14071);
xor U14378 (N_14378,N_14137,N_14142);
and U14379 (N_14379,N_14128,N_14144);
nand U14380 (N_14380,N_14133,N_14025);
nand U14381 (N_14381,N_14205,N_14184);
or U14382 (N_14382,N_14209,N_14078);
xor U14383 (N_14383,N_14140,N_14158);
xnor U14384 (N_14384,N_14245,N_14168);
xnor U14385 (N_14385,N_14201,N_14036);
xor U14386 (N_14386,N_14086,N_14061);
and U14387 (N_14387,N_14050,N_14110);
and U14388 (N_14388,N_14051,N_14165);
and U14389 (N_14389,N_14232,N_14247);
nand U14390 (N_14390,N_14234,N_14242);
nand U14391 (N_14391,N_14145,N_14015);
xnor U14392 (N_14392,N_14013,N_14043);
xnor U14393 (N_14393,N_14191,N_14168);
nor U14394 (N_14394,N_14208,N_14055);
or U14395 (N_14395,N_14110,N_14069);
xor U14396 (N_14396,N_14008,N_14081);
nor U14397 (N_14397,N_14246,N_14000);
nor U14398 (N_14398,N_14178,N_14239);
and U14399 (N_14399,N_14081,N_14007);
and U14400 (N_14400,N_14085,N_14126);
and U14401 (N_14401,N_14090,N_14217);
xnor U14402 (N_14402,N_14029,N_14004);
xnor U14403 (N_14403,N_14151,N_14019);
or U14404 (N_14404,N_14095,N_14235);
nor U14405 (N_14405,N_14124,N_14131);
nand U14406 (N_14406,N_14160,N_14004);
and U14407 (N_14407,N_14125,N_14124);
and U14408 (N_14408,N_14210,N_14103);
xnor U14409 (N_14409,N_14118,N_14141);
nand U14410 (N_14410,N_14248,N_14009);
and U14411 (N_14411,N_14116,N_14055);
nor U14412 (N_14412,N_14141,N_14249);
nor U14413 (N_14413,N_14023,N_14069);
xnor U14414 (N_14414,N_14210,N_14005);
nor U14415 (N_14415,N_14021,N_14135);
xnor U14416 (N_14416,N_14002,N_14053);
nor U14417 (N_14417,N_14039,N_14096);
nor U14418 (N_14418,N_14001,N_14164);
nand U14419 (N_14419,N_14116,N_14133);
and U14420 (N_14420,N_14017,N_14243);
nand U14421 (N_14421,N_14248,N_14232);
xor U14422 (N_14422,N_14102,N_14025);
or U14423 (N_14423,N_14229,N_14193);
nand U14424 (N_14424,N_14193,N_14198);
nand U14425 (N_14425,N_14144,N_14137);
xor U14426 (N_14426,N_14062,N_14228);
nor U14427 (N_14427,N_14076,N_14032);
or U14428 (N_14428,N_14011,N_14048);
nand U14429 (N_14429,N_14183,N_14064);
nor U14430 (N_14430,N_14173,N_14218);
or U14431 (N_14431,N_14234,N_14156);
xor U14432 (N_14432,N_14172,N_14166);
or U14433 (N_14433,N_14173,N_14044);
xnor U14434 (N_14434,N_14002,N_14010);
xnor U14435 (N_14435,N_14029,N_14063);
nor U14436 (N_14436,N_14028,N_14056);
and U14437 (N_14437,N_14185,N_14139);
and U14438 (N_14438,N_14238,N_14020);
and U14439 (N_14439,N_14024,N_14073);
or U14440 (N_14440,N_14238,N_14115);
or U14441 (N_14441,N_14043,N_14215);
and U14442 (N_14442,N_14048,N_14097);
xnor U14443 (N_14443,N_14222,N_14215);
or U14444 (N_14444,N_14003,N_14148);
or U14445 (N_14445,N_14066,N_14131);
nand U14446 (N_14446,N_14205,N_14211);
or U14447 (N_14447,N_14002,N_14192);
nand U14448 (N_14448,N_14216,N_14198);
nand U14449 (N_14449,N_14193,N_14225);
or U14450 (N_14450,N_14236,N_14165);
nand U14451 (N_14451,N_14019,N_14135);
nor U14452 (N_14452,N_14060,N_14096);
xnor U14453 (N_14453,N_14109,N_14137);
xnor U14454 (N_14454,N_14011,N_14016);
and U14455 (N_14455,N_14036,N_14115);
xnor U14456 (N_14456,N_14021,N_14234);
nand U14457 (N_14457,N_14027,N_14003);
xor U14458 (N_14458,N_14143,N_14035);
and U14459 (N_14459,N_14139,N_14012);
or U14460 (N_14460,N_14135,N_14232);
nor U14461 (N_14461,N_14222,N_14207);
nor U14462 (N_14462,N_14151,N_14041);
or U14463 (N_14463,N_14233,N_14046);
nor U14464 (N_14464,N_14153,N_14162);
and U14465 (N_14465,N_14210,N_14229);
and U14466 (N_14466,N_14023,N_14194);
nand U14467 (N_14467,N_14020,N_14170);
nor U14468 (N_14468,N_14241,N_14003);
xor U14469 (N_14469,N_14246,N_14097);
nand U14470 (N_14470,N_14169,N_14145);
nor U14471 (N_14471,N_14154,N_14144);
nor U14472 (N_14472,N_14180,N_14113);
nand U14473 (N_14473,N_14188,N_14028);
xor U14474 (N_14474,N_14123,N_14126);
or U14475 (N_14475,N_14003,N_14092);
or U14476 (N_14476,N_14141,N_14150);
or U14477 (N_14477,N_14011,N_14083);
nor U14478 (N_14478,N_14190,N_14033);
and U14479 (N_14479,N_14189,N_14050);
nor U14480 (N_14480,N_14196,N_14165);
nand U14481 (N_14481,N_14058,N_14068);
xnor U14482 (N_14482,N_14057,N_14240);
and U14483 (N_14483,N_14238,N_14015);
or U14484 (N_14484,N_14062,N_14092);
nand U14485 (N_14485,N_14122,N_14174);
or U14486 (N_14486,N_14049,N_14177);
nand U14487 (N_14487,N_14223,N_14080);
nor U14488 (N_14488,N_14045,N_14112);
or U14489 (N_14489,N_14234,N_14045);
and U14490 (N_14490,N_14185,N_14129);
nor U14491 (N_14491,N_14129,N_14126);
or U14492 (N_14492,N_14019,N_14067);
xnor U14493 (N_14493,N_14213,N_14007);
xor U14494 (N_14494,N_14048,N_14003);
or U14495 (N_14495,N_14127,N_14164);
nor U14496 (N_14496,N_14086,N_14189);
nor U14497 (N_14497,N_14240,N_14137);
or U14498 (N_14498,N_14180,N_14155);
nand U14499 (N_14499,N_14166,N_14217);
nand U14500 (N_14500,N_14309,N_14361);
nor U14501 (N_14501,N_14386,N_14308);
nand U14502 (N_14502,N_14275,N_14450);
nand U14503 (N_14503,N_14460,N_14335);
nor U14504 (N_14504,N_14458,N_14486);
nand U14505 (N_14505,N_14409,N_14349);
nor U14506 (N_14506,N_14387,N_14461);
or U14507 (N_14507,N_14397,N_14297);
and U14508 (N_14508,N_14265,N_14277);
xnor U14509 (N_14509,N_14396,N_14488);
xor U14510 (N_14510,N_14272,N_14414);
xnor U14511 (N_14511,N_14364,N_14378);
and U14512 (N_14512,N_14467,N_14348);
and U14513 (N_14513,N_14468,N_14260);
nand U14514 (N_14514,N_14324,N_14473);
or U14515 (N_14515,N_14452,N_14432);
nand U14516 (N_14516,N_14479,N_14471);
and U14517 (N_14517,N_14327,N_14415);
xnor U14518 (N_14518,N_14284,N_14384);
nand U14519 (N_14519,N_14363,N_14404);
nor U14520 (N_14520,N_14377,N_14298);
xor U14521 (N_14521,N_14395,N_14426);
and U14522 (N_14522,N_14420,N_14328);
or U14523 (N_14523,N_14489,N_14312);
and U14524 (N_14524,N_14494,N_14388);
nand U14525 (N_14525,N_14399,N_14441);
nand U14526 (N_14526,N_14398,N_14436);
nor U14527 (N_14527,N_14266,N_14339);
or U14528 (N_14528,N_14371,N_14331);
nand U14529 (N_14529,N_14394,N_14310);
nand U14530 (N_14530,N_14448,N_14251);
or U14531 (N_14531,N_14434,N_14317);
or U14532 (N_14532,N_14304,N_14342);
xnor U14533 (N_14533,N_14355,N_14367);
and U14534 (N_14534,N_14336,N_14358);
nand U14535 (N_14535,N_14411,N_14430);
nor U14536 (N_14536,N_14492,N_14465);
and U14537 (N_14537,N_14498,N_14445);
nor U14538 (N_14538,N_14282,N_14424);
nand U14539 (N_14539,N_14289,N_14259);
or U14540 (N_14540,N_14346,N_14359);
nand U14541 (N_14541,N_14290,N_14405);
xnor U14542 (N_14542,N_14319,N_14372);
nand U14543 (N_14543,N_14357,N_14279);
nor U14544 (N_14544,N_14316,N_14254);
or U14545 (N_14545,N_14439,N_14256);
nor U14546 (N_14546,N_14285,N_14446);
or U14547 (N_14547,N_14493,N_14269);
nand U14548 (N_14548,N_14354,N_14403);
nand U14549 (N_14549,N_14487,N_14470);
nand U14550 (N_14550,N_14410,N_14307);
or U14551 (N_14551,N_14318,N_14495);
xnor U14552 (N_14552,N_14286,N_14499);
nor U14553 (N_14553,N_14330,N_14255);
and U14554 (N_14554,N_14370,N_14440);
nor U14555 (N_14555,N_14303,N_14369);
nand U14556 (N_14556,N_14427,N_14345);
nor U14557 (N_14557,N_14302,N_14484);
xor U14558 (N_14558,N_14301,N_14314);
and U14559 (N_14559,N_14347,N_14428);
nand U14560 (N_14560,N_14326,N_14464);
xor U14561 (N_14561,N_14469,N_14380);
xnor U14562 (N_14562,N_14299,N_14422);
nor U14563 (N_14563,N_14274,N_14315);
xnor U14564 (N_14564,N_14273,N_14456);
nand U14565 (N_14565,N_14323,N_14338);
xor U14566 (N_14566,N_14287,N_14393);
nand U14567 (N_14567,N_14413,N_14313);
xnor U14568 (N_14568,N_14350,N_14383);
or U14569 (N_14569,N_14258,N_14360);
nor U14570 (N_14570,N_14281,N_14477);
nand U14571 (N_14571,N_14278,N_14419);
nand U14572 (N_14572,N_14423,N_14293);
xor U14573 (N_14573,N_14332,N_14344);
nor U14574 (N_14574,N_14270,N_14463);
nand U14575 (N_14575,N_14447,N_14392);
xor U14576 (N_14576,N_14276,N_14453);
and U14577 (N_14577,N_14476,N_14325);
xor U14578 (N_14578,N_14438,N_14454);
nand U14579 (N_14579,N_14267,N_14381);
nand U14580 (N_14580,N_14296,N_14262);
nand U14581 (N_14581,N_14408,N_14390);
xor U14582 (N_14582,N_14412,N_14320);
nand U14583 (N_14583,N_14472,N_14368);
xnor U14584 (N_14584,N_14362,N_14429);
xnor U14585 (N_14585,N_14300,N_14433);
nor U14586 (N_14586,N_14253,N_14379);
xor U14587 (N_14587,N_14268,N_14491);
xnor U14588 (N_14588,N_14443,N_14457);
xnor U14589 (N_14589,N_14402,N_14264);
or U14590 (N_14590,N_14329,N_14442);
nor U14591 (N_14591,N_14366,N_14341);
or U14592 (N_14592,N_14451,N_14474);
nand U14593 (N_14593,N_14466,N_14437);
and U14594 (N_14594,N_14497,N_14496);
and U14595 (N_14595,N_14425,N_14333);
nor U14596 (N_14596,N_14283,N_14340);
nor U14597 (N_14597,N_14482,N_14280);
nand U14598 (N_14598,N_14261,N_14406);
or U14599 (N_14599,N_14391,N_14421);
xor U14600 (N_14600,N_14417,N_14375);
or U14601 (N_14601,N_14455,N_14418);
xor U14602 (N_14602,N_14490,N_14311);
nor U14603 (N_14603,N_14385,N_14483);
or U14604 (N_14604,N_14294,N_14305);
nor U14605 (N_14605,N_14252,N_14356);
nand U14606 (N_14606,N_14250,N_14382);
nand U14607 (N_14607,N_14376,N_14444);
nor U14608 (N_14608,N_14352,N_14351);
or U14609 (N_14609,N_14401,N_14263);
and U14610 (N_14610,N_14389,N_14365);
xor U14611 (N_14611,N_14353,N_14373);
nand U14612 (N_14612,N_14480,N_14321);
nor U14613 (N_14613,N_14435,N_14449);
nor U14614 (N_14614,N_14306,N_14431);
and U14615 (N_14615,N_14271,N_14485);
and U14616 (N_14616,N_14462,N_14343);
xor U14617 (N_14617,N_14322,N_14475);
nor U14618 (N_14618,N_14374,N_14407);
nor U14619 (N_14619,N_14334,N_14292);
nand U14620 (N_14620,N_14459,N_14400);
nand U14621 (N_14621,N_14291,N_14481);
xnor U14622 (N_14622,N_14478,N_14416);
nor U14623 (N_14623,N_14295,N_14257);
and U14624 (N_14624,N_14288,N_14337);
nand U14625 (N_14625,N_14279,N_14257);
nor U14626 (N_14626,N_14329,N_14403);
or U14627 (N_14627,N_14425,N_14255);
or U14628 (N_14628,N_14428,N_14435);
or U14629 (N_14629,N_14485,N_14262);
nand U14630 (N_14630,N_14330,N_14399);
and U14631 (N_14631,N_14292,N_14458);
nand U14632 (N_14632,N_14437,N_14297);
or U14633 (N_14633,N_14359,N_14458);
and U14634 (N_14634,N_14283,N_14327);
xor U14635 (N_14635,N_14269,N_14351);
nor U14636 (N_14636,N_14360,N_14380);
xnor U14637 (N_14637,N_14426,N_14277);
or U14638 (N_14638,N_14342,N_14402);
xnor U14639 (N_14639,N_14306,N_14499);
nor U14640 (N_14640,N_14322,N_14447);
nand U14641 (N_14641,N_14337,N_14315);
or U14642 (N_14642,N_14384,N_14350);
nor U14643 (N_14643,N_14394,N_14399);
xor U14644 (N_14644,N_14410,N_14311);
or U14645 (N_14645,N_14323,N_14395);
nor U14646 (N_14646,N_14368,N_14284);
and U14647 (N_14647,N_14459,N_14451);
and U14648 (N_14648,N_14264,N_14449);
nand U14649 (N_14649,N_14442,N_14387);
nor U14650 (N_14650,N_14412,N_14376);
nand U14651 (N_14651,N_14466,N_14344);
nand U14652 (N_14652,N_14305,N_14359);
or U14653 (N_14653,N_14280,N_14486);
nand U14654 (N_14654,N_14271,N_14348);
or U14655 (N_14655,N_14294,N_14393);
nor U14656 (N_14656,N_14377,N_14279);
or U14657 (N_14657,N_14379,N_14366);
xnor U14658 (N_14658,N_14398,N_14250);
xor U14659 (N_14659,N_14299,N_14335);
nor U14660 (N_14660,N_14260,N_14395);
nor U14661 (N_14661,N_14422,N_14484);
or U14662 (N_14662,N_14491,N_14316);
nor U14663 (N_14663,N_14460,N_14340);
nor U14664 (N_14664,N_14280,N_14361);
nand U14665 (N_14665,N_14410,N_14288);
nand U14666 (N_14666,N_14494,N_14334);
or U14667 (N_14667,N_14365,N_14413);
nand U14668 (N_14668,N_14298,N_14336);
nand U14669 (N_14669,N_14463,N_14493);
and U14670 (N_14670,N_14279,N_14310);
and U14671 (N_14671,N_14417,N_14496);
and U14672 (N_14672,N_14296,N_14250);
or U14673 (N_14673,N_14394,N_14266);
or U14674 (N_14674,N_14433,N_14295);
nor U14675 (N_14675,N_14492,N_14329);
nor U14676 (N_14676,N_14264,N_14476);
or U14677 (N_14677,N_14272,N_14342);
nor U14678 (N_14678,N_14266,N_14383);
or U14679 (N_14679,N_14495,N_14404);
or U14680 (N_14680,N_14309,N_14392);
nand U14681 (N_14681,N_14441,N_14466);
nand U14682 (N_14682,N_14307,N_14344);
and U14683 (N_14683,N_14482,N_14394);
and U14684 (N_14684,N_14285,N_14372);
xnor U14685 (N_14685,N_14264,N_14398);
or U14686 (N_14686,N_14461,N_14310);
and U14687 (N_14687,N_14327,N_14459);
nand U14688 (N_14688,N_14411,N_14402);
or U14689 (N_14689,N_14375,N_14282);
nor U14690 (N_14690,N_14399,N_14352);
nor U14691 (N_14691,N_14418,N_14396);
nor U14692 (N_14692,N_14263,N_14460);
xor U14693 (N_14693,N_14439,N_14336);
or U14694 (N_14694,N_14338,N_14291);
nand U14695 (N_14695,N_14250,N_14420);
or U14696 (N_14696,N_14287,N_14281);
xor U14697 (N_14697,N_14265,N_14308);
nor U14698 (N_14698,N_14320,N_14493);
nor U14699 (N_14699,N_14297,N_14296);
nand U14700 (N_14700,N_14451,N_14345);
nor U14701 (N_14701,N_14488,N_14276);
xnor U14702 (N_14702,N_14457,N_14326);
and U14703 (N_14703,N_14291,N_14406);
nor U14704 (N_14704,N_14409,N_14266);
nand U14705 (N_14705,N_14405,N_14364);
nand U14706 (N_14706,N_14436,N_14256);
nor U14707 (N_14707,N_14475,N_14252);
or U14708 (N_14708,N_14433,N_14486);
nand U14709 (N_14709,N_14271,N_14434);
or U14710 (N_14710,N_14389,N_14257);
and U14711 (N_14711,N_14468,N_14374);
and U14712 (N_14712,N_14400,N_14271);
nand U14713 (N_14713,N_14406,N_14260);
and U14714 (N_14714,N_14487,N_14396);
or U14715 (N_14715,N_14430,N_14371);
xnor U14716 (N_14716,N_14279,N_14485);
nor U14717 (N_14717,N_14439,N_14416);
xnor U14718 (N_14718,N_14469,N_14473);
nand U14719 (N_14719,N_14420,N_14258);
nand U14720 (N_14720,N_14471,N_14499);
xnor U14721 (N_14721,N_14319,N_14403);
nor U14722 (N_14722,N_14494,N_14338);
nand U14723 (N_14723,N_14313,N_14489);
nand U14724 (N_14724,N_14286,N_14328);
nand U14725 (N_14725,N_14359,N_14470);
nor U14726 (N_14726,N_14304,N_14432);
and U14727 (N_14727,N_14434,N_14297);
xor U14728 (N_14728,N_14253,N_14484);
nor U14729 (N_14729,N_14379,N_14296);
or U14730 (N_14730,N_14296,N_14421);
xnor U14731 (N_14731,N_14288,N_14476);
or U14732 (N_14732,N_14497,N_14266);
nand U14733 (N_14733,N_14475,N_14355);
and U14734 (N_14734,N_14363,N_14255);
or U14735 (N_14735,N_14262,N_14269);
nor U14736 (N_14736,N_14401,N_14435);
xor U14737 (N_14737,N_14333,N_14287);
nor U14738 (N_14738,N_14303,N_14262);
nand U14739 (N_14739,N_14369,N_14318);
or U14740 (N_14740,N_14486,N_14252);
or U14741 (N_14741,N_14333,N_14382);
and U14742 (N_14742,N_14474,N_14378);
xor U14743 (N_14743,N_14320,N_14298);
and U14744 (N_14744,N_14446,N_14431);
nor U14745 (N_14745,N_14267,N_14360);
or U14746 (N_14746,N_14399,N_14375);
nor U14747 (N_14747,N_14366,N_14417);
xnor U14748 (N_14748,N_14425,N_14304);
and U14749 (N_14749,N_14319,N_14397);
or U14750 (N_14750,N_14560,N_14614);
nor U14751 (N_14751,N_14592,N_14699);
xnor U14752 (N_14752,N_14654,N_14612);
or U14753 (N_14753,N_14594,N_14563);
nor U14754 (N_14754,N_14642,N_14696);
or U14755 (N_14755,N_14675,N_14747);
nand U14756 (N_14756,N_14655,N_14625);
xnor U14757 (N_14757,N_14704,N_14566);
nand U14758 (N_14758,N_14715,N_14637);
xnor U14759 (N_14759,N_14710,N_14690);
or U14760 (N_14760,N_14595,N_14590);
and U14761 (N_14761,N_14659,N_14722);
nand U14762 (N_14762,N_14674,N_14546);
or U14763 (N_14763,N_14733,N_14552);
or U14764 (N_14764,N_14725,N_14580);
and U14765 (N_14765,N_14677,N_14685);
nor U14766 (N_14766,N_14663,N_14573);
and U14767 (N_14767,N_14711,N_14660);
nor U14768 (N_14768,N_14603,N_14732);
nor U14769 (N_14769,N_14651,N_14537);
xor U14770 (N_14770,N_14652,N_14591);
or U14771 (N_14771,N_14565,N_14553);
xnor U14772 (N_14772,N_14728,N_14604);
and U14773 (N_14773,N_14631,N_14527);
nor U14774 (N_14774,N_14640,N_14549);
xor U14775 (N_14775,N_14542,N_14691);
or U14776 (N_14776,N_14567,N_14678);
nor U14777 (N_14777,N_14624,N_14586);
and U14778 (N_14778,N_14687,N_14582);
or U14779 (N_14779,N_14708,N_14541);
nor U14780 (N_14780,N_14576,N_14686);
nand U14781 (N_14781,N_14689,N_14589);
or U14782 (N_14782,N_14536,N_14627);
nor U14783 (N_14783,N_14745,N_14535);
nand U14784 (N_14784,N_14523,N_14608);
xnor U14785 (N_14785,N_14626,N_14701);
or U14786 (N_14786,N_14602,N_14670);
and U14787 (N_14787,N_14500,N_14524);
xnor U14788 (N_14788,N_14520,N_14676);
or U14789 (N_14789,N_14667,N_14507);
and U14790 (N_14790,N_14668,N_14746);
and U14791 (N_14791,N_14538,N_14714);
or U14792 (N_14792,N_14645,N_14620);
xor U14793 (N_14793,N_14719,N_14606);
nand U14794 (N_14794,N_14729,N_14703);
nor U14795 (N_14795,N_14564,N_14741);
nand U14796 (N_14796,N_14514,N_14706);
nor U14797 (N_14797,N_14610,N_14512);
or U14798 (N_14798,N_14616,N_14588);
nand U14799 (N_14799,N_14650,N_14611);
xnor U14800 (N_14800,N_14726,N_14695);
nand U14801 (N_14801,N_14705,N_14605);
xnor U14802 (N_14802,N_14697,N_14730);
xnor U14803 (N_14803,N_14662,N_14724);
nor U14804 (N_14804,N_14585,N_14548);
and U14805 (N_14805,N_14599,N_14510);
or U14806 (N_14806,N_14633,N_14601);
and U14807 (N_14807,N_14666,N_14643);
and U14808 (N_14808,N_14577,N_14698);
nor U14809 (N_14809,N_14684,N_14534);
or U14810 (N_14810,N_14634,N_14556);
nor U14811 (N_14811,N_14615,N_14657);
xnor U14812 (N_14812,N_14557,N_14607);
and U14813 (N_14813,N_14569,N_14628);
and U14814 (N_14814,N_14740,N_14579);
xnor U14815 (N_14815,N_14646,N_14570);
xor U14816 (N_14816,N_14683,N_14700);
and U14817 (N_14817,N_14707,N_14723);
or U14818 (N_14818,N_14644,N_14619);
nand U14819 (N_14819,N_14543,N_14638);
nand U14820 (N_14820,N_14734,N_14717);
nor U14821 (N_14821,N_14679,N_14735);
xnor U14822 (N_14822,N_14503,N_14571);
xnor U14823 (N_14823,N_14544,N_14506);
xor U14824 (N_14824,N_14575,N_14622);
and U14825 (N_14825,N_14727,N_14629);
or U14826 (N_14826,N_14748,N_14617);
nand U14827 (N_14827,N_14609,N_14702);
nor U14828 (N_14828,N_14501,N_14688);
nand U14829 (N_14829,N_14630,N_14531);
and U14830 (N_14830,N_14530,N_14641);
xor U14831 (N_14831,N_14692,N_14558);
xor U14832 (N_14832,N_14731,N_14739);
nor U14833 (N_14833,N_14508,N_14561);
xor U14834 (N_14834,N_14528,N_14712);
or U14835 (N_14835,N_14653,N_14521);
xor U14836 (N_14836,N_14647,N_14658);
and U14837 (N_14837,N_14533,N_14532);
nand U14838 (N_14838,N_14738,N_14562);
nand U14839 (N_14839,N_14713,N_14550);
nor U14840 (N_14840,N_14694,N_14509);
xor U14841 (N_14841,N_14572,N_14721);
or U14842 (N_14842,N_14736,N_14669);
and U14843 (N_14843,N_14587,N_14635);
or U14844 (N_14844,N_14639,N_14665);
nor U14845 (N_14845,N_14551,N_14596);
or U14846 (N_14846,N_14743,N_14681);
nand U14847 (N_14847,N_14554,N_14584);
xnor U14848 (N_14848,N_14597,N_14623);
and U14849 (N_14849,N_14522,N_14749);
nand U14850 (N_14850,N_14671,N_14519);
nor U14851 (N_14851,N_14648,N_14621);
and U14852 (N_14852,N_14716,N_14518);
or U14853 (N_14853,N_14525,N_14540);
or U14854 (N_14854,N_14547,N_14515);
xor U14855 (N_14855,N_14664,N_14632);
nand U14856 (N_14856,N_14709,N_14613);
and U14857 (N_14857,N_14559,N_14656);
nand U14858 (N_14858,N_14737,N_14578);
and U14859 (N_14859,N_14555,N_14720);
xnor U14860 (N_14860,N_14574,N_14568);
xnor U14861 (N_14861,N_14513,N_14545);
or U14862 (N_14862,N_14583,N_14511);
xor U14863 (N_14863,N_14529,N_14517);
nand U14864 (N_14864,N_14673,N_14718);
and U14865 (N_14865,N_14618,N_14744);
nand U14866 (N_14866,N_14598,N_14682);
nor U14867 (N_14867,N_14649,N_14636);
xnor U14868 (N_14868,N_14600,N_14742);
xor U14869 (N_14869,N_14526,N_14661);
and U14870 (N_14870,N_14581,N_14680);
nor U14871 (N_14871,N_14504,N_14593);
or U14872 (N_14872,N_14693,N_14516);
nand U14873 (N_14873,N_14672,N_14505);
nand U14874 (N_14874,N_14502,N_14539);
or U14875 (N_14875,N_14745,N_14655);
and U14876 (N_14876,N_14639,N_14572);
or U14877 (N_14877,N_14728,N_14748);
or U14878 (N_14878,N_14714,N_14723);
and U14879 (N_14879,N_14539,N_14622);
nor U14880 (N_14880,N_14599,N_14584);
xnor U14881 (N_14881,N_14655,N_14512);
and U14882 (N_14882,N_14605,N_14542);
nor U14883 (N_14883,N_14567,N_14529);
or U14884 (N_14884,N_14689,N_14500);
or U14885 (N_14885,N_14537,N_14633);
nor U14886 (N_14886,N_14534,N_14630);
or U14887 (N_14887,N_14711,N_14675);
and U14888 (N_14888,N_14718,N_14627);
nand U14889 (N_14889,N_14552,N_14696);
nand U14890 (N_14890,N_14574,N_14664);
nand U14891 (N_14891,N_14674,N_14655);
or U14892 (N_14892,N_14647,N_14629);
xor U14893 (N_14893,N_14689,N_14621);
nand U14894 (N_14894,N_14721,N_14557);
and U14895 (N_14895,N_14652,N_14679);
nand U14896 (N_14896,N_14674,N_14541);
and U14897 (N_14897,N_14578,N_14630);
xor U14898 (N_14898,N_14561,N_14677);
and U14899 (N_14899,N_14678,N_14528);
or U14900 (N_14900,N_14694,N_14654);
nor U14901 (N_14901,N_14639,N_14680);
and U14902 (N_14902,N_14507,N_14648);
xnor U14903 (N_14903,N_14701,N_14505);
nor U14904 (N_14904,N_14676,N_14736);
or U14905 (N_14905,N_14604,N_14558);
nor U14906 (N_14906,N_14535,N_14596);
nor U14907 (N_14907,N_14600,N_14700);
xnor U14908 (N_14908,N_14694,N_14679);
xnor U14909 (N_14909,N_14511,N_14671);
nor U14910 (N_14910,N_14581,N_14597);
and U14911 (N_14911,N_14665,N_14687);
and U14912 (N_14912,N_14663,N_14746);
nand U14913 (N_14913,N_14583,N_14564);
xor U14914 (N_14914,N_14512,N_14564);
xnor U14915 (N_14915,N_14639,N_14645);
nor U14916 (N_14916,N_14515,N_14612);
nor U14917 (N_14917,N_14530,N_14741);
or U14918 (N_14918,N_14698,N_14700);
or U14919 (N_14919,N_14695,N_14510);
xor U14920 (N_14920,N_14656,N_14600);
and U14921 (N_14921,N_14679,N_14686);
nor U14922 (N_14922,N_14583,N_14617);
nand U14923 (N_14923,N_14591,N_14511);
and U14924 (N_14924,N_14569,N_14514);
or U14925 (N_14925,N_14500,N_14647);
and U14926 (N_14926,N_14736,N_14702);
nand U14927 (N_14927,N_14675,N_14581);
xor U14928 (N_14928,N_14513,N_14625);
xor U14929 (N_14929,N_14583,N_14508);
and U14930 (N_14930,N_14536,N_14613);
and U14931 (N_14931,N_14747,N_14503);
nand U14932 (N_14932,N_14662,N_14670);
or U14933 (N_14933,N_14631,N_14720);
or U14934 (N_14934,N_14659,N_14724);
nor U14935 (N_14935,N_14664,N_14511);
nor U14936 (N_14936,N_14583,N_14737);
nand U14937 (N_14937,N_14553,N_14519);
xnor U14938 (N_14938,N_14673,N_14699);
nor U14939 (N_14939,N_14536,N_14537);
nand U14940 (N_14940,N_14657,N_14578);
xnor U14941 (N_14941,N_14549,N_14585);
nand U14942 (N_14942,N_14581,N_14632);
and U14943 (N_14943,N_14532,N_14616);
or U14944 (N_14944,N_14695,N_14647);
xor U14945 (N_14945,N_14725,N_14648);
nor U14946 (N_14946,N_14555,N_14543);
or U14947 (N_14947,N_14617,N_14747);
xor U14948 (N_14948,N_14702,N_14685);
xor U14949 (N_14949,N_14640,N_14554);
nand U14950 (N_14950,N_14590,N_14729);
nor U14951 (N_14951,N_14633,N_14517);
xor U14952 (N_14952,N_14738,N_14619);
or U14953 (N_14953,N_14679,N_14632);
nand U14954 (N_14954,N_14682,N_14706);
and U14955 (N_14955,N_14575,N_14745);
and U14956 (N_14956,N_14688,N_14596);
or U14957 (N_14957,N_14722,N_14591);
and U14958 (N_14958,N_14726,N_14715);
nor U14959 (N_14959,N_14747,N_14632);
nand U14960 (N_14960,N_14570,N_14571);
xor U14961 (N_14961,N_14727,N_14639);
nand U14962 (N_14962,N_14652,N_14642);
nand U14963 (N_14963,N_14600,N_14602);
nor U14964 (N_14964,N_14645,N_14619);
and U14965 (N_14965,N_14571,N_14713);
or U14966 (N_14966,N_14609,N_14706);
nor U14967 (N_14967,N_14686,N_14646);
xor U14968 (N_14968,N_14569,N_14732);
or U14969 (N_14969,N_14680,N_14747);
xnor U14970 (N_14970,N_14609,N_14538);
or U14971 (N_14971,N_14536,N_14727);
nand U14972 (N_14972,N_14500,N_14650);
nor U14973 (N_14973,N_14512,N_14653);
or U14974 (N_14974,N_14557,N_14559);
xnor U14975 (N_14975,N_14709,N_14660);
and U14976 (N_14976,N_14578,N_14563);
nand U14977 (N_14977,N_14541,N_14616);
nor U14978 (N_14978,N_14516,N_14564);
or U14979 (N_14979,N_14537,N_14649);
and U14980 (N_14980,N_14596,N_14711);
or U14981 (N_14981,N_14636,N_14541);
nand U14982 (N_14982,N_14651,N_14574);
xor U14983 (N_14983,N_14610,N_14603);
and U14984 (N_14984,N_14526,N_14704);
nor U14985 (N_14985,N_14669,N_14625);
or U14986 (N_14986,N_14644,N_14670);
and U14987 (N_14987,N_14560,N_14541);
nor U14988 (N_14988,N_14624,N_14505);
xnor U14989 (N_14989,N_14680,N_14686);
nand U14990 (N_14990,N_14594,N_14622);
xnor U14991 (N_14991,N_14745,N_14626);
nand U14992 (N_14992,N_14670,N_14608);
and U14993 (N_14993,N_14575,N_14586);
xor U14994 (N_14994,N_14682,N_14672);
and U14995 (N_14995,N_14643,N_14660);
or U14996 (N_14996,N_14677,N_14530);
nor U14997 (N_14997,N_14664,N_14603);
nand U14998 (N_14998,N_14551,N_14687);
nor U14999 (N_14999,N_14722,N_14543);
or U15000 (N_15000,N_14880,N_14919);
and U15001 (N_15001,N_14862,N_14937);
and U15002 (N_15002,N_14771,N_14797);
nor U15003 (N_15003,N_14851,N_14964);
xnor U15004 (N_15004,N_14801,N_14821);
nand U15005 (N_15005,N_14840,N_14828);
xor U15006 (N_15006,N_14894,N_14820);
nor U15007 (N_15007,N_14809,N_14825);
xor U15008 (N_15008,N_14767,N_14990);
nand U15009 (N_15009,N_14939,N_14757);
xnor U15010 (N_15010,N_14965,N_14921);
xnor U15011 (N_15011,N_14788,N_14804);
xnor U15012 (N_15012,N_14925,N_14835);
or U15013 (N_15013,N_14868,N_14899);
nor U15014 (N_15014,N_14764,N_14772);
nor U15015 (N_15015,N_14885,N_14783);
and U15016 (N_15016,N_14961,N_14762);
xor U15017 (N_15017,N_14908,N_14819);
nor U15018 (N_15018,N_14888,N_14910);
or U15019 (N_15019,N_14996,N_14860);
nor U15020 (N_15020,N_14847,N_14778);
nand U15021 (N_15021,N_14872,N_14988);
or U15022 (N_15022,N_14782,N_14857);
xor U15023 (N_15023,N_14922,N_14812);
or U15024 (N_15024,N_14861,N_14789);
nor U15025 (N_15025,N_14848,N_14844);
or U15026 (N_15026,N_14752,N_14995);
and U15027 (N_15027,N_14978,N_14979);
and U15028 (N_15028,N_14830,N_14900);
or U15029 (N_15029,N_14930,N_14909);
xnor U15030 (N_15030,N_14838,N_14896);
xnor U15031 (N_15031,N_14865,N_14799);
or U15032 (N_15032,N_14776,N_14854);
nand U15033 (N_15033,N_14766,N_14876);
and U15034 (N_15034,N_14756,N_14891);
and U15035 (N_15035,N_14955,N_14813);
xnor U15036 (N_15036,N_14892,N_14856);
xor U15037 (N_15037,N_14818,N_14785);
or U15038 (N_15038,N_14981,N_14758);
or U15039 (N_15039,N_14897,N_14986);
nor U15040 (N_15040,N_14786,N_14833);
xnor U15041 (N_15041,N_14927,N_14949);
or U15042 (N_15042,N_14884,N_14975);
or U15043 (N_15043,N_14887,N_14952);
or U15044 (N_15044,N_14878,N_14976);
xnor U15045 (N_15045,N_14882,N_14792);
or U15046 (N_15046,N_14841,N_14881);
nor U15047 (N_15047,N_14761,N_14956);
xor U15048 (N_15048,N_14817,N_14893);
nor U15049 (N_15049,N_14946,N_14911);
or U15050 (N_15050,N_14784,N_14794);
or U15051 (N_15051,N_14980,N_14824);
nor U15052 (N_15052,N_14943,N_14924);
or U15053 (N_15053,N_14855,N_14798);
xor U15054 (N_15054,N_14984,N_14929);
xnor U15055 (N_15055,N_14871,N_14879);
or U15056 (N_15056,N_14834,N_14950);
nand U15057 (N_15057,N_14886,N_14958);
xnor U15058 (N_15058,N_14829,N_14987);
or U15059 (N_15059,N_14999,N_14765);
and U15060 (N_15060,N_14906,N_14807);
xor U15061 (N_15061,N_14800,N_14836);
or U15062 (N_15062,N_14947,N_14864);
xor U15063 (N_15063,N_14944,N_14973);
xnor U15064 (N_15064,N_14839,N_14898);
xor U15065 (N_15065,N_14940,N_14763);
nand U15066 (N_15066,N_14935,N_14942);
or U15067 (N_15067,N_14938,N_14869);
nand U15068 (N_15068,N_14774,N_14993);
nor U15069 (N_15069,N_14905,N_14777);
and U15070 (N_15070,N_14810,N_14754);
and U15071 (N_15071,N_14904,N_14991);
and U15072 (N_15072,N_14793,N_14941);
or U15073 (N_15073,N_14843,N_14751);
xor U15074 (N_15074,N_14823,N_14780);
nor U15075 (N_15075,N_14842,N_14907);
or U15076 (N_15076,N_14971,N_14846);
and U15077 (N_15077,N_14870,N_14845);
and U15078 (N_15078,N_14805,N_14883);
nor U15079 (N_15079,N_14994,N_14877);
and U15080 (N_15080,N_14928,N_14796);
xor U15081 (N_15081,N_14853,N_14914);
or U15082 (N_15082,N_14859,N_14968);
nor U15083 (N_15083,N_14920,N_14989);
nand U15084 (N_15084,N_14811,N_14822);
and U15085 (N_15085,N_14969,N_14992);
nand U15086 (N_15086,N_14803,N_14760);
nor U15087 (N_15087,N_14874,N_14867);
nor U15088 (N_15088,N_14970,N_14997);
nor U15089 (N_15089,N_14790,N_14837);
xnor U15090 (N_15090,N_14959,N_14918);
nor U15091 (N_15091,N_14972,N_14982);
nand U15092 (N_15092,N_14933,N_14951);
nor U15093 (N_15093,N_14781,N_14948);
or U15094 (N_15094,N_14858,N_14917);
nand U15095 (N_15095,N_14974,N_14895);
nor U15096 (N_15096,N_14902,N_14998);
xnor U15097 (N_15097,N_14966,N_14945);
or U15098 (N_15098,N_14967,N_14889);
or U15099 (N_15099,N_14806,N_14901);
or U15100 (N_15100,N_14816,N_14983);
nand U15101 (N_15101,N_14923,N_14913);
and U15102 (N_15102,N_14768,N_14926);
and U15103 (N_15103,N_14808,N_14849);
or U15104 (N_15104,N_14773,N_14831);
nand U15105 (N_15105,N_14850,N_14775);
or U15106 (N_15106,N_14815,N_14875);
or U15107 (N_15107,N_14873,N_14934);
nand U15108 (N_15108,N_14814,N_14957);
nor U15109 (N_15109,N_14932,N_14770);
or U15110 (N_15110,N_14787,N_14753);
or U15111 (N_15111,N_14827,N_14903);
nand U15112 (N_15112,N_14759,N_14866);
or U15113 (N_15113,N_14791,N_14963);
xor U15114 (N_15114,N_14750,N_14912);
and U15115 (N_15115,N_14931,N_14977);
or U15116 (N_15116,N_14852,N_14802);
xor U15117 (N_15117,N_14962,N_14832);
xnor U15118 (N_15118,N_14985,N_14916);
nand U15119 (N_15119,N_14890,N_14863);
xnor U15120 (N_15120,N_14779,N_14795);
nand U15121 (N_15121,N_14915,N_14960);
nand U15122 (N_15122,N_14936,N_14953);
xor U15123 (N_15123,N_14954,N_14755);
nand U15124 (N_15124,N_14826,N_14769);
nor U15125 (N_15125,N_14763,N_14999);
nor U15126 (N_15126,N_14858,N_14883);
nor U15127 (N_15127,N_14769,N_14946);
xor U15128 (N_15128,N_14811,N_14917);
nand U15129 (N_15129,N_14966,N_14778);
and U15130 (N_15130,N_14824,N_14926);
xor U15131 (N_15131,N_14998,N_14931);
or U15132 (N_15132,N_14819,N_14766);
or U15133 (N_15133,N_14961,N_14840);
or U15134 (N_15134,N_14977,N_14795);
xor U15135 (N_15135,N_14759,N_14813);
nor U15136 (N_15136,N_14884,N_14836);
and U15137 (N_15137,N_14822,N_14964);
and U15138 (N_15138,N_14971,N_14888);
xor U15139 (N_15139,N_14792,N_14960);
nor U15140 (N_15140,N_14782,N_14875);
nor U15141 (N_15141,N_14768,N_14998);
nand U15142 (N_15142,N_14840,N_14772);
nand U15143 (N_15143,N_14769,N_14905);
or U15144 (N_15144,N_14934,N_14931);
nand U15145 (N_15145,N_14842,N_14829);
or U15146 (N_15146,N_14766,N_14810);
or U15147 (N_15147,N_14898,N_14993);
nand U15148 (N_15148,N_14931,N_14855);
xnor U15149 (N_15149,N_14838,N_14868);
nor U15150 (N_15150,N_14935,N_14807);
and U15151 (N_15151,N_14768,N_14757);
nor U15152 (N_15152,N_14862,N_14929);
nor U15153 (N_15153,N_14821,N_14828);
xnor U15154 (N_15154,N_14883,N_14880);
and U15155 (N_15155,N_14956,N_14983);
nor U15156 (N_15156,N_14958,N_14784);
nand U15157 (N_15157,N_14900,N_14817);
nor U15158 (N_15158,N_14976,N_14760);
and U15159 (N_15159,N_14836,N_14887);
nor U15160 (N_15160,N_14972,N_14938);
nor U15161 (N_15161,N_14903,N_14816);
and U15162 (N_15162,N_14832,N_14996);
xor U15163 (N_15163,N_14831,N_14769);
or U15164 (N_15164,N_14846,N_14978);
xnor U15165 (N_15165,N_14823,N_14827);
and U15166 (N_15166,N_14885,N_14776);
nor U15167 (N_15167,N_14947,N_14903);
nand U15168 (N_15168,N_14775,N_14882);
or U15169 (N_15169,N_14844,N_14765);
xor U15170 (N_15170,N_14830,N_14907);
and U15171 (N_15171,N_14956,N_14820);
xor U15172 (N_15172,N_14798,N_14936);
or U15173 (N_15173,N_14872,N_14909);
nor U15174 (N_15174,N_14868,N_14809);
xnor U15175 (N_15175,N_14868,N_14821);
and U15176 (N_15176,N_14928,N_14993);
or U15177 (N_15177,N_14820,N_14994);
nor U15178 (N_15178,N_14992,N_14812);
and U15179 (N_15179,N_14927,N_14862);
or U15180 (N_15180,N_14852,N_14905);
nand U15181 (N_15181,N_14972,N_14986);
or U15182 (N_15182,N_14894,N_14967);
nor U15183 (N_15183,N_14949,N_14926);
nor U15184 (N_15184,N_14954,N_14964);
and U15185 (N_15185,N_14761,N_14945);
or U15186 (N_15186,N_14947,N_14834);
xor U15187 (N_15187,N_14978,N_14896);
nand U15188 (N_15188,N_14873,N_14782);
and U15189 (N_15189,N_14879,N_14926);
and U15190 (N_15190,N_14870,N_14805);
and U15191 (N_15191,N_14966,N_14906);
xnor U15192 (N_15192,N_14854,N_14890);
nor U15193 (N_15193,N_14763,N_14820);
nor U15194 (N_15194,N_14916,N_14992);
xor U15195 (N_15195,N_14960,N_14914);
xor U15196 (N_15196,N_14926,N_14756);
or U15197 (N_15197,N_14769,N_14913);
nor U15198 (N_15198,N_14754,N_14853);
nand U15199 (N_15199,N_14827,N_14995);
nor U15200 (N_15200,N_14950,N_14837);
or U15201 (N_15201,N_14880,N_14860);
nor U15202 (N_15202,N_14814,N_14766);
nand U15203 (N_15203,N_14961,N_14911);
nor U15204 (N_15204,N_14859,N_14814);
xor U15205 (N_15205,N_14817,N_14854);
xnor U15206 (N_15206,N_14996,N_14961);
and U15207 (N_15207,N_14822,N_14887);
xnor U15208 (N_15208,N_14837,N_14936);
and U15209 (N_15209,N_14955,N_14989);
and U15210 (N_15210,N_14956,N_14917);
nor U15211 (N_15211,N_14892,N_14775);
or U15212 (N_15212,N_14894,N_14803);
or U15213 (N_15213,N_14873,N_14848);
nand U15214 (N_15214,N_14759,N_14815);
and U15215 (N_15215,N_14779,N_14822);
nor U15216 (N_15216,N_14830,N_14809);
nand U15217 (N_15217,N_14925,N_14850);
xor U15218 (N_15218,N_14918,N_14899);
and U15219 (N_15219,N_14840,N_14953);
nor U15220 (N_15220,N_14986,N_14898);
or U15221 (N_15221,N_14865,N_14808);
and U15222 (N_15222,N_14826,N_14870);
nand U15223 (N_15223,N_14843,N_14785);
nand U15224 (N_15224,N_14945,N_14968);
nand U15225 (N_15225,N_14950,N_14807);
nor U15226 (N_15226,N_14771,N_14810);
nand U15227 (N_15227,N_14800,N_14780);
nor U15228 (N_15228,N_14998,N_14838);
nor U15229 (N_15229,N_14825,N_14980);
nor U15230 (N_15230,N_14911,N_14910);
and U15231 (N_15231,N_14837,N_14904);
or U15232 (N_15232,N_14926,N_14829);
and U15233 (N_15233,N_14821,N_14896);
and U15234 (N_15234,N_14943,N_14856);
and U15235 (N_15235,N_14788,N_14812);
and U15236 (N_15236,N_14942,N_14869);
and U15237 (N_15237,N_14870,N_14892);
or U15238 (N_15238,N_14982,N_14813);
nor U15239 (N_15239,N_14810,N_14996);
or U15240 (N_15240,N_14830,N_14999);
and U15241 (N_15241,N_14912,N_14781);
nor U15242 (N_15242,N_14961,N_14780);
and U15243 (N_15243,N_14991,N_14997);
and U15244 (N_15244,N_14948,N_14855);
and U15245 (N_15245,N_14877,N_14875);
nand U15246 (N_15246,N_14885,N_14829);
xor U15247 (N_15247,N_14958,N_14893);
nor U15248 (N_15248,N_14917,N_14985);
and U15249 (N_15249,N_14792,N_14994);
and U15250 (N_15250,N_15078,N_15009);
nor U15251 (N_15251,N_15221,N_15226);
nand U15252 (N_15252,N_15244,N_15243);
nor U15253 (N_15253,N_15201,N_15174);
nand U15254 (N_15254,N_15228,N_15033);
or U15255 (N_15255,N_15072,N_15093);
and U15256 (N_15256,N_15246,N_15137);
and U15257 (N_15257,N_15238,N_15140);
xnor U15258 (N_15258,N_15068,N_15112);
xnor U15259 (N_15259,N_15036,N_15186);
nand U15260 (N_15260,N_15002,N_15180);
nor U15261 (N_15261,N_15222,N_15224);
xor U15262 (N_15262,N_15022,N_15011);
xnor U15263 (N_15263,N_15107,N_15015);
xnor U15264 (N_15264,N_15017,N_15166);
nand U15265 (N_15265,N_15132,N_15215);
nor U15266 (N_15266,N_15209,N_15050);
nor U15267 (N_15267,N_15001,N_15188);
and U15268 (N_15268,N_15207,N_15142);
and U15269 (N_15269,N_15067,N_15183);
and U15270 (N_15270,N_15032,N_15120);
and U15271 (N_15271,N_15006,N_15127);
or U15272 (N_15272,N_15125,N_15021);
or U15273 (N_15273,N_15028,N_15026);
or U15274 (N_15274,N_15233,N_15217);
nand U15275 (N_15275,N_15129,N_15141);
nor U15276 (N_15276,N_15152,N_15019);
nor U15277 (N_15277,N_15045,N_15220);
or U15278 (N_15278,N_15216,N_15063);
xnor U15279 (N_15279,N_15095,N_15155);
or U15280 (N_15280,N_15007,N_15108);
nand U15281 (N_15281,N_15071,N_15172);
nand U15282 (N_15282,N_15212,N_15008);
or U15283 (N_15283,N_15121,N_15013);
nor U15284 (N_15284,N_15074,N_15100);
xor U15285 (N_15285,N_15232,N_15133);
xor U15286 (N_15286,N_15211,N_15177);
nor U15287 (N_15287,N_15138,N_15065);
or U15288 (N_15288,N_15116,N_15139);
nand U15289 (N_15289,N_15047,N_15070);
nand U15290 (N_15290,N_15175,N_15210);
or U15291 (N_15291,N_15035,N_15016);
and U15292 (N_15292,N_15156,N_15241);
or U15293 (N_15293,N_15101,N_15029);
nor U15294 (N_15294,N_15130,N_15196);
nand U15295 (N_15295,N_15225,N_15235);
nor U15296 (N_15296,N_15136,N_15088);
or U15297 (N_15297,N_15128,N_15048);
nand U15298 (N_15298,N_15058,N_15126);
xnor U15299 (N_15299,N_15024,N_15134);
xor U15300 (N_15300,N_15004,N_15037);
or U15301 (N_15301,N_15176,N_15190);
nand U15302 (N_15302,N_15154,N_15161);
xor U15303 (N_15303,N_15194,N_15023);
nor U15304 (N_15304,N_15150,N_15147);
and U15305 (N_15305,N_15083,N_15199);
nor U15306 (N_15306,N_15079,N_15014);
nand U15307 (N_15307,N_15202,N_15169);
and U15308 (N_15308,N_15146,N_15030);
xor U15309 (N_15309,N_15005,N_15179);
nor U15310 (N_15310,N_15157,N_15165);
or U15311 (N_15311,N_15053,N_15034);
xnor U15312 (N_15312,N_15236,N_15086);
xnor U15313 (N_15313,N_15105,N_15055);
xnor U15314 (N_15314,N_15111,N_15203);
and U15315 (N_15315,N_15087,N_15227);
and U15316 (N_15316,N_15162,N_15187);
and U15317 (N_15317,N_15069,N_15064);
xnor U15318 (N_15318,N_15214,N_15230);
and U15319 (N_15319,N_15145,N_15171);
nor U15320 (N_15320,N_15041,N_15080);
xnor U15321 (N_15321,N_15153,N_15219);
nand U15322 (N_15322,N_15164,N_15191);
xor U15323 (N_15323,N_15184,N_15229);
nor U15324 (N_15324,N_15049,N_15038);
or U15325 (N_15325,N_15131,N_15239);
nand U15326 (N_15326,N_15018,N_15247);
xor U15327 (N_15327,N_15237,N_15081);
nor U15328 (N_15328,N_15102,N_15057);
nand U15329 (N_15329,N_15060,N_15000);
xnor U15330 (N_15330,N_15012,N_15066);
xor U15331 (N_15331,N_15059,N_15043);
or U15332 (N_15332,N_15151,N_15122);
or U15333 (N_15333,N_15052,N_15249);
nor U15334 (N_15334,N_15091,N_15182);
xor U15335 (N_15335,N_15109,N_15103);
and U15336 (N_15336,N_15046,N_15085);
and U15337 (N_15337,N_15010,N_15106);
xor U15338 (N_15338,N_15204,N_15084);
nor U15339 (N_15339,N_15123,N_15089);
nor U15340 (N_15340,N_15025,N_15143);
nand U15341 (N_15341,N_15223,N_15159);
and U15342 (N_15342,N_15124,N_15075);
and U15343 (N_15343,N_15094,N_15040);
nand U15344 (N_15344,N_15240,N_15118);
nand U15345 (N_15345,N_15189,N_15039);
nand U15346 (N_15346,N_15061,N_15242);
and U15347 (N_15347,N_15163,N_15206);
nor U15348 (N_15348,N_15020,N_15042);
and U15349 (N_15349,N_15099,N_15077);
and U15350 (N_15350,N_15027,N_15117);
nor U15351 (N_15351,N_15062,N_15082);
nand U15352 (N_15352,N_15245,N_15218);
or U15353 (N_15353,N_15092,N_15114);
nor U15354 (N_15354,N_15231,N_15110);
nand U15355 (N_15355,N_15168,N_15051);
and U15356 (N_15356,N_15090,N_15044);
or U15357 (N_15357,N_15208,N_15003);
xnor U15358 (N_15358,N_15031,N_15054);
or U15359 (N_15359,N_15098,N_15158);
and U15360 (N_15360,N_15119,N_15144);
nand U15361 (N_15361,N_15248,N_15097);
and U15362 (N_15362,N_15076,N_15167);
xor U15363 (N_15363,N_15160,N_15205);
xnor U15364 (N_15364,N_15113,N_15192);
xnor U15365 (N_15365,N_15104,N_15200);
or U15366 (N_15366,N_15213,N_15115);
and U15367 (N_15367,N_15198,N_15170);
and U15368 (N_15368,N_15135,N_15181);
nor U15369 (N_15369,N_15148,N_15178);
or U15370 (N_15370,N_15149,N_15197);
or U15371 (N_15371,N_15185,N_15073);
nand U15372 (N_15372,N_15195,N_15096);
nand U15373 (N_15373,N_15173,N_15056);
nor U15374 (N_15374,N_15193,N_15234);
and U15375 (N_15375,N_15114,N_15233);
nor U15376 (N_15376,N_15044,N_15234);
or U15377 (N_15377,N_15220,N_15243);
nand U15378 (N_15378,N_15194,N_15143);
nor U15379 (N_15379,N_15166,N_15052);
or U15380 (N_15380,N_15107,N_15082);
nand U15381 (N_15381,N_15127,N_15135);
nand U15382 (N_15382,N_15113,N_15164);
xnor U15383 (N_15383,N_15217,N_15135);
xnor U15384 (N_15384,N_15058,N_15091);
xor U15385 (N_15385,N_15155,N_15120);
nor U15386 (N_15386,N_15034,N_15113);
nor U15387 (N_15387,N_15012,N_15233);
and U15388 (N_15388,N_15065,N_15223);
nand U15389 (N_15389,N_15018,N_15145);
and U15390 (N_15390,N_15185,N_15202);
xnor U15391 (N_15391,N_15076,N_15028);
xor U15392 (N_15392,N_15022,N_15210);
nor U15393 (N_15393,N_15182,N_15022);
or U15394 (N_15394,N_15205,N_15005);
nand U15395 (N_15395,N_15126,N_15051);
or U15396 (N_15396,N_15048,N_15081);
xnor U15397 (N_15397,N_15169,N_15004);
nor U15398 (N_15398,N_15236,N_15143);
nand U15399 (N_15399,N_15115,N_15078);
nor U15400 (N_15400,N_15223,N_15197);
or U15401 (N_15401,N_15208,N_15035);
or U15402 (N_15402,N_15155,N_15144);
nand U15403 (N_15403,N_15137,N_15093);
and U15404 (N_15404,N_15009,N_15186);
or U15405 (N_15405,N_15199,N_15192);
nor U15406 (N_15406,N_15067,N_15162);
nor U15407 (N_15407,N_15000,N_15006);
and U15408 (N_15408,N_15039,N_15056);
or U15409 (N_15409,N_15123,N_15121);
and U15410 (N_15410,N_15002,N_15118);
and U15411 (N_15411,N_15221,N_15136);
nor U15412 (N_15412,N_15224,N_15177);
and U15413 (N_15413,N_15014,N_15091);
nor U15414 (N_15414,N_15197,N_15186);
nand U15415 (N_15415,N_15043,N_15208);
nand U15416 (N_15416,N_15109,N_15026);
nor U15417 (N_15417,N_15017,N_15007);
xor U15418 (N_15418,N_15042,N_15155);
nor U15419 (N_15419,N_15119,N_15137);
nor U15420 (N_15420,N_15063,N_15215);
and U15421 (N_15421,N_15106,N_15194);
nand U15422 (N_15422,N_15145,N_15169);
nand U15423 (N_15423,N_15060,N_15124);
xor U15424 (N_15424,N_15195,N_15025);
nor U15425 (N_15425,N_15195,N_15033);
nand U15426 (N_15426,N_15172,N_15049);
nor U15427 (N_15427,N_15145,N_15111);
xnor U15428 (N_15428,N_15003,N_15170);
nand U15429 (N_15429,N_15091,N_15111);
xnor U15430 (N_15430,N_15183,N_15210);
nor U15431 (N_15431,N_15144,N_15093);
nand U15432 (N_15432,N_15065,N_15219);
nor U15433 (N_15433,N_15222,N_15199);
xnor U15434 (N_15434,N_15237,N_15114);
nor U15435 (N_15435,N_15247,N_15132);
and U15436 (N_15436,N_15021,N_15230);
xor U15437 (N_15437,N_15236,N_15062);
xor U15438 (N_15438,N_15219,N_15003);
or U15439 (N_15439,N_15234,N_15214);
or U15440 (N_15440,N_15220,N_15124);
and U15441 (N_15441,N_15090,N_15202);
xnor U15442 (N_15442,N_15027,N_15188);
or U15443 (N_15443,N_15222,N_15225);
and U15444 (N_15444,N_15231,N_15247);
nand U15445 (N_15445,N_15111,N_15081);
or U15446 (N_15446,N_15130,N_15099);
or U15447 (N_15447,N_15153,N_15122);
and U15448 (N_15448,N_15081,N_15202);
or U15449 (N_15449,N_15152,N_15149);
nand U15450 (N_15450,N_15211,N_15022);
nand U15451 (N_15451,N_15100,N_15112);
or U15452 (N_15452,N_15064,N_15131);
xnor U15453 (N_15453,N_15167,N_15145);
and U15454 (N_15454,N_15085,N_15200);
and U15455 (N_15455,N_15022,N_15227);
nand U15456 (N_15456,N_15126,N_15097);
nand U15457 (N_15457,N_15216,N_15046);
nor U15458 (N_15458,N_15044,N_15176);
xnor U15459 (N_15459,N_15111,N_15004);
or U15460 (N_15460,N_15021,N_15216);
or U15461 (N_15461,N_15004,N_15120);
nor U15462 (N_15462,N_15066,N_15001);
and U15463 (N_15463,N_15097,N_15196);
nor U15464 (N_15464,N_15088,N_15014);
xnor U15465 (N_15465,N_15036,N_15215);
nor U15466 (N_15466,N_15061,N_15105);
xor U15467 (N_15467,N_15186,N_15249);
nand U15468 (N_15468,N_15034,N_15005);
nor U15469 (N_15469,N_15140,N_15159);
and U15470 (N_15470,N_15173,N_15046);
and U15471 (N_15471,N_15026,N_15180);
xnor U15472 (N_15472,N_15184,N_15242);
or U15473 (N_15473,N_15130,N_15156);
nand U15474 (N_15474,N_15210,N_15139);
nand U15475 (N_15475,N_15157,N_15232);
and U15476 (N_15476,N_15002,N_15185);
and U15477 (N_15477,N_15228,N_15200);
xnor U15478 (N_15478,N_15063,N_15164);
nor U15479 (N_15479,N_15116,N_15107);
and U15480 (N_15480,N_15159,N_15013);
nor U15481 (N_15481,N_15214,N_15175);
xor U15482 (N_15482,N_15195,N_15082);
xnor U15483 (N_15483,N_15079,N_15217);
xnor U15484 (N_15484,N_15145,N_15217);
xor U15485 (N_15485,N_15033,N_15186);
or U15486 (N_15486,N_15192,N_15241);
nor U15487 (N_15487,N_15110,N_15184);
nand U15488 (N_15488,N_15184,N_15157);
nand U15489 (N_15489,N_15150,N_15044);
nand U15490 (N_15490,N_15238,N_15170);
or U15491 (N_15491,N_15177,N_15039);
or U15492 (N_15492,N_15126,N_15172);
or U15493 (N_15493,N_15213,N_15186);
and U15494 (N_15494,N_15224,N_15065);
nor U15495 (N_15495,N_15041,N_15038);
nand U15496 (N_15496,N_15245,N_15180);
nand U15497 (N_15497,N_15025,N_15190);
nand U15498 (N_15498,N_15246,N_15013);
xor U15499 (N_15499,N_15081,N_15103);
xor U15500 (N_15500,N_15294,N_15303);
and U15501 (N_15501,N_15401,N_15426);
xor U15502 (N_15502,N_15306,N_15457);
or U15503 (N_15503,N_15353,N_15268);
nor U15504 (N_15504,N_15283,N_15312);
and U15505 (N_15505,N_15474,N_15298);
xor U15506 (N_15506,N_15320,N_15388);
xor U15507 (N_15507,N_15321,N_15275);
nor U15508 (N_15508,N_15455,N_15450);
or U15509 (N_15509,N_15389,N_15487);
nand U15510 (N_15510,N_15324,N_15423);
xor U15511 (N_15511,N_15266,N_15296);
nor U15512 (N_15512,N_15251,N_15322);
nand U15513 (N_15513,N_15292,N_15465);
nor U15514 (N_15514,N_15365,N_15383);
and U15515 (N_15515,N_15341,N_15333);
or U15516 (N_15516,N_15387,N_15259);
and U15517 (N_15517,N_15364,N_15472);
nor U15518 (N_15518,N_15462,N_15253);
and U15519 (N_15519,N_15284,N_15269);
and U15520 (N_15520,N_15398,N_15456);
or U15521 (N_15521,N_15489,N_15278);
or U15522 (N_15522,N_15488,N_15461);
nor U15523 (N_15523,N_15434,N_15481);
xnor U15524 (N_15524,N_15412,N_15262);
or U15525 (N_15525,N_15289,N_15492);
and U15526 (N_15526,N_15453,N_15404);
nand U15527 (N_15527,N_15413,N_15368);
xnor U15528 (N_15528,N_15411,N_15491);
nor U15529 (N_15529,N_15495,N_15441);
and U15530 (N_15530,N_15343,N_15367);
or U15531 (N_15531,N_15486,N_15342);
or U15532 (N_15532,N_15274,N_15490);
xor U15533 (N_15533,N_15277,N_15280);
or U15534 (N_15534,N_15422,N_15340);
and U15535 (N_15535,N_15309,N_15403);
nor U15536 (N_15536,N_15396,N_15399);
xor U15537 (N_15537,N_15362,N_15313);
nand U15538 (N_15538,N_15419,N_15265);
and U15539 (N_15539,N_15406,N_15250);
xor U15540 (N_15540,N_15372,N_15327);
or U15541 (N_15541,N_15408,N_15484);
xnor U15542 (N_15542,N_15479,N_15332);
or U15543 (N_15543,N_15318,N_15302);
nand U15544 (N_15544,N_15410,N_15392);
and U15545 (N_15545,N_15390,N_15430);
nor U15546 (N_15546,N_15347,N_15371);
and U15547 (N_15547,N_15291,N_15370);
xnor U15548 (N_15548,N_15311,N_15409);
or U15549 (N_15549,N_15494,N_15316);
nor U15550 (N_15550,N_15468,N_15308);
and U15551 (N_15551,N_15394,N_15255);
xor U15552 (N_15552,N_15382,N_15357);
nand U15553 (N_15553,N_15436,N_15256);
or U15554 (N_15554,N_15446,N_15286);
xnor U15555 (N_15555,N_15452,N_15325);
nand U15556 (N_15556,N_15381,N_15483);
nor U15557 (N_15557,N_15421,N_15431);
or U15558 (N_15558,N_15281,N_15393);
xor U15559 (N_15559,N_15477,N_15470);
or U15560 (N_15560,N_15405,N_15380);
or U15561 (N_15561,N_15448,N_15307);
or U15562 (N_15562,N_15336,N_15438);
xor U15563 (N_15563,N_15300,N_15493);
or U15564 (N_15564,N_15440,N_15498);
xor U15565 (N_15565,N_15375,N_15350);
or U15566 (N_15566,N_15270,N_15485);
or U15567 (N_15567,N_15264,N_15334);
xor U15568 (N_15568,N_15445,N_15359);
or U15569 (N_15569,N_15499,N_15254);
xnor U15570 (N_15570,N_15418,N_15315);
nand U15571 (N_15571,N_15271,N_15344);
nand U15572 (N_15572,N_15310,N_15444);
nor U15573 (N_15573,N_15349,N_15424);
nand U15574 (N_15574,N_15263,N_15348);
and U15575 (N_15575,N_15433,N_15317);
nand U15576 (N_15576,N_15345,N_15304);
nor U15577 (N_15577,N_15369,N_15337);
and U15578 (N_15578,N_15319,N_15338);
nand U15579 (N_15579,N_15476,N_15361);
nor U15580 (N_15580,N_15407,N_15473);
nand U15581 (N_15581,N_15385,N_15466);
nor U15582 (N_15582,N_15329,N_15257);
xnor U15583 (N_15583,N_15273,N_15429);
and U15584 (N_15584,N_15414,N_15443);
nor U15585 (N_15585,N_15425,N_15467);
or U15586 (N_15586,N_15460,N_15469);
xor U15587 (N_15587,N_15261,N_15285);
or U15588 (N_15588,N_15282,N_15288);
nor U15589 (N_15589,N_15415,N_15427);
and U15590 (N_15590,N_15397,N_15475);
nor U15591 (N_15591,N_15355,N_15295);
or U15592 (N_15592,N_15379,N_15260);
or U15593 (N_15593,N_15471,N_15420);
xnor U15594 (N_15594,N_15299,N_15352);
or U15595 (N_15595,N_15331,N_15463);
nand U15596 (N_15596,N_15305,N_15416);
nor U15597 (N_15597,N_15330,N_15358);
and U15598 (N_15598,N_15464,N_15326);
nand U15599 (N_15599,N_15354,N_15439);
nand U15600 (N_15600,N_15293,N_15314);
xor U15601 (N_15601,N_15432,N_15451);
xor U15602 (N_15602,N_15374,N_15346);
xnor U15603 (N_15603,N_15378,N_15454);
nor U15604 (N_15604,N_15391,N_15335);
nor U15605 (N_15605,N_15458,N_15417);
nor U15606 (N_15606,N_15386,N_15384);
or U15607 (N_15607,N_15482,N_15287);
and U15608 (N_15608,N_15279,N_15323);
or U15609 (N_15609,N_15290,N_15328);
nor U15610 (N_15610,N_15297,N_15435);
and U15611 (N_15611,N_15360,N_15497);
and U15612 (N_15612,N_15437,N_15478);
or U15613 (N_15613,N_15376,N_15373);
nand U15614 (N_15614,N_15447,N_15449);
xor U15615 (N_15615,N_15366,N_15395);
nand U15616 (N_15616,N_15459,N_15267);
or U15617 (N_15617,N_15428,N_15356);
xor U15618 (N_15618,N_15400,N_15442);
nand U15619 (N_15619,N_15276,N_15402);
xnor U15620 (N_15620,N_15272,N_15258);
xor U15621 (N_15621,N_15301,N_15351);
or U15622 (N_15622,N_15252,N_15339);
nand U15623 (N_15623,N_15363,N_15480);
or U15624 (N_15624,N_15496,N_15377);
nand U15625 (N_15625,N_15253,N_15352);
or U15626 (N_15626,N_15252,N_15413);
and U15627 (N_15627,N_15378,N_15393);
xnor U15628 (N_15628,N_15324,N_15414);
and U15629 (N_15629,N_15414,N_15264);
and U15630 (N_15630,N_15265,N_15286);
xor U15631 (N_15631,N_15460,N_15465);
or U15632 (N_15632,N_15318,N_15253);
nor U15633 (N_15633,N_15442,N_15355);
nand U15634 (N_15634,N_15455,N_15288);
nor U15635 (N_15635,N_15328,N_15459);
nand U15636 (N_15636,N_15489,N_15384);
nor U15637 (N_15637,N_15438,N_15481);
xnor U15638 (N_15638,N_15378,N_15315);
xor U15639 (N_15639,N_15447,N_15257);
nand U15640 (N_15640,N_15273,N_15410);
and U15641 (N_15641,N_15255,N_15449);
nand U15642 (N_15642,N_15417,N_15473);
and U15643 (N_15643,N_15489,N_15298);
and U15644 (N_15644,N_15496,N_15413);
xor U15645 (N_15645,N_15394,N_15402);
nor U15646 (N_15646,N_15499,N_15365);
or U15647 (N_15647,N_15410,N_15372);
or U15648 (N_15648,N_15380,N_15300);
nand U15649 (N_15649,N_15353,N_15459);
nor U15650 (N_15650,N_15450,N_15438);
nor U15651 (N_15651,N_15467,N_15473);
nor U15652 (N_15652,N_15424,N_15310);
or U15653 (N_15653,N_15409,N_15469);
nand U15654 (N_15654,N_15380,N_15495);
nand U15655 (N_15655,N_15319,N_15408);
nor U15656 (N_15656,N_15411,N_15481);
nor U15657 (N_15657,N_15499,N_15329);
or U15658 (N_15658,N_15481,N_15329);
nor U15659 (N_15659,N_15268,N_15424);
xor U15660 (N_15660,N_15264,N_15492);
or U15661 (N_15661,N_15392,N_15295);
or U15662 (N_15662,N_15300,N_15392);
xnor U15663 (N_15663,N_15495,N_15349);
nand U15664 (N_15664,N_15291,N_15340);
or U15665 (N_15665,N_15310,N_15301);
xor U15666 (N_15666,N_15337,N_15438);
xor U15667 (N_15667,N_15461,N_15269);
or U15668 (N_15668,N_15424,N_15302);
nor U15669 (N_15669,N_15486,N_15437);
nor U15670 (N_15670,N_15413,N_15294);
xnor U15671 (N_15671,N_15364,N_15320);
and U15672 (N_15672,N_15317,N_15250);
nand U15673 (N_15673,N_15312,N_15438);
nor U15674 (N_15674,N_15325,N_15261);
nor U15675 (N_15675,N_15489,N_15365);
xnor U15676 (N_15676,N_15450,N_15269);
nor U15677 (N_15677,N_15380,N_15330);
xnor U15678 (N_15678,N_15489,N_15479);
and U15679 (N_15679,N_15486,N_15485);
nand U15680 (N_15680,N_15364,N_15259);
nor U15681 (N_15681,N_15398,N_15325);
nor U15682 (N_15682,N_15314,N_15451);
and U15683 (N_15683,N_15344,N_15457);
nor U15684 (N_15684,N_15304,N_15317);
and U15685 (N_15685,N_15367,N_15269);
or U15686 (N_15686,N_15398,N_15444);
nand U15687 (N_15687,N_15494,N_15288);
xnor U15688 (N_15688,N_15395,N_15384);
and U15689 (N_15689,N_15305,N_15485);
nand U15690 (N_15690,N_15412,N_15292);
or U15691 (N_15691,N_15354,N_15491);
nor U15692 (N_15692,N_15281,N_15459);
nand U15693 (N_15693,N_15357,N_15475);
xnor U15694 (N_15694,N_15315,N_15362);
or U15695 (N_15695,N_15253,N_15307);
and U15696 (N_15696,N_15348,N_15337);
nand U15697 (N_15697,N_15337,N_15437);
nor U15698 (N_15698,N_15367,N_15270);
nor U15699 (N_15699,N_15428,N_15474);
nor U15700 (N_15700,N_15316,N_15260);
and U15701 (N_15701,N_15418,N_15333);
xor U15702 (N_15702,N_15483,N_15374);
nand U15703 (N_15703,N_15329,N_15283);
and U15704 (N_15704,N_15445,N_15437);
xor U15705 (N_15705,N_15388,N_15275);
and U15706 (N_15706,N_15282,N_15325);
and U15707 (N_15707,N_15319,N_15300);
nor U15708 (N_15708,N_15447,N_15264);
and U15709 (N_15709,N_15445,N_15323);
nor U15710 (N_15710,N_15441,N_15267);
xnor U15711 (N_15711,N_15346,N_15385);
xor U15712 (N_15712,N_15333,N_15424);
and U15713 (N_15713,N_15343,N_15489);
xnor U15714 (N_15714,N_15351,N_15427);
or U15715 (N_15715,N_15423,N_15358);
and U15716 (N_15716,N_15371,N_15285);
or U15717 (N_15717,N_15433,N_15473);
or U15718 (N_15718,N_15255,N_15252);
or U15719 (N_15719,N_15423,N_15469);
nor U15720 (N_15720,N_15479,N_15259);
and U15721 (N_15721,N_15353,N_15483);
and U15722 (N_15722,N_15434,N_15354);
nor U15723 (N_15723,N_15465,N_15462);
xnor U15724 (N_15724,N_15341,N_15257);
or U15725 (N_15725,N_15456,N_15251);
or U15726 (N_15726,N_15359,N_15486);
xnor U15727 (N_15727,N_15341,N_15433);
or U15728 (N_15728,N_15350,N_15445);
nand U15729 (N_15729,N_15311,N_15478);
or U15730 (N_15730,N_15449,N_15287);
nand U15731 (N_15731,N_15258,N_15259);
nor U15732 (N_15732,N_15404,N_15264);
nand U15733 (N_15733,N_15337,N_15486);
nor U15734 (N_15734,N_15494,N_15456);
nor U15735 (N_15735,N_15272,N_15338);
or U15736 (N_15736,N_15280,N_15357);
xnor U15737 (N_15737,N_15381,N_15331);
nand U15738 (N_15738,N_15488,N_15499);
nand U15739 (N_15739,N_15343,N_15307);
nor U15740 (N_15740,N_15398,N_15304);
nor U15741 (N_15741,N_15319,N_15317);
nand U15742 (N_15742,N_15313,N_15383);
nor U15743 (N_15743,N_15491,N_15251);
or U15744 (N_15744,N_15256,N_15439);
or U15745 (N_15745,N_15483,N_15438);
or U15746 (N_15746,N_15428,N_15388);
or U15747 (N_15747,N_15260,N_15471);
or U15748 (N_15748,N_15480,N_15337);
nor U15749 (N_15749,N_15431,N_15367);
or U15750 (N_15750,N_15715,N_15500);
and U15751 (N_15751,N_15693,N_15584);
nand U15752 (N_15752,N_15610,N_15688);
and U15753 (N_15753,N_15506,N_15678);
or U15754 (N_15754,N_15621,N_15525);
nand U15755 (N_15755,N_15647,N_15734);
nor U15756 (N_15756,N_15563,N_15707);
and U15757 (N_15757,N_15583,N_15512);
xor U15758 (N_15758,N_15710,N_15546);
nor U15759 (N_15759,N_15545,N_15503);
and U15760 (N_15760,N_15703,N_15656);
xor U15761 (N_15761,N_15560,N_15694);
nand U15762 (N_15762,N_15697,N_15681);
or U15763 (N_15763,N_15590,N_15632);
or U15764 (N_15764,N_15711,N_15675);
nand U15765 (N_15765,N_15730,N_15731);
xor U15766 (N_15766,N_15745,N_15660);
and U15767 (N_15767,N_15573,N_15741);
or U15768 (N_15768,N_15670,N_15700);
xor U15769 (N_15769,N_15637,N_15702);
nand U15770 (N_15770,N_15732,N_15722);
nand U15771 (N_15771,N_15586,N_15704);
nand U15772 (N_15772,N_15646,N_15591);
nand U15773 (N_15773,N_15508,N_15562);
or U15774 (N_15774,N_15581,N_15659);
and U15775 (N_15775,N_15520,N_15542);
and U15776 (N_15776,N_15534,N_15528);
nor U15777 (N_15777,N_15565,N_15532);
nand U15778 (N_15778,N_15739,N_15684);
xor U15779 (N_15779,N_15719,N_15634);
or U15780 (N_15780,N_15686,N_15547);
and U15781 (N_15781,N_15533,N_15747);
nor U15782 (N_15782,N_15605,N_15724);
and U15783 (N_15783,N_15594,N_15705);
nand U15784 (N_15784,N_15564,N_15645);
or U15785 (N_15785,N_15648,N_15517);
xor U15786 (N_15786,N_15539,N_15582);
and U15787 (N_15787,N_15555,N_15602);
nand U15788 (N_15788,N_15653,N_15623);
nor U15789 (N_15789,N_15550,N_15527);
and U15790 (N_15790,N_15514,N_15551);
nor U15791 (N_15791,N_15652,N_15580);
nor U15792 (N_15792,N_15570,N_15598);
nand U15793 (N_15793,N_15556,N_15682);
nand U15794 (N_15794,N_15510,N_15631);
nor U15795 (N_15795,N_15740,N_15701);
xnor U15796 (N_15796,N_15725,N_15540);
or U15797 (N_15797,N_15572,N_15604);
nor U15798 (N_15798,N_15625,N_15685);
and U15799 (N_15799,N_15742,N_15609);
nand U15800 (N_15800,N_15672,N_15668);
and U15801 (N_15801,N_15511,N_15733);
nor U15802 (N_15802,N_15683,N_15595);
and U15803 (N_15803,N_15744,N_15530);
and U15804 (N_15804,N_15679,N_15577);
nor U15805 (N_15805,N_15677,N_15620);
nand U15806 (N_15806,N_15669,N_15735);
or U15807 (N_15807,N_15579,N_15709);
or U15808 (N_15808,N_15662,N_15521);
nand U15809 (N_15809,N_15665,N_15522);
nand U15810 (N_15810,N_15553,N_15504);
and U15811 (N_15811,N_15596,N_15619);
xor U15812 (N_15812,N_15606,N_15746);
or U15813 (N_15813,N_15657,N_15629);
nor U15814 (N_15814,N_15633,N_15699);
xor U15815 (N_15815,N_15708,N_15654);
or U15816 (N_15816,N_15554,N_15676);
nand U15817 (N_15817,N_15558,N_15523);
nand U15818 (N_15818,N_15592,N_15666);
xnor U15819 (N_15819,N_15738,N_15526);
and U15820 (N_15820,N_15593,N_15636);
or U15821 (N_15821,N_15529,N_15513);
nand U15822 (N_15822,N_15588,N_15635);
xor U15823 (N_15823,N_15651,N_15664);
or U15824 (N_15824,N_15640,N_15541);
and U15825 (N_15825,N_15568,N_15509);
nor U15826 (N_15826,N_15507,N_15691);
or U15827 (N_15827,N_15566,N_15658);
xor U15828 (N_15828,N_15692,N_15721);
nor U15829 (N_15829,N_15505,N_15650);
and U15830 (N_15830,N_15608,N_15718);
or U15831 (N_15831,N_15663,N_15728);
or U15832 (N_15832,N_15627,N_15515);
xnor U15833 (N_15833,N_15624,N_15743);
nor U15834 (N_15834,N_15599,N_15649);
nor U15835 (N_15835,N_15616,N_15706);
nand U15836 (N_15836,N_15690,N_15537);
xnor U15837 (N_15837,N_15671,N_15680);
or U15838 (N_15838,N_15587,N_15617);
and U15839 (N_15839,N_15614,N_15536);
nand U15840 (N_15840,N_15687,N_15712);
and U15841 (N_15841,N_15576,N_15524);
nor U15842 (N_15842,N_15717,N_15737);
nor U15843 (N_15843,N_15611,N_15585);
nand U15844 (N_15844,N_15552,N_15531);
nand U15845 (N_15845,N_15544,N_15689);
nor U15846 (N_15846,N_15502,N_15716);
nand U15847 (N_15847,N_15575,N_15727);
and U15848 (N_15848,N_15748,N_15622);
nor U15849 (N_15849,N_15600,N_15538);
nand U15850 (N_15850,N_15667,N_15661);
xor U15851 (N_15851,N_15557,N_15628);
xor U15852 (N_15852,N_15641,N_15639);
nor U15853 (N_15853,N_15535,N_15726);
xor U15854 (N_15854,N_15749,N_15601);
xnor U15855 (N_15855,N_15518,N_15695);
xnor U15856 (N_15856,N_15613,N_15644);
nor U15857 (N_15857,N_15638,N_15607);
or U15858 (N_15858,N_15597,N_15578);
or U15859 (N_15859,N_15655,N_15720);
nor U15860 (N_15860,N_15589,N_15519);
xnor U15861 (N_15861,N_15626,N_15574);
nor U15862 (N_15862,N_15729,N_15674);
nor U15863 (N_15863,N_15696,N_15603);
or U15864 (N_15864,N_15516,N_15618);
nor U15865 (N_15865,N_15571,N_15714);
or U15866 (N_15866,N_15561,N_15713);
xnor U15867 (N_15867,N_15567,N_15736);
and U15868 (N_15868,N_15673,N_15643);
and U15869 (N_15869,N_15501,N_15612);
xor U15870 (N_15870,N_15569,N_15642);
or U15871 (N_15871,N_15559,N_15615);
nor U15872 (N_15872,N_15698,N_15548);
nor U15873 (N_15873,N_15543,N_15723);
nand U15874 (N_15874,N_15549,N_15630);
or U15875 (N_15875,N_15583,N_15521);
or U15876 (N_15876,N_15547,N_15517);
or U15877 (N_15877,N_15603,N_15609);
nor U15878 (N_15878,N_15550,N_15610);
and U15879 (N_15879,N_15679,N_15605);
xnor U15880 (N_15880,N_15532,N_15611);
and U15881 (N_15881,N_15711,N_15633);
nor U15882 (N_15882,N_15631,N_15645);
nor U15883 (N_15883,N_15658,N_15579);
nand U15884 (N_15884,N_15616,N_15724);
nor U15885 (N_15885,N_15509,N_15667);
xnor U15886 (N_15886,N_15675,N_15655);
nand U15887 (N_15887,N_15585,N_15543);
nand U15888 (N_15888,N_15708,N_15522);
and U15889 (N_15889,N_15705,N_15669);
or U15890 (N_15890,N_15595,N_15628);
and U15891 (N_15891,N_15635,N_15625);
or U15892 (N_15892,N_15514,N_15710);
and U15893 (N_15893,N_15575,N_15518);
and U15894 (N_15894,N_15617,N_15725);
and U15895 (N_15895,N_15713,N_15522);
or U15896 (N_15896,N_15567,N_15535);
or U15897 (N_15897,N_15596,N_15721);
nor U15898 (N_15898,N_15717,N_15682);
or U15899 (N_15899,N_15689,N_15506);
and U15900 (N_15900,N_15626,N_15672);
and U15901 (N_15901,N_15734,N_15542);
nor U15902 (N_15902,N_15504,N_15678);
or U15903 (N_15903,N_15682,N_15545);
nor U15904 (N_15904,N_15721,N_15699);
xor U15905 (N_15905,N_15707,N_15700);
xor U15906 (N_15906,N_15683,N_15623);
nor U15907 (N_15907,N_15547,N_15533);
nand U15908 (N_15908,N_15686,N_15722);
nor U15909 (N_15909,N_15715,N_15726);
or U15910 (N_15910,N_15609,N_15736);
or U15911 (N_15911,N_15597,N_15535);
nand U15912 (N_15912,N_15739,N_15509);
nor U15913 (N_15913,N_15554,N_15570);
nand U15914 (N_15914,N_15675,N_15584);
nand U15915 (N_15915,N_15510,N_15591);
nand U15916 (N_15916,N_15553,N_15583);
nor U15917 (N_15917,N_15513,N_15601);
nor U15918 (N_15918,N_15545,N_15557);
xnor U15919 (N_15919,N_15745,N_15507);
and U15920 (N_15920,N_15688,N_15719);
nor U15921 (N_15921,N_15717,N_15516);
or U15922 (N_15922,N_15538,N_15693);
xor U15923 (N_15923,N_15517,N_15528);
and U15924 (N_15924,N_15729,N_15536);
nand U15925 (N_15925,N_15565,N_15587);
xnor U15926 (N_15926,N_15593,N_15581);
nand U15927 (N_15927,N_15739,N_15659);
or U15928 (N_15928,N_15670,N_15525);
or U15929 (N_15929,N_15718,N_15647);
or U15930 (N_15930,N_15583,N_15725);
and U15931 (N_15931,N_15584,N_15525);
nor U15932 (N_15932,N_15574,N_15685);
nor U15933 (N_15933,N_15681,N_15509);
nor U15934 (N_15934,N_15544,N_15542);
and U15935 (N_15935,N_15565,N_15675);
or U15936 (N_15936,N_15713,N_15533);
xnor U15937 (N_15937,N_15661,N_15745);
or U15938 (N_15938,N_15679,N_15506);
nor U15939 (N_15939,N_15714,N_15697);
nor U15940 (N_15940,N_15692,N_15630);
nand U15941 (N_15941,N_15669,N_15658);
or U15942 (N_15942,N_15583,N_15653);
or U15943 (N_15943,N_15531,N_15551);
nand U15944 (N_15944,N_15577,N_15720);
or U15945 (N_15945,N_15626,N_15508);
and U15946 (N_15946,N_15678,N_15654);
xnor U15947 (N_15947,N_15671,N_15669);
nand U15948 (N_15948,N_15602,N_15582);
and U15949 (N_15949,N_15559,N_15651);
or U15950 (N_15950,N_15621,N_15605);
and U15951 (N_15951,N_15535,N_15547);
xnor U15952 (N_15952,N_15639,N_15703);
and U15953 (N_15953,N_15514,N_15560);
nand U15954 (N_15954,N_15576,N_15688);
or U15955 (N_15955,N_15590,N_15583);
nor U15956 (N_15956,N_15525,N_15617);
nor U15957 (N_15957,N_15739,N_15632);
and U15958 (N_15958,N_15600,N_15655);
or U15959 (N_15959,N_15632,N_15622);
nor U15960 (N_15960,N_15526,N_15572);
or U15961 (N_15961,N_15586,N_15547);
xnor U15962 (N_15962,N_15629,N_15712);
nand U15963 (N_15963,N_15663,N_15673);
xnor U15964 (N_15964,N_15719,N_15708);
and U15965 (N_15965,N_15709,N_15521);
nand U15966 (N_15966,N_15608,N_15629);
or U15967 (N_15967,N_15631,N_15726);
or U15968 (N_15968,N_15574,N_15634);
nor U15969 (N_15969,N_15717,N_15508);
nor U15970 (N_15970,N_15526,N_15540);
nand U15971 (N_15971,N_15620,N_15663);
or U15972 (N_15972,N_15624,N_15742);
xnor U15973 (N_15973,N_15667,N_15573);
xor U15974 (N_15974,N_15700,N_15735);
nand U15975 (N_15975,N_15736,N_15673);
xor U15976 (N_15976,N_15642,N_15543);
nor U15977 (N_15977,N_15657,N_15569);
nand U15978 (N_15978,N_15501,N_15600);
nand U15979 (N_15979,N_15508,N_15722);
xnor U15980 (N_15980,N_15637,N_15729);
xor U15981 (N_15981,N_15647,N_15695);
nand U15982 (N_15982,N_15508,N_15563);
nor U15983 (N_15983,N_15575,N_15629);
or U15984 (N_15984,N_15586,N_15534);
nand U15985 (N_15985,N_15598,N_15542);
xor U15986 (N_15986,N_15674,N_15519);
nand U15987 (N_15987,N_15589,N_15601);
xnor U15988 (N_15988,N_15673,N_15538);
or U15989 (N_15989,N_15546,N_15746);
nor U15990 (N_15990,N_15728,N_15704);
and U15991 (N_15991,N_15552,N_15506);
nand U15992 (N_15992,N_15580,N_15744);
nand U15993 (N_15993,N_15645,N_15665);
nand U15994 (N_15994,N_15718,N_15535);
and U15995 (N_15995,N_15580,N_15505);
nand U15996 (N_15996,N_15519,N_15661);
nand U15997 (N_15997,N_15650,N_15564);
nor U15998 (N_15998,N_15665,N_15616);
xor U15999 (N_15999,N_15628,N_15555);
nor U16000 (N_16000,N_15991,N_15975);
and U16001 (N_16001,N_15802,N_15864);
xnor U16002 (N_16002,N_15755,N_15893);
and U16003 (N_16003,N_15815,N_15916);
xnor U16004 (N_16004,N_15971,N_15912);
and U16005 (N_16005,N_15931,N_15878);
nand U16006 (N_16006,N_15988,N_15918);
and U16007 (N_16007,N_15941,N_15839);
or U16008 (N_16008,N_15830,N_15958);
nor U16009 (N_16009,N_15964,N_15906);
xnor U16010 (N_16010,N_15981,N_15952);
nand U16011 (N_16011,N_15885,N_15966);
nand U16012 (N_16012,N_15969,N_15915);
or U16013 (N_16013,N_15832,N_15803);
nand U16014 (N_16014,N_15820,N_15961);
nor U16015 (N_16015,N_15833,N_15945);
nor U16016 (N_16016,N_15985,N_15978);
nor U16017 (N_16017,N_15826,N_15873);
or U16018 (N_16018,N_15756,N_15807);
and U16019 (N_16019,N_15902,N_15851);
and U16020 (N_16020,N_15750,N_15960);
nor U16021 (N_16021,N_15948,N_15977);
xnor U16022 (N_16022,N_15800,N_15859);
xnor U16023 (N_16023,N_15947,N_15974);
nand U16024 (N_16024,N_15894,N_15779);
or U16025 (N_16025,N_15796,N_15842);
nand U16026 (N_16026,N_15854,N_15816);
xor U16027 (N_16027,N_15970,N_15999);
xor U16028 (N_16028,N_15836,N_15761);
and U16029 (N_16029,N_15776,N_15812);
or U16030 (N_16030,N_15786,N_15870);
or U16031 (N_16031,N_15751,N_15879);
xor U16032 (N_16032,N_15811,N_15758);
nor U16033 (N_16033,N_15943,N_15998);
xor U16034 (N_16034,N_15899,N_15809);
nor U16035 (N_16035,N_15797,N_15858);
or U16036 (N_16036,N_15959,N_15817);
nor U16037 (N_16037,N_15869,N_15877);
or U16038 (N_16038,N_15848,N_15949);
xnor U16039 (N_16039,N_15872,N_15788);
nand U16040 (N_16040,N_15835,N_15890);
and U16041 (N_16041,N_15976,N_15767);
nand U16042 (N_16042,N_15806,N_15987);
xor U16043 (N_16043,N_15884,N_15838);
or U16044 (N_16044,N_15891,N_15940);
nand U16045 (N_16045,N_15955,N_15901);
nand U16046 (N_16046,N_15799,N_15954);
nor U16047 (N_16047,N_15930,N_15825);
and U16048 (N_16048,N_15759,N_15900);
and U16049 (N_16049,N_15917,N_15777);
nor U16050 (N_16050,N_15798,N_15925);
nor U16051 (N_16051,N_15904,N_15804);
nand U16052 (N_16052,N_15994,N_15942);
and U16053 (N_16053,N_15946,N_15793);
nor U16054 (N_16054,N_15775,N_15760);
and U16055 (N_16055,N_15914,N_15923);
nand U16056 (N_16056,N_15828,N_15920);
nand U16057 (N_16057,N_15827,N_15989);
xnor U16058 (N_16058,N_15924,N_15783);
xor U16059 (N_16059,N_15853,N_15903);
and U16060 (N_16060,N_15754,N_15782);
and U16061 (N_16061,N_15837,N_15944);
and U16062 (N_16062,N_15763,N_15973);
nor U16063 (N_16063,N_15979,N_15992);
and U16064 (N_16064,N_15822,N_15933);
nor U16065 (N_16065,N_15892,N_15932);
or U16066 (N_16066,N_15962,N_15897);
and U16067 (N_16067,N_15857,N_15913);
xor U16068 (N_16068,N_15935,N_15927);
nor U16069 (N_16069,N_15909,N_15982);
nand U16070 (N_16070,N_15773,N_15895);
and U16071 (N_16071,N_15928,N_15965);
and U16072 (N_16072,N_15846,N_15997);
xnor U16073 (N_16073,N_15937,N_15995);
or U16074 (N_16074,N_15792,N_15871);
xor U16075 (N_16075,N_15875,N_15865);
nand U16076 (N_16076,N_15910,N_15847);
xor U16077 (N_16077,N_15936,N_15785);
nand U16078 (N_16078,N_15770,N_15813);
nor U16079 (N_16079,N_15956,N_15860);
nor U16080 (N_16080,N_15907,N_15787);
nor U16081 (N_16081,N_15953,N_15823);
or U16082 (N_16082,N_15951,N_15990);
or U16083 (N_16083,N_15866,N_15929);
or U16084 (N_16084,N_15766,N_15934);
or U16085 (N_16085,N_15957,N_15810);
and U16086 (N_16086,N_15868,N_15939);
or U16087 (N_16087,N_15840,N_15852);
nor U16088 (N_16088,N_15963,N_15753);
nor U16089 (N_16089,N_15769,N_15752);
xnor U16090 (N_16090,N_15862,N_15896);
nand U16091 (N_16091,N_15790,N_15972);
or U16092 (N_16092,N_15781,N_15780);
xnor U16093 (N_16093,N_15824,N_15757);
xor U16094 (N_16094,N_15950,N_15849);
and U16095 (N_16095,N_15831,N_15794);
or U16096 (N_16096,N_15967,N_15888);
and U16097 (N_16097,N_15996,N_15808);
nor U16098 (N_16098,N_15784,N_15980);
and U16099 (N_16099,N_15887,N_15834);
or U16100 (N_16100,N_15983,N_15883);
nand U16101 (N_16101,N_15843,N_15774);
and U16102 (N_16102,N_15886,N_15771);
xnor U16103 (N_16103,N_15850,N_15986);
or U16104 (N_16104,N_15829,N_15921);
xor U16105 (N_16105,N_15889,N_15856);
and U16106 (N_16106,N_15968,N_15876);
nor U16107 (N_16107,N_15905,N_15772);
nand U16108 (N_16108,N_15993,N_15938);
nor U16109 (N_16109,N_15898,N_15765);
and U16110 (N_16110,N_15768,N_15814);
and U16111 (N_16111,N_15795,N_15762);
nand U16112 (N_16112,N_15874,N_15801);
xnor U16113 (N_16113,N_15789,N_15841);
xor U16114 (N_16114,N_15844,N_15882);
xnor U16115 (N_16115,N_15805,N_15845);
and U16116 (N_16116,N_15984,N_15791);
and U16117 (N_16117,N_15881,N_15821);
xnor U16118 (N_16118,N_15867,N_15911);
and U16119 (N_16119,N_15818,N_15764);
xor U16120 (N_16120,N_15880,N_15778);
or U16121 (N_16121,N_15926,N_15919);
xnor U16122 (N_16122,N_15861,N_15819);
and U16123 (N_16123,N_15922,N_15863);
and U16124 (N_16124,N_15855,N_15908);
and U16125 (N_16125,N_15949,N_15998);
or U16126 (N_16126,N_15840,N_15900);
xnor U16127 (N_16127,N_15980,N_15827);
nor U16128 (N_16128,N_15963,N_15785);
nor U16129 (N_16129,N_15794,N_15835);
or U16130 (N_16130,N_15876,N_15949);
and U16131 (N_16131,N_15801,N_15804);
nor U16132 (N_16132,N_15892,N_15804);
or U16133 (N_16133,N_15974,N_15753);
nor U16134 (N_16134,N_15891,N_15816);
nor U16135 (N_16135,N_15770,N_15821);
nand U16136 (N_16136,N_15982,N_15754);
xnor U16137 (N_16137,N_15759,N_15754);
and U16138 (N_16138,N_15867,N_15879);
and U16139 (N_16139,N_15781,N_15775);
and U16140 (N_16140,N_15956,N_15832);
nand U16141 (N_16141,N_15788,N_15793);
and U16142 (N_16142,N_15804,N_15888);
or U16143 (N_16143,N_15806,N_15996);
and U16144 (N_16144,N_15845,N_15797);
xor U16145 (N_16145,N_15779,N_15893);
nand U16146 (N_16146,N_15835,N_15944);
nor U16147 (N_16147,N_15768,N_15965);
nor U16148 (N_16148,N_15909,N_15854);
xnor U16149 (N_16149,N_15994,N_15988);
or U16150 (N_16150,N_15806,N_15972);
nor U16151 (N_16151,N_15888,N_15893);
or U16152 (N_16152,N_15784,N_15843);
xor U16153 (N_16153,N_15961,N_15872);
or U16154 (N_16154,N_15943,N_15781);
and U16155 (N_16155,N_15874,N_15862);
nand U16156 (N_16156,N_15909,N_15890);
nor U16157 (N_16157,N_15783,N_15816);
nor U16158 (N_16158,N_15881,N_15966);
xnor U16159 (N_16159,N_15959,N_15985);
or U16160 (N_16160,N_15912,N_15817);
nor U16161 (N_16161,N_15788,N_15996);
xor U16162 (N_16162,N_15869,N_15855);
and U16163 (N_16163,N_15910,N_15803);
xor U16164 (N_16164,N_15800,N_15816);
or U16165 (N_16165,N_15775,N_15924);
nand U16166 (N_16166,N_15843,N_15942);
or U16167 (N_16167,N_15987,N_15884);
nor U16168 (N_16168,N_15971,N_15824);
and U16169 (N_16169,N_15781,N_15886);
xnor U16170 (N_16170,N_15815,N_15773);
nor U16171 (N_16171,N_15841,N_15781);
nor U16172 (N_16172,N_15876,N_15822);
and U16173 (N_16173,N_15831,N_15869);
nand U16174 (N_16174,N_15911,N_15893);
nor U16175 (N_16175,N_15868,N_15947);
xnor U16176 (N_16176,N_15763,N_15864);
nand U16177 (N_16177,N_15978,N_15879);
and U16178 (N_16178,N_15924,N_15981);
xnor U16179 (N_16179,N_15874,N_15997);
nand U16180 (N_16180,N_15979,N_15950);
xor U16181 (N_16181,N_15897,N_15823);
and U16182 (N_16182,N_15891,N_15813);
xor U16183 (N_16183,N_15977,N_15982);
or U16184 (N_16184,N_15996,N_15945);
nor U16185 (N_16185,N_15757,N_15930);
and U16186 (N_16186,N_15782,N_15939);
nor U16187 (N_16187,N_15998,N_15906);
nand U16188 (N_16188,N_15773,N_15838);
nand U16189 (N_16189,N_15756,N_15812);
and U16190 (N_16190,N_15955,N_15840);
nand U16191 (N_16191,N_15800,N_15925);
nand U16192 (N_16192,N_15946,N_15993);
or U16193 (N_16193,N_15854,N_15765);
nand U16194 (N_16194,N_15956,N_15932);
or U16195 (N_16195,N_15922,N_15887);
xnor U16196 (N_16196,N_15990,N_15818);
nor U16197 (N_16197,N_15823,N_15847);
nor U16198 (N_16198,N_15993,N_15835);
or U16199 (N_16199,N_15775,N_15962);
or U16200 (N_16200,N_15792,N_15827);
nor U16201 (N_16201,N_15994,N_15936);
xnor U16202 (N_16202,N_15968,N_15918);
nor U16203 (N_16203,N_15831,N_15899);
nand U16204 (N_16204,N_15840,N_15918);
and U16205 (N_16205,N_15880,N_15890);
nor U16206 (N_16206,N_15835,N_15969);
or U16207 (N_16207,N_15886,N_15824);
nor U16208 (N_16208,N_15869,N_15974);
nor U16209 (N_16209,N_15958,N_15813);
and U16210 (N_16210,N_15933,N_15835);
and U16211 (N_16211,N_15981,N_15912);
and U16212 (N_16212,N_15974,N_15756);
xor U16213 (N_16213,N_15824,N_15953);
xor U16214 (N_16214,N_15910,N_15878);
or U16215 (N_16215,N_15975,N_15922);
and U16216 (N_16216,N_15775,N_15784);
or U16217 (N_16217,N_15788,N_15994);
nand U16218 (N_16218,N_15994,N_15828);
nor U16219 (N_16219,N_15806,N_15917);
nor U16220 (N_16220,N_15802,N_15792);
nand U16221 (N_16221,N_15794,N_15945);
or U16222 (N_16222,N_15758,N_15937);
and U16223 (N_16223,N_15897,N_15923);
nor U16224 (N_16224,N_15855,N_15968);
nand U16225 (N_16225,N_15807,N_15791);
nor U16226 (N_16226,N_15902,N_15993);
and U16227 (N_16227,N_15984,N_15933);
and U16228 (N_16228,N_15879,N_15939);
xnor U16229 (N_16229,N_15881,N_15847);
nor U16230 (N_16230,N_15822,N_15848);
nand U16231 (N_16231,N_15983,N_15792);
nand U16232 (N_16232,N_15870,N_15766);
nand U16233 (N_16233,N_15912,N_15851);
nand U16234 (N_16234,N_15912,N_15975);
or U16235 (N_16235,N_15872,N_15761);
and U16236 (N_16236,N_15864,N_15769);
nor U16237 (N_16237,N_15886,N_15927);
xor U16238 (N_16238,N_15857,N_15825);
xnor U16239 (N_16239,N_15941,N_15798);
xnor U16240 (N_16240,N_15857,N_15975);
xnor U16241 (N_16241,N_15908,N_15782);
xor U16242 (N_16242,N_15817,N_15973);
and U16243 (N_16243,N_15925,N_15965);
xnor U16244 (N_16244,N_15880,N_15767);
xnor U16245 (N_16245,N_15877,N_15942);
nor U16246 (N_16246,N_15794,N_15802);
nor U16247 (N_16247,N_15753,N_15773);
xor U16248 (N_16248,N_15842,N_15984);
nand U16249 (N_16249,N_15767,N_15910);
xor U16250 (N_16250,N_16191,N_16185);
nor U16251 (N_16251,N_16150,N_16121);
and U16252 (N_16252,N_16188,N_16128);
and U16253 (N_16253,N_16067,N_16011);
nand U16254 (N_16254,N_16097,N_16117);
or U16255 (N_16255,N_16171,N_16072);
or U16256 (N_16256,N_16239,N_16020);
xnor U16257 (N_16257,N_16133,N_16243);
nand U16258 (N_16258,N_16081,N_16061);
nor U16259 (N_16259,N_16194,N_16071);
xnor U16260 (N_16260,N_16079,N_16029);
or U16261 (N_16261,N_16063,N_16028);
and U16262 (N_16262,N_16051,N_16153);
xnor U16263 (N_16263,N_16147,N_16219);
xor U16264 (N_16264,N_16215,N_16232);
and U16265 (N_16265,N_16100,N_16162);
xnor U16266 (N_16266,N_16076,N_16134);
nor U16267 (N_16267,N_16013,N_16123);
and U16268 (N_16268,N_16113,N_16106);
nand U16269 (N_16269,N_16172,N_16039);
or U16270 (N_16270,N_16052,N_16196);
nor U16271 (N_16271,N_16060,N_16065);
xnor U16272 (N_16272,N_16008,N_16221);
nand U16273 (N_16273,N_16021,N_16170);
or U16274 (N_16274,N_16179,N_16057);
or U16275 (N_16275,N_16132,N_16111);
or U16276 (N_16276,N_16160,N_16098);
nand U16277 (N_16277,N_16141,N_16088);
and U16278 (N_16278,N_16032,N_16237);
nand U16279 (N_16279,N_16140,N_16165);
and U16280 (N_16280,N_16093,N_16108);
nor U16281 (N_16281,N_16030,N_16122);
nand U16282 (N_16282,N_16077,N_16037);
nor U16283 (N_16283,N_16047,N_16182);
and U16284 (N_16284,N_16145,N_16214);
and U16285 (N_16285,N_16101,N_16201);
or U16286 (N_16286,N_16027,N_16216);
nor U16287 (N_16287,N_16022,N_16238);
nor U16288 (N_16288,N_16007,N_16049);
xnor U16289 (N_16289,N_16026,N_16164);
xor U16290 (N_16290,N_16136,N_16205);
xor U16291 (N_16291,N_16228,N_16190);
and U16292 (N_16292,N_16207,N_16159);
nor U16293 (N_16293,N_16224,N_16073);
xor U16294 (N_16294,N_16249,N_16019);
or U16295 (N_16295,N_16112,N_16040);
and U16296 (N_16296,N_16070,N_16235);
xor U16297 (N_16297,N_16158,N_16035);
nor U16298 (N_16298,N_16083,N_16090);
or U16299 (N_16299,N_16233,N_16127);
xor U16300 (N_16300,N_16055,N_16208);
or U16301 (N_16301,N_16003,N_16087);
and U16302 (N_16302,N_16107,N_16034);
nor U16303 (N_16303,N_16126,N_16152);
nand U16304 (N_16304,N_16240,N_16193);
or U16305 (N_16305,N_16074,N_16069);
and U16306 (N_16306,N_16234,N_16005);
nand U16307 (N_16307,N_16018,N_16082);
and U16308 (N_16308,N_16043,N_16181);
xnor U16309 (N_16309,N_16119,N_16059);
xor U16310 (N_16310,N_16095,N_16161);
nor U16311 (N_16311,N_16062,N_16149);
nand U16312 (N_16312,N_16246,N_16050);
and U16313 (N_16313,N_16189,N_16148);
or U16314 (N_16314,N_16200,N_16016);
nand U16315 (N_16315,N_16120,N_16092);
and U16316 (N_16316,N_16010,N_16192);
and U16317 (N_16317,N_16105,N_16236);
nand U16318 (N_16318,N_16231,N_16096);
and U16319 (N_16319,N_16110,N_16064);
nand U16320 (N_16320,N_16089,N_16042);
xnor U16321 (N_16321,N_16183,N_16058);
xor U16322 (N_16322,N_16198,N_16176);
or U16323 (N_16323,N_16163,N_16229);
or U16324 (N_16324,N_16226,N_16211);
xor U16325 (N_16325,N_16230,N_16002);
nand U16326 (N_16326,N_16033,N_16178);
and U16327 (N_16327,N_16168,N_16038);
nand U16328 (N_16328,N_16156,N_16115);
and U16329 (N_16329,N_16130,N_16056);
and U16330 (N_16330,N_16180,N_16085);
nor U16331 (N_16331,N_16116,N_16080);
or U16332 (N_16332,N_16175,N_16151);
nand U16333 (N_16333,N_16166,N_16142);
and U16334 (N_16334,N_16187,N_16114);
nand U16335 (N_16335,N_16220,N_16131);
and U16336 (N_16336,N_16006,N_16066);
nor U16337 (N_16337,N_16138,N_16212);
xnor U16338 (N_16338,N_16045,N_16099);
nand U16339 (N_16339,N_16199,N_16118);
xnor U16340 (N_16340,N_16217,N_16245);
nand U16341 (N_16341,N_16014,N_16157);
or U16342 (N_16342,N_16031,N_16000);
nand U16343 (N_16343,N_16210,N_16012);
nor U16344 (N_16344,N_16203,N_16102);
and U16345 (N_16345,N_16017,N_16244);
and U16346 (N_16346,N_16004,N_16197);
and U16347 (N_16347,N_16048,N_16124);
xnor U16348 (N_16348,N_16227,N_16209);
nor U16349 (N_16349,N_16146,N_16177);
nand U16350 (N_16350,N_16125,N_16024);
or U16351 (N_16351,N_16143,N_16023);
xor U16352 (N_16352,N_16091,N_16195);
or U16353 (N_16353,N_16044,N_16103);
nor U16354 (N_16354,N_16094,N_16104);
and U16355 (N_16355,N_16222,N_16174);
and U16356 (N_16356,N_16242,N_16241);
and U16357 (N_16357,N_16129,N_16154);
nand U16358 (N_16358,N_16086,N_16025);
or U16359 (N_16359,N_16144,N_16137);
or U16360 (N_16360,N_16054,N_16202);
or U16361 (N_16361,N_16169,N_16223);
or U16362 (N_16362,N_16155,N_16213);
xnor U16363 (N_16363,N_16015,N_16218);
or U16364 (N_16364,N_16186,N_16075);
nor U16365 (N_16365,N_16247,N_16009);
and U16366 (N_16366,N_16109,N_16248);
or U16367 (N_16367,N_16184,N_16173);
xnor U16368 (N_16368,N_16046,N_16206);
and U16369 (N_16369,N_16041,N_16204);
xor U16370 (N_16370,N_16139,N_16036);
xnor U16371 (N_16371,N_16078,N_16135);
and U16372 (N_16372,N_16068,N_16167);
and U16373 (N_16373,N_16053,N_16225);
or U16374 (N_16374,N_16001,N_16084);
nor U16375 (N_16375,N_16185,N_16206);
and U16376 (N_16376,N_16239,N_16146);
and U16377 (N_16377,N_16175,N_16229);
nor U16378 (N_16378,N_16142,N_16176);
nor U16379 (N_16379,N_16242,N_16162);
nand U16380 (N_16380,N_16046,N_16218);
xnor U16381 (N_16381,N_16003,N_16114);
nor U16382 (N_16382,N_16044,N_16075);
and U16383 (N_16383,N_16076,N_16004);
or U16384 (N_16384,N_16198,N_16249);
nand U16385 (N_16385,N_16241,N_16218);
xnor U16386 (N_16386,N_16157,N_16174);
nor U16387 (N_16387,N_16073,N_16190);
and U16388 (N_16388,N_16039,N_16021);
nor U16389 (N_16389,N_16022,N_16236);
nor U16390 (N_16390,N_16108,N_16001);
and U16391 (N_16391,N_16141,N_16089);
or U16392 (N_16392,N_16105,N_16106);
or U16393 (N_16393,N_16050,N_16159);
nand U16394 (N_16394,N_16036,N_16042);
xnor U16395 (N_16395,N_16039,N_16185);
xnor U16396 (N_16396,N_16244,N_16222);
and U16397 (N_16397,N_16213,N_16144);
and U16398 (N_16398,N_16027,N_16219);
nand U16399 (N_16399,N_16172,N_16011);
nor U16400 (N_16400,N_16195,N_16124);
xor U16401 (N_16401,N_16175,N_16237);
nand U16402 (N_16402,N_16124,N_16143);
or U16403 (N_16403,N_16125,N_16011);
or U16404 (N_16404,N_16170,N_16107);
or U16405 (N_16405,N_16134,N_16077);
or U16406 (N_16406,N_16012,N_16112);
xor U16407 (N_16407,N_16104,N_16138);
xor U16408 (N_16408,N_16218,N_16003);
xor U16409 (N_16409,N_16227,N_16113);
nand U16410 (N_16410,N_16168,N_16083);
or U16411 (N_16411,N_16063,N_16102);
nand U16412 (N_16412,N_16147,N_16009);
and U16413 (N_16413,N_16019,N_16072);
xnor U16414 (N_16414,N_16171,N_16107);
or U16415 (N_16415,N_16143,N_16043);
and U16416 (N_16416,N_16076,N_16195);
xor U16417 (N_16417,N_16216,N_16190);
nand U16418 (N_16418,N_16139,N_16209);
and U16419 (N_16419,N_16165,N_16035);
or U16420 (N_16420,N_16235,N_16009);
or U16421 (N_16421,N_16053,N_16150);
nor U16422 (N_16422,N_16100,N_16171);
xor U16423 (N_16423,N_16039,N_16136);
nand U16424 (N_16424,N_16103,N_16106);
xnor U16425 (N_16425,N_16037,N_16213);
xor U16426 (N_16426,N_16212,N_16025);
nand U16427 (N_16427,N_16013,N_16146);
or U16428 (N_16428,N_16112,N_16144);
or U16429 (N_16429,N_16218,N_16226);
or U16430 (N_16430,N_16194,N_16243);
xor U16431 (N_16431,N_16027,N_16196);
nand U16432 (N_16432,N_16160,N_16244);
xor U16433 (N_16433,N_16054,N_16163);
nand U16434 (N_16434,N_16247,N_16189);
and U16435 (N_16435,N_16145,N_16042);
nand U16436 (N_16436,N_16020,N_16193);
nor U16437 (N_16437,N_16135,N_16051);
xor U16438 (N_16438,N_16249,N_16180);
xor U16439 (N_16439,N_16134,N_16200);
or U16440 (N_16440,N_16118,N_16232);
nor U16441 (N_16441,N_16109,N_16099);
nor U16442 (N_16442,N_16050,N_16121);
and U16443 (N_16443,N_16087,N_16028);
or U16444 (N_16444,N_16249,N_16101);
nand U16445 (N_16445,N_16083,N_16237);
nor U16446 (N_16446,N_16040,N_16181);
nor U16447 (N_16447,N_16179,N_16031);
nand U16448 (N_16448,N_16086,N_16083);
nor U16449 (N_16449,N_16193,N_16128);
and U16450 (N_16450,N_16149,N_16169);
xor U16451 (N_16451,N_16177,N_16032);
nor U16452 (N_16452,N_16035,N_16001);
and U16453 (N_16453,N_16225,N_16214);
and U16454 (N_16454,N_16142,N_16237);
nand U16455 (N_16455,N_16076,N_16084);
nor U16456 (N_16456,N_16101,N_16086);
xnor U16457 (N_16457,N_16178,N_16132);
and U16458 (N_16458,N_16111,N_16131);
and U16459 (N_16459,N_16182,N_16248);
and U16460 (N_16460,N_16063,N_16180);
nor U16461 (N_16461,N_16207,N_16066);
or U16462 (N_16462,N_16232,N_16177);
and U16463 (N_16463,N_16066,N_16164);
nor U16464 (N_16464,N_16110,N_16223);
nand U16465 (N_16465,N_16246,N_16227);
and U16466 (N_16466,N_16235,N_16154);
or U16467 (N_16467,N_16207,N_16187);
nor U16468 (N_16468,N_16092,N_16053);
nand U16469 (N_16469,N_16075,N_16018);
nor U16470 (N_16470,N_16096,N_16113);
or U16471 (N_16471,N_16150,N_16020);
nor U16472 (N_16472,N_16070,N_16178);
or U16473 (N_16473,N_16088,N_16169);
nor U16474 (N_16474,N_16042,N_16184);
and U16475 (N_16475,N_16026,N_16043);
and U16476 (N_16476,N_16220,N_16238);
and U16477 (N_16477,N_16230,N_16211);
xnor U16478 (N_16478,N_16109,N_16065);
and U16479 (N_16479,N_16179,N_16034);
or U16480 (N_16480,N_16134,N_16122);
xnor U16481 (N_16481,N_16104,N_16144);
and U16482 (N_16482,N_16099,N_16190);
nand U16483 (N_16483,N_16225,N_16076);
xor U16484 (N_16484,N_16242,N_16118);
nand U16485 (N_16485,N_16033,N_16224);
or U16486 (N_16486,N_16162,N_16145);
nor U16487 (N_16487,N_16146,N_16226);
nand U16488 (N_16488,N_16173,N_16103);
or U16489 (N_16489,N_16053,N_16031);
nand U16490 (N_16490,N_16190,N_16090);
nor U16491 (N_16491,N_16073,N_16229);
and U16492 (N_16492,N_16151,N_16249);
nor U16493 (N_16493,N_16141,N_16232);
or U16494 (N_16494,N_16247,N_16083);
nor U16495 (N_16495,N_16124,N_16008);
and U16496 (N_16496,N_16176,N_16155);
nand U16497 (N_16497,N_16067,N_16152);
and U16498 (N_16498,N_16015,N_16186);
or U16499 (N_16499,N_16174,N_16168);
or U16500 (N_16500,N_16315,N_16468);
nor U16501 (N_16501,N_16409,N_16440);
or U16502 (N_16502,N_16410,N_16292);
or U16503 (N_16503,N_16296,N_16284);
xnor U16504 (N_16504,N_16367,N_16434);
nand U16505 (N_16505,N_16407,N_16310);
nand U16506 (N_16506,N_16355,N_16364);
and U16507 (N_16507,N_16471,N_16452);
or U16508 (N_16508,N_16251,N_16405);
nand U16509 (N_16509,N_16335,N_16469);
or U16510 (N_16510,N_16262,N_16441);
nor U16511 (N_16511,N_16485,N_16481);
or U16512 (N_16512,N_16374,N_16337);
or U16513 (N_16513,N_16400,N_16422);
nor U16514 (N_16514,N_16454,N_16484);
and U16515 (N_16515,N_16304,N_16278);
nand U16516 (N_16516,N_16342,N_16359);
xor U16517 (N_16517,N_16276,N_16493);
or U16518 (N_16518,N_16309,N_16346);
xnor U16519 (N_16519,N_16438,N_16444);
xnor U16520 (N_16520,N_16338,N_16302);
nand U16521 (N_16521,N_16386,N_16483);
nor U16522 (N_16522,N_16428,N_16265);
nor U16523 (N_16523,N_16253,N_16482);
or U16524 (N_16524,N_16496,N_16476);
and U16525 (N_16525,N_16254,N_16344);
or U16526 (N_16526,N_16394,N_16312);
xnor U16527 (N_16527,N_16329,N_16474);
xnor U16528 (N_16528,N_16472,N_16412);
or U16529 (N_16529,N_16281,N_16420);
nand U16530 (N_16530,N_16497,N_16317);
nand U16531 (N_16531,N_16263,N_16490);
nand U16532 (N_16532,N_16361,N_16431);
xor U16533 (N_16533,N_16369,N_16383);
nand U16534 (N_16534,N_16390,N_16321);
or U16535 (N_16535,N_16343,N_16380);
xor U16536 (N_16536,N_16399,N_16358);
and U16537 (N_16537,N_16272,N_16373);
xor U16538 (N_16538,N_16453,N_16418);
xnor U16539 (N_16539,N_16379,N_16449);
xnor U16540 (N_16540,N_16271,N_16462);
or U16541 (N_16541,N_16421,N_16297);
nor U16542 (N_16542,N_16378,N_16457);
nand U16543 (N_16543,N_16425,N_16460);
nand U16544 (N_16544,N_16261,N_16356);
nor U16545 (N_16545,N_16331,N_16455);
or U16546 (N_16546,N_16280,N_16328);
nor U16547 (N_16547,N_16345,N_16387);
nor U16548 (N_16548,N_16488,N_16294);
xor U16549 (N_16549,N_16450,N_16318);
or U16550 (N_16550,N_16397,N_16432);
or U16551 (N_16551,N_16314,N_16406);
nor U16552 (N_16552,N_16436,N_16258);
nand U16553 (N_16553,N_16267,N_16316);
or U16554 (N_16554,N_16423,N_16250);
and U16555 (N_16555,N_16494,N_16486);
xnor U16556 (N_16556,N_16376,N_16442);
nor U16557 (N_16557,N_16363,N_16259);
nand U16558 (N_16558,N_16325,N_16349);
and U16559 (N_16559,N_16347,N_16333);
and U16560 (N_16560,N_16445,N_16458);
or U16561 (N_16561,N_16403,N_16323);
and U16562 (N_16562,N_16392,N_16341);
nand U16563 (N_16563,N_16368,N_16467);
and U16564 (N_16564,N_16446,N_16498);
and U16565 (N_16565,N_16275,N_16293);
or U16566 (N_16566,N_16447,N_16408);
xor U16567 (N_16567,N_16257,N_16288);
and U16568 (N_16568,N_16388,N_16464);
nand U16569 (N_16569,N_16385,N_16389);
nand U16570 (N_16570,N_16306,N_16274);
nand U16571 (N_16571,N_16300,N_16456);
and U16572 (N_16572,N_16255,N_16350);
nor U16573 (N_16573,N_16417,N_16339);
xor U16574 (N_16574,N_16366,N_16324);
nor U16575 (N_16575,N_16326,N_16360);
xnor U16576 (N_16576,N_16372,N_16279);
or U16577 (N_16577,N_16424,N_16491);
or U16578 (N_16578,N_16435,N_16396);
and U16579 (N_16579,N_16414,N_16398);
and U16580 (N_16580,N_16377,N_16473);
and U16581 (N_16581,N_16270,N_16287);
and U16582 (N_16582,N_16268,N_16426);
xnor U16583 (N_16583,N_16470,N_16283);
xnor U16584 (N_16584,N_16285,N_16336);
nor U16585 (N_16585,N_16395,N_16260);
and U16586 (N_16586,N_16439,N_16451);
or U16587 (N_16587,N_16384,N_16286);
and U16588 (N_16588,N_16340,N_16308);
and U16589 (N_16589,N_16415,N_16480);
nor U16590 (N_16590,N_16461,N_16282);
nand U16591 (N_16591,N_16419,N_16348);
or U16592 (N_16592,N_16290,N_16437);
or U16593 (N_16593,N_16269,N_16429);
nand U16594 (N_16594,N_16352,N_16273);
or U16595 (N_16595,N_16319,N_16327);
and U16596 (N_16596,N_16332,N_16463);
and U16597 (N_16597,N_16401,N_16411);
nand U16598 (N_16598,N_16365,N_16334);
xnor U16599 (N_16599,N_16459,N_16495);
nor U16600 (N_16600,N_16489,N_16322);
nor U16601 (N_16601,N_16499,N_16492);
or U16602 (N_16602,N_16382,N_16404);
nand U16603 (N_16603,N_16351,N_16354);
nand U16604 (N_16604,N_16295,N_16313);
nand U16605 (N_16605,N_16413,N_16277);
xor U16606 (N_16606,N_16370,N_16256);
or U16607 (N_16607,N_16307,N_16402);
nand U16608 (N_16608,N_16375,N_16381);
and U16609 (N_16609,N_16266,N_16448);
and U16610 (N_16610,N_16465,N_16330);
or U16611 (N_16611,N_16393,N_16291);
xor U16612 (N_16612,N_16475,N_16477);
and U16613 (N_16613,N_16391,N_16264);
nor U16614 (N_16614,N_16353,N_16478);
nand U16615 (N_16615,N_16289,N_16305);
nand U16616 (N_16616,N_16311,N_16443);
or U16617 (N_16617,N_16487,N_16320);
nor U16618 (N_16618,N_16301,N_16362);
or U16619 (N_16619,N_16252,N_16433);
and U16620 (N_16620,N_16303,N_16371);
nor U16621 (N_16621,N_16416,N_16299);
xnor U16622 (N_16622,N_16298,N_16357);
xnor U16623 (N_16623,N_16430,N_16466);
nor U16624 (N_16624,N_16427,N_16479);
xnor U16625 (N_16625,N_16413,N_16364);
and U16626 (N_16626,N_16380,N_16488);
nor U16627 (N_16627,N_16330,N_16488);
xor U16628 (N_16628,N_16475,N_16310);
xor U16629 (N_16629,N_16371,N_16333);
or U16630 (N_16630,N_16487,N_16385);
and U16631 (N_16631,N_16498,N_16251);
nand U16632 (N_16632,N_16436,N_16316);
xor U16633 (N_16633,N_16495,N_16375);
and U16634 (N_16634,N_16481,N_16261);
xor U16635 (N_16635,N_16293,N_16329);
nand U16636 (N_16636,N_16446,N_16391);
and U16637 (N_16637,N_16283,N_16497);
nand U16638 (N_16638,N_16300,N_16478);
or U16639 (N_16639,N_16477,N_16428);
xnor U16640 (N_16640,N_16412,N_16436);
nor U16641 (N_16641,N_16282,N_16356);
xnor U16642 (N_16642,N_16452,N_16352);
xor U16643 (N_16643,N_16497,N_16321);
or U16644 (N_16644,N_16364,N_16352);
nand U16645 (N_16645,N_16298,N_16385);
xnor U16646 (N_16646,N_16389,N_16416);
or U16647 (N_16647,N_16460,N_16322);
or U16648 (N_16648,N_16424,N_16310);
nor U16649 (N_16649,N_16422,N_16314);
nor U16650 (N_16650,N_16407,N_16373);
and U16651 (N_16651,N_16468,N_16365);
nand U16652 (N_16652,N_16393,N_16472);
xor U16653 (N_16653,N_16352,N_16385);
or U16654 (N_16654,N_16336,N_16408);
xor U16655 (N_16655,N_16373,N_16470);
nand U16656 (N_16656,N_16284,N_16424);
and U16657 (N_16657,N_16419,N_16287);
nand U16658 (N_16658,N_16316,N_16343);
nor U16659 (N_16659,N_16274,N_16383);
nand U16660 (N_16660,N_16376,N_16473);
nor U16661 (N_16661,N_16380,N_16489);
xor U16662 (N_16662,N_16412,N_16408);
xor U16663 (N_16663,N_16318,N_16480);
or U16664 (N_16664,N_16342,N_16290);
xor U16665 (N_16665,N_16262,N_16422);
or U16666 (N_16666,N_16472,N_16319);
nor U16667 (N_16667,N_16359,N_16270);
and U16668 (N_16668,N_16486,N_16489);
nor U16669 (N_16669,N_16346,N_16378);
nand U16670 (N_16670,N_16255,N_16320);
and U16671 (N_16671,N_16317,N_16352);
nor U16672 (N_16672,N_16440,N_16498);
xnor U16673 (N_16673,N_16312,N_16331);
nand U16674 (N_16674,N_16485,N_16461);
xor U16675 (N_16675,N_16274,N_16356);
nand U16676 (N_16676,N_16479,N_16483);
nor U16677 (N_16677,N_16398,N_16251);
nor U16678 (N_16678,N_16290,N_16333);
nand U16679 (N_16679,N_16388,N_16369);
xor U16680 (N_16680,N_16257,N_16319);
nand U16681 (N_16681,N_16320,N_16311);
and U16682 (N_16682,N_16359,N_16417);
xnor U16683 (N_16683,N_16278,N_16409);
or U16684 (N_16684,N_16449,N_16256);
or U16685 (N_16685,N_16424,N_16499);
nand U16686 (N_16686,N_16368,N_16281);
and U16687 (N_16687,N_16498,N_16403);
or U16688 (N_16688,N_16382,N_16427);
or U16689 (N_16689,N_16382,N_16472);
and U16690 (N_16690,N_16407,N_16395);
and U16691 (N_16691,N_16441,N_16473);
or U16692 (N_16692,N_16256,N_16422);
or U16693 (N_16693,N_16254,N_16322);
nand U16694 (N_16694,N_16321,N_16435);
nand U16695 (N_16695,N_16280,N_16450);
or U16696 (N_16696,N_16332,N_16466);
or U16697 (N_16697,N_16496,N_16495);
xor U16698 (N_16698,N_16483,N_16287);
xnor U16699 (N_16699,N_16359,N_16426);
or U16700 (N_16700,N_16430,N_16497);
nand U16701 (N_16701,N_16474,N_16297);
xnor U16702 (N_16702,N_16468,N_16270);
or U16703 (N_16703,N_16319,N_16348);
or U16704 (N_16704,N_16405,N_16255);
nor U16705 (N_16705,N_16345,N_16341);
or U16706 (N_16706,N_16400,N_16300);
nor U16707 (N_16707,N_16492,N_16351);
nand U16708 (N_16708,N_16446,N_16468);
and U16709 (N_16709,N_16353,N_16255);
or U16710 (N_16710,N_16370,N_16415);
xor U16711 (N_16711,N_16323,N_16400);
xor U16712 (N_16712,N_16337,N_16450);
xor U16713 (N_16713,N_16338,N_16326);
and U16714 (N_16714,N_16270,N_16301);
nor U16715 (N_16715,N_16483,N_16410);
xnor U16716 (N_16716,N_16380,N_16262);
or U16717 (N_16717,N_16414,N_16298);
nand U16718 (N_16718,N_16396,N_16374);
xor U16719 (N_16719,N_16461,N_16493);
nor U16720 (N_16720,N_16430,N_16418);
xor U16721 (N_16721,N_16329,N_16361);
or U16722 (N_16722,N_16311,N_16301);
xor U16723 (N_16723,N_16408,N_16494);
and U16724 (N_16724,N_16327,N_16488);
nand U16725 (N_16725,N_16440,N_16470);
xor U16726 (N_16726,N_16456,N_16493);
and U16727 (N_16727,N_16374,N_16392);
nand U16728 (N_16728,N_16389,N_16311);
nand U16729 (N_16729,N_16378,N_16443);
nand U16730 (N_16730,N_16278,N_16385);
xnor U16731 (N_16731,N_16440,N_16355);
and U16732 (N_16732,N_16306,N_16454);
or U16733 (N_16733,N_16488,N_16458);
nor U16734 (N_16734,N_16350,N_16409);
or U16735 (N_16735,N_16299,N_16431);
xnor U16736 (N_16736,N_16400,N_16394);
nor U16737 (N_16737,N_16460,N_16357);
and U16738 (N_16738,N_16486,N_16254);
or U16739 (N_16739,N_16335,N_16419);
or U16740 (N_16740,N_16343,N_16473);
or U16741 (N_16741,N_16307,N_16497);
or U16742 (N_16742,N_16423,N_16456);
xnor U16743 (N_16743,N_16471,N_16311);
or U16744 (N_16744,N_16267,N_16332);
xnor U16745 (N_16745,N_16483,N_16311);
xor U16746 (N_16746,N_16331,N_16304);
and U16747 (N_16747,N_16457,N_16297);
xor U16748 (N_16748,N_16304,N_16426);
and U16749 (N_16749,N_16495,N_16408);
nand U16750 (N_16750,N_16704,N_16591);
and U16751 (N_16751,N_16745,N_16729);
xor U16752 (N_16752,N_16700,N_16594);
nand U16753 (N_16753,N_16610,N_16657);
xnor U16754 (N_16754,N_16658,N_16727);
or U16755 (N_16755,N_16708,N_16736);
and U16756 (N_16756,N_16562,N_16693);
or U16757 (N_16757,N_16501,N_16692);
xor U16758 (N_16758,N_16520,N_16654);
nor U16759 (N_16759,N_16725,N_16719);
and U16760 (N_16760,N_16611,N_16712);
xnor U16761 (N_16761,N_16525,N_16601);
nor U16762 (N_16762,N_16555,N_16739);
and U16763 (N_16763,N_16643,N_16710);
xor U16764 (N_16764,N_16568,N_16662);
and U16765 (N_16765,N_16549,N_16541);
xnor U16766 (N_16766,N_16687,N_16519);
nand U16767 (N_16767,N_16733,N_16527);
nor U16768 (N_16768,N_16641,N_16617);
and U16769 (N_16769,N_16576,N_16640);
xnor U16770 (N_16770,N_16656,N_16539);
nor U16771 (N_16771,N_16633,N_16597);
xnor U16772 (N_16772,N_16655,N_16543);
xnor U16773 (N_16773,N_16577,N_16573);
and U16774 (N_16774,N_16648,N_16626);
xnor U16775 (N_16775,N_16645,N_16668);
nand U16776 (N_16776,N_16506,N_16557);
nor U16777 (N_16777,N_16697,N_16717);
and U16778 (N_16778,N_16579,N_16550);
or U16779 (N_16779,N_16533,N_16531);
nand U16780 (N_16780,N_16571,N_16653);
xor U16781 (N_16781,N_16673,N_16627);
or U16782 (N_16782,N_16628,N_16614);
nor U16783 (N_16783,N_16676,N_16570);
or U16784 (N_16784,N_16669,N_16592);
or U16785 (N_16785,N_16596,N_16583);
xnor U16786 (N_16786,N_16618,N_16607);
and U16787 (N_16787,N_16679,N_16621);
nor U16788 (N_16788,N_16584,N_16646);
or U16789 (N_16789,N_16521,N_16559);
nand U16790 (N_16790,N_16660,N_16590);
and U16791 (N_16791,N_16644,N_16706);
xnor U16792 (N_16792,N_16609,N_16623);
and U16793 (N_16793,N_16619,N_16665);
nand U16794 (N_16794,N_16613,N_16580);
nand U16795 (N_16795,N_16552,N_16691);
or U16796 (N_16796,N_16682,N_16608);
or U16797 (N_16797,N_16681,N_16723);
nor U16798 (N_16798,N_16748,N_16743);
and U16799 (N_16799,N_16650,N_16666);
xor U16800 (N_16800,N_16625,N_16566);
or U16801 (N_16801,N_16730,N_16616);
and U16802 (N_16802,N_16512,N_16538);
xor U16803 (N_16803,N_16599,N_16516);
nor U16804 (N_16804,N_16546,N_16631);
xor U16805 (N_16805,N_16651,N_16713);
nand U16806 (N_16806,N_16690,N_16556);
or U16807 (N_16807,N_16524,N_16720);
or U16808 (N_16808,N_16636,N_16718);
nor U16809 (N_16809,N_16667,N_16707);
and U16810 (N_16810,N_16548,N_16661);
nor U16811 (N_16811,N_16734,N_16528);
and U16812 (N_16812,N_16639,N_16638);
nand U16813 (N_16813,N_16737,N_16672);
nand U16814 (N_16814,N_16586,N_16675);
nand U16815 (N_16815,N_16542,N_16522);
nor U16816 (N_16816,N_16620,N_16507);
xor U16817 (N_16817,N_16513,N_16598);
or U16818 (N_16818,N_16680,N_16561);
xnor U16819 (N_16819,N_16688,N_16558);
and U16820 (N_16820,N_16551,N_16699);
and U16821 (N_16821,N_16670,N_16634);
nor U16822 (N_16822,N_16502,N_16696);
nor U16823 (N_16823,N_16744,N_16683);
xnor U16824 (N_16824,N_16685,N_16663);
or U16825 (N_16825,N_16532,N_16677);
and U16826 (N_16826,N_16671,N_16635);
and U16827 (N_16827,N_16567,N_16588);
xor U16828 (N_16828,N_16684,N_16545);
nand U16829 (N_16829,N_16536,N_16575);
nor U16830 (N_16830,N_16726,N_16716);
xnor U16831 (N_16831,N_16605,N_16518);
and U16832 (N_16832,N_16508,N_16565);
xnor U16833 (N_16833,N_16505,N_16738);
nor U16834 (N_16834,N_16735,N_16595);
and U16835 (N_16835,N_16587,N_16732);
nand U16836 (N_16836,N_16721,N_16593);
nand U16837 (N_16837,N_16740,N_16560);
nor U16838 (N_16838,N_16711,N_16741);
nand U16839 (N_16839,N_16689,N_16600);
nor U16840 (N_16840,N_16747,N_16701);
xor U16841 (N_16841,N_16746,N_16534);
and U16842 (N_16842,N_16589,N_16742);
or U16843 (N_16843,N_16615,N_16709);
or U16844 (N_16844,N_16581,N_16702);
nor U16845 (N_16845,N_16529,N_16647);
xnor U16846 (N_16846,N_16574,N_16749);
or U16847 (N_16847,N_16724,N_16523);
or U16848 (N_16848,N_16514,N_16630);
nor U16849 (N_16849,N_16585,N_16637);
nor U16850 (N_16850,N_16517,N_16731);
xnor U16851 (N_16851,N_16624,N_16632);
or U16852 (N_16852,N_16715,N_16530);
and U16853 (N_16853,N_16503,N_16629);
nand U16854 (N_16854,N_16504,N_16511);
or U16855 (N_16855,N_16604,N_16674);
and U16856 (N_16856,N_16578,N_16642);
xnor U16857 (N_16857,N_16695,N_16582);
and U16858 (N_16858,N_16537,N_16526);
and U16859 (N_16859,N_16603,N_16535);
nor U16860 (N_16860,N_16703,N_16705);
nand U16861 (N_16861,N_16547,N_16678);
nand U16862 (N_16862,N_16500,N_16659);
nand U16863 (N_16863,N_16686,N_16572);
or U16864 (N_16864,N_16649,N_16554);
xnor U16865 (N_16865,N_16714,N_16564);
xnor U16866 (N_16866,N_16509,N_16553);
and U16867 (N_16867,N_16540,N_16728);
nor U16868 (N_16868,N_16612,N_16698);
and U16869 (N_16869,N_16602,N_16515);
nand U16870 (N_16870,N_16622,N_16606);
and U16871 (N_16871,N_16569,N_16563);
or U16872 (N_16872,N_16694,N_16510);
nor U16873 (N_16873,N_16722,N_16652);
xor U16874 (N_16874,N_16664,N_16544);
xnor U16875 (N_16875,N_16540,N_16617);
nand U16876 (N_16876,N_16734,N_16673);
xnor U16877 (N_16877,N_16552,N_16667);
nor U16878 (N_16878,N_16644,N_16508);
nand U16879 (N_16879,N_16728,N_16608);
or U16880 (N_16880,N_16629,N_16567);
nor U16881 (N_16881,N_16677,N_16645);
nand U16882 (N_16882,N_16510,N_16518);
or U16883 (N_16883,N_16537,N_16559);
and U16884 (N_16884,N_16653,N_16672);
xor U16885 (N_16885,N_16584,N_16515);
xor U16886 (N_16886,N_16577,N_16711);
nand U16887 (N_16887,N_16738,N_16596);
nor U16888 (N_16888,N_16630,N_16598);
nor U16889 (N_16889,N_16544,N_16713);
xnor U16890 (N_16890,N_16657,N_16744);
nor U16891 (N_16891,N_16713,N_16571);
xor U16892 (N_16892,N_16683,N_16614);
or U16893 (N_16893,N_16572,N_16735);
and U16894 (N_16894,N_16744,N_16677);
nand U16895 (N_16895,N_16694,N_16710);
and U16896 (N_16896,N_16566,N_16501);
and U16897 (N_16897,N_16576,N_16538);
nor U16898 (N_16898,N_16681,N_16535);
nor U16899 (N_16899,N_16716,N_16649);
or U16900 (N_16900,N_16631,N_16646);
xor U16901 (N_16901,N_16695,N_16504);
and U16902 (N_16902,N_16698,N_16704);
nor U16903 (N_16903,N_16621,N_16598);
nor U16904 (N_16904,N_16589,N_16565);
or U16905 (N_16905,N_16504,N_16513);
nand U16906 (N_16906,N_16535,N_16614);
and U16907 (N_16907,N_16501,N_16629);
or U16908 (N_16908,N_16732,N_16654);
xnor U16909 (N_16909,N_16647,N_16660);
and U16910 (N_16910,N_16599,N_16692);
or U16911 (N_16911,N_16536,N_16726);
or U16912 (N_16912,N_16554,N_16720);
xnor U16913 (N_16913,N_16742,N_16509);
nand U16914 (N_16914,N_16744,N_16553);
and U16915 (N_16915,N_16508,N_16749);
and U16916 (N_16916,N_16574,N_16661);
and U16917 (N_16917,N_16507,N_16749);
and U16918 (N_16918,N_16592,N_16570);
or U16919 (N_16919,N_16682,N_16706);
xnor U16920 (N_16920,N_16620,N_16665);
nor U16921 (N_16921,N_16689,N_16651);
nor U16922 (N_16922,N_16625,N_16571);
nand U16923 (N_16923,N_16603,N_16587);
and U16924 (N_16924,N_16748,N_16684);
nor U16925 (N_16925,N_16711,N_16746);
nor U16926 (N_16926,N_16679,N_16646);
nand U16927 (N_16927,N_16545,N_16725);
nor U16928 (N_16928,N_16505,N_16527);
xor U16929 (N_16929,N_16535,N_16531);
and U16930 (N_16930,N_16577,N_16588);
nor U16931 (N_16931,N_16593,N_16695);
or U16932 (N_16932,N_16706,N_16523);
or U16933 (N_16933,N_16575,N_16520);
nand U16934 (N_16934,N_16651,N_16586);
nand U16935 (N_16935,N_16731,N_16577);
or U16936 (N_16936,N_16603,N_16632);
nand U16937 (N_16937,N_16605,N_16739);
nand U16938 (N_16938,N_16592,N_16747);
nor U16939 (N_16939,N_16684,N_16589);
nand U16940 (N_16940,N_16536,N_16747);
xnor U16941 (N_16941,N_16684,N_16713);
nor U16942 (N_16942,N_16662,N_16682);
or U16943 (N_16943,N_16564,N_16723);
xor U16944 (N_16944,N_16583,N_16667);
xor U16945 (N_16945,N_16589,N_16679);
xnor U16946 (N_16946,N_16610,N_16706);
or U16947 (N_16947,N_16547,N_16576);
nand U16948 (N_16948,N_16733,N_16560);
nand U16949 (N_16949,N_16570,N_16572);
nor U16950 (N_16950,N_16712,N_16571);
nand U16951 (N_16951,N_16636,N_16551);
nand U16952 (N_16952,N_16501,N_16536);
xor U16953 (N_16953,N_16534,N_16599);
and U16954 (N_16954,N_16712,N_16621);
xor U16955 (N_16955,N_16601,N_16557);
xor U16956 (N_16956,N_16721,N_16558);
or U16957 (N_16957,N_16687,N_16609);
or U16958 (N_16958,N_16621,N_16656);
nor U16959 (N_16959,N_16572,N_16674);
xnor U16960 (N_16960,N_16544,N_16580);
nor U16961 (N_16961,N_16728,N_16624);
and U16962 (N_16962,N_16647,N_16512);
nor U16963 (N_16963,N_16625,N_16588);
xnor U16964 (N_16964,N_16734,N_16604);
or U16965 (N_16965,N_16538,N_16637);
nor U16966 (N_16966,N_16717,N_16749);
and U16967 (N_16967,N_16563,N_16511);
nor U16968 (N_16968,N_16701,N_16604);
or U16969 (N_16969,N_16500,N_16732);
nand U16970 (N_16970,N_16533,N_16541);
xor U16971 (N_16971,N_16631,N_16597);
nand U16972 (N_16972,N_16681,N_16563);
nor U16973 (N_16973,N_16653,N_16702);
xor U16974 (N_16974,N_16679,N_16680);
nand U16975 (N_16975,N_16641,N_16674);
nand U16976 (N_16976,N_16632,N_16569);
nor U16977 (N_16977,N_16663,N_16571);
nor U16978 (N_16978,N_16518,N_16651);
nand U16979 (N_16979,N_16639,N_16701);
nor U16980 (N_16980,N_16726,N_16701);
nor U16981 (N_16981,N_16667,N_16642);
and U16982 (N_16982,N_16575,N_16640);
and U16983 (N_16983,N_16680,N_16577);
nor U16984 (N_16984,N_16739,N_16546);
nand U16985 (N_16985,N_16593,N_16741);
xor U16986 (N_16986,N_16581,N_16601);
and U16987 (N_16987,N_16743,N_16574);
xor U16988 (N_16988,N_16632,N_16690);
xor U16989 (N_16989,N_16654,N_16567);
nand U16990 (N_16990,N_16690,N_16553);
nor U16991 (N_16991,N_16610,N_16711);
nor U16992 (N_16992,N_16661,N_16706);
nor U16993 (N_16993,N_16645,N_16731);
nand U16994 (N_16994,N_16558,N_16514);
and U16995 (N_16995,N_16544,N_16566);
nor U16996 (N_16996,N_16538,N_16507);
xor U16997 (N_16997,N_16627,N_16663);
nand U16998 (N_16998,N_16500,N_16697);
nand U16999 (N_16999,N_16627,N_16613);
and U17000 (N_17000,N_16968,N_16796);
and U17001 (N_17001,N_16816,N_16778);
nand U17002 (N_17002,N_16754,N_16821);
xnor U17003 (N_17003,N_16940,N_16767);
and U17004 (N_17004,N_16989,N_16758);
xnor U17005 (N_17005,N_16880,N_16787);
nand U17006 (N_17006,N_16904,N_16813);
nor U17007 (N_17007,N_16994,N_16829);
nor U17008 (N_17008,N_16782,N_16863);
xnor U17009 (N_17009,N_16873,N_16756);
nand U17010 (N_17010,N_16885,N_16900);
and U17011 (N_17011,N_16985,N_16830);
or U17012 (N_17012,N_16814,N_16958);
xor U17013 (N_17013,N_16824,N_16927);
nand U17014 (N_17014,N_16890,N_16934);
nand U17015 (N_17015,N_16941,N_16862);
and U17016 (N_17016,N_16933,N_16954);
or U17017 (N_17017,N_16975,N_16820);
or U17018 (N_17018,N_16929,N_16801);
nor U17019 (N_17019,N_16764,N_16931);
nor U17020 (N_17020,N_16977,N_16834);
and U17021 (N_17021,N_16992,N_16779);
and U17022 (N_17022,N_16917,N_16896);
or U17023 (N_17023,N_16752,N_16938);
nand U17024 (N_17024,N_16979,N_16911);
and U17025 (N_17025,N_16916,N_16860);
and U17026 (N_17026,N_16803,N_16853);
xor U17027 (N_17027,N_16818,N_16851);
nor U17028 (N_17028,N_16867,N_16869);
and U17029 (N_17029,N_16960,N_16770);
or U17030 (N_17030,N_16969,N_16924);
xnor U17031 (N_17031,N_16875,N_16809);
nand U17032 (N_17032,N_16760,N_16769);
or U17033 (N_17033,N_16915,N_16800);
and U17034 (N_17034,N_16850,N_16783);
or U17035 (N_17035,N_16943,N_16974);
or U17036 (N_17036,N_16998,N_16855);
nor U17037 (N_17037,N_16887,N_16847);
xnor U17038 (N_17038,N_16997,N_16861);
nor U17039 (N_17039,N_16775,N_16906);
or U17040 (N_17040,N_16859,N_16806);
or U17041 (N_17041,N_16971,N_16987);
or U17042 (N_17042,N_16976,N_16799);
nor U17043 (N_17043,N_16872,N_16921);
nor U17044 (N_17044,N_16884,N_16902);
and U17045 (N_17045,N_16828,N_16955);
and U17046 (N_17046,N_16848,N_16870);
nor U17047 (N_17047,N_16939,N_16822);
nand U17048 (N_17048,N_16852,N_16983);
and U17049 (N_17049,N_16881,N_16928);
xor U17050 (N_17050,N_16889,N_16792);
or U17051 (N_17051,N_16922,N_16912);
and U17052 (N_17052,N_16951,N_16991);
xor U17053 (N_17053,N_16965,N_16837);
and U17054 (N_17054,N_16956,N_16804);
xor U17055 (N_17055,N_16914,N_16949);
nor U17056 (N_17056,N_16840,N_16894);
xor U17057 (N_17057,N_16795,N_16856);
nor U17058 (N_17058,N_16937,N_16973);
xnor U17059 (N_17059,N_16835,N_16964);
xnor U17060 (N_17060,N_16759,N_16891);
nand U17061 (N_17061,N_16948,N_16945);
and U17062 (N_17062,N_16953,N_16879);
or U17063 (N_17063,N_16751,N_16838);
nor U17064 (N_17064,N_16842,N_16959);
and U17065 (N_17065,N_16961,N_16766);
nand U17066 (N_17066,N_16926,N_16865);
or U17067 (N_17067,N_16876,N_16966);
nand U17068 (N_17068,N_16936,N_16750);
and U17069 (N_17069,N_16999,N_16993);
and U17070 (N_17070,N_16774,N_16980);
and U17071 (N_17071,N_16793,N_16810);
xor U17072 (N_17072,N_16846,N_16892);
or U17073 (N_17073,N_16918,N_16839);
or U17074 (N_17074,N_16845,N_16962);
or U17075 (N_17075,N_16836,N_16970);
or U17076 (N_17076,N_16868,N_16831);
nand U17077 (N_17077,N_16919,N_16753);
and U17078 (N_17078,N_16878,N_16942);
and U17079 (N_17079,N_16802,N_16808);
xor U17080 (N_17080,N_16909,N_16996);
xor U17081 (N_17081,N_16773,N_16776);
nor U17082 (N_17082,N_16882,N_16950);
nand U17083 (N_17083,N_16901,N_16886);
and U17084 (N_17084,N_16858,N_16826);
nand U17085 (N_17085,N_16908,N_16843);
nor U17086 (N_17086,N_16981,N_16925);
xor U17087 (N_17087,N_16898,N_16823);
and U17088 (N_17088,N_16772,N_16967);
and U17089 (N_17089,N_16986,N_16755);
nand U17090 (N_17090,N_16988,N_16794);
xor U17091 (N_17091,N_16946,N_16920);
nand U17092 (N_17092,N_16768,N_16963);
and U17093 (N_17093,N_16789,N_16893);
or U17094 (N_17094,N_16923,N_16888);
nor U17095 (N_17095,N_16947,N_16982);
xnor U17096 (N_17096,N_16930,N_16899);
nand U17097 (N_17097,N_16972,N_16952);
and U17098 (N_17098,N_16798,N_16874);
and U17099 (N_17099,N_16757,N_16788);
nor U17100 (N_17100,N_16765,N_16841);
or U17101 (N_17101,N_16871,N_16854);
nor U17102 (N_17102,N_16781,N_16815);
or U17103 (N_17103,N_16957,N_16897);
and U17104 (N_17104,N_16827,N_16784);
or U17105 (N_17105,N_16978,N_16995);
and U17106 (N_17106,N_16790,N_16812);
nor U17107 (N_17107,N_16944,N_16857);
nand U17108 (N_17108,N_16817,N_16811);
nand U17109 (N_17109,N_16797,N_16895);
xor U17110 (N_17110,N_16761,N_16913);
and U17111 (N_17111,N_16844,N_16763);
nand U17112 (N_17112,N_16990,N_16905);
xnor U17113 (N_17113,N_16805,N_16984);
nor U17114 (N_17114,N_16932,N_16849);
and U17115 (N_17115,N_16780,N_16771);
nor U17116 (N_17116,N_16762,N_16785);
xnor U17117 (N_17117,N_16825,N_16877);
xnor U17118 (N_17118,N_16864,N_16819);
nand U17119 (N_17119,N_16777,N_16903);
and U17120 (N_17120,N_16807,N_16910);
nor U17121 (N_17121,N_16935,N_16786);
or U17122 (N_17122,N_16883,N_16833);
or U17123 (N_17123,N_16866,N_16791);
xor U17124 (N_17124,N_16832,N_16907);
nor U17125 (N_17125,N_16930,N_16888);
xor U17126 (N_17126,N_16928,N_16943);
nor U17127 (N_17127,N_16874,N_16982);
and U17128 (N_17128,N_16958,N_16776);
and U17129 (N_17129,N_16794,N_16805);
nor U17130 (N_17130,N_16811,N_16786);
and U17131 (N_17131,N_16754,N_16879);
and U17132 (N_17132,N_16887,N_16896);
nand U17133 (N_17133,N_16911,N_16843);
nor U17134 (N_17134,N_16757,N_16934);
or U17135 (N_17135,N_16897,N_16969);
nor U17136 (N_17136,N_16975,N_16766);
nand U17137 (N_17137,N_16969,N_16775);
xor U17138 (N_17138,N_16812,N_16772);
or U17139 (N_17139,N_16783,N_16927);
and U17140 (N_17140,N_16998,N_16796);
xor U17141 (N_17141,N_16830,N_16906);
nand U17142 (N_17142,N_16893,N_16968);
and U17143 (N_17143,N_16983,N_16918);
nor U17144 (N_17144,N_16919,N_16956);
xnor U17145 (N_17145,N_16767,N_16952);
xnor U17146 (N_17146,N_16810,N_16775);
nand U17147 (N_17147,N_16864,N_16988);
nand U17148 (N_17148,N_16799,N_16843);
nor U17149 (N_17149,N_16947,N_16890);
nand U17150 (N_17150,N_16981,N_16800);
xor U17151 (N_17151,N_16984,N_16872);
or U17152 (N_17152,N_16842,N_16751);
nor U17153 (N_17153,N_16797,N_16838);
and U17154 (N_17154,N_16791,N_16886);
xor U17155 (N_17155,N_16798,N_16950);
or U17156 (N_17156,N_16882,N_16937);
nand U17157 (N_17157,N_16877,N_16985);
or U17158 (N_17158,N_16837,N_16970);
xnor U17159 (N_17159,N_16752,N_16967);
and U17160 (N_17160,N_16863,N_16986);
nor U17161 (N_17161,N_16846,N_16814);
nor U17162 (N_17162,N_16890,N_16832);
nor U17163 (N_17163,N_16787,N_16777);
or U17164 (N_17164,N_16767,N_16931);
or U17165 (N_17165,N_16863,N_16983);
and U17166 (N_17166,N_16935,N_16913);
xnor U17167 (N_17167,N_16816,N_16834);
nand U17168 (N_17168,N_16963,N_16829);
xor U17169 (N_17169,N_16940,N_16753);
or U17170 (N_17170,N_16868,N_16905);
or U17171 (N_17171,N_16950,N_16969);
xnor U17172 (N_17172,N_16882,N_16767);
or U17173 (N_17173,N_16766,N_16988);
nor U17174 (N_17174,N_16828,N_16807);
nand U17175 (N_17175,N_16958,N_16837);
and U17176 (N_17176,N_16973,N_16992);
and U17177 (N_17177,N_16817,N_16940);
or U17178 (N_17178,N_16977,N_16859);
nand U17179 (N_17179,N_16759,N_16933);
xor U17180 (N_17180,N_16774,N_16956);
or U17181 (N_17181,N_16797,N_16764);
nor U17182 (N_17182,N_16845,N_16820);
xor U17183 (N_17183,N_16913,N_16975);
xor U17184 (N_17184,N_16901,N_16856);
and U17185 (N_17185,N_16983,N_16822);
nor U17186 (N_17186,N_16822,N_16892);
or U17187 (N_17187,N_16829,N_16783);
and U17188 (N_17188,N_16795,N_16840);
nor U17189 (N_17189,N_16830,N_16982);
xor U17190 (N_17190,N_16868,N_16772);
nand U17191 (N_17191,N_16883,N_16917);
xnor U17192 (N_17192,N_16787,N_16973);
nor U17193 (N_17193,N_16751,N_16954);
and U17194 (N_17194,N_16880,N_16763);
xor U17195 (N_17195,N_16940,N_16802);
xnor U17196 (N_17196,N_16787,N_16955);
and U17197 (N_17197,N_16919,N_16984);
and U17198 (N_17198,N_16944,N_16962);
and U17199 (N_17199,N_16904,N_16981);
and U17200 (N_17200,N_16831,N_16810);
or U17201 (N_17201,N_16915,N_16923);
nand U17202 (N_17202,N_16839,N_16802);
xnor U17203 (N_17203,N_16952,N_16905);
xnor U17204 (N_17204,N_16853,N_16891);
or U17205 (N_17205,N_16941,N_16849);
nor U17206 (N_17206,N_16819,N_16992);
nor U17207 (N_17207,N_16792,N_16797);
and U17208 (N_17208,N_16892,N_16954);
xor U17209 (N_17209,N_16991,N_16999);
and U17210 (N_17210,N_16887,N_16784);
and U17211 (N_17211,N_16750,N_16755);
xor U17212 (N_17212,N_16756,N_16849);
and U17213 (N_17213,N_16891,N_16912);
nor U17214 (N_17214,N_16950,N_16783);
nor U17215 (N_17215,N_16990,N_16982);
nand U17216 (N_17216,N_16878,N_16876);
xnor U17217 (N_17217,N_16861,N_16880);
nor U17218 (N_17218,N_16863,N_16815);
or U17219 (N_17219,N_16832,N_16874);
xnor U17220 (N_17220,N_16940,N_16816);
or U17221 (N_17221,N_16868,N_16968);
xor U17222 (N_17222,N_16913,N_16923);
and U17223 (N_17223,N_16913,N_16942);
nor U17224 (N_17224,N_16855,N_16849);
nor U17225 (N_17225,N_16975,N_16895);
and U17226 (N_17226,N_16775,N_16926);
nor U17227 (N_17227,N_16959,N_16893);
xnor U17228 (N_17228,N_16887,N_16874);
xor U17229 (N_17229,N_16799,N_16900);
and U17230 (N_17230,N_16765,N_16896);
nand U17231 (N_17231,N_16776,N_16937);
or U17232 (N_17232,N_16996,N_16807);
nand U17233 (N_17233,N_16927,N_16847);
nand U17234 (N_17234,N_16822,N_16772);
or U17235 (N_17235,N_16846,N_16947);
nor U17236 (N_17236,N_16982,N_16993);
and U17237 (N_17237,N_16876,N_16967);
nand U17238 (N_17238,N_16989,N_16981);
nor U17239 (N_17239,N_16965,N_16808);
and U17240 (N_17240,N_16825,N_16840);
xor U17241 (N_17241,N_16821,N_16753);
xnor U17242 (N_17242,N_16950,N_16772);
or U17243 (N_17243,N_16967,N_16968);
nand U17244 (N_17244,N_16779,N_16807);
xor U17245 (N_17245,N_16898,N_16847);
and U17246 (N_17246,N_16845,N_16991);
nor U17247 (N_17247,N_16806,N_16825);
nor U17248 (N_17248,N_16767,N_16832);
and U17249 (N_17249,N_16920,N_16924);
or U17250 (N_17250,N_17130,N_17048);
or U17251 (N_17251,N_17059,N_17109);
or U17252 (N_17252,N_17168,N_17007);
or U17253 (N_17253,N_17207,N_17002);
xor U17254 (N_17254,N_17176,N_17000);
xnor U17255 (N_17255,N_17053,N_17172);
nor U17256 (N_17256,N_17067,N_17040);
nand U17257 (N_17257,N_17177,N_17061);
or U17258 (N_17258,N_17236,N_17234);
or U17259 (N_17259,N_17088,N_17156);
xnor U17260 (N_17260,N_17235,N_17232);
xnor U17261 (N_17261,N_17237,N_17108);
nor U17262 (N_17262,N_17228,N_17139);
nor U17263 (N_17263,N_17165,N_17239);
or U17264 (N_17264,N_17164,N_17016);
and U17265 (N_17265,N_17141,N_17075);
and U17266 (N_17266,N_17096,N_17204);
nor U17267 (N_17267,N_17062,N_17101);
or U17268 (N_17268,N_17205,N_17224);
xnor U17269 (N_17269,N_17153,N_17039);
nor U17270 (N_17270,N_17084,N_17032);
or U17271 (N_17271,N_17068,N_17226);
nand U17272 (N_17272,N_17098,N_17052);
or U17273 (N_17273,N_17063,N_17134);
xnor U17274 (N_17274,N_17182,N_17083);
nand U17275 (N_17275,N_17227,N_17137);
and U17276 (N_17276,N_17029,N_17217);
xor U17277 (N_17277,N_17192,N_17195);
nand U17278 (N_17278,N_17154,N_17072);
xnor U17279 (N_17279,N_17238,N_17030);
nor U17280 (N_17280,N_17222,N_17246);
or U17281 (N_17281,N_17146,N_17066);
nor U17282 (N_17282,N_17142,N_17221);
or U17283 (N_17283,N_17100,N_17200);
or U17284 (N_17284,N_17212,N_17202);
xnor U17285 (N_17285,N_17116,N_17051);
or U17286 (N_17286,N_17094,N_17206);
xnor U17287 (N_17287,N_17076,N_17189);
xor U17288 (N_17288,N_17035,N_17244);
nor U17289 (N_17289,N_17208,N_17049);
xor U17290 (N_17290,N_17071,N_17230);
and U17291 (N_17291,N_17104,N_17171);
nor U17292 (N_17292,N_17093,N_17057);
or U17293 (N_17293,N_17015,N_17211);
nand U17294 (N_17294,N_17128,N_17127);
or U17295 (N_17295,N_17080,N_17181);
xnor U17296 (N_17296,N_17201,N_17191);
xor U17297 (N_17297,N_17245,N_17106);
xor U17298 (N_17298,N_17023,N_17115);
or U17299 (N_17299,N_17214,N_17095);
or U17300 (N_17300,N_17219,N_17175);
nor U17301 (N_17301,N_17034,N_17112);
nand U17302 (N_17302,N_17097,N_17119);
and U17303 (N_17303,N_17240,N_17132);
or U17304 (N_17304,N_17033,N_17114);
nor U17305 (N_17305,N_17126,N_17113);
or U17306 (N_17306,N_17001,N_17152);
and U17307 (N_17307,N_17184,N_17046);
xnor U17308 (N_17308,N_17010,N_17183);
and U17309 (N_17309,N_17020,N_17178);
xnor U17310 (N_17310,N_17163,N_17225);
nor U17311 (N_17311,N_17055,N_17166);
nor U17312 (N_17312,N_17144,N_17121);
nand U17313 (N_17313,N_17103,N_17131);
xnor U17314 (N_17314,N_17159,N_17138);
xnor U17315 (N_17315,N_17122,N_17149);
nor U17316 (N_17316,N_17118,N_17019);
or U17317 (N_17317,N_17220,N_17092);
nor U17318 (N_17318,N_17161,N_17105);
or U17319 (N_17319,N_17042,N_17162);
nor U17320 (N_17320,N_17243,N_17120);
or U17321 (N_17321,N_17198,N_17008);
xor U17322 (N_17322,N_17107,N_17027);
nand U17323 (N_17323,N_17169,N_17054);
nor U17324 (N_17324,N_17233,N_17117);
or U17325 (N_17325,N_17194,N_17082);
nor U17326 (N_17326,N_17173,N_17148);
or U17327 (N_17327,N_17009,N_17037);
or U17328 (N_17328,N_17151,N_17188);
nand U17329 (N_17329,N_17014,N_17249);
nor U17330 (N_17330,N_17136,N_17058);
nor U17331 (N_17331,N_17036,N_17170);
or U17332 (N_17332,N_17025,N_17209);
nand U17333 (N_17333,N_17038,N_17185);
xnor U17334 (N_17334,N_17160,N_17248);
nand U17335 (N_17335,N_17077,N_17073);
xnor U17336 (N_17336,N_17060,N_17216);
nand U17337 (N_17337,N_17215,N_17099);
nand U17338 (N_17338,N_17123,N_17193);
or U17339 (N_17339,N_17087,N_17086);
or U17340 (N_17340,N_17174,N_17190);
xor U17341 (N_17341,N_17140,N_17125);
nand U17342 (N_17342,N_17223,N_17203);
xnor U17343 (N_17343,N_17158,N_17064);
nand U17344 (N_17344,N_17241,N_17069);
xor U17345 (N_17345,N_17187,N_17018);
nor U17346 (N_17346,N_17147,N_17028);
and U17347 (N_17347,N_17242,N_17213);
xnor U17348 (N_17348,N_17011,N_17089);
nor U17349 (N_17349,N_17047,N_17005);
xnor U17350 (N_17350,N_17197,N_17102);
nand U17351 (N_17351,N_17006,N_17111);
nand U17352 (N_17352,N_17085,N_17179);
xor U17353 (N_17353,N_17056,N_17031);
and U17354 (N_17354,N_17004,N_17078);
and U17355 (N_17355,N_17155,N_17091);
xor U17356 (N_17356,N_17157,N_17090);
and U17357 (N_17357,N_17045,N_17050);
nor U17358 (N_17358,N_17196,N_17145);
nand U17359 (N_17359,N_17021,N_17041);
nor U17360 (N_17360,N_17012,N_17003);
nor U17361 (N_17361,N_17167,N_17124);
xor U17362 (N_17362,N_17229,N_17065);
xnor U17363 (N_17363,N_17135,N_17210);
nand U17364 (N_17364,N_17247,N_17231);
nor U17365 (N_17365,N_17079,N_17017);
or U17366 (N_17366,N_17110,N_17143);
xnor U17367 (N_17367,N_17024,N_17180);
xor U17368 (N_17368,N_17026,N_17218);
and U17369 (N_17369,N_17044,N_17013);
nor U17370 (N_17370,N_17186,N_17129);
nor U17371 (N_17371,N_17081,N_17150);
and U17372 (N_17372,N_17022,N_17133);
and U17373 (N_17373,N_17074,N_17199);
xor U17374 (N_17374,N_17070,N_17043);
or U17375 (N_17375,N_17034,N_17131);
or U17376 (N_17376,N_17031,N_17018);
xor U17377 (N_17377,N_17089,N_17004);
nand U17378 (N_17378,N_17216,N_17011);
or U17379 (N_17379,N_17210,N_17195);
nand U17380 (N_17380,N_17245,N_17156);
xnor U17381 (N_17381,N_17135,N_17206);
xnor U17382 (N_17382,N_17209,N_17190);
nand U17383 (N_17383,N_17017,N_17084);
and U17384 (N_17384,N_17037,N_17188);
nor U17385 (N_17385,N_17125,N_17184);
nor U17386 (N_17386,N_17096,N_17244);
or U17387 (N_17387,N_17186,N_17203);
or U17388 (N_17388,N_17191,N_17104);
nand U17389 (N_17389,N_17245,N_17172);
or U17390 (N_17390,N_17211,N_17204);
and U17391 (N_17391,N_17105,N_17031);
or U17392 (N_17392,N_17233,N_17112);
and U17393 (N_17393,N_17197,N_17160);
nand U17394 (N_17394,N_17119,N_17146);
and U17395 (N_17395,N_17092,N_17182);
nor U17396 (N_17396,N_17058,N_17064);
or U17397 (N_17397,N_17006,N_17145);
and U17398 (N_17398,N_17090,N_17089);
xor U17399 (N_17399,N_17195,N_17029);
and U17400 (N_17400,N_17193,N_17243);
or U17401 (N_17401,N_17051,N_17102);
or U17402 (N_17402,N_17221,N_17062);
xor U17403 (N_17403,N_17016,N_17143);
xor U17404 (N_17404,N_17199,N_17235);
nand U17405 (N_17405,N_17219,N_17028);
or U17406 (N_17406,N_17134,N_17041);
and U17407 (N_17407,N_17125,N_17177);
and U17408 (N_17408,N_17024,N_17217);
nor U17409 (N_17409,N_17004,N_17226);
xnor U17410 (N_17410,N_17205,N_17121);
nand U17411 (N_17411,N_17214,N_17030);
nand U17412 (N_17412,N_17079,N_17225);
nor U17413 (N_17413,N_17068,N_17071);
nand U17414 (N_17414,N_17076,N_17217);
xnor U17415 (N_17415,N_17217,N_17064);
or U17416 (N_17416,N_17032,N_17015);
or U17417 (N_17417,N_17004,N_17043);
or U17418 (N_17418,N_17155,N_17172);
or U17419 (N_17419,N_17224,N_17170);
or U17420 (N_17420,N_17020,N_17068);
nor U17421 (N_17421,N_17234,N_17083);
xnor U17422 (N_17422,N_17115,N_17034);
or U17423 (N_17423,N_17240,N_17121);
nand U17424 (N_17424,N_17028,N_17048);
or U17425 (N_17425,N_17240,N_17247);
xnor U17426 (N_17426,N_17131,N_17056);
xor U17427 (N_17427,N_17044,N_17033);
and U17428 (N_17428,N_17157,N_17134);
nand U17429 (N_17429,N_17189,N_17002);
and U17430 (N_17430,N_17156,N_17030);
xor U17431 (N_17431,N_17149,N_17060);
or U17432 (N_17432,N_17190,N_17221);
and U17433 (N_17433,N_17227,N_17230);
nor U17434 (N_17434,N_17228,N_17193);
nor U17435 (N_17435,N_17129,N_17123);
nand U17436 (N_17436,N_17246,N_17217);
nand U17437 (N_17437,N_17024,N_17068);
xor U17438 (N_17438,N_17028,N_17044);
nand U17439 (N_17439,N_17116,N_17113);
nor U17440 (N_17440,N_17156,N_17145);
or U17441 (N_17441,N_17113,N_17206);
or U17442 (N_17442,N_17209,N_17073);
or U17443 (N_17443,N_17145,N_17130);
nand U17444 (N_17444,N_17123,N_17151);
and U17445 (N_17445,N_17160,N_17224);
or U17446 (N_17446,N_17010,N_17098);
or U17447 (N_17447,N_17087,N_17114);
nor U17448 (N_17448,N_17160,N_17045);
xor U17449 (N_17449,N_17177,N_17236);
nand U17450 (N_17450,N_17051,N_17153);
nand U17451 (N_17451,N_17165,N_17248);
nor U17452 (N_17452,N_17084,N_17151);
and U17453 (N_17453,N_17170,N_17181);
xor U17454 (N_17454,N_17165,N_17011);
or U17455 (N_17455,N_17189,N_17210);
nor U17456 (N_17456,N_17019,N_17032);
or U17457 (N_17457,N_17046,N_17121);
or U17458 (N_17458,N_17136,N_17104);
xor U17459 (N_17459,N_17014,N_17079);
xnor U17460 (N_17460,N_17211,N_17125);
and U17461 (N_17461,N_17144,N_17072);
or U17462 (N_17462,N_17214,N_17189);
nor U17463 (N_17463,N_17109,N_17091);
nor U17464 (N_17464,N_17034,N_17055);
and U17465 (N_17465,N_17142,N_17018);
nand U17466 (N_17466,N_17192,N_17084);
and U17467 (N_17467,N_17050,N_17065);
and U17468 (N_17468,N_17201,N_17142);
nor U17469 (N_17469,N_17028,N_17235);
or U17470 (N_17470,N_17071,N_17043);
nand U17471 (N_17471,N_17197,N_17106);
xnor U17472 (N_17472,N_17188,N_17195);
xnor U17473 (N_17473,N_17058,N_17072);
or U17474 (N_17474,N_17112,N_17244);
nand U17475 (N_17475,N_17164,N_17235);
xnor U17476 (N_17476,N_17180,N_17212);
or U17477 (N_17477,N_17043,N_17057);
nand U17478 (N_17478,N_17172,N_17147);
or U17479 (N_17479,N_17245,N_17157);
and U17480 (N_17480,N_17093,N_17030);
or U17481 (N_17481,N_17075,N_17185);
nand U17482 (N_17482,N_17051,N_17216);
nor U17483 (N_17483,N_17165,N_17023);
and U17484 (N_17484,N_17161,N_17032);
or U17485 (N_17485,N_17206,N_17127);
nand U17486 (N_17486,N_17043,N_17226);
nor U17487 (N_17487,N_17166,N_17010);
xnor U17488 (N_17488,N_17245,N_17185);
nor U17489 (N_17489,N_17153,N_17234);
and U17490 (N_17490,N_17063,N_17210);
or U17491 (N_17491,N_17213,N_17085);
xor U17492 (N_17492,N_17153,N_17049);
nor U17493 (N_17493,N_17221,N_17181);
or U17494 (N_17494,N_17045,N_17114);
nand U17495 (N_17495,N_17102,N_17156);
and U17496 (N_17496,N_17096,N_17169);
nand U17497 (N_17497,N_17115,N_17227);
or U17498 (N_17498,N_17244,N_17095);
and U17499 (N_17499,N_17178,N_17201);
or U17500 (N_17500,N_17325,N_17295);
or U17501 (N_17501,N_17265,N_17417);
nand U17502 (N_17502,N_17492,N_17474);
nor U17503 (N_17503,N_17268,N_17305);
nand U17504 (N_17504,N_17348,N_17278);
xnor U17505 (N_17505,N_17300,N_17387);
or U17506 (N_17506,N_17264,N_17297);
nand U17507 (N_17507,N_17323,N_17369);
and U17508 (N_17508,N_17448,N_17440);
nor U17509 (N_17509,N_17306,N_17280);
and U17510 (N_17510,N_17496,N_17463);
nand U17511 (N_17511,N_17490,N_17371);
nand U17512 (N_17512,N_17449,N_17415);
nor U17513 (N_17513,N_17255,N_17303);
or U17514 (N_17514,N_17324,N_17466);
nor U17515 (N_17515,N_17365,N_17291);
and U17516 (N_17516,N_17376,N_17453);
xor U17517 (N_17517,N_17311,N_17360);
nor U17518 (N_17518,N_17420,N_17361);
nor U17519 (N_17519,N_17283,N_17436);
nor U17520 (N_17520,N_17298,N_17428);
xnor U17521 (N_17521,N_17368,N_17259);
xor U17522 (N_17522,N_17335,N_17254);
or U17523 (N_17523,N_17481,N_17334);
or U17524 (N_17524,N_17251,N_17435);
and U17525 (N_17525,N_17364,N_17427);
nand U17526 (N_17526,N_17263,N_17434);
xor U17527 (N_17527,N_17310,N_17464);
or U17528 (N_17528,N_17388,N_17408);
nand U17529 (N_17529,N_17421,N_17363);
nor U17530 (N_17530,N_17358,N_17416);
xnor U17531 (N_17531,N_17478,N_17469);
xnor U17532 (N_17532,N_17273,N_17275);
and U17533 (N_17533,N_17461,N_17269);
xnor U17534 (N_17534,N_17451,N_17362);
nand U17535 (N_17535,N_17484,N_17397);
nor U17536 (N_17536,N_17431,N_17250);
or U17537 (N_17537,N_17332,N_17302);
and U17538 (N_17538,N_17320,N_17336);
or U17539 (N_17539,N_17487,N_17445);
and U17540 (N_17540,N_17344,N_17418);
nand U17541 (N_17541,N_17382,N_17472);
and U17542 (N_17542,N_17425,N_17375);
xor U17543 (N_17543,N_17411,N_17488);
nand U17544 (N_17544,N_17489,N_17292);
nand U17545 (N_17545,N_17404,N_17422);
nand U17546 (N_17546,N_17483,N_17351);
and U17547 (N_17547,N_17390,N_17491);
xnor U17548 (N_17548,N_17257,N_17341);
or U17549 (N_17549,N_17367,N_17270);
and U17550 (N_17550,N_17442,N_17424);
xnor U17551 (N_17551,N_17260,N_17477);
nor U17552 (N_17552,N_17346,N_17467);
nor U17553 (N_17553,N_17296,N_17359);
and U17554 (N_17554,N_17372,N_17252);
or U17555 (N_17555,N_17340,N_17406);
and U17556 (N_17556,N_17392,N_17389);
nor U17557 (N_17557,N_17309,N_17437);
nor U17558 (N_17558,N_17462,N_17316);
or U17559 (N_17559,N_17274,N_17498);
xnor U17560 (N_17560,N_17399,N_17284);
nand U17561 (N_17561,N_17494,N_17383);
xnor U17562 (N_17562,N_17315,N_17384);
nand U17563 (N_17563,N_17357,N_17267);
or U17564 (N_17564,N_17258,N_17379);
and U17565 (N_17565,N_17345,N_17401);
nor U17566 (N_17566,N_17452,N_17419);
nand U17567 (N_17567,N_17301,N_17285);
nand U17568 (N_17568,N_17370,N_17433);
nand U17569 (N_17569,N_17349,N_17286);
nor U17570 (N_17570,N_17398,N_17499);
xnor U17571 (N_17571,N_17331,N_17430);
xnor U17572 (N_17572,N_17454,N_17455);
xor U17573 (N_17573,N_17465,N_17410);
or U17574 (N_17574,N_17458,N_17327);
and U17575 (N_17575,N_17429,N_17308);
or U17576 (N_17576,N_17378,N_17386);
nand U17577 (N_17577,N_17480,N_17329);
or U17578 (N_17578,N_17317,N_17288);
nand U17579 (N_17579,N_17272,N_17441);
nand U17580 (N_17580,N_17266,N_17405);
nand U17581 (N_17581,N_17289,N_17460);
xor U17582 (N_17582,N_17374,N_17333);
xnor U17583 (N_17583,N_17319,N_17432);
and U17584 (N_17584,N_17328,N_17318);
nor U17585 (N_17585,N_17337,N_17281);
or U17586 (N_17586,N_17400,N_17443);
xnor U17587 (N_17587,N_17261,N_17407);
nor U17588 (N_17588,N_17380,N_17394);
nand U17589 (N_17589,N_17299,N_17256);
nand U17590 (N_17590,N_17347,N_17476);
nand U17591 (N_17591,N_17497,N_17438);
nand U17592 (N_17592,N_17343,N_17470);
and U17593 (N_17593,N_17447,N_17293);
nand U17594 (N_17594,N_17486,N_17271);
and U17595 (N_17595,N_17353,N_17444);
and U17596 (N_17596,N_17413,N_17355);
nand U17597 (N_17597,N_17356,N_17312);
nand U17598 (N_17598,N_17402,N_17450);
nor U17599 (N_17599,N_17294,N_17409);
xor U17600 (N_17600,N_17479,N_17473);
nor U17601 (N_17601,N_17457,N_17253);
nand U17602 (N_17602,N_17339,N_17373);
nand U17603 (N_17603,N_17338,N_17446);
and U17604 (N_17604,N_17262,N_17350);
xnor U17605 (N_17605,N_17352,N_17495);
nand U17606 (N_17606,N_17426,N_17314);
xnor U17607 (N_17607,N_17414,N_17482);
nor U17608 (N_17608,N_17304,N_17330);
and U17609 (N_17609,N_17468,N_17276);
nand U17610 (N_17610,N_17475,N_17485);
nand U17611 (N_17611,N_17321,N_17366);
nand U17612 (N_17612,N_17287,N_17322);
and U17613 (N_17613,N_17385,N_17423);
and U17614 (N_17614,N_17277,N_17456);
or U17615 (N_17615,N_17307,N_17396);
xor U17616 (N_17616,N_17381,N_17459);
nand U17617 (N_17617,N_17393,N_17342);
nor U17618 (N_17618,N_17471,N_17493);
nor U17619 (N_17619,N_17279,N_17412);
and U17620 (N_17620,N_17290,N_17326);
and U17621 (N_17621,N_17439,N_17282);
nand U17622 (N_17622,N_17403,N_17354);
nand U17623 (N_17623,N_17391,N_17395);
xor U17624 (N_17624,N_17313,N_17377);
xnor U17625 (N_17625,N_17387,N_17329);
or U17626 (N_17626,N_17462,N_17300);
and U17627 (N_17627,N_17320,N_17293);
and U17628 (N_17628,N_17311,N_17326);
xnor U17629 (N_17629,N_17410,N_17437);
xnor U17630 (N_17630,N_17384,N_17253);
and U17631 (N_17631,N_17261,N_17442);
nor U17632 (N_17632,N_17252,N_17431);
and U17633 (N_17633,N_17358,N_17331);
or U17634 (N_17634,N_17439,N_17322);
xor U17635 (N_17635,N_17393,N_17296);
nand U17636 (N_17636,N_17454,N_17334);
or U17637 (N_17637,N_17343,N_17429);
xnor U17638 (N_17638,N_17453,N_17284);
and U17639 (N_17639,N_17478,N_17369);
nand U17640 (N_17640,N_17326,N_17476);
nand U17641 (N_17641,N_17465,N_17463);
or U17642 (N_17642,N_17455,N_17485);
and U17643 (N_17643,N_17345,N_17272);
and U17644 (N_17644,N_17466,N_17464);
and U17645 (N_17645,N_17285,N_17394);
xnor U17646 (N_17646,N_17492,N_17264);
or U17647 (N_17647,N_17289,N_17304);
and U17648 (N_17648,N_17252,N_17257);
and U17649 (N_17649,N_17449,N_17445);
xnor U17650 (N_17650,N_17262,N_17495);
xor U17651 (N_17651,N_17250,N_17348);
xor U17652 (N_17652,N_17315,N_17480);
xnor U17653 (N_17653,N_17465,N_17260);
nand U17654 (N_17654,N_17343,N_17375);
and U17655 (N_17655,N_17399,N_17290);
or U17656 (N_17656,N_17355,N_17489);
nor U17657 (N_17657,N_17362,N_17307);
or U17658 (N_17658,N_17307,N_17489);
nor U17659 (N_17659,N_17437,N_17252);
nor U17660 (N_17660,N_17380,N_17422);
nor U17661 (N_17661,N_17323,N_17294);
or U17662 (N_17662,N_17295,N_17345);
and U17663 (N_17663,N_17312,N_17441);
or U17664 (N_17664,N_17320,N_17386);
or U17665 (N_17665,N_17263,N_17470);
nor U17666 (N_17666,N_17282,N_17497);
or U17667 (N_17667,N_17422,N_17390);
nand U17668 (N_17668,N_17499,N_17400);
nor U17669 (N_17669,N_17337,N_17346);
nor U17670 (N_17670,N_17330,N_17498);
nand U17671 (N_17671,N_17491,N_17278);
nand U17672 (N_17672,N_17415,N_17478);
xnor U17673 (N_17673,N_17276,N_17330);
nor U17674 (N_17674,N_17320,N_17481);
and U17675 (N_17675,N_17310,N_17286);
nand U17676 (N_17676,N_17455,N_17422);
nand U17677 (N_17677,N_17352,N_17485);
nor U17678 (N_17678,N_17406,N_17369);
xor U17679 (N_17679,N_17291,N_17436);
nand U17680 (N_17680,N_17404,N_17430);
xor U17681 (N_17681,N_17447,N_17423);
nand U17682 (N_17682,N_17419,N_17341);
xnor U17683 (N_17683,N_17321,N_17497);
nand U17684 (N_17684,N_17286,N_17466);
and U17685 (N_17685,N_17264,N_17326);
nand U17686 (N_17686,N_17460,N_17308);
nand U17687 (N_17687,N_17447,N_17465);
nand U17688 (N_17688,N_17476,N_17356);
xnor U17689 (N_17689,N_17427,N_17476);
and U17690 (N_17690,N_17279,N_17482);
xnor U17691 (N_17691,N_17274,N_17261);
nand U17692 (N_17692,N_17308,N_17379);
or U17693 (N_17693,N_17394,N_17474);
nand U17694 (N_17694,N_17255,N_17277);
or U17695 (N_17695,N_17284,N_17328);
and U17696 (N_17696,N_17433,N_17369);
and U17697 (N_17697,N_17460,N_17450);
nor U17698 (N_17698,N_17304,N_17251);
or U17699 (N_17699,N_17318,N_17476);
nor U17700 (N_17700,N_17412,N_17409);
or U17701 (N_17701,N_17310,N_17448);
nand U17702 (N_17702,N_17480,N_17482);
xnor U17703 (N_17703,N_17496,N_17378);
nor U17704 (N_17704,N_17459,N_17263);
or U17705 (N_17705,N_17398,N_17430);
nor U17706 (N_17706,N_17281,N_17394);
nor U17707 (N_17707,N_17270,N_17411);
nor U17708 (N_17708,N_17394,N_17298);
nand U17709 (N_17709,N_17437,N_17373);
nor U17710 (N_17710,N_17442,N_17380);
nand U17711 (N_17711,N_17437,N_17374);
or U17712 (N_17712,N_17421,N_17385);
xor U17713 (N_17713,N_17254,N_17482);
nand U17714 (N_17714,N_17309,N_17344);
xor U17715 (N_17715,N_17422,N_17376);
nor U17716 (N_17716,N_17408,N_17478);
nand U17717 (N_17717,N_17383,N_17277);
and U17718 (N_17718,N_17252,N_17282);
and U17719 (N_17719,N_17272,N_17447);
nor U17720 (N_17720,N_17282,N_17331);
nand U17721 (N_17721,N_17257,N_17387);
or U17722 (N_17722,N_17301,N_17450);
nor U17723 (N_17723,N_17481,N_17250);
nor U17724 (N_17724,N_17494,N_17296);
nand U17725 (N_17725,N_17316,N_17411);
and U17726 (N_17726,N_17349,N_17354);
and U17727 (N_17727,N_17356,N_17295);
nor U17728 (N_17728,N_17388,N_17266);
and U17729 (N_17729,N_17256,N_17400);
xor U17730 (N_17730,N_17403,N_17435);
and U17731 (N_17731,N_17377,N_17281);
and U17732 (N_17732,N_17302,N_17266);
or U17733 (N_17733,N_17361,N_17326);
nor U17734 (N_17734,N_17429,N_17446);
nor U17735 (N_17735,N_17320,N_17451);
nor U17736 (N_17736,N_17438,N_17283);
xnor U17737 (N_17737,N_17334,N_17286);
or U17738 (N_17738,N_17452,N_17329);
or U17739 (N_17739,N_17342,N_17475);
and U17740 (N_17740,N_17422,N_17442);
nor U17741 (N_17741,N_17373,N_17319);
or U17742 (N_17742,N_17255,N_17402);
xor U17743 (N_17743,N_17429,N_17404);
and U17744 (N_17744,N_17403,N_17483);
nor U17745 (N_17745,N_17306,N_17314);
and U17746 (N_17746,N_17415,N_17466);
or U17747 (N_17747,N_17282,N_17483);
nor U17748 (N_17748,N_17488,N_17349);
nor U17749 (N_17749,N_17308,N_17486);
nand U17750 (N_17750,N_17611,N_17622);
xnor U17751 (N_17751,N_17659,N_17654);
nor U17752 (N_17752,N_17679,N_17607);
or U17753 (N_17753,N_17672,N_17665);
xor U17754 (N_17754,N_17558,N_17512);
and U17755 (N_17755,N_17710,N_17734);
nor U17756 (N_17756,N_17623,N_17691);
nor U17757 (N_17757,N_17674,N_17714);
nand U17758 (N_17758,N_17618,N_17598);
xnor U17759 (N_17759,N_17636,N_17732);
and U17760 (N_17760,N_17564,N_17548);
nand U17761 (N_17761,N_17528,N_17725);
and U17762 (N_17762,N_17637,N_17695);
nor U17763 (N_17763,N_17740,N_17612);
xnor U17764 (N_17764,N_17680,N_17671);
nor U17765 (N_17765,N_17524,N_17572);
nor U17766 (N_17766,N_17509,N_17707);
nor U17767 (N_17767,N_17538,N_17583);
and U17768 (N_17768,N_17621,N_17689);
and U17769 (N_17769,N_17566,N_17660);
xor U17770 (N_17770,N_17573,N_17577);
or U17771 (N_17771,N_17617,N_17615);
nor U17772 (N_17772,N_17709,N_17711);
nor U17773 (N_17773,N_17744,N_17624);
or U17774 (N_17774,N_17690,N_17669);
nor U17775 (N_17775,N_17545,N_17597);
xor U17776 (N_17776,N_17535,N_17634);
or U17777 (N_17777,N_17543,N_17626);
nand U17778 (N_17778,N_17653,N_17556);
nor U17779 (N_17779,N_17571,N_17736);
xor U17780 (N_17780,N_17557,N_17526);
and U17781 (N_17781,N_17505,N_17640);
nor U17782 (N_17782,N_17688,N_17609);
or U17783 (N_17783,N_17718,N_17681);
nand U17784 (N_17784,N_17638,N_17602);
nor U17785 (N_17785,N_17693,N_17510);
or U17786 (N_17786,N_17601,N_17507);
nor U17787 (N_17787,N_17514,N_17614);
nand U17788 (N_17788,N_17673,N_17629);
xnor U17789 (N_17789,N_17731,N_17733);
nand U17790 (N_17790,N_17503,N_17704);
and U17791 (N_17791,N_17508,N_17519);
xnor U17792 (N_17792,N_17720,N_17668);
or U17793 (N_17793,N_17588,N_17708);
xor U17794 (N_17794,N_17747,N_17596);
and U17795 (N_17795,N_17703,N_17523);
or U17796 (N_17796,N_17527,N_17540);
or U17797 (N_17797,N_17698,N_17646);
nand U17798 (N_17798,N_17730,N_17506);
or U17799 (N_17799,N_17666,N_17518);
xor U17800 (N_17800,N_17534,N_17628);
xor U17801 (N_17801,N_17586,N_17715);
and U17802 (N_17802,N_17678,N_17530);
nor U17803 (N_17803,N_17592,N_17748);
xor U17804 (N_17804,N_17589,N_17656);
and U17805 (N_17805,N_17594,N_17677);
nand U17806 (N_17806,N_17664,N_17702);
and U17807 (N_17807,N_17726,N_17570);
and U17808 (N_17808,N_17619,N_17745);
nand U17809 (N_17809,N_17717,N_17576);
and U17810 (N_17810,N_17502,N_17737);
xnor U17811 (N_17811,N_17661,N_17608);
xor U17812 (N_17812,N_17501,N_17743);
xor U17813 (N_17813,N_17521,N_17610);
xor U17814 (N_17814,N_17712,N_17716);
and U17815 (N_17815,N_17539,N_17599);
or U17816 (N_17816,N_17560,N_17549);
xor U17817 (N_17817,N_17613,N_17699);
xor U17818 (N_17818,N_17682,N_17579);
nor U17819 (N_17819,N_17537,N_17649);
xor U17820 (N_17820,N_17705,N_17516);
nor U17821 (N_17821,N_17542,N_17605);
xor U17822 (N_17822,N_17676,N_17627);
nor U17823 (N_17823,N_17580,N_17749);
nand U17824 (N_17824,N_17544,N_17500);
and U17825 (N_17825,N_17670,N_17728);
xor U17826 (N_17826,N_17517,N_17675);
nor U17827 (N_17827,N_17722,N_17551);
nand U17828 (N_17828,N_17729,N_17727);
nor U17829 (N_17829,N_17643,N_17706);
nor U17830 (N_17830,N_17520,N_17658);
xnor U17831 (N_17831,N_17546,N_17721);
and U17832 (N_17832,N_17522,N_17569);
nand U17833 (N_17833,N_17567,N_17600);
nand U17834 (N_17834,N_17531,N_17585);
or U17835 (N_17835,N_17511,N_17581);
or U17836 (N_17836,N_17735,N_17723);
or U17837 (N_17837,N_17687,N_17562);
nand U17838 (N_17838,N_17741,N_17639);
xnor U17839 (N_17839,N_17552,N_17642);
nand U17840 (N_17840,N_17593,N_17713);
nor U17841 (N_17841,N_17697,N_17606);
xnor U17842 (N_17842,N_17561,N_17550);
xnor U17843 (N_17843,N_17700,N_17604);
nor U17844 (N_17844,N_17587,N_17515);
nand U17845 (N_17845,N_17635,N_17529);
and U17846 (N_17846,N_17686,N_17647);
nor U17847 (N_17847,N_17590,N_17625);
nor U17848 (N_17848,N_17648,N_17667);
xnor U17849 (N_17849,N_17632,N_17739);
nor U17850 (N_17850,N_17633,N_17631);
xnor U17851 (N_17851,N_17746,N_17701);
nor U17852 (N_17852,N_17504,N_17541);
nor U17853 (N_17853,N_17554,N_17692);
nor U17854 (N_17854,N_17513,N_17651);
or U17855 (N_17855,N_17652,N_17657);
or U17856 (N_17856,N_17641,N_17591);
or U17857 (N_17857,N_17582,N_17645);
and U17858 (N_17858,N_17724,N_17547);
and U17859 (N_17859,N_17655,N_17738);
nand U17860 (N_17860,N_17696,N_17663);
and U17861 (N_17861,N_17595,N_17616);
nor U17862 (N_17862,N_17650,N_17563);
or U17863 (N_17863,N_17684,N_17532);
xor U17864 (N_17864,N_17555,N_17533);
nand U17865 (N_17865,N_17630,N_17584);
nand U17866 (N_17866,N_17694,N_17685);
and U17867 (N_17867,N_17603,N_17719);
or U17868 (N_17868,N_17553,N_17620);
xor U17869 (N_17869,N_17575,N_17568);
and U17870 (N_17870,N_17536,N_17742);
and U17871 (N_17871,N_17559,N_17578);
nand U17872 (N_17872,N_17662,N_17683);
xnor U17873 (N_17873,N_17565,N_17574);
xnor U17874 (N_17874,N_17644,N_17525);
xnor U17875 (N_17875,N_17670,N_17691);
and U17876 (N_17876,N_17745,N_17567);
nor U17877 (N_17877,N_17604,N_17624);
nand U17878 (N_17878,N_17584,N_17667);
nor U17879 (N_17879,N_17592,N_17647);
nor U17880 (N_17880,N_17568,N_17620);
and U17881 (N_17881,N_17664,N_17649);
and U17882 (N_17882,N_17559,N_17560);
and U17883 (N_17883,N_17518,N_17526);
xnor U17884 (N_17884,N_17500,N_17640);
or U17885 (N_17885,N_17555,N_17621);
and U17886 (N_17886,N_17650,N_17559);
nand U17887 (N_17887,N_17589,N_17598);
or U17888 (N_17888,N_17711,N_17514);
and U17889 (N_17889,N_17606,N_17578);
nand U17890 (N_17890,N_17583,N_17533);
nand U17891 (N_17891,N_17527,N_17622);
and U17892 (N_17892,N_17668,N_17728);
and U17893 (N_17893,N_17592,N_17502);
nor U17894 (N_17894,N_17534,N_17560);
and U17895 (N_17895,N_17562,N_17538);
or U17896 (N_17896,N_17501,N_17539);
and U17897 (N_17897,N_17713,N_17536);
nor U17898 (N_17898,N_17594,N_17748);
or U17899 (N_17899,N_17731,N_17669);
nor U17900 (N_17900,N_17501,N_17708);
nor U17901 (N_17901,N_17518,N_17721);
xor U17902 (N_17902,N_17562,N_17722);
xnor U17903 (N_17903,N_17667,N_17597);
xor U17904 (N_17904,N_17741,N_17700);
nand U17905 (N_17905,N_17629,N_17687);
nand U17906 (N_17906,N_17668,N_17623);
xnor U17907 (N_17907,N_17556,N_17630);
and U17908 (N_17908,N_17666,N_17586);
nor U17909 (N_17909,N_17652,N_17656);
or U17910 (N_17910,N_17558,N_17621);
and U17911 (N_17911,N_17552,N_17578);
and U17912 (N_17912,N_17555,N_17650);
or U17913 (N_17913,N_17634,N_17626);
or U17914 (N_17914,N_17671,N_17531);
nand U17915 (N_17915,N_17679,N_17614);
or U17916 (N_17916,N_17625,N_17704);
and U17917 (N_17917,N_17596,N_17748);
and U17918 (N_17918,N_17525,N_17653);
nor U17919 (N_17919,N_17622,N_17660);
and U17920 (N_17920,N_17701,N_17691);
or U17921 (N_17921,N_17600,N_17735);
nand U17922 (N_17922,N_17733,N_17638);
nor U17923 (N_17923,N_17621,N_17533);
nor U17924 (N_17924,N_17676,N_17514);
nand U17925 (N_17925,N_17639,N_17727);
nor U17926 (N_17926,N_17547,N_17693);
nand U17927 (N_17927,N_17622,N_17733);
nor U17928 (N_17928,N_17550,N_17664);
xnor U17929 (N_17929,N_17717,N_17547);
nand U17930 (N_17930,N_17605,N_17524);
nor U17931 (N_17931,N_17589,N_17719);
nor U17932 (N_17932,N_17599,N_17679);
or U17933 (N_17933,N_17503,N_17747);
nor U17934 (N_17934,N_17651,N_17731);
and U17935 (N_17935,N_17713,N_17541);
and U17936 (N_17936,N_17575,N_17540);
or U17937 (N_17937,N_17722,N_17554);
xor U17938 (N_17938,N_17506,N_17654);
nand U17939 (N_17939,N_17729,N_17550);
or U17940 (N_17940,N_17600,N_17731);
or U17941 (N_17941,N_17536,N_17587);
xnor U17942 (N_17942,N_17649,N_17689);
or U17943 (N_17943,N_17550,N_17720);
nand U17944 (N_17944,N_17568,N_17607);
or U17945 (N_17945,N_17665,N_17685);
xor U17946 (N_17946,N_17650,N_17537);
and U17947 (N_17947,N_17661,N_17576);
nor U17948 (N_17948,N_17637,N_17743);
nor U17949 (N_17949,N_17696,N_17588);
nand U17950 (N_17950,N_17566,N_17702);
xor U17951 (N_17951,N_17564,N_17569);
nor U17952 (N_17952,N_17564,N_17743);
nand U17953 (N_17953,N_17700,N_17701);
and U17954 (N_17954,N_17552,N_17504);
or U17955 (N_17955,N_17684,N_17516);
nand U17956 (N_17956,N_17633,N_17585);
xor U17957 (N_17957,N_17746,N_17566);
or U17958 (N_17958,N_17655,N_17692);
or U17959 (N_17959,N_17702,N_17716);
xor U17960 (N_17960,N_17679,N_17556);
and U17961 (N_17961,N_17699,N_17522);
nand U17962 (N_17962,N_17501,N_17626);
and U17963 (N_17963,N_17515,N_17625);
nand U17964 (N_17964,N_17714,N_17562);
nor U17965 (N_17965,N_17626,N_17723);
nor U17966 (N_17966,N_17625,N_17725);
nand U17967 (N_17967,N_17735,N_17625);
nand U17968 (N_17968,N_17581,N_17685);
xor U17969 (N_17969,N_17557,N_17528);
or U17970 (N_17970,N_17675,N_17547);
nand U17971 (N_17971,N_17692,N_17642);
nor U17972 (N_17972,N_17541,N_17677);
nand U17973 (N_17973,N_17701,N_17594);
xnor U17974 (N_17974,N_17716,N_17744);
nor U17975 (N_17975,N_17728,N_17615);
nor U17976 (N_17976,N_17653,N_17558);
and U17977 (N_17977,N_17630,N_17501);
or U17978 (N_17978,N_17522,N_17589);
or U17979 (N_17979,N_17571,N_17574);
xor U17980 (N_17980,N_17644,N_17636);
or U17981 (N_17981,N_17547,N_17620);
or U17982 (N_17982,N_17684,N_17554);
and U17983 (N_17983,N_17512,N_17587);
nand U17984 (N_17984,N_17620,N_17515);
nor U17985 (N_17985,N_17678,N_17524);
nor U17986 (N_17986,N_17663,N_17587);
nor U17987 (N_17987,N_17724,N_17540);
nor U17988 (N_17988,N_17733,N_17739);
nor U17989 (N_17989,N_17526,N_17644);
xor U17990 (N_17990,N_17670,N_17699);
nand U17991 (N_17991,N_17632,N_17730);
and U17992 (N_17992,N_17574,N_17523);
or U17993 (N_17993,N_17506,N_17747);
or U17994 (N_17994,N_17538,N_17669);
nand U17995 (N_17995,N_17676,N_17653);
nor U17996 (N_17996,N_17702,N_17649);
nor U17997 (N_17997,N_17660,N_17507);
or U17998 (N_17998,N_17514,N_17640);
or U17999 (N_17999,N_17674,N_17552);
xor U18000 (N_18000,N_17976,N_17879);
xnor U18001 (N_18001,N_17758,N_17818);
and U18002 (N_18002,N_17851,N_17896);
nor U18003 (N_18003,N_17826,N_17905);
or U18004 (N_18004,N_17787,N_17969);
and U18005 (N_18005,N_17836,N_17858);
xor U18006 (N_18006,N_17775,N_17980);
nand U18007 (N_18007,N_17800,N_17906);
nor U18008 (N_18008,N_17952,N_17845);
nor U18009 (N_18009,N_17861,N_17856);
nand U18010 (N_18010,N_17789,N_17997);
or U18011 (N_18011,N_17982,N_17949);
nand U18012 (N_18012,N_17967,N_17784);
nand U18013 (N_18013,N_17971,N_17773);
xor U18014 (N_18014,N_17790,N_17791);
nor U18015 (N_18015,N_17860,N_17972);
and U18016 (N_18016,N_17804,N_17857);
or U18017 (N_18017,N_17943,N_17844);
xor U18018 (N_18018,N_17957,N_17958);
nand U18019 (N_18019,N_17799,N_17812);
xor U18020 (N_18020,N_17985,N_17920);
and U18021 (N_18021,N_17829,N_17961);
nor U18022 (N_18022,N_17966,N_17876);
and U18023 (N_18023,N_17869,N_17960);
and U18024 (N_18024,N_17864,N_17802);
and U18025 (N_18025,N_17898,N_17763);
nand U18026 (N_18026,N_17835,N_17877);
xor U18027 (N_18027,N_17926,N_17813);
xnor U18028 (N_18028,N_17897,N_17837);
xnor U18029 (N_18029,N_17820,N_17852);
xor U18030 (N_18030,N_17930,N_17783);
nand U18031 (N_18031,N_17965,N_17766);
or U18032 (N_18032,N_17963,N_17817);
and U18033 (N_18033,N_17811,N_17939);
xnor U18034 (N_18034,N_17995,N_17915);
nor U18035 (N_18035,N_17803,N_17979);
nand U18036 (N_18036,N_17993,N_17824);
nor U18037 (N_18037,N_17873,N_17999);
nor U18038 (N_18038,N_17848,N_17942);
xor U18039 (N_18039,N_17927,N_17987);
and U18040 (N_18040,N_17975,N_17878);
xnor U18041 (N_18041,N_17956,N_17925);
nand U18042 (N_18042,N_17941,N_17838);
xnor U18043 (N_18043,N_17889,N_17768);
or U18044 (N_18044,N_17922,N_17753);
nor U18045 (N_18045,N_17984,N_17886);
nand U18046 (N_18046,N_17797,N_17918);
xnor U18047 (N_18047,N_17761,N_17796);
xnor U18048 (N_18048,N_17947,N_17808);
or U18049 (N_18049,N_17825,N_17892);
and U18050 (N_18050,N_17940,N_17923);
xor U18051 (N_18051,N_17765,N_17929);
or U18052 (N_18052,N_17847,N_17953);
nor U18053 (N_18053,N_17759,N_17893);
xor U18054 (N_18054,N_17767,N_17973);
or U18055 (N_18055,N_17815,N_17885);
or U18056 (N_18056,N_17855,N_17854);
nor U18057 (N_18057,N_17912,N_17795);
or U18058 (N_18058,N_17901,N_17891);
nand U18059 (N_18059,N_17888,N_17793);
nor U18060 (N_18060,N_17986,N_17908);
xnor U18061 (N_18061,N_17756,N_17974);
xor U18062 (N_18062,N_17830,N_17863);
xnor U18063 (N_18063,N_17883,N_17771);
or U18064 (N_18064,N_17846,N_17895);
and U18065 (N_18065,N_17776,N_17827);
nor U18066 (N_18066,N_17798,N_17821);
nor U18067 (N_18067,N_17928,N_17868);
and U18068 (N_18068,N_17772,N_17964);
or U18069 (N_18069,N_17779,N_17792);
nor U18070 (N_18070,N_17996,N_17807);
xor U18071 (N_18071,N_17770,N_17875);
nor U18072 (N_18072,N_17809,N_17754);
xnor U18073 (N_18073,N_17992,N_17955);
nand U18074 (N_18074,N_17959,N_17932);
nor U18075 (N_18075,N_17998,N_17806);
nor U18076 (N_18076,N_17900,N_17774);
xor U18077 (N_18077,N_17833,N_17946);
and U18078 (N_18078,N_17750,N_17780);
or U18079 (N_18079,N_17801,N_17831);
or U18080 (N_18080,N_17778,N_17762);
and U18081 (N_18081,N_17884,N_17871);
xnor U18082 (N_18082,N_17755,N_17978);
nand U18083 (N_18083,N_17865,N_17840);
nand U18084 (N_18084,N_17887,N_17786);
nand U18085 (N_18085,N_17936,N_17866);
nor U18086 (N_18086,N_17769,N_17881);
and U18087 (N_18087,N_17834,N_17823);
nor U18088 (N_18088,N_17933,N_17991);
or U18089 (N_18089,N_17781,N_17909);
and U18090 (N_18090,N_17828,N_17983);
and U18091 (N_18091,N_17810,N_17910);
or U18092 (N_18092,N_17890,N_17968);
or U18093 (N_18093,N_17874,N_17822);
xor U18094 (N_18094,N_17794,N_17989);
or U18095 (N_18095,N_17819,N_17937);
xor U18096 (N_18096,N_17850,N_17950);
or U18097 (N_18097,N_17907,N_17994);
nor U18098 (N_18098,N_17945,N_17924);
nand U18099 (N_18099,N_17981,N_17751);
xnor U18100 (N_18100,N_17913,N_17904);
nor U18101 (N_18101,N_17917,N_17843);
nor U18102 (N_18102,N_17752,N_17944);
nor U18103 (N_18103,N_17816,N_17814);
nand U18104 (N_18104,N_17862,N_17880);
nor U18105 (N_18105,N_17931,N_17870);
and U18106 (N_18106,N_17951,N_17882);
or U18107 (N_18107,N_17757,N_17954);
or U18108 (N_18108,N_17859,N_17760);
xor U18109 (N_18109,N_17990,N_17988);
nor U18110 (N_18110,N_17970,N_17805);
or U18111 (N_18111,N_17934,N_17788);
nor U18112 (N_18112,N_17902,N_17867);
nor U18113 (N_18113,N_17916,N_17921);
xnor U18114 (N_18114,N_17938,N_17849);
and U18115 (N_18115,N_17899,N_17777);
nand U18116 (N_18116,N_17948,N_17903);
or U18117 (N_18117,N_17764,N_17782);
or U18118 (N_18118,N_17841,N_17962);
nand U18119 (N_18119,N_17977,N_17914);
nor U18120 (N_18120,N_17872,N_17894);
nor U18121 (N_18121,N_17832,N_17785);
or U18122 (N_18122,N_17935,N_17911);
or U18123 (N_18123,N_17839,N_17853);
or U18124 (N_18124,N_17919,N_17842);
xor U18125 (N_18125,N_17810,N_17869);
xnor U18126 (N_18126,N_17974,N_17758);
xnor U18127 (N_18127,N_17787,N_17777);
nand U18128 (N_18128,N_17964,N_17947);
nand U18129 (N_18129,N_17997,N_17895);
and U18130 (N_18130,N_17867,N_17903);
nor U18131 (N_18131,N_17941,N_17952);
or U18132 (N_18132,N_17778,N_17933);
nor U18133 (N_18133,N_17864,N_17768);
or U18134 (N_18134,N_17830,N_17896);
xor U18135 (N_18135,N_17960,N_17859);
xor U18136 (N_18136,N_17959,N_17897);
nor U18137 (N_18137,N_17790,N_17792);
and U18138 (N_18138,N_17847,N_17758);
nor U18139 (N_18139,N_17905,N_17973);
or U18140 (N_18140,N_17836,N_17942);
and U18141 (N_18141,N_17899,N_17888);
or U18142 (N_18142,N_17952,N_17887);
nor U18143 (N_18143,N_17762,N_17960);
and U18144 (N_18144,N_17858,N_17897);
or U18145 (N_18145,N_17856,N_17865);
xor U18146 (N_18146,N_17971,N_17772);
xnor U18147 (N_18147,N_17962,N_17908);
nand U18148 (N_18148,N_17984,N_17859);
or U18149 (N_18149,N_17962,N_17827);
and U18150 (N_18150,N_17942,N_17987);
nor U18151 (N_18151,N_17782,N_17852);
nand U18152 (N_18152,N_17872,N_17948);
or U18153 (N_18153,N_17774,N_17913);
and U18154 (N_18154,N_17874,N_17900);
nand U18155 (N_18155,N_17948,N_17921);
or U18156 (N_18156,N_17970,N_17996);
nor U18157 (N_18157,N_17760,N_17814);
nand U18158 (N_18158,N_17875,N_17960);
and U18159 (N_18159,N_17762,N_17860);
nor U18160 (N_18160,N_17961,N_17822);
and U18161 (N_18161,N_17812,N_17912);
and U18162 (N_18162,N_17780,N_17783);
and U18163 (N_18163,N_17798,N_17850);
xor U18164 (N_18164,N_17903,N_17854);
nor U18165 (N_18165,N_17968,N_17829);
or U18166 (N_18166,N_17884,N_17947);
nand U18167 (N_18167,N_17841,N_17964);
nand U18168 (N_18168,N_17912,N_17889);
and U18169 (N_18169,N_17994,N_17865);
nor U18170 (N_18170,N_17968,N_17778);
nand U18171 (N_18171,N_17841,N_17900);
xnor U18172 (N_18172,N_17884,N_17815);
and U18173 (N_18173,N_17803,N_17875);
nand U18174 (N_18174,N_17809,N_17923);
xor U18175 (N_18175,N_17869,N_17897);
or U18176 (N_18176,N_17763,N_17765);
and U18177 (N_18177,N_17940,N_17821);
and U18178 (N_18178,N_17809,N_17964);
and U18179 (N_18179,N_17848,N_17883);
nor U18180 (N_18180,N_17816,N_17974);
nand U18181 (N_18181,N_17883,N_17761);
and U18182 (N_18182,N_17802,N_17821);
or U18183 (N_18183,N_17844,N_17962);
xnor U18184 (N_18184,N_17887,N_17918);
xnor U18185 (N_18185,N_17832,N_17912);
and U18186 (N_18186,N_17874,N_17906);
nor U18187 (N_18187,N_17913,N_17973);
nor U18188 (N_18188,N_17873,N_17884);
and U18189 (N_18189,N_17778,N_17777);
and U18190 (N_18190,N_17927,N_17921);
xnor U18191 (N_18191,N_17905,N_17867);
or U18192 (N_18192,N_17758,N_17969);
nand U18193 (N_18193,N_17780,N_17901);
or U18194 (N_18194,N_17835,N_17947);
nor U18195 (N_18195,N_17976,N_17848);
and U18196 (N_18196,N_17899,N_17750);
nand U18197 (N_18197,N_17788,N_17789);
nor U18198 (N_18198,N_17844,N_17960);
and U18199 (N_18199,N_17850,N_17938);
nand U18200 (N_18200,N_17807,N_17775);
or U18201 (N_18201,N_17948,N_17762);
nand U18202 (N_18202,N_17790,N_17973);
or U18203 (N_18203,N_17869,N_17851);
nor U18204 (N_18204,N_17982,N_17792);
or U18205 (N_18205,N_17934,N_17812);
or U18206 (N_18206,N_17902,N_17815);
xor U18207 (N_18207,N_17865,N_17940);
and U18208 (N_18208,N_17926,N_17808);
or U18209 (N_18209,N_17870,N_17864);
nand U18210 (N_18210,N_17873,N_17975);
nand U18211 (N_18211,N_17818,N_17863);
nand U18212 (N_18212,N_17804,N_17951);
nand U18213 (N_18213,N_17896,N_17829);
or U18214 (N_18214,N_17942,N_17920);
xor U18215 (N_18215,N_17793,N_17776);
or U18216 (N_18216,N_17843,N_17964);
or U18217 (N_18217,N_17895,N_17905);
and U18218 (N_18218,N_17811,N_17785);
nor U18219 (N_18219,N_17782,N_17886);
or U18220 (N_18220,N_17939,N_17842);
nand U18221 (N_18221,N_17899,N_17844);
and U18222 (N_18222,N_17859,N_17866);
xnor U18223 (N_18223,N_17913,N_17896);
nand U18224 (N_18224,N_17780,N_17804);
or U18225 (N_18225,N_17992,N_17803);
nand U18226 (N_18226,N_17964,N_17803);
or U18227 (N_18227,N_17841,N_17820);
or U18228 (N_18228,N_17965,N_17942);
or U18229 (N_18229,N_17755,N_17758);
nand U18230 (N_18230,N_17809,N_17980);
xnor U18231 (N_18231,N_17817,N_17845);
and U18232 (N_18232,N_17860,N_17843);
nor U18233 (N_18233,N_17878,N_17960);
or U18234 (N_18234,N_17898,N_17917);
or U18235 (N_18235,N_17887,N_17873);
nor U18236 (N_18236,N_17981,N_17994);
xnor U18237 (N_18237,N_17924,N_17775);
or U18238 (N_18238,N_17940,N_17820);
nor U18239 (N_18239,N_17750,N_17910);
nand U18240 (N_18240,N_17777,N_17792);
nor U18241 (N_18241,N_17891,N_17809);
and U18242 (N_18242,N_17813,N_17859);
or U18243 (N_18243,N_17777,N_17806);
nand U18244 (N_18244,N_17971,N_17958);
or U18245 (N_18245,N_17856,N_17849);
nand U18246 (N_18246,N_17971,N_17939);
nor U18247 (N_18247,N_17883,N_17887);
xor U18248 (N_18248,N_17827,N_17983);
or U18249 (N_18249,N_17913,N_17863);
nand U18250 (N_18250,N_18203,N_18076);
or U18251 (N_18251,N_18081,N_18113);
nor U18252 (N_18252,N_18012,N_18135);
or U18253 (N_18253,N_18187,N_18048);
and U18254 (N_18254,N_18136,N_18202);
nand U18255 (N_18255,N_18063,N_18009);
and U18256 (N_18256,N_18032,N_18055);
xor U18257 (N_18257,N_18053,N_18003);
xnor U18258 (N_18258,N_18071,N_18069);
and U18259 (N_18259,N_18041,N_18130);
and U18260 (N_18260,N_18115,N_18178);
nand U18261 (N_18261,N_18153,N_18169);
nand U18262 (N_18262,N_18129,N_18212);
xor U18263 (N_18263,N_18161,N_18198);
nor U18264 (N_18264,N_18028,N_18025);
nand U18265 (N_18265,N_18029,N_18031);
and U18266 (N_18266,N_18083,N_18089);
nor U18267 (N_18267,N_18010,N_18228);
and U18268 (N_18268,N_18194,N_18121);
nor U18269 (N_18269,N_18145,N_18229);
xnor U18270 (N_18270,N_18247,N_18208);
nor U18271 (N_18271,N_18157,N_18188);
xor U18272 (N_18272,N_18051,N_18195);
xnor U18273 (N_18273,N_18215,N_18039);
and U18274 (N_18274,N_18019,N_18190);
or U18275 (N_18275,N_18101,N_18227);
or U18276 (N_18276,N_18112,N_18013);
or U18277 (N_18277,N_18074,N_18026);
and U18278 (N_18278,N_18137,N_18217);
xor U18279 (N_18279,N_18235,N_18084);
xnor U18280 (N_18280,N_18104,N_18164);
xnor U18281 (N_18281,N_18058,N_18148);
nand U18282 (N_18282,N_18160,N_18245);
nand U18283 (N_18283,N_18175,N_18100);
xor U18284 (N_18284,N_18172,N_18065);
and U18285 (N_18285,N_18177,N_18170);
xor U18286 (N_18286,N_18117,N_18222);
or U18287 (N_18287,N_18124,N_18186);
xor U18288 (N_18288,N_18033,N_18205);
nor U18289 (N_18289,N_18183,N_18180);
nand U18290 (N_18290,N_18165,N_18006);
and U18291 (N_18291,N_18036,N_18139);
or U18292 (N_18292,N_18020,N_18173);
xnor U18293 (N_18293,N_18191,N_18151);
and U18294 (N_18294,N_18163,N_18231);
xnor U18295 (N_18295,N_18192,N_18144);
nor U18296 (N_18296,N_18141,N_18056);
xor U18297 (N_18297,N_18125,N_18244);
nor U18298 (N_18298,N_18097,N_18209);
or U18299 (N_18299,N_18226,N_18054);
and U18300 (N_18300,N_18064,N_18199);
and U18301 (N_18301,N_18092,N_18220);
xor U18302 (N_18302,N_18037,N_18072);
or U18303 (N_18303,N_18118,N_18107);
nor U18304 (N_18304,N_18015,N_18088);
nand U18305 (N_18305,N_18002,N_18146);
xor U18306 (N_18306,N_18241,N_18134);
or U18307 (N_18307,N_18082,N_18147);
nand U18308 (N_18308,N_18138,N_18011);
and U18309 (N_18309,N_18197,N_18080);
nor U18310 (N_18310,N_18196,N_18149);
and U18311 (N_18311,N_18167,N_18142);
or U18312 (N_18312,N_18004,N_18182);
nor U18313 (N_18313,N_18030,N_18090);
nand U18314 (N_18314,N_18200,N_18211);
nor U18315 (N_18315,N_18075,N_18027);
and U18316 (N_18316,N_18116,N_18106);
or U18317 (N_18317,N_18174,N_18181);
or U18318 (N_18318,N_18213,N_18238);
xnor U18319 (N_18319,N_18152,N_18050);
or U18320 (N_18320,N_18007,N_18111);
nand U18321 (N_18321,N_18207,N_18038);
nor U18322 (N_18322,N_18091,N_18109);
or U18323 (N_18323,N_18201,N_18043);
or U18324 (N_18324,N_18224,N_18021);
and U18325 (N_18325,N_18000,N_18034);
nand U18326 (N_18326,N_18094,N_18171);
nand U18327 (N_18327,N_18189,N_18119);
xor U18328 (N_18328,N_18070,N_18060);
nor U18329 (N_18329,N_18122,N_18061);
nor U18330 (N_18330,N_18123,N_18114);
and U18331 (N_18331,N_18042,N_18204);
nand U18332 (N_18332,N_18035,N_18248);
and U18333 (N_18333,N_18214,N_18022);
nor U18334 (N_18334,N_18246,N_18024);
nand U18335 (N_18335,N_18128,N_18073);
nand U18336 (N_18336,N_18168,N_18166);
nand U18337 (N_18337,N_18102,N_18062);
and U18338 (N_18338,N_18159,N_18132);
xor U18339 (N_18339,N_18017,N_18018);
xor U18340 (N_18340,N_18023,N_18140);
and U18341 (N_18341,N_18242,N_18044);
or U18342 (N_18342,N_18087,N_18085);
nor U18343 (N_18343,N_18049,N_18120);
xor U18344 (N_18344,N_18218,N_18059);
or U18345 (N_18345,N_18110,N_18077);
or U18346 (N_18346,N_18068,N_18185);
nor U18347 (N_18347,N_18236,N_18105);
xnor U18348 (N_18348,N_18206,N_18216);
xnor U18349 (N_18349,N_18093,N_18233);
nor U18350 (N_18350,N_18210,N_18066);
or U18351 (N_18351,N_18096,N_18086);
and U18352 (N_18352,N_18158,N_18095);
and U18353 (N_18353,N_18040,N_18179);
nand U18354 (N_18354,N_18249,N_18219);
nor U18355 (N_18355,N_18223,N_18127);
nand U18356 (N_18356,N_18057,N_18232);
nor U18357 (N_18357,N_18240,N_18131);
and U18358 (N_18358,N_18150,N_18239);
or U18359 (N_18359,N_18243,N_18067);
or U18360 (N_18360,N_18098,N_18079);
xnor U18361 (N_18361,N_18103,N_18126);
or U18362 (N_18362,N_18225,N_18193);
nor U18363 (N_18363,N_18099,N_18001);
xor U18364 (N_18364,N_18234,N_18221);
and U18365 (N_18365,N_18155,N_18143);
nor U18366 (N_18366,N_18045,N_18230);
nand U18367 (N_18367,N_18046,N_18008);
nand U18368 (N_18368,N_18014,N_18237);
xor U18369 (N_18369,N_18176,N_18047);
nand U18370 (N_18370,N_18156,N_18133);
or U18371 (N_18371,N_18005,N_18108);
and U18372 (N_18372,N_18078,N_18016);
or U18373 (N_18373,N_18052,N_18162);
xor U18374 (N_18374,N_18154,N_18184);
and U18375 (N_18375,N_18088,N_18150);
and U18376 (N_18376,N_18089,N_18168);
nor U18377 (N_18377,N_18122,N_18088);
xor U18378 (N_18378,N_18113,N_18161);
nand U18379 (N_18379,N_18220,N_18146);
and U18380 (N_18380,N_18097,N_18084);
nand U18381 (N_18381,N_18094,N_18147);
xnor U18382 (N_18382,N_18209,N_18104);
nor U18383 (N_18383,N_18064,N_18119);
and U18384 (N_18384,N_18104,N_18062);
or U18385 (N_18385,N_18033,N_18152);
and U18386 (N_18386,N_18137,N_18239);
nand U18387 (N_18387,N_18152,N_18189);
or U18388 (N_18388,N_18094,N_18200);
and U18389 (N_18389,N_18026,N_18050);
and U18390 (N_18390,N_18210,N_18120);
and U18391 (N_18391,N_18109,N_18217);
nor U18392 (N_18392,N_18035,N_18042);
xnor U18393 (N_18393,N_18065,N_18085);
and U18394 (N_18394,N_18245,N_18191);
or U18395 (N_18395,N_18197,N_18215);
nor U18396 (N_18396,N_18201,N_18129);
nand U18397 (N_18397,N_18225,N_18177);
nor U18398 (N_18398,N_18227,N_18000);
and U18399 (N_18399,N_18066,N_18079);
and U18400 (N_18400,N_18023,N_18151);
or U18401 (N_18401,N_18158,N_18143);
or U18402 (N_18402,N_18246,N_18036);
nor U18403 (N_18403,N_18158,N_18224);
nand U18404 (N_18404,N_18100,N_18132);
xnor U18405 (N_18405,N_18086,N_18126);
or U18406 (N_18406,N_18179,N_18234);
nor U18407 (N_18407,N_18046,N_18105);
nand U18408 (N_18408,N_18045,N_18156);
xnor U18409 (N_18409,N_18128,N_18150);
nand U18410 (N_18410,N_18195,N_18233);
or U18411 (N_18411,N_18139,N_18146);
xor U18412 (N_18412,N_18052,N_18118);
nand U18413 (N_18413,N_18184,N_18085);
nor U18414 (N_18414,N_18202,N_18196);
nor U18415 (N_18415,N_18147,N_18056);
nand U18416 (N_18416,N_18082,N_18024);
xnor U18417 (N_18417,N_18132,N_18062);
nand U18418 (N_18418,N_18170,N_18060);
nor U18419 (N_18419,N_18148,N_18159);
or U18420 (N_18420,N_18089,N_18195);
xor U18421 (N_18421,N_18134,N_18102);
or U18422 (N_18422,N_18058,N_18214);
xnor U18423 (N_18423,N_18150,N_18072);
or U18424 (N_18424,N_18031,N_18183);
nor U18425 (N_18425,N_18229,N_18144);
nor U18426 (N_18426,N_18180,N_18042);
and U18427 (N_18427,N_18073,N_18239);
nand U18428 (N_18428,N_18117,N_18028);
and U18429 (N_18429,N_18087,N_18122);
nor U18430 (N_18430,N_18164,N_18076);
nand U18431 (N_18431,N_18114,N_18044);
xor U18432 (N_18432,N_18171,N_18179);
nor U18433 (N_18433,N_18199,N_18070);
nor U18434 (N_18434,N_18144,N_18000);
xor U18435 (N_18435,N_18056,N_18020);
nand U18436 (N_18436,N_18161,N_18028);
or U18437 (N_18437,N_18197,N_18213);
or U18438 (N_18438,N_18145,N_18160);
and U18439 (N_18439,N_18123,N_18089);
or U18440 (N_18440,N_18096,N_18087);
xor U18441 (N_18441,N_18118,N_18108);
nand U18442 (N_18442,N_18056,N_18163);
nor U18443 (N_18443,N_18109,N_18088);
xor U18444 (N_18444,N_18024,N_18191);
nand U18445 (N_18445,N_18222,N_18044);
or U18446 (N_18446,N_18143,N_18025);
nor U18447 (N_18447,N_18046,N_18050);
xor U18448 (N_18448,N_18041,N_18126);
xor U18449 (N_18449,N_18087,N_18040);
and U18450 (N_18450,N_18231,N_18142);
and U18451 (N_18451,N_18027,N_18157);
and U18452 (N_18452,N_18245,N_18100);
or U18453 (N_18453,N_18162,N_18087);
xnor U18454 (N_18454,N_18219,N_18241);
nand U18455 (N_18455,N_18216,N_18029);
and U18456 (N_18456,N_18214,N_18134);
and U18457 (N_18457,N_18077,N_18102);
nor U18458 (N_18458,N_18066,N_18121);
nor U18459 (N_18459,N_18014,N_18073);
and U18460 (N_18460,N_18241,N_18103);
nand U18461 (N_18461,N_18176,N_18064);
or U18462 (N_18462,N_18051,N_18102);
nand U18463 (N_18463,N_18237,N_18050);
and U18464 (N_18464,N_18131,N_18194);
xnor U18465 (N_18465,N_18070,N_18010);
xnor U18466 (N_18466,N_18025,N_18024);
xnor U18467 (N_18467,N_18096,N_18154);
xor U18468 (N_18468,N_18030,N_18244);
and U18469 (N_18469,N_18009,N_18114);
nor U18470 (N_18470,N_18158,N_18098);
nand U18471 (N_18471,N_18162,N_18204);
and U18472 (N_18472,N_18249,N_18208);
xor U18473 (N_18473,N_18242,N_18156);
nor U18474 (N_18474,N_18132,N_18239);
and U18475 (N_18475,N_18217,N_18090);
or U18476 (N_18476,N_18210,N_18087);
nand U18477 (N_18477,N_18228,N_18208);
and U18478 (N_18478,N_18167,N_18233);
nand U18479 (N_18479,N_18020,N_18210);
nand U18480 (N_18480,N_18054,N_18006);
or U18481 (N_18481,N_18098,N_18244);
and U18482 (N_18482,N_18057,N_18213);
and U18483 (N_18483,N_18131,N_18005);
or U18484 (N_18484,N_18076,N_18165);
xor U18485 (N_18485,N_18030,N_18066);
or U18486 (N_18486,N_18027,N_18235);
nor U18487 (N_18487,N_18004,N_18185);
and U18488 (N_18488,N_18190,N_18057);
and U18489 (N_18489,N_18225,N_18056);
xnor U18490 (N_18490,N_18003,N_18006);
and U18491 (N_18491,N_18084,N_18030);
xnor U18492 (N_18492,N_18018,N_18116);
and U18493 (N_18493,N_18218,N_18167);
or U18494 (N_18494,N_18225,N_18065);
or U18495 (N_18495,N_18018,N_18113);
or U18496 (N_18496,N_18176,N_18182);
or U18497 (N_18497,N_18186,N_18216);
xor U18498 (N_18498,N_18138,N_18004);
nor U18499 (N_18499,N_18219,N_18019);
or U18500 (N_18500,N_18300,N_18325);
xnor U18501 (N_18501,N_18305,N_18382);
xnor U18502 (N_18502,N_18493,N_18274);
xor U18503 (N_18503,N_18397,N_18479);
xor U18504 (N_18504,N_18335,N_18282);
and U18505 (N_18505,N_18441,N_18426);
xnor U18506 (N_18506,N_18256,N_18400);
and U18507 (N_18507,N_18492,N_18278);
xor U18508 (N_18508,N_18427,N_18338);
nor U18509 (N_18509,N_18250,N_18329);
nor U18510 (N_18510,N_18414,N_18353);
or U18511 (N_18511,N_18462,N_18350);
nor U18512 (N_18512,N_18408,N_18401);
nand U18513 (N_18513,N_18299,N_18330);
or U18514 (N_18514,N_18362,N_18336);
nand U18515 (N_18515,N_18355,N_18496);
or U18516 (N_18516,N_18402,N_18322);
and U18517 (N_18517,N_18410,N_18298);
xnor U18518 (N_18518,N_18475,N_18381);
nand U18519 (N_18519,N_18385,N_18473);
xor U18520 (N_18520,N_18415,N_18477);
xor U18521 (N_18521,N_18392,N_18471);
nand U18522 (N_18522,N_18294,N_18277);
nand U18523 (N_18523,N_18483,N_18442);
xor U18524 (N_18524,N_18478,N_18316);
nand U18525 (N_18525,N_18379,N_18433);
xor U18526 (N_18526,N_18340,N_18461);
and U18527 (N_18527,N_18369,N_18268);
xor U18528 (N_18528,N_18312,N_18365);
nand U18529 (N_18529,N_18318,N_18404);
nor U18530 (N_18530,N_18388,N_18279);
and U18531 (N_18531,N_18418,N_18284);
or U18532 (N_18532,N_18344,N_18320);
xor U18533 (N_18533,N_18425,N_18302);
xnor U18534 (N_18534,N_18292,N_18422);
nand U18535 (N_18535,N_18361,N_18390);
xnor U18536 (N_18536,N_18447,N_18384);
and U18537 (N_18537,N_18494,N_18259);
and U18538 (N_18538,N_18341,N_18393);
or U18539 (N_18539,N_18399,N_18421);
and U18540 (N_18540,N_18303,N_18458);
or U18541 (N_18541,N_18254,N_18417);
and U18542 (N_18542,N_18286,N_18367);
nor U18543 (N_18543,N_18326,N_18464);
nor U18544 (N_18544,N_18260,N_18395);
nor U18545 (N_18545,N_18272,N_18283);
nand U18546 (N_18546,N_18373,N_18364);
nor U18547 (N_18547,N_18405,N_18285);
xor U18548 (N_18548,N_18389,N_18308);
xnor U18549 (N_18549,N_18333,N_18280);
or U18550 (N_18550,N_18486,N_18370);
nand U18551 (N_18551,N_18430,N_18310);
and U18552 (N_18552,N_18440,N_18267);
xnor U18553 (N_18553,N_18484,N_18453);
nor U18554 (N_18554,N_18295,N_18387);
and U18555 (N_18555,N_18323,N_18474);
nor U18556 (N_18556,N_18363,N_18269);
or U18557 (N_18557,N_18380,N_18375);
xor U18558 (N_18558,N_18297,N_18352);
nor U18559 (N_18559,N_18281,N_18411);
nor U18560 (N_18560,N_18357,N_18327);
or U18561 (N_18561,N_18301,N_18495);
xnor U18562 (N_18562,N_18446,N_18354);
or U18563 (N_18563,N_18424,N_18386);
nand U18564 (N_18564,N_18319,N_18324);
and U18565 (N_18565,N_18288,N_18413);
or U18566 (N_18566,N_18266,N_18450);
nor U18567 (N_18567,N_18472,N_18378);
xnor U18568 (N_18568,N_18346,N_18251);
nor U18569 (N_18569,N_18255,N_18291);
and U18570 (N_18570,N_18456,N_18276);
xnor U18571 (N_18571,N_18459,N_18331);
nand U18572 (N_18572,N_18454,N_18314);
xor U18573 (N_18573,N_18396,N_18358);
or U18574 (N_18574,N_18432,N_18339);
nor U18575 (N_18575,N_18485,N_18449);
nor U18576 (N_18576,N_18368,N_18443);
nand U18577 (N_18577,N_18383,N_18293);
nand U18578 (N_18578,N_18349,N_18487);
nand U18579 (N_18579,N_18287,N_18342);
nand U18580 (N_18580,N_18271,N_18306);
and U18581 (N_18581,N_18435,N_18460);
nor U18582 (N_18582,N_18304,N_18311);
and U18583 (N_18583,N_18315,N_18409);
xor U18584 (N_18584,N_18498,N_18348);
nor U18585 (N_18585,N_18332,N_18445);
xor U18586 (N_18586,N_18434,N_18253);
and U18587 (N_18587,N_18273,N_18491);
and U18588 (N_18588,N_18419,N_18366);
or U18589 (N_18589,N_18457,N_18423);
nand U18590 (N_18590,N_18465,N_18347);
nor U18591 (N_18591,N_18489,N_18372);
or U18592 (N_18592,N_18391,N_18431);
and U18593 (N_18593,N_18394,N_18406);
or U18594 (N_18594,N_18416,N_18466);
or U18595 (N_18595,N_18463,N_18420);
xnor U18596 (N_18596,N_18448,N_18499);
nor U18597 (N_18597,N_18436,N_18261);
and U18598 (N_18598,N_18313,N_18481);
and U18599 (N_18599,N_18263,N_18343);
and U18600 (N_18600,N_18469,N_18345);
and U18601 (N_18601,N_18290,N_18403);
or U18602 (N_18602,N_18451,N_18429);
or U18603 (N_18603,N_18467,N_18480);
and U18604 (N_18604,N_18328,N_18359);
and U18605 (N_18605,N_18265,N_18490);
or U18606 (N_18606,N_18437,N_18275);
nor U18607 (N_18607,N_18371,N_18289);
nor U18608 (N_18608,N_18296,N_18252);
nand U18609 (N_18609,N_18262,N_18351);
and U18610 (N_18610,N_18376,N_18488);
nand U18611 (N_18611,N_18377,N_18309);
xor U18612 (N_18612,N_18444,N_18470);
and U18613 (N_18613,N_18476,N_18428);
nor U18614 (N_18614,N_18412,N_18334);
xnor U18615 (N_18615,N_18257,N_18337);
or U18616 (N_18616,N_18398,N_18407);
nor U18617 (N_18617,N_18438,N_18455);
and U18618 (N_18618,N_18356,N_18482);
and U18619 (N_18619,N_18258,N_18360);
xor U18620 (N_18620,N_18439,N_18264);
nor U18621 (N_18621,N_18321,N_18317);
nand U18622 (N_18622,N_18497,N_18374);
nor U18623 (N_18623,N_18468,N_18452);
and U18624 (N_18624,N_18307,N_18270);
or U18625 (N_18625,N_18297,N_18404);
and U18626 (N_18626,N_18337,N_18335);
nor U18627 (N_18627,N_18324,N_18333);
and U18628 (N_18628,N_18357,N_18273);
xor U18629 (N_18629,N_18353,N_18422);
nand U18630 (N_18630,N_18367,N_18361);
or U18631 (N_18631,N_18267,N_18449);
nand U18632 (N_18632,N_18476,N_18467);
nor U18633 (N_18633,N_18480,N_18487);
nor U18634 (N_18634,N_18355,N_18461);
or U18635 (N_18635,N_18393,N_18456);
nor U18636 (N_18636,N_18313,N_18488);
xnor U18637 (N_18637,N_18310,N_18428);
xor U18638 (N_18638,N_18290,N_18441);
nand U18639 (N_18639,N_18460,N_18413);
nand U18640 (N_18640,N_18312,N_18313);
xor U18641 (N_18641,N_18418,N_18307);
xnor U18642 (N_18642,N_18306,N_18314);
nand U18643 (N_18643,N_18423,N_18309);
nand U18644 (N_18644,N_18424,N_18266);
nor U18645 (N_18645,N_18291,N_18462);
and U18646 (N_18646,N_18260,N_18317);
and U18647 (N_18647,N_18486,N_18270);
nand U18648 (N_18648,N_18470,N_18311);
and U18649 (N_18649,N_18294,N_18314);
nor U18650 (N_18650,N_18428,N_18480);
or U18651 (N_18651,N_18263,N_18339);
and U18652 (N_18652,N_18321,N_18485);
xor U18653 (N_18653,N_18311,N_18270);
xnor U18654 (N_18654,N_18402,N_18431);
or U18655 (N_18655,N_18430,N_18323);
nor U18656 (N_18656,N_18325,N_18369);
and U18657 (N_18657,N_18388,N_18492);
nor U18658 (N_18658,N_18376,N_18335);
or U18659 (N_18659,N_18326,N_18460);
or U18660 (N_18660,N_18301,N_18298);
xnor U18661 (N_18661,N_18468,N_18410);
or U18662 (N_18662,N_18359,N_18260);
nor U18663 (N_18663,N_18341,N_18285);
xor U18664 (N_18664,N_18482,N_18328);
or U18665 (N_18665,N_18350,N_18490);
nor U18666 (N_18666,N_18336,N_18327);
or U18667 (N_18667,N_18325,N_18258);
nand U18668 (N_18668,N_18467,N_18252);
nor U18669 (N_18669,N_18275,N_18451);
nand U18670 (N_18670,N_18309,N_18254);
nand U18671 (N_18671,N_18306,N_18386);
xor U18672 (N_18672,N_18388,N_18332);
nand U18673 (N_18673,N_18300,N_18288);
or U18674 (N_18674,N_18498,N_18408);
xnor U18675 (N_18675,N_18438,N_18273);
or U18676 (N_18676,N_18373,N_18492);
and U18677 (N_18677,N_18465,N_18424);
or U18678 (N_18678,N_18283,N_18469);
nor U18679 (N_18679,N_18403,N_18348);
nand U18680 (N_18680,N_18275,N_18467);
and U18681 (N_18681,N_18352,N_18288);
or U18682 (N_18682,N_18471,N_18404);
and U18683 (N_18683,N_18314,N_18435);
xor U18684 (N_18684,N_18457,N_18372);
xnor U18685 (N_18685,N_18449,N_18386);
nor U18686 (N_18686,N_18296,N_18386);
nand U18687 (N_18687,N_18302,N_18402);
xnor U18688 (N_18688,N_18306,N_18257);
xor U18689 (N_18689,N_18477,N_18487);
nand U18690 (N_18690,N_18251,N_18322);
or U18691 (N_18691,N_18330,N_18332);
nand U18692 (N_18692,N_18363,N_18496);
and U18693 (N_18693,N_18390,N_18300);
nand U18694 (N_18694,N_18401,N_18404);
xnor U18695 (N_18695,N_18355,N_18415);
or U18696 (N_18696,N_18258,N_18394);
or U18697 (N_18697,N_18419,N_18306);
nor U18698 (N_18698,N_18499,N_18323);
nor U18699 (N_18699,N_18447,N_18354);
xor U18700 (N_18700,N_18416,N_18336);
or U18701 (N_18701,N_18379,N_18252);
nand U18702 (N_18702,N_18324,N_18426);
or U18703 (N_18703,N_18266,N_18494);
or U18704 (N_18704,N_18382,N_18494);
nand U18705 (N_18705,N_18250,N_18418);
and U18706 (N_18706,N_18471,N_18490);
or U18707 (N_18707,N_18408,N_18375);
nor U18708 (N_18708,N_18399,N_18496);
nand U18709 (N_18709,N_18495,N_18258);
nand U18710 (N_18710,N_18256,N_18480);
nor U18711 (N_18711,N_18362,N_18323);
xor U18712 (N_18712,N_18390,N_18477);
and U18713 (N_18713,N_18270,N_18313);
xnor U18714 (N_18714,N_18473,N_18465);
nand U18715 (N_18715,N_18275,N_18458);
nor U18716 (N_18716,N_18419,N_18269);
nand U18717 (N_18717,N_18495,N_18413);
or U18718 (N_18718,N_18347,N_18433);
nand U18719 (N_18719,N_18308,N_18445);
and U18720 (N_18720,N_18350,N_18423);
and U18721 (N_18721,N_18277,N_18477);
or U18722 (N_18722,N_18293,N_18399);
nand U18723 (N_18723,N_18326,N_18257);
xnor U18724 (N_18724,N_18397,N_18438);
or U18725 (N_18725,N_18461,N_18396);
nor U18726 (N_18726,N_18467,N_18388);
and U18727 (N_18727,N_18347,N_18317);
or U18728 (N_18728,N_18371,N_18417);
and U18729 (N_18729,N_18419,N_18456);
or U18730 (N_18730,N_18337,N_18322);
and U18731 (N_18731,N_18348,N_18481);
nand U18732 (N_18732,N_18336,N_18283);
and U18733 (N_18733,N_18476,N_18439);
xnor U18734 (N_18734,N_18255,N_18476);
and U18735 (N_18735,N_18449,N_18392);
or U18736 (N_18736,N_18444,N_18394);
nand U18737 (N_18737,N_18346,N_18287);
or U18738 (N_18738,N_18496,N_18386);
xnor U18739 (N_18739,N_18436,N_18277);
nor U18740 (N_18740,N_18388,N_18432);
nor U18741 (N_18741,N_18332,N_18328);
xnor U18742 (N_18742,N_18250,N_18309);
nand U18743 (N_18743,N_18352,N_18395);
nor U18744 (N_18744,N_18298,N_18494);
xnor U18745 (N_18745,N_18302,N_18471);
and U18746 (N_18746,N_18267,N_18429);
or U18747 (N_18747,N_18489,N_18304);
nor U18748 (N_18748,N_18272,N_18487);
nand U18749 (N_18749,N_18268,N_18265);
nand U18750 (N_18750,N_18557,N_18575);
xor U18751 (N_18751,N_18747,N_18717);
and U18752 (N_18752,N_18704,N_18697);
nand U18753 (N_18753,N_18698,N_18655);
nand U18754 (N_18754,N_18519,N_18706);
xnor U18755 (N_18755,N_18541,N_18691);
nor U18756 (N_18756,N_18547,N_18682);
xnor U18757 (N_18757,N_18621,N_18740);
and U18758 (N_18758,N_18700,N_18588);
or U18759 (N_18759,N_18560,N_18596);
and U18760 (N_18760,N_18561,N_18531);
nand U18761 (N_18761,N_18600,N_18720);
xor U18762 (N_18762,N_18503,N_18637);
nand U18763 (N_18763,N_18705,N_18727);
or U18764 (N_18764,N_18578,N_18728);
nor U18765 (N_18765,N_18568,N_18688);
and U18766 (N_18766,N_18741,N_18726);
or U18767 (N_18767,N_18549,N_18734);
nand U18768 (N_18768,N_18701,N_18582);
or U18769 (N_18769,N_18696,N_18533);
and U18770 (N_18770,N_18501,N_18627);
and U18771 (N_18771,N_18689,N_18632);
or U18772 (N_18772,N_18508,N_18711);
nand U18773 (N_18773,N_18748,N_18517);
nor U18774 (N_18774,N_18725,N_18749);
nand U18775 (N_18775,N_18585,N_18673);
nand U18776 (N_18776,N_18580,N_18710);
nand U18777 (N_18777,N_18545,N_18719);
nor U18778 (N_18778,N_18555,N_18647);
nor U18779 (N_18779,N_18603,N_18666);
nor U18780 (N_18780,N_18644,N_18683);
nor U18781 (N_18781,N_18724,N_18633);
nand U18782 (N_18782,N_18524,N_18614);
nand U18783 (N_18783,N_18605,N_18690);
nand U18784 (N_18784,N_18664,N_18733);
nand U18785 (N_18785,N_18675,N_18654);
xor U18786 (N_18786,N_18743,N_18732);
and U18787 (N_18787,N_18671,N_18658);
nor U18788 (N_18788,N_18572,N_18616);
or U18789 (N_18789,N_18723,N_18514);
or U18790 (N_18790,N_18507,N_18611);
and U18791 (N_18791,N_18525,N_18737);
xor U18792 (N_18792,N_18712,N_18528);
nand U18793 (N_18793,N_18601,N_18665);
nand U18794 (N_18794,N_18657,N_18692);
nor U18795 (N_18795,N_18722,N_18641);
or U18796 (N_18796,N_18521,N_18598);
nor U18797 (N_18797,N_18635,N_18684);
or U18798 (N_18798,N_18573,N_18694);
nand U18799 (N_18799,N_18579,N_18680);
nor U18800 (N_18800,N_18583,N_18615);
nand U18801 (N_18801,N_18504,N_18718);
xor U18802 (N_18802,N_18703,N_18739);
xnor U18803 (N_18803,N_18593,N_18677);
or U18804 (N_18804,N_18590,N_18708);
or U18805 (N_18805,N_18623,N_18569);
nand U18806 (N_18806,N_18513,N_18625);
xor U18807 (N_18807,N_18642,N_18558);
nand U18808 (N_18808,N_18631,N_18713);
nand U18809 (N_18809,N_18653,N_18685);
and U18810 (N_18810,N_18742,N_18744);
nor U18811 (N_18811,N_18537,N_18552);
or U18812 (N_18812,N_18538,N_18544);
and U18813 (N_18813,N_18570,N_18628);
or U18814 (N_18814,N_18648,N_18526);
and U18815 (N_18815,N_18546,N_18535);
nor U18816 (N_18816,N_18556,N_18707);
or U18817 (N_18817,N_18512,N_18656);
or U18818 (N_18818,N_18746,N_18500);
nand U18819 (N_18819,N_18553,N_18550);
nand U18820 (N_18820,N_18670,N_18702);
and U18821 (N_18821,N_18509,N_18506);
nor U18822 (N_18822,N_18629,N_18624);
nand U18823 (N_18823,N_18518,N_18599);
nand U18824 (N_18824,N_18693,N_18716);
nor U18825 (N_18825,N_18731,N_18559);
nand U18826 (N_18826,N_18645,N_18604);
or U18827 (N_18827,N_18577,N_18571);
and U18828 (N_18828,N_18714,N_18662);
xor U18829 (N_18829,N_18626,N_18668);
and U18830 (N_18830,N_18609,N_18709);
nand U18831 (N_18831,N_18715,N_18638);
or U18832 (N_18832,N_18567,N_18607);
nand U18833 (N_18833,N_18516,N_18610);
xor U18834 (N_18834,N_18563,N_18745);
nor U18835 (N_18835,N_18566,N_18548);
nor U18836 (N_18836,N_18672,N_18618);
xor U18837 (N_18837,N_18539,N_18646);
and U18838 (N_18838,N_18591,N_18620);
and U18839 (N_18839,N_18622,N_18659);
nor U18840 (N_18840,N_18640,N_18699);
xor U18841 (N_18841,N_18669,N_18520);
nor U18842 (N_18842,N_18534,N_18619);
nand U18843 (N_18843,N_18606,N_18510);
nor U18844 (N_18844,N_18595,N_18721);
nand U18845 (N_18845,N_18735,N_18634);
nor U18846 (N_18846,N_18674,N_18676);
and U18847 (N_18847,N_18586,N_18527);
or U18848 (N_18848,N_18502,N_18738);
and U18849 (N_18849,N_18695,N_18511);
and U18850 (N_18850,N_18581,N_18551);
nand U18851 (N_18851,N_18663,N_18636);
or U18852 (N_18852,N_18532,N_18729);
and U18853 (N_18853,N_18542,N_18523);
nor U18854 (N_18854,N_18613,N_18529);
and U18855 (N_18855,N_18540,N_18576);
nor U18856 (N_18856,N_18736,N_18564);
xnor U18857 (N_18857,N_18602,N_18687);
nand U18858 (N_18858,N_18565,N_18617);
nand U18859 (N_18859,N_18651,N_18587);
or U18860 (N_18860,N_18730,N_18589);
nor U18861 (N_18861,N_18543,N_18686);
or U18862 (N_18862,N_18630,N_18660);
or U18863 (N_18863,N_18679,N_18649);
or U18864 (N_18864,N_18678,N_18612);
or U18865 (N_18865,N_18650,N_18652);
or U18866 (N_18866,N_18608,N_18522);
nor U18867 (N_18867,N_18592,N_18574);
or U18868 (N_18868,N_18681,N_18584);
and U18869 (N_18869,N_18643,N_18530);
nor U18870 (N_18870,N_18536,N_18597);
or U18871 (N_18871,N_18661,N_18639);
xor U18872 (N_18872,N_18594,N_18562);
and U18873 (N_18873,N_18515,N_18667);
nor U18874 (N_18874,N_18505,N_18554);
xor U18875 (N_18875,N_18500,N_18561);
nand U18876 (N_18876,N_18655,N_18624);
nor U18877 (N_18877,N_18649,N_18595);
or U18878 (N_18878,N_18603,N_18520);
nor U18879 (N_18879,N_18557,N_18612);
nor U18880 (N_18880,N_18650,N_18564);
nor U18881 (N_18881,N_18597,N_18676);
nor U18882 (N_18882,N_18508,N_18702);
nor U18883 (N_18883,N_18719,N_18624);
nand U18884 (N_18884,N_18612,N_18665);
or U18885 (N_18885,N_18518,N_18686);
nand U18886 (N_18886,N_18699,N_18679);
or U18887 (N_18887,N_18563,N_18669);
or U18888 (N_18888,N_18693,N_18723);
or U18889 (N_18889,N_18542,N_18508);
and U18890 (N_18890,N_18639,N_18505);
or U18891 (N_18891,N_18522,N_18659);
xnor U18892 (N_18892,N_18652,N_18560);
or U18893 (N_18893,N_18585,N_18502);
or U18894 (N_18894,N_18609,N_18676);
nor U18895 (N_18895,N_18680,N_18682);
xnor U18896 (N_18896,N_18510,N_18645);
xnor U18897 (N_18897,N_18691,N_18621);
xnor U18898 (N_18898,N_18664,N_18593);
and U18899 (N_18899,N_18698,N_18662);
xnor U18900 (N_18900,N_18728,N_18535);
xnor U18901 (N_18901,N_18524,N_18673);
xnor U18902 (N_18902,N_18628,N_18555);
xnor U18903 (N_18903,N_18654,N_18557);
nor U18904 (N_18904,N_18745,N_18628);
nand U18905 (N_18905,N_18647,N_18673);
nor U18906 (N_18906,N_18592,N_18731);
nor U18907 (N_18907,N_18688,N_18500);
nor U18908 (N_18908,N_18657,N_18539);
nor U18909 (N_18909,N_18613,N_18515);
xor U18910 (N_18910,N_18743,N_18624);
nor U18911 (N_18911,N_18571,N_18608);
and U18912 (N_18912,N_18672,N_18596);
and U18913 (N_18913,N_18566,N_18663);
xnor U18914 (N_18914,N_18660,N_18648);
or U18915 (N_18915,N_18733,N_18562);
xnor U18916 (N_18916,N_18610,N_18607);
or U18917 (N_18917,N_18530,N_18573);
nor U18918 (N_18918,N_18666,N_18736);
xor U18919 (N_18919,N_18680,N_18593);
or U18920 (N_18920,N_18652,N_18595);
xnor U18921 (N_18921,N_18692,N_18552);
nand U18922 (N_18922,N_18700,N_18522);
nand U18923 (N_18923,N_18596,N_18715);
nor U18924 (N_18924,N_18500,N_18506);
xor U18925 (N_18925,N_18532,N_18564);
nand U18926 (N_18926,N_18579,N_18561);
or U18927 (N_18927,N_18543,N_18710);
nand U18928 (N_18928,N_18575,N_18709);
nand U18929 (N_18929,N_18737,N_18699);
nor U18930 (N_18930,N_18734,N_18743);
nor U18931 (N_18931,N_18565,N_18614);
or U18932 (N_18932,N_18600,N_18602);
nor U18933 (N_18933,N_18743,N_18702);
and U18934 (N_18934,N_18683,N_18500);
xnor U18935 (N_18935,N_18735,N_18704);
nor U18936 (N_18936,N_18666,N_18589);
nand U18937 (N_18937,N_18662,N_18711);
xnor U18938 (N_18938,N_18509,N_18702);
nor U18939 (N_18939,N_18556,N_18617);
nand U18940 (N_18940,N_18573,N_18510);
nor U18941 (N_18941,N_18742,N_18646);
nor U18942 (N_18942,N_18663,N_18693);
and U18943 (N_18943,N_18710,N_18614);
and U18944 (N_18944,N_18716,N_18612);
nor U18945 (N_18945,N_18636,N_18597);
xnor U18946 (N_18946,N_18743,N_18587);
and U18947 (N_18947,N_18577,N_18525);
nor U18948 (N_18948,N_18568,N_18548);
xnor U18949 (N_18949,N_18517,N_18707);
or U18950 (N_18950,N_18635,N_18674);
or U18951 (N_18951,N_18613,N_18731);
nand U18952 (N_18952,N_18737,N_18658);
xnor U18953 (N_18953,N_18500,N_18680);
xor U18954 (N_18954,N_18745,N_18642);
nand U18955 (N_18955,N_18564,N_18573);
or U18956 (N_18956,N_18595,N_18744);
or U18957 (N_18957,N_18709,N_18700);
nand U18958 (N_18958,N_18503,N_18572);
and U18959 (N_18959,N_18605,N_18679);
or U18960 (N_18960,N_18738,N_18579);
or U18961 (N_18961,N_18611,N_18627);
and U18962 (N_18962,N_18688,N_18737);
nor U18963 (N_18963,N_18603,N_18736);
nand U18964 (N_18964,N_18516,N_18705);
xor U18965 (N_18965,N_18562,N_18572);
nand U18966 (N_18966,N_18692,N_18566);
and U18967 (N_18967,N_18504,N_18722);
nor U18968 (N_18968,N_18716,N_18629);
nor U18969 (N_18969,N_18510,N_18707);
or U18970 (N_18970,N_18690,N_18671);
xnor U18971 (N_18971,N_18749,N_18662);
or U18972 (N_18972,N_18737,N_18724);
nor U18973 (N_18973,N_18710,N_18722);
nand U18974 (N_18974,N_18553,N_18660);
nor U18975 (N_18975,N_18505,N_18712);
and U18976 (N_18976,N_18651,N_18648);
and U18977 (N_18977,N_18713,N_18564);
nor U18978 (N_18978,N_18646,N_18514);
xnor U18979 (N_18979,N_18510,N_18647);
and U18980 (N_18980,N_18603,N_18514);
xor U18981 (N_18981,N_18627,N_18529);
nand U18982 (N_18982,N_18615,N_18621);
nand U18983 (N_18983,N_18684,N_18510);
and U18984 (N_18984,N_18669,N_18703);
xor U18985 (N_18985,N_18741,N_18646);
or U18986 (N_18986,N_18538,N_18679);
and U18987 (N_18987,N_18549,N_18729);
nor U18988 (N_18988,N_18612,N_18642);
xor U18989 (N_18989,N_18623,N_18696);
xor U18990 (N_18990,N_18749,N_18515);
and U18991 (N_18991,N_18665,N_18678);
nor U18992 (N_18992,N_18523,N_18630);
or U18993 (N_18993,N_18548,N_18542);
xnor U18994 (N_18994,N_18716,N_18635);
and U18995 (N_18995,N_18576,N_18730);
nand U18996 (N_18996,N_18581,N_18706);
or U18997 (N_18997,N_18600,N_18663);
and U18998 (N_18998,N_18537,N_18512);
nor U18999 (N_18999,N_18565,N_18730);
nor U19000 (N_19000,N_18869,N_18848);
and U19001 (N_19001,N_18960,N_18810);
xnor U19002 (N_19002,N_18913,N_18818);
xor U19003 (N_19003,N_18751,N_18927);
nand U19004 (N_19004,N_18846,N_18896);
nand U19005 (N_19005,N_18767,N_18882);
xnor U19006 (N_19006,N_18973,N_18897);
or U19007 (N_19007,N_18822,N_18983);
or U19008 (N_19008,N_18862,N_18889);
or U19009 (N_19009,N_18934,N_18994);
nand U19010 (N_19010,N_18984,N_18845);
or U19011 (N_19011,N_18932,N_18907);
and U19012 (N_19012,N_18881,N_18791);
nor U19013 (N_19013,N_18854,N_18860);
or U19014 (N_19014,N_18899,N_18976);
xnor U19015 (N_19015,N_18765,N_18925);
and U19016 (N_19016,N_18964,N_18774);
nor U19017 (N_19017,N_18790,N_18781);
nor U19018 (N_19018,N_18877,N_18804);
nor U19019 (N_19019,N_18966,N_18943);
nor U19020 (N_19020,N_18948,N_18884);
and U19021 (N_19021,N_18778,N_18782);
xor U19022 (N_19022,N_18937,N_18788);
xnor U19023 (N_19023,N_18800,N_18861);
or U19024 (N_19024,N_18811,N_18816);
nand U19025 (N_19025,N_18941,N_18820);
or U19026 (N_19026,N_18863,N_18777);
nand U19027 (N_19027,N_18793,N_18933);
nand U19028 (N_19028,N_18894,N_18864);
xnor U19029 (N_19029,N_18796,N_18803);
nand U19030 (N_19030,N_18761,N_18963);
nand U19031 (N_19031,N_18857,N_18829);
nor U19032 (N_19032,N_18794,N_18906);
or U19033 (N_19033,N_18752,N_18888);
nand U19034 (N_19034,N_18987,N_18988);
nand U19035 (N_19035,N_18832,N_18874);
and U19036 (N_19036,N_18850,N_18997);
and U19037 (N_19037,N_18817,N_18944);
and U19038 (N_19038,N_18945,N_18962);
xnor U19039 (N_19039,N_18768,N_18806);
or U19040 (N_19040,N_18965,N_18898);
and U19041 (N_19041,N_18931,N_18799);
and U19042 (N_19042,N_18779,N_18996);
or U19043 (N_19043,N_18904,N_18795);
or U19044 (N_19044,N_18967,N_18903);
nor U19045 (N_19045,N_18947,N_18920);
and U19046 (N_19046,N_18760,N_18910);
nand U19047 (N_19047,N_18815,N_18905);
xor U19048 (N_19048,N_18821,N_18902);
nor U19049 (N_19049,N_18784,N_18926);
nand U19050 (N_19050,N_18866,N_18989);
nor U19051 (N_19051,N_18824,N_18801);
and U19052 (N_19052,N_18823,N_18911);
and U19053 (N_19053,N_18807,N_18859);
nand U19054 (N_19054,N_18879,N_18851);
nor U19055 (N_19055,N_18993,N_18835);
xnor U19056 (N_19056,N_18878,N_18939);
nand U19057 (N_19057,N_18786,N_18827);
xor U19058 (N_19058,N_18758,N_18982);
or U19059 (N_19059,N_18951,N_18955);
nand U19060 (N_19060,N_18969,N_18843);
or U19061 (N_19061,N_18855,N_18954);
nand U19062 (N_19062,N_18938,N_18797);
nor U19063 (N_19063,N_18959,N_18764);
nor U19064 (N_19064,N_18809,N_18792);
or U19065 (N_19065,N_18930,N_18766);
nand U19066 (N_19066,N_18839,N_18756);
nor U19067 (N_19067,N_18853,N_18769);
or U19068 (N_19068,N_18956,N_18952);
nor U19069 (N_19069,N_18814,N_18819);
xor U19070 (N_19070,N_18754,N_18986);
xor U19071 (N_19071,N_18828,N_18880);
nor U19072 (N_19072,N_18841,N_18890);
and U19073 (N_19073,N_18978,N_18950);
or U19074 (N_19074,N_18914,N_18798);
nor U19075 (N_19075,N_18757,N_18928);
and U19076 (N_19076,N_18921,N_18949);
xor U19077 (N_19077,N_18875,N_18852);
xor U19078 (N_19078,N_18961,N_18883);
nor U19079 (N_19079,N_18912,N_18813);
nor U19080 (N_19080,N_18887,N_18980);
and U19081 (N_19081,N_18755,N_18901);
nand U19082 (N_19082,N_18929,N_18773);
xnor U19083 (N_19083,N_18812,N_18916);
or U19084 (N_19084,N_18972,N_18844);
xnor U19085 (N_19085,N_18831,N_18762);
or U19086 (N_19086,N_18974,N_18891);
nand U19087 (N_19087,N_18789,N_18957);
and U19088 (N_19088,N_18876,N_18776);
xor U19089 (N_19089,N_18775,N_18772);
or U19090 (N_19090,N_18856,N_18990);
xor U19091 (N_19091,N_18908,N_18958);
and U19092 (N_19092,N_18895,N_18836);
xor U19093 (N_19093,N_18915,N_18979);
nor U19094 (N_19094,N_18770,N_18942);
or U19095 (N_19095,N_18870,N_18808);
or U19096 (N_19096,N_18985,N_18837);
or U19097 (N_19097,N_18842,N_18759);
or U19098 (N_19098,N_18771,N_18783);
xor U19099 (N_19099,N_18991,N_18998);
xnor U19100 (N_19100,N_18909,N_18826);
nand U19101 (N_19101,N_18935,N_18834);
or U19102 (N_19102,N_18900,N_18873);
and U19103 (N_19103,N_18840,N_18871);
or U19104 (N_19104,N_18992,N_18892);
nor U19105 (N_19105,N_18975,N_18918);
and U19106 (N_19106,N_18886,N_18977);
xor U19107 (N_19107,N_18763,N_18885);
nor U19108 (N_19108,N_18802,N_18923);
or U19109 (N_19109,N_18924,N_18946);
and U19110 (N_19110,N_18849,N_18922);
xor U19111 (N_19111,N_18970,N_18868);
nand U19112 (N_19112,N_18787,N_18750);
nor U19113 (N_19113,N_18968,N_18753);
and U19114 (N_19114,N_18833,N_18838);
and U19115 (N_19115,N_18936,N_18981);
nor U19116 (N_19116,N_18953,N_18847);
xnor U19117 (N_19117,N_18867,N_18785);
nand U19118 (N_19118,N_18917,N_18805);
xor U19119 (N_19119,N_18999,N_18995);
xnor U19120 (N_19120,N_18780,N_18865);
nand U19121 (N_19121,N_18858,N_18893);
nor U19122 (N_19122,N_18825,N_18830);
xor U19123 (N_19123,N_18940,N_18872);
nor U19124 (N_19124,N_18919,N_18971);
and U19125 (N_19125,N_18930,N_18946);
nand U19126 (N_19126,N_18860,N_18766);
and U19127 (N_19127,N_18965,N_18933);
or U19128 (N_19128,N_18869,N_18907);
or U19129 (N_19129,N_18837,N_18884);
or U19130 (N_19130,N_18898,N_18883);
xor U19131 (N_19131,N_18951,N_18833);
nor U19132 (N_19132,N_18757,N_18763);
nor U19133 (N_19133,N_18783,N_18970);
nand U19134 (N_19134,N_18924,N_18779);
nor U19135 (N_19135,N_18974,N_18973);
xor U19136 (N_19136,N_18885,N_18975);
xnor U19137 (N_19137,N_18947,N_18850);
nand U19138 (N_19138,N_18896,N_18828);
nand U19139 (N_19139,N_18929,N_18962);
or U19140 (N_19140,N_18967,N_18843);
nor U19141 (N_19141,N_18762,N_18955);
nand U19142 (N_19142,N_18953,N_18855);
or U19143 (N_19143,N_18777,N_18928);
nand U19144 (N_19144,N_18962,N_18817);
or U19145 (N_19145,N_18835,N_18784);
nand U19146 (N_19146,N_18878,N_18861);
nand U19147 (N_19147,N_18988,N_18901);
nand U19148 (N_19148,N_18752,N_18866);
nand U19149 (N_19149,N_18890,N_18823);
or U19150 (N_19150,N_18956,N_18970);
xor U19151 (N_19151,N_18905,N_18758);
and U19152 (N_19152,N_18875,N_18766);
nand U19153 (N_19153,N_18858,N_18822);
or U19154 (N_19154,N_18766,N_18822);
nor U19155 (N_19155,N_18927,N_18805);
nor U19156 (N_19156,N_18874,N_18995);
nand U19157 (N_19157,N_18986,N_18924);
xnor U19158 (N_19158,N_18955,N_18840);
xnor U19159 (N_19159,N_18775,N_18938);
nand U19160 (N_19160,N_18925,N_18900);
xnor U19161 (N_19161,N_18799,N_18783);
and U19162 (N_19162,N_18782,N_18853);
and U19163 (N_19163,N_18848,N_18842);
and U19164 (N_19164,N_18805,N_18942);
and U19165 (N_19165,N_18798,N_18843);
xnor U19166 (N_19166,N_18964,N_18908);
and U19167 (N_19167,N_18979,N_18843);
nor U19168 (N_19168,N_18851,N_18792);
or U19169 (N_19169,N_18898,N_18938);
xor U19170 (N_19170,N_18902,N_18952);
and U19171 (N_19171,N_18787,N_18784);
or U19172 (N_19172,N_18809,N_18965);
xor U19173 (N_19173,N_18942,N_18832);
xor U19174 (N_19174,N_18753,N_18784);
nor U19175 (N_19175,N_18986,N_18943);
nand U19176 (N_19176,N_18756,N_18933);
xor U19177 (N_19177,N_18802,N_18909);
xnor U19178 (N_19178,N_18780,N_18889);
and U19179 (N_19179,N_18999,N_18964);
xor U19180 (N_19180,N_18856,N_18897);
and U19181 (N_19181,N_18825,N_18867);
nand U19182 (N_19182,N_18998,N_18931);
xnor U19183 (N_19183,N_18926,N_18855);
xnor U19184 (N_19184,N_18946,N_18879);
or U19185 (N_19185,N_18984,N_18982);
nor U19186 (N_19186,N_18803,N_18856);
nand U19187 (N_19187,N_18839,N_18877);
nand U19188 (N_19188,N_18806,N_18811);
nand U19189 (N_19189,N_18866,N_18799);
and U19190 (N_19190,N_18880,N_18898);
nand U19191 (N_19191,N_18827,N_18891);
nand U19192 (N_19192,N_18835,N_18989);
nor U19193 (N_19193,N_18828,N_18928);
and U19194 (N_19194,N_18980,N_18903);
and U19195 (N_19195,N_18792,N_18789);
or U19196 (N_19196,N_18926,N_18847);
xor U19197 (N_19197,N_18763,N_18865);
and U19198 (N_19198,N_18885,N_18753);
and U19199 (N_19199,N_18819,N_18985);
or U19200 (N_19200,N_18806,N_18794);
or U19201 (N_19201,N_18956,N_18914);
nand U19202 (N_19202,N_18948,N_18997);
and U19203 (N_19203,N_18754,N_18786);
xnor U19204 (N_19204,N_18958,N_18856);
or U19205 (N_19205,N_18800,N_18843);
nand U19206 (N_19206,N_18773,N_18778);
nand U19207 (N_19207,N_18752,N_18811);
xor U19208 (N_19208,N_18985,N_18941);
xnor U19209 (N_19209,N_18901,N_18821);
nor U19210 (N_19210,N_18875,N_18931);
nand U19211 (N_19211,N_18901,N_18886);
nor U19212 (N_19212,N_18912,N_18871);
nor U19213 (N_19213,N_18989,N_18810);
nor U19214 (N_19214,N_18868,N_18969);
xnor U19215 (N_19215,N_18924,N_18847);
or U19216 (N_19216,N_18864,N_18956);
nor U19217 (N_19217,N_18776,N_18790);
and U19218 (N_19218,N_18833,N_18811);
nor U19219 (N_19219,N_18754,N_18952);
nand U19220 (N_19220,N_18758,N_18939);
xnor U19221 (N_19221,N_18930,N_18782);
xnor U19222 (N_19222,N_18774,N_18803);
or U19223 (N_19223,N_18772,N_18999);
xnor U19224 (N_19224,N_18936,N_18818);
or U19225 (N_19225,N_18904,N_18753);
nor U19226 (N_19226,N_18920,N_18791);
xnor U19227 (N_19227,N_18782,N_18791);
xnor U19228 (N_19228,N_18938,N_18963);
or U19229 (N_19229,N_18786,N_18854);
or U19230 (N_19230,N_18802,N_18800);
or U19231 (N_19231,N_18816,N_18944);
xor U19232 (N_19232,N_18782,N_18983);
xnor U19233 (N_19233,N_18906,N_18826);
and U19234 (N_19234,N_18895,N_18969);
xor U19235 (N_19235,N_18991,N_18794);
xor U19236 (N_19236,N_18985,N_18810);
nand U19237 (N_19237,N_18992,N_18802);
or U19238 (N_19238,N_18945,N_18991);
or U19239 (N_19239,N_18932,N_18780);
and U19240 (N_19240,N_18873,N_18943);
or U19241 (N_19241,N_18768,N_18812);
or U19242 (N_19242,N_18940,N_18833);
nand U19243 (N_19243,N_18806,N_18988);
nand U19244 (N_19244,N_18910,N_18814);
and U19245 (N_19245,N_18895,N_18948);
xor U19246 (N_19246,N_18782,N_18774);
and U19247 (N_19247,N_18991,N_18976);
and U19248 (N_19248,N_18761,N_18767);
xnor U19249 (N_19249,N_18998,N_18778);
nand U19250 (N_19250,N_19197,N_19157);
xor U19251 (N_19251,N_19223,N_19145);
and U19252 (N_19252,N_19220,N_19176);
xnor U19253 (N_19253,N_19123,N_19034);
xor U19254 (N_19254,N_19066,N_19137);
nor U19255 (N_19255,N_19142,N_19160);
and U19256 (N_19256,N_19010,N_19083);
and U19257 (N_19257,N_19149,N_19241);
xnor U19258 (N_19258,N_19048,N_19165);
or U19259 (N_19259,N_19141,N_19063);
or U19260 (N_19260,N_19093,N_19042);
nor U19261 (N_19261,N_19064,N_19085);
nor U19262 (N_19262,N_19043,N_19130);
xor U19263 (N_19263,N_19051,N_19013);
nor U19264 (N_19264,N_19110,N_19174);
nor U19265 (N_19265,N_19041,N_19221);
nor U19266 (N_19266,N_19072,N_19055);
xor U19267 (N_19267,N_19001,N_19092);
or U19268 (N_19268,N_19112,N_19222);
and U19269 (N_19269,N_19074,N_19186);
nand U19270 (N_19270,N_19089,N_19070);
and U19271 (N_19271,N_19080,N_19017);
and U19272 (N_19272,N_19067,N_19114);
xnor U19273 (N_19273,N_19209,N_19007);
and U19274 (N_19274,N_19162,N_19029);
xnor U19275 (N_19275,N_19039,N_19182);
and U19276 (N_19276,N_19204,N_19213);
or U19277 (N_19277,N_19090,N_19033);
nor U19278 (N_19278,N_19062,N_19179);
nand U19279 (N_19279,N_19231,N_19103);
nor U19280 (N_19280,N_19107,N_19216);
xnor U19281 (N_19281,N_19138,N_19187);
and U19282 (N_19282,N_19206,N_19205);
nand U19283 (N_19283,N_19100,N_19075);
xnor U19284 (N_19284,N_19247,N_19242);
or U19285 (N_19285,N_19234,N_19136);
and U19286 (N_19286,N_19191,N_19022);
nor U19287 (N_19287,N_19009,N_19188);
and U19288 (N_19288,N_19069,N_19211);
xor U19289 (N_19289,N_19077,N_19170);
xor U19290 (N_19290,N_19053,N_19151);
nand U19291 (N_19291,N_19230,N_19104);
nor U19292 (N_19292,N_19208,N_19054);
xor U19293 (N_19293,N_19030,N_19134);
nand U19294 (N_19294,N_19147,N_19108);
and U19295 (N_19295,N_19203,N_19016);
nor U19296 (N_19296,N_19015,N_19046);
and U19297 (N_19297,N_19244,N_19236);
or U19298 (N_19298,N_19012,N_19228);
nand U19299 (N_19299,N_19031,N_19095);
nor U19300 (N_19300,N_19200,N_19132);
xnor U19301 (N_19301,N_19082,N_19181);
xor U19302 (N_19302,N_19225,N_19172);
or U19303 (N_19303,N_19150,N_19117);
nor U19304 (N_19304,N_19192,N_19232);
or U19305 (N_19305,N_19105,N_19018);
nand U19306 (N_19306,N_19003,N_19248);
or U19307 (N_19307,N_19180,N_19101);
and U19308 (N_19308,N_19226,N_19146);
nand U19309 (N_19309,N_19195,N_19097);
xnor U19310 (N_19310,N_19159,N_19058);
nand U19311 (N_19311,N_19037,N_19087);
or U19312 (N_19312,N_19086,N_19217);
and U19313 (N_19313,N_19128,N_19219);
nand U19314 (N_19314,N_19056,N_19027);
or U19315 (N_19315,N_19148,N_19246);
nor U19316 (N_19316,N_19189,N_19059);
nand U19317 (N_19317,N_19088,N_19040);
and U19318 (N_19318,N_19152,N_19049);
nor U19319 (N_19319,N_19238,N_19071);
or U19320 (N_19320,N_19143,N_19036);
and U19321 (N_19321,N_19073,N_19173);
nand U19322 (N_19322,N_19233,N_19032);
and U19323 (N_19323,N_19050,N_19166);
or U19324 (N_19324,N_19118,N_19155);
and U19325 (N_19325,N_19168,N_19196);
xnor U19326 (N_19326,N_19183,N_19127);
or U19327 (N_19327,N_19124,N_19091);
nand U19328 (N_19328,N_19214,N_19158);
and U19329 (N_19329,N_19115,N_19240);
xnor U19330 (N_19330,N_19178,N_19079);
nand U19331 (N_19331,N_19239,N_19135);
and U19332 (N_19332,N_19000,N_19065);
nor U19333 (N_19333,N_19212,N_19052);
and U19334 (N_19334,N_19177,N_19201);
or U19335 (N_19335,N_19153,N_19194);
xnor U19336 (N_19336,N_19119,N_19061);
nor U19337 (N_19337,N_19161,N_19154);
or U19338 (N_19338,N_19126,N_19207);
and U19339 (N_19339,N_19020,N_19035);
or U19340 (N_19340,N_19025,N_19006);
xor U19341 (N_19341,N_19129,N_19023);
xor U19342 (N_19342,N_19045,N_19109);
or U19343 (N_19343,N_19175,N_19215);
and U19344 (N_19344,N_19084,N_19004);
and U19345 (N_19345,N_19193,N_19224);
nor U19346 (N_19346,N_19106,N_19122);
nor U19347 (N_19347,N_19057,N_19199);
or U19348 (N_19348,N_19094,N_19026);
xor U19349 (N_19349,N_19229,N_19185);
nor U19350 (N_19350,N_19156,N_19008);
xnor U19351 (N_19351,N_19081,N_19198);
xnor U19352 (N_19352,N_19164,N_19005);
xnor U19353 (N_19353,N_19227,N_19171);
nand U19354 (N_19354,N_19099,N_19011);
nand U19355 (N_19355,N_19120,N_19121);
xnor U19356 (N_19356,N_19190,N_19218);
nand U19357 (N_19357,N_19014,N_19140);
or U19358 (N_19358,N_19021,N_19044);
nand U19359 (N_19359,N_19144,N_19133);
and U19360 (N_19360,N_19028,N_19169);
nand U19361 (N_19361,N_19210,N_19076);
nand U19362 (N_19362,N_19019,N_19002);
or U19363 (N_19363,N_19235,N_19111);
or U19364 (N_19364,N_19184,N_19202);
or U19365 (N_19365,N_19243,N_19131);
xnor U19366 (N_19366,N_19098,N_19024);
nand U19367 (N_19367,N_19167,N_19102);
nand U19368 (N_19368,N_19163,N_19245);
or U19369 (N_19369,N_19078,N_19116);
nor U19370 (N_19370,N_19125,N_19139);
or U19371 (N_19371,N_19047,N_19249);
nand U19372 (N_19372,N_19113,N_19038);
nand U19373 (N_19373,N_19096,N_19068);
nor U19374 (N_19374,N_19237,N_19060);
and U19375 (N_19375,N_19130,N_19236);
nand U19376 (N_19376,N_19053,N_19110);
nand U19377 (N_19377,N_19084,N_19142);
nor U19378 (N_19378,N_19065,N_19021);
and U19379 (N_19379,N_19191,N_19048);
and U19380 (N_19380,N_19125,N_19167);
or U19381 (N_19381,N_19227,N_19090);
and U19382 (N_19382,N_19116,N_19122);
nor U19383 (N_19383,N_19062,N_19204);
and U19384 (N_19384,N_19123,N_19121);
and U19385 (N_19385,N_19196,N_19215);
and U19386 (N_19386,N_19009,N_19125);
xnor U19387 (N_19387,N_19244,N_19230);
or U19388 (N_19388,N_19013,N_19088);
or U19389 (N_19389,N_19172,N_19022);
xor U19390 (N_19390,N_19132,N_19014);
nand U19391 (N_19391,N_19197,N_19076);
and U19392 (N_19392,N_19150,N_19000);
nor U19393 (N_19393,N_19107,N_19224);
and U19394 (N_19394,N_19054,N_19245);
xnor U19395 (N_19395,N_19223,N_19187);
nor U19396 (N_19396,N_19149,N_19136);
nand U19397 (N_19397,N_19146,N_19187);
nor U19398 (N_19398,N_19011,N_19133);
xor U19399 (N_19399,N_19195,N_19074);
xnor U19400 (N_19400,N_19110,N_19016);
or U19401 (N_19401,N_19155,N_19094);
nor U19402 (N_19402,N_19166,N_19002);
xnor U19403 (N_19403,N_19227,N_19099);
and U19404 (N_19404,N_19231,N_19248);
nor U19405 (N_19405,N_19143,N_19190);
and U19406 (N_19406,N_19024,N_19235);
or U19407 (N_19407,N_19055,N_19146);
nor U19408 (N_19408,N_19185,N_19006);
xnor U19409 (N_19409,N_19055,N_19086);
nor U19410 (N_19410,N_19183,N_19061);
xnor U19411 (N_19411,N_19184,N_19139);
xor U19412 (N_19412,N_19247,N_19118);
xor U19413 (N_19413,N_19234,N_19224);
xor U19414 (N_19414,N_19035,N_19091);
and U19415 (N_19415,N_19155,N_19049);
xnor U19416 (N_19416,N_19242,N_19161);
or U19417 (N_19417,N_19247,N_19094);
or U19418 (N_19418,N_19203,N_19226);
xor U19419 (N_19419,N_19039,N_19078);
or U19420 (N_19420,N_19103,N_19230);
xor U19421 (N_19421,N_19105,N_19070);
or U19422 (N_19422,N_19139,N_19156);
xor U19423 (N_19423,N_19063,N_19047);
or U19424 (N_19424,N_19168,N_19231);
or U19425 (N_19425,N_19156,N_19228);
and U19426 (N_19426,N_19208,N_19218);
nor U19427 (N_19427,N_19231,N_19242);
nand U19428 (N_19428,N_19246,N_19052);
nand U19429 (N_19429,N_19194,N_19079);
nand U19430 (N_19430,N_19090,N_19169);
and U19431 (N_19431,N_19233,N_19040);
and U19432 (N_19432,N_19112,N_19218);
xor U19433 (N_19433,N_19177,N_19056);
xnor U19434 (N_19434,N_19174,N_19225);
xnor U19435 (N_19435,N_19203,N_19009);
or U19436 (N_19436,N_19173,N_19021);
or U19437 (N_19437,N_19165,N_19238);
nand U19438 (N_19438,N_19039,N_19168);
nand U19439 (N_19439,N_19185,N_19034);
nor U19440 (N_19440,N_19229,N_19066);
and U19441 (N_19441,N_19246,N_19178);
and U19442 (N_19442,N_19010,N_19146);
nor U19443 (N_19443,N_19151,N_19107);
nor U19444 (N_19444,N_19241,N_19076);
and U19445 (N_19445,N_19243,N_19192);
nor U19446 (N_19446,N_19194,N_19138);
and U19447 (N_19447,N_19150,N_19068);
and U19448 (N_19448,N_19201,N_19127);
nand U19449 (N_19449,N_19153,N_19081);
xor U19450 (N_19450,N_19031,N_19114);
nor U19451 (N_19451,N_19125,N_19109);
or U19452 (N_19452,N_19090,N_19211);
and U19453 (N_19453,N_19065,N_19129);
or U19454 (N_19454,N_19127,N_19200);
xnor U19455 (N_19455,N_19135,N_19120);
nand U19456 (N_19456,N_19194,N_19240);
nor U19457 (N_19457,N_19197,N_19127);
nand U19458 (N_19458,N_19028,N_19208);
nor U19459 (N_19459,N_19169,N_19201);
xor U19460 (N_19460,N_19123,N_19029);
xnor U19461 (N_19461,N_19130,N_19054);
nor U19462 (N_19462,N_19094,N_19149);
or U19463 (N_19463,N_19137,N_19240);
nor U19464 (N_19464,N_19147,N_19166);
xnor U19465 (N_19465,N_19200,N_19223);
nor U19466 (N_19466,N_19206,N_19179);
or U19467 (N_19467,N_19223,N_19121);
and U19468 (N_19468,N_19088,N_19090);
nand U19469 (N_19469,N_19165,N_19002);
xor U19470 (N_19470,N_19116,N_19123);
nor U19471 (N_19471,N_19007,N_19245);
and U19472 (N_19472,N_19175,N_19134);
nor U19473 (N_19473,N_19197,N_19207);
nand U19474 (N_19474,N_19104,N_19201);
nand U19475 (N_19475,N_19113,N_19017);
xnor U19476 (N_19476,N_19049,N_19150);
or U19477 (N_19477,N_19198,N_19076);
nor U19478 (N_19478,N_19220,N_19057);
nand U19479 (N_19479,N_19233,N_19190);
xor U19480 (N_19480,N_19221,N_19084);
xnor U19481 (N_19481,N_19137,N_19207);
or U19482 (N_19482,N_19215,N_19117);
and U19483 (N_19483,N_19178,N_19222);
or U19484 (N_19484,N_19249,N_19132);
nor U19485 (N_19485,N_19197,N_19030);
xnor U19486 (N_19486,N_19042,N_19026);
nand U19487 (N_19487,N_19075,N_19172);
xor U19488 (N_19488,N_19059,N_19247);
or U19489 (N_19489,N_19010,N_19078);
or U19490 (N_19490,N_19159,N_19158);
and U19491 (N_19491,N_19157,N_19065);
xor U19492 (N_19492,N_19240,N_19015);
nand U19493 (N_19493,N_19182,N_19005);
and U19494 (N_19494,N_19234,N_19199);
xor U19495 (N_19495,N_19097,N_19247);
and U19496 (N_19496,N_19122,N_19189);
xor U19497 (N_19497,N_19031,N_19152);
and U19498 (N_19498,N_19022,N_19113);
nor U19499 (N_19499,N_19215,N_19080);
nor U19500 (N_19500,N_19459,N_19480);
and U19501 (N_19501,N_19408,N_19377);
xor U19502 (N_19502,N_19359,N_19320);
and U19503 (N_19503,N_19313,N_19469);
xnor U19504 (N_19504,N_19422,N_19447);
nand U19505 (N_19505,N_19337,N_19276);
nor U19506 (N_19506,N_19267,N_19297);
nor U19507 (N_19507,N_19454,N_19354);
nand U19508 (N_19508,N_19431,N_19277);
and U19509 (N_19509,N_19410,N_19293);
or U19510 (N_19510,N_19365,N_19371);
or U19511 (N_19511,N_19380,N_19455);
and U19512 (N_19512,N_19271,N_19258);
or U19513 (N_19513,N_19483,N_19491);
nor U19514 (N_19514,N_19304,N_19299);
and U19515 (N_19515,N_19294,N_19362);
nor U19516 (N_19516,N_19384,N_19372);
xnor U19517 (N_19517,N_19487,N_19340);
nand U19518 (N_19518,N_19460,N_19474);
and U19519 (N_19519,N_19386,N_19498);
or U19520 (N_19520,N_19291,N_19265);
nand U19521 (N_19521,N_19256,N_19451);
nor U19522 (N_19522,N_19368,N_19433);
or U19523 (N_19523,N_19301,N_19306);
nor U19524 (N_19524,N_19432,N_19349);
nand U19525 (N_19525,N_19419,N_19444);
and U19526 (N_19526,N_19441,N_19353);
or U19527 (N_19527,N_19281,N_19479);
nand U19528 (N_19528,N_19295,N_19318);
nand U19529 (N_19529,N_19466,N_19450);
and U19530 (N_19530,N_19350,N_19427);
and U19531 (N_19531,N_19457,N_19310);
nand U19532 (N_19532,N_19413,N_19486);
or U19533 (N_19533,N_19407,N_19425);
xor U19534 (N_19534,N_19328,N_19330);
xor U19535 (N_19535,N_19415,N_19379);
or U19536 (N_19536,N_19401,N_19395);
xnor U19537 (N_19537,N_19333,N_19315);
or U19538 (N_19538,N_19331,N_19387);
nand U19539 (N_19539,N_19376,N_19428);
xnor U19540 (N_19540,N_19282,N_19250);
nand U19541 (N_19541,N_19290,N_19280);
nor U19542 (N_19542,N_19437,N_19311);
nor U19543 (N_19543,N_19268,N_19373);
nor U19544 (N_19544,N_19287,N_19283);
and U19545 (N_19545,N_19251,N_19485);
and U19546 (N_19546,N_19493,N_19452);
and U19547 (N_19547,N_19322,N_19332);
nand U19548 (N_19548,N_19321,N_19495);
and U19549 (N_19549,N_19274,N_19461);
nor U19550 (N_19550,N_19292,N_19475);
or U19551 (N_19551,N_19476,N_19423);
nand U19552 (N_19552,N_19358,N_19468);
or U19553 (N_19553,N_19346,N_19388);
nor U19554 (N_19554,N_19446,N_19254);
xor U19555 (N_19555,N_19382,N_19329);
xor U19556 (N_19556,N_19352,N_19307);
nor U19557 (N_19557,N_19477,N_19343);
and U19558 (N_19558,N_19478,N_19300);
nor U19559 (N_19559,N_19393,N_19374);
and U19560 (N_19560,N_19488,N_19284);
xor U19561 (N_19561,N_19309,N_19302);
nand U19562 (N_19562,N_19490,N_19471);
nand U19563 (N_19563,N_19378,N_19449);
xor U19564 (N_19564,N_19253,N_19473);
xnor U19565 (N_19565,N_19399,N_19312);
xnor U19566 (N_19566,N_19335,N_19339);
xor U19567 (N_19567,N_19314,N_19356);
or U19568 (N_19568,N_19397,N_19308);
xnor U19569 (N_19569,N_19420,N_19484);
nand U19570 (N_19570,N_19336,N_19448);
nand U19571 (N_19571,N_19344,N_19467);
xnor U19572 (N_19572,N_19348,N_19497);
or U19573 (N_19573,N_19255,N_19443);
nand U19574 (N_19574,N_19355,N_19430);
xnor U19575 (N_19575,N_19481,N_19470);
xnor U19576 (N_19576,N_19319,N_19398);
nand U19577 (N_19577,N_19385,N_19435);
or U19578 (N_19578,N_19463,N_19416);
nor U19579 (N_19579,N_19252,N_19424);
or U19580 (N_19580,N_19275,N_19323);
or U19581 (N_19581,N_19264,N_19260);
or U19582 (N_19582,N_19496,N_19499);
and U19583 (N_19583,N_19472,N_19357);
nand U19584 (N_19584,N_19404,N_19289);
and U19585 (N_19585,N_19325,N_19278);
xor U19586 (N_19586,N_19489,N_19361);
and U19587 (N_19587,N_19341,N_19411);
or U19588 (N_19588,N_19412,N_19262);
nor U19589 (N_19589,N_19429,N_19286);
xnor U19590 (N_19590,N_19438,N_19442);
nand U19591 (N_19591,N_19381,N_19418);
nor U19592 (N_19592,N_19370,N_19279);
nor U19593 (N_19593,N_19273,N_19367);
or U19594 (N_19594,N_19270,N_19327);
or U19595 (N_19595,N_19338,N_19263);
and U19596 (N_19596,N_19400,N_19464);
and U19597 (N_19597,N_19405,N_19494);
nand U19598 (N_19598,N_19439,N_19296);
and U19599 (N_19599,N_19305,N_19363);
or U19600 (N_19600,N_19465,N_19317);
and U19601 (N_19601,N_19257,N_19414);
nor U19602 (N_19602,N_19456,N_19417);
nor U19603 (N_19603,N_19426,N_19266);
xnor U19604 (N_19604,N_19303,N_19406);
and U19605 (N_19605,N_19421,N_19326);
nand U19606 (N_19606,N_19392,N_19360);
nor U19607 (N_19607,N_19434,N_19316);
and U19608 (N_19608,N_19261,N_19403);
and U19609 (N_19609,N_19402,N_19351);
nor U19610 (N_19610,N_19334,N_19345);
xor U19611 (N_19611,N_19462,N_19285);
or U19612 (N_19612,N_19458,N_19389);
xnor U19613 (N_19613,N_19342,N_19391);
or U19614 (N_19614,N_19375,N_19269);
nand U19615 (N_19615,N_19324,N_19396);
nor U19616 (N_19616,N_19364,N_19440);
and U19617 (N_19617,N_19347,N_19453);
nor U19618 (N_19618,N_19394,N_19445);
nor U19619 (N_19619,N_19383,N_19259);
nor U19620 (N_19620,N_19409,N_19482);
and U19621 (N_19621,N_19390,N_19366);
or U19622 (N_19622,N_19436,N_19298);
nand U19623 (N_19623,N_19288,N_19369);
nand U19624 (N_19624,N_19272,N_19492);
nand U19625 (N_19625,N_19325,N_19473);
or U19626 (N_19626,N_19329,N_19412);
nand U19627 (N_19627,N_19479,N_19440);
xnor U19628 (N_19628,N_19319,N_19465);
nand U19629 (N_19629,N_19354,N_19312);
nor U19630 (N_19630,N_19302,N_19384);
nor U19631 (N_19631,N_19396,N_19379);
xnor U19632 (N_19632,N_19498,N_19450);
nor U19633 (N_19633,N_19318,N_19275);
nand U19634 (N_19634,N_19296,N_19417);
or U19635 (N_19635,N_19465,N_19254);
and U19636 (N_19636,N_19468,N_19424);
xor U19637 (N_19637,N_19341,N_19328);
nand U19638 (N_19638,N_19424,N_19410);
or U19639 (N_19639,N_19285,N_19442);
nor U19640 (N_19640,N_19349,N_19413);
xnor U19641 (N_19641,N_19368,N_19280);
or U19642 (N_19642,N_19433,N_19497);
nand U19643 (N_19643,N_19403,N_19499);
nand U19644 (N_19644,N_19379,N_19407);
nor U19645 (N_19645,N_19265,N_19407);
and U19646 (N_19646,N_19460,N_19471);
and U19647 (N_19647,N_19411,N_19396);
or U19648 (N_19648,N_19435,N_19272);
or U19649 (N_19649,N_19337,N_19427);
nor U19650 (N_19650,N_19391,N_19299);
nor U19651 (N_19651,N_19446,N_19404);
and U19652 (N_19652,N_19274,N_19325);
nand U19653 (N_19653,N_19259,N_19363);
nand U19654 (N_19654,N_19447,N_19457);
xor U19655 (N_19655,N_19485,N_19411);
nor U19656 (N_19656,N_19418,N_19368);
nor U19657 (N_19657,N_19451,N_19453);
nor U19658 (N_19658,N_19357,N_19337);
nor U19659 (N_19659,N_19316,N_19267);
and U19660 (N_19660,N_19488,N_19411);
nand U19661 (N_19661,N_19357,N_19311);
nand U19662 (N_19662,N_19410,N_19323);
xnor U19663 (N_19663,N_19277,N_19334);
or U19664 (N_19664,N_19373,N_19362);
or U19665 (N_19665,N_19358,N_19474);
nor U19666 (N_19666,N_19317,N_19488);
or U19667 (N_19667,N_19272,N_19316);
nand U19668 (N_19668,N_19281,N_19439);
and U19669 (N_19669,N_19333,N_19451);
and U19670 (N_19670,N_19446,N_19307);
nor U19671 (N_19671,N_19427,N_19381);
nor U19672 (N_19672,N_19321,N_19370);
nor U19673 (N_19673,N_19313,N_19412);
xor U19674 (N_19674,N_19457,N_19486);
nor U19675 (N_19675,N_19413,N_19423);
or U19676 (N_19676,N_19309,N_19306);
nor U19677 (N_19677,N_19297,N_19421);
or U19678 (N_19678,N_19484,N_19281);
nand U19679 (N_19679,N_19307,N_19496);
or U19680 (N_19680,N_19481,N_19401);
and U19681 (N_19681,N_19393,N_19366);
or U19682 (N_19682,N_19317,N_19478);
nor U19683 (N_19683,N_19393,N_19300);
or U19684 (N_19684,N_19419,N_19388);
nor U19685 (N_19685,N_19251,N_19347);
xnor U19686 (N_19686,N_19413,N_19497);
nand U19687 (N_19687,N_19258,N_19270);
or U19688 (N_19688,N_19435,N_19398);
xor U19689 (N_19689,N_19478,N_19437);
and U19690 (N_19690,N_19372,N_19434);
or U19691 (N_19691,N_19319,N_19493);
xnor U19692 (N_19692,N_19485,N_19358);
and U19693 (N_19693,N_19469,N_19333);
xor U19694 (N_19694,N_19470,N_19323);
and U19695 (N_19695,N_19273,N_19300);
and U19696 (N_19696,N_19343,N_19499);
nand U19697 (N_19697,N_19493,N_19398);
nand U19698 (N_19698,N_19422,N_19407);
and U19699 (N_19699,N_19431,N_19499);
nor U19700 (N_19700,N_19310,N_19288);
and U19701 (N_19701,N_19339,N_19310);
nor U19702 (N_19702,N_19376,N_19304);
xnor U19703 (N_19703,N_19363,N_19430);
and U19704 (N_19704,N_19429,N_19468);
nand U19705 (N_19705,N_19279,N_19441);
nor U19706 (N_19706,N_19485,N_19310);
nand U19707 (N_19707,N_19327,N_19401);
xor U19708 (N_19708,N_19422,N_19438);
xnor U19709 (N_19709,N_19402,N_19440);
nor U19710 (N_19710,N_19491,N_19430);
nand U19711 (N_19711,N_19342,N_19274);
xnor U19712 (N_19712,N_19448,N_19415);
nor U19713 (N_19713,N_19446,N_19286);
and U19714 (N_19714,N_19389,N_19426);
nor U19715 (N_19715,N_19254,N_19279);
xnor U19716 (N_19716,N_19294,N_19401);
xor U19717 (N_19717,N_19269,N_19378);
xor U19718 (N_19718,N_19414,N_19451);
nor U19719 (N_19719,N_19389,N_19437);
nand U19720 (N_19720,N_19309,N_19342);
nor U19721 (N_19721,N_19480,N_19428);
and U19722 (N_19722,N_19341,N_19425);
and U19723 (N_19723,N_19396,N_19361);
nand U19724 (N_19724,N_19340,N_19283);
and U19725 (N_19725,N_19441,N_19434);
nand U19726 (N_19726,N_19287,N_19265);
or U19727 (N_19727,N_19307,N_19464);
or U19728 (N_19728,N_19265,N_19331);
xor U19729 (N_19729,N_19274,N_19387);
and U19730 (N_19730,N_19316,N_19418);
nor U19731 (N_19731,N_19352,N_19390);
or U19732 (N_19732,N_19417,N_19317);
and U19733 (N_19733,N_19468,N_19386);
and U19734 (N_19734,N_19327,N_19369);
nand U19735 (N_19735,N_19437,N_19475);
nor U19736 (N_19736,N_19285,N_19465);
and U19737 (N_19737,N_19492,N_19313);
xor U19738 (N_19738,N_19375,N_19413);
or U19739 (N_19739,N_19386,N_19486);
nor U19740 (N_19740,N_19459,N_19361);
xnor U19741 (N_19741,N_19297,N_19253);
nor U19742 (N_19742,N_19369,N_19285);
and U19743 (N_19743,N_19373,N_19370);
nand U19744 (N_19744,N_19308,N_19485);
or U19745 (N_19745,N_19402,N_19379);
nor U19746 (N_19746,N_19479,N_19462);
or U19747 (N_19747,N_19401,N_19477);
xor U19748 (N_19748,N_19328,N_19308);
nand U19749 (N_19749,N_19251,N_19308);
or U19750 (N_19750,N_19694,N_19532);
and U19751 (N_19751,N_19632,N_19693);
nor U19752 (N_19752,N_19698,N_19644);
nor U19753 (N_19753,N_19583,N_19745);
nor U19754 (N_19754,N_19727,N_19623);
xor U19755 (N_19755,N_19595,N_19688);
and U19756 (N_19756,N_19502,N_19507);
xnor U19757 (N_19757,N_19548,N_19598);
and U19758 (N_19758,N_19655,N_19656);
nor U19759 (N_19759,N_19657,N_19633);
nand U19760 (N_19760,N_19530,N_19747);
nor U19761 (N_19761,N_19609,N_19631);
or U19762 (N_19762,N_19602,N_19640);
xor U19763 (N_19763,N_19738,N_19739);
and U19764 (N_19764,N_19718,N_19552);
or U19765 (N_19765,N_19550,N_19500);
nand U19766 (N_19766,N_19725,N_19549);
xor U19767 (N_19767,N_19674,N_19638);
and U19768 (N_19768,N_19586,N_19710);
nor U19769 (N_19769,N_19746,N_19707);
nand U19770 (N_19770,N_19663,N_19729);
xnor U19771 (N_19771,N_19683,N_19510);
xor U19772 (N_19772,N_19614,N_19721);
and U19773 (N_19773,N_19579,N_19506);
and U19774 (N_19774,N_19538,N_19643);
xnor U19775 (N_19775,N_19514,N_19553);
nor U19776 (N_19776,N_19679,N_19515);
nor U19777 (N_19777,N_19705,N_19650);
or U19778 (N_19778,N_19678,N_19547);
and U19779 (N_19779,N_19642,N_19733);
nand U19780 (N_19780,N_19726,N_19566);
xor U19781 (N_19781,N_19567,N_19735);
nor U19782 (N_19782,N_19607,N_19653);
nor U19783 (N_19783,N_19648,N_19513);
and U19784 (N_19784,N_19596,N_19569);
nand U19785 (N_19785,N_19749,N_19524);
nor U19786 (N_19786,N_19554,N_19531);
xnor U19787 (N_19787,N_19731,N_19691);
xnor U19788 (N_19788,N_19668,N_19543);
or U19789 (N_19789,N_19702,N_19516);
nor U19790 (N_19790,N_19520,N_19621);
or U19791 (N_19791,N_19574,N_19700);
nor U19792 (N_19792,N_19673,N_19615);
or U19793 (N_19793,N_19573,N_19564);
and U19794 (N_19794,N_19692,N_19584);
and U19795 (N_19795,N_19744,N_19723);
xor U19796 (N_19796,N_19539,N_19713);
and U19797 (N_19797,N_19684,N_19511);
nor U19798 (N_19798,N_19525,N_19551);
xnor U19799 (N_19799,N_19652,N_19536);
xor U19800 (N_19800,N_19588,N_19575);
xor U19801 (N_19801,N_19545,N_19521);
nand U19802 (N_19802,N_19740,N_19534);
nor U19803 (N_19803,N_19676,N_19568);
xor U19804 (N_19804,N_19504,N_19617);
or U19805 (N_19805,N_19533,N_19724);
or U19806 (N_19806,N_19716,N_19742);
xnor U19807 (N_19807,N_19696,N_19714);
nand U19808 (N_19808,N_19667,N_19654);
and U19809 (N_19809,N_19708,N_19730);
and U19810 (N_19810,N_19704,N_19544);
nand U19811 (N_19811,N_19701,N_19690);
nor U19812 (N_19812,N_19627,N_19581);
or U19813 (N_19813,N_19565,N_19639);
or U19814 (N_19814,N_19616,N_19618);
nor U19815 (N_19815,N_19665,N_19736);
and U19816 (N_19816,N_19529,N_19689);
and U19817 (N_19817,N_19526,N_19680);
nand U19818 (N_19818,N_19715,N_19597);
xnor U19819 (N_19819,N_19503,N_19662);
or U19820 (N_19820,N_19541,N_19560);
and U19821 (N_19821,N_19628,N_19610);
and U19822 (N_19822,N_19604,N_19608);
xor U19823 (N_19823,N_19555,N_19589);
and U19824 (N_19824,N_19572,N_19685);
xor U19825 (N_19825,N_19732,N_19634);
nor U19826 (N_19826,N_19666,N_19622);
or U19827 (N_19827,N_19658,N_19743);
nand U19828 (N_19828,N_19682,N_19587);
xnor U19829 (N_19829,N_19599,N_19508);
xnor U19830 (N_19830,N_19671,N_19590);
or U19831 (N_19831,N_19523,N_19711);
nor U19832 (N_19832,N_19647,N_19578);
nand U19833 (N_19833,N_19720,N_19687);
nor U19834 (N_19834,N_19546,N_19600);
and U19835 (N_19835,N_19585,N_19703);
nor U19836 (N_19836,N_19563,N_19636);
and U19837 (N_19837,N_19629,N_19709);
xnor U19838 (N_19838,N_19734,N_19577);
and U19839 (N_19839,N_19518,N_19637);
and U19840 (N_19840,N_19517,N_19557);
nor U19841 (N_19841,N_19645,N_19611);
nor U19842 (N_19842,N_19664,N_19501);
or U19843 (N_19843,N_19558,N_19562);
or U19844 (N_19844,N_19592,N_19624);
and U19845 (N_19845,N_19605,N_19625);
nand U19846 (N_19846,N_19661,N_19706);
and U19847 (N_19847,N_19719,N_19561);
nor U19848 (N_19848,N_19593,N_19612);
or U19849 (N_19849,N_19712,N_19699);
and U19850 (N_19850,N_19522,N_19675);
and U19851 (N_19851,N_19571,N_19519);
nor U19852 (N_19852,N_19535,N_19670);
and U19853 (N_19853,N_19559,N_19669);
or U19854 (N_19854,N_19737,N_19651);
nor U19855 (N_19855,N_19619,N_19646);
nand U19856 (N_19856,N_19603,N_19527);
nand U19857 (N_19857,N_19505,N_19641);
nand U19858 (N_19858,N_19697,N_19528);
xnor U19859 (N_19859,N_19722,N_19681);
or U19860 (N_19860,N_19613,N_19509);
xor U19861 (N_19861,N_19601,N_19556);
nand U19862 (N_19862,N_19649,N_19741);
xnor U19863 (N_19863,N_19542,N_19582);
and U19864 (N_19864,N_19672,N_19512);
xnor U19865 (N_19865,N_19686,N_19626);
nand U19866 (N_19866,N_19717,N_19630);
xnor U19867 (N_19867,N_19591,N_19576);
or U19868 (N_19868,N_19537,N_19540);
and U19869 (N_19869,N_19635,N_19660);
xnor U19870 (N_19870,N_19580,N_19677);
and U19871 (N_19871,N_19695,N_19620);
nor U19872 (N_19872,N_19606,N_19659);
nor U19873 (N_19873,N_19748,N_19594);
and U19874 (N_19874,N_19728,N_19570);
or U19875 (N_19875,N_19709,N_19711);
or U19876 (N_19876,N_19636,N_19664);
xor U19877 (N_19877,N_19564,N_19741);
xor U19878 (N_19878,N_19697,N_19741);
nor U19879 (N_19879,N_19560,N_19573);
xor U19880 (N_19880,N_19695,N_19636);
or U19881 (N_19881,N_19594,N_19583);
and U19882 (N_19882,N_19589,N_19570);
xnor U19883 (N_19883,N_19570,N_19582);
and U19884 (N_19884,N_19501,N_19605);
nand U19885 (N_19885,N_19544,N_19650);
or U19886 (N_19886,N_19641,N_19719);
or U19887 (N_19887,N_19701,N_19681);
and U19888 (N_19888,N_19629,N_19683);
and U19889 (N_19889,N_19695,N_19568);
and U19890 (N_19890,N_19711,N_19562);
or U19891 (N_19891,N_19551,N_19592);
xnor U19892 (N_19892,N_19715,N_19645);
nor U19893 (N_19893,N_19575,N_19672);
nand U19894 (N_19894,N_19705,N_19732);
and U19895 (N_19895,N_19700,N_19626);
and U19896 (N_19896,N_19659,N_19689);
nand U19897 (N_19897,N_19668,N_19506);
nor U19898 (N_19898,N_19554,N_19606);
or U19899 (N_19899,N_19652,N_19524);
nor U19900 (N_19900,N_19681,N_19596);
nor U19901 (N_19901,N_19577,N_19686);
nand U19902 (N_19902,N_19637,N_19560);
nor U19903 (N_19903,N_19625,N_19611);
nand U19904 (N_19904,N_19646,N_19582);
or U19905 (N_19905,N_19528,N_19531);
or U19906 (N_19906,N_19711,N_19648);
or U19907 (N_19907,N_19590,N_19546);
or U19908 (N_19908,N_19556,N_19704);
nand U19909 (N_19909,N_19524,N_19622);
nor U19910 (N_19910,N_19602,N_19607);
xor U19911 (N_19911,N_19736,N_19678);
or U19912 (N_19912,N_19748,N_19600);
nand U19913 (N_19913,N_19688,N_19745);
xor U19914 (N_19914,N_19622,N_19609);
nor U19915 (N_19915,N_19670,N_19594);
nor U19916 (N_19916,N_19674,N_19719);
nand U19917 (N_19917,N_19661,N_19622);
xnor U19918 (N_19918,N_19675,N_19641);
and U19919 (N_19919,N_19686,N_19678);
or U19920 (N_19920,N_19703,N_19614);
nor U19921 (N_19921,N_19584,N_19589);
nand U19922 (N_19922,N_19552,N_19741);
xnor U19923 (N_19923,N_19641,N_19713);
nand U19924 (N_19924,N_19613,N_19532);
nor U19925 (N_19925,N_19701,N_19728);
or U19926 (N_19926,N_19616,N_19682);
nand U19927 (N_19927,N_19632,N_19634);
xnor U19928 (N_19928,N_19699,N_19743);
nand U19929 (N_19929,N_19595,N_19667);
or U19930 (N_19930,N_19658,N_19527);
nor U19931 (N_19931,N_19749,N_19623);
nand U19932 (N_19932,N_19601,N_19533);
xnor U19933 (N_19933,N_19671,N_19691);
or U19934 (N_19934,N_19693,N_19734);
nor U19935 (N_19935,N_19588,N_19540);
xnor U19936 (N_19936,N_19550,N_19549);
or U19937 (N_19937,N_19585,N_19569);
nor U19938 (N_19938,N_19529,N_19570);
xor U19939 (N_19939,N_19733,N_19740);
and U19940 (N_19940,N_19575,N_19718);
nand U19941 (N_19941,N_19539,N_19634);
xnor U19942 (N_19942,N_19563,N_19602);
and U19943 (N_19943,N_19691,N_19579);
nor U19944 (N_19944,N_19745,N_19707);
and U19945 (N_19945,N_19700,N_19584);
xnor U19946 (N_19946,N_19509,N_19500);
and U19947 (N_19947,N_19656,N_19726);
and U19948 (N_19948,N_19632,N_19657);
or U19949 (N_19949,N_19674,N_19594);
nand U19950 (N_19950,N_19511,N_19641);
nor U19951 (N_19951,N_19692,N_19741);
nor U19952 (N_19952,N_19718,N_19647);
nand U19953 (N_19953,N_19747,N_19538);
or U19954 (N_19954,N_19749,N_19740);
nand U19955 (N_19955,N_19683,N_19565);
nor U19956 (N_19956,N_19649,N_19591);
nor U19957 (N_19957,N_19730,N_19585);
nand U19958 (N_19958,N_19583,N_19671);
or U19959 (N_19959,N_19631,N_19724);
xor U19960 (N_19960,N_19703,N_19586);
nor U19961 (N_19961,N_19717,N_19599);
nor U19962 (N_19962,N_19721,N_19643);
xnor U19963 (N_19963,N_19707,N_19724);
nand U19964 (N_19964,N_19738,N_19524);
nand U19965 (N_19965,N_19503,N_19724);
xor U19966 (N_19966,N_19526,N_19707);
nand U19967 (N_19967,N_19576,N_19582);
or U19968 (N_19968,N_19593,N_19661);
nand U19969 (N_19969,N_19660,N_19711);
nand U19970 (N_19970,N_19615,N_19597);
xnor U19971 (N_19971,N_19619,N_19665);
nor U19972 (N_19972,N_19685,N_19583);
and U19973 (N_19973,N_19620,N_19584);
nor U19974 (N_19974,N_19733,N_19635);
nand U19975 (N_19975,N_19610,N_19527);
nand U19976 (N_19976,N_19678,N_19748);
nand U19977 (N_19977,N_19553,N_19526);
nor U19978 (N_19978,N_19653,N_19680);
and U19979 (N_19979,N_19658,N_19735);
xor U19980 (N_19980,N_19650,N_19714);
nand U19981 (N_19981,N_19631,N_19556);
nor U19982 (N_19982,N_19535,N_19641);
and U19983 (N_19983,N_19607,N_19507);
or U19984 (N_19984,N_19693,N_19638);
and U19985 (N_19985,N_19657,N_19577);
xor U19986 (N_19986,N_19662,N_19568);
and U19987 (N_19987,N_19539,N_19706);
and U19988 (N_19988,N_19724,N_19656);
or U19989 (N_19989,N_19559,N_19649);
and U19990 (N_19990,N_19566,N_19738);
and U19991 (N_19991,N_19728,N_19675);
nor U19992 (N_19992,N_19655,N_19601);
xnor U19993 (N_19993,N_19735,N_19715);
nor U19994 (N_19994,N_19716,N_19707);
nand U19995 (N_19995,N_19555,N_19732);
or U19996 (N_19996,N_19717,N_19651);
or U19997 (N_19997,N_19665,N_19500);
and U19998 (N_19998,N_19712,N_19722);
nand U19999 (N_19999,N_19686,N_19580);
nor U20000 (N_20000,N_19992,N_19832);
nand U20001 (N_20001,N_19935,N_19809);
and U20002 (N_20002,N_19818,N_19819);
and U20003 (N_20003,N_19994,N_19954);
nand U20004 (N_20004,N_19790,N_19987);
xor U20005 (N_20005,N_19947,N_19925);
xor U20006 (N_20006,N_19808,N_19958);
nand U20007 (N_20007,N_19858,N_19782);
nand U20008 (N_20008,N_19814,N_19854);
nor U20009 (N_20009,N_19763,N_19861);
nand U20010 (N_20010,N_19974,N_19953);
and U20011 (N_20011,N_19765,N_19866);
nor U20012 (N_20012,N_19914,N_19849);
xnor U20013 (N_20013,N_19929,N_19811);
xnor U20014 (N_20014,N_19901,N_19923);
and U20015 (N_20015,N_19946,N_19840);
nand U20016 (N_20016,N_19951,N_19852);
nand U20017 (N_20017,N_19936,N_19862);
xor U20018 (N_20018,N_19909,N_19783);
nand U20019 (N_20019,N_19781,N_19881);
xor U20020 (N_20020,N_19920,N_19788);
nor U20021 (N_20021,N_19888,N_19896);
and U20022 (N_20022,N_19993,N_19856);
nand U20023 (N_20023,N_19973,N_19848);
nand U20024 (N_20024,N_19807,N_19940);
xnor U20025 (N_20025,N_19759,N_19839);
nor U20026 (N_20026,N_19859,N_19803);
nand U20027 (N_20027,N_19835,N_19756);
nor U20028 (N_20028,N_19800,N_19944);
xnor U20029 (N_20029,N_19916,N_19773);
xor U20030 (N_20030,N_19982,N_19816);
nor U20031 (N_20031,N_19879,N_19830);
and U20032 (N_20032,N_19764,N_19957);
nor U20033 (N_20033,N_19961,N_19778);
and U20034 (N_20034,N_19871,N_19952);
nor U20035 (N_20035,N_19921,N_19963);
xnor U20036 (N_20036,N_19938,N_19757);
nand U20037 (N_20037,N_19980,N_19865);
xor U20038 (N_20038,N_19872,N_19821);
or U20039 (N_20039,N_19959,N_19804);
xnor U20040 (N_20040,N_19823,N_19897);
and U20041 (N_20041,N_19842,N_19949);
nand U20042 (N_20042,N_19898,N_19831);
and U20043 (N_20043,N_19966,N_19813);
and U20044 (N_20044,N_19919,N_19899);
xor U20045 (N_20045,N_19761,N_19900);
xnor U20046 (N_20046,N_19753,N_19884);
or U20047 (N_20047,N_19945,N_19817);
nand U20048 (N_20048,N_19844,N_19754);
or U20049 (N_20049,N_19885,N_19792);
xor U20050 (N_20050,N_19863,N_19990);
or U20051 (N_20051,N_19972,N_19960);
xnor U20052 (N_20052,N_19834,N_19962);
or U20053 (N_20053,N_19853,N_19933);
xnor U20054 (N_20054,N_19796,N_19977);
xor U20055 (N_20055,N_19956,N_19995);
xnor U20056 (N_20056,N_19867,N_19822);
nor U20057 (N_20057,N_19922,N_19902);
xor U20058 (N_20058,N_19981,N_19767);
or U20059 (N_20059,N_19875,N_19786);
nor U20060 (N_20060,N_19912,N_19988);
xor U20061 (N_20061,N_19976,N_19874);
nor U20062 (N_20062,N_19969,N_19941);
and U20063 (N_20063,N_19978,N_19930);
or U20064 (N_20064,N_19843,N_19880);
and U20065 (N_20065,N_19785,N_19774);
or U20066 (N_20066,N_19975,N_19873);
nand U20067 (N_20067,N_19799,N_19998);
xnor U20068 (N_20068,N_19904,N_19762);
or U20069 (N_20069,N_19777,N_19989);
nand U20070 (N_20070,N_19893,N_19924);
or U20071 (N_20071,N_19910,N_19868);
nand U20072 (N_20072,N_19780,N_19894);
and U20073 (N_20073,N_19825,N_19967);
nor U20074 (N_20074,N_19869,N_19760);
nor U20075 (N_20075,N_19776,N_19836);
xor U20076 (N_20076,N_19791,N_19931);
xor U20077 (N_20077,N_19882,N_19928);
nand U20078 (N_20078,N_19911,N_19795);
nand U20079 (N_20079,N_19845,N_19892);
xor U20080 (N_20080,N_19805,N_19878);
nor U20081 (N_20081,N_19768,N_19758);
and U20082 (N_20082,N_19991,N_19846);
xor U20083 (N_20083,N_19769,N_19948);
and U20084 (N_20084,N_19820,N_19779);
or U20085 (N_20085,N_19999,N_19908);
or U20086 (N_20086,N_19794,N_19829);
nor U20087 (N_20087,N_19810,N_19775);
nand U20088 (N_20088,N_19841,N_19971);
and U20089 (N_20089,N_19857,N_19926);
nand U20090 (N_20090,N_19851,N_19891);
nand U20091 (N_20091,N_19877,N_19895);
nor U20092 (N_20092,N_19889,N_19855);
xnor U20093 (N_20093,N_19755,N_19907);
nand U20094 (N_20094,N_19770,N_19824);
or U20095 (N_20095,N_19751,N_19772);
and U20096 (N_20096,N_19997,N_19793);
nand U20097 (N_20097,N_19942,N_19787);
and U20098 (N_20098,N_19985,N_19905);
and U20099 (N_20099,N_19932,N_19965);
nor U20100 (N_20100,N_19801,N_19939);
or U20101 (N_20101,N_19752,N_19860);
nand U20102 (N_20102,N_19847,N_19937);
xor U20103 (N_20103,N_19955,N_19915);
nor U20104 (N_20104,N_19886,N_19917);
and U20105 (N_20105,N_19964,N_19979);
or U20106 (N_20106,N_19890,N_19918);
and U20107 (N_20107,N_19797,N_19986);
and U20108 (N_20108,N_19903,N_19789);
or U20109 (N_20109,N_19850,N_19750);
nor U20110 (N_20110,N_19883,N_19802);
or U20111 (N_20111,N_19815,N_19784);
and U20112 (N_20112,N_19876,N_19887);
or U20113 (N_20113,N_19798,N_19826);
and U20114 (N_20114,N_19864,N_19983);
nand U20115 (N_20115,N_19766,N_19968);
nand U20116 (N_20116,N_19870,N_19934);
nor U20117 (N_20117,N_19827,N_19837);
nor U20118 (N_20118,N_19950,N_19833);
xor U20119 (N_20119,N_19984,N_19812);
or U20120 (N_20120,N_19771,N_19806);
nand U20121 (N_20121,N_19943,N_19996);
and U20122 (N_20122,N_19828,N_19906);
nor U20123 (N_20123,N_19970,N_19913);
or U20124 (N_20124,N_19838,N_19927);
nand U20125 (N_20125,N_19957,N_19914);
nor U20126 (N_20126,N_19781,N_19846);
nand U20127 (N_20127,N_19890,N_19954);
nand U20128 (N_20128,N_19793,N_19764);
and U20129 (N_20129,N_19978,N_19970);
and U20130 (N_20130,N_19963,N_19813);
and U20131 (N_20131,N_19952,N_19966);
or U20132 (N_20132,N_19784,N_19962);
and U20133 (N_20133,N_19823,N_19830);
and U20134 (N_20134,N_19818,N_19850);
xor U20135 (N_20135,N_19802,N_19808);
xnor U20136 (N_20136,N_19824,N_19887);
nand U20137 (N_20137,N_19763,N_19939);
nor U20138 (N_20138,N_19777,N_19978);
xor U20139 (N_20139,N_19965,N_19896);
xor U20140 (N_20140,N_19959,N_19983);
or U20141 (N_20141,N_19897,N_19913);
and U20142 (N_20142,N_19964,N_19977);
or U20143 (N_20143,N_19811,N_19884);
nand U20144 (N_20144,N_19791,N_19778);
and U20145 (N_20145,N_19873,N_19987);
nand U20146 (N_20146,N_19818,N_19909);
nor U20147 (N_20147,N_19811,N_19824);
nor U20148 (N_20148,N_19860,N_19791);
nor U20149 (N_20149,N_19780,N_19945);
nand U20150 (N_20150,N_19815,N_19845);
or U20151 (N_20151,N_19845,N_19856);
xor U20152 (N_20152,N_19953,N_19753);
nand U20153 (N_20153,N_19981,N_19859);
or U20154 (N_20154,N_19878,N_19957);
or U20155 (N_20155,N_19991,N_19882);
nand U20156 (N_20156,N_19980,N_19809);
and U20157 (N_20157,N_19963,N_19843);
and U20158 (N_20158,N_19901,N_19910);
nor U20159 (N_20159,N_19810,N_19895);
xor U20160 (N_20160,N_19797,N_19961);
nand U20161 (N_20161,N_19832,N_19775);
and U20162 (N_20162,N_19870,N_19996);
nor U20163 (N_20163,N_19780,N_19913);
xnor U20164 (N_20164,N_19941,N_19842);
nor U20165 (N_20165,N_19824,N_19763);
or U20166 (N_20166,N_19947,N_19933);
and U20167 (N_20167,N_19868,N_19882);
and U20168 (N_20168,N_19923,N_19806);
xnor U20169 (N_20169,N_19802,N_19825);
and U20170 (N_20170,N_19911,N_19948);
xor U20171 (N_20171,N_19885,N_19804);
or U20172 (N_20172,N_19752,N_19818);
xnor U20173 (N_20173,N_19766,N_19806);
nand U20174 (N_20174,N_19814,N_19810);
or U20175 (N_20175,N_19835,N_19952);
nand U20176 (N_20176,N_19863,N_19799);
xor U20177 (N_20177,N_19845,N_19894);
nor U20178 (N_20178,N_19820,N_19913);
xnor U20179 (N_20179,N_19874,N_19865);
nor U20180 (N_20180,N_19892,N_19959);
nand U20181 (N_20181,N_19996,N_19966);
and U20182 (N_20182,N_19988,N_19822);
nor U20183 (N_20183,N_19948,N_19897);
or U20184 (N_20184,N_19888,N_19782);
nand U20185 (N_20185,N_19968,N_19830);
and U20186 (N_20186,N_19983,N_19951);
nand U20187 (N_20187,N_19967,N_19803);
nor U20188 (N_20188,N_19979,N_19807);
and U20189 (N_20189,N_19754,N_19982);
xnor U20190 (N_20190,N_19790,N_19766);
and U20191 (N_20191,N_19951,N_19944);
and U20192 (N_20192,N_19812,N_19935);
or U20193 (N_20193,N_19934,N_19941);
nor U20194 (N_20194,N_19978,N_19986);
or U20195 (N_20195,N_19874,N_19921);
nor U20196 (N_20196,N_19750,N_19964);
nor U20197 (N_20197,N_19765,N_19862);
or U20198 (N_20198,N_19880,N_19874);
and U20199 (N_20199,N_19996,N_19942);
or U20200 (N_20200,N_19919,N_19902);
xor U20201 (N_20201,N_19903,N_19887);
xnor U20202 (N_20202,N_19898,N_19932);
nor U20203 (N_20203,N_19972,N_19922);
and U20204 (N_20204,N_19783,N_19763);
or U20205 (N_20205,N_19856,N_19818);
and U20206 (N_20206,N_19852,N_19980);
and U20207 (N_20207,N_19928,N_19765);
or U20208 (N_20208,N_19776,N_19824);
nor U20209 (N_20209,N_19915,N_19788);
or U20210 (N_20210,N_19916,N_19879);
nor U20211 (N_20211,N_19793,N_19944);
nand U20212 (N_20212,N_19796,N_19946);
nand U20213 (N_20213,N_19856,N_19812);
xor U20214 (N_20214,N_19836,N_19934);
and U20215 (N_20215,N_19770,N_19774);
nand U20216 (N_20216,N_19891,N_19903);
nand U20217 (N_20217,N_19783,N_19836);
or U20218 (N_20218,N_19972,N_19763);
nor U20219 (N_20219,N_19794,N_19776);
xnor U20220 (N_20220,N_19997,N_19750);
nand U20221 (N_20221,N_19952,N_19817);
nor U20222 (N_20222,N_19788,N_19842);
and U20223 (N_20223,N_19786,N_19802);
and U20224 (N_20224,N_19761,N_19972);
nand U20225 (N_20225,N_19877,N_19813);
xor U20226 (N_20226,N_19803,N_19993);
xnor U20227 (N_20227,N_19938,N_19933);
nor U20228 (N_20228,N_19885,N_19939);
nor U20229 (N_20229,N_19898,N_19883);
and U20230 (N_20230,N_19851,N_19900);
nand U20231 (N_20231,N_19814,N_19834);
or U20232 (N_20232,N_19902,N_19874);
or U20233 (N_20233,N_19865,N_19955);
nand U20234 (N_20234,N_19763,N_19765);
xnor U20235 (N_20235,N_19954,N_19891);
or U20236 (N_20236,N_19959,N_19924);
and U20237 (N_20237,N_19802,N_19971);
and U20238 (N_20238,N_19759,N_19863);
nand U20239 (N_20239,N_19958,N_19863);
xor U20240 (N_20240,N_19921,N_19995);
and U20241 (N_20241,N_19777,N_19990);
and U20242 (N_20242,N_19870,N_19965);
nand U20243 (N_20243,N_19799,N_19964);
xor U20244 (N_20244,N_19975,N_19945);
or U20245 (N_20245,N_19955,N_19845);
and U20246 (N_20246,N_19919,N_19888);
xnor U20247 (N_20247,N_19899,N_19813);
nor U20248 (N_20248,N_19854,N_19864);
and U20249 (N_20249,N_19948,N_19949);
xnor U20250 (N_20250,N_20087,N_20101);
or U20251 (N_20251,N_20009,N_20155);
nand U20252 (N_20252,N_20083,N_20195);
xnor U20253 (N_20253,N_20134,N_20158);
or U20254 (N_20254,N_20175,N_20036);
and U20255 (N_20255,N_20047,N_20072);
nor U20256 (N_20256,N_20160,N_20075);
xnor U20257 (N_20257,N_20128,N_20200);
or U20258 (N_20258,N_20177,N_20066);
and U20259 (N_20259,N_20068,N_20185);
nor U20260 (N_20260,N_20076,N_20226);
nand U20261 (N_20261,N_20123,N_20245);
or U20262 (N_20262,N_20034,N_20107);
nand U20263 (N_20263,N_20204,N_20153);
and U20264 (N_20264,N_20082,N_20190);
or U20265 (N_20265,N_20090,N_20224);
nand U20266 (N_20266,N_20148,N_20205);
xor U20267 (N_20267,N_20130,N_20162);
nand U20268 (N_20268,N_20100,N_20013);
and U20269 (N_20269,N_20057,N_20040);
or U20270 (N_20270,N_20117,N_20042);
nand U20271 (N_20271,N_20038,N_20219);
nand U20272 (N_20272,N_20095,N_20064);
or U20273 (N_20273,N_20105,N_20189);
nor U20274 (N_20274,N_20112,N_20070);
and U20275 (N_20275,N_20007,N_20132);
nand U20276 (N_20276,N_20097,N_20152);
and U20277 (N_20277,N_20126,N_20184);
nor U20278 (N_20278,N_20046,N_20212);
and U20279 (N_20279,N_20137,N_20079);
or U20280 (N_20280,N_20139,N_20240);
and U20281 (N_20281,N_20147,N_20161);
xnor U20282 (N_20282,N_20154,N_20116);
xnor U20283 (N_20283,N_20136,N_20193);
xnor U20284 (N_20284,N_20170,N_20058);
and U20285 (N_20285,N_20209,N_20001);
xor U20286 (N_20286,N_20182,N_20180);
nor U20287 (N_20287,N_20196,N_20056);
or U20288 (N_20288,N_20230,N_20019);
xnor U20289 (N_20289,N_20225,N_20027);
and U20290 (N_20290,N_20241,N_20074);
nor U20291 (N_20291,N_20071,N_20033);
and U20292 (N_20292,N_20016,N_20211);
and U20293 (N_20293,N_20227,N_20198);
nor U20294 (N_20294,N_20050,N_20014);
nor U20295 (N_20295,N_20081,N_20049);
and U20296 (N_20296,N_20005,N_20021);
or U20297 (N_20297,N_20096,N_20231);
and U20298 (N_20298,N_20249,N_20186);
and U20299 (N_20299,N_20243,N_20088);
or U20300 (N_20300,N_20141,N_20133);
or U20301 (N_20301,N_20104,N_20159);
xor U20302 (N_20302,N_20004,N_20118);
or U20303 (N_20303,N_20106,N_20089);
nor U20304 (N_20304,N_20120,N_20208);
nor U20305 (N_20305,N_20086,N_20093);
and U20306 (N_20306,N_20011,N_20142);
nor U20307 (N_20307,N_20213,N_20145);
nand U20308 (N_20308,N_20063,N_20197);
nand U20309 (N_20309,N_20122,N_20229);
nand U20310 (N_20310,N_20077,N_20163);
xor U20311 (N_20311,N_20173,N_20022);
or U20312 (N_20312,N_20085,N_20178);
nor U20313 (N_20313,N_20234,N_20191);
xor U20314 (N_20314,N_20171,N_20084);
nand U20315 (N_20315,N_20062,N_20210);
or U20316 (N_20316,N_20244,N_20055);
xnor U20317 (N_20317,N_20149,N_20179);
nand U20318 (N_20318,N_20032,N_20232);
xor U20319 (N_20319,N_20166,N_20156);
and U20320 (N_20320,N_20024,N_20098);
nand U20321 (N_20321,N_20157,N_20165);
nand U20322 (N_20322,N_20129,N_20018);
or U20323 (N_20323,N_20080,N_20172);
nor U20324 (N_20324,N_20168,N_20201);
nor U20325 (N_20325,N_20143,N_20039);
or U20326 (N_20326,N_20020,N_20236);
nor U20327 (N_20327,N_20037,N_20217);
nor U20328 (N_20328,N_20115,N_20125);
nand U20329 (N_20329,N_20203,N_20073);
and U20330 (N_20330,N_20167,N_20029);
or U20331 (N_20331,N_20248,N_20150);
and U20332 (N_20332,N_20099,N_20017);
xnor U20333 (N_20333,N_20221,N_20003);
xor U20334 (N_20334,N_20113,N_20215);
nor U20335 (N_20335,N_20035,N_20242);
nor U20336 (N_20336,N_20045,N_20131);
and U20337 (N_20337,N_20008,N_20054);
xnor U20338 (N_20338,N_20078,N_20164);
xor U20339 (N_20339,N_20060,N_20048);
nor U20340 (N_20340,N_20119,N_20102);
nor U20341 (N_20341,N_20041,N_20202);
nor U20342 (N_20342,N_20114,N_20238);
nor U20343 (N_20343,N_20187,N_20124);
nand U20344 (N_20344,N_20065,N_20044);
xor U20345 (N_20345,N_20103,N_20006);
xnor U20346 (N_20346,N_20194,N_20218);
nor U20347 (N_20347,N_20146,N_20207);
or U20348 (N_20348,N_20181,N_20092);
or U20349 (N_20349,N_20010,N_20214);
or U20350 (N_20350,N_20091,N_20059);
xnor U20351 (N_20351,N_20199,N_20144);
xnor U20352 (N_20352,N_20216,N_20176);
or U20353 (N_20353,N_20015,N_20028);
or U20354 (N_20354,N_20043,N_20069);
and U20355 (N_20355,N_20192,N_20109);
or U20356 (N_20356,N_20222,N_20228);
xnor U20357 (N_20357,N_20206,N_20026);
nand U20358 (N_20358,N_20110,N_20247);
and U20359 (N_20359,N_20140,N_20220);
and U20360 (N_20360,N_20061,N_20000);
and U20361 (N_20361,N_20094,N_20067);
nand U20362 (N_20362,N_20030,N_20051);
xor U20363 (N_20363,N_20239,N_20121);
or U20364 (N_20364,N_20246,N_20183);
or U20365 (N_20365,N_20235,N_20188);
xor U20366 (N_20366,N_20237,N_20053);
xnor U20367 (N_20367,N_20031,N_20138);
and U20368 (N_20368,N_20012,N_20111);
or U20369 (N_20369,N_20169,N_20127);
and U20370 (N_20370,N_20025,N_20052);
nand U20371 (N_20371,N_20108,N_20233);
and U20372 (N_20372,N_20151,N_20135);
nor U20373 (N_20373,N_20174,N_20002);
nand U20374 (N_20374,N_20223,N_20023);
nor U20375 (N_20375,N_20123,N_20191);
nand U20376 (N_20376,N_20097,N_20085);
or U20377 (N_20377,N_20186,N_20141);
or U20378 (N_20378,N_20084,N_20242);
nand U20379 (N_20379,N_20220,N_20139);
or U20380 (N_20380,N_20204,N_20083);
nor U20381 (N_20381,N_20032,N_20054);
and U20382 (N_20382,N_20020,N_20029);
xnor U20383 (N_20383,N_20064,N_20242);
or U20384 (N_20384,N_20185,N_20214);
nor U20385 (N_20385,N_20141,N_20044);
nor U20386 (N_20386,N_20165,N_20065);
and U20387 (N_20387,N_20088,N_20063);
nor U20388 (N_20388,N_20234,N_20150);
xnor U20389 (N_20389,N_20199,N_20196);
and U20390 (N_20390,N_20117,N_20115);
nand U20391 (N_20391,N_20123,N_20132);
nand U20392 (N_20392,N_20008,N_20231);
nand U20393 (N_20393,N_20123,N_20084);
or U20394 (N_20394,N_20192,N_20055);
nand U20395 (N_20395,N_20218,N_20147);
nand U20396 (N_20396,N_20242,N_20096);
xor U20397 (N_20397,N_20159,N_20105);
nand U20398 (N_20398,N_20200,N_20015);
or U20399 (N_20399,N_20099,N_20210);
xor U20400 (N_20400,N_20175,N_20071);
xor U20401 (N_20401,N_20050,N_20144);
or U20402 (N_20402,N_20132,N_20231);
nor U20403 (N_20403,N_20218,N_20052);
or U20404 (N_20404,N_20236,N_20035);
xor U20405 (N_20405,N_20044,N_20221);
nand U20406 (N_20406,N_20109,N_20228);
or U20407 (N_20407,N_20129,N_20189);
nor U20408 (N_20408,N_20094,N_20111);
nor U20409 (N_20409,N_20007,N_20030);
xnor U20410 (N_20410,N_20000,N_20249);
or U20411 (N_20411,N_20133,N_20106);
and U20412 (N_20412,N_20125,N_20189);
or U20413 (N_20413,N_20040,N_20113);
and U20414 (N_20414,N_20055,N_20141);
and U20415 (N_20415,N_20196,N_20173);
or U20416 (N_20416,N_20135,N_20051);
nand U20417 (N_20417,N_20211,N_20219);
xnor U20418 (N_20418,N_20212,N_20037);
and U20419 (N_20419,N_20127,N_20059);
and U20420 (N_20420,N_20175,N_20170);
nand U20421 (N_20421,N_20212,N_20068);
nand U20422 (N_20422,N_20166,N_20072);
and U20423 (N_20423,N_20235,N_20071);
or U20424 (N_20424,N_20086,N_20092);
nor U20425 (N_20425,N_20166,N_20076);
xnor U20426 (N_20426,N_20233,N_20215);
or U20427 (N_20427,N_20083,N_20011);
and U20428 (N_20428,N_20232,N_20084);
or U20429 (N_20429,N_20118,N_20001);
xnor U20430 (N_20430,N_20176,N_20248);
xnor U20431 (N_20431,N_20030,N_20125);
nor U20432 (N_20432,N_20010,N_20136);
nand U20433 (N_20433,N_20184,N_20110);
or U20434 (N_20434,N_20198,N_20115);
xnor U20435 (N_20435,N_20113,N_20055);
nor U20436 (N_20436,N_20014,N_20002);
xor U20437 (N_20437,N_20021,N_20228);
and U20438 (N_20438,N_20113,N_20212);
or U20439 (N_20439,N_20036,N_20078);
nor U20440 (N_20440,N_20182,N_20029);
nand U20441 (N_20441,N_20237,N_20008);
and U20442 (N_20442,N_20214,N_20144);
or U20443 (N_20443,N_20207,N_20067);
xnor U20444 (N_20444,N_20119,N_20067);
xor U20445 (N_20445,N_20097,N_20019);
xnor U20446 (N_20446,N_20011,N_20028);
and U20447 (N_20447,N_20028,N_20208);
or U20448 (N_20448,N_20120,N_20019);
xor U20449 (N_20449,N_20214,N_20212);
nand U20450 (N_20450,N_20199,N_20011);
nand U20451 (N_20451,N_20048,N_20122);
or U20452 (N_20452,N_20037,N_20210);
and U20453 (N_20453,N_20223,N_20122);
nand U20454 (N_20454,N_20198,N_20034);
and U20455 (N_20455,N_20092,N_20195);
nor U20456 (N_20456,N_20115,N_20047);
nand U20457 (N_20457,N_20151,N_20016);
nor U20458 (N_20458,N_20137,N_20031);
and U20459 (N_20459,N_20099,N_20192);
nor U20460 (N_20460,N_20126,N_20225);
and U20461 (N_20461,N_20143,N_20042);
or U20462 (N_20462,N_20090,N_20245);
nand U20463 (N_20463,N_20126,N_20092);
and U20464 (N_20464,N_20184,N_20041);
or U20465 (N_20465,N_20115,N_20053);
nand U20466 (N_20466,N_20198,N_20183);
nand U20467 (N_20467,N_20089,N_20124);
and U20468 (N_20468,N_20026,N_20154);
xnor U20469 (N_20469,N_20033,N_20131);
or U20470 (N_20470,N_20161,N_20016);
nor U20471 (N_20471,N_20181,N_20031);
nand U20472 (N_20472,N_20143,N_20095);
nand U20473 (N_20473,N_20004,N_20128);
and U20474 (N_20474,N_20213,N_20200);
nand U20475 (N_20475,N_20032,N_20196);
and U20476 (N_20476,N_20057,N_20071);
and U20477 (N_20477,N_20045,N_20184);
and U20478 (N_20478,N_20116,N_20048);
nor U20479 (N_20479,N_20012,N_20039);
xnor U20480 (N_20480,N_20214,N_20033);
nand U20481 (N_20481,N_20239,N_20180);
and U20482 (N_20482,N_20236,N_20090);
and U20483 (N_20483,N_20124,N_20228);
or U20484 (N_20484,N_20078,N_20163);
nor U20485 (N_20485,N_20093,N_20122);
nor U20486 (N_20486,N_20130,N_20038);
or U20487 (N_20487,N_20026,N_20008);
nor U20488 (N_20488,N_20204,N_20070);
nand U20489 (N_20489,N_20199,N_20013);
or U20490 (N_20490,N_20004,N_20235);
and U20491 (N_20491,N_20247,N_20020);
nor U20492 (N_20492,N_20150,N_20158);
nor U20493 (N_20493,N_20030,N_20048);
nor U20494 (N_20494,N_20093,N_20230);
and U20495 (N_20495,N_20019,N_20076);
and U20496 (N_20496,N_20140,N_20000);
nand U20497 (N_20497,N_20092,N_20065);
nand U20498 (N_20498,N_20089,N_20054);
xnor U20499 (N_20499,N_20160,N_20085);
and U20500 (N_20500,N_20250,N_20260);
nand U20501 (N_20501,N_20428,N_20296);
nand U20502 (N_20502,N_20413,N_20419);
xnor U20503 (N_20503,N_20418,N_20326);
and U20504 (N_20504,N_20344,N_20405);
xnor U20505 (N_20505,N_20416,N_20396);
nand U20506 (N_20506,N_20410,N_20374);
nor U20507 (N_20507,N_20261,N_20437);
nor U20508 (N_20508,N_20290,N_20475);
and U20509 (N_20509,N_20337,N_20403);
nand U20510 (N_20510,N_20318,N_20451);
or U20511 (N_20511,N_20336,N_20386);
nor U20512 (N_20512,N_20355,N_20455);
nand U20513 (N_20513,N_20469,N_20332);
nor U20514 (N_20514,N_20280,N_20390);
xnor U20515 (N_20515,N_20361,N_20466);
nor U20516 (N_20516,N_20442,N_20480);
xnor U20517 (N_20517,N_20368,N_20497);
or U20518 (N_20518,N_20422,N_20474);
nor U20519 (N_20519,N_20458,N_20383);
nand U20520 (N_20520,N_20335,N_20263);
xor U20521 (N_20521,N_20459,N_20317);
nand U20522 (N_20522,N_20482,N_20493);
nand U20523 (N_20523,N_20434,N_20283);
nor U20524 (N_20524,N_20421,N_20301);
nor U20525 (N_20525,N_20393,N_20481);
xor U20526 (N_20526,N_20346,N_20484);
nor U20527 (N_20527,N_20398,N_20495);
nor U20528 (N_20528,N_20476,N_20275);
xnor U20529 (N_20529,N_20401,N_20310);
nand U20530 (N_20530,N_20464,N_20488);
xor U20531 (N_20531,N_20454,N_20328);
nand U20532 (N_20532,N_20417,N_20358);
xor U20533 (N_20533,N_20343,N_20460);
xor U20534 (N_20534,N_20307,N_20256);
and U20535 (N_20535,N_20433,N_20281);
or U20536 (N_20536,N_20457,N_20440);
nor U20537 (N_20537,N_20364,N_20266);
xor U20538 (N_20538,N_20282,N_20376);
nand U20539 (N_20539,N_20435,N_20365);
and U20540 (N_20540,N_20298,N_20424);
nor U20541 (N_20541,N_20449,N_20342);
xnor U20542 (N_20542,N_20378,N_20492);
or U20543 (N_20543,N_20253,N_20322);
and U20544 (N_20544,N_20465,N_20441);
nor U20545 (N_20545,N_20363,N_20284);
and U20546 (N_20546,N_20353,N_20498);
or U20547 (N_20547,N_20494,N_20379);
xnor U20548 (N_20548,N_20409,N_20399);
nand U20549 (N_20549,N_20375,N_20425);
and U20550 (N_20550,N_20321,N_20427);
nor U20551 (N_20551,N_20436,N_20351);
or U20552 (N_20552,N_20339,N_20496);
and U20553 (N_20553,N_20392,N_20308);
nand U20554 (N_20554,N_20473,N_20395);
nor U20555 (N_20555,N_20381,N_20499);
nand U20556 (N_20556,N_20286,N_20265);
and U20557 (N_20557,N_20311,N_20309);
or U20558 (N_20558,N_20432,N_20268);
and U20559 (N_20559,N_20412,N_20408);
nand U20560 (N_20560,N_20297,N_20288);
nor U20561 (N_20561,N_20420,N_20354);
nand U20562 (N_20562,N_20370,N_20262);
nand U20563 (N_20563,N_20414,N_20255);
nor U20564 (N_20564,N_20330,N_20439);
xor U20565 (N_20565,N_20257,N_20316);
nand U20566 (N_20566,N_20490,N_20264);
and U20567 (N_20567,N_20485,N_20293);
nor U20568 (N_20568,N_20299,N_20470);
xnor U20569 (N_20569,N_20334,N_20415);
xnor U20570 (N_20570,N_20357,N_20340);
xor U20571 (N_20571,N_20315,N_20366);
xnor U20572 (N_20572,N_20446,N_20259);
nand U20573 (N_20573,N_20388,N_20306);
or U20574 (N_20574,N_20252,N_20452);
or U20575 (N_20575,N_20373,N_20267);
nor U20576 (N_20576,N_20302,N_20274);
nor U20577 (N_20577,N_20312,N_20347);
nand U20578 (N_20578,N_20430,N_20448);
or U20579 (N_20579,N_20367,N_20269);
or U20580 (N_20580,N_20305,N_20477);
xnor U20581 (N_20581,N_20423,N_20345);
and U20582 (N_20582,N_20277,N_20380);
xnor U20583 (N_20583,N_20327,N_20384);
or U20584 (N_20584,N_20478,N_20483);
nor U20585 (N_20585,N_20443,N_20276);
nand U20586 (N_20586,N_20352,N_20377);
xor U20587 (N_20587,N_20406,N_20272);
nor U20588 (N_20588,N_20397,N_20453);
nand U20589 (N_20589,N_20292,N_20479);
nor U20590 (N_20590,N_20356,N_20426);
nand U20591 (N_20591,N_20438,N_20341);
or U20592 (N_20592,N_20411,N_20404);
nand U20593 (N_20593,N_20314,N_20407);
or U20594 (N_20594,N_20391,N_20319);
or U20595 (N_20595,N_20444,N_20456);
or U20596 (N_20596,N_20278,N_20271);
and U20597 (N_20597,N_20402,N_20303);
nand U20598 (N_20598,N_20313,N_20348);
or U20599 (N_20599,N_20279,N_20333);
nor U20600 (N_20600,N_20285,N_20323);
xnor U20601 (N_20601,N_20394,N_20350);
nand U20602 (N_20602,N_20371,N_20304);
or U20603 (N_20603,N_20382,N_20331);
or U20604 (N_20604,N_20287,N_20289);
xor U20605 (N_20605,N_20360,N_20429);
xor U20606 (N_20606,N_20389,N_20320);
or U20607 (N_20607,N_20295,N_20273);
and U20608 (N_20608,N_20491,N_20461);
or U20609 (N_20609,N_20254,N_20251);
nand U20610 (N_20610,N_20372,N_20359);
xnor U20611 (N_20611,N_20431,N_20468);
nand U20612 (N_20612,N_20487,N_20463);
nor U20613 (N_20613,N_20291,N_20369);
nor U20614 (N_20614,N_20400,N_20467);
and U20615 (N_20615,N_20489,N_20447);
nand U20616 (N_20616,N_20300,N_20324);
nor U20617 (N_20617,N_20258,N_20472);
nor U20618 (N_20618,N_20387,N_20338);
nor U20619 (N_20619,N_20294,N_20270);
nand U20620 (N_20620,N_20362,N_20349);
xor U20621 (N_20621,N_20471,N_20486);
nand U20622 (N_20622,N_20462,N_20385);
xor U20623 (N_20623,N_20329,N_20450);
and U20624 (N_20624,N_20325,N_20445);
nand U20625 (N_20625,N_20358,N_20287);
xnor U20626 (N_20626,N_20297,N_20284);
xnor U20627 (N_20627,N_20264,N_20402);
nor U20628 (N_20628,N_20484,N_20343);
and U20629 (N_20629,N_20332,N_20300);
xnor U20630 (N_20630,N_20372,N_20255);
xor U20631 (N_20631,N_20422,N_20392);
or U20632 (N_20632,N_20348,N_20468);
nand U20633 (N_20633,N_20441,N_20387);
or U20634 (N_20634,N_20261,N_20481);
nor U20635 (N_20635,N_20360,N_20333);
or U20636 (N_20636,N_20436,N_20280);
nand U20637 (N_20637,N_20418,N_20425);
nor U20638 (N_20638,N_20291,N_20474);
xor U20639 (N_20639,N_20488,N_20268);
and U20640 (N_20640,N_20384,N_20443);
nand U20641 (N_20641,N_20331,N_20290);
nor U20642 (N_20642,N_20494,N_20374);
and U20643 (N_20643,N_20371,N_20391);
nand U20644 (N_20644,N_20467,N_20361);
nor U20645 (N_20645,N_20457,N_20479);
nand U20646 (N_20646,N_20437,N_20409);
and U20647 (N_20647,N_20358,N_20298);
or U20648 (N_20648,N_20419,N_20357);
or U20649 (N_20649,N_20319,N_20406);
xor U20650 (N_20650,N_20465,N_20447);
and U20651 (N_20651,N_20309,N_20438);
and U20652 (N_20652,N_20410,N_20335);
nor U20653 (N_20653,N_20393,N_20352);
or U20654 (N_20654,N_20299,N_20487);
or U20655 (N_20655,N_20404,N_20418);
or U20656 (N_20656,N_20351,N_20374);
nand U20657 (N_20657,N_20342,N_20423);
xnor U20658 (N_20658,N_20468,N_20420);
xnor U20659 (N_20659,N_20481,N_20262);
and U20660 (N_20660,N_20437,N_20479);
nand U20661 (N_20661,N_20445,N_20336);
nand U20662 (N_20662,N_20279,N_20261);
and U20663 (N_20663,N_20384,N_20440);
xnor U20664 (N_20664,N_20292,N_20361);
or U20665 (N_20665,N_20270,N_20481);
and U20666 (N_20666,N_20311,N_20344);
nor U20667 (N_20667,N_20467,N_20265);
or U20668 (N_20668,N_20391,N_20479);
and U20669 (N_20669,N_20362,N_20320);
xnor U20670 (N_20670,N_20435,N_20284);
nor U20671 (N_20671,N_20285,N_20456);
and U20672 (N_20672,N_20334,N_20433);
and U20673 (N_20673,N_20430,N_20297);
or U20674 (N_20674,N_20476,N_20383);
nand U20675 (N_20675,N_20495,N_20466);
nor U20676 (N_20676,N_20468,N_20294);
nand U20677 (N_20677,N_20352,N_20397);
nand U20678 (N_20678,N_20408,N_20488);
nand U20679 (N_20679,N_20261,N_20336);
nand U20680 (N_20680,N_20270,N_20307);
or U20681 (N_20681,N_20444,N_20275);
and U20682 (N_20682,N_20262,N_20464);
nand U20683 (N_20683,N_20419,N_20327);
or U20684 (N_20684,N_20346,N_20493);
xnor U20685 (N_20685,N_20313,N_20331);
and U20686 (N_20686,N_20321,N_20399);
nand U20687 (N_20687,N_20416,N_20471);
nand U20688 (N_20688,N_20367,N_20298);
xnor U20689 (N_20689,N_20430,N_20488);
xor U20690 (N_20690,N_20450,N_20268);
xnor U20691 (N_20691,N_20303,N_20283);
nor U20692 (N_20692,N_20498,N_20373);
and U20693 (N_20693,N_20291,N_20421);
nor U20694 (N_20694,N_20396,N_20376);
and U20695 (N_20695,N_20264,N_20435);
nor U20696 (N_20696,N_20369,N_20266);
or U20697 (N_20697,N_20474,N_20373);
and U20698 (N_20698,N_20330,N_20296);
or U20699 (N_20699,N_20413,N_20274);
or U20700 (N_20700,N_20453,N_20465);
and U20701 (N_20701,N_20315,N_20424);
nor U20702 (N_20702,N_20386,N_20293);
nand U20703 (N_20703,N_20303,N_20358);
and U20704 (N_20704,N_20394,N_20286);
nor U20705 (N_20705,N_20364,N_20455);
nor U20706 (N_20706,N_20495,N_20346);
nand U20707 (N_20707,N_20462,N_20489);
or U20708 (N_20708,N_20264,N_20358);
nand U20709 (N_20709,N_20448,N_20415);
and U20710 (N_20710,N_20266,N_20296);
nand U20711 (N_20711,N_20479,N_20443);
xor U20712 (N_20712,N_20370,N_20329);
nand U20713 (N_20713,N_20472,N_20493);
nor U20714 (N_20714,N_20318,N_20443);
and U20715 (N_20715,N_20281,N_20257);
and U20716 (N_20716,N_20338,N_20407);
xnor U20717 (N_20717,N_20313,N_20310);
nand U20718 (N_20718,N_20321,N_20302);
nor U20719 (N_20719,N_20489,N_20283);
nor U20720 (N_20720,N_20297,N_20427);
or U20721 (N_20721,N_20452,N_20337);
xor U20722 (N_20722,N_20436,N_20338);
nand U20723 (N_20723,N_20426,N_20306);
and U20724 (N_20724,N_20410,N_20334);
nor U20725 (N_20725,N_20435,N_20314);
nand U20726 (N_20726,N_20327,N_20255);
or U20727 (N_20727,N_20438,N_20254);
xor U20728 (N_20728,N_20390,N_20410);
nand U20729 (N_20729,N_20357,N_20345);
and U20730 (N_20730,N_20309,N_20360);
and U20731 (N_20731,N_20284,N_20285);
or U20732 (N_20732,N_20330,N_20438);
xnor U20733 (N_20733,N_20384,N_20424);
nor U20734 (N_20734,N_20498,N_20400);
nor U20735 (N_20735,N_20316,N_20458);
nand U20736 (N_20736,N_20336,N_20347);
xnor U20737 (N_20737,N_20326,N_20336);
or U20738 (N_20738,N_20311,N_20347);
and U20739 (N_20739,N_20480,N_20435);
or U20740 (N_20740,N_20418,N_20262);
and U20741 (N_20741,N_20285,N_20480);
nor U20742 (N_20742,N_20433,N_20303);
nand U20743 (N_20743,N_20277,N_20431);
nor U20744 (N_20744,N_20322,N_20277);
and U20745 (N_20745,N_20467,N_20488);
nor U20746 (N_20746,N_20322,N_20252);
xor U20747 (N_20747,N_20251,N_20448);
nand U20748 (N_20748,N_20440,N_20408);
xor U20749 (N_20749,N_20433,N_20390);
and U20750 (N_20750,N_20682,N_20571);
or U20751 (N_20751,N_20554,N_20616);
nand U20752 (N_20752,N_20655,N_20702);
or U20753 (N_20753,N_20584,N_20660);
xor U20754 (N_20754,N_20629,N_20569);
and U20755 (N_20755,N_20739,N_20520);
nand U20756 (N_20756,N_20568,N_20661);
xor U20757 (N_20757,N_20555,N_20592);
nor U20758 (N_20758,N_20550,N_20650);
or U20759 (N_20759,N_20526,N_20675);
nor U20760 (N_20760,N_20551,N_20595);
nand U20761 (N_20761,N_20743,N_20689);
nand U20762 (N_20762,N_20742,N_20634);
nor U20763 (N_20763,N_20536,N_20722);
and U20764 (N_20764,N_20604,N_20620);
or U20765 (N_20765,N_20715,N_20635);
nor U20766 (N_20766,N_20600,N_20706);
nand U20767 (N_20767,N_20736,N_20602);
or U20768 (N_20768,N_20601,N_20565);
nand U20769 (N_20769,N_20587,N_20656);
nor U20770 (N_20770,N_20628,N_20627);
xnor U20771 (N_20771,N_20638,N_20582);
nor U20772 (N_20772,N_20547,N_20570);
or U20773 (N_20773,N_20617,N_20646);
nor U20774 (N_20774,N_20537,N_20506);
and U20775 (N_20775,N_20533,N_20531);
nand U20776 (N_20776,N_20717,N_20679);
xnor U20777 (N_20777,N_20647,N_20690);
nor U20778 (N_20778,N_20588,N_20539);
and U20779 (N_20779,N_20522,N_20718);
xor U20780 (N_20780,N_20672,N_20562);
xnor U20781 (N_20781,N_20703,N_20505);
and U20782 (N_20782,N_20503,N_20527);
and U20783 (N_20783,N_20519,N_20700);
nor U20784 (N_20784,N_20668,N_20540);
or U20785 (N_20785,N_20692,N_20603);
nor U20786 (N_20786,N_20557,N_20637);
nand U20787 (N_20787,N_20696,N_20596);
nor U20788 (N_20788,N_20662,N_20687);
and U20789 (N_20789,N_20591,N_20632);
nor U20790 (N_20790,N_20676,N_20619);
or U20791 (N_20791,N_20559,N_20701);
or U20792 (N_20792,N_20741,N_20719);
nor U20793 (N_20793,N_20524,N_20615);
xnor U20794 (N_20794,N_20525,N_20558);
nor U20795 (N_20795,N_20744,N_20724);
or U20796 (N_20796,N_20579,N_20622);
nor U20797 (N_20797,N_20633,N_20610);
or U20798 (N_20798,N_20561,N_20652);
nor U20799 (N_20799,N_20733,N_20726);
nand U20800 (N_20800,N_20653,N_20575);
nor U20801 (N_20801,N_20508,N_20658);
nand U20802 (N_20802,N_20535,N_20573);
or U20803 (N_20803,N_20698,N_20589);
nand U20804 (N_20804,N_20636,N_20654);
or U20805 (N_20805,N_20659,N_20710);
nor U20806 (N_20806,N_20734,N_20534);
or U20807 (N_20807,N_20631,N_20608);
nor U20808 (N_20808,N_20640,N_20686);
xnor U20809 (N_20809,N_20510,N_20727);
or U20810 (N_20810,N_20737,N_20688);
nand U20811 (N_20811,N_20645,N_20516);
nand U20812 (N_20812,N_20576,N_20606);
nor U20813 (N_20813,N_20748,N_20641);
or U20814 (N_20814,N_20556,N_20621);
xor U20815 (N_20815,N_20541,N_20566);
nor U20816 (N_20816,N_20552,N_20593);
nor U20817 (N_20817,N_20673,N_20712);
and U20818 (N_20818,N_20605,N_20685);
nand U20819 (N_20819,N_20648,N_20695);
xor U20820 (N_20820,N_20625,N_20528);
xor U20821 (N_20821,N_20512,N_20709);
and U20822 (N_20822,N_20511,N_20613);
or U20823 (N_20823,N_20699,N_20590);
xor U20824 (N_20824,N_20542,N_20580);
xor U20825 (N_20825,N_20732,N_20738);
nor U20826 (N_20826,N_20693,N_20609);
or U20827 (N_20827,N_20597,N_20643);
nand U20828 (N_20828,N_20714,N_20563);
nor U20829 (N_20829,N_20665,N_20572);
xor U20830 (N_20830,N_20683,N_20720);
and U20831 (N_20831,N_20543,N_20517);
and U20832 (N_20832,N_20729,N_20544);
xor U20833 (N_20833,N_20691,N_20507);
xor U20834 (N_20834,N_20730,N_20723);
nor U20835 (N_20835,N_20546,N_20716);
nand U20836 (N_20836,N_20529,N_20735);
nor U20837 (N_20837,N_20538,N_20530);
xnor U20838 (N_20838,N_20594,N_20515);
and U20839 (N_20839,N_20623,N_20514);
and U20840 (N_20840,N_20681,N_20747);
nor U20841 (N_20841,N_20746,N_20574);
or U20842 (N_20842,N_20670,N_20725);
and U20843 (N_20843,N_20721,N_20669);
nand U20844 (N_20844,N_20509,N_20618);
nor U20845 (N_20845,N_20705,N_20521);
and U20846 (N_20846,N_20671,N_20740);
or U20847 (N_20847,N_20677,N_20707);
or U20848 (N_20848,N_20586,N_20713);
and U20849 (N_20849,N_20518,N_20749);
or U20850 (N_20850,N_20664,N_20674);
nor U20851 (N_20851,N_20704,N_20642);
nor U20852 (N_20852,N_20599,N_20667);
nand U20853 (N_20853,N_20532,N_20607);
xor U20854 (N_20854,N_20626,N_20549);
nand U20855 (N_20855,N_20553,N_20614);
xnor U20856 (N_20856,N_20548,N_20624);
nand U20857 (N_20857,N_20577,N_20731);
or U20858 (N_20858,N_20630,N_20657);
xnor U20859 (N_20859,N_20678,N_20500);
nand U20860 (N_20860,N_20578,N_20523);
xnor U20861 (N_20861,N_20581,N_20502);
nand U20862 (N_20862,N_20694,N_20513);
or U20863 (N_20863,N_20560,N_20680);
or U20864 (N_20864,N_20598,N_20504);
or U20865 (N_20865,N_20611,N_20644);
and U20866 (N_20866,N_20711,N_20651);
or U20867 (N_20867,N_20612,N_20545);
and U20868 (N_20868,N_20745,N_20663);
and U20869 (N_20869,N_20666,N_20564);
and U20870 (N_20870,N_20585,N_20684);
and U20871 (N_20871,N_20567,N_20583);
nand U20872 (N_20872,N_20649,N_20501);
nor U20873 (N_20873,N_20639,N_20708);
nand U20874 (N_20874,N_20697,N_20728);
or U20875 (N_20875,N_20714,N_20651);
nor U20876 (N_20876,N_20711,N_20535);
nor U20877 (N_20877,N_20640,N_20641);
nand U20878 (N_20878,N_20518,N_20593);
xnor U20879 (N_20879,N_20701,N_20567);
xnor U20880 (N_20880,N_20641,N_20738);
or U20881 (N_20881,N_20746,N_20721);
nand U20882 (N_20882,N_20666,N_20579);
nor U20883 (N_20883,N_20550,N_20557);
or U20884 (N_20884,N_20505,N_20501);
or U20885 (N_20885,N_20510,N_20689);
and U20886 (N_20886,N_20632,N_20640);
nor U20887 (N_20887,N_20509,N_20555);
or U20888 (N_20888,N_20716,N_20647);
nor U20889 (N_20889,N_20600,N_20678);
nand U20890 (N_20890,N_20578,N_20614);
xor U20891 (N_20891,N_20566,N_20562);
xor U20892 (N_20892,N_20599,N_20614);
nor U20893 (N_20893,N_20553,N_20615);
and U20894 (N_20894,N_20503,N_20650);
xnor U20895 (N_20895,N_20576,N_20635);
and U20896 (N_20896,N_20557,N_20718);
and U20897 (N_20897,N_20535,N_20500);
nor U20898 (N_20898,N_20523,N_20589);
xnor U20899 (N_20899,N_20548,N_20629);
and U20900 (N_20900,N_20690,N_20710);
nor U20901 (N_20901,N_20702,N_20567);
nand U20902 (N_20902,N_20577,N_20729);
nor U20903 (N_20903,N_20739,N_20508);
nand U20904 (N_20904,N_20737,N_20681);
nor U20905 (N_20905,N_20518,N_20746);
and U20906 (N_20906,N_20585,N_20719);
nor U20907 (N_20907,N_20591,N_20737);
xnor U20908 (N_20908,N_20564,N_20638);
and U20909 (N_20909,N_20543,N_20639);
nor U20910 (N_20910,N_20579,N_20613);
nand U20911 (N_20911,N_20672,N_20692);
and U20912 (N_20912,N_20608,N_20509);
xor U20913 (N_20913,N_20569,N_20653);
xnor U20914 (N_20914,N_20672,N_20725);
and U20915 (N_20915,N_20637,N_20592);
nor U20916 (N_20916,N_20553,N_20603);
and U20917 (N_20917,N_20583,N_20665);
and U20918 (N_20918,N_20686,N_20545);
and U20919 (N_20919,N_20514,N_20545);
nor U20920 (N_20920,N_20500,N_20676);
and U20921 (N_20921,N_20703,N_20526);
nor U20922 (N_20922,N_20598,N_20738);
and U20923 (N_20923,N_20650,N_20608);
nor U20924 (N_20924,N_20680,N_20505);
or U20925 (N_20925,N_20577,N_20601);
xnor U20926 (N_20926,N_20553,N_20708);
and U20927 (N_20927,N_20742,N_20684);
and U20928 (N_20928,N_20668,N_20555);
xnor U20929 (N_20929,N_20671,N_20705);
and U20930 (N_20930,N_20569,N_20505);
nand U20931 (N_20931,N_20685,N_20669);
nor U20932 (N_20932,N_20567,N_20504);
nor U20933 (N_20933,N_20555,N_20733);
and U20934 (N_20934,N_20688,N_20570);
or U20935 (N_20935,N_20545,N_20580);
nor U20936 (N_20936,N_20541,N_20716);
xor U20937 (N_20937,N_20501,N_20531);
or U20938 (N_20938,N_20509,N_20506);
xor U20939 (N_20939,N_20723,N_20576);
or U20940 (N_20940,N_20657,N_20523);
nand U20941 (N_20941,N_20570,N_20551);
and U20942 (N_20942,N_20732,N_20627);
or U20943 (N_20943,N_20621,N_20731);
or U20944 (N_20944,N_20623,N_20605);
nor U20945 (N_20945,N_20692,N_20582);
nand U20946 (N_20946,N_20639,N_20531);
and U20947 (N_20947,N_20718,N_20567);
nor U20948 (N_20948,N_20716,N_20568);
xor U20949 (N_20949,N_20711,N_20724);
or U20950 (N_20950,N_20534,N_20660);
and U20951 (N_20951,N_20606,N_20731);
nor U20952 (N_20952,N_20517,N_20746);
and U20953 (N_20953,N_20745,N_20711);
and U20954 (N_20954,N_20689,N_20686);
xor U20955 (N_20955,N_20580,N_20717);
and U20956 (N_20956,N_20670,N_20716);
nand U20957 (N_20957,N_20614,N_20669);
xor U20958 (N_20958,N_20728,N_20572);
nand U20959 (N_20959,N_20513,N_20602);
nand U20960 (N_20960,N_20616,N_20578);
or U20961 (N_20961,N_20710,N_20612);
nor U20962 (N_20962,N_20626,N_20634);
nor U20963 (N_20963,N_20669,N_20528);
or U20964 (N_20964,N_20717,N_20652);
xnor U20965 (N_20965,N_20713,N_20581);
nor U20966 (N_20966,N_20662,N_20635);
or U20967 (N_20967,N_20508,N_20625);
nand U20968 (N_20968,N_20654,N_20653);
nor U20969 (N_20969,N_20634,N_20681);
nor U20970 (N_20970,N_20586,N_20725);
nor U20971 (N_20971,N_20675,N_20724);
xor U20972 (N_20972,N_20630,N_20643);
xor U20973 (N_20973,N_20541,N_20653);
nand U20974 (N_20974,N_20714,N_20613);
nand U20975 (N_20975,N_20714,N_20523);
or U20976 (N_20976,N_20590,N_20581);
nand U20977 (N_20977,N_20557,N_20597);
and U20978 (N_20978,N_20653,N_20682);
and U20979 (N_20979,N_20664,N_20517);
nand U20980 (N_20980,N_20744,N_20668);
or U20981 (N_20981,N_20725,N_20744);
or U20982 (N_20982,N_20685,N_20641);
and U20983 (N_20983,N_20560,N_20513);
and U20984 (N_20984,N_20649,N_20563);
nand U20985 (N_20985,N_20554,N_20736);
xor U20986 (N_20986,N_20500,N_20667);
or U20987 (N_20987,N_20731,N_20596);
or U20988 (N_20988,N_20564,N_20532);
or U20989 (N_20989,N_20605,N_20712);
nor U20990 (N_20990,N_20699,N_20563);
xnor U20991 (N_20991,N_20566,N_20635);
or U20992 (N_20992,N_20620,N_20605);
or U20993 (N_20993,N_20708,N_20743);
or U20994 (N_20994,N_20655,N_20520);
nor U20995 (N_20995,N_20534,N_20599);
and U20996 (N_20996,N_20717,N_20648);
and U20997 (N_20997,N_20541,N_20527);
nand U20998 (N_20998,N_20642,N_20626);
nor U20999 (N_20999,N_20671,N_20526);
or U21000 (N_21000,N_20933,N_20946);
or U21001 (N_21001,N_20878,N_20778);
and U21002 (N_21002,N_20928,N_20782);
nand U21003 (N_21003,N_20965,N_20982);
xor U21004 (N_21004,N_20823,N_20947);
nor U21005 (N_21005,N_20981,N_20858);
nand U21006 (N_21006,N_20880,N_20934);
or U21007 (N_21007,N_20884,N_20828);
nor U21008 (N_21008,N_20961,N_20786);
xnor U21009 (N_21009,N_20832,N_20830);
or U21010 (N_21010,N_20849,N_20990);
nand U21011 (N_21011,N_20795,N_20894);
xnor U21012 (N_21012,N_20789,N_20794);
and U21013 (N_21013,N_20792,N_20975);
and U21014 (N_21014,N_20954,N_20930);
nor U21015 (N_21015,N_20783,N_20963);
and U21016 (N_21016,N_20993,N_20898);
xnor U21017 (N_21017,N_20814,N_20911);
xor U21018 (N_21018,N_20809,N_20979);
nand U21019 (N_21019,N_20775,N_20756);
nor U21020 (N_21020,N_20773,N_20888);
or U21021 (N_21021,N_20970,N_20939);
xnor U21022 (N_21022,N_20781,N_20945);
nor U21023 (N_21023,N_20989,N_20905);
or U21024 (N_21024,N_20763,N_20974);
and U21025 (N_21025,N_20998,N_20863);
xnor U21026 (N_21026,N_20799,N_20811);
nand U21027 (N_21027,N_20834,N_20914);
or U21028 (N_21028,N_20772,N_20761);
and U21029 (N_21029,N_20854,N_20774);
xnor U21030 (N_21030,N_20831,N_20956);
xnor U21031 (N_21031,N_20952,N_20833);
nor U21032 (N_21032,N_20948,N_20818);
xor U21033 (N_21033,N_20983,N_20912);
nand U21034 (N_21034,N_20919,N_20779);
or U21035 (N_21035,N_20882,N_20924);
nand U21036 (N_21036,N_20867,N_20759);
and U21037 (N_21037,N_20966,N_20860);
and U21038 (N_21038,N_20904,N_20903);
nor U21039 (N_21039,N_20855,N_20829);
nor U21040 (N_21040,N_20790,N_20932);
xor U21041 (N_21041,N_20900,N_20908);
and U21042 (N_21042,N_20896,N_20796);
xnor U21043 (N_21043,N_20897,N_20845);
xnor U21044 (N_21044,N_20967,N_20870);
and U21045 (N_21045,N_20788,N_20874);
nand U21046 (N_21046,N_20943,N_20959);
nor U21047 (N_21047,N_20869,N_20899);
or U21048 (N_21048,N_20807,N_20852);
and U21049 (N_21049,N_20771,N_20913);
or U21050 (N_21050,N_20962,N_20995);
or U21051 (N_21051,N_20824,N_20950);
and U21052 (N_21052,N_20866,N_20769);
xor U21053 (N_21053,N_20978,N_20926);
nor U21054 (N_21054,N_20840,N_20889);
and U21055 (N_21055,N_20953,N_20879);
and U21056 (N_21056,N_20838,N_20992);
or U21057 (N_21057,N_20750,N_20754);
and U21058 (N_21058,N_20810,N_20784);
nand U21059 (N_21059,N_20753,N_20921);
nor U21060 (N_21060,N_20920,N_20976);
and U21061 (N_21061,N_20996,N_20909);
xor U21062 (N_21062,N_20877,N_20785);
xor U21063 (N_21063,N_20800,N_20893);
nand U21064 (N_21064,N_20910,N_20780);
xor U21065 (N_21065,N_20787,N_20836);
xnor U21066 (N_21066,N_20865,N_20891);
nor U21067 (N_21067,N_20841,N_20819);
or U21068 (N_21068,N_20940,N_20915);
and U21069 (N_21069,N_20797,N_20941);
xnor U21070 (N_21070,N_20886,N_20927);
or U21071 (N_21071,N_20951,N_20872);
nor U21072 (N_21072,N_20842,N_20890);
nor U21073 (N_21073,N_20839,N_20895);
xor U21074 (N_21074,N_20760,N_20805);
nand U21075 (N_21075,N_20881,N_20821);
or U21076 (N_21076,N_20757,N_20848);
nand U21077 (N_21077,N_20765,N_20862);
and U21078 (N_21078,N_20907,N_20885);
xor U21079 (N_21079,N_20931,N_20923);
nor U21080 (N_21080,N_20980,N_20837);
nor U21081 (N_21081,N_20850,N_20957);
nor U21082 (N_21082,N_20958,N_20851);
or U21083 (N_21083,N_20815,N_20826);
nor U21084 (N_21084,N_20917,N_20949);
and U21085 (N_21085,N_20804,N_20803);
nand U21086 (N_21086,N_20971,N_20938);
nand U21087 (N_21087,N_20857,N_20859);
xnor U21088 (N_21088,N_20770,N_20973);
nor U21089 (N_21089,N_20964,N_20856);
and U21090 (N_21090,N_20922,N_20793);
nand U21091 (N_21091,N_20752,N_20916);
nand U21092 (N_21092,N_20984,N_20843);
or U21093 (N_21093,N_20901,N_20994);
xor U21094 (N_21094,N_20798,N_20883);
nor U21095 (N_21095,N_20892,N_20827);
nor U21096 (N_21096,N_20768,N_20758);
nor U21097 (N_21097,N_20847,N_20825);
nor U21098 (N_21098,N_20813,N_20868);
or U21099 (N_21099,N_20844,N_20887);
xor U21100 (N_21100,N_20755,N_20935);
and U21101 (N_21101,N_20751,N_20861);
xor U21102 (N_21102,N_20942,N_20972);
or U21103 (N_21103,N_20846,N_20767);
xor U21104 (N_21104,N_20764,N_20816);
nor U21105 (N_21105,N_20925,N_20776);
nor U21106 (N_21106,N_20985,N_20969);
and U21107 (N_21107,N_20802,N_20968);
or U21108 (N_21108,N_20944,N_20762);
nor U21109 (N_21109,N_20929,N_20801);
nor U21110 (N_21110,N_20791,N_20937);
nand U21111 (N_21111,N_20835,N_20997);
or U21112 (N_21112,N_20875,N_20777);
xnor U21113 (N_21113,N_20999,N_20906);
xnor U21114 (N_21114,N_20808,N_20988);
and U21115 (N_21115,N_20822,N_20986);
or U21116 (N_21116,N_20960,N_20955);
or U21117 (N_21117,N_20876,N_20902);
xnor U21118 (N_21118,N_20864,N_20766);
nor U21119 (N_21119,N_20871,N_20918);
and U21120 (N_21120,N_20817,N_20812);
xnor U21121 (N_21121,N_20853,N_20987);
and U21122 (N_21122,N_20977,N_20806);
or U21123 (N_21123,N_20820,N_20991);
xor U21124 (N_21124,N_20936,N_20873);
and U21125 (N_21125,N_20894,N_20805);
xnor U21126 (N_21126,N_20903,N_20839);
and U21127 (N_21127,N_20770,N_20879);
and U21128 (N_21128,N_20949,N_20860);
nand U21129 (N_21129,N_20856,N_20928);
nor U21130 (N_21130,N_20926,N_20753);
and U21131 (N_21131,N_20879,N_20904);
xor U21132 (N_21132,N_20917,N_20934);
xnor U21133 (N_21133,N_20761,N_20988);
nor U21134 (N_21134,N_20962,N_20956);
or U21135 (N_21135,N_20760,N_20905);
or U21136 (N_21136,N_20893,N_20897);
xor U21137 (N_21137,N_20986,N_20881);
xnor U21138 (N_21138,N_20793,N_20995);
xnor U21139 (N_21139,N_20920,N_20853);
nor U21140 (N_21140,N_20955,N_20925);
nand U21141 (N_21141,N_20855,N_20769);
nand U21142 (N_21142,N_20974,N_20994);
xor U21143 (N_21143,N_20756,N_20912);
or U21144 (N_21144,N_20835,N_20828);
nor U21145 (N_21145,N_20881,N_20799);
nand U21146 (N_21146,N_20979,N_20931);
or U21147 (N_21147,N_20786,N_20964);
nor U21148 (N_21148,N_20820,N_20756);
or U21149 (N_21149,N_20892,N_20900);
xor U21150 (N_21150,N_20774,N_20938);
or U21151 (N_21151,N_20819,N_20809);
and U21152 (N_21152,N_20841,N_20875);
nand U21153 (N_21153,N_20851,N_20902);
nand U21154 (N_21154,N_20768,N_20909);
nor U21155 (N_21155,N_20750,N_20978);
xnor U21156 (N_21156,N_20786,N_20753);
or U21157 (N_21157,N_20982,N_20779);
and U21158 (N_21158,N_20951,N_20845);
xnor U21159 (N_21159,N_20843,N_20954);
nor U21160 (N_21160,N_20765,N_20809);
and U21161 (N_21161,N_20795,N_20942);
xor U21162 (N_21162,N_20986,N_20914);
nor U21163 (N_21163,N_20887,N_20847);
nand U21164 (N_21164,N_20857,N_20804);
or U21165 (N_21165,N_20919,N_20982);
and U21166 (N_21166,N_20816,N_20845);
or U21167 (N_21167,N_20911,N_20772);
nor U21168 (N_21168,N_20999,N_20893);
xor U21169 (N_21169,N_20816,N_20921);
xnor U21170 (N_21170,N_20752,N_20919);
and U21171 (N_21171,N_20797,N_20861);
nand U21172 (N_21172,N_20992,N_20965);
nor U21173 (N_21173,N_20907,N_20819);
xor U21174 (N_21174,N_20996,N_20961);
nor U21175 (N_21175,N_20799,N_20892);
and U21176 (N_21176,N_20758,N_20815);
nand U21177 (N_21177,N_20853,N_20961);
and U21178 (N_21178,N_20946,N_20863);
nand U21179 (N_21179,N_20769,N_20869);
xnor U21180 (N_21180,N_20917,N_20820);
or U21181 (N_21181,N_20760,N_20929);
or U21182 (N_21182,N_20951,N_20794);
and U21183 (N_21183,N_20819,N_20936);
or U21184 (N_21184,N_20882,N_20764);
nand U21185 (N_21185,N_20933,N_20976);
nor U21186 (N_21186,N_20764,N_20905);
and U21187 (N_21187,N_20961,N_20937);
or U21188 (N_21188,N_20973,N_20808);
nor U21189 (N_21189,N_20843,N_20811);
nand U21190 (N_21190,N_20924,N_20971);
and U21191 (N_21191,N_20768,N_20778);
nand U21192 (N_21192,N_20913,N_20884);
and U21193 (N_21193,N_20841,N_20779);
and U21194 (N_21194,N_20936,N_20803);
nor U21195 (N_21195,N_20842,N_20956);
xor U21196 (N_21196,N_20801,N_20789);
xnor U21197 (N_21197,N_20984,N_20799);
nor U21198 (N_21198,N_20906,N_20980);
and U21199 (N_21199,N_20913,N_20785);
nor U21200 (N_21200,N_20976,N_20776);
nor U21201 (N_21201,N_20853,N_20985);
or U21202 (N_21202,N_20850,N_20788);
or U21203 (N_21203,N_20761,N_20790);
or U21204 (N_21204,N_20950,N_20990);
or U21205 (N_21205,N_20829,N_20836);
or U21206 (N_21206,N_20752,N_20787);
nor U21207 (N_21207,N_20904,N_20949);
or U21208 (N_21208,N_20781,N_20857);
or U21209 (N_21209,N_20928,N_20893);
xnor U21210 (N_21210,N_20838,N_20975);
and U21211 (N_21211,N_20857,N_20807);
nand U21212 (N_21212,N_20772,N_20770);
nor U21213 (N_21213,N_20753,N_20930);
and U21214 (N_21214,N_20867,N_20970);
nor U21215 (N_21215,N_20876,N_20921);
or U21216 (N_21216,N_20865,N_20877);
xnor U21217 (N_21217,N_20831,N_20815);
nand U21218 (N_21218,N_20898,N_20781);
or U21219 (N_21219,N_20902,N_20763);
nand U21220 (N_21220,N_20909,N_20807);
xor U21221 (N_21221,N_20915,N_20883);
xnor U21222 (N_21222,N_20839,N_20784);
and U21223 (N_21223,N_20926,N_20817);
or U21224 (N_21224,N_20834,N_20930);
nor U21225 (N_21225,N_20994,N_20991);
or U21226 (N_21226,N_20991,N_20944);
or U21227 (N_21227,N_20928,N_20840);
or U21228 (N_21228,N_20997,N_20816);
xnor U21229 (N_21229,N_20861,N_20792);
nand U21230 (N_21230,N_20817,N_20802);
xor U21231 (N_21231,N_20778,N_20952);
nor U21232 (N_21232,N_20878,N_20909);
or U21233 (N_21233,N_20978,N_20903);
xor U21234 (N_21234,N_20987,N_20837);
xnor U21235 (N_21235,N_20845,N_20992);
nor U21236 (N_21236,N_20838,N_20910);
and U21237 (N_21237,N_20989,N_20916);
nand U21238 (N_21238,N_20784,N_20972);
nand U21239 (N_21239,N_20761,N_20982);
or U21240 (N_21240,N_20967,N_20992);
and U21241 (N_21241,N_20834,N_20785);
and U21242 (N_21242,N_20839,N_20984);
nor U21243 (N_21243,N_20921,N_20815);
nor U21244 (N_21244,N_20923,N_20982);
nand U21245 (N_21245,N_20973,N_20826);
nand U21246 (N_21246,N_20883,N_20937);
or U21247 (N_21247,N_20903,N_20932);
xnor U21248 (N_21248,N_20976,N_20780);
xor U21249 (N_21249,N_20820,N_20829);
or U21250 (N_21250,N_21229,N_21037);
and U21251 (N_21251,N_21227,N_21099);
nand U21252 (N_21252,N_21181,N_21092);
or U21253 (N_21253,N_21019,N_21151);
nand U21254 (N_21254,N_21248,N_21086);
nand U21255 (N_21255,N_21088,N_21035);
nor U21256 (N_21256,N_21200,N_21081);
nor U21257 (N_21257,N_21029,N_21185);
and U21258 (N_21258,N_21093,N_21196);
nor U21259 (N_21259,N_21194,N_21209);
nand U21260 (N_21260,N_21098,N_21212);
nand U21261 (N_21261,N_21144,N_21179);
or U21262 (N_21262,N_21110,N_21247);
nand U21263 (N_21263,N_21182,N_21084);
nand U21264 (N_21264,N_21188,N_21038);
and U21265 (N_21265,N_21053,N_21156);
nand U21266 (N_21266,N_21062,N_21127);
and U21267 (N_21267,N_21170,N_21136);
nand U21268 (N_21268,N_21075,N_21243);
or U21269 (N_21269,N_21071,N_21042);
or U21270 (N_21270,N_21187,N_21103);
nand U21271 (N_21271,N_21234,N_21207);
xor U21272 (N_21272,N_21108,N_21014);
xnor U21273 (N_21273,N_21007,N_21226);
and U21274 (N_21274,N_21126,N_21223);
or U21275 (N_21275,N_21246,N_21055);
or U21276 (N_21276,N_21024,N_21155);
xnor U21277 (N_21277,N_21150,N_21199);
nor U21278 (N_21278,N_21089,N_21186);
or U21279 (N_21279,N_21060,N_21013);
nor U21280 (N_21280,N_21245,N_21009);
xor U21281 (N_21281,N_21215,N_21195);
or U21282 (N_21282,N_21167,N_21090);
xor U21283 (N_21283,N_21046,N_21027);
nor U21284 (N_21284,N_21122,N_21079);
and U21285 (N_21285,N_21161,N_21074);
or U21286 (N_21286,N_21069,N_21119);
and U21287 (N_21287,N_21214,N_21201);
nor U21288 (N_21288,N_21218,N_21111);
nand U21289 (N_21289,N_21077,N_21008);
or U21290 (N_21290,N_21033,N_21238);
nand U21291 (N_21291,N_21052,N_21100);
nand U21292 (N_21292,N_21141,N_21131);
nor U21293 (N_21293,N_21034,N_21242);
xnor U21294 (N_21294,N_21070,N_21138);
and U21295 (N_21295,N_21180,N_21235);
or U21296 (N_21296,N_21130,N_21148);
nor U21297 (N_21297,N_21058,N_21220);
or U21298 (N_21298,N_21190,N_21076);
or U21299 (N_21299,N_21172,N_21010);
and U21300 (N_21300,N_21117,N_21211);
nor U21301 (N_21301,N_21085,N_21005);
nand U21302 (N_21302,N_21118,N_21178);
or U21303 (N_21303,N_21173,N_21032);
nand U21304 (N_21304,N_21073,N_21044);
or U21305 (N_21305,N_21083,N_21132);
or U21306 (N_21306,N_21232,N_21147);
xor U21307 (N_21307,N_21241,N_21031);
and U21308 (N_21308,N_21094,N_21056);
xor U21309 (N_21309,N_21221,N_21154);
and U21310 (N_21310,N_21114,N_21228);
nand U21311 (N_21311,N_21191,N_21149);
and U21312 (N_21312,N_21217,N_21137);
and U21313 (N_21313,N_21164,N_21159);
and U21314 (N_21314,N_21125,N_21050);
xor U21315 (N_21315,N_21123,N_21012);
or U21316 (N_21316,N_21080,N_21121);
xnor U21317 (N_21317,N_21171,N_21017);
and U21318 (N_21318,N_21135,N_21129);
xor U21319 (N_21319,N_21030,N_21006);
nor U21320 (N_21320,N_21061,N_21219);
nor U21321 (N_21321,N_21028,N_21249);
and U21322 (N_21322,N_21040,N_21020);
and U21323 (N_21323,N_21107,N_21018);
or U21324 (N_21324,N_21002,N_21210);
xor U21325 (N_21325,N_21021,N_21239);
xor U21326 (N_21326,N_21134,N_21054);
nand U21327 (N_21327,N_21000,N_21204);
nand U21328 (N_21328,N_21128,N_21152);
nand U21329 (N_21329,N_21183,N_21140);
and U21330 (N_21330,N_21169,N_21142);
xnor U21331 (N_21331,N_21025,N_21174);
xor U21332 (N_21332,N_21225,N_21068);
or U21333 (N_21333,N_21213,N_21015);
or U21334 (N_21334,N_21036,N_21049);
nand U21335 (N_21335,N_21115,N_21203);
xor U21336 (N_21336,N_21189,N_21166);
nor U21337 (N_21337,N_21124,N_21244);
and U21338 (N_21338,N_21096,N_21120);
nand U21339 (N_21339,N_21163,N_21116);
or U21340 (N_21340,N_21113,N_21082);
xor U21341 (N_21341,N_21157,N_21197);
nand U21342 (N_21342,N_21066,N_21063);
and U21343 (N_21343,N_21146,N_21237);
nor U21344 (N_21344,N_21177,N_21065);
nand U21345 (N_21345,N_21067,N_21139);
or U21346 (N_21346,N_21233,N_21011);
xnor U21347 (N_21347,N_21192,N_21095);
or U21348 (N_21348,N_21101,N_21160);
nor U21349 (N_21349,N_21153,N_21039);
and U21350 (N_21350,N_21087,N_21202);
nand U21351 (N_21351,N_21158,N_21236);
nor U21352 (N_21352,N_21105,N_21059);
or U21353 (N_21353,N_21003,N_21222);
and U21354 (N_21354,N_21048,N_21102);
nor U21355 (N_21355,N_21175,N_21112);
and U21356 (N_21356,N_21193,N_21057);
and U21357 (N_21357,N_21165,N_21026);
nand U21358 (N_21358,N_21184,N_21023);
or U21359 (N_21359,N_21001,N_21072);
nor U21360 (N_21360,N_21145,N_21143);
or U21361 (N_21361,N_21104,N_21043);
nor U21362 (N_21362,N_21091,N_21133);
or U21363 (N_21363,N_21047,N_21078);
nand U21364 (N_21364,N_21045,N_21162);
and U21365 (N_21365,N_21206,N_21022);
and U21366 (N_21366,N_21176,N_21231);
xnor U21367 (N_21367,N_21198,N_21064);
nor U21368 (N_21368,N_21208,N_21168);
xnor U21369 (N_21369,N_21205,N_21004);
or U21370 (N_21370,N_21230,N_21041);
nor U21371 (N_21371,N_21216,N_21109);
or U21372 (N_21372,N_21016,N_21224);
and U21373 (N_21373,N_21097,N_21051);
xor U21374 (N_21374,N_21106,N_21240);
nor U21375 (N_21375,N_21165,N_21067);
nor U21376 (N_21376,N_21018,N_21242);
and U21377 (N_21377,N_21071,N_21094);
or U21378 (N_21378,N_21042,N_21013);
and U21379 (N_21379,N_21187,N_21144);
or U21380 (N_21380,N_21038,N_21247);
nor U21381 (N_21381,N_21247,N_21065);
or U21382 (N_21382,N_21218,N_21115);
nor U21383 (N_21383,N_21041,N_21151);
nand U21384 (N_21384,N_21129,N_21068);
and U21385 (N_21385,N_21151,N_21191);
and U21386 (N_21386,N_21160,N_21038);
and U21387 (N_21387,N_21022,N_21159);
nand U21388 (N_21388,N_21238,N_21199);
and U21389 (N_21389,N_21227,N_21085);
nand U21390 (N_21390,N_21182,N_21119);
nand U21391 (N_21391,N_21236,N_21166);
or U21392 (N_21392,N_21107,N_21150);
xor U21393 (N_21393,N_21147,N_21221);
xor U21394 (N_21394,N_21017,N_21060);
nand U21395 (N_21395,N_21240,N_21019);
or U21396 (N_21396,N_21038,N_21180);
nand U21397 (N_21397,N_21031,N_21117);
nor U21398 (N_21398,N_21036,N_21007);
xnor U21399 (N_21399,N_21141,N_21201);
xnor U21400 (N_21400,N_21177,N_21132);
or U21401 (N_21401,N_21223,N_21249);
and U21402 (N_21402,N_21236,N_21244);
xor U21403 (N_21403,N_21074,N_21062);
nand U21404 (N_21404,N_21084,N_21228);
or U21405 (N_21405,N_21111,N_21139);
or U21406 (N_21406,N_21058,N_21010);
nor U21407 (N_21407,N_21090,N_21152);
xnor U21408 (N_21408,N_21058,N_21153);
xor U21409 (N_21409,N_21071,N_21234);
and U21410 (N_21410,N_21087,N_21022);
nand U21411 (N_21411,N_21187,N_21243);
nor U21412 (N_21412,N_21209,N_21000);
and U21413 (N_21413,N_21110,N_21168);
nor U21414 (N_21414,N_21067,N_21235);
and U21415 (N_21415,N_21170,N_21076);
xnor U21416 (N_21416,N_21161,N_21115);
nor U21417 (N_21417,N_21109,N_21149);
and U21418 (N_21418,N_21127,N_21189);
and U21419 (N_21419,N_21180,N_21002);
nor U21420 (N_21420,N_21140,N_21065);
nand U21421 (N_21421,N_21030,N_21144);
xnor U21422 (N_21422,N_21012,N_21181);
nor U21423 (N_21423,N_21174,N_21064);
nand U21424 (N_21424,N_21110,N_21034);
xnor U21425 (N_21425,N_21148,N_21187);
and U21426 (N_21426,N_21240,N_21014);
or U21427 (N_21427,N_21188,N_21204);
xnor U21428 (N_21428,N_21087,N_21207);
nor U21429 (N_21429,N_21175,N_21241);
xor U21430 (N_21430,N_21202,N_21126);
xnor U21431 (N_21431,N_21192,N_21104);
nor U21432 (N_21432,N_21008,N_21027);
or U21433 (N_21433,N_21206,N_21240);
or U21434 (N_21434,N_21206,N_21241);
nor U21435 (N_21435,N_21214,N_21013);
or U21436 (N_21436,N_21237,N_21236);
and U21437 (N_21437,N_21136,N_21150);
and U21438 (N_21438,N_21033,N_21160);
xnor U21439 (N_21439,N_21123,N_21161);
nor U21440 (N_21440,N_21009,N_21035);
and U21441 (N_21441,N_21027,N_21133);
and U21442 (N_21442,N_21050,N_21077);
nand U21443 (N_21443,N_21002,N_21120);
and U21444 (N_21444,N_21211,N_21183);
nor U21445 (N_21445,N_21033,N_21192);
and U21446 (N_21446,N_21164,N_21143);
nand U21447 (N_21447,N_21153,N_21070);
nor U21448 (N_21448,N_21247,N_21152);
or U21449 (N_21449,N_21006,N_21184);
xor U21450 (N_21450,N_21153,N_21071);
nor U21451 (N_21451,N_21185,N_21023);
xor U21452 (N_21452,N_21062,N_21171);
nor U21453 (N_21453,N_21152,N_21211);
nor U21454 (N_21454,N_21114,N_21238);
or U21455 (N_21455,N_21050,N_21038);
nor U21456 (N_21456,N_21152,N_21097);
nor U21457 (N_21457,N_21005,N_21104);
or U21458 (N_21458,N_21020,N_21184);
or U21459 (N_21459,N_21072,N_21174);
or U21460 (N_21460,N_21131,N_21185);
nand U21461 (N_21461,N_21181,N_21242);
and U21462 (N_21462,N_21121,N_21057);
xnor U21463 (N_21463,N_21086,N_21076);
nand U21464 (N_21464,N_21194,N_21235);
and U21465 (N_21465,N_21031,N_21171);
nand U21466 (N_21466,N_21033,N_21154);
nor U21467 (N_21467,N_21137,N_21109);
nor U21468 (N_21468,N_21239,N_21206);
nor U21469 (N_21469,N_21115,N_21193);
and U21470 (N_21470,N_21101,N_21214);
xnor U21471 (N_21471,N_21032,N_21111);
nand U21472 (N_21472,N_21227,N_21247);
xor U21473 (N_21473,N_21191,N_21115);
xnor U21474 (N_21474,N_21180,N_21059);
or U21475 (N_21475,N_21142,N_21233);
nand U21476 (N_21476,N_21211,N_21049);
and U21477 (N_21477,N_21174,N_21214);
nand U21478 (N_21478,N_21041,N_21204);
nor U21479 (N_21479,N_21141,N_21194);
nor U21480 (N_21480,N_21186,N_21130);
or U21481 (N_21481,N_21154,N_21137);
xor U21482 (N_21482,N_21092,N_21096);
and U21483 (N_21483,N_21200,N_21119);
xnor U21484 (N_21484,N_21201,N_21116);
nor U21485 (N_21485,N_21181,N_21085);
xor U21486 (N_21486,N_21028,N_21006);
xor U21487 (N_21487,N_21232,N_21166);
xnor U21488 (N_21488,N_21005,N_21067);
xnor U21489 (N_21489,N_21218,N_21173);
nand U21490 (N_21490,N_21156,N_21016);
or U21491 (N_21491,N_21105,N_21097);
nor U21492 (N_21492,N_21018,N_21073);
and U21493 (N_21493,N_21197,N_21004);
nor U21494 (N_21494,N_21085,N_21161);
nor U21495 (N_21495,N_21190,N_21219);
nor U21496 (N_21496,N_21158,N_21167);
xor U21497 (N_21497,N_21181,N_21057);
or U21498 (N_21498,N_21160,N_21234);
or U21499 (N_21499,N_21114,N_21205);
or U21500 (N_21500,N_21465,N_21455);
and U21501 (N_21501,N_21315,N_21361);
nor U21502 (N_21502,N_21440,N_21392);
xor U21503 (N_21503,N_21310,N_21384);
nor U21504 (N_21504,N_21468,N_21401);
xor U21505 (N_21505,N_21283,N_21297);
nor U21506 (N_21506,N_21447,N_21370);
and U21507 (N_21507,N_21369,N_21335);
nor U21508 (N_21508,N_21341,N_21357);
nand U21509 (N_21509,N_21489,N_21279);
xnor U21510 (N_21510,N_21433,N_21428);
nor U21511 (N_21511,N_21438,N_21343);
nand U21512 (N_21512,N_21454,N_21266);
nor U21513 (N_21513,N_21367,N_21352);
and U21514 (N_21514,N_21265,N_21309);
and U21515 (N_21515,N_21379,N_21270);
or U21516 (N_21516,N_21462,N_21368);
nor U21517 (N_21517,N_21360,N_21282);
or U21518 (N_21518,N_21486,N_21424);
xnor U21519 (N_21519,N_21364,N_21332);
or U21520 (N_21520,N_21291,N_21487);
nor U21521 (N_21521,N_21408,N_21426);
nor U21522 (N_21522,N_21432,N_21444);
and U21523 (N_21523,N_21460,N_21313);
nor U21524 (N_21524,N_21490,N_21345);
nand U21525 (N_21525,N_21481,N_21336);
and U21526 (N_21526,N_21316,N_21496);
or U21527 (N_21527,N_21308,N_21453);
xnor U21528 (N_21528,N_21268,N_21449);
nor U21529 (N_21529,N_21417,N_21331);
nand U21530 (N_21530,N_21395,N_21495);
xor U21531 (N_21531,N_21380,N_21287);
or U21532 (N_21532,N_21353,N_21302);
or U21533 (N_21533,N_21320,N_21294);
or U21534 (N_21534,N_21480,N_21328);
or U21535 (N_21535,N_21347,N_21427);
or U21536 (N_21536,N_21330,N_21418);
nand U21537 (N_21537,N_21425,N_21373);
xnor U21538 (N_21538,N_21351,N_21323);
nor U21539 (N_21539,N_21488,N_21470);
and U21540 (N_21540,N_21406,N_21419);
nor U21541 (N_21541,N_21355,N_21293);
or U21542 (N_21542,N_21333,N_21356);
or U21543 (N_21543,N_21262,N_21349);
nor U21544 (N_21544,N_21482,N_21322);
xor U21545 (N_21545,N_21376,N_21388);
nand U21546 (N_21546,N_21307,N_21327);
and U21547 (N_21547,N_21437,N_21475);
and U21548 (N_21548,N_21461,N_21259);
and U21549 (N_21549,N_21421,N_21324);
nor U21550 (N_21550,N_21387,N_21374);
nor U21551 (N_21551,N_21366,N_21340);
nor U21552 (N_21552,N_21371,N_21292);
or U21553 (N_21553,N_21415,N_21457);
and U21554 (N_21554,N_21446,N_21458);
nor U21555 (N_21555,N_21365,N_21346);
xnor U21556 (N_21556,N_21300,N_21445);
nor U21557 (N_21557,N_21338,N_21325);
or U21558 (N_21558,N_21305,N_21411);
or U21559 (N_21559,N_21251,N_21478);
xnor U21560 (N_21560,N_21312,N_21258);
nand U21561 (N_21561,N_21377,N_21381);
or U21562 (N_21562,N_21362,N_21334);
and U21563 (N_21563,N_21469,N_21255);
or U21564 (N_21564,N_21375,N_21301);
nor U21565 (N_21565,N_21275,N_21409);
and U21566 (N_21566,N_21267,N_21314);
nand U21567 (N_21567,N_21393,N_21280);
nand U21568 (N_21568,N_21382,N_21413);
xnor U21569 (N_21569,N_21286,N_21272);
xnor U21570 (N_21570,N_21386,N_21319);
or U21571 (N_21571,N_21402,N_21303);
and U21572 (N_21572,N_21442,N_21289);
nor U21573 (N_21573,N_21423,N_21483);
or U21574 (N_21574,N_21311,N_21403);
nand U21575 (N_21575,N_21463,N_21493);
nand U21576 (N_21576,N_21306,N_21288);
nor U21577 (N_21577,N_21261,N_21491);
xor U21578 (N_21578,N_21354,N_21420);
nor U21579 (N_21579,N_21430,N_21263);
xnor U21580 (N_21580,N_21396,N_21296);
xor U21581 (N_21581,N_21256,N_21295);
nand U21582 (N_21582,N_21492,N_21337);
nor U21583 (N_21583,N_21274,N_21474);
xor U21584 (N_21584,N_21476,N_21359);
xor U21585 (N_21585,N_21264,N_21344);
nand U21586 (N_21586,N_21498,N_21318);
xnor U21587 (N_21587,N_21407,N_21254);
nor U21588 (N_21588,N_21434,N_21405);
or U21589 (N_21589,N_21390,N_21435);
and U21590 (N_21590,N_21412,N_21451);
nor U21591 (N_21591,N_21383,N_21410);
nand U21592 (N_21592,N_21389,N_21276);
or U21593 (N_21593,N_21278,N_21441);
nand U21594 (N_21594,N_21404,N_21273);
xnor U21595 (N_21595,N_21277,N_21443);
nor U21596 (N_21596,N_21391,N_21342);
nor U21597 (N_21597,N_21363,N_21339);
and U21598 (N_21598,N_21416,N_21399);
xor U21599 (N_21599,N_21252,N_21271);
nand U21600 (N_21600,N_21452,N_21400);
or U21601 (N_21601,N_21350,N_21448);
nor U21602 (N_21602,N_21397,N_21281);
or U21603 (N_21603,N_21485,N_21450);
xnor U21604 (N_21604,N_21464,N_21260);
and U21605 (N_21605,N_21431,N_21253);
or U21606 (N_21606,N_21473,N_21250);
nor U21607 (N_21607,N_21467,N_21494);
or U21608 (N_21608,N_21439,N_21479);
nor U21609 (N_21609,N_21484,N_21436);
and U21610 (N_21610,N_21317,N_21459);
nor U21611 (N_21611,N_21290,N_21497);
nor U21612 (N_21612,N_21358,N_21422);
nand U21613 (N_21613,N_21348,N_21466);
xor U21614 (N_21614,N_21398,N_21329);
or U21615 (N_21615,N_21499,N_21269);
xor U21616 (N_21616,N_21429,N_21385);
nor U21617 (N_21617,N_21378,N_21372);
nand U21618 (N_21618,N_21321,N_21299);
xor U21619 (N_21619,N_21298,N_21414);
nor U21620 (N_21620,N_21326,N_21284);
or U21621 (N_21621,N_21472,N_21285);
or U21622 (N_21622,N_21471,N_21394);
nand U21623 (N_21623,N_21477,N_21257);
xor U21624 (N_21624,N_21456,N_21304);
and U21625 (N_21625,N_21331,N_21403);
or U21626 (N_21626,N_21453,N_21482);
or U21627 (N_21627,N_21322,N_21268);
and U21628 (N_21628,N_21395,N_21376);
nand U21629 (N_21629,N_21455,N_21382);
nand U21630 (N_21630,N_21479,N_21251);
nor U21631 (N_21631,N_21291,N_21258);
or U21632 (N_21632,N_21441,N_21287);
and U21633 (N_21633,N_21271,N_21284);
xor U21634 (N_21634,N_21302,N_21250);
xor U21635 (N_21635,N_21278,N_21462);
and U21636 (N_21636,N_21487,N_21370);
xnor U21637 (N_21637,N_21344,N_21255);
nor U21638 (N_21638,N_21297,N_21378);
or U21639 (N_21639,N_21476,N_21333);
and U21640 (N_21640,N_21250,N_21349);
and U21641 (N_21641,N_21464,N_21307);
nor U21642 (N_21642,N_21489,N_21470);
nor U21643 (N_21643,N_21387,N_21378);
nand U21644 (N_21644,N_21415,N_21295);
nand U21645 (N_21645,N_21432,N_21370);
xnor U21646 (N_21646,N_21371,N_21441);
nand U21647 (N_21647,N_21376,N_21251);
xor U21648 (N_21648,N_21334,N_21306);
nand U21649 (N_21649,N_21359,N_21406);
and U21650 (N_21650,N_21362,N_21253);
or U21651 (N_21651,N_21356,N_21433);
nor U21652 (N_21652,N_21430,N_21433);
nor U21653 (N_21653,N_21279,N_21477);
xnor U21654 (N_21654,N_21263,N_21393);
or U21655 (N_21655,N_21336,N_21371);
xor U21656 (N_21656,N_21290,N_21408);
and U21657 (N_21657,N_21277,N_21423);
xor U21658 (N_21658,N_21483,N_21304);
and U21659 (N_21659,N_21439,N_21462);
or U21660 (N_21660,N_21478,N_21447);
nand U21661 (N_21661,N_21385,N_21465);
nand U21662 (N_21662,N_21366,N_21387);
and U21663 (N_21663,N_21478,N_21340);
nand U21664 (N_21664,N_21384,N_21280);
nand U21665 (N_21665,N_21379,N_21346);
nor U21666 (N_21666,N_21289,N_21463);
nor U21667 (N_21667,N_21263,N_21356);
and U21668 (N_21668,N_21449,N_21361);
and U21669 (N_21669,N_21358,N_21325);
nand U21670 (N_21670,N_21373,N_21331);
nor U21671 (N_21671,N_21403,N_21423);
nor U21672 (N_21672,N_21280,N_21480);
and U21673 (N_21673,N_21470,N_21379);
nand U21674 (N_21674,N_21435,N_21413);
and U21675 (N_21675,N_21463,N_21303);
xnor U21676 (N_21676,N_21362,N_21256);
nor U21677 (N_21677,N_21475,N_21328);
xnor U21678 (N_21678,N_21302,N_21269);
nor U21679 (N_21679,N_21456,N_21412);
nand U21680 (N_21680,N_21255,N_21478);
nor U21681 (N_21681,N_21481,N_21418);
and U21682 (N_21682,N_21374,N_21370);
nand U21683 (N_21683,N_21421,N_21390);
and U21684 (N_21684,N_21441,N_21444);
nor U21685 (N_21685,N_21250,N_21293);
nand U21686 (N_21686,N_21381,N_21461);
or U21687 (N_21687,N_21390,N_21370);
xnor U21688 (N_21688,N_21270,N_21313);
and U21689 (N_21689,N_21256,N_21425);
nand U21690 (N_21690,N_21407,N_21448);
and U21691 (N_21691,N_21254,N_21290);
and U21692 (N_21692,N_21342,N_21373);
and U21693 (N_21693,N_21343,N_21251);
nor U21694 (N_21694,N_21433,N_21342);
nand U21695 (N_21695,N_21363,N_21319);
or U21696 (N_21696,N_21423,N_21324);
and U21697 (N_21697,N_21327,N_21296);
nor U21698 (N_21698,N_21366,N_21258);
xnor U21699 (N_21699,N_21490,N_21402);
and U21700 (N_21700,N_21496,N_21351);
and U21701 (N_21701,N_21461,N_21429);
nor U21702 (N_21702,N_21293,N_21331);
nand U21703 (N_21703,N_21486,N_21402);
xor U21704 (N_21704,N_21443,N_21352);
and U21705 (N_21705,N_21284,N_21289);
or U21706 (N_21706,N_21343,N_21412);
xnor U21707 (N_21707,N_21348,N_21401);
nand U21708 (N_21708,N_21405,N_21276);
nand U21709 (N_21709,N_21456,N_21323);
nand U21710 (N_21710,N_21317,N_21370);
and U21711 (N_21711,N_21313,N_21428);
xnor U21712 (N_21712,N_21446,N_21336);
nand U21713 (N_21713,N_21449,N_21428);
and U21714 (N_21714,N_21484,N_21339);
or U21715 (N_21715,N_21275,N_21450);
nand U21716 (N_21716,N_21478,N_21496);
nand U21717 (N_21717,N_21339,N_21477);
and U21718 (N_21718,N_21342,N_21431);
or U21719 (N_21719,N_21480,N_21281);
xor U21720 (N_21720,N_21454,N_21383);
nor U21721 (N_21721,N_21301,N_21293);
or U21722 (N_21722,N_21258,N_21331);
or U21723 (N_21723,N_21468,N_21489);
and U21724 (N_21724,N_21378,N_21278);
and U21725 (N_21725,N_21344,N_21383);
xnor U21726 (N_21726,N_21317,N_21435);
and U21727 (N_21727,N_21449,N_21494);
and U21728 (N_21728,N_21300,N_21463);
nand U21729 (N_21729,N_21471,N_21285);
and U21730 (N_21730,N_21479,N_21254);
and U21731 (N_21731,N_21420,N_21492);
nor U21732 (N_21732,N_21462,N_21313);
nor U21733 (N_21733,N_21487,N_21333);
or U21734 (N_21734,N_21450,N_21428);
nor U21735 (N_21735,N_21455,N_21257);
or U21736 (N_21736,N_21346,N_21289);
and U21737 (N_21737,N_21413,N_21403);
and U21738 (N_21738,N_21293,N_21405);
nand U21739 (N_21739,N_21322,N_21467);
and U21740 (N_21740,N_21268,N_21344);
or U21741 (N_21741,N_21331,N_21386);
or U21742 (N_21742,N_21292,N_21342);
and U21743 (N_21743,N_21389,N_21342);
xnor U21744 (N_21744,N_21412,N_21251);
and U21745 (N_21745,N_21466,N_21492);
xor U21746 (N_21746,N_21286,N_21375);
or U21747 (N_21747,N_21261,N_21284);
or U21748 (N_21748,N_21356,N_21369);
nand U21749 (N_21749,N_21284,N_21385);
nand U21750 (N_21750,N_21650,N_21728);
xor U21751 (N_21751,N_21627,N_21501);
and U21752 (N_21752,N_21700,N_21500);
nand U21753 (N_21753,N_21600,N_21664);
or U21754 (N_21754,N_21692,N_21599);
nand U21755 (N_21755,N_21746,N_21682);
xor U21756 (N_21756,N_21542,N_21741);
xor U21757 (N_21757,N_21663,N_21503);
nor U21758 (N_21758,N_21506,N_21694);
or U21759 (N_21759,N_21584,N_21658);
xor U21760 (N_21760,N_21651,N_21634);
nand U21761 (N_21761,N_21720,N_21564);
xnor U21762 (N_21762,N_21705,N_21677);
nor U21763 (N_21763,N_21516,N_21613);
or U21764 (N_21764,N_21661,N_21563);
xnor U21765 (N_21765,N_21518,N_21646);
or U21766 (N_21766,N_21533,N_21534);
xor U21767 (N_21767,N_21696,N_21550);
nand U21768 (N_21768,N_21636,N_21541);
and U21769 (N_21769,N_21546,N_21617);
or U21770 (N_21770,N_21568,N_21504);
and U21771 (N_21771,N_21589,N_21675);
nor U21772 (N_21772,N_21510,N_21697);
nand U21773 (N_21773,N_21521,N_21668);
and U21774 (N_21774,N_21723,N_21610);
and U21775 (N_21775,N_21508,N_21565);
or U21776 (N_21776,N_21686,N_21555);
xnor U21777 (N_21777,N_21579,N_21570);
nand U21778 (N_21778,N_21666,N_21727);
xnor U21779 (N_21779,N_21638,N_21679);
nor U21780 (N_21780,N_21701,N_21711);
and U21781 (N_21781,N_21742,N_21558);
xor U21782 (N_21782,N_21595,N_21519);
and U21783 (N_21783,N_21545,N_21547);
or U21784 (N_21784,N_21706,N_21543);
and U21785 (N_21785,N_21721,N_21735);
xnor U21786 (N_21786,N_21591,N_21635);
nand U21787 (N_21787,N_21647,N_21652);
nor U21788 (N_21788,N_21608,N_21684);
or U21789 (N_21789,N_21590,N_21629);
nor U21790 (N_21790,N_21699,N_21637);
nor U21791 (N_21791,N_21580,N_21640);
nand U21792 (N_21792,N_21578,N_21687);
xor U21793 (N_21793,N_21683,N_21734);
xnor U21794 (N_21794,N_21562,N_21744);
or U21795 (N_21795,N_21515,N_21583);
or U21796 (N_21796,N_21581,N_21615);
xor U21797 (N_21797,N_21725,N_21669);
nor U21798 (N_21798,N_21645,N_21710);
xor U21799 (N_21799,N_21724,N_21674);
nand U21800 (N_21800,N_21601,N_21680);
or U21801 (N_21801,N_21719,N_21670);
or U21802 (N_21802,N_21618,N_21739);
nand U21803 (N_21803,N_21514,N_21525);
nor U21804 (N_21804,N_21616,N_21571);
nor U21805 (N_21805,N_21573,N_21737);
xor U21806 (N_21806,N_21609,N_21553);
xor U21807 (N_21807,N_21622,N_21530);
nor U21808 (N_21808,N_21604,N_21603);
nor U21809 (N_21809,N_21654,N_21569);
nor U21810 (N_21810,N_21585,N_21621);
nand U21811 (N_21811,N_21512,N_21690);
or U21812 (N_21812,N_21567,N_21517);
and U21813 (N_21813,N_21648,N_21633);
or U21814 (N_21814,N_21631,N_21540);
and U21815 (N_21815,N_21611,N_21641);
nand U21816 (N_21816,N_21743,N_21709);
or U21817 (N_21817,N_21531,N_21704);
or U21818 (N_21818,N_21537,N_21502);
nand U21819 (N_21819,N_21532,N_21703);
xor U21820 (N_21820,N_21596,N_21643);
nand U21821 (N_21821,N_21693,N_21556);
and U21822 (N_21822,N_21708,N_21747);
or U21823 (N_21823,N_21529,N_21691);
and U21824 (N_21824,N_21509,N_21740);
nor U21825 (N_21825,N_21527,N_21685);
or U21826 (N_21826,N_21730,N_21552);
xnor U21827 (N_21827,N_21653,N_21681);
nand U21828 (N_21828,N_21513,N_21507);
xnor U21829 (N_21829,N_21707,N_21718);
nor U21830 (N_21830,N_21729,N_21749);
or U21831 (N_21831,N_21524,N_21733);
and U21832 (N_21832,N_21625,N_21657);
nor U21833 (N_21833,N_21538,N_21598);
nand U21834 (N_21834,N_21726,N_21619);
or U21835 (N_21835,N_21695,N_21628);
xor U21836 (N_21836,N_21713,N_21522);
or U21837 (N_21837,N_21689,N_21660);
nand U21838 (N_21838,N_21574,N_21505);
nor U21839 (N_21839,N_21577,N_21548);
or U21840 (N_21840,N_21678,N_21597);
or U21841 (N_21841,N_21671,N_21702);
nor U21842 (N_21842,N_21535,N_21659);
nand U21843 (N_21843,N_21624,N_21536);
nor U21844 (N_21844,N_21560,N_21667);
nand U21845 (N_21845,N_21632,N_21566);
xnor U21846 (N_21846,N_21587,N_21626);
nor U21847 (N_21847,N_21717,N_21557);
or U21848 (N_21848,N_21586,N_21528);
and U21849 (N_21849,N_21594,N_21588);
nand U21850 (N_21850,N_21520,N_21593);
nand U21851 (N_21851,N_21712,N_21732);
nor U21852 (N_21852,N_21716,N_21551);
xnor U21853 (N_21853,N_21526,N_21575);
nand U21854 (N_21854,N_21642,N_21698);
and U21855 (N_21855,N_21549,N_21602);
nor U21856 (N_21856,N_21572,N_21605);
xor U21857 (N_21857,N_21715,N_21606);
nand U21858 (N_21858,N_21662,N_21665);
and U21859 (N_21859,N_21644,N_21673);
and U21860 (N_21860,N_21612,N_21614);
nor U21861 (N_21861,N_21592,N_21688);
or U21862 (N_21862,N_21576,N_21539);
xor U21863 (N_21863,N_21554,N_21544);
or U21864 (N_21864,N_21607,N_21620);
or U21865 (N_21865,N_21639,N_21649);
nor U21866 (N_21866,N_21523,N_21714);
or U21867 (N_21867,N_21748,N_21731);
or U21868 (N_21868,N_21672,N_21738);
xor U21869 (N_21869,N_21511,N_21745);
and U21870 (N_21870,N_21655,N_21582);
or U21871 (N_21871,N_21561,N_21623);
nand U21872 (N_21872,N_21722,N_21656);
nand U21873 (N_21873,N_21736,N_21559);
nor U21874 (N_21874,N_21676,N_21630);
or U21875 (N_21875,N_21555,N_21713);
and U21876 (N_21876,N_21506,N_21691);
or U21877 (N_21877,N_21578,N_21506);
and U21878 (N_21878,N_21730,N_21731);
nor U21879 (N_21879,N_21501,N_21598);
and U21880 (N_21880,N_21747,N_21674);
nand U21881 (N_21881,N_21700,N_21585);
nor U21882 (N_21882,N_21637,N_21733);
nand U21883 (N_21883,N_21748,N_21640);
nor U21884 (N_21884,N_21661,N_21558);
xnor U21885 (N_21885,N_21748,N_21725);
nor U21886 (N_21886,N_21606,N_21702);
or U21887 (N_21887,N_21581,N_21712);
and U21888 (N_21888,N_21679,N_21662);
or U21889 (N_21889,N_21505,N_21610);
nand U21890 (N_21890,N_21536,N_21596);
xor U21891 (N_21891,N_21709,N_21501);
nor U21892 (N_21892,N_21597,N_21635);
xnor U21893 (N_21893,N_21629,N_21707);
and U21894 (N_21894,N_21703,N_21560);
or U21895 (N_21895,N_21554,N_21530);
nand U21896 (N_21896,N_21511,N_21682);
nand U21897 (N_21897,N_21587,N_21710);
and U21898 (N_21898,N_21694,N_21636);
nor U21899 (N_21899,N_21683,N_21713);
xnor U21900 (N_21900,N_21676,N_21667);
or U21901 (N_21901,N_21747,N_21608);
nor U21902 (N_21902,N_21519,N_21591);
and U21903 (N_21903,N_21720,N_21741);
or U21904 (N_21904,N_21579,N_21664);
xor U21905 (N_21905,N_21504,N_21609);
and U21906 (N_21906,N_21638,N_21732);
xor U21907 (N_21907,N_21576,N_21611);
xnor U21908 (N_21908,N_21550,N_21538);
and U21909 (N_21909,N_21663,N_21576);
nand U21910 (N_21910,N_21591,N_21564);
nand U21911 (N_21911,N_21570,N_21621);
nand U21912 (N_21912,N_21592,N_21636);
xnor U21913 (N_21913,N_21558,N_21714);
nor U21914 (N_21914,N_21587,N_21662);
nand U21915 (N_21915,N_21730,N_21622);
or U21916 (N_21916,N_21621,N_21648);
xnor U21917 (N_21917,N_21507,N_21598);
or U21918 (N_21918,N_21685,N_21726);
or U21919 (N_21919,N_21578,N_21745);
or U21920 (N_21920,N_21553,N_21731);
xnor U21921 (N_21921,N_21738,N_21535);
xnor U21922 (N_21922,N_21647,N_21738);
nor U21923 (N_21923,N_21618,N_21726);
nor U21924 (N_21924,N_21625,N_21556);
and U21925 (N_21925,N_21522,N_21749);
nand U21926 (N_21926,N_21729,N_21747);
and U21927 (N_21927,N_21604,N_21742);
nand U21928 (N_21928,N_21623,N_21639);
nor U21929 (N_21929,N_21538,N_21675);
and U21930 (N_21930,N_21536,N_21631);
nand U21931 (N_21931,N_21513,N_21504);
nand U21932 (N_21932,N_21601,N_21525);
xor U21933 (N_21933,N_21613,N_21749);
and U21934 (N_21934,N_21683,N_21548);
nor U21935 (N_21935,N_21727,N_21550);
xor U21936 (N_21936,N_21656,N_21604);
or U21937 (N_21937,N_21541,N_21683);
and U21938 (N_21938,N_21631,N_21665);
nand U21939 (N_21939,N_21612,N_21742);
nand U21940 (N_21940,N_21559,N_21561);
nand U21941 (N_21941,N_21598,N_21658);
nand U21942 (N_21942,N_21552,N_21502);
nor U21943 (N_21943,N_21729,N_21557);
and U21944 (N_21944,N_21746,N_21580);
and U21945 (N_21945,N_21588,N_21739);
nor U21946 (N_21946,N_21646,N_21714);
nor U21947 (N_21947,N_21682,N_21506);
or U21948 (N_21948,N_21572,N_21731);
and U21949 (N_21949,N_21522,N_21626);
nor U21950 (N_21950,N_21709,N_21614);
nor U21951 (N_21951,N_21578,N_21603);
xnor U21952 (N_21952,N_21526,N_21589);
and U21953 (N_21953,N_21633,N_21572);
nand U21954 (N_21954,N_21507,N_21597);
nor U21955 (N_21955,N_21504,N_21543);
xor U21956 (N_21956,N_21708,N_21633);
nand U21957 (N_21957,N_21722,N_21512);
nor U21958 (N_21958,N_21731,N_21562);
and U21959 (N_21959,N_21665,N_21703);
nor U21960 (N_21960,N_21664,N_21739);
or U21961 (N_21961,N_21565,N_21631);
and U21962 (N_21962,N_21654,N_21599);
or U21963 (N_21963,N_21617,N_21672);
or U21964 (N_21964,N_21703,N_21589);
or U21965 (N_21965,N_21620,N_21733);
and U21966 (N_21966,N_21646,N_21717);
xor U21967 (N_21967,N_21617,N_21700);
nand U21968 (N_21968,N_21578,N_21729);
and U21969 (N_21969,N_21694,N_21556);
nor U21970 (N_21970,N_21632,N_21718);
nand U21971 (N_21971,N_21593,N_21533);
and U21972 (N_21972,N_21727,N_21672);
nand U21973 (N_21973,N_21602,N_21533);
nand U21974 (N_21974,N_21718,N_21738);
nand U21975 (N_21975,N_21512,N_21728);
nand U21976 (N_21976,N_21593,N_21713);
nor U21977 (N_21977,N_21681,N_21664);
and U21978 (N_21978,N_21519,N_21649);
nand U21979 (N_21979,N_21631,N_21686);
nand U21980 (N_21980,N_21749,N_21656);
nor U21981 (N_21981,N_21688,N_21672);
xnor U21982 (N_21982,N_21693,N_21596);
or U21983 (N_21983,N_21641,N_21716);
nand U21984 (N_21984,N_21691,N_21579);
nor U21985 (N_21985,N_21581,N_21598);
nor U21986 (N_21986,N_21728,N_21613);
xnor U21987 (N_21987,N_21709,N_21556);
nand U21988 (N_21988,N_21544,N_21584);
and U21989 (N_21989,N_21531,N_21516);
or U21990 (N_21990,N_21616,N_21708);
and U21991 (N_21991,N_21536,N_21591);
and U21992 (N_21992,N_21509,N_21610);
nor U21993 (N_21993,N_21639,N_21501);
xnor U21994 (N_21994,N_21659,N_21682);
and U21995 (N_21995,N_21514,N_21593);
and U21996 (N_21996,N_21645,N_21749);
or U21997 (N_21997,N_21733,N_21531);
and U21998 (N_21998,N_21521,N_21509);
and U21999 (N_21999,N_21603,N_21605);
or U22000 (N_22000,N_21980,N_21967);
nor U22001 (N_22001,N_21853,N_21795);
or U22002 (N_22002,N_21763,N_21971);
and U22003 (N_22003,N_21886,N_21864);
xnor U22004 (N_22004,N_21903,N_21920);
nand U22005 (N_22005,N_21919,N_21925);
or U22006 (N_22006,N_21805,N_21995);
nor U22007 (N_22007,N_21750,N_21895);
nand U22008 (N_22008,N_21817,N_21877);
xor U22009 (N_22009,N_21911,N_21969);
nor U22010 (N_22010,N_21944,N_21810);
and U22011 (N_22011,N_21922,N_21783);
and U22012 (N_22012,N_21801,N_21912);
xnor U22013 (N_22013,N_21751,N_21765);
nand U22014 (N_22014,N_21955,N_21803);
and U22015 (N_22015,N_21837,N_21844);
xor U22016 (N_22016,N_21927,N_21908);
xor U22017 (N_22017,N_21889,N_21834);
xor U22018 (N_22018,N_21959,N_21778);
xor U22019 (N_22019,N_21869,N_21981);
nand U22020 (N_22020,N_21999,N_21901);
and U22021 (N_22021,N_21949,N_21769);
xnor U22022 (N_22022,N_21825,N_21781);
xnor U22023 (N_22023,N_21946,N_21872);
xnor U22024 (N_22024,N_21868,N_21929);
nor U22025 (N_22025,N_21892,N_21887);
xnor U22026 (N_22026,N_21876,N_21900);
or U22027 (N_22027,N_21847,N_21790);
nor U22028 (N_22028,N_21994,N_21802);
and U22029 (N_22029,N_21815,N_21928);
xnor U22030 (N_22030,N_21830,N_21934);
or U22031 (N_22031,N_21983,N_21849);
or U22032 (N_22032,N_21857,N_21859);
xor U22033 (N_22033,N_21986,N_21996);
and U22034 (N_22034,N_21862,N_21968);
and U22035 (N_22035,N_21898,N_21807);
nand U22036 (N_22036,N_21880,N_21787);
nand U22037 (N_22037,N_21905,N_21829);
nand U22038 (N_22038,N_21914,N_21838);
xor U22039 (N_22039,N_21789,N_21854);
nor U22040 (N_22040,N_21873,N_21942);
nor U22041 (N_22041,N_21835,N_21962);
nor U22042 (N_22042,N_21773,N_21758);
or U22043 (N_22043,N_21757,N_21806);
xor U22044 (N_22044,N_21907,N_21970);
or U22045 (N_22045,N_21819,N_21800);
nor U22046 (N_22046,N_21867,N_21974);
nor U22047 (N_22047,N_21933,N_21948);
and U22048 (N_22048,N_21760,N_21842);
and U22049 (N_22049,N_21821,N_21976);
nor U22050 (N_22050,N_21784,N_21932);
or U22051 (N_22051,N_21952,N_21984);
nor U22052 (N_22052,N_21852,N_21828);
nand U22053 (N_22053,N_21866,N_21771);
xor U22054 (N_22054,N_21782,N_21754);
and U22055 (N_22055,N_21823,N_21973);
and U22056 (N_22056,N_21752,N_21899);
xnor U22057 (N_22057,N_21768,N_21776);
and U22058 (N_22058,N_21780,N_21924);
xor U22059 (N_22059,N_21833,N_21985);
nor U22060 (N_22060,N_21918,N_21858);
and U22061 (N_22061,N_21953,N_21788);
and U22062 (N_22062,N_21843,N_21965);
nand U22063 (N_22063,N_21909,N_21756);
xor U22064 (N_22064,N_21796,N_21961);
or U22065 (N_22065,N_21874,N_21824);
nor U22066 (N_22066,N_21972,N_21767);
xnor U22067 (N_22067,N_21964,N_21863);
nand U22068 (N_22068,N_21875,N_21989);
nor U22069 (N_22069,N_21786,N_21822);
and U22070 (N_22070,N_21982,N_21832);
or U22071 (N_22071,N_21910,N_21766);
nand U22072 (N_22072,N_21936,N_21755);
xnor U22073 (N_22073,N_21891,N_21861);
nor U22074 (N_22074,N_21761,N_21977);
and U22075 (N_22075,N_21960,N_21894);
xor U22076 (N_22076,N_21818,N_21935);
xor U22077 (N_22077,N_21906,N_21770);
and U22078 (N_22078,N_21890,N_21930);
and U22079 (N_22079,N_21947,N_21848);
xnor U22080 (N_22080,N_21855,N_21814);
or U22081 (N_22081,N_21978,N_21904);
or U22082 (N_22082,N_21772,N_21811);
nand U22083 (N_22083,N_21851,N_21826);
nor U22084 (N_22084,N_21988,N_21779);
and U22085 (N_22085,N_21958,N_21813);
and U22086 (N_22086,N_21804,N_21923);
and U22087 (N_22087,N_21812,N_21951);
nor U22088 (N_22088,N_21860,N_21884);
and U22089 (N_22089,N_21831,N_21992);
nor U22090 (N_22090,N_21841,N_21998);
and U22091 (N_22091,N_21997,N_21792);
and U22092 (N_22092,N_21839,N_21963);
nor U22093 (N_22093,N_21950,N_21915);
xnor U22094 (N_22094,N_21881,N_21856);
nand U22095 (N_22095,N_21975,N_21762);
or U22096 (N_22096,N_21870,N_21865);
xnor U22097 (N_22097,N_21836,N_21850);
nand U22098 (N_22098,N_21902,N_21871);
nor U22099 (N_22099,N_21979,N_21943);
or U22100 (N_22100,N_21827,N_21799);
or U22101 (N_22101,N_21939,N_21966);
and U22102 (N_22102,N_21764,N_21921);
and U22103 (N_22103,N_21809,N_21753);
and U22104 (N_22104,N_21785,N_21993);
and U22105 (N_22105,N_21845,N_21816);
nand U22106 (N_22106,N_21897,N_21940);
and U22107 (N_22107,N_21879,N_21885);
nor U22108 (N_22108,N_21937,N_21991);
or U22109 (N_22109,N_21794,N_21896);
nand U22110 (N_22110,N_21888,N_21820);
and U22111 (N_22111,N_21945,N_21846);
xor U22112 (N_22112,N_21941,N_21882);
and U22113 (N_22113,N_21883,N_21926);
nor U22114 (N_22114,N_21777,N_21954);
nor U22115 (N_22115,N_21987,N_21797);
xor U22116 (N_22116,N_21878,N_21798);
nand U22117 (N_22117,N_21793,N_21990);
nor U22118 (N_22118,N_21791,N_21956);
xor U22119 (N_22119,N_21931,N_21916);
nor U22120 (N_22120,N_21957,N_21808);
nor U22121 (N_22121,N_21913,N_21938);
nor U22122 (N_22122,N_21775,N_21840);
xor U22123 (N_22123,N_21893,N_21917);
and U22124 (N_22124,N_21774,N_21759);
nor U22125 (N_22125,N_21915,N_21828);
and U22126 (N_22126,N_21859,N_21751);
and U22127 (N_22127,N_21822,N_21836);
or U22128 (N_22128,N_21814,N_21897);
xnor U22129 (N_22129,N_21962,N_21956);
xor U22130 (N_22130,N_21800,N_21752);
xor U22131 (N_22131,N_21891,N_21756);
and U22132 (N_22132,N_21883,N_21756);
xor U22133 (N_22133,N_21920,N_21914);
nor U22134 (N_22134,N_21875,N_21891);
nand U22135 (N_22135,N_21801,N_21992);
or U22136 (N_22136,N_21776,N_21933);
nand U22137 (N_22137,N_21835,N_21815);
nand U22138 (N_22138,N_21891,N_21938);
and U22139 (N_22139,N_21898,N_21793);
nand U22140 (N_22140,N_21919,N_21933);
nand U22141 (N_22141,N_21893,N_21847);
nor U22142 (N_22142,N_21917,N_21786);
or U22143 (N_22143,N_21952,N_21756);
or U22144 (N_22144,N_21843,N_21880);
and U22145 (N_22145,N_21756,N_21865);
and U22146 (N_22146,N_21788,N_21950);
or U22147 (N_22147,N_21956,N_21991);
nand U22148 (N_22148,N_21925,N_21859);
nand U22149 (N_22149,N_21761,N_21876);
or U22150 (N_22150,N_21969,N_21940);
xnor U22151 (N_22151,N_21935,N_21913);
nor U22152 (N_22152,N_21803,N_21878);
or U22153 (N_22153,N_21831,N_21884);
xor U22154 (N_22154,N_21996,N_21982);
xnor U22155 (N_22155,N_21958,N_21887);
or U22156 (N_22156,N_21859,N_21839);
xor U22157 (N_22157,N_21972,N_21928);
and U22158 (N_22158,N_21778,N_21873);
nor U22159 (N_22159,N_21867,N_21933);
nand U22160 (N_22160,N_21910,N_21986);
or U22161 (N_22161,N_21872,N_21989);
and U22162 (N_22162,N_21990,N_21905);
nor U22163 (N_22163,N_21840,N_21918);
nor U22164 (N_22164,N_21768,N_21978);
and U22165 (N_22165,N_21924,N_21982);
nor U22166 (N_22166,N_21787,N_21890);
xor U22167 (N_22167,N_21782,N_21906);
xnor U22168 (N_22168,N_21998,N_21994);
xnor U22169 (N_22169,N_21921,N_21770);
and U22170 (N_22170,N_21769,N_21828);
xor U22171 (N_22171,N_21837,N_21804);
or U22172 (N_22172,N_21795,N_21845);
and U22173 (N_22173,N_21862,N_21781);
nand U22174 (N_22174,N_21956,N_21944);
or U22175 (N_22175,N_21886,N_21923);
nand U22176 (N_22176,N_21969,N_21977);
nor U22177 (N_22177,N_21884,N_21963);
and U22178 (N_22178,N_21941,N_21965);
nand U22179 (N_22179,N_21959,N_21819);
or U22180 (N_22180,N_21874,N_21983);
or U22181 (N_22181,N_21800,N_21755);
nor U22182 (N_22182,N_21978,N_21844);
and U22183 (N_22183,N_21997,N_21957);
or U22184 (N_22184,N_21753,N_21834);
or U22185 (N_22185,N_21841,N_21801);
nor U22186 (N_22186,N_21808,N_21900);
nor U22187 (N_22187,N_21836,N_21919);
nand U22188 (N_22188,N_21791,N_21858);
xor U22189 (N_22189,N_21856,N_21828);
nand U22190 (N_22190,N_21835,N_21915);
nor U22191 (N_22191,N_21812,N_21981);
nor U22192 (N_22192,N_21771,N_21803);
or U22193 (N_22193,N_21817,N_21780);
and U22194 (N_22194,N_21754,N_21900);
or U22195 (N_22195,N_21856,N_21911);
and U22196 (N_22196,N_21908,N_21843);
or U22197 (N_22197,N_21812,N_21873);
nand U22198 (N_22198,N_21977,N_21781);
nand U22199 (N_22199,N_21901,N_21987);
and U22200 (N_22200,N_21997,N_21867);
or U22201 (N_22201,N_21891,N_21951);
and U22202 (N_22202,N_21793,N_21930);
or U22203 (N_22203,N_21998,N_21925);
and U22204 (N_22204,N_21821,N_21943);
nand U22205 (N_22205,N_21895,N_21977);
or U22206 (N_22206,N_21967,N_21812);
or U22207 (N_22207,N_21875,N_21993);
and U22208 (N_22208,N_21763,N_21815);
nor U22209 (N_22209,N_21856,N_21919);
xnor U22210 (N_22210,N_21919,N_21862);
nor U22211 (N_22211,N_21889,N_21784);
and U22212 (N_22212,N_21875,N_21765);
nor U22213 (N_22213,N_21762,N_21974);
nand U22214 (N_22214,N_21839,N_21955);
or U22215 (N_22215,N_21833,N_21960);
nor U22216 (N_22216,N_21958,N_21891);
nor U22217 (N_22217,N_21954,N_21916);
nor U22218 (N_22218,N_21982,N_21799);
xnor U22219 (N_22219,N_21866,N_21954);
or U22220 (N_22220,N_21938,N_21932);
nor U22221 (N_22221,N_21890,N_21753);
xnor U22222 (N_22222,N_21777,N_21921);
and U22223 (N_22223,N_21863,N_21967);
or U22224 (N_22224,N_21926,N_21879);
xnor U22225 (N_22225,N_21966,N_21814);
xor U22226 (N_22226,N_21850,N_21964);
and U22227 (N_22227,N_21990,N_21975);
nor U22228 (N_22228,N_21895,N_21821);
nand U22229 (N_22229,N_21842,N_21985);
or U22230 (N_22230,N_21897,N_21982);
and U22231 (N_22231,N_21946,N_21910);
nor U22232 (N_22232,N_21757,N_21755);
nand U22233 (N_22233,N_21827,N_21858);
xor U22234 (N_22234,N_21982,N_21892);
and U22235 (N_22235,N_21806,N_21811);
nor U22236 (N_22236,N_21936,N_21932);
nand U22237 (N_22237,N_21997,N_21849);
xor U22238 (N_22238,N_21895,N_21941);
and U22239 (N_22239,N_21853,N_21868);
xnor U22240 (N_22240,N_21839,N_21910);
and U22241 (N_22241,N_21784,N_21956);
nand U22242 (N_22242,N_21942,N_21783);
or U22243 (N_22243,N_21873,N_21931);
and U22244 (N_22244,N_21768,N_21793);
nand U22245 (N_22245,N_21849,N_21888);
nor U22246 (N_22246,N_21860,N_21985);
xnor U22247 (N_22247,N_21914,N_21987);
xor U22248 (N_22248,N_21750,N_21933);
nor U22249 (N_22249,N_21823,N_21951);
xnor U22250 (N_22250,N_22038,N_22113);
nand U22251 (N_22251,N_22142,N_22068);
and U22252 (N_22252,N_22048,N_22001);
nor U22253 (N_22253,N_22059,N_22181);
and U22254 (N_22254,N_22117,N_22140);
nand U22255 (N_22255,N_22215,N_22209);
nand U22256 (N_22256,N_22018,N_22146);
and U22257 (N_22257,N_22096,N_22151);
nand U22258 (N_22258,N_22171,N_22021);
or U22259 (N_22259,N_22026,N_22029);
nand U22260 (N_22260,N_22226,N_22243);
or U22261 (N_22261,N_22086,N_22046);
xnor U22262 (N_22262,N_22075,N_22201);
xor U22263 (N_22263,N_22193,N_22164);
nand U22264 (N_22264,N_22237,N_22187);
xnor U22265 (N_22265,N_22159,N_22000);
and U22266 (N_22266,N_22074,N_22189);
or U22267 (N_22267,N_22139,N_22025);
and U22268 (N_22268,N_22121,N_22120);
and U22269 (N_22269,N_22114,N_22055);
nand U22270 (N_22270,N_22103,N_22248);
xor U22271 (N_22271,N_22175,N_22180);
nand U22272 (N_22272,N_22003,N_22172);
nand U22273 (N_22273,N_22112,N_22109);
and U22274 (N_22274,N_22101,N_22198);
nor U22275 (N_22275,N_22174,N_22110);
xor U22276 (N_22276,N_22182,N_22232);
and U22277 (N_22277,N_22061,N_22154);
nor U22278 (N_22278,N_22013,N_22153);
or U22279 (N_22279,N_22093,N_22083);
and U22280 (N_22280,N_22124,N_22242);
nand U22281 (N_22281,N_22145,N_22078);
xor U22282 (N_22282,N_22183,N_22168);
nor U22283 (N_22283,N_22091,N_22156);
nand U22284 (N_22284,N_22207,N_22123);
and U22285 (N_22285,N_22066,N_22245);
or U22286 (N_22286,N_22220,N_22058);
nor U22287 (N_22287,N_22130,N_22057);
xnor U22288 (N_22288,N_22213,N_22053);
nor U22289 (N_22289,N_22116,N_22167);
or U22290 (N_22290,N_22221,N_22197);
xor U22291 (N_22291,N_22014,N_22206);
or U22292 (N_22292,N_22065,N_22076);
and U22293 (N_22293,N_22227,N_22240);
xnor U22294 (N_22294,N_22234,N_22188);
nor U22295 (N_22295,N_22138,N_22104);
or U22296 (N_22296,N_22229,N_22235);
nand U22297 (N_22297,N_22119,N_22185);
and U22298 (N_22298,N_22081,N_22122);
nand U22299 (N_22299,N_22077,N_22158);
or U22300 (N_22300,N_22236,N_22202);
nor U22301 (N_22301,N_22196,N_22039);
xnor U22302 (N_22302,N_22070,N_22106);
and U22303 (N_22303,N_22247,N_22218);
nand U22304 (N_22304,N_22173,N_22143);
or U22305 (N_22305,N_22090,N_22099);
nor U22306 (N_22306,N_22085,N_22062);
or U22307 (N_22307,N_22246,N_22179);
or U22308 (N_22308,N_22073,N_22056);
or U22309 (N_22309,N_22087,N_22163);
and U22310 (N_22310,N_22203,N_22225);
or U22311 (N_22311,N_22233,N_22031);
nor U22312 (N_22312,N_22042,N_22052);
nand U22313 (N_22313,N_22088,N_22005);
or U22314 (N_22314,N_22214,N_22137);
or U22315 (N_22315,N_22222,N_22069);
or U22316 (N_22316,N_22148,N_22115);
or U22317 (N_22317,N_22244,N_22129);
nor U22318 (N_22318,N_22204,N_22043);
xnor U22319 (N_22319,N_22238,N_22002);
nor U22320 (N_22320,N_22060,N_22131);
or U22321 (N_22321,N_22210,N_22044);
nand U22322 (N_22322,N_22010,N_22064);
nor U22323 (N_22323,N_22249,N_22191);
xnor U22324 (N_22324,N_22105,N_22144);
xor U22325 (N_22325,N_22147,N_22212);
nand U22326 (N_22326,N_22040,N_22107);
or U22327 (N_22327,N_22133,N_22160);
or U22328 (N_22328,N_22155,N_22136);
nand U22329 (N_22329,N_22192,N_22027);
nand U22330 (N_22330,N_22205,N_22127);
and U22331 (N_22331,N_22230,N_22125);
xor U22332 (N_22332,N_22016,N_22012);
nor U22333 (N_22333,N_22080,N_22011);
nand U22334 (N_22334,N_22132,N_22186);
or U22335 (N_22335,N_22071,N_22111);
or U22336 (N_22336,N_22211,N_22035);
and U22337 (N_22337,N_22200,N_22092);
or U22338 (N_22338,N_22007,N_22184);
nor U22339 (N_22339,N_22228,N_22047);
nor U22340 (N_22340,N_22084,N_22100);
and U22341 (N_22341,N_22161,N_22030);
xnor U22342 (N_22342,N_22223,N_22176);
xor U22343 (N_22343,N_22195,N_22208);
xor U22344 (N_22344,N_22022,N_22063);
or U22345 (N_22345,N_22241,N_22045);
xnor U22346 (N_22346,N_22162,N_22128);
xor U22347 (N_22347,N_22067,N_22165);
xnor U22348 (N_22348,N_22141,N_22082);
nor U22349 (N_22349,N_22008,N_22149);
xor U22350 (N_22350,N_22004,N_22023);
nand U22351 (N_22351,N_22006,N_22054);
and U22352 (N_22352,N_22019,N_22152);
nor U22353 (N_22353,N_22095,N_22102);
nand U22354 (N_22354,N_22034,N_22169);
xor U22355 (N_22355,N_22177,N_22009);
xor U22356 (N_22356,N_22072,N_22015);
and U22357 (N_22357,N_22178,N_22089);
nor U22358 (N_22358,N_22051,N_22135);
nand U22359 (N_22359,N_22032,N_22134);
and U22360 (N_22360,N_22079,N_22219);
xnor U22361 (N_22361,N_22041,N_22097);
nand U22362 (N_22362,N_22239,N_22118);
nand U22363 (N_22363,N_22020,N_22050);
xnor U22364 (N_22364,N_22098,N_22166);
or U22365 (N_22365,N_22224,N_22126);
nand U22366 (N_22366,N_22049,N_22028);
xor U22367 (N_22367,N_22150,N_22217);
nor U22368 (N_22368,N_22017,N_22216);
or U22369 (N_22369,N_22037,N_22108);
nor U22370 (N_22370,N_22033,N_22231);
or U22371 (N_22371,N_22024,N_22199);
nor U22372 (N_22372,N_22170,N_22194);
nor U22373 (N_22373,N_22036,N_22094);
nand U22374 (N_22374,N_22190,N_22157);
or U22375 (N_22375,N_22036,N_22016);
xor U22376 (N_22376,N_22207,N_22152);
and U22377 (N_22377,N_22011,N_22083);
nand U22378 (N_22378,N_22167,N_22078);
nand U22379 (N_22379,N_22061,N_22249);
nor U22380 (N_22380,N_22073,N_22160);
nand U22381 (N_22381,N_22235,N_22224);
or U22382 (N_22382,N_22128,N_22217);
nor U22383 (N_22383,N_22095,N_22019);
nor U22384 (N_22384,N_22095,N_22163);
nor U22385 (N_22385,N_22166,N_22225);
and U22386 (N_22386,N_22166,N_22094);
or U22387 (N_22387,N_22225,N_22219);
xor U22388 (N_22388,N_22186,N_22036);
or U22389 (N_22389,N_22167,N_22082);
and U22390 (N_22390,N_22119,N_22183);
nor U22391 (N_22391,N_22025,N_22101);
nand U22392 (N_22392,N_22171,N_22223);
nor U22393 (N_22393,N_22104,N_22083);
nand U22394 (N_22394,N_22187,N_22017);
nand U22395 (N_22395,N_22040,N_22227);
and U22396 (N_22396,N_22075,N_22244);
nand U22397 (N_22397,N_22246,N_22193);
xor U22398 (N_22398,N_22008,N_22164);
nand U22399 (N_22399,N_22176,N_22094);
and U22400 (N_22400,N_22107,N_22131);
xor U22401 (N_22401,N_22196,N_22080);
and U22402 (N_22402,N_22139,N_22114);
and U22403 (N_22403,N_22154,N_22053);
nor U22404 (N_22404,N_22193,N_22100);
or U22405 (N_22405,N_22141,N_22197);
nor U22406 (N_22406,N_22077,N_22239);
nor U22407 (N_22407,N_22069,N_22130);
or U22408 (N_22408,N_22224,N_22170);
xnor U22409 (N_22409,N_22102,N_22120);
xnor U22410 (N_22410,N_22101,N_22033);
and U22411 (N_22411,N_22000,N_22247);
xor U22412 (N_22412,N_22118,N_22219);
nand U22413 (N_22413,N_22219,N_22213);
or U22414 (N_22414,N_22152,N_22161);
nor U22415 (N_22415,N_22163,N_22143);
and U22416 (N_22416,N_22080,N_22010);
or U22417 (N_22417,N_22044,N_22246);
xnor U22418 (N_22418,N_22247,N_22186);
and U22419 (N_22419,N_22065,N_22057);
and U22420 (N_22420,N_22172,N_22224);
xor U22421 (N_22421,N_22187,N_22002);
nand U22422 (N_22422,N_22198,N_22242);
nand U22423 (N_22423,N_22122,N_22151);
or U22424 (N_22424,N_22043,N_22154);
nand U22425 (N_22425,N_22074,N_22154);
xor U22426 (N_22426,N_22120,N_22157);
or U22427 (N_22427,N_22236,N_22138);
and U22428 (N_22428,N_22181,N_22246);
nor U22429 (N_22429,N_22008,N_22133);
nor U22430 (N_22430,N_22220,N_22031);
xnor U22431 (N_22431,N_22198,N_22009);
xor U22432 (N_22432,N_22199,N_22167);
or U22433 (N_22433,N_22209,N_22028);
xnor U22434 (N_22434,N_22063,N_22092);
nor U22435 (N_22435,N_22051,N_22245);
and U22436 (N_22436,N_22062,N_22226);
and U22437 (N_22437,N_22045,N_22099);
and U22438 (N_22438,N_22096,N_22199);
nand U22439 (N_22439,N_22065,N_22009);
or U22440 (N_22440,N_22088,N_22222);
or U22441 (N_22441,N_22079,N_22191);
nand U22442 (N_22442,N_22211,N_22046);
or U22443 (N_22443,N_22193,N_22021);
xor U22444 (N_22444,N_22016,N_22171);
nor U22445 (N_22445,N_22127,N_22154);
nand U22446 (N_22446,N_22175,N_22137);
xnor U22447 (N_22447,N_22083,N_22102);
or U22448 (N_22448,N_22024,N_22118);
or U22449 (N_22449,N_22026,N_22010);
nand U22450 (N_22450,N_22170,N_22102);
nor U22451 (N_22451,N_22039,N_22160);
xnor U22452 (N_22452,N_22225,N_22043);
and U22453 (N_22453,N_22176,N_22215);
and U22454 (N_22454,N_22143,N_22184);
nand U22455 (N_22455,N_22059,N_22097);
nor U22456 (N_22456,N_22090,N_22147);
xor U22457 (N_22457,N_22071,N_22023);
xnor U22458 (N_22458,N_22120,N_22057);
nand U22459 (N_22459,N_22023,N_22215);
nand U22460 (N_22460,N_22186,N_22239);
nor U22461 (N_22461,N_22173,N_22202);
xor U22462 (N_22462,N_22196,N_22059);
nand U22463 (N_22463,N_22016,N_22052);
or U22464 (N_22464,N_22216,N_22180);
xnor U22465 (N_22465,N_22067,N_22248);
nand U22466 (N_22466,N_22012,N_22061);
nand U22467 (N_22467,N_22026,N_22028);
nand U22468 (N_22468,N_22111,N_22097);
nor U22469 (N_22469,N_22020,N_22010);
and U22470 (N_22470,N_22119,N_22147);
or U22471 (N_22471,N_22243,N_22069);
nor U22472 (N_22472,N_22130,N_22243);
nand U22473 (N_22473,N_22184,N_22181);
nor U22474 (N_22474,N_22048,N_22241);
or U22475 (N_22475,N_22019,N_22028);
nand U22476 (N_22476,N_22179,N_22166);
nand U22477 (N_22477,N_22159,N_22160);
nor U22478 (N_22478,N_22194,N_22066);
or U22479 (N_22479,N_22164,N_22188);
nand U22480 (N_22480,N_22008,N_22136);
nand U22481 (N_22481,N_22056,N_22174);
and U22482 (N_22482,N_22221,N_22209);
nand U22483 (N_22483,N_22138,N_22109);
xnor U22484 (N_22484,N_22037,N_22120);
nor U22485 (N_22485,N_22180,N_22150);
or U22486 (N_22486,N_22178,N_22032);
nor U22487 (N_22487,N_22103,N_22073);
or U22488 (N_22488,N_22114,N_22059);
and U22489 (N_22489,N_22031,N_22171);
nand U22490 (N_22490,N_22078,N_22097);
or U22491 (N_22491,N_22192,N_22066);
nand U22492 (N_22492,N_22039,N_22154);
and U22493 (N_22493,N_22242,N_22176);
nand U22494 (N_22494,N_22218,N_22141);
and U22495 (N_22495,N_22175,N_22085);
and U22496 (N_22496,N_22114,N_22024);
nand U22497 (N_22497,N_22072,N_22180);
and U22498 (N_22498,N_22211,N_22094);
and U22499 (N_22499,N_22196,N_22218);
nand U22500 (N_22500,N_22430,N_22497);
nor U22501 (N_22501,N_22406,N_22384);
and U22502 (N_22502,N_22401,N_22467);
nor U22503 (N_22503,N_22433,N_22268);
nor U22504 (N_22504,N_22456,N_22377);
xnor U22505 (N_22505,N_22445,N_22293);
xnor U22506 (N_22506,N_22319,N_22416);
xnor U22507 (N_22507,N_22251,N_22345);
xor U22508 (N_22508,N_22465,N_22343);
nand U22509 (N_22509,N_22302,N_22423);
xor U22510 (N_22510,N_22470,N_22352);
nor U22511 (N_22511,N_22420,N_22386);
or U22512 (N_22512,N_22385,N_22476);
and U22513 (N_22513,N_22388,N_22375);
and U22514 (N_22514,N_22298,N_22295);
nor U22515 (N_22515,N_22400,N_22483);
xnor U22516 (N_22516,N_22273,N_22276);
and U22517 (N_22517,N_22315,N_22362);
nand U22518 (N_22518,N_22279,N_22370);
nor U22519 (N_22519,N_22374,N_22355);
nand U22520 (N_22520,N_22324,N_22277);
nor U22521 (N_22521,N_22414,N_22421);
or U22522 (N_22522,N_22429,N_22307);
and U22523 (N_22523,N_22346,N_22264);
nor U22524 (N_22524,N_22335,N_22284);
or U22525 (N_22525,N_22272,N_22418);
nand U22526 (N_22526,N_22359,N_22271);
or U22527 (N_22527,N_22487,N_22457);
or U22528 (N_22528,N_22296,N_22441);
nand U22529 (N_22529,N_22313,N_22321);
nand U22530 (N_22530,N_22468,N_22274);
or U22531 (N_22531,N_22287,N_22499);
and U22532 (N_22532,N_22305,N_22495);
nand U22533 (N_22533,N_22297,N_22455);
and U22534 (N_22534,N_22471,N_22344);
nor U22535 (N_22535,N_22444,N_22327);
nand U22536 (N_22536,N_22435,N_22424);
or U22537 (N_22537,N_22283,N_22338);
nor U22538 (N_22538,N_22451,N_22267);
nand U22539 (N_22539,N_22348,N_22481);
nor U22540 (N_22540,N_22411,N_22285);
and U22541 (N_22541,N_22387,N_22383);
and U22542 (N_22542,N_22361,N_22312);
or U22543 (N_22543,N_22294,N_22360);
xor U22544 (N_22544,N_22265,N_22378);
nand U22545 (N_22545,N_22405,N_22252);
nor U22546 (N_22546,N_22309,N_22341);
nor U22547 (N_22547,N_22316,N_22395);
and U22548 (N_22548,N_22280,N_22475);
nand U22549 (N_22549,N_22389,N_22261);
or U22550 (N_22550,N_22270,N_22317);
and U22551 (N_22551,N_22437,N_22320);
xnor U22552 (N_22552,N_22301,N_22308);
nand U22553 (N_22553,N_22484,N_22492);
or U22554 (N_22554,N_22460,N_22459);
xnor U22555 (N_22555,N_22336,N_22478);
and U22556 (N_22556,N_22286,N_22466);
and U22557 (N_22557,N_22486,N_22480);
and U22558 (N_22558,N_22402,N_22376);
and U22559 (N_22559,N_22407,N_22256);
xor U22560 (N_22560,N_22263,N_22454);
and U22561 (N_22561,N_22303,N_22472);
nand U22562 (N_22562,N_22432,N_22282);
nor U22563 (N_22563,N_22419,N_22477);
nor U22564 (N_22564,N_22381,N_22371);
and U22565 (N_22565,N_22431,N_22289);
xor U22566 (N_22566,N_22390,N_22314);
and U22567 (N_22567,N_22448,N_22469);
nor U22568 (N_22568,N_22258,N_22417);
nor U22569 (N_22569,N_22290,N_22250);
nand U22570 (N_22570,N_22413,N_22447);
nor U22571 (N_22571,N_22255,N_22372);
xnor U22572 (N_22572,N_22439,N_22422);
xor U22573 (N_22573,N_22408,N_22349);
nand U22574 (N_22574,N_22334,N_22354);
or U22575 (N_22575,N_22412,N_22329);
nand U22576 (N_22576,N_22260,N_22365);
nand U22577 (N_22577,N_22485,N_22496);
or U22578 (N_22578,N_22398,N_22452);
and U22579 (N_22579,N_22373,N_22382);
or U22580 (N_22580,N_22333,N_22392);
nand U22581 (N_22581,N_22356,N_22328);
xor U22582 (N_22582,N_22325,N_22489);
nor U22583 (N_22583,N_22369,N_22288);
xnor U22584 (N_22584,N_22266,N_22330);
xor U22585 (N_22585,N_22403,N_22347);
xor U22586 (N_22586,N_22391,N_22351);
and U22587 (N_22587,N_22350,N_22253);
xnor U22588 (N_22588,N_22326,N_22306);
xor U22589 (N_22589,N_22443,N_22257);
nand U22590 (N_22590,N_22438,N_22453);
nor U22591 (N_22591,N_22310,N_22363);
nand U22592 (N_22592,N_22458,N_22463);
nor U22593 (N_22593,N_22462,N_22357);
or U22594 (N_22594,N_22300,N_22269);
or U22595 (N_22595,N_22342,N_22474);
nand U22596 (N_22596,N_22259,N_22366);
or U22597 (N_22597,N_22323,N_22367);
and U22598 (N_22598,N_22380,N_22358);
nand U22599 (N_22599,N_22482,N_22493);
nand U22600 (N_22600,N_22353,N_22331);
and U22601 (N_22601,N_22396,N_22337);
or U22602 (N_22602,N_22473,N_22461);
or U22603 (N_22603,N_22488,N_22434);
or U22604 (N_22604,N_22339,N_22449);
xor U22605 (N_22605,N_22368,N_22275);
nor U22606 (N_22606,N_22364,N_22446);
nor U22607 (N_22607,N_22410,N_22393);
or U22608 (N_22608,N_22464,N_22254);
nor U22609 (N_22609,N_22404,N_22427);
and U22610 (N_22610,N_22399,N_22262);
or U22611 (N_22611,N_22426,N_22278);
xnor U22612 (N_22612,N_22425,N_22440);
or U22613 (N_22613,N_22428,N_22397);
or U22614 (N_22614,N_22491,N_22379);
xor U22615 (N_22615,N_22450,N_22479);
nor U22616 (N_22616,N_22409,N_22415);
nand U22617 (N_22617,N_22436,N_22311);
nand U22618 (N_22618,N_22490,N_22494);
nor U22619 (N_22619,N_22340,N_22318);
nand U22620 (N_22620,N_22442,N_22292);
or U22621 (N_22621,N_22304,N_22322);
or U22622 (N_22622,N_22291,N_22394);
and U22623 (N_22623,N_22498,N_22281);
nor U22624 (N_22624,N_22332,N_22299);
or U22625 (N_22625,N_22340,N_22351);
xor U22626 (N_22626,N_22275,N_22421);
and U22627 (N_22627,N_22412,N_22333);
nand U22628 (N_22628,N_22256,N_22325);
or U22629 (N_22629,N_22339,N_22363);
nand U22630 (N_22630,N_22370,N_22301);
nand U22631 (N_22631,N_22290,N_22377);
or U22632 (N_22632,N_22427,N_22340);
and U22633 (N_22633,N_22388,N_22426);
and U22634 (N_22634,N_22374,N_22440);
nand U22635 (N_22635,N_22281,N_22443);
xor U22636 (N_22636,N_22389,N_22329);
and U22637 (N_22637,N_22265,N_22337);
xnor U22638 (N_22638,N_22375,N_22279);
nor U22639 (N_22639,N_22362,N_22330);
nor U22640 (N_22640,N_22429,N_22367);
nand U22641 (N_22641,N_22406,N_22409);
and U22642 (N_22642,N_22275,N_22498);
xor U22643 (N_22643,N_22285,N_22260);
nand U22644 (N_22644,N_22253,N_22382);
xor U22645 (N_22645,N_22498,N_22373);
xor U22646 (N_22646,N_22381,N_22410);
or U22647 (N_22647,N_22461,N_22293);
or U22648 (N_22648,N_22458,N_22378);
xnor U22649 (N_22649,N_22486,N_22339);
nand U22650 (N_22650,N_22493,N_22275);
or U22651 (N_22651,N_22365,N_22405);
or U22652 (N_22652,N_22432,N_22490);
or U22653 (N_22653,N_22467,N_22289);
nor U22654 (N_22654,N_22307,N_22367);
nor U22655 (N_22655,N_22453,N_22263);
or U22656 (N_22656,N_22385,N_22269);
or U22657 (N_22657,N_22293,N_22337);
or U22658 (N_22658,N_22312,N_22435);
and U22659 (N_22659,N_22368,N_22252);
nand U22660 (N_22660,N_22430,N_22496);
nand U22661 (N_22661,N_22369,N_22392);
xor U22662 (N_22662,N_22303,N_22325);
xnor U22663 (N_22663,N_22303,N_22342);
nor U22664 (N_22664,N_22374,N_22390);
and U22665 (N_22665,N_22308,N_22441);
nand U22666 (N_22666,N_22405,N_22436);
nor U22667 (N_22667,N_22405,N_22364);
and U22668 (N_22668,N_22448,N_22425);
and U22669 (N_22669,N_22326,N_22392);
or U22670 (N_22670,N_22349,N_22338);
and U22671 (N_22671,N_22406,N_22349);
nor U22672 (N_22672,N_22272,N_22253);
xor U22673 (N_22673,N_22328,N_22467);
xor U22674 (N_22674,N_22251,N_22436);
and U22675 (N_22675,N_22251,N_22382);
nand U22676 (N_22676,N_22447,N_22264);
xnor U22677 (N_22677,N_22297,N_22284);
xor U22678 (N_22678,N_22421,N_22278);
and U22679 (N_22679,N_22330,N_22284);
or U22680 (N_22680,N_22270,N_22363);
and U22681 (N_22681,N_22498,N_22371);
or U22682 (N_22682,N_22359,N_22263);
nor U22683 (N_22683,N_22354,N_22273);
nor U22684 (N_22684,N_22258,N_22486);
nand U22685 (N_22685,N_22340,N_22415);
or U22686 (N_22686,N_22489,N_22477);
or U22687 (N_22687,N_22391,N_22472);
or U22688 (N_22688,N_22395,N_22317);
or U22689 (N_22689,N_22427,N_22489);
and U22690 (N_22690,N_22283,N_22259);
xnor U22691 (N_22691,N_22289,N_22386);
and U22692 (N_22692,N_22265,N_22452);
nand U22693 (N_22693,N_22386,N_22434);
nor U22694 (N_22694,N_22287,N_22414);
xor U22695 (N_22695,N_22474,N_22280);
xnor U22696 (N_22696,N_22310,N_22452);
xnor U22697 (N_22697,N_22332,N_22259);
xnor U22698 (N_22698,N_22380,N_22302);
nor U22699 (N_22699,N_22310,N_22319);
and U22700 (N_22700,N_22359,N_22495);
nand U22701 (N_22701,N_22390,N_22391);
nand U22702 (N_22702,N_22295,N_22387);
nor U22703 (N_22703,N_22367,N_22283);
or U22704 (N_22704,N_22334,N_22309);
nor U22705 (N_22705,N_22251,N_22283);
xnor U22706 (N_22706,N_22450,N_22414);
xor U22707 (N_22707,N_22489,N_22483);
xnor U22708 (N_22708,N_22431,N_22285);
nand U22709 (N_22709,N_22327,N_22437);
xnor U22710 (N_22710,N_22458,N_22372);
xor U22711 (N_22711,N_22420,N_22382);
xor U22712 (N_22712,N_22304,N_22417);
nand U22713 (N_22713,N_22422,N_22262);
or U22714 (N_22714,N_22273,N_22326);
nand U22715 (N_22715,N_22426,N_22428);
nand U22716 (N_22716,N_22428,N_22323);
nor U22717 (N_22717,N_22367,N_22462);
xnor U22718 (N_22718,N_22267,N_22279);
nand U22719 (N_22719,N_22254,N_22457);
nand U22720 (N_22720,N_22352,N_22332);
nand U22721 (N_22721,N_22411,N_22335);
xnor U22722 (N_22722,N_22497,N_22346);
xor U22723 (N_22723,N_22284,N_22371);
nor U22724 (N_22724,N_22479,N_22408);
xnor U22725 (N_22725,N_22414,N_22259);
xnor U22726 (N_22726,N_22499,N_22477);
nand U22727 (N_22727,N_22429,N_22296);
or U22728 (N_22728,N_22460,N_22322);
nor U22729 (N_22729,N_22447,N_22407);
nor U22730 (N_22730,N_22450,N_22261);
nor U22731 (N_22731,N_22416,N_22252);
nand U22732 (N_22732,N_22372,N_22278);
and U22733 (N_22733,N_22442,N_22402);
nand U22734 (N_22734,N_22484,N_22270);
nor U22735 (N_22735,N_22492,N_22289);
xnor U22736 (N_22736,N_22398,N_22488);
nand U22737 (N_22737,N_22409,N_22493);
xnor U22738 (N_22738,N_22365,N_22324);
or U22739 (N_22739,N_22453,N_22306);
nor U22740 (N_22740,N_22433,N_22392);
nor U22741 (N_22741,N_22369,N_22318);
xnor U22742 (N_22742,N_22310,N_22494);
or U22743 (N_22743,N_22462,N_22477);
and U22744 (N_22744,N_22264,N_22355);
xor U22745 (N_22745,N_22342,N_22480);
and U22746 (N_22746,N_22300,N_22371);
nor U22747 (N_22747,N_22494,N_22314);
xor U22748 (N_22748,N_22362,N_22269);
xor U22749 (N_22749,N_22382,N_22426);
nand U22750 (N_22750,N_22538,N_22707);
xor U22751 (N_22751,N_22719,N_22599);
xnor U22752 (N_22752,N_22747,N_22603);
nor U22753 (N_22753,N_22665,N_22597);
nand U22754 (N_22754,N_22674,N_22559);
or U22755 (N_22755,N_22574,N_22615);
nand U22756 (N_22756,N_22726,N_22557);
or U22757 (N_22757,N_22681,N_22701);
xnor U22758 (N_22758,N_22589,N_22714);
xnor U22759 (N_22759,N_22717,N_22667);
nor U22760 (N_22760,N_22639,N_22725);
nor U22761 (N_22761,N_22602,N_22541);
nor U22762 (N_22762,N_22694,N_22700);
or U22763 (N_22763,N_22630,N_22676);
nand U22764 (N_22764,N_22572,N_22678);
nor U22765 (N_22765,N_22688,N_22735);
nand U22766 (N_22766,N_22617,N_22584);
or U22767 (N_22767,N_22518,N_22622);
and U22768 (N_22768,N_22739,N_22661);
nand U22769 (N_22769,N_22643,N_22534);
xor U22770 (N_22770,N_22675,N_22660);
and U22771 (N_22771,N_22601,N_22659);
xor U22772 (N_22772,N_22642,N_22501);
xor U22773 (N_22773,N_22586,N_22535);
xor U22774 (N_22774,N_22621,N_22682);
or U22775 (N_22775,N_22712,N_22690);
xor U22776 (N_22776,N_22632,N_22656);
or U22777 (N_22777,N_22608,N_22531);
or U22778 (N_22778,N_22598,N_22703);
nand U22779 (N_22779,N_22588,N_22595);
xor U22780 (N_22780,N_22724,N_22650);
xnor U22781 (N_22781,N_22552,N_22649);
nor U22782 (N_22782,N_22610,N_22540);
or U22783 (N_22783,N_22549,N_22663);
and U22784 (N_22784,N_22502,N_22532);
nor U22785 (N_22785,N_22748,N_22685);
nor U22786 (N_22786,N_22503,N_22715);
and U22787 (N_22787,N_22723,N_22583);
or U22788 (N_22788,N_22525,N_22738);
nand U22789 (N_22789,N_22593,N_22514);
nor U22790 (N_22790,N_22744,N_22569);
nor U22791 (N_22791,N_22580,N_22628);
nand U22792 (N_22792,N_22594,N_22516);
and U22793 (N_22793,N_22728,N_22507);
nand U22794 (N_22794,N_22536,N_22581);
xnor U22795 (N_22795,N_22737,N_22533);
nor U22796 (N_22796,N_22616,N_22528);
nor U22797 (N_22797,N_22582,N_22670);
nor U22798 (N_22798,N_22696,N_22713);
nor U22799 (N_22799,N_22560,N_22691);
or U22800 (N_22800,N_22699,N_22671);
nand U22801 (N_22801,N_22596,N_22504);
nor U22802 (N_22802,N_22524,N_22645);
or U22803 (N_22803,N_22606,N_22526);
nand U22804 (N_22804,N_22658,N_22539);
xnor U22805 (N_22805,N_22720,N_22657);
nor U22806 (N_22806,N_22637,N_22677);
and U22807 (N_22807,N_22565,N_22508);
nand U22808 (N_22808,N_22662,N_22687);
nor U22809 (N_22809,N_22679,N_22561);
nand U22810 (N_22810,N_22500,N_22544);
and U22811 (N_22811,N_22579,N_22578);
and U22812 (N_22812,N_22668,N_22710);
or U22813 (N_22813,N_22680,N_22548);
nand U22814 (N_22814,N_22545,N_22550);
or U22815 (N_22815,N_22689,N_22631);
and U22816 (N_22816,N_22666,N_22510);
nor U22817 (N_22817,N_22730,N_22566);
or U22818 (N_22818,N_22743,N_22695);
and U22819 (N_22819,N_22709,N_22587);
xnor U22820 (N_22820,N_22556,N_22722);
nor U22821 (N_22821,N_22612,N_22519);
nand U22822 (N_22822,N_22605,N_22635);
nand U22823 (N_22823,N_22530,N_22633);
or U22824 (N_22824,N_22692,N_22734);
and U22825 (N_22825,N_22537,N_22638);
nand U22826 (N_22826,N_22651,N_22506);
and U22827 (N_22827,N_22664,N_22693);
and U22828 (N_22828,N_22505,N_22686);
and U22829 (N_22829,N_22527,N_22563);
nor U22830 (N_22830,N_22729,N_22684);
xor U22831 (N_22831,N_22646,N_22577);
and U22832 (N_22832,N_22513,N_22623);
xor U22833 (N_22833,N_22547,N_22585);
xnor U22834 (N_22834,N_22555,N_22512);
or U22835 (N_22835,N_22620,N_22683);
and U22836 (N_22836,N_22740,N_22607);
xor U22837 (N_22837,N_22626,N_22745);
nor U22838 (N_22838,N_22613,N_22716);
and U22839 (N_22839,N_22641,N_22571);
or U22840 (N_22840,N_22522,N_22749);
nand U22841 (N_22841,N_22564,N_22543);
nor U22842 (N_22842,N_22672,N_22509);
nand U22843 (N_22843,N_22746,N_22542);
or U22844 (N_22844,N_22721,N_22570);
and U22845 (N_22845,N_22611,N_22708);
nor U22846 (N_22846,N_22551,N_22647);
or U22847 (N_22847,N_22697,N_22733);
xnor U22848 (N_22848,N_22629,N_22614);
nand U22849 (N_22849,N_22648,N_22634);
xor U22850 (N_22850,N_22640,N_22736);
and U22851 (N_22851,N_22627,N_22576);
xor U22852 (N_22852,N_22573,N_22625);
xnor U22853 (N_22853,N_22673,N_22704);
and U22854 (N_22854,N_22702,N_22529);
nor U22855 (N_22855,N_22705,N_22520);
and U22856 (N_22856,N_22609,N_22567);
xnor U22857 (N_22857,N_22523,N_22592);
nor U22858 (N_22858,N_22742,N_22652);
and U22859 (N_22859,N_22618,N_22653);
or U22860 (N_22860,N_22590,N_22521);
xor U22861 (N_22861,N_22562,N_22558);
nand U22862 (N_22862,N_22600,N_22636);
nand U22863 (N_22863,N_22706,N_22718);
or U22864 (N_22864,N_22741,N_22575);
xnor U22865 (N_22865,N_22711,N_22553);
and U22866 (N_22866,N_22554,N_22591);
nand U22867 (N_22867,N_22619,N_22669);
and U22868 (N_22868,N_22624,N_22654);
xnor U22869 (N_22869,N_22515,N_22604);
or U22870 (N_22870,N_22698,N_22731);
xor U22871 (N_22871,N_22511,N_22546);
or U22872 (N_22872,N_22568,N_22727);
nand U22873 (N_22873,N_22517,N_22732);
nand U22874 (N_22874,N_22644,N_22655);
nor U22875 (N_22875,N_22502,N_22681);
or U22876 (N_22876,N_22550,N_22640);
nor U22877 (N_22877,N_22609,N_22738);
or U22878 (N_22878,N_22723,N_22652);
xnor U22879 (N_22879,N_22647,N_22652);
nand U22880 (N_22880,N_22686,N_22749);
nand U22881 (N_22881,N_22512,N_22513);
and U22882 (N_22882,N_22622,N_22510);
xor U22883 (N_22883,N_22580,N_22656);
nand U22884 (N_22884,N_22686,N_22572);
or U22885 (N_22885,N_22656,N_22602);
nor U22886 (N_22886,N_22574,N_22747);
and U22887 (N_22887,N_22504,N_22613);
nand U22888 (N_22888,N_22651,N_22640);
nand U22889 (N_22889,N_22666,N_22584);
xnor U22890 (N_22890,N_22659,N_22517);
and U22891 (N_22891,N_22659,N_22693);
xor U22892 (N_22892,N_22616,N_22564);
nand U22893 (N_22893,N_22640,N_22644);
nand U22894 (N_22894,N_22524,N_22532);
or U22895 (N_22895,N_22616,N_22735);
xnor U22896 (N_22896,N_22743,N_22609);
or U22897 (N_22897,N_22731,N_22599);
nor U22898 (N_22898,N_22538,N_22716);
xor U22899 (N_22899,N_22721,N_22639);
xnor U22900 (N_22900,N_22581,N_22689);
nand U22901 (N_22901,N_22622,N_22548);
xor U22902 (N_22902,N_22651,N_22733);
and U22903 (N_22903,N_22629,N_22585);
nor U22904 (N_22904,N_22506,N_22576);
nor U22905 (N_22905,N_22516,N_22717);
nand U22906 (N_22906,N_22687,N_22724);
xor U22907 (N_22907,N_22686,N_22599);
nand U22908 (N_22908,N_22590,N_22709);
and U22909 (N_22909,N_22516,N_22545);
nand U22910 (N_22910,N_22581,N_22644);
or U22911 (N_22911,N_22678,N_22570);
xnor U22912 (N_22912,N_22712,N_22560);
nand U22913 (N_22913,N_22707,N_22726);
nor U22914 (N_22914,N_22571,N_22730);
nor U22915 (N_22915,N_22670,N_22700);
nor U22916 (N_22916,N_22617,N_22517);
nor U22917 (N_22917,N_22560,N_22503);
nand U22918 (N_22918,N_22555,N_22572);
nand U22919 (N_22919,N_22589,N_22605);
nand U22920 (N_22920,N_22662,N_22725);
nor U22921 (N_22921,N_22645,N_22604);
nand U22922 (N_22922,N_22604,N_22692);
nor U22923 (N_22923,N_22725,N_22716);
nand U22924 (N_22924,N_22520,N_22677);
or U22925 (N_22925,N_22553,N_22540);
xor U22926 (N_22926,N_22545,N_22535);
nor U22927 (N_22927,N_22569,N_22517);
nor U22928 (N_22928,N_22719,N_22734);
xnor U22929 (N_22929,N_22687,N_22590);
xnor U22930 (N_22930,N_22620,N_22717);
xor U22931 (N_22931,N_22630,N_22723);
xnor U22932 (N_22932,N_22745,N_22688);
and U22933 (N_22933,N_22514,N_22645);
nor U22934 (N_22934,N_22555,N_22566);
or U22935 (N_22935,N_22729,N_22718);
or U22936 (N_22936,N_22565,N_22710);
nor U22937 (N_22937,N_22546,N_22727);
xor U22938 (N_22938,N_22720,N_22709);
or U22939 (N_22939,N_22557,N_22569);
nand U22940 (N_22940,N_22540,N_22645);
and U22941 (N_22941,N_22611,N_22707);
nor U22942 (N_22942,N_22627,N_22581);
nand U22943 (N_22943,N_22622,N_22717);
xor U22944 (N_22944,N_22585,N_22572);
or U22945 (N_22945,N_22732,N_22614);
xor U22946 (N_22946,N_22711,N_22661);
nor U22947 (N_22947,N_22531,N_22677);
nand U22948 (N_22948,N_22721,N_22615);
nand U22949 (N_22949,N_22700,N_22741);
xor U22950 (N_22950,N_22510,N_22566);
nand U22951 (N_22951,N_22740,N_22695);
nor U22952 (N_22952,N_22511,N_22624);
xor U22953 (N_22953,N_22707,N_22517);
nand U22954 (N_22954,N_22695,N_22616);
xnor U22955 (N_22955,N_22745,N_22741);
or U22956 (N_22956,N_22674,N_22739);
or U22957 (N_22957,N_22672,N_22743);
nand U22958 (N_22958,N_22726,N_22620);
nor U22959 (N_22959,N_22672,N_22544);
or U22960 (N_22960,N_22547,N_22627);
nor U22961 (N_22961,N_22627,N_22738);
or U22962 (N_22962,N_22578,N_22647);
and U22963 (N_22963,N_22635,N_22726);
xor U22964 (N_22964,N_22534,N_22564);
nand U22965 (N_22965,N_22534,N_22633);
and U22966 (N_22966,N_22622,N_22724);
or U22967 (N_22967,N_22576,N_22702);
nand U22968 (N_22968,N_22670,N_22714);
or U22969 (N_22969,N_22702,N_22533);
nor U22970 (N_22970,N_22689,N_22503);
xor U22971 (N_22971,N_22521,N_22721);
xor U22972 (N_22972,N_22669,N_22569);
nand U22973 (N_22973,N_22649,N_22726);
nor U22974 (N_22974,N_22747,N_22707);
nand U22975 (N_22975,N_22584,N_22743);
or U22976 (N_22976,N_22552,N_22602);
xor U22977 (N_22977,N_22719,N_22555);
or U22978 (N_22978,N_22646,N_22721);
xor U22979 (N_22979,N_22626,N_22707);
or U22980 (N_22980,N_22649,N_22624);
and U22981 (N_22981,N_22567,N_22570);
and U22982 (N_22982,N_22704,N_22634);
nand U22983 (N_22983,N_22508,N_22649);
xor U22984 (N_22984,N_22719,N_22735);
or U22985 (N_22985,N_22745,N_22735);
nand U22986 (N_22986,N_22595,N_22549);
xor U22987 (N_22987,N_22523,N_22599);
and U22988 (N_22988,N_22518,N_22665);
and U22989 (N_22989,N_22736,N_22625);
and U22990 (N_22990,N_22607,N_22668);
and U22991 (N_22991,N_22702,N_22627);
nor U22992 (N_22992,N_22537,N_22709);
and U22993 (N_22993,N_22501,N_22517);
nor U22994 (N_22994,N_22724,N_22531);
nor U22995 (N_22995,N_22570,N_22629);
and U22996 (N_22996,N_22594,N_22513);
nand U22997 (N_22997,N_22526,N_22715);
or U22998 (N_22998,N_22509,N_22745);
and U22999 (N_22999,N_22639,N_22509);
and U23000 (N_23000,N_22772,N_22857);
nand U23001 (N_23001,N_22967,N_22753);
xnor U23002 (N_23002,N_22890,N_22852);
nand U23003 (N_23003,N_22929,N_22790);
xnor U23004 (N_23004,N_22818,N_22797);
nor U23005 (N_23005,N_22898,N_22900);
or U23006 (N_23006,N_22986,N_22950);
or U23007 (N_23007,N_22939,N_22905);
nor U23008 (N_23008,N_22845,N_22993);
nand U23009 (N_23009,N_22844,N_22766);
nor U23010 (N_23010,N_22904,N_22817);
nand U23011 (N_23011,N_22769,N_22867);
or U23012 (N_23012,N_22834,N_22851);
nand U23013 (N_23013,N_22914,N_22935);
xor U23014 (N_23014,N_22975,N_22938);
and U23015 (N_23015,N_22759,N_22868);
or U23016 (N_23016,N_22962,N_22850);
nor U23017 (N_23017,N_22765,N_22873);
or U23018 (N_23018,N_22983,N_22903);
nand U23019 (N_23019,N_22936,N_22785);
nand U23020 (N_23020,N_22922,N_22944);
nor U23021 (N_23021,N_22970,N_22913);
nand U23022 (N_23022,N_22948,N_22994);
nand U23023 (N_23023,N_22872,N_22840);
xnor U23024 (N_23024,N_22837,N_22763);
and U23025 (N_23025,N_22902,N_22919);
xnor U23026 (N_23026,N_22953,N_22965);
and U23027 (N_23027,N_22931,N_22980);
xnor U23028 (N_23028,N_22781,N_22760);
nand U23029 (N_23029,N_22943,N_22964);
xnor U23030 (N_23030,N_22816,N_22961);
nor U23031 (N_23031,N_22883,N_22791);
nand U23032 (N_23032,N_22752,N_22786);
nand U23033 (N_23033,N_22966,N_22784);
nand U23034 (N_23034,N_22884,N_22896);
nand U23035 (N_23035,N_22787,N_22798);
and U23036 (N_23036,N_22841,N_22924);
nor U23037 (N_23037,N_22881,N_22799);
nand U23038 (N_23038,N_22888,N_22848);
xnor U23039 (N_23039,N_22991,N_22773);
and U23040 (N_23040,N_22930,N_22978);
xnor U23041 (N_23041,N_22908,N_22774);
and U23042 (N_23042,N_22849,N_22972);
nand U23043 (N_23043,N_22822,N_22916);
nand U23044 (N_23044,N_22937,N_22968);
nand U23045 (N_23045,N_22831,N_22775);
xor U23046 (N_23046,N_22877,N_22928);
and U23047 (N_23047,N_22992,N_22767);
or U23048 (N_23048,N_22814,N_22982);
nor U23049 (N_23049,N_22771,N_22940);
nor U23050 (N_23050,N_22863,N_22979);
and U23051 (N_23051,N_22751,N_22942);
nand U23052 (N_23052,N_22941,N_22889);
nand U23053 (N_23053,N_22754,N_22792);
nor U23054 (N_23054,N_22894,N_22853);
xnor U23055 (N_23055,N_22846,N_22995);
or U23056 (N_23056,N_22807,N_22990);
nor U23057 (N_23057,N_22906,N_22985);
nor U23058 (N_23058,N_22880,N_22907);
xnor U23059 (N_23059,N_22825,N_22912);
nor U23060 (N_23060,N_22915,N_22954);
or U23061 (N_23061,N_22777,N_22882);
and U23062 (N_23062,N_22758,N_22836);
xnor U23063 (N_23063,N_22959,N_22976);
or U23064 (N_23064,N_22886,N_22819);
nor U23065 (N_23065,N_22803,N_22901);
xor U23066 (N_23066,N_22764,N_22805);
or U23067 (N_23067,N_22874,N_22780);
and U23068 (N_23068,N_22789,N_22897);
xnor U23069 (N_23069,N_22804,N_22839);
and U23070 (N_23070,N_22932,N_22909);
nor U23071 (N_23071,N_22933,N_22999);
nor U23072 (N_23072,N_22830,N_22957);
nand U23073 (N_23073,N_22911,N_22815);
nand U23074 (N_23074,N_22963,N_22800);
and U23075 (N_23075,N_22864,N_22843);
xnor U23076 (N_23076,N_22810,N_22768);
or U23077 (N_23077,N_22783,N_22951);
nand U23078 (N_23078,N_22826,N_22885);
or U23079 (N_23079,N_22876,N_22899);
and U23080 (N_23080,N_22947,N_22782);
xor U23081 (N_23081,N_22776,N_22750);
nor U23082 (N_23082,N_22824,N_22757);
xor U23083 (N_23083,N_22862,N_22820);
nor U23084 (N_23084,N_22969,N_22833);
xor U23085 (N_23085,N_22762,N_22971);
or U23086 (N_23086,N_22960,N_22808);
nor U23087 (N_23087,N_22977,N_22921);
xnor U23088 (N_23088,N_22855,N_22756);
nand U23089 (N_23089,N_22871,N_22893);
nand U23090 (N_23090,N_22981,N_22988);
nor U23091 (N_23091,N_22801,N_22956);
xor U23092 (N_23092,N_22794,N_22865);
and U23093 (N_23093,N_22829,N_22895);
nand U23094 (N_23094,N_22770,N_22989);
nor U23095 (N_23095,N_22925,N_22934);
xor U23096 (N_23096,N_22847,N_22984);
xor U23097 (N_23097,N_22779,N_22854);
or U23098 (N_23098,N_22974,N_22793);
xnor U23099 (N_23099,N_22892,N_22809);
nor U23100 (N_23100,N_22955,N_22761);
and U23101 (N_23101,N_22927,N_22869);
and U23102 (N_23102,N_22802,N_22866);
nor U23103 (N_23103,N_22917,N_22910);
or U23104 (N_23104,N_22821,N_22859);
and U23105 (N_23105,N_22823,N_22778);
xnor U23106 (N_23106,N_22952,N_22958);
nor U23107 (N_23107,N_22891,N_22813);
or U23108 (N_23108,N_22861,N_22998);
or U23109 (N_23109,N_22856,N_22926);
and U23110 (N_23110,N_22997,N_22832);
nor U23111 (N_23111,N_22996,N_22949);
and U23112 (N_23112,N_22838,N_22946);
xnor U23113 (N_23113,N_22827,N_22828);
xor U23114 (N_23114,N_22945,N_22920);
or U23115 (N_23115,N_22806,N_22795);
or U23116 (N_23116,N_22858,N_22860);
and U23117 (N_23117,N_22796,N_22755);
nand U23118 (N_23118,N_22878,N_22835);
nand U23119 (N_23119,N_22811,N_22923);
or U23120 (N_23120,N_22973,N_22870);
and U23121 (N_23121,N_22812,N_22842);
nor U23122 (N_23122,N_22918,N_22875);
nand U23123 (N_23123,N_22879,N_22887);
and U23124 (N_23124,N_22987,N_22788);
and U23125 (N_23125,N_22871,N_22922);
nand U23126 (N_23126,N_22816,N_22929);
xnor U23127 (N_23127,N_22762,N_22881);
nor U23128 (N_23128,N_22816,N_22850);
nor U23129 (N_23129,N_22907,N_22765);
nand U23130 (N_23130,N_22758,N_22938);
xor U23131 (N_23131,N_22886,N_22801);
or U23132 (N_23132,N_22909,N_22822);
and U23133 (N_23133,N_22849,N_22956);
and U23134 (N_23134,N_22886,N_22778);
or U23135 (N_23135,N_22840,N_22892);
nor U23136 (N_23136,N_22946,N_22855);
or U23137 (N_23137,N_22820,N_22855);
and U23138 (N_23138,N_22995,N_22889);
and U23139 (N_23139,N_22963,N_22783);
xor U23140 (N_23140,N_22760,N_22814);
nor U23141 (N_23141,N_22773,N_22844);
nor U23142 (N_23142,N_22943,N_22997);
or U23143 (N_23143,N_22787,N_22825);
nor U23144 (N_23144,N_22939,N_22971);
xor U23145 (N_23145,N_22842,N_22896);
nand U23146 (N_23146,N_22893,N_22884);
or U23147 (N_23147,N_22764,N_22856);
nand U23148 (N_23148,N_22942,N_22757);
nand U23149 (N_23149,N_22751,N_22770);
xnor U23150 (N_23150,N_22920,N_22804);
nor U23151 (N_23151,N_22752,N_22869);
nor U23152 (N_23152,N_22820,N_22993);
xnor U23153 (N_23153,N_22774,N_22957);
nor U23154 (N_23154,N_22884,N_22823);
and U23155 (N_23155,N_22942,N_22801);
or U23156 (N_23156,N_22937,N_22877);
nand U23157 (N_23157,N_22831,N_22990);
nor U23158 (N_23158,N_22852,N_22783);
nor U23159 (N_23159,N_22886,N_22848);
nand U23160 (N_23160,N_22830,N_22970);
xor U23161 (N_23161,N_22889,N_22780);
nor U23162 (N_23162,N_22812,N_22860);
nor U23163 (N_23163,N_22873,N_22908);
xnor U23164 (N_23164,N_22813,N_22986);
or U23165 (N_23165,N_22836,N_22880);
xor U23166 (N_23166,N_22828,N_22888);
and U23167 (N_23167,N_22932,N_22891);
nand U23168 (N_23168,N_22961,N_22926);
nand U23169 (N_23169,N_22784,N_22969);
or U23170 (N_23170,N_22913,N_22982);
nor U23171 (N_23171,N_22934,N_22814);
and U23172 (N_23172,N_22828,N_22842);
nor U23173 (N_23173,N_22772,N_22916);
nand U23174 (N_23174,N_22800,N_22915);
nor U23175 (N_23175,N_22962,N_22763);
or U23176 (N_23176,N_22757,N_22887);
or U23177 (N_23177,N_22786,N_22797);
nand U23178 (N_23178,N_22840,N_22806);
xnor U23179 (N_23179,N_22840,N_22895);
nor U23180 (N_23180,N_22961,N_22927);
xor U23181 (N_23181,N_22941,N_22911);
nor U23182 (N_23182,N_22956,N_22998);
xnor U23183 (N_23183,N_22863,N_22934);
xor U23184 (N_23184,N_22761,N_22846);
xnor U23185 (N_23185,N_22784,N_22846);
or U23186 (N_23186,N_22981,N_22931);
and U23187 (N_23187,N_22890,N_22858);
and U23188 (N_23188,N_22800,N_22988);
or U23189 (N_23189,N_22802,N_22792);
nor U23190 (N_23190,N_22756,N_22814);
xnor U23191 (N_23191,N_22938,N_22884);
nand U23192 (N_23192,N_22901,N_22854);
and U23193 (N_23193,N_22930,N_22953);
xor U23194 (N_23194,N_22971,N_22768);
and U23195 (N_23195,N_22819,N_22872);
or U23196 (N_23196,N_22934,N_22856);
or U23197 (N_23197,N_22971,N_22993);
nand U23198 (N_23198,N_22800,N_22778);
nor U23199 (N_23199,N_22753,N_22867);
nor U23200 (N_23200,N_22770,N_22986);
and U23201 (N_23201,N_22784,N_22829);
xnor U23202 (N_23202,N_22789,N_22883);
nand U23203 (N_23203,N_22860,N_22923);
or U23204 (N_23204,N_22879,N_22869);
nand U23205 (N_23205,N_22976,N_22999);
xnor U23206 (N_23206,N_22766,N_22976);
or U23207 (N_23207,N_22857,N_22879);
and U23208 (N_23208,N_22996,N_22971);
nand U23209 (N_23209,N_22952,N_22765);
or U23210 (N_23210,N_22858,N_22817);
or U23211 (N_23211,N_22920,N_22791);
and U23212 (N_23212,N_22764,N_22954);
nor U23213 (N_23213,N_22771,N_22754);
or U23214 (N_23214,N_22936,N_22913);
xor U23215 (N_23215,N_22775,N_22842);
nand U23216 (N_23216,N_22863,N_22819);
xor U23217 (N_23217,N_22979,N_22770);
xnor U23218 (N_23218,N_22820,N_22812);
nor U23219 (N_23219,N_22966,N_22811);
or U23220 (N_23220,N_22849,N_22918);
nor U23221 (N_23221,N_22770,N_22863);
nand U23222 (N_23222,N_22763,N_22877);
or U23223 (N_23223,N_22822,N_22802);
xnor U23224 (N_23224,N_22941,N_22752);
nor U23225 (N_23225,N_22934,N_22817);
xnor U23226 (N_23226,N_22758,N_22765);
and U23227 (N_23227,N_22869,N_22823);
nand U23228 (N_23228,N_22886,N_22882);
and U23229 (N_23229,N_22821,N_22996);
and U23230 (N_23230,N_22781,N_22908);
and U23231 (N_23231,N_22795,N_22918);
nor U23232 (N_23232,N_22984,N_22899);
and U23233 (N_23233,N_22953,N_22927);
xnor U23234 (N_23234,N_22994,N_22878);
and U23235 (N_23235,N_22940,N_22866);
or U23236 (N_23236,N_22962,N_22891);
xnor U23237 (N_23237,N_22865,N_22928);
nor U23238 (N_23238,N_22887,N_22972);
nor U23239 (N_23239,N_22765,N_22754);
and U23240 (N_23240,N_22882,N_22829);
or U23241 (N_23241,N_22771,N_22902);
nor U23242 (N_23242,N_22755,N_22875);
nand U23243 (N_23243,N_22795,N_22997);
nor U23244 (N_23244,N_22753,N_22940);
xnor U23245 (N_23245,N_22839,N_22847);
and U23246 (N_23246,N_22790,N_22889);
nand U23247 (N_23247,N_22824,N_22825);
and U23248 (N_23248,N_22868,N_22862);
and U23249 (N_23249,N_22956,N_22871);
or U23250 (N_23250,N_23010,N_23244);
and U23251 (N_23251,N_23232,N_23173);
xnor U23252 (N_23252,N_23129,N_23153);
nor U23253 (N_23253,N_23145,N_23030);
nand U23254 (N_23254,N_23006,N_23159);
nor U23255 (N_23255,N_23230,N_23065);
xnor U23256 (N_23256,N_23052,N_23091);
nor U23257 (N_23257,N_23190,N_23122);
or U23258 (N_23258,N_23083,N_23020);
nand U23259 (N_23259,N_23124,N_23073);
and U23260 (N_23260,N_23092,N_23204);
xor U23261 (N_23261,N_23031,N_23007);
and U23262 (N_23262,N_23101,N_23016);
xnor U23263 (N_23263,N_23000,N_23189);
or U23264 (N_23264,N_23053,N_23021);
nand U23265 (N_23265,N_23067,N_23044);
nor U23266 (N_23266,N_23150,N_23085);
nand U23267 (N_23267,N_23050,N_23027);
and U23268 (N_23268,N_23017,N_23100);
nor U23269 (N_23269,N_23117,N_23034);
xnor U23270 (N_23270,N_23076,N_23161);
nand U23271 (N_23271,N_23055,N_23127);
xor U23272 (N_23272,N_23023,N_23011);
nand U23273 (N_23273,N_23208,N_23082);
nand U23274 (N_23274,N_23164,N_23035);
nand U23275 (N_23275,N_23206,N_23107);
nor U23276 (N_23276,N_23186,N_23063);
xnor U23277 (N_23277,N_23046,N_23132);
nand U23278 (N_23278,N_23248,N_23199);
and U23279 (N_23279,N_23247,N_23049);
nor U23280 (N_23280,N_23152,N_23013);
and U23281 (N_23281,N_23115,N_23123);
and U23282 (N_23282,N_23181,N_23172);
or U23283 (N_23283,N_23151,N_23227);
nor U23284 (N_23284,N_23045,N_23138);
xor U23285 (N_23285,N_23079,N_23070);
and U23286 (N_23286,N_23165,N_23249);
and U23287 (N_23287,N_23125,N_23059);
and U23288 (N_23288,N_23155,N_23216);
or U23289 (N_23289,N_23141,N_23048);
nor U23290 (N_23290,N_23116,N_23245);
and U23291 (N_23291,N_23109,N_23080);
or U23292 (N_23292,N_23194,N_23197);
nor U23293 (N_23293,N_23179,N_23233);
nor U23294 (N_23294,N_23126,N_23196);
or U23295 (N_23295,N_23191,N_23225);
and U23296 (N_23296,N_23009,N_23108);
nand U23297 (N_23297,N_23043,N_23193);
or U23298 (N_23298,N_23180,N_23195);
and U23299 (N_23299,N_23056,N_23236);
and U23300 (N_23300,N_23111,N_23143);
or U23301 (N_23301,N_23094,N_23240);
xor U23302 (N_23302,N_23157,N_23064);
and U23303 (N_23303,N_23119,N_23062);
or U23304 (N_23304,N_23042,N_23176);
xnor U23305 (N_23305,N_23211,N_23088);
or U23306 (N_23306,N_23201,N_23029);
xnor U23307 (N_23307,N_23170,N_23128);
xnor U23308 (N_23308,N_23096,N_23015);
or U23309 (N_23309,N_23003,N_23239);
and U23310 (N_23310,N_23147,N_23139);
nor U23311 (N_23311,N_23205,N_23198);
nand U23312 (N_23312,N_23051,N_23175);
nand U23313 (N_23313,N_23148,N_23024);
nand U23314 (N_23314,N_23218,N_23058);
xor U23315 (N_23315,N_23037,N_23118);
xnor U23316 (N_23316,N_23113,N_23149);
and U23317 (N_23317,N_23177,N_23078);
nand U23318 (N_23318,N_23033,N_23112);
nand U23319 (N_23319,N_23235,N_23014);
nor U23320 (N_23320,N_23040,N_23209);
or U23321 (N_23321,N_23086,N_23184);
or U23322 (N_23322,N_23140,N_23168);
nand U23323 (N_23323,N_23008,N_23238);
xnor U23324 (N_23324,N_23104,N_23217);
xnor U23325 (N_23325,N_23222,N_23133);
nand U23326 (N_23326,N_23137,N_23039);
nor U23327 (N_23327,N_23054,N_23095);
nand U23328 (N_23328,N_23134,N_23087);
and U23329 (N_23329,N_23019,N_23005);
nor U23330 (N_23330,N_23167,N_23229);
nand U23331 (N_23331,N_23213,N_23012);
or U23332 (N_23332,N_23038,N_23068);
nor U23333 (N_23333,N_23242,N_23142);
nor U23334 (N_23334,N_23243,N_23188);
nor U23335 (N_23335,N_23098,N_23163);
nand U23336 (N_23336,N_23219,N_23146);
and U23337 (N_23337,N_23081,N_23075);
and U23338 (N_23338,N_23071,N_23202);
xnor U23339 (N_23339,N_23099,N_23032);
nand U23340 (N_23340,N_23131,N_23121);
nand U23341 (N_23341,N_23212,N_23136);
xor U23342 (N_23342,N_23077,N_23097);
nor U23343 (N_23343,N_23187,N_23215);
or U23344 (N_23344,N_23018,N_23234);
and U23345 (N_23345,N_23025,N_23154);
and U23346 (N_23346,N_23174,N_23102);
and U23347 (N_23347,N_23069,N_23090);
and U23348 (N_23348,N_23185,N_23061);
and U23349 (N_23349,N_23057,N_23114);
and U23350 (N_23350,N_23047,N_23120);
nor U23351 (N_23351,N_23200,N_23210);
nand U23352 (N_23352,N_23220,N_23093);
or U23353 (N_23353,N_23169,N_23171);
and U23354 (N_23354,N_23158,N_23226);
nand U23355 (N_23355,N_23036,N_23026);
or U23356 (N_23356,N_23178,N_23130);
xnor U23357 (N_23357,N_23074,N_23066);
nor U23358 (N_23358,N_23041,N_23084);
nor U23359 (N_23359,N_23089,N_23228);
nor U23360 (N_23360,N_23192,N_23221);
and U23361 (N_23361,N_23002,N_23223);
or U23362 (N_23362,N_23182,N_23231);
and U23363 (N_23363,N_23022,N_23203);
or U23364 (N_23364,N_23241,N_23183);
nand U23365 (N_23365,N_23166,N_23060);
xor U23366 (N_23366,N_23001,N_23144);
nor U23367 (N_23367,N_23207,N_23105);
and U23368 (N_23368,N_23162,N_23224);
and U23369 (N_23369,N_23028,N_23237);
nor U23370 (N_23370,N_23135,N_23072);
nor U23371 (N_23371,N_23004,N_23214);
and U23372 (N_23372,N_23110,N_23103);
nand U23373 (N_23373,N_23106,N_23246);
nand U23374 (N_23374,N_23156,N_23160);
or U23375 (N_23375,N_23181,N_23013);
nand U23376 (N_23376,N_23035,N_23143);
and U23377 (N_23377,N_23214,N_23185);
and U23378 (N_23378,N_23181,N_23146);
nor U23379 (N_23379,N_23031,N_23192);
xor U23380 (N_23380,N_23147,N_23184);
nor U23381 (N_23381,N_23054,N_23000);
nand U23382 (N_23382,N_23193,N_23023);
nor U23383 (N_23383,N_23107,N_23217);
xnor U23384 (N_23384,N_23089,N_23138);
and U23385 (N_23385,N_23028,N_23232);
xnor U23386 (N_23386,N_23047,N_23152);
and U23387 (N_23387,N_23101,N_23067);
and U23388 (N_23388,N_23197,N_23071);
and U23389 (N_23389,N_23221,N_23059);
nand U23390 (N_23390,N_23008,N_23103);
nand U23391 (N_23391,N_23025,N_23108);
or U23392 (N_23392,N_23000,N_23178);
and U23393 (N_23393,N_23120,N_23192);
xnor U23394 (N_23394,N_23158,N_23141);
nand U23395 (N_23395,N_23139,N_23179);
xnor U23396 (N_23396,N_23114,N_23140);
or U23397 (N_23397,N_23167,N_23204);
and U23398 (N_23398,N_23238,N_23126);
or U23399 (N_23399,N_23203,N_23146);
and U23400 (N_23400,N_23204,N_23189);
xor U23401 (N_23401,N_23065,N_23042);
xor U23402 (N_23402,N_23104,N_23060);
nand U23403 (N_23403,N_23126,N_23204);
and U23404 (N_23404,N_23030,N_23083);
and U23405 (N_23405,N_23105,N_23059);
xnor U23406 (N_23406,N_23022,N_23239);
nand U23407 (N_23407,N_23063,N_23119);
nor U23408 (N_23408,N_23181,N_23122);
or U23409 (N_23409,N_23037,N_23175);
and U23410 (N_23410,N_23200,N_23069);
xor U23411 (N_23411,N_23212,N_23243);
xnor U23412 (N_23412,N_23062,N_23047);
or U23413 (N_23413,N_23128,N_23076);
or U23414 (N_23414,N_23108,N_23150);
and U23415 (N_23415,N_23167,N_23184);
nand U23416 (N_23416,N_23195,N_23152);
and U23417 (N_23417,N_23238,N_23110);
and U23418 (N_23418,N_23145,N_23033);
and U23419 (N_23419,N_23067,N_23104);
and U23420 (N_23420,N_23137,N_23028);
nor U23421 (N_23421,N_23243,N_23230);
or U23422 (N_23422,N_23073,N_23007);
xnor U23423 (N_23423,N_23133,N_23239);
nand U23424 (N_23424,N_23043,N_23179);
xor U23425 (N_23425,N_23095,N_23112);
or U23426 (N_23426,N_23144,N_23215);
or U23427 (N_23427,N_23095,N_23058);
xnor U23428 (N_23428,N_23235,N_23207);
nor U23429 (N_23429,N_23042,N_23158);
and U23430 (N_23430,N_23001,N_23038);
or U23431 (N_23431,N_23146,N_23051);
nand U23432 (N_23432,N_23041,N_23175);
and U23433 (N_23433,N_23092,N_23129);
and U23434 (N_23434,N_23165,N_23123);
nor U23435 (N_23435,N_23219,N_23054);
nor U23436 (N_23436,N_23142,N_23136);
nand U23437 (N_23437,N_23139,N_23005);
and U23438 (N_23438,N_23012,N_23088);
nor U23439 (N_23439,N_23034,N_23188);
or U23440 (N_23440,N_23182,N_23084);
nand U23441 (N_23441,N_23205,N_23025);
xor U23442 (N_23442,N_23197,N_23147);
xnor U23443 (N_23443,N_23071,N_23106);
nor U23444 (N_23444,N_23126,N_23149);
or U23445 (N_23445,N_23181,N_23174);
or U23446 (N_23446,N_23087,N_23222);
and U23447 (N_23447,N_23239,N_23113);
and U23448 (N_23448,N_23075,N_23203);
or U23449 (N_23449,N_23177,N_23226);
xnor U23450 (N_23450,N_23236,N_23043);
and U23451 (N_23451,N_23134,N_23143);
nand U23452 (N_23452,N_23158,N_23208);
xnor U23453 (N_23453,N_23206,N_23104);
and U23454 (N_23454,N_23219,N_23237);
nand U23455 (N_23455,N_23006,N_23148);
and U23456 (N_23456,N_23194,N_23028);
nor U23457 (N_23457,N_23217,N_23180);
nor U23458 (N_23458,N_23102,N_23085);
nor U23459 (N_23459,N_23166,N_23001);
or U23460 (N_23460,N_23175,N_23085);
and U23461 (N_23461,N_23249,N_23116);
nor U23462 (N_23462,N_23249,N_23172);
nand U23463 (N_23463,N_23151,N_23176);
nor U23464 (N_23464,N_23134,N_23034);
xor U23465 (N_23465,N_23205,N_23019);
nand U23466 (N_23466,N_23015,N_23105);
xor U23467 (N_23467,N_23200,N_23055);
or U23468 (N_23468,N_23089,N_23034);
nand U23469 (N_23469,N_23111,N_23176);
and U23470 (N_23470,N_23001,N_23215);
and U23471 (N_23471,N_23109,N_23009);
and U23472 (N_23472,N_23243,N_23220);
nand U23473 (N_23473,N_23044,N_23021);
or U23474 (N_23474,N_23052,N_23097);
and U23475 (N_23475,N_23229,N_23237);
or U23476 (N_23476,N_23073,N_23110);
xnor U23477 (N_23477,N_23213,N_23124);
or U23478 (N_23478,N_23078,N_23215);
or U23479 (N_23479,N_23050,N_23161);
nand U23480 (N_23480,N_23096,N_23091);
nor U23481 (N_23481,N_23180,N_23193);
xor U23482 (N_23482,N_23073,N_23027);
or U23483 (N_23483,N_23063,N_23031);
nand U23484 (N_23484,N_23001,N_23180);
and U23485 (N_23485,N_23107,N_23157);
and U23486 (N_23486,N_23024,N_23017);
nor U23487 (N_23487,N_23016,N_23204);
nand U23488 (N_23488,N_23068,N_23183);
nand U23489 (N_23489,N_23159,N_23019);
nor U23490 (N_23490,N_23207,N_23145);
and U23491 (N_23491,N_23202,N_23181);
nand U23492 (N_23492,N_23119,N_23243);
and U23493 (N_23493,N_23168,N_23232);
xnor U23494 (N_23494,N_23151,N_23146);
nor U23495 (N_23495,N_23046,N_23084);
or U23496 (N_23496,N_23081,N_23071);
and U23497 (N_23497,N_23131,N_23164);
or U23498 (N_23498,N_23198,N_23035);
xnor U23499 (N_23499,N_23229,N_23067);
and U23500 (N_23500,N_23358,N_23283);
xor U23501 (N_23501,N_23479,N_23343);
nor U23502 (N_23502,N_23381,N_23452);
xnor U23503 (N_23503,N_23350,N_23386);
or U23504 (N_23504,N_23314,N_23433);
or U23505 (N_23505,N_23254,N_23422);
nand U23506 (N_23506,N_23404,N_23408);
or U23507 (N_23507,N_23388,N_23366);
xor U23508 (N_23508,N_23423,N_23313);
xor U23509 (N_23509,N_23345,N_23458);
nand U23510 (N_23510,N_23259,N_23490);
or U23511 (N_23511,N_23496,N_23330);
nand U23512 (N_23512,N_23383,N_23339);
and U23513 (N_23513,N_23453,N_23435);
or U23514 (N_23514,N_23438,N_23318);
xor U23515 (N_23515,N_23307,N_23364);
nand U23516 (N_23516,N_23252,N_23402);
and U23517 (N_23517,N_23323,N_23424);
or U23518 (N_23518,N_23338,N_23352);
nand U23519 (N_23519,N_23387,N_23341);
nor U23520 (N_23520,N_23380,N_23297);
or U23521 (N_23521,N_23480,N_23414);
and U23522 (N_23522,N_23348,N_23489);
nor U23523 (N_23523,N_23329,N_23403);
nor U23524 (N_23524,N_23442,N_23264);
or U23525 (N_23525,N_23346,N_23320);
and U23526 (N_23526,N_23400,N_23434);
and U23527 (N_23527,N_23494,N_23472);
nand U23528 (N_23528,N_23287,N_23253);
or U23529 (N_23529,N_23260,N_23405);
nand U23530 (N_23530,N_23284,N_23272);
nor U23531 (N_23531,N_23411,N_23292);
or U23532 (N_23532,N_23270,N_23427);
xor U23533 (N_23533,N_23310,N_23406);
xor U23534 (N_23534,N_23371,N_23436);
xor U23535 (N_23535,N_23362,N_23293);
or U23536 (N_23536,N_23360,N_23456);
or U23537 (N_23537,N_23258,N_23356);
nor U23538 (N_23538,N_23332,N_23417);
or U23539 (N_23539,N_23275,N_23291);
nor U23540 (N_23540,N_23466,N_23491);
or U23541 (N_23541,N_23482,N_23476);
xnor U23542 (N_23542,N_23295,N_23263);
and U23543 (N_23543,N_23398,N_23429);
and U23544 (N_23544,N_23495,N_23333);
xor U23545 (N_23545,N_23484,N_23374);
nand U23546 (N_23546,N_23385,N_23394);
xnor U23547 (N_23547,N_23474,N_23445);
xnor U23548 (N_23548,N_23357,N_23301);
nand U23549 (N_23549,N_23493,N_23447);
or U23550 (N_23550,N_23267,N_23441);
or U23551 (N_23551,N_23271,N_23351);
nand U23552 (N_23552,N_23321,N_23342);
and U23553 (N_23553,N_23379,N_23296);
xnor U23554 (N_23554,N_23355,N_23288);
xnor U23555 (N_23555,N_23334,N_23281);
and U23556 (N_23556,N_23390,N_23431);
nor U23557 (N_23557,N_23274,N_23426);
or U23558 (N_23558,N_23328,N_23409);
nand U23559 (N_23559,N_23319,N_23309);
and U23560 (N_23560,N_23378,N_23460);
xor U23561 (N_23561,N_23285,N_23444);
or U23562 (N_23562,N_23266,N_23468);
nand U23563 (N_23563,N_23459,N_23365);
nor U23564 (N_23564,N_23473,N_23485);
xnor U23565 (N_23565,N_23377,N_23265);
or U23566 (N_23566,N_23420,N_23477);
or U23567 (N_23567,N_23298,N_23389);
nand U23568 (N_23568,N_23488,N_23337);
nor U23569 (N_23569,N_23478,N_23467);
or U23570 (N_23570,N_23425,N_23443);
xnor U23571 (N_23571,N_23449,N_23277);
nor U23572 (N_23572,N_23311,N_23457);
nor U23573 (N_23573,N_23269,N_23363);
nand U23574 (N_23574,N_23344,N_23373);
and U23575 (N_23575,N_23497,N_23289);
nand U23576 (N_23576,N_23483,N_23300);
and U23577 (N_23577,N_23372,N_23354);
and U23578 (N_23578,N_23439,N_23499);
or U23579 (N_23579,N_23440,N_23450);
and U23580 (N_23580,N_23303,N_23257);
and U23581 (N_23581,N_23463,N_23279);
nor U23582 (N_23582,N_23273,N_23261);
nand U23583 (N_23583,N_23325,N_23401);
xor U23584 (N_23584,N_23384,N_23294);
nor U23585 (N_23585,N_23268,N_23396);
nor U23586 (N_23586,N_23286,N_23306);
nand U23587 (N_23587,N_23397,N_23481);
nand U23588 (N_23588,N_23349,N_23308);
nor U23589 (N_23589,N_23317,N_23461);
xor U23590 (N_23590,N_23305,N_23369);
nor U23591 (N_23591,N_23471,N_23340);
and U23592 (N_23592,N_23312,N_23486);
xnor U23593 (N_23593,N_23280,N_23421);
nor U23594 (N_23594,N_23399,N_23392);
xnor U23595 (N_23595,N_23262,N_23324);
nor U23596 (N_23596,N_23415,N_23469);
nand U23597 (N_23597,N_23492,N_23335);
nor U23598 (N_23598,N_23454,N_23498);
xor U23599 (N_23599,N_23278,N_23451);
or U23600 (N_23600,N_23455,N_23282);
xnor U23601 (N_23601,N_23418,N_23250);
nand U23602 (N_23602,N_23375,N_23465);
nand U23603 (N_23603,N_23487,N_23470);
xor U23604 (N_23604,N_23251,N_23410);
and U23605 (N_23605,N_23327,N_23464);
and U23606 (N_23606,N_23322,N_23462);
xnor U23607 (N_23607,N_23382,N_23367);
xnor U23608 (N_23608,N_23448,N_23419);
xor U23609 (N_23609,N_23368,N_23437);
nand U23610 (N_23610,N_23412,N_23428);
nor U23611 (N_23611,N_23413,N_23255);
xnor U23612 (N_23612,N_23370,N_23316);
nor U23613 (N_23613,N_23331,N_23347);
and U23614 (N_23614,N_23299,N_23407);
or U23615 (N_23615,N_23376,N_23315);
xnor U23616 (N_23616,N_23290,N_23276);
xor U23617 (N_23617,N_23336,N_23446);
nor U23618 (N_23618,N_23416,N_23430);
or U23619 (N_23619,N_23361,N_23304);
nor U23620 (N_23620,N_23395,N_23302);
and U23621 (N_23621,N_23359,N_23326);
or U23622 (N_23622,N_23353,N_23475);
nor U23623 (N_23623,N_23432,N_23256);
nor U23624 (N_23624,N_23391,N_23393);
or U23625 (N_23625,N_23468,N_23301);
nand U23626 (N_23626,N_23336,N_23442);
or U23627 (N_23627,N_23348,N_23331);
nand U23628 (N_23628,N_23278,N_23478);
nand U23629 (N_23629,N_23404,N_23323);
or U23630 (N_23630,N_23283,N_23378);
and U23631 (N_23631,N_23327,N_23370);
nand U23632 (N_23632,N_23260,N_23457);
or U23633 (N_23633,N_23273,N_23435);
xnor U23634 (N_23634,N_23467,N_23338);
xor U23635 (N_23635,N_23293,N_23447);
nand U23636 (N_23636,N_23364,N_23292);
xor U23637 (N_23637,N_23444,N_23365);
xnor U23638 (N_23638,N_23256,N_23409);
nand U23639 (N_23639,N_23488,N_23254);
xor U23640 (N_23640,N_23251,N_23384);
xor U23641 (N_23641,N_23348,N_23342);
nor U23642 (N_23642,N_23438,N_23417);
nor U23643 (N_23643,N_23310,N_23283);
nand U23644 (N_23644,N_23393,N_23296);
xnor U23645 (N_23645,N_23474,N_23471);
xor U23646 (N_23646,N_23475,N_23489);
nor U23647 (N_23647,N_23337,N_23301);
nor U23648 (N_23648,N_23416,N_23485);
nor U23649 (N_23649,N_23431,N_23479);
or U23650 (N_23650,N_23443,N_23499);
nor U23651 (N_23651,N_23387,N_23452);
nand U23652 (N_23652,N_23334,N_23484);
and U23653 (N_23653,N_23371,N_23275);
or U23654 (N_23654,N_23294,N_23275);
nand U23655 (N_23655,N_23459,N_23445);
nand U23656 (N_23656,N_23341,N_23421);
nor U23657 (N_23657,N_23442,N_23363);
or U23658 (N_23658,N_23456,N_23413);
or U23659 (N_23659,N_23348,N_23285);
xnor U23660 (N_23660,N_23374,N_23467);
xnor U23661 (N_23661,N_23417,N_23327);
and U23662 (N_23662,N_23465,N_23371);
xnor U23663 (N_23663,N_23276,N_23412);
nor U23664 (N_23664,N_23442,N_23439);
nor U23665 (N_23665,N_23441,N_23474);
nor U23666 (N_23666,N_23383,N_23438);
and U23667 (N_23667,N_23444,N_23463);
nor U23668 (N_23668,N_23354,N_23498);
and U23669 (N_23669,N_23332,N_23290);
or U23670 (N_23670,N_23315,N_23445);
or U23671 (N_23671,N_23412,N_23274);
or U23672 (N_23672,N_23364,N_23282);
nand U23673 (N_23673,N_23418,N_23273);
nand U23674 (N_23674,N_23257,N_23345);
nor U23675 (N_23675,N_23403,N_23327);
and U23676 (N_23676,N_23456,N_23400);
and U23677 (N_23677,N_23440,N_23466);
nor U23678 (N_23678,N_23270,N_23328);
or U23679 (N_23679,N_23376,N_23387);
or U23680 (N_23680,N_23425,N_23259);
nor U23681 (N_23681,N_23469,N_23291);
or U23682 (N_23682,N_23394,N_23266);
nand U23683 (N_23683,N_23470,N_23476);
xnor U23684 (N_23684,N_23375,N_23478);
nand U23685 (N_23685,N_23340,N_23427);
and U23686 (N_23686,N_23377,N_23376);
nor U23687 (N_23687,N_23447,N_23281);
nor U23688 (N_23688,N_23278,N_23316);
nand U23689 (N_23689,N_23412,N_23283);
nand U23690 (N_23690,N_23295,N_23494);
nor U23691 (N_23691,N_23467,N_23335);
or U23692 (N_23692,N_23462,N_23438);
and U23693 (N_23693,N_23325,N_23307);
and U23694 (N_23694,N_23349,N_23454);
nor U23695 (N_23695,N_23457,N_23324);
or U23696 (N_23696,N_23295,N_23275);
or U23697 (N_23697,N_23412,N_23347);
nor U23698 (N_23698,N_23386,N_23276);
or U23699 (N_23699,N_23283,N_23417);
and U23700 (N_23700,N_23408,N_23479);
xnor U23701 (N_23701,N_23402,N_23329);
and U23702 (N_23702,N_23430,N_23277);
and U23703 (N_23703,N_23340,N_23435);
xnor U23704 (N_23704,N_23492,N_23424);
or U23705 (N_23705,N_23336,N_23448);
nor U23706 (N_23706,N_23429,N_23484);
or U23707 (N_23707,N_23392,N_23413);
nor U23708 (N_23708,N_23334,N_23476);
and U23709 (N_23709,N_23287,N_23399);
nor U23710 (N_23710,N_23364,N_23263);
nand U23711 (N_23711,N_23491,N_23323);
nand U23712 (N_23712,N_23402,N_23470);
nand U23713 (N_23713,N_23334,N_23348);
nor U23714 (N_23714,N_23498,N_23378);
or U23715 (N_23715,N_23289,N_23302);
xnor U23716 (N_23716,N_23495,N_23270);
nand U23717 (N_23717,N_23268,N_23455);
xnor U23718 (N_23718,N_23377,N_23430);
xor U23719 (N_23719,N_23435,N_23357);
nand U23720 (N_23720,N_23392,N_23254);
or U23721 (N_23721,N_23474,N_23253);
nand U23722 (N_23722,N_23263,N_23303);
or U23723 (N_23723,N_23376,N_23378);
or U23724 (N_23724,N_23305,N_23379);
xor U23725 (N_23725,N_23284,N_23400);
and U23726 (N_23726,N_23487,N_23421);
nor U23727 (N_23727,N_23330,N_23285);
xnor U23728 (N_23728,N_23343,N_23275);
nand U23729 (N_23729,N_23494,N_23359);
nand U23730 (N_23730,N_23494,N_23366);
nor U23731 (N_23731,N_23447,N_23291);
nand U23732 (N_23732,N_23257,N_23454);
and U23733 (N_23733,N_23250,N_23363);
and U23734 (N_23734,N_23440,N_23448);
and U23735 (N_23735,N_23295,N_23344);
nor U23736 (N_23736,N_23366,N_23459);
xnor U23737 (N_23737,N_23314,N_23343);
or U23738 (N_23738,N_23337,N_23485);
nand U23739 (N_23739,N_23435,N_23382);
nand U23740 (N_23740,N_23258,N_23372);
and U23741 (N_23741,N_23299,N_23386);
nand U23742 (N_23742,N_23441,N_23329);
nand U23743 (N_23743,N_23498,N_23251);
and U23744 (N_23744,N_23277,N_23396);
nor U23745 (N_23745,N_23361,N_23268);
xnor U23746 (N_23746,N_23321,N_23388);
nor U23747 (N_23747,N_23461,N_23337);
nand U23748 (N_23748,N_23277,N_23303);
xnor U23749 (N_23749,N_23489,N_23377);
xor U23750 (N_23750,N_23507,N_23679);
nand U23751 (N_23751,N_23608,N_23590);
or U23752 (N_23752,N_23605,N_23640);
nand U23753 (N_23753,N_23637,N_23621);
xor U23754 (N_23754,N_23558,N_23514);
nor U23755 (N_23755,N_23681,N_23606);
nor U23756 (N_23756,N_23645,N_23740);
and U23757 (N_23757,N_23564,N_23698);
or U23758 (N_23758,N_23529,N_23643);
nor U23759 (N_23759,N_23734,N_23589);
xnor U23760 (N_23760,N_23594,N_23631);
or U23761 (N_23761,N_23647,N_23702);
nor U23762 (N_23762,N_23569,N_23708);
or U23763 (N_23763,N_23713,N_23718);
nand U23764 (N_23764,N_23554,N_23584);
or U23765 (N_23765,N_23692,N_23635);
nand U23766 (N_23766,N_23559,N_23628);
nand U23767 (N_23767,N_23693,N_23676);
or U23768 (N_23768,N_23524,N_23501);
nor U23769 (N_23769,N_23662,N_23537);
nor U23770 (N_23770,N_23700,N_23639);
xor U23771 (N_23771,N_23502,N_23688);
nor U23772 (N_23772,N_23603,N_23579);
xor U23773 (N_23773,N_23586,N_23585);
xor U23774 (N_23774,N_23611,N_23598);
and U23775 (N_23775,N_23632,N_23546);
nor U23776 (N_23776,N_23595,N_23733);
or U23777 (N_23777,N_23601,N_23675);
nor U23778 (N_23778,N_23684,N_23654);
or U23779 (N_23779,N_23682,N_23660);
and U23780 (N_23780,N_23642,N_23604);
and U23781 (N_23781,N_23510,N_23687);
and U23782 (N_23782,N_23691,N_23652);
xor U23783 (N_23783,N_23587,N_23553);
nand U23784 (N_23784,N_23661,N_23739);
or U23785 (N_23785,N_23532,N_23509);
nand U23786 (N_23786,N_23591,N_23508);
nand U23787 (N_23787,N_23746,N_23527);
xnor U23788 (N_23788,N_23549,N_23505);
or U23789 (N_23789,N_23671,N_23523);
nand U23790 (N_23790,N_23748,N_23503);
nand U23791 (N_23791,N_23607,N_23724);
or U23792 (N_23792,N_23511,N_23578);
or U23793 (N_23793,N_23583,N_23539);
or U23794 (N_23794,N_23519,N_23528);
or U23795 (N_23795,N_23720,N_23582);
or U23796 (N_23796,N_23737,N_23612);
or U23797 (N_23797,N_23735,N_23525);
or U23798 (N_23798,N_23518,N_23536);
xor U23799 (N_23799,N_23513,N_23592);
nand U23800 (N_23800,N_23540,N_23723);
nand U23801 (N_23801,N_23575,N_23573);
xor U23802 (N_23802,N_23663,N_23580);
or U23803 (N_23803,N_23581,N_23609);
nor U23804 (N_23804,N_23618,N_23747);
nor U23805 (N_23805,N_23659,N_23665);
nor U23806 (N_23806,N_23664,N_23516);
xnor U23807 (N_23807,N_23650,N_23577);
and U23808 (N_23808,N_23726,N_23567);
or U23809 (N_23809,N_23701,N_23695);
and U23810 (N_23810,N_23504,N_23556);
nor U23811 (N_23811,N_23534,N_23562);
nor U23812 (N_23812,N_23619,N_23657);
xor U23813 (N_23813,N_23576,N_23615);
or U23814 (N_23814,N_23714,N_23593);
nand U23815 (N_23815,N_23625,N_23543);
and U23816 (N_23816,N_23669,N_23568);
xor U23817 (N_23817,N_23703,N_23709);
nor U23818 (N_23818,N_23636,N_23743);
nand U23819 (N_23819,N_23694,N_23614);
nor U23820 (N_23820,N_23570,N_23638);
nor U23821 (N_23821,N_23715,N_23633);
or U23822 (N_23822,N_23599,N_23732);
nor U23823 (N_23823,N_23544,N_23566);
and U23824 (N_23824,N_23533,N_23626);
and U23825 (N_23825,N_23613,N_23744);
xnor U23826 (N_23826,N_23706,N_23572);
and U23827 (N_23827,N_23600,N_23722);
nor U23828 (N_23828,N_23646,N_23641);
nor U23829 (N_23829,N_23565,N_23571);
nor U23830 (N_23830,N_23506,N_23712);
and U23831 (N_23831,N_23547,N_23710);
nor U23832 (N_23832,N_23531,N_23538);
nor U23833 (N_23833,N_23542,N_23648);
xnor U23834 (N_23834,N_23629,N_23597);
nor U23835 (N_23835,N_23749,N_23500);
and U23836 (N_23836,N_23670,N_23727);
nor U23837 (N_23837,N_23574,N_23742);
or U23838 (N_23838,N_23725,N_23563);
nor U23839 (N_23839,N_23736,N_23738);
nand U23840 (N_23840,N_23627,N_23535);
or U23841 (N_23841,N_23686,N_23551);
and U23842 (N_23842,N_23696,N_23655);
or U23843 (N_23843,N_23561,N_23690);
xor U23844 (N_23844,N_23677,N_23674);
nand U23845 (N_23845,N_23719,N_23624);
and U23846 (N_23846,N_23711,N_23699);
or U23847 (N_23847,N_23522,N_23666);
nor U23848 (N_23848,N_23667,N_23517);
xnor U23849 (N_23849,N_23588,N_23515);
and U23850 (N_23850,N_23704,N_23680);
and U23851 (N_23851,N_23512,N_23545);
nand U23852 (N_23852,N_23602,N_23745);
and U23853 (N_23853,N_23634,N_23555);
nand U23854 (N_23854,N_23685,N_23521);
xor U23855 (N_23855,N_23649,N_23707);
or U23856 (N_23856,N_23731,N_23717);
nor U23857 (N_23857,N_23530,N_23689);
nand U23858 (N_23858,N_23610,N_23653);
nor U23859 (N_23859,N_23651,N_23596);
or U23860 (N_23860,N_23644,N_23673);
nand U23861 (N_23861,N_23520,N_23658);
or U23862 (N_23862,N_23620,N_23541);
nand U23863 (N_23863,N_23622,N_23630);
nand U23864 (N_23864,N_23557,N_23552);
nand U23865 (N_23865,N_23697,N_23668);
or U23866 (N_23866,N_23729,N_23728);
xor U23867 (N_23867,N_23616,N_23716);
nor U23868 (N_23868,N_23721,N_23548);
and U23869 (N_23869,N_23526,N_23678);
nor U23870 (N_23870,N_23550,N_23705);
or U23871 (N_23871,N_23730,N_23560);
nand U23872 (N_23872,N_23683,N_23617);
or U23873 (N_23873,N_23741,N_23656);
nand U23874 (N_23874,N_23623,N_23672);
nand U23875 (N_23875,N_23563,N_23542);
xor U23876 (N_23876,N_23611,N_23536);
xnor U23877 (N_23877,N_23598,N_23575);
xor U23878 (N_23878,N_23633,N_23553);
nor U23879 (N_23879,N_23744,N_23694);
xor U23880 (N_23880,N_23686,N_23748);
nor U23881 (N_23881,N_23733,N_23582);
nor U23882 (N_23882,N_23579,N_23634);
and U23883 (N_23883,N_23552,N_23748);
and U23884 (N_23884,N_23597,N_23683);
nand U23885 (N_23885,N_23631,N_23709);
xnor U23886 (N_23886,N_23742,N_23617);
nor U23887 (N_23887,N_23656,N_23565);
nand U23888 (N_23888,N_23717,N_23687);
nor U23889 (N_23889,N_23528,N_23572);
nand U23890 (N_23890,N_23583,N_23525);
nand U23891 (N_23891,N_23660,N_23703);
or U23892 (N_23892,N_23727,N_23592);
xnor U23893 (N_23893,N_23595,N_23743);
and U23894 (N_23894,N_23503,N_23537);
xor U23895 (N_23895,N_23679,N_23628);
or U23896 (N_23896,N_23548,N_23709);
nor U23897 (N_23897,N_23698,N_23546);
or U23898 (N_23898,N_23502,N_23728);
xor U23899 (N_23899,N_23692,N_23671);
nor U23900 (N_23900,N_23745,N_23646);
nand U23901 (N_23901,N_23582,N_23682);
xnor U23902 (N_23902,N_23696,N_23539);
nand U23903 (N_23903,N_23625,N_23584);
or U23904 (N_23904,N_23524,N_23547);
and U23905 (N_23905,N_23667,N_23576);
xor U23906 (N_23906,N_23631,N_23511);
nor U23907 (N_23907,N_23552,N_23671);
and U23908 (N_23908,N_23515,N_23586);
or U23909 (N_23909,N_23731,N_23707);
and U23910 (N_23910,N_23676,N_23734);
or U23911 (N_23911,N_23712,N_23743);
nor U23912 (N_23912,N_23604,N_23645);
and U23913 (N_23913,N_23747,N_23571);
nand U23914 (N_23914,N_23629,N_23639);
and U23915 (N_23915,N_23706,N_23560);
nor U23916 (N_23916,N_23572,N_23657);
nand U23917 (N_23917,N_23578,N_23625);
or U23918 (N_23918,N_23547,N_23546);
xor U23919 (N_23919,N_23517,N_23607);
and U23920 (N_23920,N_23536,N_23519);
nand U23921 (N_23921,N_23696,N_23693);
and U23922 (N_23922,N_23684,N_23578);
nand U23923 (N_23923,N_23626,N_23552);
xnor U23924 (N_23924,N_23652,N_23540);
xor U23925 (N_23925,N_23512,N_23747);
nor U23926 (N_23926,N_23592,N_23735);
xor U23927 (N_23927,N_23745,N_23678);
or U23928 (N_23928,N_23678,N_23638);
nand U23929 (N_23929,N_23520,N_23608);
xnor U23930 (N_23930,N_23705,N_23749);
nor U23931 (N_23931,N_23517,N_23707);
and U23932 (N_23932,N_23743,N_23500);
xor U23933 (N_23933,N_23590,N_23558);
or U23934 (N_23934,N_23506,N_23519);
nor U23935 (N_23935,N_23557,N_23601);
xor U23936 (N_23936,N_23601,N_23654);
and U23937 (N_23937,N_23621,N_23665);
and U23938 (N_23938,N_23621,N_23652);
or U23939 (N_23939,N_23647,N_23540);
xnor U23940 (N_23940,N_23507,N_23516);
nand U23941 (N_23941,N_23620,N_23717);
and U23942 (N_23942,N_23624,N_23503);
xor U23943 (N_23943,N_23742,N_23584);
and U23944 (N_23944,N_23622,N_23688);
and U23945 (N_23945,N_23730,N_23505);
nor U23946 (N_23946,N_23621,N_23526);
and U23947 (N_23947,N_23536,N_23689);
nor U23948 (N_23948,N_23507,N_23648);
nand U23949 (N_23949,N_23619,N_23744);
nand U23950 (N_23950,N_23695,N_23721);
and U23951 (N_23951,N_23703,N_23735);
nand U23952 (N_23952,N_23513,N_23502);
xnor U23953 (N_23953,N_23669,N_23733);
nor U23954 (N_23954,N_23738,N_23516);
xor U23955 (N_23955,N_23621,N_23506);
and U23956 (N_23956,N_23659,N_23680);
or U23957 (N_23957,N_23539,N_23632);
nor U23958 (N_23958,N_23746,N_23614);
nor U23959 (N_23959,N_23563,N_23651);
nand U23960 (N_23960,N_23540,N_23581);
nand U23961 (N_23961,N_23714,N_23656);
and U23962 (N_23962,N_23636,N_23631);
nor U23963 (N_23963,N_23715,N_23703);
nand U23964 (N_23964,N_23558,N_23552);
and U23965 (N_23965,N_23559,N_23526);
or U23966 (N_23966,N_23703,N_23540);
or U23967 (N_23967,N_23705,N_23650);
xor U23968 (N_23968,N_23678,N_23620);
or U23969 (N_23969,N_23581,N_23656);
and U23970 (N_23970,N_23525,N_23720);
xnor U23971 (N_23971,N_23628,N_23568);
nand U23972 (N_23972,N_23624,N_23590);
nor U23973 (N_23973,N_23590,N_23695);
nand U23974 (N_23974,N_23529,N_23541);
nor U23975 (N_23975,N_23690,N_23639);
nor U23976 (N_23976,N_23621,N_23684);
nand U23977 (N_23977,N_23649,N_23570);
nand U23978 (N_23978,N_23536,N_23610);
xnor U23979 (N_23979,N_23617,N_23734);
xnor U23980 (N_23980,N_23663,N_23529);
nor U23981 (N_23981,N_23615,N_23742);
nor U23982 (N_23982,N_23561,N_23570);
xnor U23983 (N_23983,N_23540,N_23667);
nand U23984 (N_23984,N_23548,N_23692);
or U23985 (N_23985,N_23554,N_23538);
nand U23986 (N_23986,N_23612,N_23662);
or U23987 (N_23987,N_23612,N_23719);
or U23988 (N_23988,N_23653,N_23656);
or U23989 (N_23989,N_23615,N_23546);
xor U23990 (N_23990,N_23689,N_23741);
and U23991 (N_23991,N_23588,N_23584);
nor U23992 (N_23992,N_23747,N_23578);
nand U23993 (N_23993,N_23597,N_23617);
and U23994 (N_23994,N_23707,N_23662);
and U23995 (N_23995,N_23664,N_23660);
and U23996 (N_23996,N_23567,N_23583);
xnor U23997 (N_23997,N_23721,N_23618);
nand U23998 (N_23998,N_23625,N_23666);
and U23999 (N_23999,N_23603,N_23518);
or U24000 (N_24000,N_23889,N_23957);
and U24001 (N_24001,N_23997,N_23795);
nor U24002 (N_24002,N_23877,N_23875);
nand U24003 (N_24003,N_23930,N_23979);
and U24004 (N_24004,N_23782,N_23755);
and U24005 (N_24005,N_23760,N_23922);
and U24006 (N_24006,N_23793,N_23887);
and U24007 (N_24007,N_23882,N_23884);
nor U24008 (N_24008,N_23892,N_23822);
xor U24009 (N_24009,N_23871,N_23973);
nor U24010 (N_24010,N_23932,N_23766);
xnor U24011 (N_24011,N_23791,N_23975);
nor U24012 (N_24012,N_23903,N_23978);
xor U24013 (N_24013,N_23984,N_23832);
and U24014 (N_24014,N_23919,N_23788);
nor U24015 (N_24015,N_23968,N_23856);
nand U24016 (N_24016,N_23989,N_23777);
or U24017 (N_24017,N_23939,N_23977);
and U24018 (N_24018,N_23776,N_23836);
or U24019 (N_24019,N_23878,N_23900);
xor U24020 (N_24020,N_23881,N_23915);
nor U24021 (N_24021,N_23969,N_23998);
xor U24022 (N_24022,N_23931,N_23965);
and U24023 (N_24023,N_23762,N_23865);
or U24024 (N_24024,N_23792,N_23988);
nand U24025 (N_24025,N_23753,N_23918);
xnor U24026 (N_24026,N_23954,N_23775);
nand U24027 (N_24027,N_23950,N_23808);
or U24028 (N_24028,N_23761,N_23789);
xnor U24029 (N_24029,N_23839,N_23976);
and U24030 (N_24030,N_23858,N_23940);
and U24031 (N_24031,N_23847,N_23826);
nor U24032 (N_24032,N_23912,N_23840);
or U24033 (N_24033,N_23914,N_23750);
xor U24034 (N_24034,N_23809,N_23929);
nor U24035 (N_24035,N_23859,N_23860);
xnor U24036 (N_24036,N_23981,N_23904);
or U24037 (N_24037,N_23964,N_23765);
or U24038 (N_24038,N_23816,N_23815);
nand U24039 (N_24039,N_23800,N_23888);
nor U24040 (N_24040,N_23879,N_23838);
and U24041 (N_24041,N_23999,N_23995);
xor U24042 (N_24042,N_23925,N_23783);
nand U24043 (N_24043,N_23885,N_23756);
xor U24044 (N_24044,N_23844,N_23828);
or U24045 (N_24045,N_23935,N_23771);
and U24046 (N_24046,N_23786,N_23894);
and U24047 (N_24047,N_23824,N_23947);
nand U24048 (N_24048,N_23764,N_23810);
nand U24049 (N_24049,N_23936,N_23767);
nor U24050 (N_24050,N_23802,N_23942);
nand U24051 (N_24051,N_23993,N_23870);
xnor U24052 (N_24052,N_23779,N_23827);
or U24053 (N_24053,N_23924,N_23905);
or U24054 (N_24054,N_23785,N_23851);
or U24055 (N_24055,N_23898,N_23962);
or U24056 (N_24056,N_23849,N_23913);
xnor U24057 (N_24057,N_23866,N_23841);
nand U24058 (N_24058,N_23814,N_23861);
nand U24059 (N_24059,N_23843,N_23953);
nand U24060 (N_24060,N_23768,N_23926);
nor U24061 (N_24061,N_23946,N_23850);
xor U24062 (N_24062,N_23862,N_23944);
nor U24063 (N_24063,N_23829,N_23857);
or U24064 (N_24064,N_23897,N_23781);
or U24065 (N_24065,N_23833,N_23959);
and U24066 (N_24066,N_23980,N_23807);
nand U24067 (N_24067,N_23896,N_23854);
and U24068 (N_24068,N_23759,N_23992);
and U24069 (N_24069,N_23906,N_23971);
nor U24070 (N_24070,N_23873,N_23958);
and U24071 (N_24071,N_23907,N_23891);
and U24072 (N_24072,N_23769,N_23798);
nand U24073 (N_24073,N_23778,N_23961);
or U24074 (N_24074,N_23917,N_23960);
and U24075 (N_24075,N_23823,N_23845);
nor U24076 (N_24076,N_23982,N_23805);
and U24077 (N_24077,N_23763,N_23880);
nand U24078 (N_24078,N_23830,N_23883);
xor U24079 (N_24079,N_23927,N_23835);
xor U24080 (N_24080,N_23825,N_23899);
or U24081 (N_24081,N_23974,N_23752);
and U24082 (N_24082,N_23970,N_23911);
and U24083 (N_24083,N_23943,N_23801);
nor U24084 (N_24084,N_23920,N_23872);
nor U24085 (N_24085,N_23754,N_23956);
and U24086 (N_24086,N_23972,N_23901);
xnor U24087 (N_24087,N_23928,N_23831);
or U24088 (N_24088,N_23933,N_23996);
xor U24089 (N_24089,N_23908,N_23784);
or U24090 (N_24090,N_23952,N_23949);
or U24091 (N_24091,N_23987,N_23804);
nor U24092 (N_24092,N_23910,N_23813);
nand U24093 (N_24093,N_23916,N_23945);
and U24094 (N_24094,N_23853,N_23855);
and U24095 (N_24095,N_23967,N_23934);
nand U24096 (N_24096,N_23893,N_23948);
and U24097 (N_24097,N_23890,N_23821);
nand U24098 (N_24098,N_23811,N_23848);
xnor U24099 (N_24099,N_23803,N_23963);
nand U24100 (N_24100,N_23796,N_23868);
nand U24101 (N_24101,N_23797,N_23852);
xnor U24102 (N_24102,N_23770,N_23869);
and U24103 (N_24103,N_23938,N_23991);
and U24104 (N_24104,N_23990,N_23923);
xnor U24105 (N_24105,N_23909,N_23817);
or U24106 (N_24106,N_23842,N_23818);
nor U24107 (N_24107,N_23966,N_23834);
nand U24108 (N_24108,N_23955,N_23986);
nor U24109 (N_24109,N_23902,N_23864);
nand U24110 (N_24110,N_23772,N_23876);
nand U24111 (N_24111,N_23819,N_23780);
nand U24112 (N_24112,N_23794,N_23757);
xor U24113 (N_24113,N_23846,N_23874);
nand U24114 (N_24114,N_23886,N_23837);
or U24115 (N_24115,N_23773,N_23994);
xnor U24116 (N_24116,N_23895,N_23951);
nand U24117 (N_24117,N_23941,N_23774);
nor U24118 (N_24118,N_23867,N_23799);
xor U24119 (N_24119,N_23812,N_23983);
or U24120 (N_24120,N_23863,N_23751);
nor U24121 (N_24121,N_23937,N_23758);
nor U24122 (N_24122,N_23820,N_23806);
and U24123 (N_24123,N_23787,N_23790);
and U24124 (N_24124,N_23921,N_23985);
or U24125 (N_24125,N_23847,N_23810);
and U24126 (N_24126,N_23873,N_23859);
and U24127 (N_24127,N_23807,N_23996);
nand U24128 (N_24128,N_23762,N_23764);
nand U24129 (N_24129,N_23795,N_23820);
and U24130 (N_24130,N_23886,N_23852);
or U24131 (N_24131,N_23943,N_23797);
nor U24132 (N_24132,N_23836,N_23821);
nand U24133 (N_24133,N_23992,N_23954);
or U24134 (N_24134,N_23828,N_23805);
and U24135 (N_24135,N_23920,N_23834);
xor U24136 (N_24136,N_23861,N_23940);
nor U24137 (N_24137,N_23917,N_23859);
or U24138 (N_24138,N_23984,N_23943);
nor U24139 (N_24139,N_23910,N_23973);
nand U24140 (N_24140,N_23930,N_23865);
or U24141 (N_24141,N_23919,N_23902);
xor U24142 (N_24142,N_23798,N_23814);
nand U24143 (N_24143,N_23844,N_23888);
and U24144 (N_24144,N_23770,N_23971);
nor U24145 (N_24145,N_23922,N_23878);
and U24146 (N_24146,N_23794,N_23838);
xor U24147 (N_24147,N_23895,N_23884);
or U24148 (N_24148,N_23925,N_23915);
xor U24149 (N_24149,N_23919,N_23836);
xor U24150 (N_24150,N_23791,N_23950);
xor U24151 (N_24151,N_23864,N_23877);
or U24152 (N_24152,N_23982,N_23966);
and U24153 (N_24153,N_23784,N_23889);
or U24154 (N_24154,N_23831,N_23815);
and U24155 (N_24155,N_23806,N_23882);
and U24156 (N_24156,N_23832,N_23861);
nand U24157 (N_24157,N_23946,N_23860);
and U24158 (N_24158,N_23832,N_23812);
nor U24159 (N_24159,N_23891,N_23857);
nor U24160 (N_24160,N_23995,N_23784);
nand U24161 (N_24161,N_23975,N_23941);
nor U24162 (N_24162,N_23993,N_23846);
and U24163 (N_24163,N_23821,N_23790);
nor U24164 (N_24164,N_23759,N_23795);
xor U24165 (N_24165,N_23752,N_23985);
or U24166 (N_24166,N_23885,N_23769);
xor U24167 (N_24167,N_23921,N_23888);
nand U24168 (N_24168,N_23785,N_23786);
and U24169 (N_24169,N_23941,N_23845);
or U24170 (N_24170,N_23761,N_23930);
or U24171 (N_24171,N_23817,N_23778);
nor U24172 (N_24172,N_23905,N_23879);
nand U24173 (N_24173,N_23955,N_23989);
nor U24174 (N_24174,N_23944,N_23874);
nor U24175 (N_24175,N_23926,N_23850);
xor U24176 (N_24176,N_23971,N_23902);
nor U24177 (N_24177,N_23939,N_23984);
or U24178 (N_24178,N_23977,N_23761);
or U24179 (N_24179,N_23997,N_23822);
nand U24180 (N_24180,N_23778,N_23857);
and U24181 (N_24181,N_23886,N_23870);
or U24182 (N_24182,N_23796,N_23840);
nand U24183 (N_24183,N_23799,N_23939);
nor U24184 (N_24184,N_23871,N_23917);
xnor U24185 (N_24185,N_23839,N_23984);
or U24186 (N_24186,N_23818,N_23973);
nor U24187 (N_24187,N_23834,N_23757);
nand U24188 (N_24188,N_23832,N_23843);
nand U24189 (N_24189,N_23922,N_23959);
xor U24190 (N_24190,N_23774,N_23913);
xnor U24191 (N_24191,N_23986,N_23896);
or U24192 (N_24192,N_23775,N_23839);
xnor U24193 (N_24193,N_23824,N_23969);
nand U24194 (N_24194,N_23765,N_23848);
and U24195 (N_24195,N_23798,N_23927);
or U24196 (N_24196,N_23893,N_23787);
or U24197 (N_24197,N_23905,N_23883);
nor U24198 (N_24198,N_23887,N_23927);
or U24199 (N_24199,N_23886,N_23922);
nor U24200 (N_24200,N_23830,N_23944);
nor U24201 (N_24201,N_23833,N_23851);
and U24202 (N_24202,N_23821,N_23999);
and U24203 (N_24203,N_23787,N_23933);
nor U24204 (N_24204,N_23781,N_23923);
or U24205 (N_24205,N_23862,N_23890);
and U24206 (N_24206,N_23940,N_23793);
xor U24207 (N_24207,N_23814,N_23875);
nor U24208 (N_24208,N_23920,N_23919);
nor U24209 (N_24209,N_23907,N_23757);
nand U24210 (N_24210,N_23996,N_23928);
nand U24211 (N_24211,N_23899,N_23927);
xor U24212 (N_24212,N_23978,N_23913);
xnor U24213 (N_24213,N_23778,N_23982);
nor U24214 (N_24214,N_23818,N_23984);
nand U24215 (N_24215,N_23759,N_23758);
nor U24216 (N_24216,N_23862,N_23840);
or U24217 (N_24217,N_23829,N_23984);
nor U24218 (N_24218,N_23981,N_23840);
nand U24219 (N_24219,N_23768,N_23933);
or U24220 (N_24220,N_23810,N_23808);
xor U24221 (N_24221,N_23959,N_23798);
or U24222 (N_24222,N_23972,N_23898);
xor U24223 (N_24223,N_23949,N_23782);
and U24224 (N_24224,N_23973,N_23860);
nand U24225 (N_24225,N_23794,N_23961);
and U24226 (N_24226,N_23993,N_23904);
or U24227 (N_24227,N_23808,N_23932);
or U24228 (N_24228,N_23835,N_23894);
nor U24229 (N_24229,N_23910,N_23902);
nand U24230 (N_24230,N_23866,N_23752);
nand U24231 (N_24231,N_23847,N_23889);
nand U24232 (N_24232,N_23950,N_23883);
nor U24233 (N_24233,N_23954,N_23938);
nand U24234 (N_24234,N_23940,N_23758);
nand U24235 (N_24235,N_23923,N_23989);
nand U24236 (N_24236,N_23764,N_23812);
nor U24237 (N_24237,N_23763,N_23885);
xnor U24238 (N_24238,N_23795,N_23842);
or U24239 (N_24239,N_23768,N_23991);
or U24240 (N_24240,N_23806,N_23841);
nor U24241 (N_24241,N_23807,N_23816);
and U24242 (N_24242,N_23965,N_23766);
nor U24243 (N_24243,N_23808,N_23846);
and U24244 (N_24244,N_23924,N_23833);
nor U24245 (N_24245,N_23888,N_23808);
xor U24246 (N_24246,N_23922,N_23993);
nand U24247 (N_24247,N_23835,N_23869);
nand U24248 (N_24248,N_23817,N_23797);
nor U24249 (N_24249,N_23784,N_23926);
and U24250 (N_24250,N_24168,N_24078);
xnor U24251 (N_24251,N_24170,N_24045);
xor U24252 (N_24252,N_24100,N_24040);
and U24253 (N_24253,N_24212,N_24208);
nand U24254 (N_24254,N_24183,N_24176);
or U24255 (N_24255,N_24088,N_24214);
nor U24256 (N_24256,N_24188,N_24080);
nor U24257 (N_24257,N_24181,N_24167);
or U24258 (N_24258,N_24207,N_24008);
or U24259 (N_24259,N_24013,N_24115);
nor U24260 (N_24260,N_24159,N_24020);
xnor U24261 (N_24261,N_24089,N_24229);
nand U24262 (N_24262,N_24187,N_24097);
nand U24263 (N_24263,N_24099,N_24102);
nand U24264 (N_24264,N_24247,N_24063);
xor U24265 (N_24265,N_24131,N_24121);
nand U24266 (N_24266,N_24071,N_24043);
and U24267 (N_24267,N_24192,N_24226);
nand U24268 (N_24268,N_24012,N_24175);
nor U24269 (N_24269,N_24238,N_24231);
or U24270 (N_24270,N_24166,N_24036);
nor U24271 (N_24271,N_24101,N_24149);
nor U24272 (N_24272,N_24221,N_24010);
nand U24273 (N_24273,N_24191,N_24157);
nand U24274 (N_24274,N_24092,N_24179);
and U24275 (N_24275,N_24235,N_24035);
nor U24276 (N_24276,N_24246,N_24103);
nor U24277 (N_24277,N_24178,N_24085);
or U24278 (N_24278,N_24206,N_24119);
xor U24279 (N_24279,N_24185,N_24062);
or U24280 (N_24280,N_24098,N_24053);
and U24281 (N_24281,N_24233,N_24051);
or U24282 (N_24282,N_24037,N_24059);
and U24283 (N_24283,N_24054,N_24120);
nor U24284 (N_24284,N_24049,N_24032);
nor U24285 (N_24285,N_24030,N_24027);
or U24286 (N_24286,N_24164,N_24123);
xnor U24287 (N_24287,N_24160,N_24005);
nand U24288 (N_24288,N_24016,N_24107);
xor U24289 (N_24289,N_24061,N_24109);
xor U24290 (N_24290,N_24234,N_24248);
xnor U24291 (N_24291,N_24224,N_24232);
nor U24292 (N_24292,N_24028,N_24114);
and U24293 (N_24293,N_24242,N_24219);
xor U24294 (N_24294,N_24064,N_24236);
xnor U24295 (N_24295,N_24173,N_24171);
nor U24296 (N_24296,N_24111,N_24217);
nor U24297 (N_24297,N_24084,N_24155);
and U24298 (N_24298,N_24150,N_24169);
nor U24299 (N_24299,N_24218,N_24152);
or U24300 (N_24300,N_24143,N_24090);
nand U24301 (N_24301,N_24031,N_24186);
nand U24302 (N_24302,N_24108,N_24091);
xor U24303 (N_24303,N_24142,N_24244);
and U24304 (N_24304,N_24210,N_24198);
and U24305 (N_24305,N_24087,N_24135);
nand U24306 (N_24306,N_24130,N_24156);
nand U24307 (N_24307,N_24116,N_24015);
nand U24308 (N_24308,N_24237,N_24145);
nand U24309 (N_24309,N_24216,N_24113);
and U24310 (N_24310,N_24245,N_24194);
xnor U24311 (N_24311,N_24134,N_24086);
nor U24312 (N_24312,N_24039,N_24195);
or U24313 (N_24313,N_24073,N_24041);
nor U24314 (N_24314,N_24122,N_24146);
and U24315 (N_24315,N_24007,N_24048);
nor U24316 (N_24316,N_24220,N_24228);
xnor U24317 (N_24317,N_24047,N_24211);
xor U24318 (N_24318,N_24034,N_24106);
or U24319 (N_24319,N_24067,N_24069);
and U24320 (N_24320,N_24112,N_24060);
or U24321 (N_24321,N_24029,N_24204);
nor U24322 (N_24322,N_24126,N_24025);
nand U24323 (N_24323,N_24065,N_24222);
and U24324 (N_24324,N_24068,N_24105);
nor U24325 (N_24325,N_24141,N_24104);
nand U24326 (N_24326,N_24137,N_24075);
xor U24327 (N_24327,N_24074,N_24009);
nor U24328 (N_24328,N_24004,N_24243);
xor U24329 (N_24329,N_24138,N_24144);
nor U24330 (N_24330,N_24019,N_24230);
nand U24331 (N_24331,N_24077,N_24209);
nand U24332 (N_24332,N_24193,N_24096);
nor U24333 (N_24333,N_24172,N_24124);
nor U24334 (N_24334,N_24046,N_24066);
and U24335 (N_24335,N_24148,N_24021);
xor U24336 (N_24336,N_24002,N_24177);
and U24337 (N_24337,N_24117,N_24205);
and U24338 (N_24338,N_24001,N_24128);
or U24339 (N_24339,N_24165,N_24003);
and U24340 (N_24340,N_24129,N_24057);
nor U24341 (N_24341,N_24070,N_24125);
xnor U24342 (N_24342,N_24174,N_24052);
nand U24343 (N_24343,N_24038,N_24147);
and U24344 (N_24344,N_24162,N_24215);
nand U24345 (N_24345,N_24072,N_24180);
or U24346 (N_24346,N_24133,N_24026);
nand U24347 (N_24347,N_24056,N_24022);
or U24348 (N_24348,N_24095,N_24081);
nand U24349 (N_24349,N_24050,N_24190);
or U24350 (N_24350,N_24044,N_24202);
and U24351 (N_24351,N_24058,N_24240);
xor U24352 (N_24352,N_24055,N_24213);
or U24353 (N_24353,N_24163,N_24132);
or U24354 (N_24354,N_24153,N_24127);
and U24355 (N_24355,N_24024,N_24093);
xnor U24356 (N_24356,N_24000,N_24154);
xnor U24357 (N_24357,N_24158,N_24241);
xor U24358 (N_24358,N_24161,N_24201);
nor U24359 (N_24359,N_24184,N_24189);
xor U24360 (N_24360,N_24136,N_24014);
and U24361 (N_24361,N_24200,N_24006);
nor U24362 (N_24362,N_24011,N_24018);
xor U24363 (N_24363,N_24082,N_24239);
and U24364 (N_24364,N_24203,N_24023);
nand U24365 (N_24365,N_24042,N_24118);
nand U24366 (N_24366,N_24249,N_24151);
nand U24367 (N_24367,N_24140,N_24199);
and U24368 (N_24368,N_24196,N_24079);
nor U24369 (N_24369,N_24017,N_24033);
xor U24370 (N_24370,N_24110,N_24139);
nand U24371 (N_24371,N_24182,N_24227);
nor U24372 (N_24372,N_24076,N_24094);
nand U24373 (N_24373,N_24225,N_24083);
nor U24374 (N_24374,N_24197,N_24223);
xnor U24375 (N_24375,N_24152,N_24109);
and U24376 (N_24376,N_24096,N_24185);
and U24377 (N_24377,N_24167,N_24102);
xnor U24378 (N_24378,N_24138,N_24166);
nand U24379 (N_24379,N_24201,N_24002);
xor U24380 (N_24380,N_24056,N_24153);
and U24381 (N_24381,N_24180,N_24172);
nand U24382 (N_24382,N_24005,N_24067);
nand U24383 (N_24383,N_24105,N_24024);
and U24384 (N_24384,N_24096,N_24091);
and U24385 (N_24385,N_24072,N_24091);
nand U24386 (N_24386,N_24064,N_24119);
nand U24387 (N_24387,N_24129,N_24009);
and U24388 (N_24388,N_24089,N_24007);
nor U24389 (N_24389,N_24185,N_24159);
xor U24390 (N_24390,N_24133,N_24224);
nor U24391 (N_24391,N_24101,N_24238);
or U24392 (N_24392,N_24056,N_24180);
xnor U24393 (N_24393,N_24214,N_24096);
xnor U24394 (N_24394,N_24188,N_24106);
and U24395 (N_24395,N_24018,N_24006);
nand U24396 (N_24396,N_24014,N_24143);
nand U24397 (N_24397,N_24031,N_24000);
nand U24398 (N_24398,N_24151,N_24177);
nor U24399 (N_24399,N_24153,N_24052);
and U24400 (N_24400,N_24058,N_24060);
nand U24401 (N_24401,N_24146,N_24012);
and U24402 (N_24402,N_24053,N_24173);
or U24403 (N_24403,N_24152,N_24233);
and U24404 (N_24404,N_24098,N_24140);
or U24405 (N_24405,N_24080,N_24038);
nand U24406 (N_24406,N_24201,N_24179);
or U24407 (N_24407,N_24018,N_24085);
xor U24408 (N_24408,N_24131,N_24129);
nor U24409 (N_24409,N_24057,N_24218);
nand U24410 (N_24410,N_24195,N_24058);
and U24411 (N_24411,N_24064,N_24086);
nand U24412 (N_24412,N_24148,N_24245);
nand U24413 (N_24413,N_24008,N_24041);
or U24414 (N_24414,N_24237,N_24021);
nand U24415 (N_24415,N_24053,N_24236);
or U24416 (N_24416,N_24108,N_24203);
or U24417 (N_24417,N_24210,N_24161);
xnor U24418 (N_24418,N_24161,N_24079);
and U24419 (N_24419,N_24018,N_24238);
or U24420 (N_24420,N_24037,N_24089);
xnor U24421 (N_24421,N_24049,N_24201);
and U24422 (N_24422,N_24173,N_24141);
nand U24423 (N_24423,N_24242,N_24001);
and U24424 (N_24424,N_24006,N_24050);
nand U24425 (N_24425,N_24067,N_24135);
and U24426 (N_24426,N_24162,N_24013);
nand U24427 (N_24427,N_24133,N_24035);
nor U24428 (N_24428,N_24034,N_24063);
nand U24429 (N_24429,N_24101,N_24095);
xor U24430 (N_24430,N_24066,N_24074);
xnor U24431 (N_24431,N_24198,N_24021);
nand U24432 (N_24432,N_24244,N_24121);
or U24433 (N_24433,N_24062,N_24114);
or U24434 (N_24434,N_24162,N_24077);
and U24435 (N_24435,N_24241,N_24165);
nor U24436 (N_24436,N_24205,N_24149);
or U24437 (N_24437,N_24013,N_24136);
nand U24438 (N_24438,N_24177,N_24056);
xor U24439 (N_24439,N_24229,N_24230);
and U24440 (N_24440,N_24165,N_24206);
nor U24441 (N_24441,N_24024,N_24192);
and U24442 (N_24442,N_24144,N_24135);
or U24443 (N_24443,N_24173,N_24088);
and U24444 (N_24444,N_24051,N_24110);
and U24445 (N_24445,N_24115,N_24071);
or U24446 (N_24446,N_24116,N_24131);
xnor U24447 (N_24447,N_24162,N_24203);
nand U24448 (N_24448,N_24048,N_24163);
and U24449 (N_24449,N_24058,N_24026);
and U24450 (N_24450,N_24101,N_24147);
or U24451 (N_24451,N_24113,N_24139);
and U24452 (N_24452,N_24054,N_24180);
and U24453 (N_24453,N_24134,N_24103);
xnor U24454 (N_24454,N_24058,N_24150);
nand U24455 (N_24455,N_24221,N_24204);
xor U24456 (N_24456,N_24126,N_24240);
or U24457 (N_24457,N_24166,N_24230);
xor U24458 (N_24458,N_24049,N_24186);
and U24459 (N_24459,N_24071,N_24215);
nor U24460 (N_24460,N_24233,N_24178);
xor U24461 (N_24461,N_24241,N_24181);
or U24462 (N_24462,N_24090,N_24191);
nor U24463 (N_24463,N_24067,N_24073);
and U24464 (N_24464,N_24174,N_24198);
nor U24465 (N_24465,N_24205,N_24192);
xnor U24466 (N_24466,N_24132,N_24069);
nand U24467 (N_24467,N_24116,N_24207);
nor U24468 (N_24468,N_24036,N_24126);
or U24469 (N_24469,N_24022,N_24122);
nand U24470 (N_24470,N_24161,N_24119);
xor U24471 (N_24471,N_24217,N_24129);
and U24472 (N_24472,N_24140,N_24091);
nor U24473 (N_24473,N_24167,N_24205);
or U24474 (N_24474,N_24163,N_24055);
nand U24475 (N_24475,N_24008,N_24191);
or U24476 (N_24476,N_24168,N_24057);
or U24477 (N_24477,N_24229,N_24078);
nand U24478 (N_24478,N_24160,N_24072);
or U24479 (N_24479,N_24200,N_24182);
xnor U24480 (N_24480,N_24159,N_24142);
or U24481 (N_24481,N_24247,N_24157);
and U24482 (N_24482,N_24154,N_24242);
xnor U24483 (N_24483,N_24143,N_24066);
nand U24484 (N_24484,N_24033,N_24154);
nor U24485 (N_24485,N_24144,N_24229);
xor U24486 (N_24486,N_24116,N_24081);
nand U24487 (N_24487,N_24020,N_24049);
xor U24488 (N_24488,N_24228,N_24218);
xor U24489 (N_24489,N_24047,N_24232);
and U24490 (N_24490,N_24153,N_24140);
and U24491 (N_24491,N_24160,N_24135);
xor U24492 (N_24492,N_24237,N_24075);
and U24493 (N_24493,N_24071,N_24002);
nand U24494 (N_24494,N_24168,N_24035);
nand U24495 (N_24495,N_24010,N_24183);
nor U24496 (N_24496,N_24011,N_24075);
nand U24497 (N_24497,N_24219,N_24199);
nand U24498 (N_24498,N_24219,N_24094);
or U24499 (N_24499,N_24138,N_24049);
xor U24500 (N_24500,N_24422,N_24295);
nor U24501 (N_24501,N_24363,N_24250);
nand U24502 (N_24502,N_24388,N_24392);
nand U24503 (N_24503,N_24453,N_24302);
xor U24504 (N_24504,N_24452,N_24298);
nor U24505 (N_24505,N_24275,N_24371);
and U24506 (N_24506,N_24297,N_24360);
nand U24507 (N_24507,N_24425,N_24324);
nor U24508 (N_24508,N_24351,N_24310);
nor U24509 (N_24509,N_24433,N_24346);
or U24510 (N_24510,N_24447,N_24283);
and U24511 (N_24511,N_24274,N_24350);
nand U24512 (N_24512,N_24399,N_24336);
nand U24513 (N_24513,N_24349,N_24304);
and U24514 (N_24514,N_24429,N_24410);
and U24515 (N_24515,N_24467,N_24320);
and U24516 (N_24516,N_24378,N_24373);
nand U24517 (N_24517,N_24270,N_24389);
and U24518 (N_24518,N_24315,N_24454);
nand U24519 (N_24519,N_24375,N_24362);
nor U24520 (N_24520,N_24342,N_24427);
nor U24521 (N_24521,N_24394,N_24461);
or U24522 (N_24522,N_24480,N_24367);
nor U24523 (N_24523,N_24344,N_24305);
nor U24524 (N_24524,N_24299,N_24478);
or U24525 (N_24525,N_24400,N_24423);
or U24526 (N_24526,N_24280,N_24317);
nand U24527 (N_24527,N_24311,N_24476);
xnor U24528 (N_24528,N_24457,N_24323);
xor U24529 (N_24529,N_24261,N_24474);
xnor U24530 (N_24530,N_24420,N_24277);
nand U24531 (N_24531,N_24340,N_24377);
nand U24532 (N_24532,N_24408,N_24443);
and U24533 (N_24533,N_24449,N_24446);
or U24534 (N_24534,N_24286,N_24273);
nand U24535 (N_24535,N_24354,N_24418);
or U24536 (N_24536,N_24258,N_24300);
or U24537 (N_24537,N_24468,N_24257);
xnor U24538 (N_24538,N_24475,N_24495);
nor U24539 (N_24539,N_24353,N_24253);
xor U24540 (N_24540,N_24471,N_24376);
xor U24541 (N_24541,N_24439,N_24285);
or U24542 (N_24542,N_24440,N_24455);
xor U24543 (N_24543,N_24485,N_24308);
xnor U24544 (N_24544,N_24329,N_24352);
and U24545 (N_24545,N_24409,N_24290);
nand U24546 (N_24546,N_24450,N_24374);
or U24547 (N_24547,N_24322,N_24309);
nand U24548 (N_24548,N_24398,N_24364);
or U24549 (N_24549,N_24293,N_24415);
xor U24550 (N_24550,N_24251,N_24442);
nor U24551 (N_24551,N_24259,N_24424);
and U24552 (N_24552,N_24318,N_24421);
nand U24553 (N_24553,N_24490,N_24325);
or U24554 (N_24554,N_24493,N_24412);
nor U24555 (N_24555,N_24434,N_24338);
nor U24556 (N_24556,N_24444,N_24437);
xor U24557 (N_24557,N_24395,N_24460);
nand U24558 (N_24558,N_24347,N_24438);
xnor U24559 (N_24559,N_24255,N_24262);
nor U24560 (N_24560,N_24481,N_24459);
or U24561 (N_24561,N_24370,N_24428);
or U24562 (N_24562,N_24498,N_24252);
nand U24563 (N_24563,N_24432,N_24335);
xnor U24564 (N_24564,N_24333,N_24483);
nor U24565 (N_24565,N_24458,N_24281);
or U24566 (N_24566,N_24314,N_24387);
or U24567 (N_24567,N_24484,N_24489);
xor U24568 (N_24568,N_24445,N_24272);
and U24569 (N_24569,N_24345,N_24284);
nand U24570 (N_24570,N_24343,N_24355);
and U24571 (N_24571,N_24441,N_24366);
and U24572 (N_24572,N_24266,N_24403);
or U24573 (N_24573,N_24465,N_24368);
nor U24574 (N_24574,N_24451,N_24384);
nand U24575 (N_24575,N_24379,N_24321);
nor U24576 (N_24576,N_24301,N_24472);
and U24577 (N_24577,N_24369,N_24282);
and U24578 (N_24578,N_24256,N_24417);
nand U24579 (N_24579,N_24462,N_24397);
xnor U24580 (N_24580,N_24291,N_24313);
and U24581 (N_24581,N_24380,N_24276);
and U24582 (N_24582,N_24271,N_24306);
nor U24583 (N_24583,N_24348,N_24456);
nand U24584 (N_24584,N_24426,N_24341);
or U24585 (N_24585,N_24466,N_24337);
xor U24586 (N_24586,N_24332,N_24396);
or U24587 (N_24587,N_24365,N_24401);
nor U24588 (N_24588,N_24382,N_24413);
and U24589 (N_24589,N_24328,N_24307);
or U24590 (N_24590,N_24381,N_24431);
nor U24591 (N_24591,N_24269,N_24294);
xor U24592 (N_24592,N_24496,N_24319);
xnor U24593 (N_24593,N_24486,N_24267);
nor U24594 (N_24594,N_24416,N_24334);
and U24595 (N_24595,N_24435,N_24464);
or U24596 (N_24596,N_24278,N_24402);
xor U24597 (N_24597,N_24327,N_24279);
or U24598 (N_24598,N_24265,N_24386);
or U24599 (N_24599,N_24331,N_24494);
xnor U24600 (N_24600,N_24357,N_24473);
or U24601 (N_24601,N_24414,N_24470);
or U24602 (N_24602,N_24419,N_24492);
and U24603 (N_24603,N_24260,N_24263);
or U24604 (N_24604,N_24288,N_24358);
xnor U24605 (N_24605,N_24268,N_24292);
or U24606 (N_24606,N_24448,N_24463);
or U24607 (N_24607,N_24477,N_24393);
and U24608 (N_24608,N_24497,N_24296);
xor U24609 (N_24609,N_24356,N_24383);
or U24610 (N_24610,N_24287,N_24491);
nor U24611 (N_24611,N_24390,N_24482);
and U24612 (N_24612,N_24391,N_24330);
xnor U24613 (N_24613,N_24339,N_24430);
nand U24614 (N_24614,N_24479,N_24289);
and U24615 (N_24615,N_24359,N_24316);
nor U24616 (N_24616,N_24411,N_24469);
or U24617 (N_24617,N_24499,N_24436);
and U24618 (N_24618,N_24407,N_24406);
xor U24619 (N_24619,N_24404,N_24385);
nor U24620 (N_24620,N_24487,N_24488);
xor U24621 (N_24621,N_24361,N_24405);
nand U24622 (N_24622,N_24303,N_24312);
xnor U24623 (N_24623,N_24264,N_24326);
or U24624 (N_24624,N_24254,N_24372);
nor U24625 (N_24625,N_24297,N_24346);
nor U24626 (N_24626,N_24352,N_24298);
xor U24627 (N_24627,N_24420,N_24275);
or U24628 (N_24628,N_24352,N_24296);
nor U24629 (N_24629,N_24292,N_24298);
nand U24630 (N_24630,N_24404,N_24382);
and U24631 (N_24631,N_24401,N_24278);
and U24632 (N_24632,N_24409,N_24480);
nand U24633 (N_24633,N_24361,N_24444);
nor U24634 (N_24634,N_24464,N_24483);
or U24635 (N_24635,N_24336,N_24339);
and U24636 (N_24636,N_24428,N_24444);
xnor U24637 (N_24637,N_24463,N_24421);
and U24638 (N_24638,N_24497,N_24442);
and U24639 (N_24639,N_24453,N_24299);
xnor U24640 (N_24640,N_24454,N_24253);
xnor U24641 (N_24641,N_24300,N_24254);
nand U24642 (N_24642,N_24319,N_24470);
xnor U24643 (N_24643,N_24311,N_24285);
nor U24644 (N_24644,N_24472,N_24260);
and U24645 (N_24645,N_24378,N_24414);
and U24646 (N_24646,N_24317,N_24480);
xnor U24647 (N_24647,N_24278,N_24260);
nand U24648 (N_24648,N_24452,N_24279);
nor U24649 (N_24649,N_24356,N_24376);
nor U24650 (N_24650,N_24316,N_24417);
nand U24651 (N_24651,N_24350,N_24331);
nand U24652 (N_24652,N_24258,N_24432);
and U24653 (N_24653,N_24263,N_24416);
and U24654 (N_24654,N_24310,N_24343);
nand U24655 (N_24655,N_24339,N_24448);
nand U24656 (N_24656,N_24490,N_24430);
xnor U24657 (N_24657,N_24250,N_24301);
nor U24658 (N_24658,N_24324,N_24420);
and U24659 (N_24659,N_24364,N_24463);
and U24660 (N_24660,N_24421,N_24382);
nor U24661 (N_24661,N_24483,N_24365);
nand U24662 (N_24662,N_24361,N_24309);
xnor U24663 (N_24663,N_24419,N_24449);
and U24664 (N_24664,N_24471,N_24351);
and U24665 (N_24665,N_24385,N_24392);
xor U24666 (N_24666,N_24282,N_24422);
nor U24667 (N_24667,N_24494,N_24485);
or U24668 (N_24668,N_24427,N_24479);
and U24669 (N_24669,N_24434,N_24302);
nand U24670 (N_24670,N_24331,N_24455);
xor U24671 (N_24671,N_24425,N_24337);
xnor U24672 (N_24672,N_24498,N_24276);
or U24673 (N_24673,N_24391,N_24387);
nand U24674 (N_24674,N_24451,N_24443);
xnor U24675 (N_24675,N_24329,N_24414);
nand U24676 (N_24676,N_24462,N_24438);
nand U24677 (N_24677,N_24329,N_24319);
or U24678 (N_24678,N_24468,N_24370);
or U24679 (N_24679,N_24397,N_24442);
xor U24680 (N_24680,N_24440,N_24276);
and U24681 (N_24681,N_24465,N_24303);
nand U24682 (N_24682,N_24271,N_24433);
or U24683 (N_24683,N_24419,N_24381);
or U24684 (N_24684,N_24284,N_24441);
nor U24685 (N_24685,N_24335,N_24375);
nand U24686 (N_24686,N_24414,N_24440);
or U24687 (N_24687,N_24404,N_24486);
nor U24688 (N_24688,N_24444,N_24319);
and U24689 (N_24689,N_24474,N_24276);
and U24690 (N_24690,N_24417,N_24294);
nor U24691 (N_24691,N_24460,N_24492);
and U24692 (N_24692,N_24256,N_24345);
nand U24693 (N_24693,N_24302,N_24489);
nor U24694 (N_24694,N_24329,N_24362);
nand U24695 (N_24695,N_24447,N_24432);
or U24696 (N_24696,N_24354,N_24421);
or U24697 (N_24697,N_24274,N_24348);
xor U24698 (N_24698,N_24349,N_24412);
or U24699 (N_24699,N_24251,N_24277);
and U24700 (N_24700,N_24394,N_24299);
nor U24701 (N_24701,N_24497,N_24488);
or U24702 (N_24702,N_24482,N_24270);
nor U24703 (N_24703,N_24497,N_24313);
and U24704 (N_24704,N_24345,N_24496);
and U24705 (N_24705,N_24283,N_24411);
nor U24706 (N_24706,N_24350,N_24478);
and U24707 (N_24707,N_24411,N_24330);
nand U24708 (N_24708,N_24354,N_24287);
xnor U24709 (N_24709,N_24466,N_24263);
nand U24710 (N_24710,N_24253,N_24297);
or U24711 (N_24711,N_24333,N_24343);
and U24712 (N_24712,N_24254,N_24319);
nor U24713 (N_24713,N_24365,N_24441);
xnor U24714 (N_24714,N_24374,N_24386);
or U24715 (N_24715,N_24349,N_24404);
and U24716 (N_24716,N_24466,N_24256);
nand U24717 (N_24717,N_24394,N_24469);
xor U24718 (N_24718,N_24426,N_24342);
or U24719 (N_24719,N_24384,N_24402);
and U24720 (N_24720,N_24484,N_24375);
xor U24721 (N_24721,N_24253,N_24342);
and U24722 (N_24722,N_24332,N_24353);
nor U24723 (N_24723,N_24499,N_24450);
or U24724 (N_24724,N_24377,N_24338);
xor U24725 (N_24725,N_24369,N_24351);
and U24726 (N_24726,N_24416,N_24253);
nand U24727 (N_24727,N_24481,N_24494);
xnor U24728 (N_24728,N_24347,N_24293);
xor U24729 (N_24729,N_24271,N_24445);
nand U24730 (N_24730,N_24447,N_24442);
nand U24731 (N_24731,N_24349,N_24484);
or U24732 (N_24732,N_24349,N_24464);
and U24733 (N_24733,N_24382,N_24488);
nand U24734 (N_24734,N_24422,N_24318);
and U24735 (N_24735,N_24432,N_24459);
or U24736 (N_24736,N_24420,N_24364);
nand U24737 (N_24737,N_24399,N_24294);
or U24738 (N_24738,N_24439,N_24459);
or U24739 (N_24739,N_24357,N_24265);
nand U24740 (N_24740,N_24426,N_24430);
xnor U24741 (N_24741,N_24439,N_24485);
and U24742 (N_24742,N_24380,N_24385);
and U24743 (N_24743,N_24344,N_24312);
or U24744 (N_24744,N_24483,N_24454);
nor U24745 (N_24745,N_24287,N_24385);
nor U24746 (N_24746,N_24434,N_24489);
and U24747 (N_24747,N_24255,N_24315);
and U24748 (N_24748,N_24265,N_24346);
nor U24749 (N_24749,N_24295,N_24364);
or U24750 (N_24750,N_24561,N_24639);
or U24751 (N_24751,N_24592,N_24522);
or U24752 (N_24752,N_24564,N_24580);
and U24753 (N_24753,N_24654,N_24513);
and U24754 (N_24754,N_24733,N_24736);
or U24755 (N_24755,N_24610,N_24653);
nor U24756 (N_24756,N_24669,N_24576);
and U24757 (N_24757,N_24646,N_24525);
xnor U24758 (N_24758,N_24658,N_24611);
and U24759 (N_24759,N_24667,N_24633);
nor U24760 (N_24760,N_24625,N_24688);
nand U24761 (N_24761,N_24632,N_24702);
xor U24762 (N_24762,N_24503,N_24511);
xnor U24763 (N_24763,N_24683,N_24630);
xnor U24764 (N_24764,N_24607,N_24705);
xor U24765 (N_24765,N_24744,N_24699);
xor U24766 (N_24766,N_24675,N_24541);
or U24767 (N_24767,N_24520,N_24536);
nand U24768 (N_24768,N_24739,N_24720);
and U24769 (N_24769,N_24597,N_24652);
or U24770 (N_24770,N_24507,N_24602);
nor U24771 (N_24771,N_24565,N_24731);
nand U24772 (N_24772,N_24636,N_24659);
and U24773 (N_24773,N_24508,N_24663);
nand U24774 (N_24774,N_24600,N_24728);
nor U24775 (N_24775,N_24635,N_24515);
or U24776 (N_24776,N_24500,N_24505);
and U24777 (N_24777,N_24722,N_24604);
xor U24778 (N_24778,N_24535,N_24555);
xnor U24779 (N_24779,N_24634,N_24725);
xnor U24780 (N_24780,N_24714,N_24601);
xnor U24781 (N_24781,N_24517,N_24681);
xor U24782 (N_24782,N_24509,N_24599);
and U24783 (N_24783,N_24530,N_24504);
xnor U24784 (N_24784,N_24542,N_24627);
nor U24785 (N_24785,N_24587,N_24551);
and U24786 (N_24786,N_24608,N_24534);
and U24787 (N_24787,N_24672,N_24571);
nand U24788 (N_24788,N_24606,N_24735);
or U24789 (N_24789,N_24645,N_24603);
xor U24790 (N_24790,N_24543,N_24605);
nor U24791 (N_24791,N_24664,N_24749);
nor U24792 (N_24792,N_24547,N_24642);
and U24793 (N_24793,N_24506,N_24570);
nor U24794 (N_24794,N_24539,N_24510);
xnor U24795 (N_24795,N_24718,N_24629);
xor U24796 (N_24796,N_24689,N_24747);
nor U24797 (N_24797,N_24549,N_24682);
nand U24798 (N_24798,N_24719,N_24647);
and U24799 (N_24799,N_24706,N_24711);
nor U24800 (N_24800,N_24695,N_24616);
or U24801 (N_24801,N_24676,N_24540);
and U24802 (N_24802,N_24662,N_24521);
nand U24803 (N_24803,N_24566,N_24586);
and U24804 (N_24804,N_24693,N_24575);
and U24805 (N_24805,N_24697,N_24524);
nor U24806 (N_24806,N_24572,N_24716);
or U24807 (N_24807,N_24655,N_24563);
nor U24808 (N_24808,N_24648,N_24591);
nor U24809 (N_24809,N_24612,N_24643);
xor U24810 (N_24810,N_24656,N_24588);
nand U24811 (N_24811,N_24526,N_24708);
nand U24812 (N_24812,N_24567,N_24631);
xor U24813 (N_24813,N_24614,N_24569);
nor U24814 (N_24814,N_24590,N_24677);
or U24815 (N_24815,N_24723,N_24746);
or U24816 (N_24816,N_24559,N_24527);
nand U24817 (N_24817,N_24568,N_24737);
nand U24818 (N_24818,N_24637,N_24618);
nor U24819 (N_24819,N_24578,N_24715);
nand U24820 (N_24820,N_24532,N_24562);
nor U24821 (N_24821,N_24680,N_24717);
xnor U24822 (N_24822,N_24707,N_24670);
nor U24823 (N_24823,N_24742,N_24512);
or U24824 (N_24824,N_24732,N_24615);
xor U24825 (N_24825,N_24558,N_24712);
and U24826 (N_24826,N_24613,N_24721);
xnor U24827 (N_24827,N_24685,N_24514);
and U24828 (N_24828,N_24698,N_24729);
nor U24829 (N_24829,N_24640,N_24585);
and U24830 (N_24830,N_24650,N_24595);
nor U24831 (N_24831,N_24528,N_24548);
xor U24832 (N_24832,N_24589,N_24554);
and U24833 (N_24833,N_24537,N_24502);
and U24834 (N_24834,N_24665,N_24673);
xnor U24835 (N_24835,N_24678,N_24704);
nor U24836 (N_24836,N_24596,N_24727);
nand U24837 (N_24837,N_24620,N_24748);
xor U24838 (N_24838,N_24622,N_24686);
and U24839 (N_24839,N_24516,N_24560);
xor U24840 (N_24840,N_24550,N_24546);
or U24841 (N_24841,N_24734,N_24738);
nor U24842 (N_24842,N_24657,N_24660);
xor U24843 (N_24843,N_24574,N_24691);
or U24844 (N_24844,N_24726,N_24730);
nor U24845 (N_24845,N_24690,N_24679);
and U24846 (N_24846,N_24609,N_24741);
or U24847 (N_24847,N_24553,N_24619);
xnor U24848 (N_24848,N_24573,N_24649);
xor U24849 (N_24849,N_24583,N_24694);
nand U24850 (N_24850,N_24628,N_24529);
nor U24851 (N_24851,N_24556,N_24701);
nor U24852 (N_24852,N_24692,N_24696);
or U24853 (N_24853,N_24593,N_24641);
and U24854 (N_24854,N_24584,N_24724);
and U24855 (N_24855,N_24531,N_24581);
xnor U24856 (N_24856,N_24501,N_24674);
nor U24857 (N_24857,N_24661,N_24544);
and U24858 (N_24858,N_24557,N_24621);
or U24859 (N_24859,N_24617,N_24552);
xnor U24860 (N_24860,N_24709,N_24594);
or U24861 (N_24861,N_24533,N_24666);
nor U24862 (N_24862,N_24545,N_24623);
nor U24863 (N_24863,N_24644,N_24518);
xor U24864 (N_24864,N_24687,N_24638);
nand U24865 (N_24865,N_24668,N_24700);
xnor U24866 (N_24866,N_24713,N_24710);
nor U24867 (N_24867,N_24624,N_24684);
or U24868 (N_24868,N_24671,N_24582);
nand U24869 (N_24869,N_24743,N_24745);
nand U24870 (N_24870,N_24523,N_24598);
nand U24871 (N_24871,N_24651,N_24538);
and U24872 (N_24872,N_24577,N_24703);
xor U24873 (N_24873,N_24579,N_24626);
xnor U24874 (N_24874,N_24740,N_24519);
nand U24875 (N_24875,N_24736,N_24655);
nor U24876 (N_24876,N_24588,N_24684);
or U24877 (N_24877,N_24591,N_24665);
or U24878 (N_24878,N_24735,N_24585);
nand U24879 (N_24879,N_24703,N_24679);
xor U24880 (N_24880,N_24589,N_24571);
xnor U24881 (N_24881,N_24559,N_24740);
and U24882 (N_24882,N_24648,N_24596);
or U24883 (N_24883,N_24525,N_24530);
or U24884 (N_24884,N_24583,N_24607);
nand U24885 (N_24885,N_24718,N_24562);
xnor U24886 (N_24886,N_24553,N_24658);
and U24887 (N_24887,N_24612,N_24525);
or U24888 (N_24888,N_24557,N_24709);
or U24889 (N_24889,N_24675,N_24614);
nand U24890 (N_24890,N_24738,N_24697);
xnor U24891 (N_24891,N_24743,N_24541);
nand U24892 (N_24892,N_24506,N_24662);
and U24893 (N_24893,N_24526,N_24706);
nor U24894 (N_24894,N_24608,N_24570);
nor U24895 (N_24895,N_24529,N_24727);
nand U24896 (N_24896,N_24709,N_24570);
nor U24897 (N_24897,N_24523,N_24514);
or U24898 (N_24898,N_24595,N_24530);
nand U24899 (N_24899,N_24526,N_24517);
xnor U24900 (N_24900,N_24527,N_24639);
nor U24901 (N_24901,N_24735,N_24531);
and U24902 (N_24902,N_24613,N_24682);
xnor U24903 (N_24903,N_24642,N_24574);
xor U24904 (N_24904,N_24707,N_24550);
and U24905 (N_24905,N_24641,N_24736);
and U24906 (N_24906,N_24637,N_24663);
nor U24907 (N_24907,N_24719,N_24594);
nor U24908 (N_24908,N_24700,N_24592);
nor U24909 (N_24909,N_24554,N_24519);
nor U24910 (N_24910,N_24539,N_24591);
nand U24911 (N_24911,N_24647,N_24726);
xnor U24912 (N_24912,N_24521,N_24659);
nor U24913 (N_24913,N_24652,N_24593);
and U24914 (N_24914,N_24648,N_24738);
xnor U24915 (N_24915,N_24659,N_24510);
nand U24916 (N_24916,N_24642,N_24679);
or U24917 (N_24917,N_24728,N_24515);
nor U24918 (N_24918,N_24741,N_24579);
nand U24919 (N_24919,N_24726,N_24515);
nand U24920 (N_24920,N_24686,N_24541);
and U24921 (N_24921,N_24747,N_24741);
nand U24922 (N_24922,N_24502,N_24548);
and U24923 (N_24923,N_24740,N_24642);
nor U24924 (N_24924,N_24521,N_24503);
or U24925 (N_24925,N_24562,N_24545);
nand U24926 (N_24926,N_24503,N_24691);
xnor U24927 (N_24927,N_24619,N_24514);
and U24928 (N_24928,N_24568,N_24552);
or U24929 (N_24929,N_24677,N_24739);
nor U24930 (N_24930,N_24588,N_24686);
nand U24931 (N_24931,N_24522,N_24571);
and U24932 (N_24932,N_24606,N_24672);
nor U24933 (N_24933,N_24564,N_24577);
xnor U24934 (N_24934,N_24541,N_24611);
and U24935 (N_24935,N_24509,N_24733);
or U24936 (N_24936,N_24597,N_24647);
nand U24937 (N_24937,N_24686,N_24603);
nor U24938 (N_24938,N_24687,N_24553);
and U24939 (N_24939,N_24573,N_24633);
xor U24940 (N_24940,N_24526,N_24638);
xor U24941 (N_24941,N_24692,N_24520);
and U24942 (N_24942,N_24561,N_24581);
or U24943 (N_24943,N_24633,N_24719);
xor U24944 (N_24944,N_24656,N_24531);
and U24945 (N_24945,N_24706,N_24622);
xnor U24946 (N_24946,N_24591,N_24663);
and U24947 (N_24947,N_24725,N_24560);
xor U24948 (N_24948,N_24700,N_24559);
nor U24949 (N_24949,N_24593,N_24630);
and U24950 (N_24950,N_24612,N_24534);
or U24951 (N_24951,N_24624,N_24565);
or U24952 (N_24952,N_24524,N_24501);
or U24953 (N_24953,N_24583,N_24639);
nor U24954 (N_24954,N_24621,N_24588);
nor U24955 (N_24955,N_24742,N_24738);
xor U24956 (N_24956,N_24606,N_24656);
and U24957 (N_24957,N_24510,N_24742);
nor U24958 (N_24958,N_24654,N_24548);
and U24959 (N_24959,N_24577,N_24717);
and U24960 (N_24960,N_24582,N_24732);
or U24961 (N_24961,N_24579,N_24534);
or U24962 (N_24962,N_24670,N_24630);
and U24963 (N_24963,N_24500,N_24638);
xor U24964 (N_24964,N_24675,N_24660);
and U24965 (N_24965,N_24516,N_24670);
nand U24966 (N_24966,N_24689,N_24677);
nand U24967 (N_24967,N_24656,N_24591);
nor U24968 (N_24968,N_24713,N_24598);
xnor U24969 (N_24969,N_24632,N_24687);
or U24970 (N_24970,N_24645,N_24679);
and U24971 (N_24971,N_24547,N_24515);
nand U24972 (N_24972,N_24548,N_24730);
nand U24973 (N_24973,N_24697,N_24708);
nor U24974 (N_24974,N_24628,N_24566);
or U24975 (N_24975,N_24654,N_24581);
xnor U24976 (N_24976,N_24500,N_24561);
nand U24977 (N_24977,N_24520,N_24626);
xor U24978 (N_24978,N_24557,N_24715);
nand U24979 (N_24979,N_24599,N_24557);
nor U24980 (N_24980,N_24593,N_24639);
and U24981 (N_24981,N_24577,N_24649);
or U24982 (N_24982,N_24575,N_24556);
nand U24983 (N_24983,N_24549,N_24603);
nor U24984 (N_24984,N_24698,N_24533);
nor U24985 (N_24985,N_24674,N_24724);
and U24986 (N_24986,N_24726,N_24547);
nor U24987 (N_24987,N_24707,N_24526);
xnor U24988 (N_24988,N_24730,N_24538);
and U24989 (N_24989,N_24640,N_24708);
nor U24990 (N_24990,N_24542,N_24582);
xnor U24991 (N_24991,N_24694,N_24554);
and U24992 (N_24992,N_24721,N_24515);
or U24993 (N_24993,N_24614,N_24680);
nor U24994 (N_24994,N_24747,N_24677);
and U24995 (N_24995,N_24701,N_24564);
nand U24996 (N_24996,N_24748,N_24555);
and U24997 (N_24997,N_24749,N_24557);
xor U24998 (N_24998,N_24534,N_24516);
nor U24999 (N_24999,N_24749,N_24640);
or U25000 (N_25000,N_24990,N_24960);
xor U25001 (N_25001,N_24771,N_24870);
or U25002 (N_25002,N_24831,N_24933);
and U25003 (N_25003,N_24911,N_24854);
xnor U25004 (N_25004,N_24972,N_24801);
nand U25005 (N_25005,N_24765,N_24868);
or U25006 (N_25006,N_24837,N_24763);
nand U25007 (N_25007,N_24808,N_24813);
nor U25008 (N_25008,N_24910,N_24946);
and U25009 (N_25009,N_24828,N_24934);
nor U25010 (N_25010,N_24764,N_24793);
or U25011 (N_25011,N_24907,N_24884);
or U25012 (N_25012,N_24768,N_24751);
or U25013 (N_25013,N_24887,N_24973);
nand U25014 (N_25014,N_24791,N_24888);
or U25015 (N_25015,N_24799,N_24780);
xor U25016 (N_25016,N_24785,N_24878);
or U25017 (N_25017,N_24955,N_24775);
nor U25018 (N_25018,N_24805,N_24874);
xnor U25019 (N_25019,N_24957,N_24994);
or U25020 (N_25020,N_24758,N_24974);
and U25021 (N_25021,N_24985,N_24998);
xor U25022 (N_25022,N_24925,N_24851);
nand U25023 (N_25023,N_24869,N_24860);
or U25024 (N_25024,N_24915,N_24849);
or U25025 (N_25025,N_24966,N_24961);
or U25026 (N_25026,N_24850,N_24846);
xnor U25027 (N_25027,N_24830,N_24969);
nand U25028 (N_25028,N_24941,N_24761);
nor U25029 (N_25029,N_24924,N_24886);
nor U25030 (N_25030,N_24829,N_24815);
xor U25031 (N_25031,N_24893,N_24922);
nand U25032 (N_25032,N_24827,N_24783);
and U25033 (N_25033,N_24792,N_24965);
and U25034 (N_25034,N_24766,N_24947);
xor U25035 (N_25035,N_24982,N_24867);
xor U25036 (N_25036,N_24826,N_24822);
nor U25037 (N_25037,N_24920,N_24858);
and U25038 (N_25038,N_24953,N_24963);
or U25039 (N_25039,N_24834,N_24855);
or U25040 (N_25040,N_24937,N_24996);
xnor U25041 (N_25041,N_24898,N_24770);
nor U25042 (N_25042,N_24995,N_24767);
and U25043 (N_25043,N_24839,N_24984);
xor U25044 (N_25044,N_24823,N_24753);
and U25045 (N_25045,N_24916,N_24825);
xnor U25046 (N_25046,N_24913,N_24853);
and U25047 (N_25047,N_24863,N_24804);
and U25048 (N_25048,N_24809,N_24774);
nor U25049 (N_25049,N_24759,N_24890);
xnor U25050 (N_25050,N_24811,N_24781);
or U25051 (N_25051,N_24787,N_24999);
nand U25052 (N_25052,N_24824,N_24782);
or U25053 (N_25053,N_24810,N_24821);
or U25054 (N_25054,N_24776,N_24844);
and U25055 (N_25055,N_24836,N_24795);
or U25056 (N_25056,N_24798,N_24818);
nand U25057 (N_25057,N_24988,N_24896);
nor U25058 (N_25058,N_24861,N_24895);
nor U25059 (N_25059,N_24938,N_24843);
nor U25060 (N_25060,N_24772,N_24948);
and U25061 (N_25061,N_24940,N_24777);
and U25062 (N_25062,N_24908,N_24897);
and U25063 (N_25063,N_24894,N_24820);
xor U25064 (N_25064,N_24816,N_24790);
nor U25065 (N_25065,N_24930,N_24975);
nand U25066 (N_25066,N_24902,N_24891);
nor U25067 (N_25067,N_24794,N_24932);
or U25068 (N_25068,N_24862,N_24859);
or U25069 (N_25069,N_24901,N_24959);
xor U25070 (N_25070,N_24952,N_24942);
or U25071 (N_25071,N_24847,N_24812);
nor U25072 (N_25072,N_24784,N_24814);
nand U25073 (N_25073,N_24857,N_24778);
nand U25074 (N_25074,N_24904,N_24871);
or U25075 (N_25075,N_24978,N_24889);
or U25076 (N_25076,N_24944,N_24864);
nor U25077 (N_25077,N_24879,N_24945);
nor U25078 (N_25078,N_24936,N_24757);
or U25079 (N_25079,N_24865,N_24921);
or U25080 (N_25080,N_24838,N_24832);
nand U25081 (N_25081,N_24882,N_24964);
xor U25082 (N_25082,N_24866,N_24797);
xor U25083 (N_25083,N_24840,N_24773);
and U25084 (N_25084,N_24819,N_24983);
or U25085 (N_25085,N_24752,N_24923);
and U25086 (N_25086,N_24789,N_24880);
nand U25087 (N_25087,N_24873,N_24881);
nand U25088 (N_25088,N_24845,N_24992);
and U25089 (N_25089,N_24856,N_24817);
and U25090 (N_25090,N_24807,N_24926);
nor U25091 (N_25091,N_24755,N_24906);
and U25092 (N_25092,N_24919,N_24929);
or U25093 (N_25093,N_24872,N_24756);
xor U25094 (N_25094,N_24899,N_24779);
nand U25095 (N_25095,N_24842,N_24967);
nor U25096 (N_25096,N_24754,N_24962);
nand U25097 (N_25097,N_24762,N_24903);
xor U25098 (N_25098,N_24956,N_24914);
nand U25099 (N_25099,N_24987,N_24980);
xor U25100 (N_25100,N_24928,N_24788);
xnor U25101 (N_25101,N_24876,N_24769);
nand U25102 (N_25102,N_24954,N_24927);
or U25103 (N_25103,N_24917,N_24958);
or U25104 (N_25104,N_24803,N_24833);
nor U25105 (N_25105,N_24939,N_24796);
or U25106 (N_25106,N_24949,N_24993);
or U25107 (N_25107,N_24841,N_24918);
xor U25108 (N_25108,N_24935,N_24806);
xnor U25109 (N_25109,N_24883,N_24976);
xnor U25110 (N_25110,N_24981,N_24900);
and U25111 (N_25111,N_24968,N_24943);
or U25112 (N_25112,N_24802,N_24852);
and U25113 (N_25113,N_24786,N_24750);
nor U25114 (N_25114,N_24997,N_24971);
nand U25115 (N_25115,N_24931,N_24912);
or U25116 (N_25116,N_24950,N_24760);
and U25117 (N_25117,N_24892,N_24979);
xor U25118 (N_25118,N_24977,N_24877);
nor U25119 (N_25119,N_24885,N_24835);
xor U25120 (N_25120,N_24951,N_24986);
nand U25121 (N_25121,N_24991,N_24875);
nor U25122 (N_25122,N_24848,N_24909);
nand U25123 (N_25123,N_24989,N_24800);
or U25124 (N_25124,N_24905,N_24970);
and U25125 (N_25125,N_24927,N_24975);
and U25126 (N_25126,N_24938,N_24874);
or U25127 (N_25127,N_24981,N_24846);
and U25128 (N_25128,N_24795,N_24978);
xnor U25129 (N_25129,N_24837,N_24980);
and U25130 (N_25130,N_24754,N_24899);
xor U25131 (N_25131,N_24751,N_24954);
nand U25132 (N_25132,N_24913,N_24942);
xnor U25133 (N_25133,N_24810,N_24900);
xnor U25134 (N_25134,N_24932,N_24785);
xnor U25135 (N_25135,N_24816,N_24758);
nand U25136 (N_25136,N_24750,N_24963);
xnor U25137 (N_25137,N_24986,N_24791);
xnor U25138 (N_25138,N_24855,N_24753);
and U25139 (N_25139,N_24962,N_24796);
nor U25140 (N_25140,N_24763,N_24988);
nor U25141 (N_25141,N_24873,N_24867);
and U25142 (N_25142,N_24960,N_24897);
xor U25143 (N_25143,N_24828,N_24827);
nand U25144 (N_25144,N_24831,N_24949);
nor U25145 (N_25145,N_24761,N_24793);
or U25146 (N_25146,N_24766,N_24770);
nand U25147 (N_25147,N_24848,N_24870);
and U25148 (N_25148,N_24890,N_24931);
or U25149 (N_25149,N_24949,N_24862);
and U25150 (N_25150,N_24907,N_24857);
xnor U25151 (N_25151,N_24879,N_24859);
xor U25152 (N_25152,N_24968,N_24804);
nor U25153 (N_25153,N_24904,N_24984);
nand U25154 (N_25154,N_24944,N_24857);
or U25155 (N_25155,N_24975,N_24950);
and U25156 (N_25156,N_24802,N_24909);
nand U25157 (N_25157,N_24824,N_24833);
nor U25158 (N_25158,N_24940,N_24814);
nor U25159 (N_25159,N_24982,N_24781);
or U25160 (N_25160,N_24761,N_24864);
nor U25161 (N_25161,N_24779,N_24975);
nor U25162 (N_25162,N_24920,N_24905);
xnor U25163 (N_25163,N_24843,N_24785);
and U25164 (N_25164,N_24895,N_24960);
and U25165 (N_25165,N_24865,N_24824);
or U25166 (N_25166,N_24965,N_24969);
or U25167 (N_25167,N_24848,N_24759);
nor U25168 (N_25168,N_24892,N_24916);
and U25169 (N_25169,N_24922,N_24802);
nor U25170 (N_25170,N_24865,N_24840);
nor U25171 (N_25171,N_24905,N_24848);
or U25172 (N_25172,N_24995,N_24916);
nor U25173 (N_25173,N_24938,N_24924);
nor U25174 (N_25174,N_24928,N_24797);
or U25175 (N_25175,N_24954,N_24777);
and U25176 (N_25176,N_24782,N_24793);
or U25177 (N_25177,N_24865,N_24780);
or U25178 (N_25178,N_24844,N_24974);
xor U25179 (N_25179,N_24769,N_24967);
or U25180 (N_25180,N_24830,N_24825);
or U25181 (N_25181,N_24871,N_24828);
nor U25182 (N_25182,N_24917,N_24786);
nand U25183 (N_25183,N_24848,N_24802);
nor U25184 (N_25184,N_24945,N_24821);
xor U25185 (N_25185,N_24895,N_24849);
and U25186 (N_25186,N_24818,N_24885);
xor U25187 (N_25187,N_24911,N_24812);
or U25188 (N_25188,N_24844,N_24772);
xor U25189 (N_25189,N_24846,N_24921);
or U25190 (N_25190,N_24924,N_24819);
or U25191 (N_25191,N_24758,N_24959);
nor U25192 (N_25192,N_24846,N_24999);
nand U25193 (N_25193,N_24797,N_24910);
and U25194 (N_25194,N_24909,N_24884);
nand U25195 (N_25195,N_24903,N_24884);
xor U25196 (N_25196,N_24857,N_24906);
or U25197 (N_25197,N_24760,N_24955);
or U25198 (N_25198,N_24837,N_24784);
xor U25199 (N_25199,N_24826,N_24815);
nand U25200 (N_25200,N_24974,N_24755);
xor U25201 (N_25201,N_24922,N_24946);
or U25202 (N_25202,N_24877,N_24923);
or U25203 (N_25203,N_24802,N_24913);
or U25204 (N_25204,N_24775,N_24989);
nor U25205 (N_25205,N_24779,N_24823);
and U25206 (N_25206,N_24882,N_24948);
and U25207 (N_25207,N_24955,N_24773);
or U25208 (N_25208,N_24902,N_24787);
and U25209 (N_25209,N_24956,N_24766);
nor U25210 (N_25210,N_24771,N_24931);
nand U25211 (N_25211,N_24820,N_24987);
or U25212 (N_25212,N_24836,N_24883);
or U25213 (N_25213,N_24793,N_24972);
or U25214 (N_25214,N_24801,N_24960);
xnor U25215 (N_25215,N_24755,N_24891);
and U25216 (N_25216,N_24765,N_24931);
nand U25217 (N_25217,N_24957,N_24866);
nand U25218 (N_25218,N_24788,N_24885);
xor U25219 (N_25219,N_24833,N_24926);
nand U25220 (N_25220,N_24802,N_24882);
xor U25221 (N_25221,N_24908,N_24793);
or U25222 (N_25222,N_24758,N_24837);
nor U25223 (N_25223,N_24998,N_24756);
nand U25224 (N_25224,N_24899,N_24862);
or U25225 (N_25225,N_24887,N_24967);
or U25226 (N_25226,N_24985,N_24995);
and U25227 (N_25227,N_24922,N_24980);
nor U25228 (N_25228,N_24910,N_24866);
nand U25229 (N_25229,N_24951,N_24948);
and U25230 (N_25230,N_24925,N_24967);
or U25231 (N_25231,N_24997,N_24778);
nor U25232 (N_25232,N_24830,N_24918);
or U25233 (N_25233,N_24770,N_24821);
nand U25234 (N_25234,N_24887,N_24879);
and U25235 (N_25235,N_24888,N_24986);
or U25236 (N_25236,N_24760,N_24953);
xor U25237 (N_25237,N_24905,N_24786);
or U25238 (N_25238,N_24801,N_24906);
and U25239 (N_25239,N_24848,N_24977);
and U25240 (N_25240,N_24963,N_24767);
or U25241 (N_25241,N_24837,N_24805);
nor U25242 (N_25242,N_24751,N_24870);
nand U25243 (N_25243,N_24805,N_24959);
and U25244 (N_25244,N_24807,N_24769);
nand U25245 (N_25245,N_24970,N_24996);
nand U25246 (N_25246,N_24791,N_24991);
and U25247 (N_25247,N_24968,N_24967);
xor U25248 (N_25248,N_24785,N_24771);
xnor U25249 (N_25249,N_24924,N_24867);
or U25250 (N_25250,N_25007,N_25162);
or U25251 (N_25251,N_25102,N_25136);
and U25252 (N_25252,N_25079,N_25222);
xor U25253 (N_25253,N_25229,N_25129);
or U25254 (N_25254,N_25012,N_25183);
or U25255 (N_25255,N_25247,N_25072);
or U25256 (N_25256,N_25110,N_25185);
nand U25257 (N_25257,N_25161,N_25023);
xor U25258 (N_25258,N_25216,N_25074);
and U25259 (N_25259,N_25249,N_25061);
xnor U25260 (N_25260,N_25186,N_25071);
and U25261 (N_25261,N_25088,N_25121);
or U25262 (N_25262,N_25180,N_25039);
and U25263 (N_25263,N_25105,N_25215);
nor U25264 (N_25264,N_25008,N_25131);
and U25265 (N_25265,N_25073,N_25077);
xnor U25266 (N_25266,N_25067,N_25244);
xor U25267 (N_25267,N_25202,N_25094);
and U25268 (N_25268,N_25005,N_25098);
or U25269 (N_25269,N_25158,N_25238);
nand U25270 (N_25270,N_25204,N_25182);
xnor U25271 (N_25271,N_25033,N_25198);
xor U25272 (N_25272,N_25032,N_25169);
or U25273 (N_25273,N_25029,N_25047);
nand U25274 (N_25274,N_25118,N_25184);
and U25275 (N_25275,N_25196,N_25108);
and U25276 (N_25276,N_25245,N_25148);
nor U25277 (N_25277,N_25192,N_25164);
xor U25278 (N_25278,N_25209,N_25167);
xor U25279 (N_25279,N_25101,N_25201);
nor U25280 (N_25280,N_25189,N_25248);
or U25281 (N_25281,N_25052,N_25124);
xor U25282 (N_25282,N_25024,N_25165);
nor U25283 (N_25283,N_25230,N_25219);
nand U25284 (N_25284,N_25157,N_25084);
and U25285 (N_25285,N_25146,N_25078);
xnor U25286 (N_25286,N_25235,N_25090);
xnor U25287 (N_25287,N_25070,N_25091);
nor U25288 (N_25288,N_25212,N_25112);
nor U25289 (N_25289,N_25224,N_25038);
nand U25290 (N_25290,N_25120,N_25082);
xnor U25291 (N_25291,N_25087,N_25064);
xnor U25292 (N_25292,N_25114,N_25147);
nor U25293 (N_25293,N_25119,N_25065);
nor U25294 (N_25294,N_25228,N_25036);
and U25295 (N_25295,N_25031,N_25170);
xor U25296 (N_25296,N_25221,N_25037);
xor U25297 (N_25297,N_25197,N_25066);
nand U25298 (N_25298,N_25178,N_25111);
or U25299 (N_25299,N_25117,N_25203);
xnor U25300 (N_25300,N_25127,N_25016);
and U25301 (N_25301,N_25100,N_25044);
or U25302 (N_25302,N_25207,N_25188);
and U25303 (N_25303,N_25001,N_25200);
or U25304 (N_25304,N_25223,N_25145);
and U25305 (N_25305,N_25057,N_25132);
nand U25306 (N_25306,N_25050,N_25075);
nor U25307 (N_25307,N_25010,N_25191);
nand U25308 (N_25308,N_25058,N_25174);
nand U25309 (N_25309,N_25092,N_25063);
nand U25310 (N_25310,N_25195,N_25172);
or U25311 (N_25311,N_25142,N_25042);
nor U25312 (N_25312,N_25139,N_25220);
nor U25313 (N_25313,N_25159,N_25144);
and U25314 (N_25314,N_25210,N_25236);
nor U25315 (N_25315,N_25017,N_25000);
xor U25316 (N_25316,N_25237,N_25143);
and U25317 (N_25317,N_25095,N_25106);
and U25318 (N_25318,N_25034,N_25171);
or U25319 (N_25319,N_25234,N_25217);
and U25320 (N_25320,N_25128,N_25187);
nor U25321 (N_25321,N_25046,N_25243);
nor U25322 (N_25322,N_25081,N_25190);
and U25323 (N_25323,N_25014,N_25232);
xnor U25324 (N_25324,N_25048,N_25122);
xor U25325 (N_25325,N_25069,N_25151);
and U25326 (N_25326,N_25040,N_25154);
or U25327 (N_25327,N_25096,N_25093);
and U25328 (N_25328,N_25116,N_25193);
nand U25329 (N_25329,N_25126,N_25019);
xnor U25330 (N_25330,N_25076,N_25004);
nor U25331 (N_25331,N_25194,N_25115);
or U25332 (N_25332,N_25022,N_25080);
nor U25333 (N_25333,N_25213,N_25035);
nor U25334 (N_25334,N_25134,N_25242);
or U25335 (N_25335,N_25225,N_25214);
nand U25336 (N_25336,N_25059,N_25173);
nor U25337 (N_25337,N_25231,N_25141);
nand U25338 (N_25338,N_25181,N_25054);
nor U25339 (N_25339,N_25123,N_25103);
nor U25340 (N_25340,N_25113,N_25149);
or U25341 (N_25341,N_25026,N_25055);
xor U25342 (N_25342,N_25218,N_25206);
xor U25343 (N_25343,N_25138,N_25049);
or U25344 (N_25344,N_25086,N_25018);
nor U25345 (N_25345,N_25041,N_25211);
xor U25346 (N_25346,N_25099,N_25135);
xor U25347 (N_25347,N_25013,N_25163);
or U25348 (N_25348,N_25125,N_25166);
and U25349 (N_25349,N_25179,N_25107);
or U25350 (N_25350,N_25053,N_25045);
and U25351 (N_25351,N_25030,N_25227);
nor U25352 (N_25352,N_25062,N_25003);
or U25353 (N_25353,N_25177,N_25006);
nand U25354 (N_25354,N_25152,N_25085);
nand U25355 (N_25355,N_25068,N_25009);
and U25356 (N_25356,N_25020,N_25002);
nand U25357 (N_25357,N_25233,N_25025);
nand U25358 (N_25358,N_25153,N_25175);
and U25359 (N_25359,N_25137,N_25028);
or U25360 (N_25360,N_25155,N_25060);
or U25361 (N_25361,N_25130,N_25083);
nor U25362 (N_25362,N_25097,N_25109);
nor U25363 (N_25363,N_25160,N_25150);
nand U25364 (N_25364,N_25240,N_25133);
and U25365 (N_25365,N_25051,N_25241);
and U25366 (N_25366,N_25199,N_25011);
and U25367 (N_25367,N_25226,N_25089);
or U25368 (N_25368,N_25021,N_25015);
nand U25369 (N_25369,N_25027,N_25208);
nor U25370 (N_25370,N_25104,N_25140);
or U25371 (N_25371,N_25156,N_25239);
or U25372 (N_25372,N_25168,N_25043);
xor U25373 (N_25373,N_25205,N_25246);
and U25374 (N_25374,N_25176,N_25056);
and U25375 (N_25375,N_25225,N_25188);
xnor U25376 (N_25376,N_25161,N_25078);
or U25377 (N_25377,N_25055,N_25140);
xnor U25378 (N_25378,N_25235,N_25025);
and U25379 (N_25379,N_25059,N_25079);
and U25380 (N_25380,N_25056,N_25227);
and U25381 (N_25381,N_25084,N_25125);
and U25382 (N_25382,N_25122,N_25245);
nor U25383 (N_25383,N_25052,N_25160);
or U25384 (N_25384,N_25224,N_25223);
nor U25385 (N_25385,N_25101,N_25153);
and U25386 (N_25386,N_25104,N_25000);
xnor U25387 (N_25387,N_25085,N_25163);
xor U25388 (N_25388,N_25112,N_25168);
and U25389 (N_25389,N_25194,N_25183);
and U25390 (N_25390,N_25122,N_25036);
nand U25391 (N_25391,N_25150,N_25122);
xor U25392 (N_25392,N_25210,N_25212);
nand U25393 (N_25393,N_25013,N_25066);
or U25394 (N_25394,N_25139,N_25150);
nor U25395 (N_25395,N_25176,N_25061);
nand U25396 (N_25396,N_25241,N_25001);
and U25397 (N_25397,N_25115,N_25134);
xnor U25398 (N_25398,N_25050,N_25087);
and U25399 (N_25399,N_25186,N_25138);
nand U25400 (N_25400,N_25132,N_25215);
nand U25401 (N_25401,N_25225,N_25095);
nor U25402 (N_25402,N_25064,N_25117);
and U25403 (N_25403,N_25119,N_25048);
or U25404 (N_25404,N_25167,N_25058);
and U25405 (N_25405,N_25203,N_25163);
or U25406 (N_25406,N_25216,N_25200);
or U25407 (N_25407,N_25194,N_25042);
or U25408 (N_25408,N_25133,N_25002);
xnor U25409 (N_25409,N_25013,N_25237);
nand U25410 (N_25410,N_25202,N_25148);
or U25411 (N_25411,N_25056,N_25223);
and U25412 (N_25412,N_25246,N_25147);
or U25413 (N_25413,N_25005,N_25061);
or U25414 (N_25414,N_25135,N_25078);
and U25415 (N_25415,N_25243,N_25157);
and U25416 (N_25416,N_25194,N_25076);
or U25417 (N_25417,N_25248,N_25222);
nand U25418 (N_25418,N_25070,N_25128);
or U25419 (N_25419,N_25121,N_25076);
and U25420 (N_25420,N_25017,N_25068);
or U25421 (N_25421,N_25181,N_25006);
nand U25422 (N_25422,N_25070,N_25060);
nor U25423 (N_25423,N_25113,N_25026);
or U25424 (N_25424,N_25119,N_25033);
or U25425 (N_25425,N_25027,N_25047);
and U25426 (N_25426,N_25238,N_25046);
nor U25427 (N_25427,N_25174,N_25140);
or U25428 (N_25428,N_25040,N_25048);
nand U25429 (N_25429,N_25179,N_25140);
xor U25430 (N_25430,N_25023,N_25110);
nor U25431 (N_25431,N_25225,N_25099);
and U25432 (N_25432,N_25207,N_25198);
nand U25433 (N_25433,N_25130,N_25094);
or U25434 (N_25434,N_25241,N_25032);
xor U25435 (N_25435,N_25181,N_25095);
and U25436 (N_25436,N_25006,N_25079);
and U25437 (N_25437,N_25166,N_25049);
xnor U25438 (N_25438,N_25118,N_25139);
nand U25439 (N_25439,N_25095,N_25147);
nand U25440 (N_25440,N_25227,N_25168);
or U25441 (N_25441,N_25122,N_25038);
and U25442 (N_25442,N_25248,N_25054);
or U25443 (N_25443,N_25156,N_25021);
nor U25444 (N_25444,N_25204,N_25113);
nand U25445 (N_25445,N_25000,N_25119);
nand U25446 (N_25446,N_25045,N_25131);
nor U25447 (N_25447,N_25200,N_25218);
or U25448 (N_25448,N_25169,N_25083);
xnor U25449 (N_25449,N_25052,N_25240);
or U25450 (N_25450,N_25058,N_25020);
xor U25451 (N_25451,N_25102,N_25194);
nor U25452 (N_25452,N_25011,N_25239);
or U25453 (N_25453,N_25105,N_25003);
and U25454 (N_25454,N_25130,N_25098);
and U25455 (N_25455,N_25174,N_25033);
nor U25456 (N_25456,N_25161,N_25108);
xor U25457 (N_25457,N_25082,N_25123);
nor U25458 (N_25458,N_25210,N_25015);
xor U25459 (N_25459,N_25157,N_25223);
and U25460 (N_25460,N_25127,N_25086);
xor U25461 (N_25461,N_25092,N_25045);
or U25462 (N_25462,N_25055,N_25062);
nand U25463 (N_25463,N_25131,N_25117);
xnor U25464 (N_25464,N_25143,N_25153);
nor U25465 (N_25465,N_25141,N_25225);
and U25466 (N_25466,N_25084,N_25107);
or U25467 (N_25467,N_25187,N_25070);
nor U25468 (N_25468,N_25122,N_25151);
and U25469 (N_25469,N_25234,N_25205);
nor U25470 (N_25470,N_25115,N_25023);
nor U25471 (N_25471,N_25189,N_25007);
xnor U25472 (N_25472,N_25120,N_25046);
nor U25473 (N_25473,N_25220,N_25056);
nor U25474 (N_25474,N_25202,N_25161);
or U25475 (N_25475,N_25191,N_25144);
nor U25476 (N_25476,N_25078,N_25029);
nor U25477 (N_25477,N_25073,N_25186);
xor U25478 (N_25478,N_25047,N_25026);
nor U25479 (N_25479,N_25171,N_25138);
xor U25480 (N_25480,N_25144,N_25114);
xnor U25481 (N_25481,N_25085,N_25141);
nand U25482 (N_25482,N_25194,N_25054);
xor U25483 (N_25483,N_25052,N_25175);
xor U25484 (N_25484,N_25222,N_25197);
and U25485 (N_25485,N_25031,N_25216);
nor U25486 (N_25486,N_25023,N_25240);
nand U25487 (N_25487,N_25052,N_25008);
nor U25488 (N_25488,N_25089,N_25245);
nor U25489 (N_25489,N_25090,N_25007);
nor U25490 (N_25490,N_25092,N_25224);
xor U25491 (N_25491,N_25137,N_25175);
nand U25492 (N_25492,N_25206,N_25249);
and U25493 (N_25493,N_25024,N_25197);
or U25494 (N_25494,N_25006,N_25062);
nand U25495 (N_25495,N_25249,N_25023);
xor U25496 (N_25496,N_25088,N_25078);
xnor U25497 (N_25497,N_25124,N_25109);
or U25498 (N_25498,N_25019,N_25246);
and U25499 (N_25499,N_25094,N_25027);
or U25500 (N_25500,N_25337,N_25385);
xnor U25501 (N_25501,N_25396,N_25281);
xor U25502 (N_25502,N_25355,N_25300);
nand U25503 (N_25503,N_25394,N_25305);
nor U25504 (N_25504,N_25349,N_25313);
nor U25505 (N_25505,N_25301,N_25443);
nor U25506 (N_25506,N_25436,N_25321);
nand U25507 (N_25507,N_25272,N_25354);
xor U25508 (N_25508,N_25324,N_25418);
or U25509 (N_25509,N_25253,N_25452);
or U25510 (N_25510,N_25286,N_25306);
nand U25511 (N_25511,N_25378,N_25490);
nand U25512 (N_25512,N_25271,N_25402);
xor U25513 (N_25513,N_25362,N_25296);
nand U25514 (N_25514,N_25339,N_25345);
nand U25515 (N_25515,N_25414,N_25471);
and U25516 (N_25516,N_25417,N_25426);
nor U25517 (N_25517,N_25343,N_25450);
nor U25518 (N_25518,N_25404,N_25274);
nand U25519 (N_25519,N_25309,N_25425);
nand U25520 (N_25520,N_25423,N_25477);
xor U25521 (N_25521,N_25461,N_25468);
or U25522 (N_25522,N_25327,N_25481);
or U25523 (N_25523,N_25469,N_25416);
nor U25524 (N_25524,N_25380,N_25252);
or U25525 (N_25525,N_25428,N_25370);
xnor U25526 (N_25526,N_25392,N_25284);
or U25527 (N_25527,N_25486,N_25429);
nor U25528 (N_25528,N_25265,N_25434);
xor U25529 (N_25529,N_25475,N_25444);
or U25530 (N_25530,N_25361,N_25371);
nor U25531 (N_25531,N_25283,N_25441);
xor U25532 (N_25532,N_25270,N_25479);
xor U25533 (N_25533,N_25432,N_25433);
xor U25534 (N_25534,N_25364,N_25328);
or U25535 (N_25535,N_25374,N_25420);
or U25536 (N_25536,N_25269,N_25334);
nor U25537 (N_25537,N_25310,N_25470);
nand U25538 (N_25538,N_25408,N_25489);
nor U25539 (N_25539,N_25323,N_25366);
or U25540 (N_25540,N_25464,N_25255);
nand U25541 (N_25541,N_25393,N_25480);
nand U25542 (N_25542,N_25390,N_25297);
and U25543 (N_25543,N_25340,N_25491);
xnor U25544 (N_25544,N_25291,N_25250);
xnor U25545 (N_25545,N_25344,N_25400);
and U25546 (N_25546,N_25497,N_25419);
xnor U25547 (N_25547,N_25303,N_25256);
and U25548 (N_25548,N_25446,N_25280);
and U25549 (N_25549,N_25311,N_25463);
or U25550 (N_25550,N_25412,N_25482);
nor U25551 (N_25551,N_25391,N_25381);
xor U25552 (N_25552,N_25346,N_25267);
nand U25553 (N_25553,N_25478,N_25290);
nand U25554 (N_25554,N_25424,N_25447);
or U25555 (N_25555,N_25262,N_25317);
nor U25556 (N_25556,N_25437,N_25495);
xnor U25557 (N_25557,N_25473,N_25388);
xnor U25558 (N_25558,N_25263,N_25466);
and U25559 (N_25559,N_25496,N_25278);
or U25560 (N_25560,N_25294,N_25376);
or U25561 (N_25561,N_25457,N_25401);
and U25562 (N_25562,N_25445,N_25435);
nor U25563 (N_25563,N_25289,N_25360);
and U25564 (N_25564,N_25372,N_25282);
nand U25565 (N_25565,N_25389,N_25483);
or U25566 (N_25566,N_25375,N_25329);
and U25567 (N_25567,N_25422,N_25460);
xor U25568 (N_25568,N_25409,N_25314);
and U25569 (N_25569,N_25369,N_25459);
xnor U25570 (N_25570,N_25356,N_25330);
xor U25571 (N_25571,N_25405,N_25277);
nand U25572 (N_25572,N_25476,N_25387);
and U25573 (N_25573,N_25413,N_25307);
and U25574 (N_25574,N_25279,N_25285);
and U25575 (N_25575,N_25302,N_25351);
xor U25576 (N_25576,N_25308,N_25273);
nor U25577 (N_25577,N_25384,N_25421);
nor U25578 (N_25578,N_25295,N_25315);
nor U25579 (N_25579,N_25368,N_25318);
nand U25580 (N_25580,N_25411,N_25275);
nand U25581 (N_25581,N_25465,N_25451);
xnor U25582 (N_25582,N_25403,N_25431);
nand U25583 (N_25583,N_25494,N_25347);
xnor U25584 (N_25584,N_25427,N_25298);
nor U25585 (N_25585,N_25454,N_25304);
nor U25586 (N_25586,N_25474,N_25485);
xor U25587 (N_25587,N_25292,N_25325);
or U25588 (N_25588,N_25397,N_25365);
nor U25589 (N_25589,N_25348,N_25493);
or U25590 (N_25590,N_25319,N_25449);
xnor U25591 (N_25591,N_25350,N_25439);
nor U25592 (N_25592,N_25326,N_25410);
xnor U25593 (N_25593,N_25462,N_25373);
nand U25594 (N_25594,N_25382,N_25257);
nor U25595 (N_25595,N_25498,N_25320);
or U25596 (N_25596,N_25288,N_25338);
or U25597 (N_25597,N_25442,N_25342);
or U25598 (N_25598,N_25287,N_25458);
xnor U25599 (N_25599,N_25331,N_25430);
xnor U25600 (N_25600,N_25448,N_25259);
and U25601 (N_25601,N_25359,N_25335);
nand U25602 (N_25602,N_25264,N_25488);
or U25603 (N_25603,N_25261,N_25332);
and U25604 (N_25604,N_25336,N_25440);
and U25605 (N_25605,N_25484,N_25316);
or U25606 (N_25606,N_25386,N_25254);
or U25607 (N_25607,N_25299,N_25398);
nor U25608 (N_25608,N_25455,N_25341);
nand U25609 (N_25609,N_25453,N_25438);
or U25610 (N_25610,N_25492,N_25415);
nand U25611 (N_25611,N_25352,N_25467);
nor U25612 (N_25612,N_25456,N_25333);
nor U25613 (N_25613,N_25487,N_25395);
nor U25614 (N_25614,N_25251,N_25268);
and U25615 (N_25615,N_25358,N_25406);
nand U25616 (N_25616,N_25363,N_25399);
xor U25617 (N_25617,N_25322,N_25499);
nor U25618 (N_25618,N_25377,N_25353);
nand U25619 (N_25619,N_25293,N_25312);
or U25620 (N_25620,N_25472,N_25266);
and U25621 (N_25621,N_25379,N_25367);
nand U25622 (N_25622,N_25276,N_25407);
and U25623 (N_25623,N_25383,N_25258);
or U25624 (N_25624,N_25260,N_25357);
xnor U25625 (N_25625,N_25448,N_25306);
xor U25626 (N_25626,N_25367,N_25343);
or U25627 (N_25627,N_25461,N_25276);
and U25628 (N_25628,N_25366,N_25339);
nand U25629 (N_25629,N_25451,N_25476);
nand U25630 (N_25630,N_25420,N_25284);
xnor U25631 (N_25631,N_25364,N_25393);
xnor U25632 (N_25632,N_25302,N_25257);
or U25633 (N_25633,N_25281,N_25440);
nor U25634 (N_25634,N_25342,N_25304);
or U25635 (N_25635,N_25402,N_25277);
nand U25636 (N_25636,N_25311,N_25280);
xor U25637 (N_25637,N_25326,N_25313);
and U25638 (N_25638,N_25449,N_25365);
or U25639 (N_25639,N_25429,N_25319);
xnor U25640 (N_25640,N_25329,N_25382);
xnor U25641 (N_25641,N_25277,N_25471);
or U25642 (N_25642,N_25406,N_25467);
nor U25643 (N_25643,N_25483,N_25373);
xnor U25644 (N_25644,N_25259,N_25378);
xnor U25645 (N_25645,N_25328,N_25411);
nand U25646 (N_25646,N_25371,N_25496);
or U25647 (N_25647,N_25313,N_25280);
or U25648 (N_25648,N_25470,N_25442);
and U25649 (N_25649,N_25371,N_25440);
and U25650 (N_25650,N_25322,N_25430);
nand U25651 (N_25651,N_25322,N_25425);
nand U25652 (N_25652,N_25319,N_25361);
xor U25653 (N_25653,N_25388,N_25307);
nor U25654 (N_25654,N_25410,N_25370);
or U25655 (N_25655,N_25457,N_25267);
and U25656 (N_25656,N_25343,N_25428);
and U25657 (N_25657,N_25262,N_25320);
xnor U25658 (N_25658,N_25371,N_25336);
or U25659 (N_25659,N_25377,N_25432);
xor U25660 (N_25660,N_25330,N_25416);
or U25661 (N_25661,N_25373,N_25411);
nand U25662 (N_25662,N_25343,N_25290);
or U25663 (N_25663,N_25298,N_25287);
and U25664 (N_25664,N_25477,N_25262);
nand U25665 (N_25665,N_25472,N_25455);
nand U25666 (N_25666,N_25379,N_25486);
nand U25667 (N_25667,N_25468,N_25449);
and U25668 (N_25668,N_25265,N_25303);
nand U25669 (N_25669,N_25336,N_25294);
nor U25670 (N_25670,N_25323,N_25441);
or U25671 (N_25671,N_25298,N_25381);
and U25672 (N_25672,N_25265,N_25332);
and U25673 (N_25673,N_25490,N_25390);
or U25674 (N_25674,N_25444,N_25326);
nand U25675 (N_25675,N_25432,N_25471);
nor U25676 (N_25676,N_25367,N_25336);
nand U25677 (N_25677,N_25445,N_25358);
nor U25678 (N_25678,N_25265,N_25496);
or U25679 (N_25679,N_25419,N_25305);
xnor U25680 (N_25680,N_25470,N_25297);
nand U25681 (N_25681,N_25474,N_25267);
and U25682 (N_25682,N_25302,N_25316);
nand U25683 (N_25683,N_25428,N_25306);
or U25684 (N_25684,N_25277,N_25279);
xnor U25685 (N_25685,N_25457,N_25279);
nor U25686 (N_25686,N_25487,N_25255);
xor U25687 (N_25687,N_25350,N_25289);
and U25688 (N_25688,N_25494,N_25453);
or U25689 (N_25689,N_25466,N_25403);
nand U25690 (N_25690,N_25472,N_25262);
xnor U25691 (N_25691,N_25340,N_25324);
and U25692 (N_25692,N_25447,N_25340);
xnor U25693 (N_25693,N_25303,N_25458);
and U25694 (N_25694,N_25266,N_25256);
and U25695 (N_25695,N_25468,N_25392);
nor U25696 (N_25696,N_25383,N_25302);
nor U25697 (N_25697,N_25283,N_25285);
nand U25698 (N_25698,N_25490,N_25412);
nand U25699 (N_25699,N_25388,N_25341);
nand U25700 (N_25700,N_25452,N_25377);
nand U25701 (N_25701,N_25299,N_25447);
and U25702 (N_25702,N_25397,N_25377);
nand U25703 (N_25703,N_25443,N_25409);
xor U25704 (N_25704,N_25447,N_25423);
nor U25705 (N_25705,N_25453,N_25327);
nor U25706 (N_25706,N_25338,N_25401);
and U25707 (N_25707,N_25497,N_25465);
nor U25708 (N_25708,N_25363,N_25264);
and U25709 (N_25709,N_25403,N_25470);
or U25710 (N_25710,N_25461,N_25273);
and U25711 (N_25711,N_25308,N_25361);
and U25712 (N_25712,N_25363,N_25270);
or U25713 (N_25713,N_25418,N_25290);
and U25714 (N_25714,N_25352,N_25460);
nor U25715 (N_25715,N_25436,N_25294);
nand U25716 (N_25716,N_25432,N_25498);
or U25717 (N_25717,N_25322,N_25361);
nor U25718 (N_25718,N_25384,N_25372);
nand U25719 (N_25719,N_25305,N_25351);
and U25720 (N_25720,N_25365,N_25373);
and U25721 (N_25721,N_25269,N_25407);
or U25722 (N_25722,N_25372,N_25278);
xor U25723 (N_25723,N_25263,N_25287);
or U25724 (N_25724,N_25497,N_25476);
nor U25725 (N_25725,N_25339,N_25484);
nand U25726 (N_25726,N_25387,N_25440);
xnor U25727 (N_25727,N_25298,N_25499);
xor U25728 (N_25728,N_25432,N_25282);
xor U25729 (N_25729,N_25369,N_25350);
xnor U25730 (N_25730,N_25342,N_25298);
nand U25731 (N_25731,N_25438,N_25345);
xor U25732 (N_25732,N_25449,N_25273);
nand U25733 (N_25733,N_25443,N_25355);
and U25734 (N_25734,N_25478,N_25408);
nor U25735 (N_25735,N_25339,N_25388);
nand U25736 (N_25736,N_25326,N_25403);
and U25737 (N_25737,N_25251,N_25451);
xor U25738 (N_25738,N_25324,N_25300);
nor U25739 (N_25739,N_25387,N_25366);
and U25740 (N_25740,N_25483,N_25319);
nand U25741 (N_25741,N_25494,N_25378);
nor U25742 (N_25742,N_25478,N_25293);
or U25743 (N_25743,N_25431,N_25251);
and U25744 (N_25744,N_25250,N_25483);
or U25745 (N_25745,N_25332,N_25443);
nand U25746 (N_25746,N_25444,N_25262);
and U25747 (N_25747,N_25393,N_25427);
xor U25748 (N_25748,N_25364,N_25322);
nor U25749 (N_25749,N_25403,N_25284);
and U25750 (N_25750,N_25619,N_25692);
nand U25751 (N_25751,N_25641,N_25521);
xnor U25752 (N_25752,N_25588,N_25600);
or U25753 (N_25753,N_25735,N_25640);
or U25754 (N_25754,N_25550,N_25651);
xnor U25755 (N_25755,N_25517,N_25618);
xor U25756 (N_25756,N_25511,N_25516);
xor U25757 (N_25757,N_25504,N_25734);
or U25758 (N_25758,N_25644,N_25688);
and U25759 (N_25759,N_25732,N_25746);
xnor U25760 (N_25760,N_25663,N_25534);
nand U25761 (N_25761,N_25599,N_25646);
xnor U25762 (N_25762,N_25724,N_25675);
xor U25763 (N_25763,N_25537,N_25706);
and U25764 (N_25764,N_25736,N_25636);
or U25765 (N_25765,N_25514,N_25681);
nor U25766 (N_25766,N_25500,N_25566);
nor U25767 (N_25767,N_25728,N_25507);
and U25768 (N_25768,N_25505,N_25589);
xnor U25769 (N_25769,N_25623,N_25743);
and U25770 (N_25770,N_25551,N_25571);
nor U25771 (N_25771,N_25614,N_25567);
and U25772 (N_25772,N_25520,N_25649);
xnor U25773 (N_25773,N_25526,N_25601);
and U25774 (N_25774,N_25635,N_25607);
or U25775 (N_25775,N_25669,N_25563);
and U25776 (N_25776,N_25524,N_25535);
nor U25777 (N_25777,N_25695,N_25667);
nor U25778 (N_25778,N_25683,N_25592);
and U25779 (N_25779,N_25586,N_25522);
nand U25780 (N_25780,N_25654,N_25733);
xor U25781 (N_25781,N_25596,N_25605);
and U25782 (N_25782,N_25701,N_25593);
nor U25783 (N_25783,N_25525,N_25530);
xor U25784 (N_25784,N_25506,N_25615);
and U25785 (N_25785,N_25647,N_25634);
nand U25786 (N_25786,N_25538,N_25722);
or U25787 (N_25787,N_25559,N_25719);
nor U25788 (N_25788,N_25503,N_25708);
nor U25789 (N_25789,N_25632,N_25591);
and U25790 (N_25790,N_25590,N_25747);
nor U25791 (N_25791,N_25502,N_25631);
nor U25792 (N_25792,N_25715,N_25568);
xnor U25793 (N_25793,N_25740,N_25585);
and U25794 (N_25794,N_25533,N_25532);
or U25795 (N_25795,N_25622,N_25693);
nand U25796 (N_25796,N_25687,N_25717);
or U25797 (N_25797,N_25513,N_25528);
or U25798 (N_25798,N_25529,N_25670);
xnor U25799 (N_25799,N_25645,N_25575);
nor U25800 (N_25800,N_25677,N_25749);
or U25801 (N_25801,N_25540,N_25582);
nand U25802 (N_25802,N_25612,N_25531);
or U25803 (N_25803,N_25725,N_25512);
and U25804 (N_25804,N_25657,N_25579);
nor U25805 (N_25805,N_25737,N_25527);
and U25806 (N_25806,N_25674,N_25616);
nor U25807 (N_25807,N_25698,N_25696);
nand U25808 (N_25808,N_25709,N_25625);
nor U25809 (N_25809,N_25628,N_25546);
xor U25810 (N_25810,N_25689,N_25569);
or U25811 (N_25811,N_25672,N_25621);
xor U25812 (N_25812,N_25574,N_25630);
nand U25813 (N_25813,N_25656,N_25572);
nor U25814 (N_25814,N_25597,N_25738);
or U25815 (N_25815,N_25665,N_25716);
and U25816 (N_25816,N_25523,N_25509);
nand U25817 (N_25817,N_25552,N_25661);
nor U25818 (N_25818,N_25720,N_25570);
or U25819 (N_25819,N_25565,N_25730);
or U25820 (N_25820,N_25723,N_25686);
xnor U25821 (N_25821,N_25518,N_25560);
and U25822 (N_25822,N_25648,N_25680);
xnor U25823 (N_25823,N_25668,N_25684);
xor U25824 (N_25824,N_25658,N_25713);
nand U25825 (N_25825,N_25594,N_25595);
nand U25826 (N_25826,N_25555,N_25633);
or U25827 (N_25827,N_25745,N_25620);
and U25828 (N_25828,N_25710,N_25554);
and U25829 (N_25829,N_25690,N_25659);
nand U25830 (N_25830,N_25598,N_25515);
xnor U25831 (N_25831,N_25548,N_25697);
nor U25832 (N_25832,N_25731,N_25627);
nand U25833 (N_25833,N_25671,N_25610);
xnor U25834 (N_25834,N_25536,N_25666);
xor U25835 (N_25835,N_25539,N_25583);
nand U25836 (N_25836,N_25662,N_25682);
or U25837 (N_25837,N_25609,N_25573);
or U25838 (N_25838,N_25545,N_25718);
xnor U25839 (N_25839,N_25603,N_25748);
and U25840 (N_25840,N_25653,N_25660);
nand U25841 (N_25841,N_25557,N_25700);
or U25842 (N_25842,N_25519,N_25711);
xnor U25843 (N_25843,N_25544,N_25727);
xor U25844 (N_25844,N_25637,N_25744);
xor U25845 (N_25845,N_25562,N_25664);
xnor U25846 (N_25846,N_25611,N_25650);
and U25847 (N_25847,N_25705,N_25655);
or U25848 (N_25848,N_25608,N_25542);
nor U25849 (N_25849,N_25587,N_25606);
or U25850 (N_25850,N_25564,N_25577);
and U25851 (N_25851,N_25617,N_25604);
xnor U25852 (N_25852,N_25629,N_25742);
nor U25853 (N_25853,N_25643,N_25676);
nand U25854 (N_25854,N_25741,N_25613);
or U25855 (N_25855,N_25576,N_25626);
nor U25856 (N_25856,N_25549,N_25714);
nand U25857 (N_25857,N_25624,N_25602);
nor U25858 (N_25858,N_25510,N_25699);
nand U25859 (N_25859,N_25556,N_25721);
nand U25860 (N_25860,N_25561,N_25726);
nand U25861 (N_25861,N_25691,N_25679);
or U25862 (N_25862,N_25642,N_25580);
and U25863 (N_25863,N_25547,N_25685);
nor U25864 (N_25864,N_25673,N_25678);
or U25865 (N_25865,N_25543,N_25652);
and U25866 (N_25866,N_25541,N_25704);
or U25867 (N_25867,N_25578,N_25553);
nand U25868 (N_25868,N_25739,N_25729);
nor U25869 (N_25869,N_25638,N_25584);
or U25870 (N_25870,N_25712,N_25702);
nor U25871 (N_25871,N_25508,N_25501);
or U25872 (N_25872,N_25581,N_25639);
nand U25873 (N_25873,N_25558,N_25703);
and U25874 (N_25874,N_25694,N_25707);
and U25875 (N_25875,N_25683,N_25710);
xor U25876 (N_25876,N_25514,N_25672);
or U25877 (N_25877,N_25736,N_25540);
and U25878 (N_25878,N_25505,N_25610);
or U25879 (N_25879,N_25687,N_25748);
nand U25880 (N_25880,N_25521,N_25522);
nand U25881 (N_25881,N_25641,N_25704);
and U25882 (N_25882,N_25683,N_25680);
or U25883 (N_25883,N_25679,N_25573);
nand U25884 (N_25884,N_25573,N_25731);
xor U25885 (N_25885,N_25505,N_25515);
nand U25886 (N_25886,N_25597,N_25630);
or U25887 (N_25887,N_25589,N_25748);
xor U25888 (N_25888,N_25655,N_25547);
xnor U25889 (N_25889,N_25558,N_25571);
and U25890 (N_25890,N_25683,N_25724);
nor U25891 (N_25891,N_25609,N_25743);
and U25892 (N_25892,N_25627,N_25684);
and U25893 (N_25893,N_25748,N_25647);
nor U25894 (N_25894,N_25688,N_25571);
xor U25895 (N_25895,N_25661,N_25601);
nand U25896 (N_25896,N_25639,N_25524);
xor U25897 (N_25897,N_25546,N_25722);
xor U25898 (N_25898,N_25587,N_25650);
nand U25899 (N_25899,N_25606,N_25558);
nand U25900 (N_25900,N_25587,N_25749);
or U25901 (N_25901,N_25701,N_25559);
xnor U25902 (N_25902,N_25552,N_25684);
xnor U25903 (N_25903,N_25665,N_25545);
nor U25904 (N_25904,N_25573,N_25621);
nand U25905 (N_25905,N_25661,N_25707);
xor U25906 (N_25906,N_25622,N_25696);
or U25907 (N_25907,N_25615,N_25719);
nand U25908 (N_25908,N_25571,N_25722);
xor U25909 (N_25909,N_25557,N_25609);
or U25910 (N_25910,N_25553,N_25741);
nand U25911 (N_25911,N_25651,N_25571);
nand U25912 (N_25912,N_25625,N_25679);
nand U25913 (N_25913,N_25611,N_25627);
nand U25914 (N_25914,N_25564,N_25586);
nand U25915 (N_25915,N_25696,N_25584);
xor U25916 (N_25916,N_25719,N_25500);
xor U25917 (N_25917,N_25710,N_25690);
xor U25918 (N_25918,N_25538,N_25646);
nor U25919 (N_25919,N_25653,N_25534);
or U25920 (N_25920,N_25671,N_25605);
nor U25921 (N_25921,N_25621,N_25583);
nand U25922 (N_25922,N_25630,N_25563);
nand U25923 (N_25923,N_25693,N_25666);
and U25924 (N_25924,N_25634,N_25729);
nor U25925 (N_25925,N_25540,N_25618);
xnor U25926 (N_25926,N_25742,N_25544);
nor U25927 (N_25927,N_25604,N_25566);
or U25928 (N_25928,N_25676,N_25647);
and U25929 (N_25929,N_25668,N_25674);
or U25930 (N_25930,N_25542,N_25678);
nor U25931 (N_25931,N_25572,N_25662);
xnor U25932 (N_25932,N_25631,N_25671);
nor U25933 (N_25933,N_25544,N_25716);
and U25934 (N_25934,N_25605,N_25638);
or U25935 (N_25935,N_25604,N_25511);
nand U25936 (N_25936,N_25734,N_25506);
nor U25937 (N_25937,N_25540,N_25524);
and U25938 (N_25938,N_25643,N_25633);
nor U25939 (N_25939,N_25561,N_25679);
xor U25940 (N_25940,N_25716,N_25641);
nand U25941 (N_25941,N_25621,N_25535);
nor U25942 (N_25942,N_25596,N_25581);
or U25943 (N_25943,N_25651,N_25609);
or U25944 (N_25944,N_25538,N_25674);
xnor U25945 (N_25945,N_25573,N_25702);
nor U25946 (N_25946,N_25544,N_25539);
or U25947 (N_25947,N_25706,N_25500);
nand U25948 (N_25948,N_25552,N_25633);
nor U25949 (N_25949,N_25651,N_25542);
xor U25950 (N_25950,N_25510,N_25690);
xor U25951 (N_25951,N_25534,N_25705);
nand U25952 (N_25952,N_25585,N_25744);
nor U25953 (N_25953,N_25670,N_25729);
xnor U25954 (N_25954,N_25521,N_25500);
xnor U25955 (N_25955,N_25546,N_25619);
nor U25956 (N_25956,N_25688,N_25702);
xor U25957 (N_25957,N_25614,N_25508);
and U25958 (N_25958,N_25675,N_25733);
xnor U25959 (N_25959,N_25684,N_25590);
nand U25960 (N_25960,N_25725,N_25619);
xor U25961 (N_25961,N_25713,N_25673);
or U25962 (N_25962,N_25660,N_25718);
or U25963 (N_25963,N_25714,N_25558);
xor U25964 (N_25964,N_25527,N_25536);
xor U25965 (N_25965,N_25617,N_25686);
xnor U25966 (N_25966,N_25687,N_25633);
and U25967 (N_25967,N_25586,N_25693);
and U25968 (N_25968,N_25670,N_25568);
nand U25969 (N_25969,N_25582,N_25703);
nor U25970 (N_25970,N_25725,N_25624);
or U25971 (N_25971,N_25673,N_25724);
xor U25972 (N_25972,N_25703,N_25674);
nor U25973 (N_25973,N_25633,N_25623);
nor U25974 (N_25974,N_25585,N_25550);
and U25975 (N_25975,N_25679,N_25513);
xor U25976 (N_25976,N_25721,N_25697);
or U25977 (N_25977,N_25660,N_25647);
nor U25978 (N_25978,N_25702,N_25568);
nor U25979 (N_25979,N_25730,N_25533);
nor U25980 (N_25980,N_25579,N_25630);
nand U25981 (N_25981,N_25666,N_25707);
and U25982 (N_25982,N_25523,N_25582);
and U25983 (N_25983,N_25553,N_25529);
and U25984 (N_25984,N_25713,N_25684);
xor U25985 (N_25985,N_25551,N_25682);
xor U25986 (N_25986,N_25710,N_25505);
nand U25987 (N_25987,N_25643,N_25663);
nand U25988 (N_25988,N_25654,N_25667);
nor U25989 (N_25989,N_25608,N_25706);
and U25990 (N_25990,N_25701,N_25580);
nor U25991 (N_25991,N_25587,N_25571);
nor U25992 (N_25992,N_25704,N_25731);
nand U25993 (N_25993,N_25732,N_25590);
xnor U25994 (N_25994,N_25645,N_25729);
nor U25995 (N_25995,N_25595,N_25637);
xor U25996 (N_25996,N_25605,N_25609);
nor U25997 (N_25997,N_25682,N_25703);
nor U25998 (N_25998,N_25578,N_25513);
nor U25999 (N_25999,N_25506,N_25511);
or U26000 (N_26000,N_25837,N_25883);
nor U26001 (N_26001,N_25864,N_25998);
nand U26002 (N_26002,N_25834,N_25875);
or U26003 (N_26003,N_25935,N_25750);
nor U26004 (N_26004,N_25787,N_25758);
xor U26005 (N_26005,N_25905,N_25775);
xnor U26006 (N_26006,N_25889,N_25845);
and U26007 (N_26007,N_25922,N_25958);
nand U26008 (N_26008,N_25955,N_25893);
nor U26009 (N_26009,N_25959,N_25851);
nand U26010 (N_26010,N_25916,N_25980);
xor U26011 (N_26011,N_25961,N_25838);
or U26012 (N_26012,N_25924,N_25826);
nand U26013 (N_26013,N_25840,N_25937);
or U26014 (N_26014,N_25800,N_25901);
or U26015 (N_26015,N_25978,N_25966);
or U26016 (N_26016,N_25963,N_25863);
or U26017 (N_26017,N_25928,N_25880);
and U26018 (N_26018,N_25830,N_25898);
or U26019 (N_26019,N_25825,N_25982);
and U26020 (N_26020,N_25939,N_25964);
xor U26021 (N_26021,N_25938,N_25862);
nor U26022 (N_26022,N_25979,N_25984);
or U26023 (N_26023,N_25781,N_25842);
or U26024 (N_26024,N_25848,N_25989);
nor U26025 (N_26025,N_25890,N_25786);
nand U26026 (N_26026,N_25932,N_25900);
or U26027 (N_26027,N_25917,N_25913);
nor U26028 (N_26028,N_25789,N_25983);
or U26029 (N_26029,N_25934,N_25799);
nor U26030 (N_26030,N_25812,N_25814);
nor U26031 (N_26031,N_25999,N_25952);
xor U26032 (N_26032,N_25856,N_25828);
and U26033 (N_26033,N_25841,N_25765);
or U26034 (N_26034,N_25993,N_25776);
or U26035 (N_26035,N_25754,N_25931);
or U26036 (N_26036,N_25791,N_25761);
nand U26037 (N_26037,N_25910,N_25891);
or U26038 (N_26038,N_25827,N_25899);
and U26039 (N_26039,N_25763,N_25801);
and U26040 (N_26040,N_25764,N_25804);
xnor U26041 (N_26041,N_25779,N_25947);
or U26042 (N_26042,N_25783,N_25879);
nor U26043 (N_26043,N_25884,N_25855);
nand U26044 (N_26044,N_25925,N_25756);
nand U26045 (N_26045,N_25994,N_25824);
or U26046 (N_26046,N_25906,N_25751);
nand U26047 (N_26047,N_25829,N_25792);
nand U26048 (N_26048,N_25936,N_25759);
nand U26049 (N_26049,N_25967,N_25985);
or U26050 (N_26050,N_25909,N_25768);
nand U26051 (N_26051,N_25914,N_25852);
or U26052 (N_26052,N_25844,N_25974);
and U26053 (N_26053,N_25861,N_25992);
nor U26054 (N_26054,N_25810,N_25871);
or U26055 (N_26055,N_25849,N_25923);
nand U26056 (N_26056,N_25805,N_25941);
xor U26057 (N_26057,N_25954,N_25986);
nor U26058 (N_26058,N_25946,N_25797);
or U26059 (N_26059,N_25927,N_25990);
or U26060 (N_26060,N_25881,N_25802);
and U26061 (N_26061,N_25772,N_25873);
xnor U26062 (N_26062,N_25908,N_25854);
xnor U26063 (N_26063,N_25762,N_25995);
and U26064 (N_26064,N_25874,N_25817);
nand U26065 (N_26065,N_25876,N_25766);
nor U26066 (N_26066,N_25926,N_25971);
and U26067 (N_26067,N_25780,N_25944);
xnor U26068 (N_26068,N_25798,N_25897);
or U26069 (N_26069,N_25940,N_25987);
xnor U26070 (N_26070,N_25996,N_25953);
or U26071 (N_26071,N_25843,N_25972);
nand U26072 (N_26072,N_25870,N_25853);
nand U26073 (N_26073,N_25811,N_25755);
nor U26074 (N_26074,N_25808,N_25930);
or U26075 (N_26075,N_25820,N_25823);
nand U26076 (N_26076,N_25767,N_25833);
xor U26077 (N_26077,N_25882,N_25784);
nand U26078 (N_26078,N_25950,N_25809);
nand U26079 (N_26079,N_25933,N_25872);
and U26080 (N_26080,N_25771,N_25894);
xnor U26081 (N_26081,N_25857,N_25760);
and U26082 (N_26082,N_25877,N_25774);
or U26083 (N_26083,N_25973,N_25885);
and U26084 (N_26084,N_25782,N_25806);
nor U26085 (N_26085,N_25970,N_25821);
xor U26086 (N_26086,N_25788,N_25836);
and U26087 (N_26087,N_25991,N_25822);
nor U26088 (N_26088,N_25907,N_25943);
nor U26089 (N_26089,N_25831,N_25847);
nand U26090 (N_26090,N_25865,N_25949);
xnor U26091 (N_26091,N_25929,N_25859);
and U26092 (N_26092,N_25886,N_25957);
and U26093 (N_26093,N_25868,N_25895);
nor U26094 (N_26094,N_25951,N_25918);
nor U26095 (N_26095,N_25752,N_25911);
or U26096 (N_26096,N_25896,N_25919);
and U26097 (N_26097,N_25807,N_25832);
and U26098 (N_26098,N_25818,N_25869);
and U26099 (N_26099,N_25915,N_25904);
xor U26100 (N_26100,N_25778,N_25976);
nor U26101 (N_26101,N_25793,N_25813);
xnor U26102 (N_26102,N_25977,N_25794);
xnor U26103 (N_26103,N_25815,N_25892);
nor U26104 (N_26104,N_25887,N_25968);
and U26105 (N_26105,N_25850,N_25753);
nand U26106 (N_26106,N_25816,N_25858);
or U26107 (N_26107,N_25757,N_25773);
or U26108 (N_26108,N_25988,N_25795);
nor U26109 (N_26109,N_25846,N_25902);
xnor U26110 (N_26110,N_25965,N_25921);
nor U26111 (N_26111,N_25867,N_25790);
or U26112 (N_26112,N_25956,N_25981);
nor U26113 (N_26113,N_25948,N_25796);
and U26114 (N_26114,N_25942,N_25777);
nor U26115 (N_26115,N_25962,N_25997);
nand U26116 (N_26116,N_25969,N_25819);
and U26117 (N_26117,N_25866,N_25769);
nor U26118 (N_26118,N_25960,N_25975);
nor U26119 (N_26119,N_25803,N_25903);
or U26120 (N_26120,N_25878,N_25770);
nand U26121 (N_26121,N_25888,N_25920);
or U26122 (N_26122,N_25912,N_25835);
nor U26123 (N_26123,N_25785,N_25945);
and U26124 (N_26124,N_25860,N_25839);
xor U26125 (N_26125,N_25892,N_25883);
or U26126 (N_26126,N_25800,N_25874);
or U26127 (N_26127,N_25904,N_25941);
or U26128 (N_26128,N_25807,N_25976);
nor U26129 (N_26129,N_25778,N_25781);
or U26130 (N_26130,N_25887,N_25963);
nand U26131 (N_26131,N_25970,N_25949);
nor U26132 (N_26132,N_25819,N_25959);
nand U26133 (N_26133,N_25999,N_25850);
or U26134 (N_26134,N_25870,N_25821);
nand U26135 (N_26135,N_25949,N_25827);
nor U26136 (N_26136,N_25867,N_25942);
and U26137 (N_26137,N_25867,N_25898);
nand U26138 (N_26138,N_25870,N_25963);
nor U26139 (N_26139,N_25815,N_25759);
nor U26140 (N_26140,N_25999,N_25786);
or U26141 (N_26141,N_25842,N_25899);
xor U26142 (N_26142,N_25875,N_25890);
xnor U26143 (N_26143,N_25753,N_25773);
and U26144 (N_26144,N_25791,N_25989);
and U26145 (N_26145,N_25786,N_25936);
or U26146 (N_26146,N_25778,N_25825);
nor U26147 (N_26147,N_25840,N_25842);
xnor U26148 (N_26148,N_25767,N_25816);
or U26149 (N_26149,N_25927,N_25799);
nand U26150 (N_26150,N_25886,N_25872);
xnor U26151 (N_26151,N_25775,N_25757);
or U26152 (N_26152,N_25785,N_25910);
or U26153 (N_26153,N_25815,N_25751);
or U26154 (N_26154,N_25922,N_25962);
or U26155 (N_26155,N_25939,N_25893);
and U26156 (N_26156,N_25985,N_25819);
nand U26157 (N_26157,N_25963,N_25880);
and U26158 (N_26158,N_25903,N_25974);
nand U26159 (N_26159,N_25881,N_25920);
nand U26160 (N_26160,N_25908,N_25848);
nand U26161 (N_26161,N_25924,N_25862);
nand U26162 (N_26162,N_25854,N_25987);
and U26163 (N_26163,N_25909,N_25811);
nor U26164 (N_26164,N_25808,N_25789);
or U26165 (N_26165,N_25790,N_25760);
nor U26166 (N_26166,N_25978,N_25869);
xnor U26167 (N_26167,N_25769,N_25853);
or U26168 (N_26168,N_25941,N_25912);
or U26169 (N_26169,N_25937,N_25897);
and U26170 (N_26170,N_25754,N_25869);
nand U26171 (N_26171,N_25953,N_25985);
xnor U26172 (N_26172,N_25833,N_25860);
or U26173 (N_26173,N_25767,N_25994);
nor U26174 (N_26174,N_25750,N_25911);
or U26175 (N_26175,N_25938,N_25844);
nand U26176 (N_26176,N_25890,N_25986);
and U26177 (N_26177,N_25977,N_25801);
nand U26178 (N_26178,N_25811,N_25895);
xor U26179 (N_26179,N_25844,N_25904);
nand U26180 (N_26180,N_25812,N_25811);
nor U26181 (N_26181,N_25956,N_25959);
or U26182 (N_26182,N_25799,N_25892);
nand U26183 (N_26183,N_25762,N_25849);
xnor U26184 (N_26184,N_25778,N_25828);
or U26185 (N_26185,N_25752,N_25770);
and U26186 (N_26186,N_25826,N_25901);
nor U26187 (N_26187,N_25904,N_25896);
or U26188 (N_26188,N_25774,N_25908);
xor U26189 (N_26189,N_25906,N_25774);
nor U26190 (N_26190,N_25768,N_25966);
and U26191 (N_26191,N_25942,N_25991);
nand U26192 (N_26192,N_25854,N_25912);
xnor U26193 (N_26193,N_25942,N_25812);
and U26194 (N_26194,N_25842,N_25866);
nand U26195 (N_26195,N_25908,N_25777);
xnor U26196 (N_26196,N_25924,N_25810);
nand U26197 (N_26197,N_25988,N_25766);
or U26198 (N_26198,N_25761,N_25917);
nor U26199 (N_26199,N_25895,N_25798);
and U26200 (N_26200,N_25875,N_25792);
nor U26201 (N_26201,N_25877,N_25798);
or U26202 (N_26202,N_25831,N_25947);
xnor U26203 (N_26203,N_25843,N_25847);
nand U26204 (N_26204,N_25909,N_25951);
and U26205 (N_26205,N_25887,N_25976);
nand U26206 (N_26206,N_25841,N_25993);
and U26207 (N_26207,N_25989,N_25801);
and U26208 (N_26208,N_25802,N_25974);
and U26209 (N_26209,N_25891,N_25853);
and U26210 (N_26210,N_25813,N_25945);
nand U26211 (N_26211,N_25931,N_25936);
nor U26212 (N_26212,N_25940,N_25900);
and U26213 (N_26213,N_25898,N_25848);
nand U26214 (N_26214,N_25945,N_25957);
nor U26215 (N_26215,N_25869,N_25867);
nor U26216 (N_26216,N_25757,N_25999);
and U26217 (N_26217,N_25868,N_25830);
xor U26218 (N_26218,N_25775,N_25795);
or U26219 (N_26219,N_25847,N_25868);
or U26220 (N_26220,N_25981,N_25769);
xnor U26221 (N_26221,N_25993,N_25797);
or U26222 (N_26222,N_25775,N_25927);
and U26223 (N_26223,N_25893,N_25774);
nand U26224 (N_26224,N_25866,N_25750);
nor U26225 (N_26225,N_25834,N_25902);
and U26226 (N_26226,N_25930,N_25756);
nor U26227 (N_26227,N_25781,N_25925);
nand U26228 (N_26228,N_25892,N_25877);
and U26229 (N_26229,N_25992,N_25844);
xor U26230 (N_26230,N_25762,N_25844);
or U26231 (N_26231,N_25955,N_25820);
and U26232 (N_26232,N_25869,N_25847);
and U26233 (N_26233,N_25931,N_25840);
or U26234 (N_26234,N_25885,N_25881);
xor U26235 (N_26235,N_25820,N_25785);
and U26236 (N_26236,N_25938,N_25812);
or U26237 (N_26237,N_25863,N_25920);
and U26238 (N_26238,N_25883,N_25906);
or U26239 (N_26239,N_25891,N_25788);
nor U26240 (N_26240,N_25868,N_25985);
and U26241 (N_26241,N_25934,N_25792);
or U26242 (N_26242,N_25774,N_25843);
and U26243 (N_26243,N_25904,N_25947);
nor U26244 (N_26244,N_25992,N_25795);
and U26245 (N_26245,N_25848,N_25982);
or U26246 (N_26246,N_25760,N_25807);
xnor U26247 (N_26247,N_25977,N_25855);
nor U26248 (N_26248,N_25942,N_25994);
nor U26249 (N_26249,N_25809,N_25857);
or U26250 (N_26250,N_26126,N_26116);
nand U26251 (N_26251,N_26073,N_26137);
or U26252 (N_26252,N_26081,N_26158);
xor U26253 (N_26253,N_26037,N_26071);
and U26254 (N_26254,N_26140,N_26106);
xnor U26255 (N_26255,N_26231,N_26066);
nand U26256 (N_26256,N_26136,N_26090);
xor U26257 (N_26257,N_26228,N_26076);
xor U26258 (N_26258,N_26006,N_26117);
xor U26259 (N_26259,N_26060,N_26186);
and U26260 (N_26260,N_26220,N_26139);
and U26261 (N_26261,N_26230,N_26043);
and U26262 (N_26262,N_26233,N_26063);
nor U26263 (N_26263,N_26131,N_26078);
xnor U26264 (N_26264,N_26122,N_26172);
nand U26265 (N_26265,N_26061,N_26000);
or U26266 (N_26266,N_26130,N_26207);
or U26267 (N_26267,N_26183,N_26123);
nor U26268 (N_26268,N_26248,N_26166);
xor U26269 (N_26269,N_26086,N_26149);
or U26270 (N_26270,N_26191,N_26121);
or U26271 (N_26271,N_26211,N_26144);
and U26272 (N_26272,N_26215,N_26160);
and U26273 (N_26273,N_26092,N_26185);
nor U26274 (N_26274,N_26038,N_26177);
nor U26275 (N_26275,N_26030,N_26011);
nor U26276 (N_26276,N_26194,N_26142);
nand U26277 (N_26277,N_26145,N_26197);
and U26278 (N_26278,N_26104,N_26135);
nor U26279 (N_26279,N_26196,N_26102);
nor U26280 (N_26280,N_26132,N_26067);
and U26281 (N_26281,N_26048,N_26202);
nand U26282 (N_26282,N_26157,N_26027);
xor U26283 (N_26283,N_26239,N_26069);
nand U26284 (N_26284,N_26174,N_26193);
or U26285 (N_26285,N_26124,N_26129);
and U26286 (N_26286,N_26064,N_26013);
nand U26287 (N_26287,N_26162,N_26082);
or U26288 (N_26288,N_26107,N_26068);
and U26289 (N_26289,N_26216,N_26009);
nor U26290 (N_26290,N_26008,N_26209);
nor U26291 (N_26291,N_26178,N_26190);
xnor U26292 (N_26292,N_26079,N_26055);
nor U26293 (N_26293,N_26148,N_26222);
nand U26294 (N_26294,N_26115,N_26242);
nand U26295 (N_26295,N_26152,N_26023);
nand U26296 (N_26296,N_26088,N_26112);
and U26297 (N_26297,N_26187,N_26065);
xnor U26298 (N_26298,N_26022,N_26025);
or U26299 (N_26299,N_26002,N_26192);
or U26300 (N_26300,N_26143,N_26159);
and U26301 (N_26301,N_26085,N_26175);
or U26302 (N_26302,N_26109,N_26015);
and U26303 (N_26303,N_26113,N_26164);
xnor U26304 (N_26304,N_26099,N_26094);
xnor U26305 (N_26305,N_26212,N_26206);
xnor U26306 (N_26306,N_26234,N_26053);
nor U26307 (N_26307,N_26161,N_26057);
or U26308 (N_26308,N_26077,N_26007);
nand U26309 (N_26309,N_26198,N_26236);
nand U26310 (N_26310,N_26244,N_26074);
nor U26311 (N_26311,N_26054,N_26173);
nor U26312 (N_26312,N_26133,N_26169);
nand U26313 (N_26313,N_26029,N_26203);
nor U26314 (N_26314,N_26155,N_26032);
nand U26315 (N_26315,N_26110,N_26020);
nor U26316 (N_26316,N_26018,N_26049);
or U26317 (N_26317,N_26217,N_26232);
xor U26318 (N_26318,N_26091,N_26195);
nand U26319 (N_26319,N_26201,N_26051);
nand U26320 (N_26320,N_26040,N_26039);
and U26321 (N_26321,N_26100,N_26229);
or U26322 (N_26322,N_26223,N_26056);
nand U26323 (N_26323,N_26147,N_26058);
nand U26324 (N_26324,N_26243,N_26050);
and U26325 (N_26325,N_26062,N_26014);
or U26326 (N_26326,N_26012,N_26010);
or U26327 (N_26327,N_26028,N_26189);
nand U26328 (N_26328,N_26214,N_26219);
or U26329 (N_26329,N_26045,N_26182);
or U26330 (N_26330,N_26240,N_26036);
nor U26331 (N_26331,N_26165,N_26033);
nand U26332 (N_26332,N_26095,N_26070);
nor U26333 (N_26333,N_26084,N_26105);
nor U26334 (N_26334,N_26150,N_26208);
or U26335 (N_26335,N_26151,N_26249);
xor U26336 (N_26336,N_26141,N_26019);
nor U26337 (N_26337,N_26052,N_26041);
nor U26338 (N_26338,N_26127,N_26103);
xnor U26339 (N_26339,N_26200,N_26180);
nor U26340 (N_26340,N_26238,N_26227);
nand U26341 (N_26341,N_26075,N_26237);
nor U26342 (N_26342,N_26096,N_26093);
nand U26343 (N_26343,N_26046,N_26245);
nor U26344 (N_26344,N_26026,N_26024);
and U26345 (N_26345,N_26163,N_26179);
nor U26346 (N_26346,N_26226,N_26246);
xor U26347 (N_26347,N_26235,N_26080);
nand U26348 (N_26348,N_26042,N_26120);
nor U26349 (N_26349,N_26047,N_26114);
and U26350 (N_26350,N_26221,N_26044);
xor U26351 (N_26351,N_26098,N_26146);
or U26352 (N_26352,N_26154,N_26168);
or U26353 (N_26353,N_26031,N_26205);
nand U26354 (N_26354,N_26003,N_26119);
or U26355 (N_26355,N_26097,N_26108);
or U26356 (N_26356,N_26035,N_26171);
or U26357 (N_26357,N_26224,N_26059);
nand U26358 (N_26358,N_26021,N_26089);
nor U26359 (N_26359,N_26004,N_26138);
nand U26360 (N_26360,N_26153,N_26204);
xnor U26361 (N_26361,N_26218,N_26083);
and U26362 (N_26362,N_26199,N_26213);
or U26363 (N_26363,N_26181,N_26034);
nand U26364 (N_26364,N_26167,N_26017);
and U26365 (N_26365,N_26101,N_26170);
nor U26366 (N_26366,N_26241,N_26001);
and U26367 (N_26367,N_26125,N_26184);
or U26368 (N_26368,N_26188,N_26128);
nand U26369 (N_26369,N_26225,N_26247);
nand U26370 (N_26370,N_26118,N_26176);
or U26371 (N_26371,N_26111,N_26210);
xor U26372 (N_26372,N_26072,N_26087);
xor U26373 (N_26373,N_26134,N_26156);
or U26374 (N_26374,N_26016,N_26005);
or U26375 (N_26375,N_26144,N_26115);
xor U26376 (N_26376,N_26156,N_26197);
xor U26377 (N_26377,N_26059,N_26179);
nand U26378 (N_26378,N_26065,N_26233);
nand U26379 (N_26379,N_26104,N_26064);
and U26380 (N_26380,N_26230,N_26092);
nand U26381 (N_26381,N_26193,N_26067);
nand U26382 (N_26382,N_26176,N_26181);
nand U26383 (N_26383,N_26117,N_26249);
xor U26384 (N_26384,N_26071,N_26143);
nor U26385 (N_26385,N_26244,N_26071);
nand U26386 (N_26386,N_26153,N_26214);
xnor U26387 (N_26387,N_26069,N_26214);
nand U26388 (N_26388,N_26020,N_26019);
xnor U26389 (N_26389,N_26240,N_26225);
and U26390 (N_26390,N_26109,N_26045);
xor U26391 (N_26391,N_26163,N_26120);
or U26392 (N_26392,N_26211,N_26019);
nor U26393 (N_26393,N_26165,N_26233);
and U26394 (N_26394,N_26159,N_26037);
and U26395 (N_26395,N_26219,N_26096);
and U26396 (N_26396,N_26050,N_26208);
nand U26397 (N_26397,N_26040,N_26147);
nand U26398 (N_26398,N_26143,N_26221);
nand U26399 (N_26399,N_26015,N_26224);
nor U26400 (N_26400,N_26237,N_26142);
xor U26401 (N_26401,N_26244,N_26199);
and U26402 (N_26402,N_26230,N_26205);
nor U26403 (N_26403,N_26181,N_26227);
xor U26404 (N_26404,N_26118,N_26203);
nand U26405 (N_26405,N_26077,N_26200);
and U26406 (N_26406,N_26112,N_26077);
nand U26407 (N_26407,N_26221,N_26158);
or U26408 (N_26408,N_26212,N_26027);
xnor U26409 (N_26409,N_26115,N_26222);
xor U26410 (N_26410,N_26063,N_26012);
nand U26411 (N_26411,N_26058,N_26005);
nor U26412 (N_26412,N_26213,N_26223);
or U26413 (N_26413,N_26084,N_26159);
xor U26414 (N_26414,N_26007,N_26191);
and U26415 (N_26415,N_26201,N_26203);
xor U26416 (N_26416,N_26186,N_26051);
xnor U26417 (N_26417,N_26138,N_26057);
xnor U26418 (N_26418,N_26121,N_26146);
xnor U26419 (N_26419,N_26102,N_26140);
nand U26420 (N_26420,N_26017,N_26239);
nor U26421 (N_26421,N_26016,N_26232);
xnor U26422 (N_26422,N_26204,N_26017);
nor U26423 (N_26423,N_26162,N_26165);
and U26424 (N_26424,N_26115,N_26070);
and U26425 (N_26425,N_26230,N_26028);
or U26426 (N_26426,N_26040,N_26246);
nor U26427 (N_26427,N_26170,N_26063);
and U26428 (N_26428,N_26109,N_26132);
nand U26429 (N_26429,N_26114,N_26008);
nor U26430 (N_26430,N_26141,N_26167);
or U26431 (N_26431,N_26246,N_26138);
xor U26432 (N_26432,N_26101,N_26020);
or U26433 (N_26433,N_26088,N_26226);
nor U26434 (N_26434,N_26075,N_26177);
or U26435 (N_26435,N_26101,N_26224);
or U26436 (N_26436,N_26199,N_26004);
nand U26437 (N_26437,N_26092,N_26010);
and U26438 (N_26438,N_26213,N_26112);
xor U26439 (N_26439,N_26234,N_26095);
xor U26440 (N_26440,N_26077,N_26139);
xnor U26441 (N_26441,N_26249,N_26089);
or U26442 (N_26442,N_26145,N_26170);
nand U26443 (N_26443,N_26231,N_26169);
xor U26444 (N_26444,N_26054,N_26216);
nor U26445 (N_26445,N_26092,N_26201);
and U26446 (N_26446,N_26238,N_26163);
and U26447 (N_26447,N_26165,N_26116);
xnor U26448 (N_26448,N_26219,N_26127);
nand U26449 (N_26449,N_26110,N_26024);
xor U26450 (N_26450,N_26119,N_26014);
nand U26451 (N_26451,N_26127,N_26076);
and U26452 (N_26452,N_26007,N_26067);
nor U26453 (N_26453,N_26009,N_26017);
nand U26454 (N_26454,N_26083,N_26235);
nor U26455 (N_26455,N_26060,N_26231);
xnor U26456 (N_26456,N_26234,N_26187);
or U26457 (N_26457,N_26193,N_26166);
xor U26458 (N_26458,N_26035,N_26109);
xor U26459 (N_26459,N_26134,N_26057);
and U26460 (N_26460,N_26161,N_26064);
xor U26461 (N_26461,N_26203,N_26015);
or U26462 (N_26462,N_26039,N_26227);
xor U26463 (N_26463,N_26165,N_26218);
or U26464 (N_26464,N_26154,N_26145);
or U26465 (N_26465,N_26228,N_26167);
nor U26466 (N_26466,N_26230,N_26158);
and U26467 (N_26467,N_26207,N_26020);
nand U26468 (N_26468,N_26200,N_26055);
xnor U26469 (N_26469,N_26213,N_26006);
nand U26470 (N_26470,N_26148,N_26133);
nor U26471 (N_26471,N_26110,N_26074);
xnor U26472 (N_26472,N_26027,N_26122);
nor U26473 (N_26473,N_26025,N_26037);
nor U26474 (N_26474,N_26171,N_26039);
and U26475 (N_26475,N_26062,N_26067);
or U26476 (N_26476,N_26129,N_26150);
and U26477 (N_26477,N_26093,N_26141);
or U26478 (N_26478,N_26165,N_26140);
nor U26479 (N_26479,N_26115,N_26189);
nand U26480 (N_26480,N_26243,N_26236);
and U26481 (N_26481,N_26060,N_26177);
xnor U26482 (N_26482,N_26041,N_26170);
nor U26483 (N_26483,N_26138,N_26012);
or U26484 (N_26484,N_26082,N_26077);
nand U26485 (N_26485,N_26101,N_26089);
nor U26486 (N_26486,N_26049,N_26107);
or U26487 (N_26487,N_26010,N_26221);
nand U26488 (N_26488,N_26111,N_26156);
nand U26489 (N_26489,N_26168,N_26111);
or U26490 (N_26490,N_26107,N_26011);
nand U26491 (N_26491,N_26006,N_26150);
and U26492 (N_26492,N_26207,N_26146);
nand U26493 (N_26493,N_26109,N_26115);
and U26494 (N_26494,N_26112,N_26193);
and U26495 (N_26495,N_26127,N_26218);
and U26496 (N_26496,N_26074,N_26088);
xor U26497 (N_26497,N_26224,N_26225);
and U26498 (N_26498,N_26212,N_26196);
nor U26499 (N_26499,N_26129,N_26123);
and U26500 (N_26500,N_26331,N_26472);
nand U26501 (N_26501,N_26286,N_26317);
nor U26502 (N_26502,N_26346,N_26363);
or U26503 (N_26503,N_26291,N_26493);
xnor U26504 (N_26504,N_26392,N_26250);
xor U26505 (N_26505,N_26399,N_26470);
or U26506 (N_26506,N_26297,N_26453);
nand U26507 (N_26507,N_26483,N_26336);
and U26508 (N_26508,N_26474,N_26365);
nor U26509 (N_26509,N_26339,N_26435);
and U26510 (N_26510,N_26454,N_26449);
nand U26511 (N_26511,N_26411,N_26316);
nand U26512 (N_26512,N_26420,N_26348);
or U26513 (N_26513,N_26325,N_26429);
and U26514 (N_26514,N_26359,N_26342);
or U26515 (N_26515,N_26387,N_26440);
nand U26516 (N_26516,N_26409,N_26284);
and U26517 (N_26517,N_26477,N_26289);
nor U26518 (N_26518,N_26455,N_26353);
nand U26519 (N_26519,N_26322,N_26438);
or U26520 (N_26520,N_26285,N_26329);
nand U26521 (N_26521,N_26378,N_26356);
xnor U26522 (N_26522,N_26290,N_26441);
and U26523 (N_26523,N_26256,N_26255);
xor U26524 (N_26524,N_26360,N_26313);
nand U26525 (N_26525,N_26442,N_26432);
nand U26526 (N_26526,N_26361,N_26478);
nand U26527 (N_26527,N_26371,N_26309);
and U26528 (N_26528,N_26415,N_26495);
or U26529 (N_26529,N_26480,N_26304);
xnor U26530 (N_26530,N_26287,N_26425);
xor U26531 (N_26531,N_26462,N_26376);
nand U26532 (N_26532,N_26266,N_26447);
xor U26533 (N_26533,N_26347,N_26315);
nor U26534 (N_26534,N_26251,N_26367);
or U26535 (N_26535,N_26412,N_26273);
or U26536 (N_26536,N_26271,N_26482);
xor U26537 (N_26537,N_26384,N_26253);
nand U26538 (N_26538,N_26254,N_26364);
nor U26539 (N_26539,N_26294,N_26445);
nand U26540 (N_26540,N_26321,N_26397);
or U26541 (N_26541,N_26252,N_26373);
nor U26542 (N_26542,N_26340,N_26421);
or U26543 (N_26543,N_26265,N_26401);
or U26544 (N_26544,N_26439,N_26452);
xor U26545 (N_26545,N_26333,N_26486);
nor U26546 (N_26546,N_26451,N_26269);
and U26547 (N_26547,N_26338,N_26281);
nand U26548 (N_26548,N_26385,N_26260);
or U26549 (N_26549,N_26417,N_26487);
nand U26550 (N_26550,N_26276,N_26264);
nor U26551 (N_26551,N_26407,N_26406);
nor U26552 (N_26552,N_26334,N_26295);
nand U26553 (N_26553,N_26377,N_26302);
nand U26554 (N_26554,N_26354,N_26464);
nand U26555 (N_26555,N_26418,N_26357);
xnor U26556 (N_26556,N_26259,N_26461);
nor U26557 (N_26557,N_26426,N_26390);
and U26558 (N_26558,N_26381,N_26282);
or U26559 (N_26559,N_26341,N_26436);
xnor U26560 (N_26560,N_26410,N_26328);
or U26561 (N_26561,N_26319,N_26278);
nor U26562 (N_26562,N_26383,N_26484);
nor U26563 (N_26563,N_26430,N_26386);
or U26564 (N_26564,N_26337,N_26498);
xnor U26565 (N_26565,N_26391,N_26293);
xnor U26566 (N_26566,N_26301,N_26431);
xnor U26567 (N_26567,N_26489,N_26450);
and U26568 (N_26568,N_26396,N_26463);
xor U26569 (N_26569,N_26326,N_26330);
nand U26570 (N_26570,N_26362,N_26292);
xor U26571 (N_26571,N_26497,N_26267);
or U26572 (N_26572,N_26270,N_26437);
nand U26573 (N_26573,N_26314,N_26469);
nand U26574 (N_26574,N_26475,N_26380);
and U26575 (N_26575,N_26444,N_26471);
nand U26576 (N_26576,N_26261,N_26344);
nor U26577 (N_26577,N_26283,N_26456);
xor U26578 (N_26578,N_26490,N_26466);
and U26579 (N_26579,N_26369,N_26358);
and U26580 (N_26580,N_26257,N_26300);
xnor U26581 (N_26581,N_26258,N_26379);
and U26582 (N_26582,N_26303,N_26388);
and U26583 (N_26583,N_26274,N_26479);
nor U26584 (N_26584,N_26288,N_26405);
xnor U26585 (N_26585,N_26395,N_26394);
and U26586 (N_26586,N_26398,N_26308);
or U26587 (N_26587,N_26476,N_26492);
nor U26588 (N_26588,N_26263,N_26370);
nor U26589 (N_26589,N_26446,N_26413);
and U26590 (N_26590,N_26467,N_26327);
nand U26591 (N_26591,N_26458,N_26296);
and U26592 (N_26592,N_26298,N_26488);
or U26593 (N_26593,N_26349,N_26481);
and U26594 (N_26594,N_26485,N_26355);
xnor U26595 (N_26595,N_26424,N_26311);
nand U26596 (N_26596,N_26414,N_26375);
or U26597 (N_26597,N_26368,N_26448);
nand U26598 (N_26598,N_26473,N_26468);
nor U26599 (N_26599,N_26280,N_26268);
and U26600 (N_26600,N_26345,N_26324);
nand U26601 (N_26601,N_26494,N_26419);
nor U26602 (N_26602,N_26277,N_26343);
and U26603 (N_26603,N_26307,N_26305);
nand U26604 (N_26604,N_26335,N_26496);
or U26605 (N_26605,N_26312,N_26404);
and U26606 (N_26606,N_26318,N_26306);
or U26607 (N_26607,N_26457,N_26389);
nand U26608 (N_26608,N_26427,N_26402);
nand U26609 (N_26609,N_26323,N_26272);
and U26610 (N_26610,N_26262,N_26299);
xnor U26611 (N_26611,N_26408,N_26393);
nor U26612 (N_26612,N_26416,N_26352);
nand U26613 (N_26613,N_26275,N_26433);
nor U26614 (N_26614,N_26372,N_26465);
and U26615 (N_26615,N_26374,N_26423);
or U26616 (N_26616,N_26310,N_26434);
nand U26617 (N_26617,N_26351,N_26400);
nor U26618 (N_26618,N_26403,N_26422);
and U26619 (N_26619,N_26332,N_26459);
and U26620 (N_26620,N_26460,N_26491);
nor U26621 (N_26621,N_26279,N_26499);
nor U26622 (N_26622,N_26366,N_26382);
or U26623 (N_26623,N_26443,N_26350);
nand U26624 (N_26624,N_26320,N_26428);
and U26625 (N_26625,N_26479,N_26337);
xor U26626 (N_26626,N_26325,N_26400);
nand U26627 (N_26627,N_26374,N_26416);
nand U26628 (N_26628,N_26455,N_26395);
and U26629 (N_26629,N_26387,N_26464);
or U26630 (N_26630,N_26265,N_26264);
nor U26631 (N_26631,N_26294,N_26311);
and U26632 (N_26632,N_26479,N_26324);
nand U26633 (N_26633,N_26339,N_26365);
xor U26634 (N_26634,N_26425,N_26276);
nand U26635 (N_26635,N_26369,N_26495);
nand U26636 (N_26636,N_26257,N_26425);
and U26637 (N_26637,N_26474,N_26482);
or U26638 (N_26638,N_26287,N_26310);
nand U26639 (N_26639,N_26412,N_26387);
and U26640 (N_26640,N_26402,N_26285);
nor U26641 (N_26641,N_26288,N_26362);
nor U26642 (N_26642,N_26373,N_26332);
or U26643 (N_26643,N_26289,N_26427);
nor U26644 (N_26644,N_26426,N_26499);
nand U26645 (N_26645,N_26468,N_26308);
and U26646 (N_26646,N_26293,N_26319);
xnor U26647 (N_26647,N_26396,N_26325);
xor U26648 (N_26648,N_26347,N_26364);
nor U26649 (N_26649,N_26257,N_26361);
and U26650 (N_26650,N_26263,N_26319);
and U26651 (N_26651,N_26462,N_26425);
xor U26652 (N_26652,N_26452,N_26358);
nor U26653 (N_26653,N_26385,N_26386);
xor U26654 (N_26654,N_26301,N_26375);
or U26655 (N_26655,N_26261,N_26378);
xor U26656 (N_26656,N_26355,N_26412);
or U26657 (N_26657,N_26437,N_26352);
nand U26658 (N_26658,N_26279,N_26371);
xnor U26659 (N_26659,N_26343,N_26424);
nor U26660 (N_26660,N_26259,N_26498);
or U26661 (N_26661,N_26457,N_26497);
or U26662 (N_26662,N_26324,N_26442);
and U26663 (N_26663,N_26265,N_26313);
nor U26664 (N_26664,N_26440,N_26317);
nor U26665 (N_26665,N_26307,N_26334);
or U26666 (N_26666,N_26434,N_26420);
nand U26667 (N_26667,N_26420,N_26334);
or U26668 (N_26668,N_26340,N_26454);
and U26669 (N_26669,N_26396,N_26400);
xor U26670 (N_26670,N_26354,N_26301);
or U26671 (N_26671,N_26293,N_26347);
and U26672 (N_26672,N_26465,N_26384);
nor U26673 (N_26673,N_26331,N_26357);
or U26674 (N_26674,N_26339,N_26473);
or U26675 (N_26675,N_26374,N_26262);
or U26676 (N_26676,N_26363,N_26325);
nand U26677 (N_26677,N_26452,N_26356);
nor U26678 (N_26678,N_26494,N_26283);
nand U26679 (N_26679,N_26336,N_26426);
nor U26680 (N_26680,N_26438,N_26497);
and U26681 (N_26681,N_26436,N_26477);
or U26682 (N_26682,N_26367,N_26352);
xnor U26683 (N_26683,N_26326,N_26443);
or U26684 (N_26684,N_26457,N_26436);
and U26685 (N_26685,N_26423,N_26464);
xor U26686 (N_26686,N_26308,N_26263);
xor U26687 (N_26687,N_26375,N_26464);
xor U26688 (N_26688,N_26290,N_26323);
nand U26689 (N_26689,N_26487,N_26284);
nor U26690 (N_26690,N_26357,N_26425);
or U26691 (N_26691,N_26300,N_26477);
nor U26692 (N_26692,N_26498,N_26494);
nand U26693 (N_26693,N_26295,N_26403);
nor U26694 (N_26694,N_26251,N_26486);
and U26695 (N_26695,N_26281,N_26326);
or U26696 (N_26696,N_26382,N_26334);
and U26697 (N_26697,N_26272,N_26314);
nand U26698 (N_26698,N_26478,N_26320);
nor U26699 (N_26699,N_26352,N_26294);
and U26700 (N_26700,N_26470,N_26476);
and U26701 (N_26701,N_26470,N_26461);
nor U26702 (N_26702,N_26495,N_26496);
and U26703 (N_26703,N_26319,N_26355);
nand U26704 (N_26704,N_26383,N_26268);
xnor U26705 (N_26705,N_26329,N_26347);
nor U26706 (N_26706,N_26443,N_26401);
or U26707 (N_26707,N_26426,N_26471);
nor U26708 (N_26708,N_26387,N_26471);
or U26709 (N_26709,N_26317,N_26355);
and U26710 (N_26710,N_26347,N_26264);
xnor U26711 (N_26711,N_26264,N_26457);
nor U26712 (N_26712,N_26301,N_26309);
nor U26713 (N_26713,N_26309,N_26479);
nor U26714 (N_26714,N_26460,N_26462);
or U26715 (N_26715,N_26466,N_26478);
nor U26716 (N_26716,N_26417,N_26319);
nor U26717 (N_26717,N_26294,N_26350);
nor U26718 (N_26718,N_26333,N_26384);
and U26719 (N_26719,N_26308,N_26342);
nand U26720 (N_26720,N_26271,N_26287);
or U26721 (N_26721,N_26327,N_26312);
xor U26722 (N_26722,N_26379,N_26358);
nand U26723 (N_26723,N_26394,N_26397);
nand U26724 (N_26724,N_26286,N_26453);
or U26725 (N_26725,N_26276,N_26300);
or U26726 (N_26726,N_26397,N_26468);
or U26727 (N_26727,N_26491,N_26263);
and U26728 (N_26728,N_26496,N_26398);
nor U26729 (N_26729,N_26414,N_26351);
or U26730 (N_26730,N_26496,N_26415);
nand U26731 (N_26731,N_26326,N_26459);
and U26732 (N_26732,N_26476,N_26325);
nor U26733 (N_26733,N_26250,N_26270);
or U26734 (N_26734,N_26329,N_26499);
and U26735 (N_26735,N_26311,N_26261);
nor U26736 (N_26736,N_26420,N_26357);
nand U26737 (N_26737,N_26472,N_26250);
and U26738 (N_26738,N_26252,N_26485);
or U26739 (N_26739,N_26435,N_26436);
nor U26740 (N_26740,N_26350,N_26357);
and U26741 (N_26741,N_26496,N_26372);
or U26742 (N_26742,N_26333,N_26412);
or U26743 (N_26743,N_26290,N_26309);
xor U26744 (N_26744,N_26380,N_26337);
xor U26745 (N_26745,N_26358,N_26340);
and U26746 (N_26746,N_26258,N_26431);
xor U26747 (N_26747,N_26326,N_26482);
nand U26748 (N_26748,N_26297,N_26444);
xnor U26749 (N_26749,N_26307,N_26379);
xor U26750 (N_26750,N_26622,N_26526);
nor U26751 (N_26751,N_26522,N_26555);
xnor U26752 (N_26752,N_26676,N_26675);
xnor U26753 (N_26753,N_26544,N_26645);
nor U26754 (N_26754,N_26562,N_26697);
xor U26755 (N_26755,N_26701,N_26742);
nand U26756 (N_26756,N_26573,N_26712);
or U26757 (N_26757,N_26745,N_26729);
nand U26758 (N_26758,N_26515,N_26629);
or U26759 (N_26759,N_26572,N_26633);
or U26760 (N_26760,N_26710,N_26648);
or U26761 (N_26761,N_26631,N_26530);
and U26762 (N_26762,N_26501,N_26593);
and U26763 (N_26763,N_26595,N_26692);
nand U26764 (N_26764,N_26743,N_26596);
nand U26765 (N_26765,N_26549,N_26610);
nand U26766 (N_26766,N_26619,N_26558);
and U26767 (N_26767,N_26539,N_26550);
nor U26768 (N_26768,N_26680,N_26685);
xnor U26769 (N_26769,N_26519,N_26630);
nand U26770 (N_26770,N_26649,N_26514);
nand U26771 (N_26771,N_26568,N_26646);
nor U26772 (N_26772,N_26554,N_26711);
and U26773 (N_26773,N_26528,N_26669);
nor U26774 (N_26774,N_26571,N_26563);
or U26775 (N_26775,N_26635,N_26664);
nand U26776 (N_26776,N_26683,N_26588);
and U26777 (N_26777,N_26704,N_26557);
and U26778 (N_26778,N_26658,N_26500);
or U26779 (N_26779,N_26678,N_26654);
xnor U26780 (N_26780,N_26735,N_26628);
nand U26781 (N_26781,N_26505,N_26607);
or U26782 (N_26782,N_26691,N_26731);
nor U26783 (N_26783,N_26749,N_26569);
or U26784 (N_26784,N_26653,N_26627);
xor U26785 (N_26785,N_26724,N_26707);
and U26786 (N_26786,N_26527,N_26617);
xnor U26787 (N_26787,N_26699,N_26686);
and U26788 (N_26788,N_26739,N_26723);
nor U26789 (N_26789,N_26728,N_26620);
nor U26790 (N_26790,N_26529,N_26706);
nand U26791 (N_26791,N_26661,N_26537);
nand U26792 (N_26792,N_26581,N_26662);
and U26793 (N_26793,N_26727,N_26615);
xor U26794 (N_26794,N_26637,N_26643);
xnor U26795 (N_26795,N_26541,N_26740);
nand U26796 (N_26796,N_26632,N_26726);
nor U26797 (N_26797,N_26682,N_26533);
xnor U26798 (N_26798,N_26679,N_26674);
nor U26799 (N_26799,N_26580,N_26538);
nand U26800 (N_26800,N_26564,N_26652);
nor U26801 (N_26801,N_26552,N_26657);
xor U26802 (N_26802,N_26513,N_26709);
nor U26803 (N_26803,N_26732,N_26576);
and U26804 (N_26804,N_26561,N_26520);
and U26805 (N_26805,N_26639,N_26598);
or U26806 (N_26806,N_26601,N_26696);
and U26807 (N_26807,N_26618,N_26695);
and U26808 (N_26808,N_26672,N_26665);
xnor U26809 (N_26809,N_26604,N_26603);
and U26810 (N_26810,N_26502,N_26606);
nor U26811 (N_26811,N_26730,N_26725);
and U26812 (N_26812,N_26738,N_26681);
and U26813 (N_26813,N_26720,N_26690);
or U26814 (N_26814,N_26602,N_26504);
or U26815 (N_26815,N_26574,N_26640);
and U26816 (N_26816,N_26542,N_26694);
nor U26817 (N_26817,N_26650,N_26600);
nor U26818 (N_26818,N_26715,N_26660);
nand U26819 (N_26819,N_26744,N_26616);
nor U26820 (N_26820,N_26584,N_26689);
xnor U26821 (N_26821,N_26659,N_26510);
nor U26822 (N_26822,N_26612,N_26677);
and U26823 (N_26823,N_26688,N_26516);
nand U26824 (N_26824,N_26547,N_26719);
xor U26825 (N_26825,N_26636,N_26548);
xor U26826 (N_26826,N_26546,N_26587);
and U26827 (N_26827,N_26668,N_26585);
nor U26828 (N_26828,N_26578,N_26582);
and U26829 (N_26829,N_26508,N_26590);
nand U26830 (N_26830,N_26718,N_26623);
and U26831 (N_26831,N_26666,N_26734);
or U26832 (N_26832,N_26553,N_26642);
xnor U26833 (N_26833,N_26722,N_26663);
or U26834 (N_26834,N_26577,N_26673);
nand U26835 (N_26835,N_26518,N_26524);
nand U26836 (N_26836,N_26703,N_26586);
or U26837 (N_26837,N_26608,N_26693);
nand U26838 (N_26838,N_26667,N_26656);
nand U26839 (N_26839,N_26507,N_26746);
and U26840 (N_26840,N_26736,N_26716);
nor U26841 (N_26841,N_26594,N_26567);
nor U26842 (N_26842,N_26540,N_26517);
nor U26843 (N_26843,N_26698,N_26741);
nor U26844 (N_26844,N_26647,N_26713);
and U26845 (N_26845,N_26613,N_26511);
xnor U26846 (N_26846,N_26575,N_26624);
and U26847 (N_26847,N_26525,N_26535);
nor U26848 (N_26848,N_26733,N_26621);
nor U26849 (N_26849,N_26625,N_26545);
and U26850 (N_26850,N_26609,N_26700);
xnor U26851 (N_26851,N_26626,N_26521);
xor U26852 (N_26852,N_26714,N_26737);
xor U26853 (N_26853,N_26560,N_26684);
and U26854 (N_26854,N_26747,N_26597);
xor U26855 (N_26855,N_26532,N_26579);
and U26856 (N_26856,N_26565,N_26512);
nand U26857 (N_26857,N_26705,N_26570);
nor U26858 (N_26858,N_26592,N_26634);
and U26859 (N_26859,N_26534,N_26671);
nand U26860 (N_26860,N_26536,N_26566);
xor U26861 (N_26861,N_26748,N_26644);
nor U26862 (N_26862,N_26641,N_26531);
nor U26863 (N_26863,N_26614,N_26611);
nand U26864 (N_26864,N_26599,N_26605);
xnor U26865 (N_26865,N_26589,N_26503);
nor U26866 (N_26866,N_26551,N_26702);
xnor U26867 (N_26867,N_26583,N_26687);
nor U26868 (N_26868,N_26523,N_26543);
nor U26869 (N_26869,N_26708,N_26591);
nand U26870 (N_26870,N_26506,N_26717);
and U26871 (N_26871,N_26651,N_26509);
nor U26872 (N_26872,N_26559,N_26556);
or U26873 (N_26873,N_26655,N_26638);
and U26874 (N_26874,N_26670,N_26721);
and U26875 (N_26875,N_26507,N_26528);
and U26876 (N_26876,N_26544,N_26667);
nand U26877 (N_26877,N_26726,N_26682);
nand U26878 (N_26878,N_26722,N_26649);
nand U26879 (N_26879,N_26647,N_26610);
and U26880 (N_26880,N_26633,N_26529);
and U26881 (N_26881,N_26660,N_26684);
nor U26882 (N_26882,N_26541,N_26688);
nand U26883 (N_26883,N_26702,N_26710);
nor U26884 (N_26884,N_26738,N_26587);
or U26885 (N_26885,N_26654,N_26538);
and U26886 (N_26886,N_26541,N_26731);
or U26887 (N_26887,N_26500,N_26547);
and U26888 (N_26888,N_26578,N_26600);
nor U26889 (N_26889,N_26612,N_26562);
nor U26890 (N_26890,N_26620,N_26554);
xor U26891 (N_26891,N_26702,N_26743);
and U26892 (N_26892,N_26572,N_26747);
nor U26893 (N_26893,N_26654,N_26748);
nand U26894 (N_26894,N_26547,N_26531);
nor U26895 (N_26895,N_26591,N_26715);
nor U26896 (N_26896,N_26666,N_26531);
or U26897 (N_26897,N_26734,N_26506);
nor U26898 (N_26898,N_26625,N_26610);
or U26899 (N_26899,N_26600,N_26726);
or U26900 (N_26900,N_26548,N_26722);
xnor U26901 (N_26901,N_26522,N_26625);
and U26902 (N_26902,N_26559,N_26583);
and U26903 (N_26903,N_26713,N_26537);
and U26904 (N_26904,N_26560,N_26727);
and U26905 (N_26905,N_26681,N_26585);
nor U26906 (N_26906,N_26542,N_26635);
xor U26907 (N_26907,N_26513,N_26722);
xnor U26908 (N_26908,N_26626,N_26501);
xor U26909 (N_26909,N_26676,N_26722);
nor U26910 (N_26910,N_26644,N_26742);
and U26911 (N_26911,N_26564,N_26724);
or U26912 (N_26912,N_26640,N_26538);
xnor U26913 (N_26913,N_26649,N_26690);
or U26914 (N_26914,N_26640,N_26680);
or U26915 (N_26915,N_26683,N_26678);
nand U26916 (N_26916,N_26739,N_26662);
xor U26917 (N_26917,N_26505,N_26584);
or U26918 (N_26918,N_26665,N_26609);
nand U26919 (N_26919,N_26740,N_26640);
xnor U26920 (N_26920,N_26635,N_26574);
nor U26921 (N_26921,N_26507,N_26533);
nor U26922 (N_26922,N_26680,N_26669);
or U26923 (N_26923,N_26672,N_26664);
or U26924 (N_26924,N_26568,N_26694);
nand U26925 (N_26925,N_26749,N_26627);
xnor U26926 (N_26926,N_26718,N_26568);
nor U26927 (N_26927,N_26502,N_26614);
xnor U26928 (N_26928,N_26666,N_26573);
xnor U26929 (N_26929,N_26581,N_26585);
nand U26930 (N_26930,N_26583,N_26712);
and U26931 (N_26931,N_26691,N_26664);
or U26932 (N_26932,N_26550,N_26587);
or U26933 (N_26933,N_26550,N_26712);
nor U26934 (N_26934,N_26516,N_26617);
xnor U26935 (N_26935,N_26624,N_26513);
or U26936 (N_26936,N_26531,N_26635);
or U26937 (N_26937,N_26711,N_26572);
or U26938 (N_26938,N_26665,N_26685);
nand U26939 (N_26939,N_26586,N_26623);
and U26940 (N_26940,N_26644,N_26578);
nand U26941 (N_26941,N_26630,N_26651);
xor U26942 (N_26942,N_26546,N_26725);
and U26943 (N_26943,N_26607,N_26733);
nand U26944 (N_26944,N_26625,N_26702);
nand U26945 (N_26945,N_26737,N_26580);
nand U26946 (N_26946,N_26745,N_26682);
or U26947 (N_26947,N_26524,N_26691);
and U26948 (N_26948,N_26602,N_26624);
or U26949 (N_26949,N_26563,N_26650);
xnor U26950 (N_26950,N_26572,N_26581);
nor U26951 (N_26951,N_26729,N_26504);
and U26952 (N_26952,N_26676,N_26617);
nor U26953 (N_26953,N_26723,N_26575);
nor U26954 (N_26954,N_26639,N_26679);
and U26955 (N_26955,N_26690,N_26702);
nor U26956 (N_26956,N_26690,N_26709);
or U26957 (N_26957,N_26636,N_26723);
xnor U26958 (N_26958,N_26563,N_26507);
xor U26959 (N_26959,N_26574,N_26667);
nand U26960 (N_26960,N_26723,N_26736);
and U26961 (N_26961,N_26609,N_26538);
nand U26962 (N_26962,N_26706,N_26704);
or U26963 (N_26963,N_26723,N_26605);
nor U26964 (N_26964,N_26703,N_26696);
or U26965 (N_26965,N_26645,N_26708);
or U26966 (N_26966,N_26583,N_26576);
nor U26967 (N_26967,N_26617,N_26618);
or U26968 (N_26968,N_26631,N_26533);
nor U26969 (N_26969,N_26712,N_26619);
nand U26970 (N_26970,N_26542,N_26699);
and U26971 (N_26971,N_26708,N_26588);
nand U26972 (N_26972,N_26680,N_26517);
and U26973 (N_26973,N_26587,N_26655);
or U26974 (N_26974,N_26570,N_26502);
nand U26975 (N_26975,N_26522,N_26505);
or U26976 (N_26976,N_26639,N_26569);
and U26977 (N_26977,N_26590,N_26643);
nor U26978 (N_26978,N_26553,N_26500);
or U26979 (N_26979,N_26689,N_26736);
nor U26980 (N_26980,N_26524,N_26603);
xor U26981 (N_26981,N_26587,N_26507);
nor U26982 (N_26982,N_26580,N_26729);
nor U26983 (N_26983,N_26637,N_26556);
or U26984 (N_26984,N_26609,N_26559);
xnor U26985 (N_26985,N_26505,N_26635);
xnor U26986 (N_26986,N_26667,N_26724);
or U26987 (N_26987,N_26697,N_26722);
xnor U26988 (N_26988,N_26502,N_26666);
nand U26989 (N_26989,N_26694,N_26579);
or U26990 (N_26990,N_26738,N_26613);
nor U26991 (N_26991,N_26609,N_26561);
xor U26992 (N_26992,N_26553,N_26725);
xor U26993 (N_26993,N_26515,N_26552);
xor U26994 (N_26994,N_26582,N_26627);
nor U26995 (N_26995,N_26594,N_26677);
or U26996 (N_26996,N_26568,N_26613);
nor U26997 (N_26997,N_26535,N_26627);
xnor U26998 (N_26998,N_26527,N_26593);
and U26999 (N_26999,N_26749,N_26582);
and U27000 (N_27000,N_26918,N_26907);
or U27001 (N_27001,N_26917,N_26922);
or U27002 (N_27002,N_26937,N_26798);
xnor U27003 (N_27003,N_26867,N_26945);
xnor U27004 (N_27004,N_26924,N_26964);
nor U27005 (N_27005,N_26985,N_26794);
or U27006 (N_27006,N_26797,N_26815);
nand U27007 (N_27007,N_26994,N_26851);
or U27008 (N_27008,N_26951,N_26900);
nor U27009 (N_27009,N_26824,N_26774);
xnor U27010 (N_27010,N_26857,N_26939);
nor U27011 (N_27011,N_26829,N_26868);
xor U27012 (N_27012,N_26811,N_26973);
nor U27013 (N_27013,N_26760,N_26799);
and U27014 (N_27014,N_26997,N_26856);
xor U27015 (N_27015,N_26795,N_26986);
nand U27016 (N_27016,N_26974,N_26770);
and U27017 (N_27017,N_26814,N_26825);
nor U27018 (N_27018,N_26771,N_26959);
or U27019 (N_27019,N_26948,N_26883);
xor U27020 (N_27020,N_26834,N_26887);
and U27021 (N_27021,N_26775,N_26776);
nor U27022 (N_27022,N_26992,N_26884);
nor U27023 (N_27023,N_26822,N_26835);
or U27024 (N_27024,N_26808,N_26925);
and U27025 (N_27025,N_26999,N_26763);
nor U27026 (N_27026,N_26979,N_26967);
nor U27027 (N_27027,N_26810,N_26832);
nand U27028 (N_27028,N_26898,N_26827);
nor U27029 (N_27029,N_26759,N_26903);
xnor U27030 (N_27030,N_26843,N_26919);
nand U27031 (N_27031,N_26773,N_26845);
xnor U27032 (N_27032,N_26984,N_26993);
or U27033 (N_27033,N_26929,N_26860);
or U27034 (N_27034,N_26879,N_26969);
nor U27035 (N_27035,N_26863,N_26846);
nor U27036 (N_27036,N_26899,N_26788);
nand U27037 (N_27037,N_26869,N_26823);
or U27038 (N_27038,N_26840,N_26910);
nand U27039 (N_27039,N_26765,N_26809);
and U27040 (N_27040,N_26978,N_26980);
and U27041 (N_27041,N_26752,N_26976);
or U27042 (N_27042,N_26878,N_26826);
xnor U27043 (N_27043,N_26895,N_26987);
nand U27044 (N_27044,N_26871,N_26833);
or U27045 (N_27045,N_26839,N_26762);
nor U27046 (N_27046,N_26963,N_26906);
or U27047 (N_27047,N_26880,N_26831);
nand U27048 (N_27048,N_26806,N_26933);
nand U27049 (N_27049,N_26865,N_26782);
nand U27050 (N_27050,N_26926,N_26761);
nor U27051 (N_27051,N_26975,N_26920);
nand U27052 (N_27052,N_26838,N_26891);
nor U27053 (N_27053,N_26781,N_26989);
and U27054 (N_27054,N_26772,N_26946);
nand U27055 (N_27055,N_26940,N_26909);
nand U27056 (N_27056,N_26934,N_26807);
nor U27057 (N_27057,N_26755,N_26875);
nand U27058 (N_27058,N_26777,N_26952);
and U27059 (N_27059,N_26971,N_26753);
xor U27060 (N_27060,N_26897,N_26791);
xor U27061 (N_27061,N_26876,N_26914);
and U27062 (N_27062,N_26894,N_26961);
or U27063 (N_27063,N_26977,N_26873);
nand U27064 (N_27064,N_26881,N_26938);
and U27065 (N_27065,N_26958,N_26836);
xnor U27066 (N_27066,N_26830,N_26996);
nand U27067 (N_27067,N_26872,N_26941);
or U27068 (N_27068,N_26988,N_26818);
and U27069 (N_27069,N_26803,N_26982);
xnor U27070 (N_27070,N_26885,N_26923);
or U27071 (N_27071,N_26842,N_26882);
nand U27072 (N_27072,N_26904,N_26844);
or U27073 (N_27073,N_26886,N_26805);
and U27074 (N_27074,N_26936,N_26849);
nand U27075 (N_27075,N_26750,N_26852);
nor U27076 (N_27076,N_26931,N_26796);
and U27077 (N_27077,N_26890,N_26790);
and U27078 (N_27078,N_26751,N_26889);
and U27079 (N_27079,N_26991,N_26932);
nand U27080 (N_27080,N_26780,N_26870);
nor U27081 (N_27081,N_26841,N_26850);
xor U27082 (N_27082,N_26928,N_26949);
nand U27083 (N_27083,N_26921,N_26864);
nor U27084 (N_27084,N_26764,N_26957);
nor U27085 (N_27085,N_26802,N_26966);
xnor U27086 (N_27086,N_26858,N_26828);
nand U27087 (N_27087,N_26854,N_26947);
or U27088 (N_27088,N_26960,N_26968);
and U27089 (N_27089,N_26908,N_26816);
or U27090 (N_27090,N_26962,N_26956);
or U27091 (N_27091,N_26965,N_26848);
nor U27092 (N_27092,N_26754,N_26787);
or U27093 (N_27093,N_26896,N_26855);
nand U27094 (N_27094,N_26756,N_26970);
nor U27095 (N_27095,N_26778,N_26915);
and U27096 (N_27096,N_26758,N_26786);
xnor U27097 (N_27097,N_26998,N_26813);
nand U27098 (N_27098,N_26766,N_26866);
and U27099 (N_27099,N_26950,N_26804);
and U27100 (N_27100,N_26821,N_26767);
nor U27101 (N_27101,N_26943,N_26955);
or U27102 (N_27102,N_26847,N_26944);
or U27103 (N_27103,N_26792,N_26893);
and U27104 (N_27104,N_26981,N_26859);
nor U27105 (N_27105,N_26877,N_26935);
nand U27106 (N_27106,N_26912,N_26853);
nor U27107 (N_27107,N_26793,N_26819);
or U27108 (N_27108,N_26954,N_26862);
nand U27109 (N_27109,N_26905,N_26911);
and U27110 (N_27110,N_26837,N_26785);
and U27111 (N_27111,N_26990,N_26801);
nand U27112 (N_27112,N_26892,N_26784);
nand U27113 (N_27113,N_26812,N_26874);
and U27114 (N_27114,N_26768,N_26972);
or U27115 (N_27115,N_26983,N_26888);
and U27116 (N_27116,N_26817,N_26789);
nor U27117 (N_27117,N_26927,N_26953);
nor U27118 (N_27118,N_26769,N_26995);
nor U27119 (N_27119,N_26916,N_26757);
or U27120 (N_27120,N_26930,N_26902);
nor U27121 (N_27121,N_26783,N_26820);
nor U27122 (N_27122,N_26861,N_26901);
or U27123 (N_27123,N_26800,N_26942);
nor U27124 (N_27124,N_26913,N_26779);
nor U27125 (N_27125,N_26879,N_26984);
nand U27126 (N_27126,N_26819,N_26925);
xnor U27127 (N_27127,N_26830,N_26977);
xnor U27128 (N_27128,N_26956,N_26961);
nand U27129 (N_27129,N_26841,N_26826);
nor U27130 (N_27130,N_26968,N_26995);
nor U27131 (N_27131,N_26935,N_26956);
or U27132 (N_27132,N_26986,N_26848);
and U27133 (N_27133,N_26823,N_26888);
nor U27134 (N_27134,N_26785,N_26757);
xor U27135 (N_27135,N_26897,N_26846);
or U27136 (N_27136,N_26834,N_26842);
xnor U27137 (N_27137,N_26974,N_26900);
and U27138 (N_27138,N_26975,N_26894);
nand U27139 (N_27139,N_26875,N_26966);
or U27140 (N_27140,N_26964,N_26906);
nand U27141 (N_27141,N_26824,N_26860);
xnor U27142 (N_27142,N_26965,N_26881);
and U27143 (N_27143,N_26846,N_26921);
xnor U27144 (N_27144,N_26838,N_26790);
nand U27145 (N_27145,N_26762,N_26894);
nor U27146 (N_27146,N_26894,N_26956);
or U27147 (N_27147,N_26751,N_26855);
nor U27148 (N_27148,N_26774,N_26950);
xnor U27149 (N_27149,N_26770,N_26825);
nor U27150 (N_27150,N_26947,N_26967);
xnor U27151 (N_27151,N_26868,N_26792);
xor U27152 (N_27152,N_26968,N_26869);
nand U27153 (N_27153,N_26811,N_26976);
nor U27154 (N_27154,N_26782,N_26947);
or U27155 (N_27155,N_26815,N_26983);
nand U27156 (N_27156,N_26854,N_26802);
and U27157 (N_27157,N_26776,N_26781);
xnor U27158 (N_27158,N_26997,N_26818);
xor U27159 (N_27159,N_26800,N_26825);
and U27160 (N_27160,N_26894,N_26939);
nor U27161 (N_27161,N_26800,N_26999);
or U27162 (N_27162,N_26750,N_26980);
xor U27163 (N_27163,N_26868,N_26994);
nor U27164 (N_27164,N_26877,N_26810);
or U27165 (N_27165,N_26783,N_26793);
nor U27166 (N_27166,N_26818,N_26764);
and U27167 (N_27167,N_26756,N_26780);
nor U27168 (N_27168,N_26805,N_26787);
nand U27169 (N_27169,N_26795,N_26929);
and U27170 (N_27170,N_26948,N_26873);
nand U27171 (N_27171,N_26830,N_26760);
or U27172 (N_27172,N_26949,N_26947);
xor U27173 (N_27173,N_26792,N_26789);
or U27174 (N_27174,N_26882,N_26823);
nand U27175 (N_27175,N_26852,N_26999);
xor U27176 (N_27176,N_26998,N_26866);
and U27177 (N_27177,N_26894,N_26998);
and U27178 (N_27178,N_26815,N_26867);
and U27179 (N_27179,N_26966,N_26832);
nor U27180 (N_27180,N_26916,N_26974);
or U27181 (N_27181,N_26904,N_26849);
and U27182 (N_27182,N_26963,N_26994);
nor U27183 (N_27183,N_26836,N_26912);
xnor U27184 (N_27184,N_26919,N_26994);
nor U27185 (N_27185,N_26999,N_26838);
xor U27186 (N_27186,N_26842,N_26867);
or U27187 (N_27187,N_26862,N_26754);
and U27188 (N_27188,N_26917,N_26774);
and U27189 (N_27189,N_26989,N_26839);
or U27190 (N_27190,N_26897,N_26908);
nand U27191 (N_27191,N_26802,N_26998);
nand U27192 (N_27192,N_26899,N_26936);
nand U27193 (N_27193,N_26924,N_26911);
nand U27194 (N_27194,N_26816,N_26751);
nand U27195 (N_27195,N_26938,N_26809);
or U27196 (N_27196,N_26757,N_26946);
nor U27197 (N_27197,N_26831,N_26762);
nor U27198 (N_27198,N_26820,N_26854);
or U27199 (N_27199,N_26903,N_26845);
nand U27200 (N_27200,N_26862,N_26762);
or U27201 (N_27201,N_26761,N_26870);
and U27202 (N_27202,N_26992,N_26797);
or U27203 (N_27203,N_26770,N_26978);
or U27204 (N_27204,N_26761,N_26911);
nor U27205 (N_27205,N_26818,N_26883);
or U27206 (N_27206,N_26919,N_26936);
xor U27207 (N_27207,N_26809,N_26859);
nor U27208 (N_27208,N_26825,N_26955);
or U27209 (N_27209,N_26933,N_26894);
nand U27210 (N_27210,N_26824,N_26983);
or U27211 (N_27211,N_26775,N_26913);
nor U27212 (N_27212,N_26926,N_26778);
or U27213 (N_27213,N_26894,N_26891);
and U27214 (N_27214,N_26946,N_26790);
and U27215 (N_27215,N_26808,N_26806);
or U27216 (N_27216,N_26921,N_26973);
nand U27217 (N_27217,N_26842,N_26778);
xor U27218 (N_27218,N_26802,N_26954);
and U27219 (N_27219,N_26824,N_26922);
and U27220 (N_27220,N_26947,N_26785);
nor U27221 (N_27221,N_26794,N_26809);
nand U27222 (N_27222,N_26834,N_26809);
and U27223 (N_27223,N_26909,N_26901);
or U27224 (N_27224,N_26808,N_26910);
nor U27225 (N_27225,N_26992,N_26979);
or U27226 (N_27226,N_26835,N_26979);
nand U27227 (N_27227,N_26961,N_26759);
nor U27228 (N_27228,N_26782,N_26881);
nor U27229 (N_27229,N_26761,N_26810);
xor U27230 (N_27230,N_26803,N_26826);
or U27231 (N_27231,N_26750,N_26910);
or U27232 (N_27232,N_26948,N_26930);
nand U27233 (N_27233,N_26989,N_26832);
or U27234 (N_27234,N_26780,N_26820);
nor U27235 (N_27235,N_26933,N_26905);
nand U27236 (N_27236,N_26807,N_26760);
and U27237 (N_27237,N_26848,N_26798);
and U27238 (N_27238,N_26851,N_26919);
or U27239 (N_27239,N_26750,N_26929);
or U27240 (N_27240,N_26763,N_26945);
xor U27241 (N_27241,N_26868,N_26914);
nor U27242 (N_27242,N_26981,N_26995);
nor U27243 (N_27243,N_26979,N_26851);
and U27244 (N_27244,N_26808,N_26878);
nand U27245 (N_27245,N_26969,N_26979);
nand U27246 (N_27246,N_26963,N_26957);
and U27247 (N_27247,N_26801,N_26854);
and U27248 (N_27248,N_26896,N_26890);
nor U27249 (N_27249,N_26931,N_26885);
nor U27250 (N_27250,N_27006,N_27075);
or U27251 (N_27251,N_27168,N_27091);
nor U27252 (N_27252,N_27154,N_27137);
or U27253 (N_27253,N_27041,N_27231);
nand U27254 (N_27254,N_27080,N_27119);
nor U27255 (N_27255,N_27032,N_27082);
nor U27256 (N_27256,N_27205,N_27000);
or U27257 (N_27257,N_27239,N_27203);
or U27258 (N_27258,N_27051,N_27210);
or U27259 (N_27259,N_27083,N_27113);
and U27260 (N_27260,N_27027,N_27107);
xnor U27261 (N_27261,N_27202,N_27044);
or U27262 (N_27262,N_27040,N_27053);
nand U27263 (N_27263,N_27180,N_27090);
xnor U27264 (N_27264,N_27070,N_27166);
nor U27265 (N_27265,N_27224,N_27173);
xnor U27266 (N_27266,N_27214,N_27245);
xor U27267 (N_27267,N_27114,N_27140);
xnor U27268 (N_27268,N_27028,N_27208);
or U27269 (N_27269,N_27133,N_27085);
xor U27270 (N_27270,N_27153,N_27159);
xor U27271 (N_27271,N_27209,N_27073);
nand U27272 (N_27272,N_27045,N_27042);
nand U27273 (N_27273,N_27177,N_27020);
or U27274 (N_27274,N_27055,N_27235);
nand U27275 (N_27275,N_27122,N_27030);
or U27276 (N_27276,N_27188,N_27128);
or U27277 (N_27277,N_27181,N_27217);
nand U27278 (N_27278,N_27111,N_27233);
or U27279 (N_27279,N_27194,N_27244);
nand U27280 (N_27280,N_27127,N_27050);
nor U27281 (N_27281,N_27211,N_27232);
xnor U27282 (N_27282,N_27236,N_27029);
and U27283 (N_27283,N_27184,N_27062);
nand U27284 (N_27284,N_27206,N_27198);
or U27285 (N_27285,N_27079,N_27015);
nor U27286 (N_27286,N_27019,N_27216);
nor U27287 (N_27287,N_27157,N_27187);
xnor U27288 (N_27288,N_27234,N_27148);
nand U27289 (N_27289,N_27242,N_27246);
nor U27290 (N_27290,N_27013,N_27192);
and U27291 (N_27291,N_27221,N_27021);
nor U27292 (N_27292,N_27117,N_27213);
nor U27293 (N_27293,N_27047,N_27056);
or U27294 (N_27294,N_27212,N_27098);
nand U27295 (N_27295,N_27176,N_27152);
xor U27296 (N_27296,N_27186,N_27109);
nand U27297 (N_27297,N_27238,N_27125);
nand U27298 (N_27298,N_27046,N_27200);
and U27299 (N_27299,N_27072,N_27165);
xor U27300 (N_27300,N_27035,N_27110);
xor U27301 (N_27301,N_27018,N_27199);
nand U27302 (N_27302,N_27066,N_27031);
xor U27303 (N_27303,N_27179,N_27061);
and U27304 (N_27304,N_27022,N_27220);
xor U27305 (N_27305,N_27141,N_27241);
nand U27306 (N_27306,N_27077,N_27131);
and U27307 (N_27307,N_27025,N_27093);
nand U27308 (N_27308,N_27100,N_27024);
or U27309 (N_27309,N_27003,N_27150);
nor U27310 (N_27310,N_27011,N_27116);
nand U27311 (N_27311,N_27139,N_27197);
and U27312 (N_27312,N_27215,N_27191);
nor U27313 (N_27313,N_27014,N_27078);
xnor U27314 (N_27314,N_27249,N_27060);
or U27315 (N_27315,N_27204,N_27099);
or U27316 (N_27316,N_27120,N_27071);
or U27317 (N_27317,N_27016,N_27145);
nand U27318 (N_27318,N_27057,N_27174);
or U27319 (N_27319,N_27196,N_27089);
and U27320 (N_27320,N_27178,N_27143);
nor U27321 (N_27321,N_27185,N_27147);
xnor U27322 (N_27322,N_27086,N_27026);
and U27323 (N_27323,N_27048,N_27115);
nand U27324 (N_27324,N_27130,N_27222);
or U27325 (N_27325,N_27049,N_27237);
and U27326 (N_27326,N_27182,N_27158);
nor U27327 (N_27327,N_27063,N_27229);
xor U27328 (N_27328,N_27189,N_27149);
or U27329 (N_27329,N_27005,N_27193);
and U27330 (N_27330,N_27167,N_27169);
and U27331 (N_27331,N_27081,N_27102);
xor U27332 (N_27332,N_27007,N_27171);
nor U27333 (N_27333,N_27039,N_27144);
nor U27334 (N_27334,N_27074,N_27160);
nor U27335 (N_27335,N_27069,N_27036);
and U27336 (N_27336,N_27067,N_27190);
and U27337 (N_27337,N_27170,N_27201);
and U27338 (N_27338,N_27009,N_27162);
or U27339 (N_27339,N_27088,N_27136);
xor U27340 (N_27340,N_27092,N_27138);
nor U27341 (N_27341,N_27002,N_27132);
nor U27342 (N_27342,N_27155,N_27175);
and U27343 (N_27343,N_27124,N_27248);
nand U27344 (N_27344,N_27096,N_27004);
nor U27345 (N_27345,N_27076,N_27033);
xor U27346 (N_27346,N_27121,N_27163);
or U27347 (N_27347,N_27104,N_27043);
nor U27348 (N_27348,N_27094,N_27183);
xnor U27349 (N_27349,N_27243,N_27106);
nor U27350 (N_27350,N_27103,N_27038);
nor U27351 (N_27351,N_27023,N_27223);
nor U27352 (N_27352,N_27012,N_27225);
and U27353 (N_27353,N_27226,N_27195);
nor U27354 (N_27354,N_27108,N_27095);
xor U27355 (N_27355,N_27219,N_27129);
and U27356 (N_27356,N_27001,N_27010);
xnor U27357 (N_27357,N_27037,N_27161);
or U27358 (N_27358,N_27112,N_27156);
xor U27359 (N_27359,N_27084,N_27087);
or U27360 (N_27360,N_27126,N_27228);
xor U27361 (N_27361,N_27146,N_27142);
nor U27362 (N_27362,N_27058,N_27230);
xnor U27363 (N_27363,N_27034,N_27207);
nand U27364 (N_27364,N_27123,N_27105);
xor U27365 (N_27365,N_27064,N_27052);
nand U27366 (N_27366,N_27164,N_27134);
nand U27367 (N_27367,N_27017,N_27135);
nor U27368 (N_27368,N_27065,N_27054);
and U27369 (N_27369,N_27008,N_27151);
or U27370 (N_27370,N_27068,N_27097);
nor U27371 (N_27371,N_27059,N_27247);
nand U27372 (N_27372,N_27118,N_27240);
nor U27373 (N_27373,N_27101,N_27218);
or U27374 (N_27374,N_27227,N_27172);
or U27375 (N_27375,N_27177,N_27229);
or U27376 (N_27376,N_27039,N_27142);
nand U27377 (N_27377,N_27036,N_27160);
or U27378 (N_27378,N_27053,N_27144);
nand U27379 (N_27379,N_27137,N_27181);
or U27380 (N_27380,N_27182,N_27030);
nand U27381 (N_27381,N_27219,N_27196);
and U27382 (N_27382,N_27052,N_27063);
and U27383 (N_27383,N_27122,N_27006);
or U27384 (N_27384,N_27145,N_27082);
nor U27385 (N_27385,N_27206,N_27165);
nand U27386 (N_27386,N_27061,N_27103);
nor U27387 (N_27387,N_27199,N_27154);
nor U27388 (N_27388,N_27088,N_27233);
or U27389 (N_27389,N_27067,N_27163);
xnor U27390 (N_27390,N_27173,N_27198);
or U27391 (N_27391,N_27218,N_27243);
xnor U27392 (N_27392,N_27009,N_27082);
xnor U27393 (N_27393,N_27170,N_27122);
xnor U27394 (N_27394,N_27053,N_27243);
nand U27395 (N_27395,N_27168,N_27078);
and U27396 (N_27396,N_27166,N_27017);
nor U27397 (N_27397,N_27202,N_27099);
nor U27398 (N_27398,N_27094,N_27082);
nand U27399 (N_27399,N_27044,N_27124);
and U27400 (N_27400,N_27169,N_27050);
xor U27401 (N_27401,N_27082,N_27177);
or U27402 (N_27402,N_27192,N_27115);
and U27403 (N_27403,N_27054,N_27176);
nor U27404 (N_27404,N_27110,N_27166);
or U27405 (N_27405,N_27109,N_27151);
nor U27406 (N_27406,N_27033,N_27069);
or U27407 (N_27407,N_27022,N_27016);
xor U27408 (N_27408,N_27203,N_27244);
or U27409 (N_27409,N_27182,N_27153);
and U27410 (N_27410,N_27183,N_27002);
or U27411 (N_27411,N_27011,N_27204);
or U27412 (N_27412,N_27051,N_27182);
and U27413 (N_27413,N_27217,N_27007);
nand U27414 (N_27414,N_27233,N_27173);
xnor U27415 (N_27415,N_27175,N_27187);
or U27416 (N_27416,N_27182,N_27167);
and U27417 (N_27417,N_27169,N_27091);
xnor U27418 (N_27418,N_27108,N_27130);
nand U27419 (N_27419,N_27018,N_27160);
xor U27420 (N_27420,N_27033,N_27105);
xor U27421 (N_27421,N_27147,N_27050);
xor U27422 (N_27422,N_27011,N_27048);
xor U27423 (N_27423,N_27227,N_27148);
or U27424 (N_27424,N_27238,N_27090);
nor U27425 (N_27425,N_27198,N_27088);
and U27426 (N_27426,N_27226,N_27188);
xor U27427 (N_27427,N_27221,N_27056);
or U27428 (N_27428,N_27184,N_27013);
and U27429 (N_27429,N_27061,N_27115);
or U27430 (N_27430,N_27226,N_27172);
xnor U27431 (N_27431,N_27094,N_27214);
and U27432 (N_27432,N_27061,N_27207);
nor U27433 (N_27433,N_27173,N_27006);
or U27434 (N_27434,N_27172,N_27059);
nand U27435 (N_27435,N_27075,N_27050);
and U27436 (N_27436,N_27121,N_27140);
xnor U27437 (N_27437,N_27190,N_27021);
nand U27438 (N_27438,N_27028,N_27111);
and U27439 (N_27439,N_27185,N_27076);
and U27440 (N_27440,N_27073,N_27231);
nor U27441 (N_27441,N_27240,N_27166);
and U27442 (N_27442,N_27247,N_27157);
and U27443 (N_27443,N_27103,N_27195);
nor U27444 (N_27444,N_27170,N_27220);
nor U27445 (N_27445,N_27195,N_27116);
nand U27446 (N_27446,N_27110,N_27029);
and U27447 (N_27447,N_27148,N_27186);
or U27448 (N_27448,N_27003,N_27079);
nor U27449 (N_27449,N_27222,N_27029);
and U27450 (N_27450,N_27038,N_27077);
and U27451 (N_27451,N_27198,N_27116);
nor U27452 (N_27452,N_27062,N_27103);
or U27453 (N_27453,N_27167,N_27177);
nor U27454 (N_27454,N_27143,N_27141);
xnor U27455 (N_27455,N_27055,N_27129);
or U27456 (N_27456,N_27209,N_27079);
and U27457 (N_27457,N_27180,N_27245);
nor U27458 (N_27458,N_27096,N_27214);
xor U27459 (N_27459,N_27184,N_27229);
nand U27460 (N_27460,N_27023,N_27064);
xnor U27461 (N_27461,N_27169,N_27040);
and U27462 (N_27462,N_27241,N_27119);
xor U27463 (N_27463,N_27069,N_27080);
or U27464 (N_27464,N_27083,N_27034);
nor U27465 (N_27465,N_27167,N_27042);
nor U27466 (N_27466,N_27172,N_27204);
and U27467 (N_27467,N_27203,N_27182);
and U27468 (N_27468,N_27164,N_27198);
nand U27469 (N_27469,N_27116,N_27246);
nand U27470 (N_27470,N_27239,N_27097);
or U27471 (N_27471,N_27141,N_27229);
or U27472 (N_27472,N_27115,N_27229);
nand U27473 (N_27473,N_27164,N_27140);
xnor U27474 (N_27474,N_27075,N_27062);
and U27475 (N_27475,N_27070,N_27206);
nand U27476 (N_27476,N_27109,N_27028);
or U27477 (N_27477,N_27096,N_27031);
xnor U27478 (N_27478,N_27205,N_27054);
xnor U27479 (N_27479,N_27043,N_27200);
xor U27480 (N_27480,N_27106,N_27079);
and U27481 (N_27481,N_27158,N_27201);
nor U27482 (N_27482,N_27176,N_27030);
nand U27483 (N_27483,N_27118,N_27049);
and U27484 (N_27484,N_27090,N_27239);
and U27485 (N_27485,N_27186,N_27228);
or U27486 (N_27486,N_27162,N_27056);
or U27487 (N_27487,N_27200,N_27018);
or U27488 (N_27488,N_27142,N_27099);
xnor U27489 (N_27489,N_27130,N_27080);
nand U27490 (N_27490,N_27040,N_27140);
nand U27491 (N_27491,N_27040,N_27227);
nand U27492 (N_27492,N_27104,N_27222);
nand U27493 (N_27493,N_27220,N_27224);
nor U27494 (N_27494,N_27030,N_27069);
nor U27495 (N_27495,N_27140,N_27134);
nand U27496 (N_27496,N_27196,N_27020);
nor U27497 (N_27497,N_27020,N_27171);
nand U27498 (N_27498,N_27200,N_27215);
nand U27499 (N_27499,N_27219,N_27076);
and U27500 (N_27500,N_27408,N_27355);
nand U27501 (N_27501,N_27489,N_27498);
nor U27502 (N_27502,N_27478,N_27343);
nor U27503 (N_27503,N_27474,N_27416);
and U27504 (N_27504,N_27379,N_27310);
nor U27505 (N_27505,N_27324,N_27461);
and U27506 (N_27506,N_27447,N_27365);
nor U27507 (N_27507,N_27280,N_27340);
nor U27508 (N_27508,N_27465,N_27357);
and U27509 (N_27509,N_27286,N_27313);
nand U27510 (N_27510,N_27263,N_27305);
and U27511 (N_27511,N_27336,N_27428);
or U27512 (N_27512,N_27493,N_27346);
nor U27513 (N_27513,N_27470,N_27414);
xnor U27514 (N_27514,N_27393,N_27253);
or U27515 (N_27515,N_27496,N_27326);
nor U27516 (N_27516,N_27267,N_27377);
nand U27517 (N_27517,N_27456,N_27257);
and U27518 (N_27518,N_27306,N_27403);
nand U27519 (N_27519,N_27252,N_27469);
nor U27520 (N_27520,N_27423,N_27283);
and U27521 (N_27521,N_27468,N_27415);
xor U27522 (N_27522,N_27272,N_27471);
nor U27523 (N_27523,N_27342,N_27341);
nor U27524 (N_27524,N_27251,N_27400);
or U27525 (N_27525,N_27301,N_27499);
xnor U27526 (N_27526,N_27320,N_27360);
nor U27527 (N_27527,N_27262,N_27392);
and U27528 (N_27528,N_27318,N_27347);
nand U27529 (N_27529,N_27276,N_27450);
and U27530 (N_27530,N_27376,N_27390);
nand U27531 (N_27531,N_27487,N_27366);
xor U27532 (N_27532,N_27273,N_27304);
and U27533 (N_27533,N_27380,N_27473);
xor U27534 (N_27534,N_27386,N_27296);
xor U27535 (N_27535,N_27453,N_27345);
nand U27536 (N_27536,N_27282,N_27375);
xnor U27537 (N_27537,N_27410,N_27373);
and U27538 (N_27538,N_27278,N_27488);
nor U27539 (N_27539,N_27451,N_27431);
or U27540 (N_27540,N_27367,N_27307);
nand U27541 (N_27541,N_27481,N_27425);
or U27542 (N_27542,N_27427,N_27314);
nor U27543 (N_27543,N_27300,N_27391);
and U27544 (N_27544,N_27406,N_27316);
and U27545 (N_27545,N_27261,N_27479);
and U27546 (N_27546,N_27445,N_27467);
or U27547 (N_27547,N_27434,N_27435);
xor U27548 (N_27548,N_27385,N_27463);
and U27549 (N_27549,N_27363,N_27331);
nand U27550 (N_27550,N_27250,N_27480);
nor U27551 (N_27551,N_27281,N_27457);
or U27552 (N_27552,N_27420,N_27460);
xnor U27553 (N_27553,N_27477,N_27458);
xor U27554 (N_27554,N_27497,N_27402);
or U27555 (N_27555,N_27388,N_27275);
and U27556 (N_27556,N_27359,N_27309);
nor U27557 (N_27557,N_27319,N_27407);
nand U27558 (N_27558,N_27398,N_27432);
xor U27559 (N_27559,N_27449,N_27356);
xnor U27560 (N_27560,N_27344,N_27370);
nor U27561 (N_27561,N_27448,N_27285);
or U27562 (N_27562,N_27475,N_27332);
xnor U27563 (N_27563,N_27486,N_27294);
nor U27564 (N_27564,N_27494,N_27372);
and U27565 (N_27565,N_27354,N_27362);
xor U27566 (N_27566,N_27413,N_27438);
xnor U27567 (N_27567,N_27382,N_27397);
xor U27568 (N_27568,N_27446,N_27269);
and U27569 (N_27569,N_27439,N_27254);
nor U27570 (N_27570,N_27274,N_27299);
nand U27571 (N_27571,N_27312,N_27277);
xor U27572 (N_27572,N_27311,N_27337);
and U27573 (N_27573,N_27290,N_27308);
and U27574 (N_27574,N_27256,N_27315);
nor U27575 (N_27575,N_27368,N_27260);
nand U27576 (N_27576,N_27433,N_27298);
nor U27577 (N_27577,N_27335,N_27325);
and U27578 (N_27578,N_27452,N_27454);
nand U27579 (N_27579,N_27395,N_27462);
or U27580 (N_27580,N_27303,N_27411);
or U27581 (N_27581,N_27321,N_27371);
and U27582 (N_27582,N_27284,N_27255);
and U27583 (N_27583,N_27292,N_27436);
nor U27584 (N_27584,N_27264,N_27401);
and U27585 (N_27585,N_27430,N_27483);
and U27586 (N_27586,N_27327,N_27437);
xnor U27587 (N_27587,N_27330,N_27383);
or U27588 (N_27588,N_27381,N_27426);
or U27589 (N_27589,N_27492,N_27374);
nand U27590 (N_27590,N_27387,N_27389);
nor U27591 (N_27591,N_27419,N_27484);
nand U27592 (N_27592,N_27329,N_27364);
xor U27593 (N_27593,N_27418,N_27455);
nor U27594 (N_27594,N_27412,N_27409);
nand U27595 (N_27595,N_27490,N_27421);
nand U27596 (N_27596,N_27268,N_27293);
xor U27597 (N_27597,N_27287,N_27353);
and U27598 (N_27598,N_27476,N_27422);
and U27599 (N_27599,N_27482,N_27323);
and U27600 (N_27600,N_27443,N_27271);
nor U27601 (N_27601,N_27328,N_27259);
or U27602 (N_27602,N_27378,N_27350);
xor U27603 (N_27603,N_27459,N_27352);
xnor U27604 (N_27604,N_27348,N_27266);
nor U27605 (N_27605,N_27270,N_27295);
xnor U27606 (N_27606,N_27317,N_27429);
nand U27607 (N_27607,N_27440,N_27358);
and U27608 (N_27608,N_27444,N_27424);
nor U27609 (N_27609,N_27291,N_27279);
and U27610 (N_27610,N_27334,N_27495);
xor U27611 (N_27611,N_27405,N_27361);
xnor U27612 (N_27612,N_27404,N_27351);
xnor U27613 (N_27613,N_27491,N_27466);
or U27614 (N_27614,N_27265,N_27289);
or U27615 (N_27615,N_27333,N_27472);
or U27616 (N_27616,N_27384,N_27302);
or U27617 (N_27617,N_27369,N_27442);
xnor U27618 (N_27618,N_27288,N_27394);
or U27619 (N_27619,N_27485,N_27441);
xnor U27620 (N_27620,N_27297,N_27396);
or U27621 (N_27621,N_27417,N_27349);
nor U27622 (N_27622,N_27464,N_27322);
nand U27623 (N_27623,N_27338,N_27399);
or U27624 (N_27624,N_27258,N_27339);
xor U27625 (N_27625,N_27485,N_27275);
or U27626 (N_27626,N_27442,N_27379);
nand U27627 (N_27627,N_27352,N_27413);
or U27628 (N_27628,N_27399,N_27373);
nand U27629 (N_27629,N_27278,N_27344);
or U27630 (N_27630,N_27378,N_27360);
nand U27631 (N_27631,N_27434,N_27333);
nor U27632 (N_27632,N_27305,N_27416);
nor U27633 (N_27633,N_27377,N_27283);
nand U27634 (N_27634,N_27331,N_27378);
nor U27635 (N_27635,N_27432,N_27319);
nor U27636 (N_27636,N_27453,N_27315);
nor U27637 (N_27637,N_27422,N_27493);
xor U27638 (N_27638,N_27298,N_27333);
nand U27639 (N_27639,N_27305,N_27370);
nor U27640 (N_27640,N_27310,N_27485);
nand U27641 (N_27641,N_27290,N_27375);
or U27642 (N_27642,N_27288,N_27458);
nor U27643 (N_27643,N_27260,N_27349);
and U27644 (N_27644,N_27365,N_27496);
xor U27645 (N_27645,N_27410,N_27331);
nor U27646 (N_27646,N_27446,N_27252);
xor U27647 (N_27647,N_27358,N_27293);
or U27648 (N_27648,N_27255,N_27336);
nor U27649 (N_27649,N_27421,N_27315);
and U27650 (N_27650,N_27277,N_27257);
nor U27651 (N_27651,N_27492,N_27380);
nand U27652 (N_27652,N_27360,N_27329);
or U27653 (N_27653,N_27394,N_27370);
and U27654 (N_27654,N_27424,N_27490);
or U27655 (N_27655,N_27488,N_27304);
xor U27656 (N_27656,N_27442,N_27360);
nor U27657 (N_27657,N_27453,N_27357);
nand U27658 (N_27658,N_27364,N_27277);
nand U27659 (N_27659,N_27360,N_27399);
and U27660 (N_27660,N_27342,N_27302);
nor U27661 (N_27661,N_27450,N_27269);
and U27662 (N_27662,N_27333,N_27331);
or U27663 (N_27663,N_27300,N_27485);
nor U27664 (N_27664,N_27302,N_27325);
xnor U27665 (N_27665,N_27420,N_27263);
xor U27666 (N_27666,N_27307,N_27303);
xor U27667 (N_27667,N_27379,N_27346);
nor U27668 (N_27668,N_27305,N_27457);
or U27669 (N_27669,N_27381,N_27334);
or U27670 (N_27670,N_27277,N_27483);
or U27671 (N_27671,N_27353,N_27424);
nor U27672 (N_27672,N_27462,N_27307);
nand U27673 (N_27673,N_27430,N_27329);
xor U27674 (N_27674,N_27396,N_27272);
or U27675 (N_27675,N_27414,N_27467);
or U27676 (N_27676,N_27291,N_27488);
nor U27677 (N_27677,N_27356,N_27485);
nor U27678 (N_27678,N_27363,N_27277);
and U27679 (N_27679,N_27250,N_27449);
xnor U27680 (N_27680,N_27429,N_27383);
or U27681 (N_27681,N_27349,N_27409);
xnor U27682 (N_27682,N_27389,N_27470);
and U27683 (N_27683,N_27284,N_27360);
xnor U27684 (N_27684,N_27451,N_27372);
nor U27685 (N_27685,N_27403,N_27277);
and U27686 (N_27686,N_27367,N_27281);
and U27687 (N_27687,N_27381,N_27276);
xor U27688 (N_27688,N_27328,N_27422);
nor U27689 (N_27689,N_27460,N_27390);
nand U27690 (N_27690,N_27286,N_27341);
and U27691 (N_27691,N_27292,N_27460);
or U27692 (N_27692,N_27468,N_27402);
nand U27693 (N_27693,N_27445,N_27419);
or U27694 (N_27694,N_27253,N_27436);
nand U27695 (N_27695,N_27279,N_27495);
nor U27696 (N_27696,N_27268,N_27381);
or U27697 (N_27697,N_27497,N_27326);
or U27698 (N_27698,N_27441,N_27351);
or U27699 (N_27699,N_27387,N_27327);
or U27700 (N_27700,N_27320,N_27393);
xnor U27701 (N_27701,N_27255,N_27408);
and U27702 (N_27702,N_27377,N_27397);
nand U27703 (N_27703,N_27306,N_27276);
nand U27704 (N_27704,N_27453,N_27426);
or U27705 (N_27705,N_27439,N_27318);
nor U27706 (N_27706,N_27425,N_27309);
xnor U27707 (N_27707,N_27364,N_27428);
or U27708 (N_27708,N_27485,N_27403);
or U27709 (N_27709,N_27381,N_27285);
and U27710 (N_27710,N_27251,N_27463);
nor U27711 (N_27711,N_27359,N_27331);
nor U27712 (N_27712,N_27281,N_27371);
or U27713 (N_27713,N_27313,N_27447);
nor U27714 (N_27714,N_27418,N_27370);
nor U27715 (N_27715,N_27492,N_27293);
xnor U27716 (N_27716,N_27455,N_27272);
nand U27717 (N_27717,N_27483,N_27257);
and U27718 (N_27718,N_27286,N_27480);
or U27719 (N_27719,N_27441,N_27271);
nand U27720 (N_27720,N_27417,N_27467);
xor U27721 (N_27721,N_27483,N_27276);
nor U27722 (N_27722,N_27414,N_27297);
nand U27723 (N_27723,N_27295,N_27329);
nor U27724 (N_27724,N_27489,N_27406);
xor U27725 (N_27725,N_27467,N_27463);
nor U27726 (N_27726,N_27341,N_27321);
or U27727 (N_27727,N_27461,N_27378);
or U27728 (N_27728,N_27418,N_27428);
nand U27729 (N_27729,N_27269,N_27259);
nor U27730 (N_27730,N_27398,N_27285);
or U27731 (N_27731,N_27457,N_27465);
or U27732 (N_27732,N_27429,N_27389);
nor U27733 (N_27733,N_27412,N_27320);
xnor U27734 (N_27734,N_27378,N_27439);
xnor U27735 (N_27735,N_27408,N_27335);
nand U27736 (N_27736,N_27455,N_27372);
nor U27737 (N_27737,N_27422,N_27453);
xor U27738 (N_27738,N_27483,N_27269);
or U27739 (N_27739,N_27254,N_27441);
xor U27740 (N_27740,N_27425,N_27344);
xnor U27741 (N_27741,N_27484,N_27361);
and U27742 (N_27742,N_27270,N_27391);
and U27743 (N_27743,N_27315,N_27293);
and U27744 (N_27744,N_27423,N_27276);
xnor U27745 (N_27745,N_27324,N_27348);
and U27746 (N_27746,N_27478,N_27327);
xnor U27747 (N_27747,N_27466,N_27478);
and U27748 (N_27748,N_27271,N_27477);
nor U27749 (N_27749,N_27453,N_27255);
and U27750 (N_27750,N_27555,N_27669);
or U27751 (N_27751,N_27559,N_27735);
or U27752 (N_27752,N_27617,N_27534);
nand U27753 (N_27753,N_27725,N_27544);
and U27754 (N_27754,N_27740,N_27588);
nand U27755 (N_27755,N_27715,N_27631);
or U27756 (N_27756,N_27604,N_27550);
nor U27757 (N_27757,N_27719,N_27670);
or U27758 (N_27758,N_27639,N_27695);
and U27759 (N_27759,N_27523,N_27681);
and U27760 (N_27760,N_27628,N_27598);
xor U27761 (N_27761,N_27717,N_27543);
xor U27762 (N_27762,N_27612,N_27510);
and U27763 (N_27763,N_27622,N_27594);
and U27764 (N_27764,N_27660,N_27633);
xor U27765 (N_27765,N_27691,N_27658);
nor U27766 (N_27766,N_27656,N_27706);
and U27767 (N_27767,N_27745,N_27541);
and U27768 (N_27768,N_27601,N_27562);
and U27769 (N_27769,N_27698,N_27697);
nand U27770 (N_27770,N_27518,N_27565);
xnor U27771 (N_27771,N_27547,N_27690);
nor U27772 (N_27772,N_27718,N_27521);
xor U27773 (N_27773,N_27629,N_27640);
and U27774 (N_27774,N_27665,N_27539);
and U27775 (N_27775,N_27738,N_27621);
xnor U27776 (N_27776,N_27610,N_27522);
nand U27777 (N_27777,N_27636,N_27668);
and U27778 (N_27778,N_27692,N_27578);
xor U27779 (N_27779,N_27630,N_27603);
or U27780 (N_27780,N_27654,N_27552);
and U27781 (N_27781,N_27537,N_27609);
xnor U27782 (N_27782,N_27568,N_27564);
and U27783 (N_27783,N_27646,N_27508);
nor U27784 (N_27784,N_27626,N_27580);
xnor U27785 (N_27785,N_27586,N_27703);
nor U27786 (N_27786,N_27592,N_27579);
or U27787 (N_27787,N_27714,N_27666);
and U27788 (N_27788,N_27529,N_27554);
nand U27789 (N_27789,N_27584,N_27587);
nand U27790 (N_27790,N_27506,N_27701);
xnor U27791 (N_27791,N_27619,N_27672);
or U27792 (N_27792,N_27533,N_27616);
xnor U27793 (N_27793,N_27685,N_27577);
nor U27794 (N_27794,N_27595,N_27618);
and U27795 (N_27795,N_27731,N_27657);
nand U27796 (N_27796,N_27560,N_27641);
nand U27797 (N_27797,N_27608,N_27570);
nor U27798 (N_27798,N_27540,N_27737);
nand U27799 (N_27799,N_27536,N_27749);
xnor U27800 (N_27800,N_27707,N_27642);
and U27801 (N_27801,N_27556,N_27591);
nand U27802 (N_27802,N_27661,N_27596);
nor U27803 (N_27803,N_27553,N_27651);
nor U27804 (N_27804,N_27652,N_27676);
nand U27805 (N_27805,N_27500,N_27585);
nor U27806 (N_27806,N_27513,N_27509);
xnor U27807 (N_27807,N_27730,N_27746);
or U27808 (N_27808,N_27597,N_27527);
xor U27809 (N_27809,N_27512,N_27615);
nand U27810 (N_27810,N_27627,N_27671);
nor U27811 (N_27811,N_27674,N_27732);
nand U27812 (N_27812,N_27687,N_27572);
and U27813 (N_27813,N_27503,N_27724);
nor U27814 (N_27814,N_27741,N_27748);
and U27815 (N_27815,N_27611,N_27590);
nand U27816 (N_27816,N_27520,N_27542);
xnor U27817 (N_27817,N_27699,N_27532);
nand U27818 (N_27818,N_27624,N_27727);
nand U27819 (N_27819,N_27643,N_27678);
nand U27820 (N_27820,N_27736,N_27721);
xnor U27821 (N_27821,N_27659,N_27515);
or U27822 (N_27822,N_27504,N_27632);
xor U27823 (N_27823,N_27589,N_27593);
nor U27824 (N_27824,N_27648,N_27729);
and U27825 (N_27825,N_27647,N_27655);
xor U27826 (N_27826,N_27667,N_27576);
or U27827 (N_27827,N_27720,N_27525);
or U27828 (N_27828,N_27742,N_27571);
nand U27829 (N_27829,N_27583,N_27519);
or U27830 (N_27830,N_27558,N_27623);
xor U27831 (N_27831,N_27514,N_27682);
or U27832 (N_27832,N_27602,N_27502);
nor U27833 (N_27833,N_27634,N_27511);
xor U27834 (N_27834,N_27620,N_27705);
and U27835 (N_27835,N_27600,N_27744);
nor U27836 (N_27836,N_27694,N_27528);
nand U27837 (N_27837,N_27650,N_27723);
nor U27838 (N_27838,N_27644,N_27574);
and U27839 (N_27839,N_27722,N_27702);
nor U27840 (N_27840,N_27675,N_27734);
nand U27841 (N_27841,N_27739,N_27551);
and U27842 (N_27842,N_27563,N_27663);
nor U27843 (N_27843,N_27505,N_27566);
and U27844 (N_27844,N_27517,N_27747);
and U27845 (N_27845,N_27613,N_27726);
xor U27846 (N_27846,N_27545,N_27662);
nor U27847 (N_27847,N_27581,N_27743);
nor U27848 (N_27848,N_27653,N_27625);
nor U27849 (N_27849,N_27501,N_27546);
nor U27850 (N_27850,N_27686,N_27649);
nor U27851 (N_27851,N_27688,N_27689);
nor U27852 (N_27852,N_27716,N_27683);
nand U27853 (N_27853,N_27679,N_27607);
and U27854 (N_27854,N_27549,N_27704);
and U27855 (N_27855,N_27561,N_27645);
and U27856 (N_27856,N_27709,N_27713);
or U27857 (N_27857,N_27733,N_27573);
nand U27858 (N_27858,N_27516,N_27684);
xor U27859 (N_27859,N_27728,N_27567);
nand U27860 (N_27860,N_27524,N_27693);
and U27861 (N_27861,N_27538,N_27664);
and U27862 (N_27862,N_27531,N_27548);
xor U27863 (N_27863,N_27526,N_27535);
nand U27864 (N_27864,N_27614,N_27599);
or U27865 (N_27865,N_27530,N_27708);
xor U27866 (N_27866,N_27710,N_27673);
nor U27867 (N_27867,N_27637,N_27569);
or U27868 (N_27868,N_27696,N_27680);
xnor U27869 (N_27869,N_27635,N_27557);
or U27870 (N_27870,N_27711,N_27638);
nand U27871 (N_27871,N_27712,N_27677);
and U27872 (N_27872,N_27507,N_27700);
xnor U27873 (N_27873,N_27582,N_27605);
xnor U27874 (N_27874,N_27575,N_27606);
or U27875 (N_27875,N_27708,N_27652);
or U27876 (N_27876,N_27504,N_27558);
and U27877 (N_27877,N_27708,N_27589);
nand U27878 (N_27878,N_27708,N_27580);
nor U27879 (N_27879,N_27673,N_27669);
nand U27880 (N_27880,N_27679,N_27684);
or U27881 (N_27881,N_27580,N_27733);
xor U27882 (N_27882,N_27571,N_27525);
xor U27883 (N_27883,N_27621,N_27629);
xnor U27884 (N_27884,N_27603,N_27614);
nor U27885 (N_27885,N_27630,N_27730);
nand U27886 (N_27886,N_27534,N_27667);
and U27887 (N_27887,N_27544,N_27683);
and U27888 (N_27888,N_27571,N_27660);
nand U27889 (N_27889,N_27605,N_27667);
or U27890 (N_27890,N_27609,N_27579);
xnor U27891 (N_27891,N_27552,N_27500);
xnor U27892 (N_27892,N_27579,N_27634);
xor U27893 (N_27893,N_27597,N_27653);
and U27894 (N_27894,N_27654,N_27723);
nand U27895 (N_27895,N_27523,N_27717);
xor U27896 (N_27896,N_27711,N_27512);
or U27897 (N_27897,N_27562,N_27549);
nand U27898 (N_27898,N_27737,N_27588);
nor U27899 (N_27899,N_27673,N_27571);
and U27900 (N_27900,N_27679,N_27500);
xor U27901 (N_27901,N_27710,N_27593);
nor U27902 (N_27902,N_27514,N_27619);
nor U27903 (N_27903,N_27643,N_27670);
and U27904 (N_27904,N_27730,N_27609);
and U27905 (N_27905,N_27701,N_27681);
xor U27906 (N_27906,N_27626,N_27514);
nor U27907 (N_27907,N_27535,N_27656);
nor U27908 (N_27908,N_27531,N_27684);
nand U27909 (N_27909,N_27696,N_27748);
and U27910 (N_27910,N_27701,N_27626);
nor U27911 (N_27911,N_27748,N_27673);
nand U27912 (N_27912,N_27662,N_27694);
nor U27913 (N_27913,N_27651,N_27704);
and U27914 (N_27914,N_27694,N_27651);
nand U27915 (N_27915,N_27731,N_27622);
xor U27916 (N_27916,N_27533,N_27571);
or U27917 (N_27917,N_27554,N_27503);
or U27918 (N_27918,N_27611,N_27648);
and U27919 (N_27919,N_27627,N_27696);
nor U27920 (N_27920,N_27549,N_27729);
nand U27921 (N_27921,N_27664,N_27644);
xor U27922 (N_27922,N_27601,N_27650);
nor U27923 (N_27923,N_27719,N_27749);
and U27924 (N_27924,N_27574,N_27714);
nor U27925 (N_27925,N_27584,N_27515);
nor U27926 (N_27926,N_27737,N_27677);
and U27927 (N_27927,N_27700,N_27593);
nor U27928 (N_27928,N_27574,N_27576);
or U27929 (N_27929,N_27609,N_27572);
nor U27930 (N_27930,N_27635,N_27680);
nand U27931 (N_27931,N_27706,N_27725);
and U27932 (N_27932,N_27553,N_27732);
or U27933 (N_27933,N_27690,N_27733);
nand U27934 (N_27934,N_27615,N_27721);
or U27935 (N_27935,N_27578,N_27665);
nor U27936 (N_27936,N_27556,N_27580);
nor U27937 (N_27937,N_27676,N_27506);
xor U27938 (N_27938,N_27574,N_27564);
nand U27939 (N_27939,N_27528,N_27633);
nand U27940 (N_27940,N_27647,N_27508);
nand U27941 (N_27941,N_27710,N_27713);
nand U27942 (N_27942,N_27503,N_27647);
or U27943 (N_27943,N_27744,N_27523);
xor U27944 (N_27944,N_27503,N_27588);
nand U27945 (N_27945,N_27546,N_27631);
and U27946 (N_27946,N_27719,N_27524);
nand U27947 (N_27947,N_27716,N_27583);
xor U27948 (N_27948,N_27626,N_27670);
or U27949 (N_27949,N_27669,N_27693);
and U27950 (N_27950,N_27645,N_27743);
or U27951 (N_27951,N_27562,N_27604);
nor U27952 (N_27952,N_27550,N_27514);
xnor U27953 (N_27953,N_27733,N_27689);
nand U27954 (N_27954,N_27716,N_27561);
nor U27955 (N_27955,N_27675,N_27580);
xnor U27956 (N_27956,N_27743,N_27561);
and U27957 (N_27957,N_27537,N_27740);
nand U27958 (N_27958,N_27734,N_27569);
and U27959 (N_27959,N_27718,N_27596);
or U27960 (N_27960,N_27573,N_27575);
nand U27961 (N_27961,N_27733,N_27560);
or U27962 (N_27962,N_27577,N_27523);
nor U27963 (N_27963,N_27536,N_27532);
and U27964 (N_27964,N_27576,N_27562);
and U27965 (N_27965,N_27546,N_27542);
xnor U27966 (N_27966,N_27582,N_27718);
nand U27967 (N_27967,N_27696,N_27573);
xor U27968 (N_27968,N_27632,N_27591);
nor U27969 (N_27969,N_27643,N_27558);
nor U27970 (N_27970,N_27721,N_27700);
nand U27971 (N_27971,N_27569,N_27668);
or U27972 (N_27972,N_27556,N_27699);
xor U27973 (N_27973,N_27632,N_27661);
nor U27974 (N_27974,N_27696,N_27584);
nand U27975 (N_27975,N_27553,N_27500);
or U27976 (N_27976,N_27576,N_27523);
and U27977 (N_27977,N_27652,N_27581);
and U27978 (N_27978,N_27726,N_27619);
or U27979 (N_27979,N_27686,N_27522);
and U27980 (N_27980,N_27598,N_27679);
and U27981 (N_27981,N_27607,N_27650);
nand U27982 (N_27982,N_27556,N_27734);
xnor U27983 (N_27983,N_27539,N_27675);
nand U27984 (N_27984,N_27649,N_27527);
and U27985 (N_27985,N_27719,N_27744);
or U27986 (N_27986,N_27583,N_27504);
nor U27987 (N_27987,N_27683,N_27545);
and U27988 (N_27988,N_27559,N_27523);
or U27989 (N_27989,N_27576,N_27578);
or U27990 (N_27990,N_27582,N_27586);
or U27991 (N_27991,N_27711,N_27618);
nand U27992 (N_27992,N_27665,N_27561);
nor U27993 (N_27993,N_27599,N_27717);
and U27994 (N_27994,N_27533,N_27635);
nand U27995 (N_27995,N_27622,N_27521);
or U27996 (N_27996,N_27660,N_27723);
or U27997 (N_27997,N_27577,N_27520);
nor U27998 (N_27998,N_27730,N_27739);
xnor U27999 (N_27999,N_27616,N_27600);
nand U28000 (N_28000,N_27966,N_27932);
nand U28001 (N_28001,N_27829,N_27839);
nand U28002 (N_28002,N_27833,N_27888);
nor U28003 (N_28003,N_27838,N_27946);
nor U28004 (N_28004,N_27837,N_27766);
nor U28005 (N_28005,N_27930,N_27952);
and U28006 (N_28006,N_27773,N_27830);
nor U28007 (N_28007,N_27910,N_27974);
nor U28008 (N_28008,N_27863,N_27812);
nand U28009 (N_28009,N_27769,N_27789);
nand U28010 (N_28010,N_27751,N_27827);
and U28011 (N_28011,N_27855,N_27750);
xor U28012 (N_28012,N_27818,N_27921);
and U28013 (N_28013,N_27851,N_27931);
xor U28014 (N_28014,N_27872,N_27788);
or U28015 (N_28015,N_27896,N_27879);
nand U28016 (N_28016,N_27997,N_27983);
and U28017 (N_28017,N_27858,N_27962);
nor U28018 (N_28018,N_27850,N_27980);
nand U28019 (N_28019,N_27813,N_27984);
nor U28020 (N_28020,N_27893,N_27913);
xnor U28021 (N_28021,N_27860,N_27944);
nand U28022 (N_28022,N_27982,N_27809);
and U28023 (N_28023,N_27808,N_27897);
and U28024 (N_28024,N_27757,N_27903);
or U28025 (N_28025,N_27994,N_27935);
nor U28026 (N_28026,N_27759,N_27940);
nor U28027 (N_28027,N_27906,N_27995);
nand U28028 (N_28028,N_27965,N_27802);
nand U28029 (N_28029,N_27928,N_27968);
xor U28030 (N_28030,N_27760,N_27848);
nor U28031 (N_28031,N_27817,N_27895);
nand U28032 (N_28032,N_27753,N_27991);
nor U28033 (N_28033,N_27956,N_27794);
or U28034 (N_28034,N_27902,N_27987);
or U28035 (N_28035,N_27894,N_27937);
xnor U28036 (N_28036,N_27876,N_27811);
or U28037 (N_28037,N_27779,N_27970);
xnor U28038 (N_28038,N_27865,N_27887);
nor U28039 (N_28039,N_27907,N_27804);
xnor U28040 (N_28040,N_27862,N_27852);
nor U28041 (N_28041,N_27960,N_27972);
nor U28042 (N_28042,N_27923,N_27803);
or U28043 (N_28043,N_27990,N_27824);
nand U28044 (N_28044,N_27868,N_27800);
and U28045 (N_28045,N_27986,N_27786);
xor U28046 (N_28046,N_27909,N_27853);
or U28047 (N_28047,N_27752,N_27978);
nand U28048 (N_28048,N_27774,N_27880);
nand U28049 (N_28049,N_27927,N_27941);
nor U28050 (N_28050,N_27875,N_27967);
and U28051 (N_28051,N_27775,N_27840);
nor U28052 (N_28052,N_27924,N_27768);
nand U28053 (N_28053,N_27918,N_27951);
and U28054 (N_28054,N_27831,N_27975);
nor U28055 (N_28055,N_27976,N_27754);
xor U28056 (N_28056,N_27806,N_27797);
nand U28057 (N_28057,N_27943,N_27816);
and U28058 (N_28058,N_27771,N_27917);
or U28059 (N_28059,N_27993,N_27845);
nor U28060 (N_28060,N_27796,N_27825);
xnor U28061 (N_28061,N_27905,N_27864);
xnor U28062 (N_28062,N_27799,N_27959);
or U28063 (N_28063,N_27755,N_27866);
and U28064 (N_28064,N_27847,N_27820);
or U28065 (N_28065,N_27792,N_27949);
nand U28066 (N_28066,N_27871,N_27869);
and U28067 (N_28067,N_27971,N_27836);
nand U28068 (N_28068,N_27947,N_27914);
nor U28069 (N_28069,N_27762,N_27882);
xor U28070 (N_28070,N_27964,N_27929);
and U28071 (N_28071,N_27989,N_27841);
nand U28072 (N_28072,N_27854,N_27878);
and U28073 (N_28073,N_27898,N_27822);
or U28074 (N_28074,N_27828,N_27890);
nand U28075 (N_28075,N_27843,N_27857);
or U28076 (N_28076,N_27870,N_27798);
and U28077 (N_28077,N_27916,N_27778);
and U28078 (N_28078,N_27973,N_27945);
or U28079 (N_28079,N_27958,N_27790);
nand U28080 (N_28080,N_27874,N_27992);
xor U28081 (N_28081,N_27933,N_27904);
and U28082 (N_28082,N_27784,N_27996);
and U28083 (N_28083,N_27957,N_27782);
nand U28084 (N_28084,N_27919,N_27846);
nand U28085 (N_28085,N_27781,N_27849);
nand U28086 (N_28086,N_27998,N_27892);
and U28087 (N_28087,N_27787,N_27765);
or U28088 (N_28088,N_27805,N_27908);
nand U28089 (N_28089,N_27936,N_27891);
nand U28090 (N_28090,N_27915,N_27777);
nor U28091 (N_28091,N_27901,N_27793);
and U28092 (N_28092,N_27954,N_27770);
nand U28093 (N_28093,N_27810,N_27939);
or U28094 (N_28094,N_27884,N_27926);
nand U28095 (N_28095,N_27867,N_27819);
nand U28096 (N_28096,N_27785,N_27912);
nand U28097 (N_28097,N_27881,N_27856);
xnor U28098 (N_28098,N_27934,N_27823);
and U28099 (N_28099,N_27969,N_27885);
or U28100 (N_28100,N_27981,N_27938);
or U28101 (N_28101,N_27767,N_27756);
or U28102 (N_28102,N_27999,N_27859);
or U28103 (N_28103,N_27795,N_27955);
nor U28104 (N_28104,N_27801,N_27977);
or U28105 (N_28105,N_27776,N_27780);
xnor U28106 (N_28106,N_27889,N_27950);
nand U28107 (N_28107,N_27861,N_27922);
nor U28108 (N_28108,N_27758,N_27988);
and U28109 (N_28109,N_27883,N_27835);
or U28110 (N_28110,N_27900,N_27772);
nand U28111 (N_28111,N_27807,N_27844);
xnor U28112 (N_28112,N_27832,N_27783);
xnor U28113 (N_28113,N_27826,N_27764);
or U28114 (N_28114,N_27877,N_27985);
nand U28115 (N_28115,N_27961,N_27791);
and U28116 (N_28116,N_27979,N_27815);
xnor U28117 (N_28117,N_27761,N_27821);
nand U28118 (N_28118,N_27814,N_27873);
xor U28119 (N_28119,N_27963,N_27911);
or U28120 (N_28120,N_27899,N_27834);
and U28121 (N_28121,N_27925,N_27842);
nand U28122 (N_28122,N_27948,N_27942);
nor U28123 (N_28123,N_27920,N_27886);
and U28124 (N_28124,N_27953,N_27763);
and U28125 (N_28125,N_27884,N_27851);
xnor U28126 (N_28126,N_27933,N_27993);
and U28127 (N_28127,N_27891,N_27947);
or U28128 (N_28128,N_27844,N_27952);
xor U28129 (N_28129,N_27942,N_27930);
xor U28130 (N_28130,N_27906,N_27985);
or U28131 (N_28131,N_27965,N_27817);
and U28132 (N_28132,N_27827,N_27934);
and U28133 (N_28133,N_27834,N_27752);
nand U28134 (N_28134,N_27977,N_27850);
nand U28135 (N_28135,N_27836,N_27819);
nand U28136 (N_28136,N_27861,N_27984);
xnor U28137 (N_28137,N_27908,N_27968);
nand U28138 (N_28138,N_27792,N_27804);
and U28139 (N_28139,N_27924,N_27993);
and U28140 (N_28140,N_27874,N_27894);
or U28141 (N_28141,N_27835,N_27937);
and U28142 (N_28142,N_27996,N_27852);
nand U28143 (N_28143,N_27996,N_27878);
nand U28144 (N_28144,N_27792,N_27955);
nand U28145 (N_28145,N_27849,N_27895);
or U28146 (N_28146,N_27950,N_27847);
nand U28147 (N_28147,N_27955,N_27866);
nand U28148 (N_28148,N_27924,N_27873);
nor U28149 (N_28149,N_27875,N_27937);
or U28150 (N_28150,N_27881,N_27953);
xor U28151 (N_28151,N_27809,N_27902);
and U28152 (N_28152,N_27960,N_27881);
xnor U28153 (N_28153,N_27903,N_27800);
nand U28154 (N_28154,N_27768,N_27834);
xnor U28155 (N_28155,N_27765,N_27866);
xor U28156 (N_28156,N_27783,N_27889);
nor U28157 (N_28157,N_27969,N_27953);
or U28158 (N_28158,N_27773,N_27763);
nor U28159 (N_28159,N_27930,N_27884);
or U28160 (N_28160,N_27816,N_27837);
nor U28161 (N_28161,N_27886,N_27797);
nor U28162 (N_28162,N_27983,N_27757);
nor U28163 (N_28163,N_27811,N_27895);
nor U28164 (N_28164,N_27988,N_27857);
nor U28165 (N_28165,N_27892,N_27994);
xnor U28166 (N_28166,N_27917,N_27915);
nand U28167 (N_28167,N_27759,N_27805);
xor U28168 (N_28168,N_27935,N_27980);
nor U28169 (N_28169,N_27779,N_27842);
nand U28170 (N_28170,N_27986,N_27824);
xnor U28171 (N_28171,N_27900,N_27783);
nor U28172 (N_28172,N_27834,N_27925);
nor U28173 (N_28173,N_27754,N_27931);
and U28174 (N_28174,N_27752,N_27842);
nand U28175 (N_28175,N_27954,N_27898);
and U28176 (N_28176,N_27941,N_27979);
nand U28177 (N_28177,N_27842,N_27977);
nand U28178 (N_28178,N_27978,N_27831);
xor U28179 (N_28179,N_27829,N_27959);
or U28180 (N_28180,N_27897,N_27856);
and U28181 (N_28181,N_27856,N_27981);
and U28182 (N_28182,N_27965,N_27933);
nor U28183 (N_28183,N_27839,N_27999);
xor U28184 (N_28184,N_27917,N_27859);
nor U28185 (N_28185,N_27796,N_27858);
nand U28186 (N_28186,N_27832,N_27828);
nand U28187 (N_28187,N_27798,N_27889);
nand U28188 (N_28188,N_27819,N_27782);
and U28189 (N_28189,N_27971,N_27876);
and U28190 (N_28190,N_27849,N_27753);
or U28191 (N_28191,N_27989,N_27894);
and U28192 (N_28192,N_27802,N_27969);
and U28193 (N_28193,N_27790,N_27872);
nand U28194 (N_28194,N_27778,N_27858);
xor U28195 (N_28195,N_27972,N_27916);
nor U28196 (N_28196,N_27900,N_27940);
nor U28197 (N_28197,N_27801,N_27872);
and U28198 (N_28198,N_27880,N_27833);
and U28199 (N_28199,N_27889,N_27870);
nor U28200 (N_28200,N_27848,N_27926);
xnor U28201 (N_28201,N_27868,N_27792);
nand U28202 (N_28202,N_27906,N_27996);
or U28203 (N_28203,N_27847,N_27845);
xor U28204 (N_28204,N_27837,N_27998);
xnor U28205 (N_28205,N_27872,N_27844);
nand U28206 (N_28206,N_27937,N_27887);
or U28207 (N_28207,N_27796,N_27775);
or U28208 (N_28208,N_27934,N_27926);
nor U28209 (N_28209,N_27915,N_27997);
and U28210 (N_28210,N_27883,N_27804);
nand U28211 (N_28211,N_27992,N_27865);
nor U28212 (N_28212,N_27819,N_27854);
xnor U28213 (N_28213,N_27953,N_27884);
xor U28214 (N_28214,N_27971,N_27870);
and U28215 (N_28215,N_27862,N_27835);
nor U28216 (N_28216,N_27958,N_27767);
xor U28217 (N_28217,N_27921,N_27879);
xnor U28218 (N_28218,N_27762,N_27890);
xnor U28219 (N_28219,N_27845,N_27967);
nor U28220 (N_28220,N_27780,N_27900);
xor U28221 (N_28221,N_27875,N_27793);
xnor U28222 (N_28222,N_27900,N_27998);
nand U28223 (N_28223,N_27943,N_27768);
and U28224 (N_28224,N_27937,N_27782);
and U28225 (N_28225,N_27935,N_27813);
xor U28226 (N_28226,N_27958,N_27934);
nor U28227 (N_28227,N_27873,N_27825);
or U28228 (N_28228,N_27987,N_27977);
nand U28229 (N_28229,N_27838,N_27790);
nor U28230 (N_28230,N_27777,N_27782);
and U28231 (N_28231,N_27878,N_27881);
nor U28232 (N_28232,N_27859,N_27900);
nor U28233 (N_28233,N_27808,N_27757);
nand U28234 (N_28234,N_27829,N_27882);
nor U28235 (N_28235,N_27917,N_27890);
nand U28236 (N_28236,N_27901,N_27915);
xnor U28237 (N_28237,N_27946,N_27992);
or U28238 (N_28238,N_27997,N_27932);
or U28239 (N_28239,N_27965,N_27832);
nor U28240 (N_28240,N_27921,N_27892);
and U28241 (N_28241,N_27967,N_27784);
xor U28242 (N_28242,N_27803,N_27886);
and U28243 (N_28243,N_27836,N_27974);
nand U28244 (N_28244,N_27964,N_27838);
nor U28245 (N_28245,N_27852,N_27887);
nor U28246 (N_28246,N_27845,N_27823);
and U28247 (N_28247,N_27981,N_27926);
nand U28248 (N_28248,N_27814,N_27933);
xnor U28249 (N_28249,N_27982,N_27750);
xor U28250 (N_28250,N_28039,N_28058);
nor U28251 (N_28251,N_28127,N_28089);
or U28252 (N_28252,N_28168,N_28050);
nor U28253 (N_28253,N_28170,N_28204);
nor U28254 (N_28254,N_28099,N_28003);
nor U28255 (N_28255,N_28198,N_28147);
xnor U28256 (N_28256,N_28228,N_28231);
or U28257 (N_28257,N_28104,N_28017);
nand U28258 (N_28258,N_28229,N_28012);
xor U28259 (N_28259,N_28035,N_28100);
nand U28260 (N_28260,N_28013,N_28016);
xnor U28261 (N_28261,N_28019,N_28116);
and U28262 (N_28262,N_28227,N_28194);
or U28263 (N_28263,N_28059,N_28037);
nand U28264 (N_28264,N_28180,N_28062);
nor U28265 (N_28265,N_28021,N_28165);
nor U28266 (N_28266,N_28000,N_28036);
xnor U28267 (N_28267,N_28055,N_28191);
and U28268 (N_28268,N_28072,N_28075);
nand U28269 (N_28269,N_28189,N_28232);
xor U28270 (N_28270,N_28132,N_28096);
nor U28271 (N_28271,N_28137,N_28034);
or U28272 (N_28272,N_28225,N_28217);
and U28273 (N_28273,N_28131,N_28077);
and U28274 (N_28274,N_28084,N_28029);
and U28275 (N_28275,N_28094,N_28120);
nand U28276 (N_28276,N_28209,N_28106);
xnor U28277 (N_28277,N_28242,N_28134);
nor U28278 (N_28278,N_28133,N_28230);
nor U28279 (N_28279,N_28161,N_28074);
or U28280 (N_28280,N_28102,N_28219);
or U28281 (N_28281,N_28244,N_28070);
or U28282 (N_28282,N_28163,N_28175);
nand U28283 (N_28283,N_28157,N_28066);
xor U28284 (N_28284,N_28117,N_28093);
nor U28285 (N_28285,N_28090,N_28152);
xor U28286 (N_28286,N_28248,N_28026);
and U28287 (N_28287,N_28042,N_28060);
nor U28288 (N_28288,N_28190,N_28142);
nor U28289 (N_28289,N_28164,N_28174);
or U28290 (N_28290,N_28202,N_28136);
nand U28291 (N_28291,N_28140,N_28171);
xor U28292 (N_28292,N_28154,N_28101);
nor U28293 (N_28293,N_28078,N_28246);
nand U28294 (N_28294,N_28008,N_28226);
nand U28295 (N_28295,N_28151,N_28193);
xor U28296 (N_28296,N_28109,N_28239);
or U28297 (N_28297,N_28129,N_28097);
or U28298 (N_28298,N_28192,N_28179);
nand U28299 (N_28299,N_28150,N_28218);
nand U28300 (N_28300,N_28088,N_28201);
nor U28301 (N_28301,N_28033,N_28169);
xnor U28302 (N_28302,N_28085,N_28023);
nand U28303 (N_28303,N_28153,N_28046);
nand U28304 (N_28304,N_28249,N_28022);
and U28305 (N_28305,N_28122,N_28160);
nand U28306 (N_28306,N_28095,N_28119);
nor U28307 (N_28307,N_28025,N_28213);
nor U28308 (N_28308,N_28079,N_28112);
nor U28309 (N_28309,N_28144,N_28172);
and U28310 (N_28310,N_28222,N_28238);
and U28311 (N_28311,N_28098,N_28240);
xor U28312 (N_28312,N_28107,N_28203);
nand U28313 (N_28313,N_28032,N_28247);
or U28314 (N_28314,N_28123,N_28241);
nand U28315 (N_28315,N_28148,N_28138);
nor U28316 (N_28316,N_28212,N_28205);
nor U28317 (N_28317,N_28155,N_28080);
nand U28318 (N_28318,N_28235,N_28038);
or U28319 (N_28319,N_28221,N_28063);
and U28320 (N_28320,N_28141,N_28052);
xnor U28321 (N_28321,N_28182,N_28068);
and U28322 (N_28322,N_28234,N_28001);
or U28323 (N_28323,N_28159,N_28224);
or U28324 (N_28324,N_28030,N_28043);
or U28325 (N_28325,N_28196,N_28002);
nand U28326 (N_28326,N_28158,N_28197);
or U28327 (N_28327,N_28200,N_28214);
or U28328 (N_28328,N_28211,N_28091);
and U28329 (N_28329,N_28236,N_28128);
or U28330 (N_28330,N_28135,N_28092);
nor U28331 (N_28331,N_28048,N_28215);
xor U28332 (N_28332,N_28114,N_28024);
nand U28333 (N_28333,N_28031,N_28208);
xor U28334 (N_28334,N_28108,N_28071);
nand U28335 (N_28335,N_28145,N_28040);
nand U28336 (N_28336,N_28124,N_28139);
xor U28337 (N_28337,N_28210,N_28005);
nor U28338 (N_28338,N_28207,N_28081);
xnor U28339 (N_28339,N_28020,N_28176);
and U28340 (N_28340,N_28177,N_28199);
or U28341 (N_28341,N_28045,N_28105);
nand U28342 (N_28342,N_28237,N_28186);
nand U28343 (N_28343,N_28167,N_28121);
and U28344 (N_28344,N_28110,N_28014);
nor U28345 (N_28345,N_28166,N_28051);
or U28346 (N_28346,N_28028,N_28067);
xnor U28347 (N_28347,N_28007,N_28056);
xor U28348 (N_28348,N_28027,N_28156);
nor U28349 (N_28349,N_28216,N_28183);
and U28350 (N_28350,N_28018,N_28086);
or U28351 (N_28351,N_28126,N_28004);
and U28352 (N_28352,N_28125,N_28206);
and U28353 (N_28353,N_28130,N_28041);
or U28354 (N_28354,N_28184,N_28223);
nand U28355 (N_28355,N_28069,N_28220);
nor U28356 (N_28356,N_28149,N_28015);
nand U28357 (N_28357,N_28173,N_28009);
and U28358 (N_28358,N_28233,N_28178);
nand U28359 (N_28359,N_28083,N_28087);
nand U28360 (N_28360,N_28073,N_28162);
and U28361 (N_28361,N_28195,N_28187);
and U28362 (N_28362,N_28011,N_28061);
nand U28363 (N_28363,N_28054,N_28245);
or U28364 (N_28364,N_28146,N_28113);
nor U28365 (N_28365,N_28006,N_28053);
or U28366 (N_28366,N_28057,N_28044);
or U28367 (N_28367,N_28143,N_28185);
nor U28368 (N_28368,N_28064,N_28010);
and U28369 (N_28369,N_28047,N_28111);
nand U28370 (N_28370,N_28181,N_28103);
or U28371 (N_28371,N_28082,N_28115);
xnor U28372 (N_28372,N_28188,N_28243);
xnor U28373 (N_28373,N_28049,N_28076);
or U28374 (N_28374,N_28118,N_28065);
xnor U28375 (N_28375,N_28138,N_28025);
or U28376 (N_28376,N_28029,N_28088);
and U28377 (N_28377,N_28168,N_28146);
nand U28378 (N_28378,N_28182,N_28106);
xnor U28379 (N_28379,N_28073,N_28185);
nand U28380 (N_28380,N_28107,N_28102);
nand U28381 (N_28381,N_28196,N_28058);
or U28382 (N_28382,N_28009,N_28000);
or U28383 (N_28383,N_28194,N_28043);
nand U28384 (N_28384,N_28097,N_28062);
nor U28385 (N_28385,N_28224,N_28032);
or U28386 (N_28386,N_28179,N_28199);
nor U28387 (N_28387,N_28229,N_28241);
nand U28388 (N_28388,N_28037,N_28109);
nor U28389 (N_28389,N_28089,N_28167);
xor U28390 (N_28390,N_28089,N_28079);
nor U28391 (N_28391,N_28098,N_28018);
and U28392 (N_28392,N_28014,N_28177);
nand U28393 (N_28393,N_28119,N_28237);
and U28394 (N_28394,N_28007,N_28145);
and U28395 (N_28395,N_28112,N_28039);
xnor U28396 (N_28396,N_28202,N_28192);
nor U28397 (N_28397,N_28097,N_28005);
or U28398 (N_28398,N_28075,N_28013);
and U28399 (N_28399,N_28163,N_28136);
nand U28400 (N_28400,N_28222,N_28105);
nor U28401 (N_28401,N_28136,N_28074);
or U28402 (N_28402,N_28052,N_28233);
nor U28403 (N_28403,N_28098,N_28211);
or U28404 (N_28404,N_28161,N_28118);
nor U28405 (N_28405,N_28067,N_28021);
xnor U28406 (N_28406,N_28128,N_28000);
or U28407 (N_28407,N_28186,N_28006);
or U28408 (N_28408,N_28111,N_28172);
nand U28409 (N_28409,N_28036,N_28016);
nor U28410 (N_28410,N_28239,N_28002);
and U28411 (N_28411,N_28108,N_28122);
and U28412 (N_28412,N_28125,N_28024);
nand U28413 (N_28413,N_28089,N_28006);
or U28414 (N_28414,N_28147,N_28163);
nand U28415 (N_28415,N_28211,N_28170);
and U28416 (N_28416,N_28180,N_28079);
nor U28417 (N_28417,N_28051,N_28160);
nor U28418 (N_28418,N_28159,N_28049);
or U28419 (N_28419,N_28083,N_28217);
nor U28420 (N_28420,N_28006,N_28084);
nand U28421 (N_28421,N_28134,N_28104);
and U28422 (N_28422,N_28119,N_28142);
nand U28423 (N_28423,N_28045,N_28102);
xnor U28424 (N_28424,N_28109,N_28107);
xor U28425 (N_28425,N_28221,N_28001);
xnor U28426 (N_28426,N_28089,N_28107);
nor U28427 (N_28427,N_28067,N_28043);
xnor U28428 (N_28428,N_28196,N_28104);
or U28429 (N_28429,N_28136,N_28125);
xnor U28430 (N_28430,N_28016,N_28018);
and U28431 (N_28431,N_28171,N_28041);
or U28432 (N_28432,N_28111,N_28144);
xnor U28433 (N_28433,N_28088,N_28152);
or U28434 (N_28434,N_28086,N_28181);
or U28435 (N_28435,N_28147,N_28041);
or U28436 (N_28436,N_28237,N_28219);
or U28437 (N_28437,N_28096,N_28231);
or U28438 (N_28438,N_28068,N_28032);
xnor U28439 (N_28439,N_28036,N_28149);
nand U28440 (N_28440,N_28144,N_28016);
nor U28441 (N_28441,N_28017,N_28088);
xor U28442 (N_28442,N_28020,N_28195);
nor U28443 (N_28443,N_28192,N_28152);
nand U28444 (N_28444,N_28176,N_28075);
nor U28445 (N_28445,N_28088,N_28037);
nand U28446 (N_28446,N_28058,N_28164);
nor U28447 (N_28447,N_28065,N_28000);
and U28448 (N_28448,N_28019,N_28122);
and U28449 (N_28449,N_28118,N_28159);
or U28450 (N_28450,N_28244,N_28117);
or U28451 (N_28451,N_28157,N_28162);
nor U28452 (N_28452,N_28242,N_28109);
and U28453 (N_28453,N_28026,N_28139);
nand U28454 (N_28454,N_28049,N_28160);
and U28455 (N_28455,N_28209,N_28079);
nand U28456 (N_28456,N_28173,N_28225);
and U28457 (N_28457,N_28097,N_28244);
or U28458 (N_28458,N_28114,N_28029);
xor U28459 (N_28459,N_28057,N_28125);
and U28460 (N_28460,N_28042,N_28090);
nor U28461 (N_28461,N_28056,N_28228);
and U28462 (N_28462,N_28102,N_28161);
or U28463 (N_28463,N_28102,N_28072);
nor U28464 (N_28464,N_28151,N_28095);
nand U28465 (N_28465,N_28104,N_28248);
or U28466 (N_28466,N_28077,N_28014);
or U28467 (N_28467,N_28162,N_28116);
and U28468 (N_28468,N_28198,N_28186);
or U28469 (N_28469,N_28054,N_28136);
nand U28470 (N_28470,N_28025,N_28112);
xnor U28471 (N_28471,N_28216,N_28151);
xor U28472 (N_28472,N_28214,N_28194);
xnor U28473 (N_28473,N_28239,N_28048);
xor U28474 (N_28474,N_28211,N_28122);
nor U28475 (N_28475,N_28129,N_28191);
nor U28476 (N_28476,N_28075,N_28167);
nand U28477 (N_28477,N_28019,N_28200);
or U28478 (N_28478,N_28209,N_28014);
nand U28479 (N_28479,N_28226,N_28227);
xor U28480 (N_28480,N_28156,N_28187);
nand U28481 (N_28481,N_28179,N_28163);
nand U28482 (N_28482,N_28076,N_28099);
and U28483 (N_28483,N_28150,N_28187);
nor U28484 (N_28484,N_28173,N_28031);
nor U28485 (N_28485,N_28002,N_28153);
and U28486 (N_28486,N_28091,N_28081);
nor U28487 (N_28487,N_28060,N_28216);
nand U28488 (N_28488,N_28085,N_28220);
nand U28489 (N_28489,N_28018,N_28171);
and U28490 (N_28490,N_28116,N_28171);
or U28491 (N_28491,N_28206,N_28085);
and U28492 (N_28492,N_28048,N_28218);
and U28493 (N_28493,N_28195,N_28178);
xnor U28494 (N_28494,N_28220,N_28110);
and U28495 (N_28495,N_28181,N_28118);
xor U28496 (N_28496,N_28143,N_28053);
nand U28497 (N_28497,N_28056,N_28217);
nand U28498 (N_28498,N_28184,N_28032);
and U28499 (N_28499,N_28180,N_28104);
and U28500 (N_28500,N_28360,N_28438);
or U28501 (N_28501,N_28459,N_28380);
nor U28502 (N_28502,N_28485,N_28398);
nor U28503 (N_28503,N_28257,N_28314);
and U28504 (N_28504,N_28357,N_28392);
and U28505 (N_28505,N_28287,N_28431);
and U28506 (N_28506,N_28325,N_28426);
nand U28507 (N_28507,N_28283,N_28267);
and U28508 (N_28508,N_28490,N_28331);
nor U28509 (N_28509,N_28302,N_28341);
and U28510 (N_28510,N_28338,N_28400);
and U28511 (N_28511,N_28448,N_28407);
or U28512 (N_28512,N_28434,N_28273);
xor U28513 (N_28513,N_28411,N_28296);
xor U28514 (N_28514,N_28297,N_28252);
xnor U28515 (N_28515,N_28362,N_28498);
nand U28516 (N_28516,N_28343,N_28479);
and U28517 (N_28517,N_28387,N_28437);
nand U28518 (N_28518,N_28310,N_28488);
or U28519 (N_28519,N_28424,N_28404);
and U28520 (N_28520,N_28394,N_28429);
nand U28521 (N_28521,N_28332,N_28319);
or U28522 (N_28522,N_28378,N_28369);
xnor U28523 (N_28523,N_28250,N_28290);
nor U28524 (N_28524,N_28337,N_28251);
and U28525 (N_28525,N_28432,N_28408);
xnor U28526 (N_28526,N_28323,N_28457);
nand U28527 (N_28527,N_28427,N_28326);
xnor U28528 (N_28528,N_28266,N_28307);
and U28529 (N_28529,N_28300,N_28350);
or U28530 (N_28530,N_28253,N_28286);
nand U28531 (N_28531,N_28476,N_28306);
and U28532 (N_28532,N_28414,N_28347);
and U28533 (N_28533,N_28418,N_28329);
nand U28534 (N_28534,N_28409,N_28368);
nor U28535 (N_28535,N_28288,N_28340);
or U28536 (N_28536,N_28475,N_28322);
nand U28537 (N_28537,N_28358,N_28452);
or U28538 (N_28538,N_28443,N_28393);
nor U28539 (N_28539,N_28342,N_28352);
and U28540 (N_28540,N_28416,N_28367);
xor U28541 (N_28541,N_28487,N_28374);
and U28542 (N_28542,N_28395,N_28466);
or U28543 (N_28543,N_28497,N_28399);
xor U28544 (N_28544,N_28462,N_28481);
nor U28545 (N_28545,N_28436,N_28413);
and U28546 (N_28546,N_28441,N_28385);
nor U28547 (N_28547,N_28363,N_28349);
or U28548 (N_28548,N_28495,N_28335);
nand U28549 (N_28549,N_28269,N_28460);
xnor U28550 (N_28550,N_28461,N_28280);
xnor U28551 (N_28551,N_28346,N_28327);
or U28552 (N_28552,N_28276,N_28491);
nor U28553 (N_28553,N_28318,N_28405);
nand U28554 (N_28554,N_28447,N_28486);
nor U28555 (N_28555,N_28333,N_28410);
xnor U28556 (N_28556,N_28371,N_28263);
xor U28557 (N_28557,N_28305,N_28469);
nand U28558 (N_28558,N_28451,N_28417);
nor U28559 (N_28559,N_28389,N_28454);
nor U28560 (N_28560,N_28477,N_28388);
and U28561 (N_28561,N_28391,N_28463);
xor U28562 (N_28562,N_28375,N_28428);
nor U28563 (N_28563,N_28317,N_28261);
nor U28564 (N_28564,N_28401,N_28474);
nor U28565 (N_28565,N_28382,N_28489);
nor U28566 (N_28566,N_28284,N_28456);
or U28567 (N_28567,N_28278,N_28311);
and U28568 (N_28568,N_28468,N_28397);
nand U28569 (N_28569,N_28402,N_28336);
nor U28570 (N_28570,N_28364,N_28258);
nor U28571 (N_28571,N_28376,N_28422);
or U28572 (N_28572,N_28496,N_28270);
nor U28573 (N_28573,N_28442,N_28445);
nor U28574 (N_28574,N_28262,N_28268);
xnor U28575 (N_28575,N_28455,N_28361);
xnor U28576 (N_28576,N_28282,N_28366);
nand U28577 (N_28577,N_28379,N_28386);
and U28578 (N_28578,N_28419,N_28472);
nor U28579 (N_28579,N_28345,N_28499);
and U28580 (N_28580,N_28313,N_28420);
nor U28581 (N_28581,N_28471,N_28449);
and U28582 (N_28582,N_28274,N_28493);
or U28583 (N_28583,N_28275,N_28298);
and U28584 (N_28584,N_28315,N_28285);
nor U28585 (N_28585,N_28467,N_28439);
xnor U28586 (N_28586,N_28295,N_28265);
and U28587 (N_28587,N_28425,N_28264);
and U28588 (N_28588,N_28355,N_28435);
nand U28589 (N_28589,N_28450,N_28309);
or U28590 (N_28590,N_28464,N_28365);
or U28591 (N_28591,N_28301,N_28272);
nor U28592 (N_28592,N_28377,N_28344);
and U28593 (N_28593,N_28421,N_28255);
nand U28594 (N_28594,N_28321,N_28293);
nand U28595 (N_28595,N_28353,N_28312);
xor U28596 (N_28596,N_28444,N_28390);
nand U28597 (N_28597,N_28415,N_28440);
nor U28598 (N_28598,N_28348,N_28470);
nand U28599 (N_28599,N_28383,N_28292);
or U28600 (N_28600,N_28354,N_28433);
and U28601 (N_28601,N_28289,N_28316);
and U28602 (N_28602,N_28494,N_28423);
nand U28603 (N_28603,N_28484,N_28320);
nor U28604 (N_28604,N_28473,N_28372);
xor U28605 (N_28605,N_28370,N_28330);
or U28606 (N_28606,N_28373,N_28359);
nor U28607 (N_28607,N_28254,N_28328);
or U28608 (N_28608,N_28351,N_28304);
xnor U28609 (N_28609,N_28483,N_28446);
nand U28610 (N_28610,N_28277,N_28256);
xnor U28611 (N_28611,N_28260,N_28406);
or U28612 (N_28612,N_28403,N_28279);
nor U28613 (N_28613,N_28412,N_28381);
and U28614 (N_28614,N_28356,N_28465);
or U28615 (N_28615,N_28339,N_28281);
xor U28616 (N_28616,N_28430,N_28259);
or U28617 (N_28617,N_28396,N_28482);
xnor U28618 (N_28618,N_28303,N_28308);
xnor U28619 (N_28619,N_28384,N_28299);
and U28620 (N_28620,N_28291,N_28453);
nand U28621 (N_28621,N_28294,N_28480);
or U28622 (N_28622,N_28478,N_28334);
xor U28623 (N_28623,N_28271,N_28324);
nor U28624 (N_28624,N_28458,N_28492);
nand U28625 (N_28625,N_28468,N_28364);
xor U28626 (N_28626,N_28306,N_28360);
or U28627 (N_28627,N_28257,N_28450);
or U28628 (N_28628,N_28318,N_28280);
and U28629 (N_28629,N_28482,N_28498);
nor U28630 (N_28630,N_28281,N_28407);
or U28631 (N_28631,N_28287,N_28456);
and U28632 (N_28632,N_28479,N_28282);
or U28633 (N_28633,N_28367,N_28344);
nor U28634 (N_28634,N_28323,N_28483);
and U28635 (N_28635,N_28481,N_28463);
nand U28636 (N_28636,N_28356,N_28358);
and U28637 (N_28637,N_28454,N_28395);
xor U28638 (N_28638,N_28258,N_28450);
nor U28639 (N_28639,N_28433,N_28490);
xnor U28640 (N_28640,N_28433,N_28349);
nand U28641 (N_28641,N_28414,N_28389);
nor U28642 (N_28642,N_28443,N_28403);
xor U28643 (N_28643,N_28445,N_28463);
or U28644 (N_28644,N_28392,N_28340);
and U28645 (N_28645,N_28355,N_28338);
or U28646 (N_28646,N_28286,N_28469);
xnor U28647 (N_28647,N_28417,N_28325);
xnor U28648 (N_28648,N_28486,N_28265);
nor U28649 (N_28649,N_28315,N_28293);
or U28650 (N_28650,N_28375,N_28265);
or U28651 (N_28651,N_28367,N_28345);
or U28652 (N_28652,N_28299,N_28456);
nand U28653 (N_28653,N_28497,N_28335);
or U28654 (N_28654,N_28474,N_28266);
or U28655 (N_28655,N_28437,N_28313);
or U28656 (N_28656,N_28450,N_28268);
and U28657 (N_28657,N_28463,N_28323);
and U28658 (N_28658,N_28447,N_28309);
nor U28659 (N_28659,N_28360,N_28434);
xnor U28660 (N_28660,N_28390,N_28328);
nor U28661 (N_28661,N_28307,N_28377);
and U28662 (N_28662,N_28254,N_28401);
nand U28663 (N_28663,N_28488,N_28397);
or U28664 (N_28664,N_28323,N_28462);
nand U28665 (N_28665,N_28429,N_28473);
xor U28666 (N_28666,N_28433,N_28420);
nor U28667 (N_28667,N_28315,N_28494);
nand U28668 (N_28668,N_28285,N_28499);
nor U28669 (N_28669,N_28305,N_28395);
nand U28670 (N_28670,N_28470,N_28489);
nor U28671 (N_28671,N_28399,N_28362);
xor U28672 (N_28672,N_28289,N_28352);
nor U28673 (N_28673,N_28289,N_28357);
nor U28674 (N_28674,N_28407,N_28464);
or U28675 (N_28675,N_28350,N_28452);
and U28676 (N_28676,N_28315,N_28307);
xnor U28677 (N_28677,N_28486,N_28433);
or U28678 (N_28678,N_28306,N_28334);
and U28679 (N_28679,N_28281,N_28253);
xor U28680 (N_28680,N_28458,N_28392);
and U28681 (N_28681,N_28342,N_28443);
or U28682 (N_28682,N_28367,N_28458);
and U28683 (N_28683,N_28285,N_28376);
nand U28684 (N_28684,N_28397,N_28395);
xnor U28685 (N_28685,N_28347,N_28279);
nor U28686 (N_28686,N_28252,N_28473);
and U28687 (N_28687,N_28327,N_28267);
xnor U28688 (N_28688,N_28293,N_28260);
and U28689 (N_28689,N_28373,N_28409);
or U28690 (N_28690,N_28457,N_28313);
nand U28691 (N_28691,N_28261,N_28376);
or U28692 (N_28692,N_28262,N_28336);
or U28693 (N_28693,N_28458,N_28356);
and U28694 (N_28694,N_28381,N_28255);
xor U28695 (N_28695,N_28301,N_28407);
or U28696 (N_28696,N_28362,N_28471);
nand U28697 (N_28697,N_28294,N_28298);
nor U28698 (N_28698,N_28379,N_28253);
nand U28699 (N_28699,N_28494,N_28400);
nand U28700 (N_28700,N_28380,N_28392);
xnor U28701 (N_28701,N_28324,N_28346);
and U28702 (N_28702,N_28421,N_28277);
and U28703 (N_28703,N_28420,N_28456);
nand U28704 (N_28704,N_28380,N_28353);
xnor U28705 (N_28705,N_28430,N_28484);
and U28706 (N_28706,N_28341,N_28254);
nand U28707 (N_28707,N_28329,N_28430);
nor U28708 (N_28708,N_28375,N_28330);
or U28709 (N_28709,N_28470,N_28313);
nand U28710 (N_28710,N_28259,N_28418);
xor U28711 (N_28711,N_28465,N_28289);
nand U28712 (N_28712,N_28427,N_28296);
and U28713 (N_28713,N_28419,N_28380);
nor U28714 (N_28714,N_28476,N_28316);
xnor U28715 (N_28715,N_28420,N_28414);
xor U28716 (N_28716,N_28270,N_28426);
xor U28717 (N_28717,N_28343,N_28364);
or U28718 (N_28718,N_28445,N_28430);
and U28719 (N_28719,N_28320,N_28409);
or U28720 (N_28720,N_28358,N_28460);
or U28721 (N_28721,N_28337,N_28472);
nand U28722 (N_28722,N_28253,N_28304);
nor U28723 (N_28723,N_28278,N_28369);
xnor U28724 (N_28724,N_28360,N_28333);
nor U28725 (N_28725,N_28300,N_28416);
nand U28726 (N_28726,N_28269,N_28376);
nor U28727 (N_28727,N_28405,N_28257);
or U28728 (N_28728,N_28471,N_28381);
nand U28729 (N_28729,N_28368,N_28353);
and U28730 (N_28730,N_28417,N_28391);
or U28731 (N_28731,N_28270,N_28389);
xnor U28732 (N_28732,N_28428,N_28440);
and U28733 (N_28733,N_28474,N_28353);
nand U28734 (N_28734,N_28479,N_28482);
nand U28735 (N_28735,N_28479,N_28347);
nor U28736 (N_28736,N_28408,N_28472);
or U28737 (N_28737,N_28426,N_28342);
nand U28738 (N_28738,N_28471,N_28371);
nor U28739 (N_28739,N_28474,N_28461);
nand U28740 (N_28740,N_28341,N_28261);
or U28741 (N_28741,N_28482,N_28345);
or U28742 (N_28742,N_28308,N_28425);
xor U28743 (N_28743,N_28261,N_28365);
xor U28744 (N_28744,N_28387,N_28289);
or U28745 (N_28745,N_28420,N_28378);
or U28746 (N_28746,N_28345,N_28469);
and U28747 (N_28747,N_28463,N_28300);
xor U28748 (N_28748,N_28328,N_28303);
or U28749 (N_28749,N_28287,N_28408);
nand U28750 (N_28750,N_28646,N_28636);
nand U28751 (N_28751,N_28552,N_28549);
nor U28752 (N_28752,N_28654,N_28740);
xnor U28753 (N_28753,N_28745,N_28672);
or U28754 (N_28754,N_28650,N_28719);
xnor U28755 (N_28755,N_28603,N_28660);
nand U28756 (N_28756,N_28706,N_28592);
or U28757 (N_28757,N_28517,N_28583);
or U28758 (N_28758,N_28553,N_28689);
and U28759 (N_28759,N_28716,N_28604);
and U28760 (N_28760,N_28627,N_28713);
or U28761 (N_28761,N_28653,N_28561);
or U28762 (N_28762,N_28584,N_28743);
nor U28763 (N_28763,N_28709,N_28649);
or U28764 (N_28764,N_28500,N_28548);
nor U28765 (N_28765,N_28718,N_28564);
nand U28766 (N_28766,N_28593,N_28519);
nor U28767 (N_28767,N_28511,N_28566);
and U28768 (N_28768,N_28739,N_28568);
nor U28769 (N_28769,N_28712,N_28622);
or U28770 (N_28770,N_28619,N_28656);
nor U28771 (N_28771,N_28736,N_28687);
or U28772 (N_28772,N_28645,N_28721);
xor U28773 (N_28773,N_28682,N_28608);
nand U28774 (N_28774,N_28698,N_28557);
xor U28775 (N_28775,N_28697,N_28588);
nand U28776 (N_28776,N_28547,N_28641);
nand U28777 (N_28777,N_28741,N_28554);
nor U28778 (N_28778,N_28711,N_28628);
nor U28779 (N_28779,N_28731,N_28556);
xor U28780 (N_28780,N_28727,N_28528);
and U28781 (N_28781,N_28701,N_28675);
nand U28782 (N_28782,N_28642,N_28742);
xnor U28783 (N_28783,N_28532,N_28668);
and U28784 (N_28784,N_28691,N_28508);
xor U28785 (N_28785,N_28598,N_28550);
xor U28786 (N_28786,N_28633,N_28587);
xor U28787 (N_28787,N_28722,N_28522);
nor U28788 (N_28788,N_28529,N_28572);
nor U28789 (N_28789,N_28504,N_28678);
and U28790 (N_28790,N_28509,N_28733);
and U28791 (N_28791,N_28600,N_28667);
xnor U28792 (N_28792,N_28664,N_28541);
xnor U28793 (N_28793,N_28501,N_28703);
and U28794 (N_28794,N_28670,N_28637);
nor U28795 (N_28795,N_28720,N_28735);
nor U28796 (N_28796,N_28558,N_28662);
nor U28797 (N_28797,N_28589,N_28734);
nor U28798 (N_28798,N_28574,N_28702);
or U28799 (N_28799,N_28674,N_28505);
or U28800 (N_28800,N_28624,N_28671);
xnor U28801 (N_28801,N_28611,N_28516);
and U28802 (N_28802,N_28643,N_28575);
nand U28803 (N_28803,N_28616,N_28669);
nor U28804 (N_28804,N_28620,N_28638);
and U28805 (N_28805,N_28591,N_28676);
and U28806 (N_28806,N_28684,N_28730);
nand U28807 (N_28807,N_28699,N_28596);
nand U28808 (N_28808,N_28614,N_28537);
or U28809 (N_28809,N_28565,N_28524);
or U28810 (N_28810,N_28714,N_28521);
and U28811 (N_28811,N_28673,N_28573);
or U28812 (N_28812,N_28530,N_28729);
xor U28813 (N_28813,N_28724,N_28681);
xnor U28814 (N_28814,N_28562,N_28690);
nor U28815 (N_28815,N_28635,N_28526);
nand U28816 (N_28816,N_28748,N_28700);
nand U28817 (N_28817,N_28694,N_28749);
or U28818 (N_28818,N_28594,N_28560);
nor U28819 (N_28819,N_28546,N_28513);
nor U28820 (N_28820,N_28514,N_28567);
nand U28821 (N_28821,N_28677,N_28686);
nand U28822 (N_28822,N_28580,N_28585);
xor U28823 (N_28823,N_28531,N_28538);
nor U28824 (N_28824,N_28602,N_28696);
nand U28825 (N_28825,N_28606,N_28577);
nand U28826 (N_28826,N_28520,N_28655);
and U28827 (N_28827,N_28623,N_28680);
or U28828 (N_28828,N_28540,N_28597);
or U28829 (N_28829,N_28595,N_28502);
nand U28830 (N_28830,N_28579,N_28618);
xnor U28831 (N_28831,N_28648,N_28609);
xor U28832 (N_28832,N_28640,N_28551);
xor U28833 (N_28833,N_28525,N_28617);
nand U28834 (N_28834,N_28651,N_28578);
or U28835 (N_28835,N_28659,N_28663);
or U28836 (N_28836,N_28527,N_28570);
and U28837 (N_28837,N_28576,N_28536);
or U28838 (N_28838,N_28679,N_28738);
nor U28839 (N_28839,N_28644,N_28632);
and U28840 (N_28840,N_28705,N_28590);
nand U28841 (N_28841,N_28657,N_28661);
nor U28842 (N_28842,N_28539,N_28605);
nor U28843 (N_28843,N_28555,N_28544);
nor U28844 (N_28844,N_28563,N_28685);
and U28845 (N_28845,N_28518,N_28629);
nor U28846 (N_28846,N_28732,N_28723);
xnor U28847 (N_28847,N_28746,N_28559);
or U28848 (N_28848,N_28631,N_28535);
and U28849 (N_28849,N_28634,N_28613);
and U28850 (N_28850,N_28639,N_28692);
or U28851 (N_28851,N_28545,N_28515);
nor U28852 (N_28852,N_28652,N_28534);
nand U28853 (N_28853,N_28601,N_28510);
xnor U28854 (N_28854,N_28704,N_28610);
nor U28855 (N_28855,N_28630,N_28715);
nor U28856 (N_28856,N_28728,N_28647);
xor U28857 (N_28857,N_28542,N_28665);
and U28858 (N_28858,N_28621,N_28581);
xor U28859 (N_28859,N_28717,N_28708);
or U28860 (N_28860,N_28737,N_28707);
and U28861 (N_28861,N_28666,N_28512);
or U28862 (N_28862,N_28658,N_28543);
and U28863 (N_28863,N_28607,N_28582);
xnor U28864 (N_28864,N_28693,N_28725);
or U28865 (N_28865,N_28710,N_28506);
nor U28866 (N_28866,N_28683,N_28586);
xnor U28867 (N_28867,N_28571,N_28695);
and U28868 (N_28868,N_28747,N_28744);
nor U28869 (N_28869,N_28507,N_28726);
nor U28870 (N_28870,N_28625,N_28523);
xnor U28871 (N_28871,N_28569,N_28599);
nand U28872 (N_28872,N_28533,N_28612);
xor U28873 (N_28873,N_28688,N_28615);
nand U28874 (N_28874,N_28503,N_28626);
nand U28875 (N_28875,N_28690,N_28522);
or U28876 (N_28876,N_28536,N_28654);
and U28877 (N_28877,N_28544,N_28521);
nor U28878 (N_28878,N_28569,N_28543);
or U28879 (N_28879,N_28594,N_28651);
xor U28880 (N_28880,N_28503,N_28642);
nand U28881 (N_28881,N_28589,N_28651);
nor U28882 (N_28882,N_28698,N_28614);
and U28883 (N_28883,N_28666,N_28709);
nand U28884 (N_28884,N_28717,N_28605);
nor U28885 (N_28885,N_28704,N_28506);
nor U28886 (N_28886,N_28738,N_28653);
nand U28887 (N_28887,N_28503,N_28545);
nor U28888 (N_28888,N_28566,N_28707);
nor U28889 (N_28889,N_28613,N_28688);
and U28890 (N_28890,N_28573,N_28694);
nand U28891 (N_28891,N_28714,N_28548);
and U28892 (N_28892,N_28652,N_28708);
nor U28893 (N_28893,N_28639,N_28663);
nand U28894 (N_28894,N_28673,N_28592);
or U28895 (N_28895,N_28743,N_28533);
nor U28896 (N_28896,N_28714,N_28713);
xnor U28897 (N_28897,N_28533,N_28666);
nor U28898 (N_28898,N_28678,N_28684);
nand U28899 (N_28899,N_28720,N_28541);
xor U28900 (N_28900,N_28699,N_28728);
and U28901 (N_28901,N_28559,N_28715);
xor U28902 (N_28902,N_28747,N_28626);
nor U28903 (N_28903,N_28748,N_28743);
or U28904 (N_28904,N_28744,N_28688);
and U28905 (N_28905,N_28544,N_28700);
nor U28906 (N_28906,N_28567,N_28624);
nor U28907 (N_28907,N_28589,N_28574);
or U28908 (N_28908,N_28678,N_28523);
xnor U28909 (N_28909,N_28525,N_28539);
or U28910 (N_28910,N_28645,N_28742);
nor U28911 (N_28911,N_28563,N_28648);
nand U28912 (N_28912,N_28727,N_28510);
xnor U28913 (N_28913,N_28723,N_28617);
xnor U28914 (N_28914,N_28639,N_28657);
and U28915 (N_28915,N_28621,N_28559);
xnor U28916 (N_28916,N_28632,N_28525);
nor U28917 (N_28917,N_28518,N_28538);
nor U28918 (N_28918,N_28653,N_28733);
nand U28919 (N_28919,N_28700,N_28737);
xor U28920 (N_28920,N_28734,N_28745);
and U28921 (N_28921,N_28576,N_28574);
and U28922 (N_28922,N_28704,N_28740);
and U28923 (N_28923,N_28672,N_28636);
nor U28924 (N_28924,N_28518,N_28708);
or U28925 (N_28925,N_28535,N_28528);
nand U28926 (N_28926,N_28635,N_28601);
nor U28927 (N_28927,N_28580,N_28723);
nor U28928 (N_28928,N_28712,N_28602);
or U28929 (N_28929,N_28503,N_28676);
and U28930 (N_28930,N_28562,N_28747);
xnor U28931 (N_28931,N_28593,N_28635);
xor U28932 (N_28932,N_28720,N_28501);
xnor U28933 (N_28933,N_28640,N_28694);
and U28934 (N_28934,N_28508,N_28521);
and U28935 (N_28935,N_28726,N_28584);
nor U28936 (N_28936,N_28531,N_28657);
nand U28937 (N_28937,N_28521,N_28560);
xor U28938 (N_28938,N_28634,N_28704);
xor U28939 (N_28939,N_28691,N_28619);
and U28940 (N_28940,N_28743,N_28687);
xnor U28941 (N_28941,N_28506,N_28562);
nand U28942 (N_28942,N_28671,N_28676);
or U28943 (N_28943,N_28502,N_28684);
or U28944 (N_28944,N_28560,N_28554);
nand U28945 (N_28945,N_28692,N_28674);
nor U28946 (N_28946,N_28613,N_28578);
xor U28947 (N_28947,N_28578,N_28518);
and U28948 (N_28948,N_28615,N_28691);
and U28949 (N_28949,N_28718,N_28532);
or U28950 (N_28950,N_28660,N_28512);
nor U28951 (N_28951,N_28530,N_28747);
nand U28952 (N_28952,N_28666,N_28653);
nand U28953 (N_28953,N_28710,N_28741);
xnor U28954 (N_28954,N_28561,N_28615);
and U28955 (N_28955,N_28695,N_28685);
or U28956 (N_28956,N_28743,N_28645);
and U28957 (N_28957,N_28585,N_28597);
xnor U28958 (N_28958,N_28556,N_28597);
or U28959 (N_28959,N_28622,N_28583);
and U28960 (N_28960,N_28543,N_28699);
xor U28961 (N_28961,N_28698,N_28584);
or U28962 (N_28962,N_28616,N_28576);
nor U28963 (N_28963,N_28682,N_28525);
or U28964 (N_28964,N_28592,N_28650);
nor U28965 (N_28965,N_28514,N_28706);
or U28966 (N_28966,N_28619,N_28566);
nor U28967 (N_28967,N_28633,N_28563);
nor U28968 (N_28968,N_28665,N_28534);
or U28969 (N_28969,N_28654,N_28557);
and U28970 (N_28970,N_28574,N_28689);
nand U28971 (N_28971,N_28508,N_28503);
nand U28972 (N_28972,N_28549,N_28675);
nor U28973 (N_28973,N_28593,N_28569);
and U28974 (N_28974,N_28608,N_28620);
nand U28975 (N_28975,N_28636,N_28551);
and U28976 (N_28976,N_28718,N_28597);
or U28977 (N_28977,N_28714,N_28747);
nand U28978 (N_28978,N_28518,N_28568);
nor U28979 (N_28979,N_28623,N_28660);
nand U28980 (N_28980,N_28573,N_28514);
nand U28981 (N_28981,N_28544,N_28708);
or U28982 (N_28982,N_28627,N_28563);
xnor U28983 (N_28983,N_28653,N_28622);
xnor U28984 (N_28984,N_28725,N_28673);
xnor U28985 (N_28985,N_28666,N_28544);
nand U28986 (N_28986,N_28700,N_28720);
xnor U28987 (N_28987,N_28663,N_28556);
xor U28988 (N_28988,N_28652,N_28624);
nor U28989 (N_28989,N_28590,N_28701);
xnor U28990 (N_28990,N_28653,N_28690);
and U28991 (N_28991,N_28509,N_28660);
nand U28992 (N_28992,N_28522,N_28540);
and U28993 (N_28993,N_28503,N_28528);
and U28994 (N_28994,N_28743,N_28529);
xnor U28995 (N_28995,N_28637,N_28690);
or U28996 (N_28996,N_28718,N_28639);
and U28997 (N_28997,N_28729,N_28748);
nand U28998 (N_28998,N_28629,N_28685);
xor U28999 (N_28999,N_28592,N_28652);
nand U29000 (N_29000,N_28990,N_28834);
and U29001 (N_29001,N_28765,N_28924);
nand U29002 (N_29002,N_28968,N_28867);
or U29003 (N_29003,N_28768,N_28777);
nor U29004 (N_29004,N_28947,N_28987);
nor U29005 (N_29005,N_28852,N_28979);
nor U29006 (N_29006,N_28848,N_28950);
or U29007 (N_29007,N_28815,N_28915);
and U29008 (N_29008,N_28778,N_28920);
and U29009 (N_29009,N_28873,N_28955);
nand U29010 (N_29010,N_28750,N_28788);
or U29011 (N_29011,N_28994,N_28981);
or U29012 (N_29012,N_28818,N_28829);
nor U29013 (N_29013,N_28830,N_28996);
xnor U29014 (N_29014,N_28886,N_28881);
nand U29015 (N_29015,N_28930,N_28806);
or U29016 (N_29016,N_28808,N_28801);
nand U29017 (N_29017,N_28870,N_28980);
xnor U29018 (N_29018,N_28841,N_28842);
and U29019 (N_29019,N_28856,N_28911);
nand U29020 (N_29020,N_28913,N_28900);
nor U29021 (N_29021,N_28902,N_28962);
and U29022 (N_29022,N_28876,N_28995);
or U29023 (N_29023,N_28901,N_28991);
or U29024 (N_29024,N_28757,N_28763);
xnor U29025 (N_29025,N_28928,N_28916);
nor U29026 (N_29026,N_28820,N_28756);
nor U29027 (N_29027,N_28824,N_28932);
or U29028 (N_29028,N_28758,N_28957);
xnor U29029 (N_29029,N_28967,N_28851);
nand U29030 (N_29030,N_28847,N_28940);
or U29031 (N_29031,N_28944,N_28952);
and U29032 (N_29032,N_28893,N_28988);
xor U29033 (N_29033,N_28906,N_28759);
nor U29034 (N_29034,N_28752,N_28878);
xor U29035 (N_29035,N_28896,N_28821);
xnor U29036 (N_29036,N_28754,N_28814);
nor U29037 (N_29037,N_28840,N_28976);
or U29038 (N_29038,N_28838,N_28882);
xor U29039 (N_29039,N_28927,N_28983);
nor U29040 (N_29040,N_28938,N_28942);
nor U29041 (N_29041,N_28799,N_28890);
or U29042 (N_29042,N_28796,N_28800);
nand U29043 (N_29043,N_28850,N_28958);
nand U29044 (N_29044,N_28827,N_28934);
nand U29045 (N_29045,N_28992,N_28953);
xor U29046 (N_29046,N_28753,N_28889);
or U29047 (N_29047,N_28937,N_28964);
nor U29048 (N_29048,N_28929,N_28872);
nor U29049 (N_29049,N_28833,N_28959);
nor U29050 (N_29050,N_28971,N_28977);
or U29051 (N_29051,N_28898,N_28844);
xor U29052 (N_29052,N_28855,N_28899);
nand U29053 (N_29053,N_28892,N_28935);
nand U29054 (N_29054,N_28787,N_28772);
or U29055 (N_29055,N_28868,N_28897);
and U29056 (N_29056,N_28776,N_28779);
or U29057 (N_29057,N_28880,N_28925);
nor U29058 (N_29058,N_28907,N_28963);
nand U29059 (N_29059,N_28939,N_28862);
or U29060 (N_29060,N_28807,N_28773);
xnor U29061 (N_29061,N_28861,N_28798);
xor U29062 (N_29062,N_28770,N_28978);
nor U29063 (N_29063,N_28946,N_28780);
and U29064 (N_29064,N_28914,N_28917);
and U29065 (N_29065,N_28970,N_28831);
or U29066 (N_29066,N_28982,N_28986);
nor U29067 (N_29067,N_28943,N_28822);
nand U29068 (N_29068,N_28909,N_28767);
or U29069 (N_29069,N_28766,N_28974);
and U29070 (N_29070,N_28854,N_28999);
nor U29071 (N_29071,N_28904,N_28972);
and U29072 (N_29072,N_28954,N_28863);
xor U29073 (N_29073,N_28797,N_28812);
or U29074 (N_29074,N_28866,N_28793);
and U29075 (N_29075,N_28794,N_28837);
nor U29076 (N_29076,N_28804,N_28966);
and U29077 (N_29077,N_28923,N_28858);
xnor U29078 (N_29078,N_28984,N_28998);
or U29079 (N_29079,N_28997,N_28823);
xor U29080 (N_29080,N_28985,N_28951);
or U29081 (N_29081,N_28921,N_28805);
or U29082 (N_29082,N_28956,N_28771);
xor U29083 (N_29083,N_28884,N_28869);
xor U29084 (N_29084,N_28859,N_28933);
nor U29085 (N_29085,N_28762,N_28922);
nand U29086 (N_29086,N_28769,N_28993);
or U29087 (N_29087,N_28908,N_28912);
xor U29088 (N_29088,N_28816,N_28857);
nand U29089 (N_29089,N_28883,N_28860);
xor U29090 (N_29090,N_28751,N_28784);
or U29091 (N_29091,N_28969,N_28755);
and U29092 (N_29092,N_28760,N_28948);
nor U29093 (N_29093,N_28960,N_28845);
and U29094 (N_29094,N_28775,N_28918);
xor U29095 (N_29095,N_28973,N_28802);
nand U29096 (N_29096,N_28817,N_28828);
nand U29097 (N_29097,N_28903,N_28782);
xor U29098 (N_29098,N_28864,N_28809);
nand U29099 (N_29099,N_28891,N_28910);
nor U29100 (N_29100,N_28888,N_28961);
xnor U29101 (N_29101,N_28849,N_28803);
nand U29102 (N_29102,N_28786,N_28781);
nor U29103 (N_29103,N_28894,N_28832);
nand U29104 (N_29104,N_28792,N_28810);
or U29105 (N_29105,N_28871,N_28989);
nand U29106 (N_29106,N_28783,N_28791);
xnor U29107 (N_29107,N_28811,N_28965);
or U29108 (N_29108,N_28785,N_28879);
or U29109 (N_29109,N_28761,N_28835);
and U29110 (N_29110,N_28795,N_28764);
nor U29111 (N_29111,N_28919,N_28895);
or U29112 (N_29112,N_28885,N_28926);
xor U29113 (N_29113,N_28789,N_28941);
or U29114 (N_29114,N_28875,N_28836);
and U29115 (N_29115,N_28975,N_28826);
nor U29116 (N_29116,N_28819,N_28945);
and U29117 (N_29117,N_28843,N_28853);
and U29118 (N_29118,N_28877,N_28774);
nor U29119 (N_29119,N_28949,N_28813);
or U29120 (N_29120,N_28874,N_28887);
nand U29121 (N_29121,N_28865,N_28905);
and U29122 (N_29122,N_28825,N_28936);
xnor U29123 (N_29123,N_28846,N_28790);
nor U29124 (N_29124,N_28839,N_28931);
xnor U29125 (N_29125,N_28877,N_28925);
or U29126 (N_29126,N_28979,N_28981);
or U29127 (N_29127,N_28775,N_28820);
nor U29128 (N_29128,N_28757,N_28909);
nor U29129 (N_29129,N_28877,N_28762);
nand U29130 (N_29130,N_28980,N_28908);
or U29131 (N_29131,N_28785,N_28893);
nor U29132 (N_29132,N_28949,N_28866);
nor U29133 (N_29133,N_28983,N_28982);
or U29134 (N_29134,N_28937,N_28796);
and U29135 (N_29135,N_28756,N_28881);
xnor U29136 (N_29136,N_28800,N_28993);
nor U29137 (N_29137,N_28927,N_28788);
xnor U29138 (N_29138,N_28882,N_28917);
nor U29139 (N_29139,N_28773,N_28864);
and U29140 (N_29140,N_28855,N_28829);
xor U29141 (N_29141,N_28803,N_28755);
xor U29142 (N_29142,N_28989,N_28819);
xnor U29143 (N_29143,N_28782,N_28976);
or U29144 (N_29144,N_28880,N_28958);
and U29145 (N_29145,N_28866,N_28940);
nand U29146 (N_29146,N_28776,N_28859);
xor U29147 (N_29147,N_28827,N_28989);
xnor U29148 (N_29148,N_28767,N_28971);
nor U29149 (N_29149,N_28766,N_28834);
nand U29150 (N_29150,N_28859,N_28971);
xnor U29151 (N_29151,N_28751,N_28959);
nand U29152 (N_29152,N_28790,N_28809);
nor U29153 (N_29153,N_28754,N_28954);
nand U29154 (N_29154,N_28901,N_28784);
and U29155 (N_29155,N_28871,N_28996);
nand U29156 (N_29156,N_28930,N_28839);
nor U29157 (N_29157,N_28915,N_28925);
xnor U29158 (N_29158,N_28906,N_28754);
and U29159 (N_29159,N_28913,N_28929);
xnor U29160 (N_29160,N_28867,N_28974);
and U29161 (N_29161,N_28896,N_28787);
and U29162 (N_29162,N_28781,N_28913);
or U29163 (N_29163,N_28864,N_28877);
nand U29164 (N_29164,N_28898,N_28996);
or U29165 (N_29165,N_28820,N_28977);
or U29166 (N_29166,N_28954,N_28819);
nor U29167 (N_29167,N_28911,N_28879);
or U29168 (N_29168,N_28906,N_28985);
or U29169 (N_29169,N_28991,N_28795);
nor U29170 (N_29170,N_28954,N_28844);
nand U29171 (N_29171,N_28833,N_28966);
nor U29172 (N_29172,N_28923,N_28914);
and U29173 (N_29173,N_28894,N_28983);
xor U29174 (N_29174,N_28997,N_28985);
nand U29175 (N_29175,N_28863,N_28815);
nor U29176 (N_29176,N_28990,N_28778);
and U29177 (N_29177,N_28992,N_28769);
and U29178 (N_29178,N_28852,N_28856);
nand U29179 (N_29179,N_28961,N_28958);
xor U29180 (N_29180,N_28885,N_28897);
or U29181 (N_29181,N_28870,N_28808);
xor U29182 (N_29182,N_28926,N_28894);
or U29183 (N_29183,N_28945,N_28809);
or U29184 (N_29184,N_28993,N_28844);
and U29185 (N_29185,N_28835,N_28910);
or U29186 (N_29186,N_28893,N_28973);
or U29187 (N_29187,N_28945,N_28889);
nand U29188 (N_29188,N_28906,N_28934);
nand U29189 (N_29189,N_28929,N_28828);
and U29190 (N_29190,N_28754,N_28815);
and U29191 (N_29191,N_28948,N_28776);
xor U29192 (N_29192,N_28886,N_28918);
and U29193 (N_29193,N_28826,N_28869);
or U29194 (N_29194,N_28765,N_28890);
nor U29195 (N_29195,N_28811,N_28891);
xnor U29196 (N_29196,N_28831,N_28967);
nor U29197 (N_29197,N_28970,N_28994);
nor U29198 (N_29198,N_28937,N_28847);
xnor U29199 (N_29199,N_28972,N_28926);
and U29200 (N_29200,N_28968,N_28784);
and U29201 (N_29201,N_28825,N_28868);
xnor U29202 (N_29202,N_28911,N_28811);
nor U29203 (N_29203,N_28978,N_28959);
and U29204 (N_29204,N_28903,N_28823);
and U29205 (N_29205,N_28948,N_28830);
or U29206 (N_29206,N_28942,N_28902);
nand U29207 (N_29207,N_28844,N_28931);
nand U29208 (N_29208,N_28785,N_28951);
nand U29209 (N_29209,N_28776,N_28830);
or U29210 (N_29210,N_28926,N_28830);
or U29211 (N_29211,N_28992,N_28935);
and U29212 (N_29212,N_28982,N_28781);
nand U29213 (N_29213,N_28983,N_28849);
nand U29214 (N_29214,N_28910,N_28926);
or U29215 (N_29215,N_28913,N_28895);
or U29216 (N_29216,N_28904,N_28760);
nor U29217 (N_29217,N_28755,N_28857);
nor U29218 (N_29218,N_28819,N_28839);
nand U29219 (N_29219,N_28830,N_28853);
nor U29220 (N_29220,N_28842,N_28786);
nor U29221 (N_29221,N_28969,N_28986);
nor U29222 (N_29222,N_28837,N_28967);
or U29223 (N_29223,N_28820,N_28915);
nand U29224 (N_29224,N_28912,N_28914);
nand U29225 (N_29225,N_28890,N_28944);
and U29226 (N_29226,N_28839,N_28750);
nand U29227 (N_29227,N_28804,N_28832);
or U29228 (N_29228,N_28892,N_28881);
or U29229 (N_29229,N_28839,N_28929);
xor U29230 (N_29230,N_28927,N_28829);
xnor U29231 (N_29231,N_28962,N_28813);
xor U29232 (N_29232,N_28773,N_28777);
or U29233 (N_29233,N_28780,N_28869);
or U29234 (N_29234,N_28848,N_28990);
nor U29235 (N_29235,N_28816,N_28890);
xnor U29236 (N_29236,N_28771,N_28829);
and U29237 (N_29237,N_28956,N_28841);
nor U29238 (N_29238,N_28774,N_28913);
xnor U29239 (N_29239,N_28806,N_28953);
and U29240 (N_29240,N_28985,N_28768);
or U29241 (N_29241,N_28839,N_28832);
xor U29242 (N_29242,N_28863,N_28823);
nor U29243 (N_29243,N_28774,N_28970);
nand U29244 (N_29244,N_28758,N_28843);
or U29245 (N_29245,N_28821,N_28941);
or U29246 (N_29246,N_28778,N_28941);
and U29247 (N_29247,N_28966,N_28895);
nand U29248 (N_29248,N_28907,N_28854);
and U29249 (N_29249,N_28770,N_28976);
or U29250 (N_29250,N_29072,N_29137);
and U29251 (N_29251,N_29138,N_29199);
and U29252 (N_29252,N_29140,N_29102);
and U29253 (N_29253,N_29161,N_29209);
or U29254 (N_29254,N_29083,N_29112);
nor U29255 (N_29255,N_29003,N_29187);
or U29256 (N_29256,N_29103,N_29226);
xor U29257 (N_29257,N_29213,N_29149);
and U29258 (N_29258,N_29046,N_29135);
xor U29259 (N_29259,N_29236,N_29203);
xor U29260 (N_29260,N_29095,N_29120);
xnor U29261 (N_29261,N_29008,N_29181);
nand U29262 (N_29262,N_29192,N_29228);
xnor U29263 (N_29263,N_29150,N_29220);
xnor U29264 (N_29264,N_29234,N_29133);
or U29265 (N_29265,N_29128,N_29110);
nand U29266 (N_29266,N_29195,N_29009);
or U29267 (N_29267,N_29170,N_29020);
and U29268 (N_29268,N_29247,N_29074);
or U29269 (N_29269,N_29145,N_29023);
or U29270 (N_29270,N_29036,N_29176);
nand U29271 (N_29271,N_29058,N_29179);
xor U29272 (N_29272,N_29193,N_29249);
nand U29273 (N_29273,N_29001,N_29157);
or U29274 (N_29274,N_29092,N_29132);
nand U29275 (N_29275,N_29186,N_29017);
xnor U29276 (N_29276,N_29109,N_29224);
or U29277 (N_29277,N_29211,N_29159);
nor U29278 (N_29278,N_29002,N_29073);
or U29279 (N_29279,N_29094,N_29107);
and U29280 (N_29280,N_29118,N_29049);
nand U29281 (N_29281,N_29246,N_29063);
nor U29282 (N_29282,N_29231,N_29087);
or U29283 (N_29283,N_29027,N_29096);
and U29284 (N_29284,N_29196,N_29183);
nand U29285 (N_29285,N_29204,N_29162);
xnor U29286 (N_29286,N_29153,N_29142);
or U29287 (N_29287,N_29164,N_29067);
or U29288 (N_29288,N_29218,N_29048);
nand U29289 (N_29289,N_29194,N_29050);
nor U29290 (N_29290,N_29034,N_29075);
nand U29291 (N_29291,N_29175,N_29028);
xnor U29292 (N_29292,N_29114,N_29007);
nor U29293 (N_29293,N_29084,N_29184);
or U29294 (N_29294,N_29033,N_29171);
nand U29295 (N_29295,N_29156,N_29198);
nand U29296 (N_29296,N_29155,N_29089);
or U29297 (N_29297,N_29006,N_29031);
or U29298 (N_29298,N_29071,N_29214);
and U29299 (N_29299,N_29223,N_29116);
nand U29300 (N_29300,N_29151,N_29126);
xnor U29301 (N_29301,N_29051,N_29052);
xor U29302 (N_29302,N_29243,N_29113);
xnor U29303 (N_29303,N_29127,N_29066);
nor U29304 (N_29304,N_29158,N_29222);
xor U29305 (N_29305,N_29144,N_29022);
nand U29306 (N_29306,N_29099,N_29202);
and U29307 (N_29307,N_29177,N_29160);
and U29308 (N_29308,N_29111,N_29244);
nand U29309 (N_29309,N_29121,N_29038);
nor U29310 (N_29310,N_29143,N_29225);
nand U29311 (N_29311,N_29069,N_29201);
nand U29312 (N_29312,N_29131,N_29217);
xnor U29313 (N_29313,N_29188,N_29080);
nand U29314 (N_29314,N_29189,N_29108);
nor U29315 (N_29315,N_29129,N_29146);
and U29316 (N_29316,N_29206,N_29029);
xnor U29317 (N_29317,N_29185,N_29011);
xnor U29318 (N_29318,N_29154,N_29088);
nand U29319 (N_29319,N_29212,N_29235);
and U29320 (N_29320,N_29064,N_29014);
nor U29321 (N_29321,N_29115,N_29056);
nor U29322 (N_29322,N_29182,N_29173);
xnor U29323 (N_29323,N_29062,N_29141);
xnor U29324 (N_29324,N_29136,N_29041);
and U29325 (N_29325,N_29172,N_29123);
or U29326 (N_29326,N_29237,N_29169);
nand U29327 (N_29327,N_29000,N_29122);
xnor U29328 (N_29328,N_29208,N_29079);
xor U29329 (N_29329,N_29037,N_29091);
and U29330 (N_29330,N_29019,N_29012);
xnor U29331 (N_29331,N_29104,N_29215);
nand U29332 (N_29332,N_29085,N_29016);
or U29333 (N_29333,N_29242,N_29239);
nand U29334 (N_29334,N_29004,N_29054);
nand U29335 (N_29335,N_29018,N_29174);
nor U29336 (N_29336,N_29232,N_29119);
nand U29337 (N_29337,N_29229,N_29125);
xor U29338 (N_29338,N_29100,N_29178);
and U29339 (N_29339,N_29032,N_29191);
nand U29340 (N_29340,N_29026,N_29039);
xnor U29341 (N_29341,N_29055,N_29227);
nor U29342 (N_29342,N_29238,N_29165);
or U29343 (N_29343,N_29190,N_29043);
xor U29344 (N_29344,N_29010,N_29219);
and U29345 (N_29345,N_29124,N_29082);
nor U29346 (N_29346,N_29086,N_29106);
xnor U29347 (N_29347,N_29076,N_29248);
nand U29348 (N_29348,N_29059,N_29139);
nor U29349 (N_29349,N_29167,N_29025);
nand U29350 (N_29350,N_29180,N_29030);
and U29351 (N_29351,N_29068,N_29134);
and U29352 (N_29352,N_29047,N_29035);
nand U29353 (N_29353,N_29221,N_29101);
or U29354 (N_29354,N_29207,N_29245);
or U29355 (N_29355,N_29065,N_29152);
nor U29356 (N_29356,N_29210,N_29057);
nor U29357 (N_29357,N_29015,N_29044);
and U29358 (N_29358,N_29078,N_29205);
nor U29359 (N_29359,N_29105,N_29166);
xor U29360 (N_29360,N_29053,N_29024);
or U29361 (N_29361,N_29168,N_29240);
and U29362 (N_29362,N_29077,N_29097);
and U29363 (N_29363,N_29061,N_29090);
or U29364 (N_29364,N_29148,N_29042);
nand U29365 (N_29365,N_29070,N_29013);
and U29366 (N_29366,N_29147,N_29045);
and U29367 (N_29367,N_29098,N_29216);
and U29368 (N_29368,N_29081,N_29230);
xor U29369 (N_29369,N_29117,N_29005);
nor U29370 (N_29370,N_29130,N_29163);
or U29371 (N_29371,N_29093,N_29197);
or U29372 (N_29372,N_29241,N_29021);
nor U29373 (N_29373,N_29060,N_29040);
and U29374 (N_29374,N_29200,N_29233);
and U29375 (N_29375,N_29141,N_29068);
nand U29376 (N_29376,N_29060,N_29144);
xnor U29377 (N_29377,N_29222,N_29165);
nor U29378 (N_29378,N_29090,N_29160);
or U29379 (N_29379,N_29133,N_29095);
nor U29380 (N_29380,N_29004,N_29022);
nand U29381 (N_29381,N_29225,N_29088);
nand U29382 (N_29382,N_29092,N_29002);
nor U29383 (N_29383,N_29048,N_29029);
or U29384 (N_29384,N_29236,N_29212);
nor U29385 (N_29385,N_29060,N_29237);
nand U29386 (N_29386,N_29020,N_29172);
xnor U29387 (N_29387,N_29128,N_29017);
and U29388 (N_29388,N_29120,N_29171);
xor U29389 (N_29389,N_29142,N_29075);
nor U29390 (N_29390,N_29108,N_29039);
or U29391 (N_29391,N_29223,N_29233);
or U29392 (N_29392,N_29046,N_29195);
and U29393 (N_29393,N_29214,N_29086);
or U29394 (N_29394,N_29038,N_29009);
nand U29395 (N_29395,N_29098,N_29213);
nor U29396 (N_29396,N_29162,N_29083);
nor U29397 (N_29397,N_29227,N_29102);
xor U29398 (N_29398,N_29147,N_29121);
or U29399 (N_29399,N_29073,N_29072);
nor U29400 (N_29400,N_29063,N_29192);
and U29401 (N_29401,N_29078,N_29143);
nor U29402 (N_29402,N_29102,N_29016);
or U29403 (N_29403,N_29077,N_29095);
or U29404 (N_29404,N_29152,N_29122);
nor U29405 (N_29405,N_29037,N_29056);
and U29406 (N_29406,N_29114,N_29154);
and U29407 (N_29407,N_29126,N_29195);
nor U29408 (N_29408,N_29112,N_29027);
nand U29409 (N_29409,N_29071,N_29197);
xnor U29410 (N_29410,N_29195,N_29120);
nand U29411 (N_29411,N_29081,N_29091);
nor U29412 (N_29412,N_29192,N_29013);
and U29413 (N_29413,N_29111,N_29086);
xor U29414 (N_29414,N_29060,N_29200);
nand U29415 (N_29415,N_29047,N_29097);
or U29416 (N_29416,N_29238,N_29214);
and U29417 (N_29417,N_29143,N_29192);
xnor U29418 (N_29418,N_29169,N_29155);
nor U29419 (N_29419,N_29042,N_29001);
or U29420 (N_29420,N_29127,N_29162);
nand U29421 (N_29421,N_29106,N_29006);
nor U29422 (N_29422,N_29162,N_29199);
xor U29423 (N_29423,N_29206,N_29130);
xnor U29424 (N_29424,N_29131,N_29241);
nand U29425 (N_29425,N_29204,N_29167);
xnor U29426 (N_29426,N_29101,N_29166);
or U29427 (N_29427,N_29204,N_29097);
nor U29428 (N_29428,N_29212,N_29003);
xnor U29429 (N_29429,N_29109,N_29036);
nand U29430 (N_29430,N_29076,N_29224);
and U29431 (N_29431,N_29091,N_29125);
or U29432 (N_29432,N_29126,N_29208);
nor U29433 (N_29433,N_29043,N_29169);
or U29434 (N_29434,N_29089,N_29184);
xor U29435 (N_29435,N_29012,N_29008);
and U29436 (N_29436,N_29195,N_29131);
xnor U29437 (N_29437,N_29096,N_29005);
xor U29438 (N_29438,N_29017,N_29075);
xnor U29439 (N_29439,N_29228,N_29034);
or U29440 (N_29440,N_29102,N_29069);
nor U29441 (N_29441,N_29244,N_29083);
xnor U29442 (N_29442,N_29219,N_29164);
nor U29443 (N_29443,N_29097,N_29057);
xnor U29444 (N_29444,N_29107,N_29059);
nor U29445 (N_29445,N_29096,N_29022);
nand U29446 (N_29446,N_29006,N_29199);
xor U29447 (N_29447,N_29156,N_29016);
and U29448 (N_29448,N_29061,N_29180);
and U29449 (N_29449,N_29089,N_29137);
xor U29450 (N_29450,N_29051,N_29244);
nand U29451 (N_29451,N_29178,N_29098);
or U29452 (N_29452,N_29041,N_29123);
xnor U29453 (N_29453,N_29240,N_29236);
or U29454 (N_29454,N_29144,N_29108);
or U29455 (N_29455,N_29074,N_29202);
xnor U29456 (N_29456,N_29074,N_29194);
or U29457 (N_29457,N_29050,N_29090);
or U29458 (N_29458,N_29215,N_29205);
nand U29459 (N_29459,N_29031,N_29216);
nor U29460 (N_29460,N_29041,N_29208);
and U29461 (N_29461,N_29001,N_29028);
xor U29462 (N_29462,N_29003,N_29174);
nor U29463 (N_29463,N_29199,N_29024);
nor U29464 (N_29464,N_29199,N_29100);
nand U29465 (N_29465,N_29079,N_29249);
and U29466 (N_29466,N_29196,N_29233);
or U29467 (N_29467,N_29209,N_29177);
xor U29468 (N_29468,N_29024,N_29183);
nand U29469 (N_29469,N_29155,N_29158);
nor U29470 (N_29470,N_29215,N_29030);
xnor U29471 (N_29471,N_29194,N_29062);
xnor U29472 (N_29472,N_29249,N_29039);
nand U29473 (N_29473,N_29118,N_29122);
and U29474 (N_29474,N_29133,N_29083);
nand U29475 (N_29475,N_29118,N_29181);
nand U29476 (N_29476,N_29049,N_29236);
xnor U29477 (N_29477,N_29050,N_29144);
nor U29478 (N_29478,N_29233,N_29139);
or U29479 (N_29479,N_29205,N_29108);
nor U29480 (N_29480,N_29190,N_29084);
or U29481 (N_29481,N_29043,N_29056);
or U29482 (N_29482,N_29130,N_29121);
and U29483 (N_29483,N_29150,N_29131);
nor U29484 (N_29484,N_29235,N_29030);
or U29485 (N_29485,N_29178,N_29123);
nand U29486 (N_29486,N_29127,N_29216);
and U29487 (N_29487,N_29054,N_29114);
xnor U29488 (N_29488,N_29235,N_29070);
nor U29489 (N_29489,N_29160,N_29202);
nand U29490 (N_29490,N_29011,N_29039);
or U29491 (N_29491,N_29068,N_29095);
nor U29492 (N_29492,N_29208,N_29210);
nand U29493 (N_29493,N_29027,N_29243);
nand U29494 (N_29494,N_29214,N_29151);
nand U29495 (N_29495,N_29089,N_29203);
nand U29496 (N_29496,N_29073,N_29141);
and U29497 (N_29497,N_29245,N_29227);
nor U29498 (N_29498,N_29132,N_29070);
xor U29499 (N_29499,N_29134,N_29237);
and U29500 (N_29500,N_29347,N_29441);
nor U29501 (N_29501,N_29410,N_29279);
or U29502 (N_29502,N_29264,N_29321);
nand U29503 (N_29503,N_29397,N_29260);
and U29504 (N_29504,N_29431,N_29409);
nand U29505 (N_29505,N_29391,N_29303);
and U29506 (N_29506,N_29446,N_29459);
or U29507 (N_29507,N_29407,N_29285);
or U29508 (N_29508,N_29396,N_29301);
nand U29509 (N_29509,N_29394,N_29402);
or U29510 (N_29510,N_29480,N_29349);
nor U29511 (N_29511,N_29418,N_29448);
nor U29512 (N_29512,N_29414,N_29469);
nand U29513 (N_29513,N_29430,N_29463);
or U29514 (N_29514,N_29284,N_29287);
xnor U29515 (N_29515,N_29438,N_29375);
nand U29516 (N_29516,N_29497,N_29356);
xnor U29517 (N_29517,N_29283,N_29265);
nor U29518 (N_29518,N_29316,N_29363);
or U29519 (N_29519,N_29372,N_29432);
nor U29520 (N_29520,N_29352,N_29496);
xor U29521 (N_29521,N_29368,N_29381);
and U29522 (N_29522,N_29378,N_29401);
and U29523 (N_29523,N_29434,N_29296);
nor U29524 (N_29524,N_29299,N_29488);
and U29525 (N_29525,N_29289,N_29456);
or U29526 (N_29526,N_29481,N_29393);
and U29527 (N_29527,N_29346,N_29433);
or U29528 (N_29528,N_29293,N_29367);
and U29529 (N_29529,N_29436,N_29404);
or U29530 (N_29530,N_29455,N_29440);
xnor U29531 (N_29531,N_29315,N_29450);
nor U29532 (N_29532,N_29318,N_29443);
and U29533 (N_29533,N_29335,N_29261);
and U29534 (N_29534,N_29345,N_29474);
nand U29535 (N_29535,N_29462,N_29408);
nand U29536 (N_29536,N_29442,N_29251);
and U29537 (N_29537,N_29371,N_29483);
xor U29538 (N_29538,N_29473,N_29376);
nor U29539 (N_29539,N_29353,N_29498);
or U29540 (N_29540,N_29340,N_29451);
xor U29541 (N_29541,N_29277,N_29460);
nor U29542 (N_29542,N_29270,N_29271);
xnor U29543 (N_29543,N_29332,N_29317);
xor U29544 (N_29544,N_29373,N_29281);
and U29545 (N_29545,N_29382,N_29314);
and U29546 (N_29546,N_29257,N_29383);
nor U29547 (N_29547,N_29369,N_29252);
nand U29548 (N_29548,N_29364,N_29411);
and U29549 (N_29549,N_29419,N_29406);
nor U29550 (N_29550,N_29254,N_29491);
nand U29551 (N_29551,N_29256,N_29266);
nor U29552 (N_29552,N_29466,N_29415);
nor U29553 (N_29553,N_29494,N_29472);
or U29554 (N_29554,N_29297,N_29392);
nand U29555 (N_29555,N_29422,N_29398);
or U29556 (N_29556,N_29272,N_29477);
and U29557 (N_29557,N_29276,N_29290);
nor U29558 (N_29558,N_29490,N_29333);
or U29559 (N_29559,N_29311,N_29467);
nor U29560 (N_29560,N_29395,N_29275);
nor U29561 (N_29561,N_29478,N_29258);
and U29562 (N_29562,N_29319,N_29457);
xor U29563 (N_29563,N_29310,N_29278);
nor U29564 (N_29564,N_29471,N_29428);
nor U29565 (N_29565,N_29309,N_29482);
nor U29566 (N_29566,N_29294,N_29361);
xor U29567 (N_29567,N_29464,N_29334);
nor U29568 (N_29568,N_29273,N_29322);
or U29569 (N_29569,N_29458,N_29348);
nor U29570 (N_29570,N_29427,N_29326);
nor U29571 (N_29571,N_29304,N_29313);
xnor U29572 (N_29572,N_29403,N_29475);
nand U29573 (N_29573,N_29262,N_29250);
or U29574 (N_29574,N_29307,N_29439);
nand U29575 (N_29575,N_29465,N_29413);
nand U29576 (N_29576,N_29339,N_29389);
or U29577 (N_29577,N_29416,N_29417);
xor U29578 (N_29578,N_29486,N_29282);
or U29579 (N_29579,N_29302,N_29385);
or U29580 (N_29580,N_29424,N_29253);
and U29581 (N_29581,N_29390,N_29343);
or U29582 (N_29582,N_29336,N_29429);
nand U29583 (N_29583,N_29421,N_29337);
nand U29584 (N_29584,N_29495,N_29454);
and U29585 (N_29585,N_29341,N_29298);
and U29586 (N_29586,N_29476,N_29329);
and U29587 (N_29587,N_29362,N_29485);
or U29588 (N_29588,N_29445,N_29499);
xor U29589 (N_29589,N_29342,N_29288);
xnor U29590 (N_29590,N_29399,N_29327);
nor U29591 (N_29591,N_29305,N_29366);
and U29592 (N_29592,N_29453,N_29461);
or U29593 (N_29593,N_29295,N_29350);
or U29594 (N_29594,N_29374,N_29357);
or U29595 (N_29595,N_29330,N_29358);
xor U29596 (N_29596,N_29312,N_29420);
or U29597 (N_29597,N_29386,N_29405);
nand U29598 (N_29598,N_29351,N_29355);
xnor U29599 (N_29599,N_29359,N_29365);
and U29600 (N_29600,N_29425,N_29400);
nand U29601 (N_29601,N_29268,N_29447);
xor U29602 (N_29602,N_29344,N_29324);
and U29603 (N_29603,N_29377,N_29479);
or U29604 (N_29604,N_29267,N_29323);
xnor U29605 (N_29605,N_29489,N_29331);
or U29606 (N_29606,N_29387,N_29308);
nor U29607 (N_29607,N_29484,N_29370);
nor U29608 (N_29608,N_29380,N_29452);
xor U29609 (N_29609,N_29360,N_29437);
xor U29610 (N_29610,N_29280,N_29354);
nand U29611 (N_29611,N_29470,N_29468);
nor U29612 (N_29612,N_29255,N_29426);
xor U29613 (N_29613,N_29259,N_29291);
nand U29614 (N_29614,N_29263,N_29423);
nor U29615 (N_29615,N_29292,N_29300);
and U29616 (N_29616,N_29320,N_29493);
nor U29617 (N_29617,N_29449,N_29412);
xnor U29618 (N_29618,N_29325,N_29435);
and U29619 (N_29619,N_29487,N_29328);
nor U29620 (N_29620,N_29492,N_29384);
and U29621 (N_29621,N_29306,N_29388);
nand U29622 (N_29622,N_29286,N_29444);
nand U29623 (N_29623,N_29338,N_29274);
nand U29624 (N_29624,N_29269,N_29379);
or U29625 (N_29625,N_29449,N_29390);
nor U29626 (N_29626,N_29273,N_29444);
and U29627 (N_29627,N_29268,N_29492);
and U29628 (N_29628,N_29287,N_29322);
or U29629 (N_29629,N_29404,N_29368);
or U29630 (N_29630,N_29287,N_29446);
and U29631 (N_29631,N_29409,N_29327);
and U29632 (N_29632,N_29380,N_29485);
nand U29633 (N_29633,N_29396,N_29338);
nor U29634 (N_29634,N_29411,N_29373);
and U29635 (N_29635,N_29395,N_29414);
nor U29636 (N_29636,N_29460,N_29441);
xnor U29637 (N_29637,N_29386,N_29439);
nand U29638 (N_29638,N_29471,N_29452);
nand U29639 (N_29639,N_29454,N_29326);
xor U29640 (N_29640,N_29262,N_29311);
nand U29641 (N_29641,N_29482,N_29285);
nor U29642 (N_29642,N_29446,N_29468);
nor U29643 (N_29643,N_29270,N_29396);
xnor U29644 (N_29644,N_29290,N_29339);
xnor U29645 (N_29645,N_29421,N_29474);
nor U29646 (N_29646,N_29434,N_29300);
nand U29647 (N_29647,N_29275,N_29326);
and U29648 (N_29648,N_29490,N_29296);
and U29649 (N_29649,N_29397,N_29270);
nand U29650 (N_29650,N_29358,N_29289);
or U29651 (N_29651,N_29478,N_29488);
nor U29652 (N_29652,N_29464,N_29372);
nand U29653 (N_29653,N_29307,N_29365);
nand U29654 (N_29654,N_29456,N_29313);
and U29655 (N_29655,N_29429,N_29288);
nor U29656 (N_29656,N_29433,N_29284);
nand U29657 (N_29657,N_29348,N_29432);
and U29658 (N_29658,N_29381,N_29282);
xor U29659 (N_29659,N_29407,N_29358);
or U29660 (N_29660,N_29347,N_29275);
nand U29661 (N_29661,N_29479,N_29422);
nor U29662 (N_29662,N_29489,N_29314);
and U29663 (N_29663,N_29276,N_29403);
or U29664 (N_29664,N_29413,N_29337);
and U29665 (N_29665,N_29323,N_29378);
and U29666 (N_29666,N_29264,N_29361);
nand U29667 (N_29667,N_29346,N_29471);
nand U29668 (N_29668,N_29434,N_29382);
nor U29669 (N_29669,N_29332,N_29439);
nor U29670 (N_29670,N_29466,N_29279);
and U29671 (N_29671,N_29452,N_29275);
nor U29672 (N_29672,N_29320,N_29494);
xnor U29673 (N_29673,N_29466,N_29473);
nor U29674 (N_29674,N_29398,N_29366);
and U29675 (N_29675,N_29337,N_29294);
or U29676 (N_29676,N_29493,N_29423);
and U29677 (N_29677,N_29299,N_29330);
or U29678 (N_29678,N_29479,N_29260);
or U29679 (N_29679,N_29430,N_29494);
xnor U29680 (N_29680,N_29419,N_29314);
and U29681 (N_29681,N_29397,N_29259);
nand U29682 (N_29682,N_29261,N_29449);
and U29683 (N_29683,N_29361,N_29317);
or U29684 (N_29684,N_29347,N_29418);
nor U29685 (N_29685,N_29473,N_29355);
or U29686 (N_29686,N_29358,N_29309);
xnor U29687 (N_29687,N_29448,N_29345);
xor U29688 (N_29688,N_29439,N_29489);
nor U29689 (N_29689,N_29491,N_29365);
or U29690 (N_29690,N_29337,N_29443);
and U29691 (N_29691,N_29339,N_29334);
or U29692 (N_29692,N_29451,N_29463);
or U29693 (N_29693,N_29497,N_29390);
and U29694 (N_29694,N_29397,N_29468);
and U29695 (N_29695,N_29383,N_29326);
nor U29696 (N_29696,N_29482,N_29337);
and U29697 (N_29697,N_29269,N_29404);
nand U29698 (N_29698,N_29274,N_29442);
nor U29699 (N_29699,N_29453,N_29415);
nand U29700 (N_29700,N_29363,N_29310);
nand U29701 (N_29701,N_29307,N_29356);
xnor U29702 (N_29702,N_29295,N_29308);
xnor U29703 (N_29703,N_29377,N_29478);
xnor U29704 (N_29704,N_29386,N_29443);
or U29705 (N_29705,N_29459,N_29387);
or U29706 (N_29706,N_29285,N_29382);
and U29707 (N_29707,N_29438,N_29489);
or U29708 (N_29708,N_29291,N_29288);
xor U29709 (N_29709,N_29459,N_29467);
nand U29710 (N_29710,N_29493,N_29352);
xor U29711 (N_29711,N_29471,N_29349);
or U29712 (N_29712,N_29473,N_29454);
and U29713 (N_29713,N_29424,N_29399);
and U29714 (N_29714,N_29477,N_29372);
nor U29715 (N_29715,N_29354,N_29334);
or U29716 (N_29716,N_29484,N_29499);
xor U29717 (N_29717,N_29299,N_29499);
nand U29718 (N_29718,N_29472,N_29362);
xor U29719 (N_29719,N_29335,N_29371);
and U29720 (N_29720,N_29271,N_29400);
and U29721 (N_29721,N_29275,N_29457);
nor U29722 (N_29722,N_29438,N_29433);
nor U29723 (N_29723,N_29446,N_29457);
nor U29724 (N_29724,N_29302,N_29391);
nor U29725 (N_29725,N_29357,N_29345);
or U29726 (N_29726,N_29255,N_29347);
or U29727 (N_29727,N_29393,N_29374);
or U29728 (N_29728,N_29442,N_29362);
xor U29729 (N_29729,N_29398,N_29424);
or U29730 (N_29730,N_29387,N_29342);
nor U29731 (N_29731,N_29363,N_29389);
or U29732 (N_29732,N_29450,N_29329);
nor U29733 (N_29733,N_29493,N_29250);
nor U29734 (N_29734,N_29327,N_29377);
nor U29735 (N_29735,N_29404,N_29310);
or U29736 (N_29736,N_29265,N_29454);
xnor U29737 (N_29737,N_29328,N_29291);
nand U29738 (N_29738,N_29440,N_29431);
nand U29739 (N_29739,N_29304,N_29411);
nand U29740 (N_29740,N_29375,N_29415);
and U29741 (N_29741,N_29281,N_29334);
nor U29742 (N_29742,N_29347,N_29352);
xnor U29743 (N_29743,N_29307,N_29260);
xor U29744 (N_29744,N_29298,N_29306);
nand U29745 (N_29745,N_29252,N_29432);
xor U29746 (N_29746,N_29365,N_29456);
xor U29747 (N_29747,N_29442,N_29322);
and U29748 (N_29748,N_29365,N_29384);
nor U29749 (N_29749,N_29488,N_29425);
nand U29750 (N_29750,N_29747,N_29643);
and U29751 (N_29751,N_29624,N_29616);
nand U29752 (N_29752,N_29519,N_29592);
and U29753 (N_29753,N_29546,N_29650);
xnor U29754 (N_29754,N_29608,N_29701);
nor U29755 (N_29755,N_29500,N_29695);
or U29756 (N_29756,N_29518,N_29594);
xor U29757 (N_29757,N_29567,N_29683);
nor U29758 (N_29758,N_29628,N_29692);
and U29759 (N_29759,N_29606,N_29506);
and U29760 (N_29760,N_29671,N_29525);
xnor U29761 (N_29761,N_29723,N_29618);
xnor U29762 (N_29762,N_29741,N_29609);
and U29763 (N_29763,N_29742,N_29548);
xnor U29764 (N_29764,N_29542,N_29703);
xnor U29765 (N_29765,N_29731,N_29659);
or U29766 (N_29766,N_29673,N_29635);
xor U29767 (N_29767,N_29712,N_29543);
or U29768 (N_29768,N_29709,N_29558);
or U29769 (N_29769,N_29682,N_29740);
and U29770 (N_29770,N_29666,N_29721);
nand U29771 (N_29771,N_29585,N_29621);
nor U29772 (N_29772,N_29664,N_29602);
or U29773 (N_29773,N_29568,N_29647);
nand U29774 (N_29774,N_29582,N_29502);
or U29775 (N_29775,N_29719,N_29679);
or U29776 (N_29776,N_29577,N_29575);
nor U29777 (N_29777,N_29738,N_29541);
nor U29778 (N_29778,N_29644,N_29574);
or U29779 (N_29779,N_29601,N_29586);
and U29780 (N_29780,N_29604,N_29711);
or U29781 (N_29781,N_29564,N_29596);
and U29782 (N_29782,N_29615,N_29654);
xnor U29783 (N_29783,N_29524,N_29613);
xnor U29784 (N_29784,N_29539,N_29600);
and U29785 (N_29785,N_29674,N_29708);
xor U29786 (N_29786,N_29545,N_29736);
xor U29787 (N_29787,N_29552,N_29579);
and U29788 (N_29788,N_29717,N_29680);
and U29789 (N_29789,N_29704,N_29535);
nand U29790 (N_29790,N_29630,N_29527);
nor U29791 (N_29791,N_29528,N_29540);
or U29792 (N_29792,N_29713,N_29663);
or U29793 (N_29793,N_29515,N_29556);
or U29794 (N_29794,N_29684,N_29728);
nand U29795 (N_29795,N_29587,N_29634);
nor U29796 (N_29796,N_29660,N_29639);
nor U29797 (N_29797,N_29529,N_29732);
nand U29798 (N_29798,N_29531,N_29536);
nand U29799 (N_29799,N_29633,N_29503);
or U29800 (N_29800,N_29559,N_29672);
xor U29801 (N_29801,N_29589,N_29566);
nand U29802 (N_29802,N_29593,N_29676);
and U29803 (N_29803,N_29668,N_29642);
nor U29804 (N_29804,N_29510,N_29513);
nand U29805 (N_29805,N_29538,N_29534);
nor U29806 (N_29806,N_29549,N_29745);
nor U29807 (N_29807,N_29658,N_29572);
xor U29808 (N_29808,N_29688,N_29565);
and U29809 (N_29809,N_29746,N_29521);
nor U29810 (N_29810,N_29687,N_29509);
xor U29811 (N_29811,N_29661,N_29652);
and U29812 (N_29812,N_29699,N_29649);
or U29813 (N_29813,N_29669,N_29690);
and U29814 (N_29814,N_29603,N_29610);
nor U29815 (N_29815,N_29743,N_29675);
nand U29816 (N_29816,N_29697,N_29581);
and U29817 (N_29817,N_29599,N_29700);
nor U29818 (N_29818,N_29722,N_29627);
or U29819 (N_29819,N_29710,N_29707);
nand U29820 (N_29820,N_29507,N_29748);
xor U29821 (N_29821,N_29694,N_29725);
xnor U29822 (N_29822,N_29514,N_29641);
xor U29823 (N_29823,N_29526,N_29504);
or U29824 (N_29824,N_29714,N_29590);
and U29825 (N_29825,N_29583,N_29533);
xnor U29826 (N_29826,N_29648,N_29667);
and U29827 (N_29827,N_29677,N_29622);
nand U29828 (N_29828,N_29544,N_29555);
nor U29829 (N_29829,N_29656,N_29576);
nor U29830 (N_29830,N_29715,N_29637);
nor U29831 (N_29831,N_29705,N_29595);
nand U29832 (N_29832,N_29691,N_29625);
nor U29833 (N_29833,N_29571,N_29569);
xor U29834 (N_29834,N_29580,N_29597);
and U29835 (N_29835,N_29720,N_29523);
nand U29836 (N_29836,N_29640,N_29716);
xor U29837 (N_29837,N_29584,N_29517);
or U29838 (N_29838,N_29665,N_29629);
nand U29839 (N_29839,N_29591,N_29520);
or U29840 (N_29840,N_29729,N_29578);
nand U29841 (N_29841,N_29638,N_29588);
xnor U29842 (N_29842,N_29550,N_29657);
xnor U29843 (N_29843,N_29607,N_29611);
and U29844 (N_29844,N_29557,N_29561);
xor U29845 (N_29845,N_29646,N_29718);
or U29846 (N_29846,N_29532,N_29653);
nor U29847 (N_29847,N_29511,N_29744);
nand U29848 (N_29848,N_29730,N_29733);
or U29849 (N_29849,N_29686,N_29547);
nor U29850 (N_29850,N_29560,N_29617);
or U29851 (N_29851,N_29614,N_29620);
or U29852 (N_29852,N_29670,N_29505);
xor U29853 (N_29853,N_29689,N_29573);
xor U29854 (N_29854,N_29554,N_29735);
nor U29855 (N_29855,N_29698,N_29706);
xnor U29856 (N_29856,N_29626,N_29512);
and U29857 (N_29857,N_29749,N_29655);
xor U29858 (N_29858,N_29662,N_29508);
or U29859 (N_29859,N_29632,N_29598);
and U29860 (N_29860,N_29734,N_29696);
nor U29861 (N_29861,N_29501,N_29737);
xnor U29862 (N_29862,N_29562,N_29563);
and U29863 (N_29863,N_29702,N_29530);
and U29864 (N_29864,N_29693,N_29551);
nor U29865 (N_29865,N_29726,N_29516);
nor U29866 (N_29866,N_29724,N_29651);
or U29867 (N_29867,N_29612,N_29681);
nand U29868 (N_29868,N_29605,N_29537);
nor U29869 (N_29869,N_29623,N_29522);
nor U29870 (N_29870,N_29619,N_29636);
nand U29871 (N_29871,N_29645,N_29570);
xnor U29872 (N_29872,N_29727,N_29739);
nor U29873 (N_29873,N_29678,N_29685);
nor U29874 (N_29874,N_29553,N_29631);
nor U29875 (N_29875,N_29631,N_29519);
or U29876 (N_29876,N_29691,N_29579);
nand U29877 (N_29877,N_29599,N_29639);
nand U29878 (N_29878,N_29506,N_29647);
nor U29879 (N_29879,N_29512,N_29586);
or U29880 (N_29880,N_29639,N_29573);
nand U29881 (N_29881,N_29708,N_29645);
or U29882 (N_29882,N_29726,N_29684);
nand U29883 (N_29883,N_29512,N_29676);
nand U29884 (N_29884,N_29699,N_29700);
nor U29885 (N_29885,N_29727,N_29686);
xnor U29886 (N_29886,N_29646,N_29721);
or U29887 (N_29887,N_29683,N_29559);
nor U29888 (N_29888,N_29568,N_29562);
or U29889 (N_29889,N_29564,N_29700);
or U29890 (N_29890,N_29583,N_29553);
or U29891 (N_29891,N_29608,N_29523);
nor U29892 (N_29892,N_29707,N_29618);
or U29893 (N_29893,N_29657,N_29717);
xor U29894 (N_29894,N_29688,N_29584);
and U29895 (N_29895,N_29583,N_29601);
nor U29896 (N_29896,N_29615,N_29556);
and U29897 (N_29897,N_29715,N_29699);
xnor U29898 (N_29898,N_29566,N_29513);
nor U29899 (N_29899,N_29561,N_29559);
nand U29900 (N_29900,N_29740,N_29666);
and U29901 (N_29901,N_29684,N_29531);
or U29902 (N_29902,N_29656,N_29589);
xnor U29903 (N_29903,N_29703,N_29604);
and U29904 (N_29904,N_29658,N_29651);
or U29905 (N_29905,N_29658,N_29655);
and U29906 (N_29906,N_29590,N_29671);
nor U29907 (N_29907,N_29631,N_29534);
nor U29908 (N_29908,N_29542,N_29593);
xor U29909 (N_29909,N_29734,N_29591);
and U29910 (N_29910,N_29501,N_29715);
and U29911 (N_29911,N_29709,N_29740);
or U29912 (N_29912,N_29529,N_29590);
or U29913 (N_29913,N_29554,N_29567);
or U29914 (N_29914,N_29654,N_29664);
and U29915 (N_29915,N_29674,N_29604);
nor U29916 (N_29916,N_29688,N_29569);
nand U29917 (N_29917,N_29529,N_29569);
or U29918 (N_29918,N_29604,N_29664);
and U29919 (N_29919,N_29742,N_29738);
nor U29920 (N_29920,N_29661,N_29749);
and U29921 (N_29921,N_29659,N_29500);
nand U29922 (N_29922,N_29521,N_29609);
nor U29923 (N_29923,N_29537,N_29691);
and U29924 (N_29924,N_29556,N_29612);
and U29925 (N_29925,N_29523,N_29684);
or U29926 (N_29926,N_29598,N_29634);
and U29927 (N_29927,N_29614,N_29505);
nor U29928 (N_29928,N_29693,N_29703);
or U29929 (N_29929,N_29655,N_29643);
nor U29930 (N_29930,N_29660,N_29589);
nor U29931 (N_29931,N_29697,N_29639);
nand U29932 (N_29932,N_29726,N_29567);
nor U29933 (N_29933,N_29720,N_29600);
nand U29934 (N_29934,N_29591,N_29575);
and U29935 (N_29935,N_29714,N_29690);
or U29936 (N_29936,N_29592,N_29564);
nand U29937 (N_29937,N_29712,N_29692);
and U29938 (N_29938,N_29685,N_29718);
or U29939 (N_29939,N_29643,N_29563);
nor U29940 (N_29940,N_29627,N_29727);
nand U29941 (N_29941,N_29532,N_29674);
or U29942 (N_29942,N_29656,N_29705);
nor U29943 (N_29943,N_29732,N_29530);
and U29944 (N_29944,N_29583,N_29568);
and U29945 (N_29945,N_29612,N_29714);
or U29946 (N_29946,N_29559,N_29613);
nor U29947 (N_29947,N_29740,N_29503);
or U29948 (N_29948,N_29537,N_29566);
and U29949 (N_29949,N_29582,N_29586);
or U29950 (N_29950,N_29515,N_29550);
nor U29951 (N_29951,N_29606,N_29622);
or U29952 (N_29952,N_29660,N_29598);
nor U29953 (N_29953,N_29554,N_29573);
nor U29954 (N_29954,N_29550,N_29631);
nand U29955 (N_29955,N_29623,N_29650);
nand U29956 (N_29956,N_29592,N_29673);
or U29957 (N_29957,N_29624,N_29645);
nand U29958 (N_29958,N_29636,N_29667);
or U29959 (N_29959,N_29556,N_29504);
or U29960 (N_29960,N_29584,N_29743);
or U29961 (N_29961,N_29602,N_29727);
or U29962 (N_29962,N_29541,N_29548);
and U29963 (N_29963,N_29518,N_29535);
or U29964 (N_29964,N_29587,N_29561);
xnor U29965 (N_29965,N_29699,N_29510);
nand U29966 (N_29966,N_29504,N_29661);
nor U29967 (N_29967,N_29582,N_29629);
nand U29968 (N_29968,N_29528,N_29738);
nand U29969 (N_29969,N_29511,N_29740);
or U29970 (N_29970,N_29689,N_29735);
and U29971 (N_29971,N_29710,N_29745);
or U29972 (N_29972,N_29745,N_29679);
nand U29973 (N_29973,N_29557,N_29726);
or U29974 (N_29974,N_29588,N_29729);
xor U29975 (N_29975,N_29684,N_29638);
or U29976 (N_29976,N_29661,N_29565);
or U29977 (N_29977,N_29502,N_29670);
nand U29978 (N_29978,N_29720,N_29672);
xnor U29979 (N_29979,N_29736,N_29704);
or U29980 (N_29980,N_29542,N_29560);
and U29981 (N_29981,N_29673,N_29552);
nand U29982 (N_29982,N_29695,N_29622);
or U29983 (N_29983,N_29736,N_29534);
xor U29984 (N_29984,N_29693,N_29508);
and U29985 (N_29985,N_29677,N_29535);
nor U29986 (N_29986,N_29578,N_29680);
or U29987 (N_29987,N_29720,N_29617);
and U29988 (N_29988,N_29541,N_29672);
nor U29989 (N_29989,N_29743,N_29535);
nor U29990 (N_29990,N_29725,N_29744);
and U29991 (N_29991,N_29607,N_29602);
xnor U29992 (N_29992,N_29571,N_29535);
or U29993 (N_29993,N_29518,N_29720);
xnor U29994 (N_29994,N_29581,N_29504);
or U29995 (N_29995,N_29630,N_29691);
nor U29996 (N_29996,N_29577,N_29539);
or U29997 (N_29997,N_29510,N_29659);
xor U29998 (N_29998,N_29687,N_29619);
xor U29999 (N_29999,N_29598,N_29710);
nor U30000 (N_30000,N_29855,N_29844);
xnor U30001 (N_30001,N_29797,N_29991);
nand U30002 (N_30002,N_29775,N_29881);
and U30003 (N_30003,N_29793,N_29928);
and U30004 (N_30004,N_29986,N_29875);
and U30005 (N_30005,N_29895,N_29988);
and U30006 (N_30006,N_29958,N_29940);
xnor U30007 (N_30007,N_29789,N_29764);
nand U30008 (N_30008,N_29939,N_29766);
and U30009 (N_30009,N_29984,N_29791);
or U30010 (N_30010,N_29901,N_29930);
nor U30011 (N_30011,N_29880,N_29981);
nand U30012 (N_30012,N_29929,N_29985);
or U30013 (N_30013,N_29759,N_29942);
nor U30014 (N_30014,N_29811,N_29921);
and U30015 (N_30015,N_29851,N_29932);
nor U30016 (N_30016,N_29836,N_29820);
or U30017 (N_30017,N_29804,N_29805);
nor U30018 (N_30018,N_29935,N_29831);
and U30019 (N_30019,N_29852,N_29987);
or U30020 (N_30020,N_29989,N_29924);
or U30021 (N_30021,N_29946,N_29848);
and U30022 (N_30022,N_29808,N_29955);
or U30023 (N_30023,N_29916,N_29968);
or U30024 (N_30024,N_29756,N_29891);
nand U30025 (N_30025,N_29798,N_29780);
nand U30026 (N_30026,N_29967,N_29779);
or U30027 (N_30027,N_29956,N_29976);
xnor U30028 (N_30028,N_29778,N_29949);
xnor U30029 (N_30029,N_29937,N_29918);
and U30030 (N_30030,N_29890,N_29963);
nand U30031 (N_30031,N_29951,N_29898);
or U30032 (N_30032,N_29903,N_29973);
and U30033 (N_30033,N_29873,N_29944);
and U30034 (N_30034,N_29962,N_29751);
nor U30035 (N_30035,N_29977,N_29769);
and U30036 (N_30036,N_29900,N_29894);
nand U30037 (N_30037,N_29876,N_29862);
or U30038 (N_30038,N_29994,N_29752);
or U30039 (N_30039,N_29763,N_29799);
and U30040 (N_30040,N_29982,N_29992);
and U30041 (N_30041,N_29767,N_29838);
nand U30042 (N_30042,N_29867,N_29919);
nor U30043 (N_30043,N_29966,N_29926);
xnor U30044 (N_30044,N_29814,N_29801);
nand U30045 (N_30045,N_29933,N_29845);
nor U30046 (N_30046,N_29856,N_29802);
or U30047 (N_30047,N_29835,N_29923);
and U30048 (N_30048,N_29948,N_29980);
and U30049 (N_30049,N_29996,N_29888);
nand U30050 (N_30050,N_29872,N_29861);
xor U30051 (N_30051,N_29854,N_29889);
nor U30052 (N_30052,N_29765,N_29783);
or U30053 (N_30053,N_29952,N_29990);
or U30054 (N_30054,N_29897,N_29896);
or U30055 (N_30055,N_29753,N_29899);
nor U30056 (N_30056,N_29837,N_29885);
nand U30057 (N_30057,N_29817,N_29849);
or U30058 (N_30058,N_29998,N_29909);
and U30059 (N_30059,N_29954,N_29886);
and U30060 (N_30060,N_29773,N_29965);
nand U30061 (N_30061,N_29784,N_29884);
nand U30062 (N_30062,N_29863,N_29970);
nor U30063 (N_30063,N_29859,N_29761);
nor U30064 (N_30064,N_29941,N_29860);
xnor U30065 (N_30065,N_29795,N_29959);
and U30066 (N_30066,N_29882,N_29818);
nand U30067 (N_30067,N_29812,N_29813);
and U30068 (N_30068,N_29922,N_29758);
nor U30069 (N_30069,N_29830,N_29978);
nor U30070 (N_30070,N_29869,N_29853);
and U30071 (N_30071,N_29816,N_29878);
nor U30072 (N_30072,N_29822,N_29796);
and U30073 (N_30073,N_29883,N_29829);
xnor U30074 (N_30074,N_29803,N_29995);
nor U30075 (N_30075,N_29794,N_29768);
nand U30076 (N_30076,N_29931,N_29917);
xnor U30077 (N_30077,N_29842,N_29815);
xnor U30078 (N_30078,N_29999,N_29771);
or U30079 (N_30079,N_29912,N_29910);
nand U30080 (N_30080,N_29834,N_29906);
nor U30081 (N_30081,N_29866,N_29936);
nor U30082 (N_30082,N_29754,N_29927);
xor U30083 (N_30083,N_29893,N_29819);
and U30084 (N_30084,N_29925,N_29833);
nor U30085 (N_30085,N_29757,N_29902);
xnor U30086 (N_30086,N_29907,N_29774);
nand U30087 (N_30087,N_29979,N_29960);
nor U30088 (N_30088,N_29969,N_29826);
nor U30089 (N_30089,N_29915,N_29786);
nor U30090 (N_30090,N_29905,N_29957);
nor U30091 (N_30091,N_29790,N_29945);
and U30092 (N_30092,N_29892,N_29781);
nor U30093 (N_30093,N_29972,N_29950);
and U30094 (N_30094,N_29871,N_29840);
nand U30095 (N_30095,N_29839,N_29943);
nand U30096 (N_30096,N_29823,N_29810);
xor U30097 (N_30097,N_29870,N_29920);
or U30098 (N_30098,N_29914,N_29961);
or U30099 (N_30099,N_29911,N_29997);
and U30100 (N_30100,N_29755,N_29782);
xor U30101 (N_30101,N_29938,N_29843);
nor U30102 (N_30102,N_29762,N_29846);
nor U30103 (N_30103,N_29879,N_29828);
nand U30104 (N_30104,N_29864,N_29770);
xnor U30105 (N_30105,N_29953,N_29847);
and U30106 (N_30106,N_29975,N_29908);
nand U30107 (N_30107,N_29772,N_29993);
nand U30108 (N_30108,N_29787,N_29800);
and U30109 (N_30109,N_29865,N_29857);
and U30110 (N_30110,N_29964,N_29809);
xnor U30111 (N_30111,N_29841,N_29874);
xor U30112 (N_30112,N_29887,N_29974);
nand U30113 (N_30113,N_29858,N_29877);
or U30114 (N_30114,N_29850,N_29821);
nand U30115 (N_30115,N_29983,N_29760);
xor U30116 (N_30116,N_29934,N_29806);
or U30117 (N_30117,N_29785,N_29971);
or U30118 (N_30118,N_29824,N_29807);
nand U30119 (N_30119,N_29750,N_29868);
or U30120 (N_30120,N_29827,N_29777);
nor U30121 (N_30121,N_29825,N_29913);
nand U30122 (N_30122,N_29788,N_29947);
or U30123 (N_30123,N_29792,N_29832);
nand U30124 (N_30124,N_29776,N_29904);
or U30125 (N_30125,N_29836,N_29910);
nor U30126 (N_30126,N_29849,N_29959);
nand U30127 (N_30127,N_29921,N_29925);
and U30128 (N_30128,N_29782,N_29941);
xor U30129 (N_30129,N_29811,N_29764);
nand U30130 (N_30130,N_29773,N_29814);
xor U30131 (N_30131,N_29874,N_29916);
xnor U30132 (N_30132,N_29844,N_29817);
or U30133 (N_30133,N_29951,N_29786);
and U30134 (N_30134,N_29887,N_29891);
xor U30135 (N_30135,N_29825,N_29778);
and U30136 (N_30136,N_29768,N_29764);
and U30137 (N_30137,N_29763,N_29935);
and U30138 (N_30138,N_29945,N_29775);
nand U30139 (N_30139,N_29834,N_29802);
or U30140 (N_30140,N_29844,N_29979);
xor U30141 (N_30141,N_29772,N_29947);
xnor U30142 (N_30142,N_29921,N_29832);
nand U30143 (N_30143,N_29765,N_29948);
or U30144 (N_30144,N_29972,N_29828);
or U30145 (N_30145,N_29973,N_29891);
and U30146 (N_30146,N_29805,N_29771);
nand U30147 (N_30147,N_29824,N_29922);
and U30148 (N_30148,N_29760,N_29815);
nor U30149 (N_30149,N_29876,N_29844);
xor U30150 (N_30150,N_29987,N_29843);
nor U30151 (N_30151,N_29765,N_29896);
or U30152 (N_30152,N_29953,N_29932);
nand U30153 (N_30153,N_29953,N_29788);
nor U30154 (N_30154,N_29772,N_29920);
nand U30155 (N_30155,N_29802,N_29982);
and U30156 (N_30156,N_29969,N_29840);
and U30157 (N_30157,N_29797,N_29992);
and U30158 (N_30158,N_29825,N_29889);
nor U30159 (N_30159,N_29845,N_29876);
and U30160 (N_30160,N_29828,N_29795);
xnor U30161 (N_30161,N_29763,N_29936);
nand U30162 (N_30162,N_29925,N_29934);
nor U30163 (N_30163,N_29814,N_29791);
and U30164 (N_30164,N_29965,N_29971);
nor U30165 (N_30165,N_29852,N_29851);
or U30166 (N_30166,N_29971,N_29918);
xor U30167 (N_30167,N_29931,N_29839);
xnor U30168 (N_30168,N_29816,N_29897);
or U30169 (N_30169,N_29966,N_29860);
or U30170 (N_30170,N_29878,N_29822);
nor U30171 (N_30171,N_29813,N_29991);
nand U30172 (N_30172,N_29838,N_29904);
xor U30173 (N_30173,N_29821,N_29996);
or U30174 (N_30174,N_29953,N_29780);
xnor U30175 (N_30175,N_29814,N_29883);
and U30176 (N_30176,N_29876,N_29978);
nor U30177 (N_30177,N_29800,N_29900);
and U30178 (N_30178,N_29829,N_29985);
nor U30179 (N_30179,N_29805,N_29836);
xor U30180 (N_30180,N_29821,N_29893);
and U30181 (N_30181,N_29960,N_29892);
or U30182 (N_30182,N_29967,N_29914);
and U30183 (N_30183,N_29841,N_29916);
nor U30184 (N_30184,N_29753,N_29837);
xor U30185 (N_30185,N_29873,N_29789);
or U30186 (N_30186,N_29764,N_29966);
nor U30187 (N_30187,N_29846,N_29811);
nand U30188 (N_30188,N_29751,N_29920);
nand U30189 (N_30189,N_29885,N_29879);
xnor U30190 (N_30190,N_29911,N_29757);
xnor U30191 (N_30191,N_29880,N_29771);
xor U30192 (N_30192,N_29974,N_29944);
and U30193 (N_30193,N_29922,N_29994);
nor U30194 (N_30194,N_29772,N_29926);
xor U30195 (N_30195,N_29857,N_29983);
and U30196 (N_30196,N_29853,N_29911);
xnor U30197 (N_30197,N_29945,N_29802);
xnor U30198 (N_30198,N_29873,N_29959);
nand U30199 (N_30199,N_29812,N_29882);
or U30200 (N_30200,N_29813,N_29832);
nand U30201 (N_30201,N_29803,N_29989);
nand U30202 (N_30202,N_29806,N_29840);
and U30203 (N_30203,N_29760,N_29819);
or U30204 (N_30204,N_29820,N_29992);
or U30205 (N_30205,N_29850,N_29965);
xor U30206 (N_30206,N_29896,N_29941);
nand U30207 (N_30207,N_29882,N_29753);
nor U30208 (N_30208,N_29953,N_29991);
or U30209 (N_30209,N_29795,N_29767);
nor U30210 (N_30210,N_29798,N_29793);
and U30211 (N_30211,N_29953,N_29762);
xnor U30212 (N_30212,N_29861,N_29761);
xor U30213 (N_30213,N_29913,N_29789);
and U30214 (N_30214,N_29923,N_29836);
xor U30215 (N_30215,N_29862,N_29973);
and U30216 (N_30216,N_29856,N_29890);
and U30217 (N_30217,N_29806,N_29857);
xor U30218 (N_30218,N_29847,N_29931);
nand U30219 (N_30219,N_29817,N_29838);
xnor U30220 (N_30220,N_29762,N_29898);
nor U30221 (N_30221,N_29860,N_29962);
nor U30222 (N_30222,N_29884,N_29956);
xor U30223 (N_30223,N_29961,N_29897);
xor U30224 (N_30224,N_29945,N_29981);
xor U30225 (N_30225,N_29917,N_29879);
xor U30226 (N_30226,N_29938,N_29947);
xor U30227 (N_30227,N_29811,N_29892);
xor U30228 (N_30228,N_29929,N_29885);
nor U30229 (N_30229,N_29908,N_29940);
and U30230 (N_30230,N_29764,N_29833);
and U30231 (N_30231,N_29943,N_29940);
nand U30232 (N_30232,N_29860,N_29914);
nand U30233 (N_30233,N_29920,N_29951);
nand U30234 (N_30234,N_29752,N_29964);
xnor U30235 (N_30235,N_29798,N_29751);
or U30236 (N_30236,N_29818,N_29830);
or U30237 (N_30237,N_29777,N_29791);
and U30238 (N_30238,N_29954,N_29930);
nand U30239 (N_30239,N_29909,N_29981);
xnor U30240 (N_30240,N_29958,N_29925);
nor U30241 (N_30241,N_29913,N_29808);
nand U30242 (N_30242,N_29880,N_29787);
nand U30243 (N_30243,N_29934,N_29797);
nand U30244 (N_30244,N_29941,N_29870);
and U30245 (N_30245,N_29978,N_29937);
or U30246 (N_30246,N_29995,N_29836);
or U30247 (N_30247,N_29951,N_29794);
or U30248 (N_30248,N_29809,N_29958);
nand U30249 (N_30249,N_29762,N_29927);
nand U30250 (N_30250,N_30243,N_30146);
and U30251 (N_30251,N_30054,N_30018);
and U30252 (N_30252,N_30182,N_30229);
xnor U30253 (N_30253,N_30239,N_30069);
nor U30254 (N_30254,N_30209,N_30196);
nand U30255 (N_30255,N_30217,N_30019);
and U30256 (N_30256,N_30166,N_30142);
or U30257 (N_30257,N_30023,N_30130);
nor U30258 (N_30258,N_30074,N_30076);
or U30259 (N_30259,N_30103,N_30248);
xor U30260 (N_30260,N_30068,N_30035);
nand U30261 (N_30261,N_30043,N_30013);
and U30262 (N_30262,N_30227,N_30240);
xnor U30263 (N_30263,N_30159,N_30040);
and U30264 (N_30264,N_30057,N_30150);
nor U30265 (N_30265,N_30176,N_30101);
nor U30266 (N_30266,N_30145,N_30088);
or U30267 (N_30267,N_30049,N_30156);
xnor U30268 (N_30268,N_30056,N_30032);
nor U30269 (N_30269,N_30026,N_30093);
or U30270 (N_30270,N_30098,N_30090);
or U30271 (N_30271,N_30204,N_30216);
and U30272 (N_30272,N_30014,N_30131);
or U30273 (N_30273,N_30165,N_30155);
xnor U30274 (N_30274,N_30108,N_30121);
nand U30275 (N_30275,N_30010,N_30061);
xnor U30276 (N_30276,N_30081,N_30193);
nand U30277 (N_30277,N_30022,N_30021);
nor U30278 (N_30278,N_30089,N_30137);
nand U30279 (N_30279,N_30042,N_30200);
nand U30280 (N_30280,N_30122,N_30083);
nor U30281 (N_30281,N_30114,N_30214);
nor U30282 (N_30282,N_30100,N_30207);
and U30283 (N_30283,N_30141,N_30181);
nor U30284 (N_30284,N_30194,N_30231);
or U30285 (N_30285,N_30185,N_30084);
and U30286 (N_30286,N_30167,N_30027);
and U30287 (N_30287,N_30161,N_30197);
or U30288 (N_30288,N_30188,N_30147);
or U30289 (N_30289,N_30051,N_30012);
nand U30290 (N_30290,N_30111,N_30191);
or U30291 (N_30291,N_30139,N_30078);
nand U30292 (N_30292,N_30199,N_30091);
xor U30293 (N_30293,N_30170,N_30039);
nand U30294 (N_30294,N_30237,N_30112);
and U30295 (N_30295,N_30046,N_30065);
nor U30296 (N_30296,N_30143,N_30002);
nand U30297 (N_30297,N_30151,N_30205);
nand U30298 (N_30298,N_30158,N_30235);
xor U30299 (N_30299,N_30006,N_30082);
xnor U30300 (N_30300,N_30080,N_30183);
and U30301 (N_30301,N_30228,N_30178);
nor U30302 (N_30302,N_30236,N_30241);
and U30303 (N_30303,N_30055,N_30050);
and U30304 (N_30304,N_30126,N_30104);
nor U30305 (N_30305,N_30160,N_30172);
or U30306 (N_30306,N_30038,N_30109);
nand U30307 (N_30307,N_30123,N_30226);
and U30308 (N_30308,N_30168,N_30249);
and U30309 (N_30309,N_30025,N_30059);
xnor U30310 (N_30310,N_30000,N_30222);
nand U30311 (N_30311,N_30071,N_30174);
xnor U30312 (N_30312,N_30186,N_30127);
nor U30313 (N_30313,N_30015,N_30052);
nor U30314 (N_30314,N_30060,N_30175);
and U30315 (N_30315,N_30187,N_30233);
and U30316 (N_30316,N_30219,N_30213);
xor U30317 (N_30317,N_30230,N_30223);
and U30318 (N_30318,N_30198,N_30140);
xnor U30319 (N_30319,N_30184,N_30124);
xnor U30320 (N_30320,N_30009,N_30007);
or U30321 (N_30321,N_30134,N_30117);
nand U30322 (N_30322,N_30144,N_30220);
nand U30323 (N_30323,N_30244,N_30033);
xor U30324 (N_30324,N_30095,N_30164);
and U30325 (N_30325,N_30116,N_30031);
xor U30326 (N_30326,N_30092,N_30148);
and U30327 (N_30327,N_30062,N_30138);
nor U30328 (N_30328,N_30099,N_30173);
nor U30329 (N_30329,N_30149,N_30005);
nand U30330 (N_30330,N_30096,N_30129);
nand U30331 (N_30331,N_30118,N_30047);
or U30332 (N_30332,N_30058,N_30232);
nor U30333 (N_30333,N_30133,N_30105);
or U30334 (N_30334,N_30064,N_30215);
nor U30335 (N_30335,N_30041,N_30119);
and U30336 (N_30336,N_30020,N_30211);
xor U30337 (N_30337,N_30208,N_30177);
and U30338 (N_30338,N_30189,N_30135);
xor U30339 (N_30339,N_30048,N_30086);
nand U30340 (N_30340,N_30073,N_30245);
xnor U30341 (N_30341,N_30094,N_30224);
or U30342 (N_30342,N_30028,N_30106);
nand U30343 (N_30343,N_30218,N_30045);
nor U30344 (N_30344,N_30179,N_30037);
or U30345 (N_30345,N_30210,N_30132);
nand U30346 (N_30346,N_30008,N_30153);
nand U30347 (N_30347,N_30225,N_30075);
xnor U30348 (N_30348,N_30169,N_30072);
or U30349 (N_30349,N_30034,N_30003);
xor U30350 (N_30350,N_30180,N_30085);
xor U30351 (N_30351,N_30162,N_30202);
and U30352 (N_30352,N_30011,N_30201);
xnor U30353 (N_30353,N_30001,N_30163);
nor U30354 (N_30354,N_30125,N_30113);
xnor U30355 (N_30355,N_30238,N_30077);
and U30356 (N_30356,N_30203,N_30044);
and U30357 (N_30357,N_30154,N_30053);
nand U30358 (N_30358,N_30120,N_30017);
nor U30359 (N_30359,N_30004,N_30107);
nor U30360 (N_30360,N_30136,N_30016);
nor U30361 (N_30361,N_30206,N_30171);
nor U30362 (N_30362,N_30190,N_30128);
or U30363 (N_30363,N_30102,N_30087);
and U30364 (N_30364,N_30242,N_30212);
and U30365 (N_30365,N_30115,N_30070);
xnor U30366 (N_30366,N_30221,N_30192);
xor U30367 (N_30367,N_30029,N_30067);
nor U30368 (N_30368,N_30036,N_30234);
nor U30369 (N_30369,N_30030,N_30097);
nand U30370 (N_30370,N_30063,N_30024);
xnor U30371 (N_30371,N_30195,N_30157);
and U30372 (N_30372,N_30079,N_30152);
nand U30373 (N_30373,N_30066,N_30110);
and U30374 (N_30374,N_30246,N_30247);
nand U30375 (N_30375,N_30017,N_30091);
and U30376 (N_30376,N_30230,N_30175);
nand U30377 (N_30377,N_30199,N_30154);
nand U30378 (N_30378,N_30169,N_30173);
nand U30379 (N_30379,N_30010,N_30024);
nand U30380 (N_30380,N_30030,N_30163);
nand U30381 (N_30381,N_30088,N_30034);
or U30382 (N_30382,N_30060,N_30189);
and U30383 (N_30383,N_30239,N_30042);
and U30384 (N_30384,N_30230,N_30106);
nand U30385 (N_30385,N_30239,N_30116);
nand U30386 (N_30386,N_30063,N_30030);
and U30387 (N_30387,N_30106,N_30022);
nor U30388 (N_30388,N_30231,N_30040);
and U30389 (N_30389,N_30125,N_30115);
or U30390 (N_30390,N_30134,N_30129);
nor U30391 (N_30391,N_30193,N_30098);
xor U30392 (N_30392,N_30174,N_30059);
xor U30393 (N_30393,N_30237,N_30024);
or U30394 (N_30394,N_30196,N_30174);
nand U30395 (N_30395,N_30129,N_30070);
and U30396 (N_30396,N_30074,N_30133);
or U30397 (N_30397,N_30188,N_30149);
nor U30398 (N_30398,N_30100,N_30203);
and U30399 (N_30399,N_30038,N_30176);
xnor U30400 (N_30400,N_30244,N_30211);
nand U30401 (N_30401,N_30024,N_30176);
nand U30402 (N_30402,N_30059,N_30183);
or U30403 (N_30403,N_30026,N_30168);
nor U30404 (N_30404,N_30161,N_30014);
nor U30405 (N_30405,N_30146,N_30178);
xor U30406 (N_30406,N_30032,N_30074);
nor U30407 (N_30407,N_30037,N_30043);
or U30408 (N_30408,N_30233,N_30096);
nor U30409 (N_30409,N_30110,N_30130);
nor U30410 (N_30410,N_30137,N_30173);
nand U30411 (N_30411,N_30033,N_30173);
and U30412 (N_30412,N_30143,N_30249);
nor U30413 (N_30413,N_30119,N_30182);
nor U30414 (N_30414,N_30119,N_30155);
nand U30415 (N_30415,N_30148,N_30201);
nor U30416 (N_30416,N_30101,N_30113);
or U30417 (N_30417,N_30011,N_30086);
and U30418 (N_30418,N_30127,N_30245);
nor U30419 (N_30419,N_30153,N_30036);
or U30420 (N_30420,N_30089,N_30093);
and U30421 (N_30421,N_30186,N_30102);
or U30422 (N_30422,N_30094,N_30095);
nand U30423 (N_30423,N_30191,N_30070);
xor U30424 (N_30424,N_30097,N_30022);
nor U30425 (N_30425,N_30216,N_30173);
or U30426 (N_30426,N_30198,N_30154);
xnor U30427 (N_30427,N_30087,N_30030);
or U30428 (N_30428,N_30158,N_30048);
or U30429 (N_30429,N_30199,N_30202);
nand U30430 (N_30430,N_30209,N_30083);
xor U30431 (N_30431,N_30097,N_30001);
nand U30432 (N_30432,N_30244,N_30128);
and U30433 (N_30433,N_30002,N_30068);
nor U30434 (N_30434,N_30071,N_30175);
xnor U30435 (N_30435,N_30206,N_30055);
nand U30436 (N_30436,N_30038,N_30187);
or U30437 (N_30437,N_30245,N_30106);
and U30438 (N_30438,N_30062,N_30038);
and U30439 (N_30439,N_30227,N_30226);
xnor U30440 (N_30440,N_30120,N_30007);
or U30441 (N_30441,N_30217,N_30146);
nor U30442 (N_30442,N_30222,N_30149);
nand U30443 (N_30443,N_30159,N_30056);
or U30444 (N_30444,N_30047,N_30083);
and U30445 (N_30445,N_30124,N_30214);
or U30446 (N_30446,N_30079,N_30198);
nand U30447 (N_30447,N_30074,N_30185);
nor U30448 (N_30448,N_30246,N_30023);
nand U30449 (N_30449,N_30238,N_30088);
nand U30450 (N_30450,N_30115,N_30121);
or U30451 (N_30451,N_30000,N_30089);
nor U30452 (N_30452,N_30208,N_30022);
nand U30453 (N_30453,N_30175,N_30134);
nand U30454 (N_30454,N_30126,N_30057);
and U30455 (N_30455,N_30020,N_30142);
nand U30456 (N_30456,N_30017,N_30149);
xor U30457 (N_30457,N_30099,N_30165);
xor U30458 (N_30458,N_30144,N_30047);
and U30459 (N_30459,N_30118,N_30044);
and U30460 (N_30460,N_30154,N_30086);
xnor U30461 (N_30461,N_30077,N_30065);
nor U30462 (N_30462,N_30110,N_30207);
or U30463 (N_30463,N_30157,N_30087);
nand U30464 (N_30464,N_30230,N_30082);
or U30465 (N_30465,N_30052,N_30173);
xnor U30466 (N_30466,N_30159,N_30051);
or U30467 (N_30467,N_30008,N_30137);
or U30468 (N_30468,N_30236,N_30026);
xnor U30469 (N_30469,N_30179,N_30124);
nand U30470 (N_30470,N_30094,N_30017);
or U30471 (N_30471,N_30113,N_30190);
nand U30472 (N_30472,N_30199,N_30120);
nor U30473 (N_30473,N_30219,N_30093);
xor U30474 (N_30474,N_30116,N_30242);
and U30475 (N_30475,N_30222,N_30154);
nand U30476 (N_30476,N_30014,N_30008);
nor U30477 (N_30477,N_30212,N_30109);
and U30478 (N_30478,N_30049,N_30103);
nand U30479 (N_30479,N_30083,N_30193);
or U30480 (N_30480,N_30205,N_30193);
xor U30481 (N_30481,N_30161,N_30003);
or U30482 (N_30482,N_30210,N_30088);
and U30483 (N_30483,N_30207,N_30172);
nor U30484 (N_30484,N_30153,N_30193);
or U30485 (N_30485,N_30025,N_30249);
or U30486 (N_30486,N_30039,N_30200);
nand U30487 (N_30487,N_30091,N_30055);
or U30488 (N_30488,N_30011,N_30089);
xor U30489 (N_30489,N_30011,N_30120);
nand U30490 (N_30490,N_30191,N_30073);
nor U30491 (N_30491,N_30145,N_30004);
nor U30492 (N_30492,N_30123,N_30239);
or U30493 (N_30493,N_30201,N_30178);
or U30494 (N_30494,N_30002,N_30185);
xnor U30495 (N_30495,N_30219,N_30031);
nor U30496 (N_30496,N_30039,N_30161);
or U30497 (N_30497,N_30066,N_30206);
nand U30498 (N_30498,N_30133,N_30207);
nor U30499 (N_30499,N_30111,N_30161);
xor U30500 (N_30500,N_30301,N_30302);
or U30501 (N_30501,N_30273,N_30438);
and U30502 (N_30502,N_30381,N_30360);
xnor U30503 (N_30503,N_30480,N_30303);
nor U30504 (N_30504,N_30370,N_30473);
nor U30505 (N_30505,N_30464,N_30304);
and U30506 (N_30506,N_30433,N_30478);
or U30507 (N_30507,N_30293,N_30452);
nand U30508 (N_30508,N_30449,N_30476);
nor U30509 (N_30509,N_30368,N_30295);
and U30510 (N_30510,N_30484,N_30399);
xnor U30511 (N_30511,N_30494,N_30441);
nor U30512 (N_30512,N_30489,N_30471);
nor U30513 (N_30513,N_30405,N_30474);
nor U30514 (N_30514,N_30428,N_30364);
and U30515 (N_30515,N_30340,N_30400);
and U30516 (N_30516,N_30334,N_30435);
and U30517 (N_30517,N_30416,N_30406);
nand U30518 (N_30518,N_30289,N_30493);
nor U30519 (N_30519,N_30294,N_30342);
nor U30520 (N_30520,N_30292,N_30350);
and U30521 (N_30521,N_30475,N_30425);
or U30522 (N_30522,N_30314,N_30357);
or U30523 (N_30523,N_30419,N_30491);
nor U30524 (N_30524,N_30281,N_30412);
nand U30525 (N_30525,N_30498,N_30254);
xor U30526 (N_30526,N_30403,N_30444);
nand U30527 (N_30527,N_30311,N_30422);
xor U30528 (N_30528,N_30366,N_30454);
and U30529 (N_30529,N_30459,N_30321);
nor U30530 (N_30530,N_30417,N_30277);
nor U30531 (N_30531,N_30495,N_30255);
or U30532 (N_30532,N_30279,N_30287);
or U30533 (N_30533,N_30466,N_30401);
nor U30534 (N_30534,N_30414,N_30463);
nor U30535 (N_30535,N_30477,N_30358);
nor U30536 (N_30536,N_30354,N_30308);
nor U30537 (N_30537,N_30367,N_30392);
nor U30538 (N_30538,N_30499,N_30420);
nor U30539 (N_30539,N_30413,N_30408);
or U30540 (N_30540,N_30250,N_30424);
or U30541 (N_30541,N_30300,N_30356);
and U30542 (N_30542,N_30305,N_30266);
or U30543 (N_30543,N_30252,N_30329);
nor U30544 (N_30544,N_30487,N_30256);
nor U30545 (N_30545,N_30497,N_30430);
nand U30546 (N_30546,N_30389,N_30328);
and U30547 (N_30547,N_30258,N_30393);
or U30548 (N_30548,N_30415,N_30343);
nor U30549 (N_30549,N_30299,N_30421);
or U30550 (N_30550,N_30330,N_30376);
and U30551 (N_30551,N_30359,N_30468);
nand U30552 (N_30552,N_30317,N_30465);
or U30553 (N_30553,N_30355,N_30398);
or U30554 (N_30554,N_30410,N_30351);
nand U30555 (N_30555,N_30327,N_30490);
xor U30556 (N_30556,N_30352,N_30492);
xor U30557 (N_30557,N_30427,N_30275);
nand U30558 (N_30558,N_30479,N_30390);
or U30559 (N_30559,N_30386,N_30269);
or U30560 (N_30560,N_30482,N_30278);
nand U30561 (N_30561,N_30394,N_30335);
or U30562 (N_30562,N_30396,N_30439);
nand U30563 (N_30563,N_30318,N_30272);
and U30564 (N_30564,N_30257,N_30338);
xor U30565 (N_30565,N_30387,N_30319);
nor U30566 (N_30566,N_30467,N_30402);
nor U30567 (N_30567,N_30426,N_30455);
or U30568 (N_30568,N_30333,N_30409);
and U30569 (N_30569,N_30280,N_30320);
xor U30570 (N_30570,N_30253,N_30445);
and U30571 (N_30571,N_30375,N_30404);
or U30572 (N_30572,N_30259,N_30348);
xor U30573 (N_30573,N_30397,N_30458);
and U30574 (N_30574,N_30462,N_30418);
or U30575 (N_30575,N_30361,N_30378);
nor U30576 (N_30576,N_30431,N_30460);
nand U30577 (N_30577,N_30344,N_30251);
xor U30578 (N_30578,N_30310,N_30411);
xor U30579 (N_30579,N_30331,N_30461);
xnor U30580 (N_30580,N_30285,N_30345);
nand U30581 (N_30581,N_30385,N_30353);
nor U30582 (N_30582,N_30380,N_30496);
nand U30583 (N_30583,N_30263,N_30347);
or U30584 (N_30584,N_30296,N_30270);
nand U30585 (N_30585,N_30339,N_30432);
nand U30586 (N_30586,N_30325,N_30448);
xnor U30587 (N_30587,N_30288,N_30264);
nand U30588 (N_30588,N_30434,N_30332);
nor U30589 (N_30589,N_30260,N_30282);
xnor U30590 (N_30590,N_30450,N_30324);
nand U30591 (N_30591,N_30261,N_30442);
xor U30592 (N_30592,N_30483,N_30383);
xnor U30593 (N_30593,N_30322,N_30436);
xnor U30594 (N_30594,N_30371,N_30395);
xnor U30595 (N_30595,N_30446,N_30374);
xor U30596 (N_30596,N_30312,N_30323);
or U30597 (N_30597,N_30429,N_30309);
or U30598 (N_30598,N_30265,N_30382);
and U30599 (N_30599,N_30336,N_30365);
nor U30600 (N_30600,N_30341,N_30457);
nand U30601 (N_30601,N_30298,N_30407);
xor U30602 (N_30602,N_30326,N_30362);
nand U30603 (N_30603,N_30440,N_30262);
nand U30604 (N_30604,N_30349,N_30486);
nor U30605 (N_30605,N_30451,N_30276);
nand U30606 (N_30606,N_30391,N_30469);
nand U30607 (N_30607,N_30286,N_30373);
xor U30608 (N_30608,N_30297,N_30268);
nand U30609 (N_30609,N_30337,N_30423);
nor U30610 (N_30610,N_30372,N_30447);
nand U30611 (N_30611,N_30346,N_30316);
or U30612 (N_30612,N_30488,N_30437);
nor U30613 (N_30613,N_30384,N_30290);
nand U30614 (N_30614,N_30481,N_30313);
xnor U30615 (N_30615,N_30388,N_30470);
nand U30616 (N_30616,N_30291,N_30271);
nand U30617 (N_30617,N_30307,N_30369);
and U30618 (N_30618,N_30443,N_30306);
xnor U30619 (N_30619,N_30274,N_30315);
or U30620 (N_30620,N_30283,N_30472);
or U30621 (N_30621,N_30284,N_30453);
nor U30622 (N_30622,N_30379,N_30363);
or U30623 (N_30623,N_30377,N_30267);
nor U30624 (N_30624,N_30485,N_30456);
nor U30625 (N_30625,N_30288,N_30458);
nand U30626 (N_30626,N_30297,N_30481);
nor U30627 (N_30627,N_30473,N_30493);
nor U30628 (N_30628,N_30280,N_30495);
xnor U30629 (N_30629,N_30270,N_30416);
and U30630 (N_30630,N_30451,N_30492);
or U30631 (N_30631,N_30289,N_30309);
or U30632 (N_30632,N_30292,N_30373);
and U30633 (N_30633,N_30299,N_30481);
nor U30634 (N_30634,N_30321,N_30414);
xor U30635 (N_30635,N_30407,N_30272);
and U30636 (N_30636,N_30368,N_30346);
or U30637 (N_30637,N_30382,N_30307);
and U30638 (N_30638,N_30458,N_30363);
and U30639 (N_30639,N_30341,N_30266);
nor U30640 (N_30640,N_30262,N_30453);
or U30641 (N_30641,N_30329,N_30493);
or U30642 (N_30642,N_30395,N_30269);
and U30643 (N_30643,N_30341,N_30290);
nor U30644 (N_30644,N_30298,N_30270);
nand U30645 (N_30645,N_30316,N_30286);
and U30646 (N_30646,N_30334,N_30419);
xor U30647 (N_30647,N_30326,N_30374);
nor U30648 (N_30648,N_30266,N_30461);
nor U30649 (N_30649,N_30260,N_30372);
and U30650 (N_30650,N_30315,N_30445);
nor U30651 (N_30651,N_30321,N_30419);
xnor U30652 (N_30652,N_30473,N_30338);
xnor U30653 (N_30653,N_30484,N_30461);
nand U30654 (N_30654,N_30389,N_30448);
or U30655 (N_30655,N_30482,N_30345);
nor U30656 (N_30656,N_30429,N_30380);
nand U30657 (N_30657,N_30416,N_30374);
or U30658 (N_30658,N_30300,N_30373);
nand U30659 (N_30659,N_30491,N_30396);
or U30660 (N_30660,N_30396,N_30473);
xnor U30661 (N_30661,N_30447,N_30260);
nor U30662 (N_30662,N_30385,N_30427);
nor U30663 (N_30663,N_30301,N_30291);
nand U30664 (N_30664,N_30400,N_30421);
nand U30665 (N_30665,N_30403,N_30339);
and U30666 (N_30666,N_30336,N_30300);
xnor U30667 (N_30667,N_30409,N_30441);
nand U30668 (N_30668,N_30393,N_30353);
or U30669 (N_30669,N_30420,N_30326);
nor U30670 (N_30670,N_30267,N_30378);
nor U30671 (N_30671,N_30335,N_30329);
xnor U30672 (N_30672,N_30328,N_30482);
and U30673 (N_30673,N_30492,N_30440);
or U30674 (N_30674,N_30471,N_30441);
xor U30675 (N_30675,N_30473,N_30293);
or U30676 (N_30676,N_30436,N_30420);
nor U30677 (N_30677,N_30367,N_30458);
and U30678 (N_30678,N_30432,N_30411);
xnor U30679 (N_30679,N_30270,N_30407);
or U30680 (N_30680,N_30419,N_30429);
nor U30681 (N_30681,N_30445,N_30313);
xor U30682 (N_30682,N_30338,N_30460);
xor U30683 (N_30683,N_30313,N_30419);
and U30684 (N_30684,N_30426,N_30261);
nor U30685 (N_30685,N_30348,N_30415);
nand U30686 (N_30686,N_30451,N_30266);
or U30687 (N_30687,N_30465,N_30439);
nand U30688 (N_30688,N_30293,N_30366);
and U30689 (N_30689,N_30408,N_30299);
or U30690 (N_30690,N_30254,N_30343);
nor U30691 (N_30691,N_30308,N_30421);
nor U30692 (N_30692,N_30348,N_30464);
nand U30693 (N_30693,N_30436,N_30287);
xnor U30694 (N_30694,N_30396,N_30379);
nor U30695 (N_30695,N_30459,N_30427);
and U30696 (N_30696,N_30278,N_30415);
nor U30697 (N_30697,N_30452,N_30346);
nor U30698 (N_30698,N_30431,N_30351);
and U30699 (N_30699,N_30459,N_30378);
nand U30700 (N_30700,N_30407,N_30263);
xnor U30701 (N_30701,N_30308,N_30418);
or U30702 (N_30702,N_30423,N_30334);
or U30703 (N_30703,N_30388,N_30400);
nor U30704 (N_30704,N_30384,N_30335);
nor U30705 (N_30705,N_30368,N_30366);
nor U30706 (N_30706,N_30331,N_30362);
nor U30707 (N_30707,N_30466,N_30408);
xor U30708 (N_30708,N_30381,N_30435);
or U30709 (N_30709,N_30293,N_30291);
nor U30710 (N_30710,N_30258,N_30282);
and U30711 (N_30711,N_30404,N_30406);
nor U30712 (N_30712,N_30293,N_30257);
or U30713 (N_30713,N_30342,N_30419);
xor U30714 (N_30714,N_30305,N_30435);
nor U30715 (N_30715,N_30435,N_30491);
xnor U30716 (N_30716,N_30256,N_30322);
or U30717 (N_30717,N_30306,N_30402);
or U30718 (N_30718,N_30486,N_30353);
and U30719 (N_30719,N_30403,N_30475);
xnor U30720 (N_30720,N_30278,N_30419);
xnor U30721 (N_30721,N_30399,N_30451);
and U30722 (N_30722,N_30301,N_30492);
nor U30723 (N_30723,N_30387,N_30415);
nor U30724 (N_30724,N_30282,N_30273);
nand U30725 (N_30725,N_30336,N_30324);
or U30726 (N_30726,N_30406,N_30278);
xnor U30727 (N_30727,N_30266,N_30286);
nor U30728 (N_30728,N_30399,N_30302);
or U30729 (N_30729,N_30418,N_30324);
and U30730 (N_30730,N_30293,N_30381);
and U30731 (N_30731,N_30312,N_30353);
or U30732 (N_30732,N_30354,N_30360);
nand U30733 (N_30733,N_30363,N_30494);
xnor U30734 (N_30734,N_30493,N_30453);
nor U30735 (N_30735,N_30374,N_30396);
xnor U30736 (N_30736,N_30429,N_30310);
and U30737 (N_30737,N_30377,N_30435);
or U30738 (N_30738,N_30433,N_30332);
nand U30739 (N_30739,N_30466,N_30361);
nand U30740 (N_30740,N_30385,N_30361);
xnor U30741 (N_30741,N_30396,N_30291);
nor U30742 (N_30742,N_30486,N_30442);
nor U30743 (N_30743,N_30263,N_30404);
nand U30744 (N_30744,N_30332,N_30290);
nor U30745 (N_30745,N_30391,N_30296);
nand U30746 (N_30746,N_30472,N_30420);
nor U30747 (N_30747,N_30487,N_30291);
nor U30748 (N_30748,N_30279,N_30476);
or U30749 (N_30749,N_30255,N_30471);
nand U30750 (N_30750,N_30655,N_30637);
xor U30751 (N_30751,N_30679,N_30500);
and U30752 (N_30752,N_30591,N_30505);
nand U30753 (N_30753,N_30544,N_30690);
xnor U30754 (N_30754,N_30718,N_30576);
nor U30755 (N_30755,N_30732,N_30636);
nor U30756 (N_30756,N_30543,N_30578);
and U30757 (N_30757,N_30736,N_30553);
xnor U30758 (N_30758,N_30541,N_30599);
or U30759 (N_30759,N_30532,N_30564);
nand U30760 (N_30760,N_30714,N_30733);
nor U30761 (N_30761,N_30674,N_30625);
and U30762 (N_30762,N_30740,N_30744);
and U30763 (N_30763,N_30589,N_30725);
and U30764 (N_30764,N_30535,N_30582);
and U30765 (N_30765,N_30600,N_30608);
and U30766 (N_30766,N_30570,N_30552);
and U30767 (N_30767,N_30703,N_30648);
nand U30768 (N_30768,N_30723,N_30737);
and U30769 (N_30769,N_30709,N_30601);
and U30770 (N_30770,N_30594,N_30524);
or U30771 (N_30771,N_30663,N_30638);
or U30772 (N_30772,N_30503,N_30537);
xor U30773 (N_30773,N_30707,N_30610);
nand U30774 (N_30774,N_30516,N_30701);
and U30775 (N_30775,N_30745,N_30586);
and U30776 (N_30776,N_30743,N_30502);
xnor U30777 (N_30777,N_30706,N_30595);
or U30778 (N_30778,N_30699,N_30546);
nor U30779 (N_30779,N_30661,N_30548);
and U30780 (N_30780,N_30504,N_30583);
nor U30781 (N_30781,N_30569,N_30649);
nand U30782 (N_30782,N_30641,N_30566);
nand U30783 (N_30783,N_30635,N_30511);
and U30784 (N_30784,N_30673,N_30710);
xnor U30785 (N_30785,N_30551,N_30726);
or U30786 (N_30786,N_30689,N_30572);
nor U30787 (N_30787,N_30550,N_30685);
or U30788 (N_30788,N_30514,N_30588);
or U30789 (N_30789,N_30618,N_30518);
and U30790 (N_30790,N_30529,N_30691);
xor U30791 (N_30791,N_30603,N_30615);
and U30792 (N_30792,N_30507,N_30696);
xor U30793 (N_30793,N_30560,N_30510);
nor U30794 (N_30794,N_30687,N_30509);
or U30795 (N_30795,N_30640,N_30590);
nor U30796 (N_30796,N_30680,N_30688);
or U30797 (N_30797,N_30693,N_30735);
xnor U30798 (N_30798,N_30580,N_30659);
nor U30799 (N_30799,N_30665,N_30587);
and U30800 (N_30800,N_30530,N_30712);
xnor U30801 (N_30801,N_30538,N_30585);
nor U30802 (N_30802,N_30719,N_30660);
nand U30803 (N_30803,N_30644,N_30748);
nor U30804 (N_30804,N_30639,N_30656);
and U30805 (N_30805,N_30547,N_30683);
nand U30806 (N_30806,N_30645,N_30624);
nor U30807 (N_30807,N_30506,N_30562);
xnor U30808 (N_30808,N_30720,N_30556);
or U30809 (N_30809,N_30702,N_30728);
and U30810 (N_30810,N_30670,N_30571);
and U30811 (N_30811,N_30606,N_30573);
nand U30812 (N_30812,N_30676,N_30581);
or U30813 (N_30813,N_30746,N_30626);
xnor U30814 (N_30814,N_30558,N_30682);
nor U30815 (N_30815,N_30686,N_30633);
nand U30816 (N_30816,N_30597,N_30575);
and U30817 (N_30817,N_30731,N_30631);
or U30818 (N_30818,N_30721,N_30708);
xnor U30819 (N_30819,N_30651,N_30675);
or U30820 (N_30820,N_30711,N_30646);
xnor U30821 (N_30821,N_30695,N_30577);
xor U30822 (N_30822,N_30684,N_30734);
or U30823 (N_30823,N_30523,N_30525);
and U30824 (N_30824,N_30555,N_30559);
and U30825 (N_30825,N_30724,N_30527);
or U30826 (N_30826,N_30579,N_30628);
and U30827 (N_30827,N_30658,N_30622);
nor U30828 (N_30828,N_30747,N_30704);
nand U30829 (N_30829,N_30602,N_30520);
or U30830 (N_30830,N_30643,N_30522);
nor U30831 (N_30831,N_30654,N_30619);
and U30832 (N_30832,N_30632,N_30738);
and U30833 (N_30833,N_30700,N_30604);
nand U30834 (N_30834,N_30713,N_30554);
or U30835 (N_30835,N_30681,N_30705);
nand U30836 (N_30836,N_30526,N_30672);
nor U30837 (N_30837,N_30533,N_30607);
xor U30838 (N_30838,N_30563,N_30508);
or U30839 (N_30839,N_30664,N_30501);
xor U30840 (N_30840,N_30513,N_30741);
and U30841 (N_30841,N_30671,N_30630);
or U30842 (N_30842,N_30561,N_30519);
nand U30843 (N_30843,N_30652,N_30534);
nor U30844 (N_30844,N_30715,N_30621);
and U30845 (N_30845,N_30574,N_30609);
xnor U30846 (N_30846,N_30598,N_30568);
and U30847 (N_30847,N_30565,N_30549);
nand U30848 (N_30848,N_30545,N_30634);
or U30849 (N_30849,N_30627,N_30666);
nand U30850 (N_30850,N_30727,N_30730);
xnor U30851 (N_30851,N_30722,N_30647);
nor U30852 (N_30852,N_30616,N_30642);
and U30853 (N_30853,N_30739,N_30620);
and U30854 (N_30854,N_30694,N_30669);
xor U30855 (N_30855,N_30677,N_30584);
xor U30856 (N_30856,N_30742,N_30528);
nand U30857 (N_30857,N_30567,N_30539);
nand U30858 (N_30858,N_30612,N_30531);
nor U30859 (N_30859,N_30697,N_30662);
and U30860 (N_30860,N_30668,N_30716);
nand U30861 (N_30861,N_30650,N_30593);
or U30862 (N_30862,N_30749,N_30692);
and U30863 (N_30863,N_30605,N_30596);
or U30864 (N_30864,N_30521,N_30517);
xnor U30865 (N_30865,N_30629,N_30623);
and U30866 (N_30866,N_30540,N_30536);
nand U30867 (N_30867,N_30515,N_30592);
nand U30868 (N_30868,N_30729,N_30557);
nand U30869 (N_30869,N_30653,N_30542);
nor U30870 (N_30870,N_30667,N_30614);
nor U30871 (N_30871,N_30512,N_30611);
and U30872 (N_30872,N_30657,N_30717);
or U30873 (N_30873,N_30617,N_30613);
xor U30874 (N_30874,N_30698,N_30678);
and U30875 (N_30875,N_30579,N_30645);
xnor U30876 (N_30876,N_30742,N_30648);
xnor U30877 (N_30877,N_30519,N_30686);
and U30878 (N_30878,N_30734,N_30676);
and U30879 (N_30879,N_30556,N_30677);
nand U30880 (N_30880,N_30714,N_30651);
xor U30881 (N_30881,N_30672,N_30644);
and U30882 (N_30882,N_30523,N_30566);
or U30883 (N_30883,N_30728,N_30692);
nor U30884 (N_30884,N_30707,N_30612);
and U30885 (N_30885,N_30648,N_30512);
nor U30886 (N_30886,N_30685,N_30677);
or U30887 (N_30887,N_30578,N_30670);
and U30888 (N_30888,N_30593,N_30626);
nand U30889 (N_30889,N_30676,N_30577);
and U30890 (N_30890,N_30721,N_30745);
xnor U30891 (N_30891,N_30528,N_30611);
xnor U30892 (N_30892,N_30685,N_30522);
nor U30893 (N_30893,N_30519,N_30723);
nand U30894 (N_30894,N_30736,N_30514);
and U30895 (N_30895,N_30596,N_30702);
nand U30896 (N_30896,N_30560,N_30710);
and U30897 (N_30897,N_30739,N_30682);
and U30898 (N_30898,N_30625,N_30508);
xor U30899 (N_30899,N_30655,N_30516);
xnor U30900 (N_30900,N_30715,N_30530);
or U30901 (N_30901,N_30507,N_30710);
or U30902 (N_30902,N_30553,N_30649);
xnor U30903 (N_30903,N_30548,N_30584);
nand U30904 (N_30904,N_30741,N_30596);
or U30905 (N_30905,N_30670,N_30582);
and U30906 (N_30906,N_30512,N_30563);
or U30907 (N_30907,N_30604,N_30665);
nand U30908 (N_30908,N_30545,N_30622);
or U30909 (N_30909,N_30660,N_30573);
xnor U30910 (N_30910,N_30667,N_30734);
xnor U30911 (N_30911,N_30747,N_30514);
xor U30912 (N_30912,N_30604,N_30577);
or U30913 (N_30913,N_30621,N_30569);
nor U30914 (N_30914,N_30725,N_30628);
and U30915 (N_30915,N_30703,N_30579);
and U30916 (N_30916,N_30685,N_30674);
and U30917 (N_30917,N_30700,N_30505);
nor U30918 (N_30918,N_30629,N_30681);
xnor U30919 (N_30919,N_30678,N_30545);
and U30920 (N_30920,N_30647,N_30723);
or U30921 (N_30921,N_30732,N_30675);
xor U30922 (N_30922,N_30647,N_30712);
or U30923 (N_30923,N_30702,N_30699);
or U30924 (N_30924,N_30543,N_30555);
nor U30925 (N_30925,N_30593,N_30514);
nand U30926 (N_30926,N_30739,N_30626);
nand U30927 (N_30927,N_30710,N_30723);
nor U30928 (N_30928,N_30744,N_30642);
xnor U30929 (N_30929,N_30728,N_30629);
or U30930 (N_30930,N_30586,N_30510);
xor U30931 (N_30931,N_30598,N_30668);
xnor U30932 (N_30932,N_30508,N_30564);
xnor U30933 (N_30933,N_30590,N_30507);
nand U30934 (N_30934,N_30536,N_30713);
nor U30935 (N_30935,N_30721,N_30582);
nor U30936 (N_30936,N_30625,N_30667);
xnor U30937 (N_30937,N_30699,N_30605);
xnor U30938 (N_30938,N_30604,N_30588);
and U30939 (N_30939,N_30551,N_30711);
and U30940 (N_30940,N_30651,N_30620);
xnor U30941 (N_30941,N_30549,N_30503);
nand U30942 (N_30942,N_30554,N_30690);
nor U30943 (N_30943,N_30741,N_30529);
and U30944 (N_30944,N_30646,N_30635);
or U30945 (N_30945,N_30675,N_30694);
nor U30946 (N_30946,N_30506,N_30707);
nor U30947 (N_30947,N_30539,N_30509);
and U30948 (N_30948,N_30599,N_30549);
or U30949 (N_30949,N_30735,N_30722);
nand U30950 (N_30950,N_30541,N_30662);
nand U30951 (N_30951,N_30639,N_30609);
nor U30952 (N_30952,N_30677,N_30610);
nand U30953 (N_30953,N_30639,N_30680);
nand U30954 (N_30954,N_30511,N_30742);
nor U30955 (N_30955,N_30560,N_30725);
nand U30956 (N_30956,N_30524,N_30609);
or U30957 (N_30957,N_30654,N_30556);
nor U30958 (N_30958,N_30510,N_30729);
and U30959 (N_30959,N_30612,N_30606);
xor U30960 (N_30960,N_30695,N_30654);
nand U30961 (N_30961,N_30723,N_30517);
xor U30962 (N_30962,N_30685,N_30621);
and U30963 (N_30963,N_30679,N_30634);
or U30964 (N_30964,N_30525,N_30672);
nand U30965 (N_30965,N_30749,N_30539);
or U30966 (N_30966,N_30696,N_30612);
nor U30967 (N_30967,N_30591,N_30708);
or U30968 (N_30968,N_30704,N_30630);
nor U30969 (N_30969,N_30533,N_30725);
xor U30970 (N_30970,N_30556,N_30557);
nand U30971 (N_30971,N_30724,N_30613);
nand U30972 (N_30972,N_30566,N_30516);
xnor U30973 (N_30973,N_30634,N_30698);
nand U30974 (N_30974,N_30736,N_30595);
or U30975 (N_30975,N_30517,N_30667);
nor U30976 (N_30976,N_30547,N_30534);
nor U30977 (N_30977,N_30685,N_30520);
and U30978 (N_30978,N_30679,N_30630);
and U30979 (N_30979,N_30723,N_30539);
xor U30980 (N_30980,N_30604,N_30531);
and U30981 (N_30981,N_30517,N_30525);
nand U30982 (N_30982,N_30503,N_30715);
nand U30983 (N_30983,N_30717,N_30523);
nor U30984 (N_30984,N_30747,N_30550);
or U30985 (N_30985,N_30628,N_30546);
nand U30986 (N_30986,N_30562,N_30551);
nor U30987 (N_30987,N_30748,N_30631);
or U30988 (N_30988,N_30713,N_30603);
xor U30989 (N_30989,N_30713,N_30680);
nand U30990 (N_30990,N_30690,N_30658);
nand U30991 (N_30991,N_30579,N_30608);
xor U30992 (N_30992,N_30548,N_30541);
or U30993 (N_30993,N_30582,N_30704);
nand U30994 (N_30994,N_30651,N_30632);
nand U30995 (N_30995,N_30576,N_30549);
xnor U30996 (N_30996,N_30568,N_30601);
xnor U30997 (N_30997,N_30726,N_30688);
nand U30998 (N_30998,N_30564,N_30725);
and U30999 (N_30999,N_30609,N_30528);
nor U31000 (N_31000,N_30995,N_30941);
nor U31001 (N_31001,N_30786,N_30817);
nand U31002 (N_31002,N_30963,N_30989);
or U31003 (N_31003,N_30801,N_30916);
or U31004 (N_31004,N_30901,N_30818);
or U31005 (N_31005,N_30803,N_30954);
and U31006 (N_31006,N_30829,N_30885);
nor U31007 (N_31007,N_30971,N_30940);
nand U31008 (N_31008,N_30925,N_30804);
nor U31009 (N_31009,N_30810,N_30837);
xor U31010 (N_31010,N_30765,N_30951);
nor U31011 (N_31011,N_30939,N_30929);
xnor U31012 (N_31012,N_30996,N_30898);
or U31013 (N_31013,N_30998,N_30934);
nor U31014 (N_31014,N_30864,N_30968);
nor U31015 (N_31015,N_30766,N_30798);
and U31016 (N_31016,N_30838,N_30792);
xor U31017 (N_31017,N_30896,N_30947);
or U31018 (N_31018,N_30815,N_30867);
nor U31019 (N_31019,N_30774,N_30877);
nor U31020 (N_31020,N_30851,N_30983);
or U31021 (N_31021,N_30930,N_30843);
nor U31022 (N_31022,N_30936,N_30831);
xnor U31023 (N_31023,N_30790,N_30993);
xnor U31024 (N_31024,N_30952,N_30924);
nor U31025 (N_31025,N_30911,N_30844);
nor U31026 (N_31026,N_30763,N_30797);
nand U31027 (N_31027,N_30891,N_30835);
and U31028 (N_31028,N_30791,N_30985);
and U31029 (N_31029,N_30894,N_30767);
xnor U31030 (N_31030,N_30895,N_30781);
and U31031 (N_31031,N_30892,N_30955);
xor U31032 (N_31032,N_30990,N_30872);
nand U31033 (N_31033,N_30874,N_30821);
or U31034 (N_31034,N_30771,N_30958);
or U31035 (N_31035,N_30943,N_30977);
nand U31036 (N_31036,N_30863,N_30793);
nor U31037 (N_31037,N_30976,N_30762);
or U31038 (N_31038,N_30927,N_30915);
and U31039 (N_31039,N_30773,N_30845);
or U31040 (N_31040,N_30782,N_30753);
and U31041 (N_31041,N_30922,N_30827);
or U31042 (N_31042,N_30808,N_30964);
nor U31043 (N_31043,N_30897,N_30812);
and U31044 (N_31044,N_30910,N_30862);
or U31045 (N_31045,N_30933,N_30778);
or U31046 (N_31046,N_30884,N_30984);
and U31047 (N_31047,N_30972,N_30914);
and U31048 (N_31048,N_30973,N_30881);
xor U31049 (N_31049,N_30866,N_30776);
xnor U31050 (N_31050,N_30772,N_30834);
and U31051 (N_31051,N_30823,N_30883);
nand U31052 (N_31052,N_30919,N_30775);
xor U31053 (N_31053,N_30979,N_30967);
and U31054 (N_31054,N_30893,N_30852);
or U31055 (N_31055,N_30926,N_30928);
xor U31056 (N_31056,N_30820,N_30899);
xnor U31057 (N_31057,N_30799,N_30950);
and U31058 (N_31058,N_30906,N_30856);
or U31059 (N_31059,N_30917,N_30980);
nor U31060 (N_31060,N_30873,N_30994);
and U31061 (N_31061,N_30949,N_30878);
nand U31062 (N_31062,N_30758,N_30904);
nand U31063 (N_31063,N_30847,N_30900);
and U31064 (N_31064,N_30828,N_30953);
nand U31065 (N_31065,N_30854,N_30978);
xor U31066 (N_31066,N_30777,N_30935);
nor U31067 (N_31067,N_30859,N_30987);
and U31068 (N_31068,N_30841,N_30944);
xnor U31069 (N_31069,N_30846,N_30870);
nand U31070 (N_31070,N_30921,N_30764);
xnor U31071 (N_31071,N_30751,N_30920);
nor U31072 (N_31072,N_30875,N_30805);
and U31073 (N_31073,N_30768,N_30965);
or U31074 (N_31074,N_30902,N_30796);
and U31075 (N_31075,N_30752,N_30962);
nor U31076 (N_31076,N_30975,N_30876);
xor U31077 (N_31077,N_30853,N_30986);
xnor U31078 (N_31078,N_30890,N_30833);
xnor U31079 (N_31079,N_30869,N_30755);
nor U31080 (N_31080,N_30966,N_30988);
or U31081 (N_31081,N_30991,N_30750);
nor U31082 (N_31082,N_30780,N_30819);
or U31083 (N_31083,N_30840,N_30825);
or U31084 (N_31084,N_30759,N_30889);
nand U31085 (N_31085,N_30842,N_30932);
and U31086 (N_31086,N_30788,N_30826);
nand U31087 (N_31087,N_30787,N_30938);
nor U31088 (N_31088,N_30981,N_30999);
nor U31089 (N_31089,N_30769,N_30830);
xor U31090 (N_31090,N_30931,N_30970);
nand U31091 (N_31091,N_30946,N_30886);
nor U31092 (N_31092,N_30770,N_30784);
nor U31093 (N_31093,N_30905,N_30942);
xor U31094 (N_31094,N_30945,N_30809);
and U31095 (N_31095,N_30909,N_30822);
and U31096 (N_31096,N_30802,N_30888);
xnor U31097 (N_31097,N_30760,N_30879);
and U31098 (N_31098,N_30789,N_30868);
nand U31099 (N_31099,N_30779,N_30807);
xor U31100 (N_31100,N_30957,N_30754);
nand U31101 (N_31101,N_30813,N_30855);
nor U31102 (N_31102,N_30857,N_30961);
xnor U31103 (N_31103,N_30811,N_30858);
xnor U31104 (N_31104,N_30907,N_30997);
nand U31105 (N_31105,N_30887,N_30956);
and U31106 (N_31106,N_30860,N_30913);
nand U31107 (N_31107,N_30795,N_30912);
nand U31108 (N_31108,N_30918,N_30923);
nand U31109 (N_31109,N_30850,N_30849);
xor U31110 (N_31110,N_30783,N_30836);
nand U31111 (N_31111,N_30974,N_30882);
and U31112 (N_31112,N_30848,N_30756);
xor U31113 (N_31113,N_30880,N_30992);
xor U31114 (N_31114,N_30937,N_30982);
nor U31115 (N_31115,N_30757,N_30871);
or U31116 (N_31116,N_30959,N_30948);
or U31117 (N_31117,N_30832,N_30800);
and U31118 (N_31118,N_30960,N_30785);
and U31119 (N_31119,N_30794,N_30806);
nand U31120 (N_31120,N_30761,N_30861);
and U31121 (N_31121,N_30865,N_30814);
nand U31122 (N_31122,N_30824,N_30908);
nor U31123 (N_31123,N_30903,N_30816);
or U31124 (N_31124,N_30839,N_30969);
or U31125 (N_31125,N_30991,N_30864);
or U31126 (N_31126,N_30844,N_30878);
xnor U31127 (N_31127,N_30826,N_30829);
xor U31128 (N_31128,N_30825,N_30891);
nor U31129 (N_31129,N_30918,N_30959);
xnor U31130 (N_31130,N_30951,N_30953);
or U31131 (N_31131,N_30944,N_30755);
xor U31132 (N_31132,N_30982,N_30903);
xor U31133 (N_31133,N_30901,N_30935);
xor U31134 (N_31134,N_30858,N_30797);
and U31135 (N_31135,N_30852,N_30780);
or U31136 (N_31136,N_30974,N_30887);
and U31137 (N_31137,N_30868,N_30986);
xnor U31138 (N_31138,N_30787,N_30933);
or U31139 (N_31139,N_30862,N_30824);
and U31140 (N_31140,N_30805,N_30992);
xnor U31141 (N_31141,N_30964,N_30849);
xnor U31142 (N_31142,N_30794,N_30859);
nand U31143 (N_31143,N_30771,N_30794);
xor U31144 (N_31144,N_30901,N_30921);
and U31145 (N_31145,N_30918,N_30895);
xnor U31146 (N_31146,N_30878,N_30975);
or U31147 (N_31147,N_30857,N_30856);
xnor U31148 (N_31148,N_30825,N_30760);
xor U31149 (N_31149,N_30980,N_30767);
xnor U31150 (N_31150,N_30955,N_30942);
xor U31151 (N_31151,N_30935,N_30987);
nand U31152 (N_31152,N_30990,N_30798);
nor U31153 (N_31153,N_30880,N_30983);
or U31154 (N_31154,N_30916,N_30833);
xor U31155 (N_31155,N_30865,N_30970);
nand U31156 (N_31156,N_30976,N_30922);
or U31157 (N_31157,N_30991,N_30840);
xnor U31158 (N_31158,N_30996,N_30923);
xnor U31159 (N_31159,N_30970,N_30765);
nand U31160 (N_31160,N_30787,N_30822);
nor U31161 (N_31161,N_30971,N_30847);
nor U31162 (N_31162,N_30854,N_30982);
xnor U31163 (N_31163,N_30972,N_30913);
or U31164 (N_31164,N_30768,N_30876);
nor U31165 (N_31165,N_30837,N_30755);
or U31166 (N_31166,N_30923,N_30836);
and U31167 (N_31167,N_30926,N_30809);
or U31168 (N_31168,N_30819,N_30859);
nand U31169 (N_31169,N_30787,N_30920);
nor U31170 (N_31170,N_30834,N_30980);
and U31171 (N_31171,N_30974,N_30912);
xnor U31172 (N_31172,N_30786,N_30852);
nand U31173 (N_31173,N_30829,N_30776);
nor U31174 (N_31174,N_30796,N_30895);
or U31175 (N_31175,N_30824,N_30777);
xor U31176 (N_31176,N_30934,N_30865);
nand U31177 (N_31177,N_30965,N_30834);
nand U31178 (N_31178,N_30812,N_30753);
nor U31179 (N_31179,N_30959,N_30977);
xnor U31180 (N_31180,N_30913,N_30878);
and U31181 (N_31181,N_30886,N_30914);
and U31182 (N_31182,N_30846,N_30886);
or U31183 (N_31183,N_30796,N_30991);
nor U31184 (N_31184,N_30810,N_30935);
and U31185 (N_31185,N_30776,N_30996);
nor U31186 (N_31186,N_30861,N_30803);
nand U31187 (N_31187,N_30815,N_30819);
or U31188 (N_31188,N_30872,N_30850);
nand U31189 (N_31189,N_30801,N_30789);
xor U31190 (N_31190,N_30910,N_30917);
or U31191 (N_31191,N_30762,N_30809);
nand U31192 (N_31192,N_30946,N_30794);
nor U31193 (N_31193,N_30931,N_30865);
or U31194 (N_31194,N_30904,N_30888);
nand U31195 (N_31195,N_30778,N_30849);
xnor U31196 (N_31196,N_30951,N_30924);
nand U31197 (N_31197,N_30917,N_30973);
nand U31198 (N_31198,N_30878,N_30972);
nor U31199 (N_31199,N_30809,N_30980);
nor U31200 (N_31200,N_30767,N_30780);
nor U31201 (N_31201,N_30870,N_30834);
nand U31202 (N_31202,N_30971,N_30844);
nand U31203 (N_31203,N_30836,N_30828);
and U31204 (N_31204,N_30887,N_30996);
xor U31205 (N_31205,N_30751,N_30836);
and U31206 (N_31206,N_30782,N_30932);
or U31207 (N_31207,N_30808,N_30770);
xor U31208 (N_31208,N_30937,N_30944);
nor U31209 (N_31209,N_30845,N_30866);
nor U31210 (N_31210,N_30858,N_30919);
or U31211 (N_31211,N_30929,N_30951);
xnor U31212 (N_31212,N_30918,N_30789);
and U31213 (N_31213,N_30962,N_30862);
nor U31214 (N_31214,N_30941,N_30967);
nand U31215 (N_31215,N_30844,N_30760);
nor U31216 (N_31216,N_30791,N_30995);
nand U31217 (N_31217,N_30776,N_30784);
or U31218 (N_31218,N_30839,N_30922);
and U31219 (N_31219,N_30885,N_30763);
nor U31220 (N_31220,N_30756,N_30804);
xor U31221 (N_31221,N_30895,N_30751);
xnor U31222 (N_31222,N_30933,N_30801);
nor U31223 (N_31223,N_30902,N_30855);
nand U31224 (N_31224,N_30998,N_30837);
or U31225 (N_31225,N_30809,N_30815);
and U31226 (N_31226,N_30943,N_30771);
nor U31227 (N_31227,N_30795,N_30897);
xor U31228 (N_31228,N_30999,N_30930);
xor U31229 (N_31229,N_30996,N_30952);
xor U31230 (N_31230,N_30758,N_30921);
nor U31231 (N_31231,N_30982,N_30827);
or U31232 (N_31232,N_30947,N_30902);
nand U31233 (N_31233,N_30914,N_30980);
xor U31234 (N_31234,N_30949,N_30769);
nand U31235 (N_31235,N_30976,N_30995);
and U31236 (N_31236,N_30763,N_30857);
or U31237 (N_31237,N_30856,N_30959);
xnor U31238 (N_31238,N_30828,N_30921);
and U31239 (N_31239,N_30762,N_30926);
and U31240 (N_31240,N_30785,N_30762);
or U31241 (N_31241,N_30984,N_30944);
and U31242 (N_31242,N_30781,N_30885);
xnor U31243 (N_31243,N_30967,N_30884);
nor U31244 (N_31244,N_30821,N_30991);
nor U31245 (N_31245,N_30822,N_30936);
or U31246 (N_31246,N_30877,N_30908);
nor U31247 (N_31247,N_30809,N_30935);
nor U31248 (N_31248,N_30934,N_30761);
nor U31249 (N_31249,N_30930,N_30791);
and U31250 (N_31250,N_31042,N_31208);
and U31251 (N_31251,N_31061,N_31196);
nor U31252 (N_31252,N_31011,N_31136);
and U31253 (N_31253,N_31179,N_31166);
xnor U31254 (N_31254,N_31048,N_31160);
xnor U31255 (N_31255,N_31059,N_31038);
or U31256 (N_31256,N_31068,N_31033);
nand U31257 (N_31257,N_31095,N_31105);
or U31258 (N_31258,N_31226,N_31007);
or U31259 (N_31259,N_31125,N_31178);
and U31260 (N_31260,N_31213,N_31232);
xor U31261 (N_31261,N_31171,N_31220);
nand U31262 (N_31262,N_31066,N_31015);
nor U31263 (N_31263,N_31083,N_31205);
nand U31264 (N_31264,N_31106,N_31189);
nor U31265 (N_31265,N_31089,N_31122);
nand U31266 (N_31266,N_31004,N_31096);
nor U31267 (N_31267,N_31147,N_31151);
and U31268 (N_31268,N_31010,N_31020);
or U31269 (N_31269,N_31234,N_31139);
nand U31270 (N_31270,N_31037,N_31173);
xnor U31271 (N_31271,N_31019,N_31014);
nand U31272 (N_31272,N_31193,N_31135);
nand U31273 (N_31273,N_31243,N_31009);
and U31274 (N_31274,N_31070,N_31204);
or U31275 (N_31275,N_31176,N_31163);
or U31276 (N_31276,N_31215,N_31023);
or U31277 (N_31277,N_31209,N_31127);
or U31278 (N_31278,N_31236,N_31081);
and U31279 (N_31279,N_31067,N_31210);
or U31280 (N_31280,N_31074,N_31118);
and U31281 (N_31281,N_31041,N_31058);
nand U31282 (N_31282,N_31072,N_31156);
nor U31283 (N_31283,N_31113,N_31085);
or U31284 (N_31284,N_31060,N_31018);
nand U31285 (N_31285,N_31143,N_31071);
nand U31286 (N_31286,N_31036,N_31065);
and U31287 (N_31287,N_31076,N_31190);
xor U31288 (N_31288,N_31195,N_31031);
xnor U31289 (N_31289,N_31230,N_31245);
nor U31290 (N_31290,N_31152,N_31248);
nor U31291 (N_31291,N_31141,N_31172);
or U31292 (N_31292,N_31055,N_31078);
and U31293 (N_31293,N_31246,N_31027);
and U31294 (N_31294,N_31093,N_31006);
nand U31295 (N_31295,N_31169,N_31188);
or U31296 (N_31296,N_31221,N_31064);
nand U31297 (N_31297,N_31170,N_31021);
nor U31298 (N_31298,N_31040,N_31079);
xor U31299 (N_31299,N_31003,N_31137);
or U31300 (N_31300,N_31167,N_31133);
and U31301 (N_31301,N_31235,N_31244);
nor U31302 (N_31302,N_31107,N_31063);
or U31303 (N_31303,N_31116,N_31239);
nand U31304 (N_31304,N_31092,N_31029);
xor U31305 (N_31305,N_31108,N_31161);
nand U31306 (N_31306,N_31197,N_31043);
nand U31307 (N_31307,N_31026,N_31094);
nor U31308 (N_31308,N_31087,N_31162);
or U31309 (N_31309,N_31191,N_31102);
and U31310 (N_31310,N_31025,N_31168);
nor U31311 (N_31311,N_31097,N_31002);
nand U31312 (N_31312,N_31073,N_31185);
or U31313 (N_31313,N_31080,N_31211);
nor U31314 (N_31314,N_31000,N_31053);
xor U31315 (N_31315,N_31242,N_31099);
nand U31316 (N_31316,N_31201,N_31240);
xnor U31317 (N_31317,N_31184,N_31198);
nand U31318 (N_31318,N_31249,N_31199);
and U31319 (N_31319,N_31192,N_31138);
xor U31320 (N_31320,N_31123,N_31049);
xnor U31321 (N_31321,N_31008,N_31030);
and U31322 (N_31322,N_31149,N_31181);
nor U31323 (N_31323,N_31069,N_31154);
nor U31324 (N_31324,N_31104,N_31229);
xnor U31325 (N_31325,N_31134,N_31117);
nand U31326 (N_31326,N_31088,N_31109);
nand U31327 (N_31327,N_31005,N_31180);
or U31328 (N_31328,N_31091,N_31022);
xor U31329 (N_31329,N_31124,N_31032);
or U31330 (N_31330,N_31062,N_31013);
nor U31331 (N_31331,N_31050,N_31155);
nor U31332 (N_31332,N_31084,N_31121);
or U31333 (N_31333,N_31129,N_31206);
and U31334 (N_31334,N_31142,N_31183);
and U31335 (N_31335,N_31132,N_31207);
xnor U31336 (N_31336,N_31148,N_31114);
xor U31337 (N_31337,N_31144,N_31233);
xor U31338 (N_31338,N_31186,N_31140);
or U31339 (N_31339,N_31238,N_31187);
nor U31340 (N_31340,N_31057,N_31086);
or U31341 (N_31341,N_31214,N_31247);
and U31342 (N_31342,N_31090,N_31024);
and U31343 (N_31343,N_31054,N_31034);
nand U31344 (N_31344,N_31110,N_31146);
and U31345 (N_31345,N_31120,N_31111);
or U31346 (N_31346,N_31101,N_31212);
nor U31347 (N_31347,N_31159,N_31227);
or U31348 (N_31348,N_31241,N_31044);
or U31349 (N_31349,N_31001,N_31115);
and U31350 (N_31350,N_31222,N_31174);
and U31351 (N_31351,N_31035,N_31175);
xor U31352 (N_31352,N_31158,N_31177);
or U31353 (N_31353,N_31218,N_31228);
or U31354 (N_31354,N_31051,N_31119);
nand U31355 (N_31355,N_31103,N_31164);
and U31356 (N_31356,N_31082,N_31165);
xor U31357 (N_31357,N_31012,N_31052);
nand U31358 (N_31358,N_31047,N_31077);
and U31359 (N_31359,N_31157,N_31126);
nand U31360 (N_31360,N_31224,N_31145);
nor U31361 (N_31361,N_31225,N_31131);
nand U31362 (N_31362,N_31231,N_31039);
xnor U31363 (N_31363,N_31216,N_31182);
or U31364 (N_31364,N_31046,N_31045);
and U31365 (N_31365,N_31219,N_31075);
xnor U31366 (N_31366,N_31202,N_31130);
nor U31367 (N_31367,N_31203,N_31016);
nor U31368 (N_31368,N_31153,N_31223);
or U31369 (N_31369,N_31098,N_31056);
xnor U31370 (N_31370,N_31100,N_31200);
xnor U31371 (N_31371,N_31028,N_31217);
nor U31372 (N_31372,N_31017,N_31194);
or U31373 (N_31373,N_31128,N_31237);
nor U31374 (N_31374,N_31150,N_31112);
or U31375 (N_31375,N_31113,N_31173);
or U31376 (N_31376,N_31180,N_31085);
and U31377 (N_31377,N_31106,N_31036);
nor U31378 (N_31378,N_31126,N_31115);
or U31379 (N_31379,N_31084,N_31182);
nor U31380 (N_31380,N_31141,N_31137);
or U31381 (N_31381,N_31107,N_31188);
or U31382 (N_31382,N_31165,N_31075);
and U31383 (N_31383,N_31067,N_31118);
nor U31384 (N_31384,N_31134,N_31213);
xnor U31385 (N_31385,N_31142,N_31154);
xnor U31386 (N_31386,N_31093,N_31242);
and U31387 (N_31387,N_31165,N_31112);
and U31388 (N_31388,N_31041,N_31230);
xnor U31389 (N_31389,N_31015,N_31105);
xor U31390 (N_31390,N_31062,N_31143);
nor U31391 (N_31391,N_31227,N_31232);
and U31392 (N_31392,N_31052,N_31163);
nand U31393 (N_31393,N_31043,N_31116);
nor U31394 (N_31394,N_31005,N_31217);
and U31395 (N_31395,N_31248,N_31162);
xor U31396 (N_31396,N_31246,N_31099);
or U31397 (N_31397,N_31122,N_31037);
and U31398 (N_31398,N_31027,N_31240);
nor U31399 (N_31399,N_31235,N_31144);
nor U31400 (N_31400,N_31115,N_31086);
nand U31401 (N_31401,N_31109,N_31103);
and U31402 (N_31402,N_31146,N_31207);
nand U31403 (N_31403,N_31118,N_31026);
or U31404 (N_31404,N_31079,N_31022);
nand U31405 (N_31405,N_31087,N_31077);
xnor U31406 (N_31406,N_31209,N_31053);
xor U31407 (N_31407,N_31030,N_31052);
xor U31408 (N_31408,N_31115,N_31152);
or U31409 (N_31409,N_31088,N_31076);
nand U31410 (N_31410,N_31178,N_31232);
nor U31411 (N_31411,N_31247,N_31223);
nand U31412 (N_31412,N_31109,N_31019);
or U31413 (N_31413,N_31134,N_31177);
nand U31414 (N_31414,N_31155,N_31239);
or U31415 (N_31415,N_31101,N_31180);
xnor U31416 (N_31416,N_31226,N_31124);
xnor U31417 (N_31417,N_31247,N_31189);
or U31418 (N_31418,N_31215,N_31011);
nor U31419 (N_31419,N_31092,N_31051);
nand U31420 (N_31420,N_31088,N_31057);
or U31421 (N_31421,N_31033,N_31169);
or U31422 (N_31422,N_31233,N_31064);
nor U31423 (N_31423,N_31185,N_31147);
nand U31424 (N_31424,N_31201,N_31185);
nand U31425 (N_31425,N_31012,N_31186);
nand U31426 (N_31426,N_31035,N_31190);
xnor U31427 (N_31427,N_31066,N_31100);
nand U31428 (N_31428,N_31223,N_31208);
and U31429 (N_31429,N_31001,N_31219);
and U31430 (N_31430,N_31053,N_31105);
and U31431 (N_31431,N_31045,N_31172);
xnor U31432 (N_31432,N_31109,N_31091);
xor U31433 (N_31433,N_31089,N_31113);
or U31434 (N_31434,N_31203,N_31218);
nor U31435 (N_31435,N_31082,N_31177);
and U31436 (N_31436,N_31022,N_31243);
nor U31437 (N_31437,N_31234,N_31209);
xor U31438 (N_31438,N_31232,N_31140);
xor U31439 (N_31439,N_31006,N_31235);
and U31440 (N_31440,N_31101,N_31003);
or U31441 (N_31441,N_31152,N_31064);
and U31442 (N_31442,N_31045,N_31025);
or U31443 (N_31443,N_31084,N_31234);
xor U31444 (N_31444,N_31205,N_31154);
and U31445 (N_31445,N_31095,N_31135);
nand U31446 (N_31446,N_31230,N_31009);
nor U31447 (N_31447,N_31001,N_31245);
or U31448 (N_31448,N_31006,N_31107);
or U31449 (N_31449,N_31181,N_31038);
xor U31450 (N_31450,N_31037,N_31083);
nand U31451 (N_31451,N_31212,N_31079);
xnor U31452 (N_31452,N_31134,N_31244);
nor U31453 (N_31453,N_31235,N_31193);
nand U31454 (N_31454,N_31051,N_31018);
or U31455 (N_31455,N_31174,N_31054);
or U31456 (N_31456,N_31137,N_31189);
nand U31457 (N_31457,N_31194,N_31130);
and U31458 (N_31458,N_31009,N_31155);
nor U31459 (N_31459,N_31169,N_31001);
nor U31460 (N_31460,N_31216,N_31143);
nand U31461 (N_31461,N_31129,N_31220);
nand U31462 (N_31462,N_31234,N_31157);
nand U31463 (N_31463,N_31085,N_31083);
xor U31464 (N_31464,N_31047,N_31200);
or U31465 (N_31465,N_31234,N_31078);
nor U31466 (N_31466,N_31121,N_31222);
xor U31467 (N_31467,N_31069,N_31041);
or U31468 (N_31468,N_31060,N_31231);
nand U31469 (N_31469,N_31020,N_31012);
nor U31470 (N_31470,N_31024,N_31083);
xnor U31471 (N_31471,N_31230,N_31248);
xor U31472 (N_31472,N_31027,N_31029);
or U31473 (N_31473,N_31114,N_31222);
and U31474 (N_31474,N_31157,N_31147);
nand U31475 (N_31475,N_31123,N_31116);
or U31476 (N_31476,N_31112,N_31058);
xnor U31477 (N_31477,N_31151,N_31169);
nand U31478 (N_31478,N_31114,N_31246);
xnor U31479 (N_31479,N_31098,N_31153);
nor U31480 (N_31480,N_31055,N_31104);
nor U31481 (N_31481,N_31238,N_31037);
or U31482 (N_31482,N_31032,N_31249);
xor U31483 (N_31483,N_31166,N_31018);
nor U31484 (N_31484,N_31028,N_31006);
nand U31485 (N_31485,N_31142,N_31033);
nor U31486 (N_31486,N_31024,N_31201);
xor U31487 (N_31487,N_31039,N_31073);
or U31488 (N_31488,N_31034,N_31008);
or U31489 (N_31489,N_31010,N_31030);
xor U31490 (N_31490,N_31137,N_31112);
nand U31491 (N_31491,N_31185,N_31232);
nand U31492 (N_31492,N_31098,N_31245);
nand U31493 (N_31493,N_31224,N_31226);
nand U31494 (N_31494,N_31118,N_31247);
nor U31495 (N_31495,N_31079,N_31058);
nor U31496 (N_31496,N_31104,N_31048);
nand U31497 (N_31497,N_31071,N_31153);
or U31498 (N_31498,N_31044,N_31161);
and U31499 (N_31499,N_31118,N_31021);
nand U31500 (N_31500,N_31377,N_31486);
xor U31501 (N_31501,N_31307,N_31360);
and U31502 (N_31502,N_31272,N_31294);
nor U31503 (N_31503,N_31278,N_31257);
or U31504 (N_31504,N_31372,N_31286);
and U31505 (N_31505,N_31346,N_31491);
nor U31506 (N_31506,N_31270,N_31354);
nand U31507 (N_31507,N_31406,N_31471);
xor U31508 (N_31508,N_31284,N_31323);
xor U31509 (N_31509,N_31321,N_31364);
or U31510 (N_31510,N_31253,N_31319);
or U31511 (N_31511,N_31483,N_31317);
nand U31512 (N_31512,N_31403,N_31353);
or U31513 (N_31513,N_31350,N_31448);
nand U31514 (N_31514,N_31488,N_31477);
xor U31515 (N_31515,N_31256,N_31260);
nor U31516 (N_31516,N_31454,N_31297);
nand U31517 (N_31517,N_31280,N_31309);
nor U31518 (N_31518,N_31250,N_31274);
or U31519 (N_31519,N_31409,N_31410);
nor U31520 (N_31520,N_31443,N_31262);
nor U31521 (N_31521,N_31355,N_31402);
and U31522 (N_31522,N_31283,N_31405);
xnor U31523 (N_31523,N_31332,N_31484);
and U31524 (N_31524,N_31322,N_31324);
and U31525 (N_31525,N_31418,N_31386);
and U31526 (N_31526,N_31493,N_31387);
or U31527 (N_31527,N_31389,N_31475);
or U31528 (N_31528,N_31441,N_31325);
xor U31529 (N_31529,N_31255,N_31427);
nand U31530 (N_31530,N_31339,N_31492);
nand U31531 (N_31531,N_31466,N_31430);
nor U31532 (N_31532,N_31445,N_31335);
nor U31533 (N_31533,N_31267,N_31370);
xnor U31534 (N_31534,N_31293,N_31407);
and U31535 (N_31535,N_31404,N_31398);
nand U31536 (N_31536,N_31397,N_31380);
xnor U31537 (N_31537,N_31452,N_31392);
and U31538 (N_31538,N_31334,N_31295);
or U31539 (N_31539,N_31450,N_31391);
and U31540 (N_31540,N_31428,N_31374);
nor U31541 (N_31541,N_31433,N_31490);
nor U31542 (N_31542,N_31436,N_31447);
or U31543 (N_31543,N_31331,N_31328);
and U31544 (N_31544,N_31282,N_31435);
nor U31545 (N_31545,N_31381,N_31432);
nand U31546 (N_31546,N_31358,N_31489);
and U31547 (N_31547,N_31470,N_31480);
nor U31548 (N_31548,N_31473,N_31365);
nor U31549 (N_31549,N_31393,N_31340);
and U31550 (N_31550,N_31288,N_31485);
nand U31551 (N_31551,N_31499,N_31251);
or U31552 (N_31552,N_31261,N_31465);
or U31553 (N_31553,N_31349,N_31361);
or U31554 (N_31554,N_31498,N_31275);
and U31555 (N_31555,N_31474,N_31449);
or U31556 (N_31556,N_31273,N_31451);
or U31557 (N_31557,N_31412,N_31347);
or U31558 (N_31558,N_31265,N_31298);
nor U31559 (N_31559,N_31378,N_31287);
nand U31560 (N_31560,N_31312,N_31400);
or U31561 (N_31561,N_31442,N_31399);
or U31562 (N_31562,N_31276,N_31422);
nor U31563 (N_31563,N_31424,N_31254);
or U31564 (N_31564,N_31396,N_31411);
and U31565 (N_31565,N_31496,N_31338);
or U31566 (N_31566,N_31277,N_31415);
and U31567 (N_31567,N_31423,N_31444);
nor U31568 (N_31568,N_31458,N_31421);
nand U31569 (N_31569,N_31476,N_31303);
or U31570 (N_31570,N_31314,N_31356);
nand U31571 (N_31571,N_31494,N_31271);
nor U31572 (N_31572,N_31413,N_31497);
or U31573 (N_31573,N_31371,N_31281);
nor U31574 (N_31574,N_31495,N_31351);
xnor U31575 (N_31575,N_31388,N_31367);
or U31576 (N_31576,N_31279,N_31459);
nor U31577 (N_31577,N_31320,N_31362);
and U31578 (N_31578,N_31363,N_31299);
xnor U31579 (N_31579,N_31327,N_31359);
nand U31580 (N_31580,N_31468,N_31341);
nand U31581 (N_31581,N_31292,N_31268);
or U31582 (N_31582,N_31382,N_31395);
or U31583 (N_31583,N_31414,N_31481);
and U31584 (N_31584,N_31318,N_31330);
or U31585 (N_31585,N_31383,N_31376);
xnor U31586 (N_31586,N_31357,N_31315);
nand U31587 (N_31587,N_31302,N_31345);
or U31588 (N_31588,N_31310,N_31416);
or U31589 (N_31589,N_31462,N_31301);
xnor U31590 (N_31590,N_31308,N_31326);
or U31591 (N_31591,N_31478,N_31296);
and U31592 (N_31592,N_31469,N_31329);
and U31593 (N_31593,N_31384,N_31348);
nand U31594 (N_31594,N_31482,N_31344);
nand U31595 (N_31595,N_31290,N_31460);
nand U31596 (N_31596,N_31291,N_31439);
and U31597 (N_31597,N_31305,N_31426);
or U31598 (N_31598,N_31479,N_31419);
and U31599 (N_31599,N_31438,N_31263);
xnor U31600 (N_31600,N_31456,N_31368);
nand U31601 (N_31601,N_31420,N_31463);
xnor U31602 (N_31602,N_31311,N_31313);
xnor U31603 (N_31603,N_31289,N_31455);
nor U31604 (N_31604,N_31457,N_31342);
or U31605 (N_31605,N_31269,N_31304);
and U31606 (N_31606,N_31472,N_31461);
nor U31607 (N_31607,N_31352,N_31467);
nor U31608 (N_31608,N_31259,N_31366);
or U31609 (N_31609,N_31453,N_31417);
nor U31610 (N_31610,N_31431,N_31285);
nand U31611 (N_31611,N_31252,N_31401);
or U31612 (N_31612,N_31343,N_31390);
nand U31613 (N_31613,N_31337,N_31408);
xnor U31614 (N_31614,N_31437,N_31487);
xnor U31615 (N_31615,N_31306,N_31440);
or U31616 (N_31616,N_31385,N_31316);
xnor U31617 (N_31617,N_31266,N_31394);
nor U31618 (N_31618,N_31425,N_31375);
and U31619 (N_31619,N_31300,N_31369);
nand U31620 (N_31620,N_31258,N_31464);
and U31621 (N_31621,N_31264,N_31446);
xor U31622 (N_31622,N_31379,N_31429);
nor U31623 (N_31623,N_31373,N_31333);
xor U31624 (N_31624,N_31336,N_31434);
or U31625 (N_31625,N_31479,N_31312);
xor U31626 (N_31626,N_31251,N_31436);
nand U31627 (N_31627,N_31269,N_31397);
and U31628 (N_31628,N_31432,N_31421);
nand U31629 (N_31629,N_31440,N_31433);
nor U31630 (N_31630,N_31256,N_31334);
nor U31631 (N_31631,N_31327,N_31367);
and U31632 (N_31632,N_31394,N_31420);
xor U31633 (N_31633,N_31344,N_31339);
nand U31634 (N_31634,N_31445,N_31375);
or U31635 (N_31635,N_31460,N_31444);
and U31636 (N_31636,N_31348,N_31415);
or U31637 (N_31637,N_31415,N_31256);
or U31638 (N_31638,N_31403,N_31271);
or U31639 (N_31639,N_31454,N_31453);
or U31640 (N_31640,N_31458,N_31278);
xnor U31641 (N_31641,N_31275,N_31353);
nor U31642 (N_31642,N_31317,N_31302);
nor U31643 (N_31643,N_31405,N_31414);
xnor U31644 (N_31644,N_31341,N_31316);
and U31645 (N_31645,N_31313,N_31350);
xnor U31646 (N_31646,N_31466,N_31351);
or U31647 (N_31647,N_31349,N_31328);
and U31648 (N_31648,N_31415,N_31319);
nand U31649 (N_31649,N_31465,N_31280);
xnor U31650 (N_31650,N_31346,N_31425);
nor U31651 (N_31651,N_31491,N_31357);
or U31652 (N_31652,N_31448,N_31453);
or U31653 (N_31653,N_31409,N_31400);
and U31654 (N_31654,N_31256,N_31402);
or U31655 (N_31655,N_31250,N_31286);
xor U31656 (N_31656,N_31329,N_31286);
or U31657 (N_31657,N_31425,N_31331);
nand U31658 (N_31658,N_31443,N_31263);
xor U31659 (N_31659,N_31252,N_31406);
nor U31660 (N_31660,N_31298,N_31308);
nor U31661 (N_31661,N_31325,N_31496);
xor U31662 (N_31662,N_31437,N_31326);
nor U31663 (N_31663,N_31446,N_31471);
or U31664 (N_31664,N_31407,N_31349);
xor U31665 (N_31665,N_31464,N_31301);
nor U31666 (N_31666,N_31479,N_31305);
or U31667 (N_31667,N_31304,N_31452);
xor U31668 (N_31668,N_31330,N_31478);
xnor U31669 (N_31669,N_31314,N_31340);
and U31670 (N_31670,N_31261,N_31459);
nor U31671 (N_31671,N_31457,N_31378);
xor U31672 (N_31672,N_31400,N_31495);
and U31673 (N_31673,N_31276,N_31274);
xor U31674 (N_31674,N_31404,N_31382);
or U31675 (N_31675,N_31273,N_31417);
nor U31676 (N_31676,N_31339,N_31283);
xor U31677 (N_31677,N_31361,N_31309);
nand U31678 (N_31678,N_31369,N_31326);
xor U31679 (N_31679,N_31426,N_31319);
nand U31680 (N_31680,N_31293,N_31289);
nand U31681 (N_31681,N_31286,N_31255);
or U31682 (N_31682,N_31483,N_31475);
nor U31683 (N_31683,N_31252,N_31446);
or U31684 (N_31684,N_31371,N_31382);
xnor U31685 (N_31685,N_31437,N_31322);
or U31686 (N_31686,N_31325,N_31482);
or U31687 (N_31687,N_31467,N_31456);
or U31688 (N_31688,N_31264,N_31477);
xnor U31689 (N_31689,N_31273,N_31331);
xnor U31690 (N_31690,N_31429,N_31263);
or U31691 (N_31691,N_31285,N_31272);
nand U31692 (N_31692,N_31406,N_31478);
and U31693 (N_31693,N_31287,N_31426);
nor U31694 (N_31694,N_31450,N_31456);
nor U31695 (N_31695,N_31477,N_31317);
xnor U31696 (N_31696,N_31260,N_31336);
nor U31697 (N_31697,N_31352,N_31278);
nor U31698 (N_31698,N_31474,N_31392);
and U31699 (N_31699,N_31390,N_31364);
or U31700 (N_31700,N_31280,N_31430);
xor U31701 (N_31701,N_31381,N_31414);
nand U31702 (N_31702,N_31357,N_31412);
or U31703 (N_31703,N_31380,N_31327);
nor U31704 (N_31704,N_31381,N_31404);
or U31705 (N_31705,N_31351,N_31473);
xor U31706 (N_31706,N_31297,N_31468);
and U31707 (N_31707,N_31431,N_31316);
nand U31708 (N_31708,N_31338,N_31398);
nand U31709 (N_31709,N_31389,N_31385);
or U31710 (N_31710,N_31452,N_31453);
nor U31711 (N_31711,N_31469,N_31269);
nand U31712 (N_31712,N_31372,N_31379);
and U31713 (N_31713,N_31393,N_31304);
xnor U31714 (N_31714,N_31335,N_31326);
or U31715 (N_31715,N_31257,N_31441);
or U31716 (N_31716,N_31315,N_31449);
or U31717 (N_31717,N_31296,N_31339);
or U31718 (N_31718,N_31264,N_31368);
and U31719 (N_31719,N_31312,N_31433);
nor U31720 (N_31720,N_31358,N_31371);
and U31721 (N_31721,N_31462,N_31386);
and U31722 (N_31722,N_31413,N_31312);
nor U31723 (N_31723,N_31388,N_31346);
nand U31724 (N_31724,N_31446,N_31341);
nor U31725 (N_31725,N_31276,N_31477);
xor U31726 (N_31726,N_31487,N_31443);
xnor U31727 (N_31727,N_31281,N_31421);
xnor U31728 (N_31728,N_31406,N_31357);
nand U31729 (N_31729,N_31415,N_31409);
or U31730 (N_31730,N_31269,N_31372);
or U31731 (N_31731,N_31483,N_31495);
or U31732 (N_31732,N_31307,N_31287);
or U31733 (N_31733,N_31433,N_31302);
nand U31734 (N_31734,N_31486,N_31361);
xnor U31735 (N_31735,N_31380,N_31418);
and U31736 (N_31736,N_31334,N_31292);
nor U31737 (N_31737,N_31291,N_31481);
nor U31738 (N_31738,N_31279,N_31351);
or U31739 (N_31739,N_31375,N_31261);
xor U31740 (N_31740,N_31386,N_31423);
nor U31741 (N_31741,N_31316,N_31416);
xor U31742 (N_31742,N_31375,N_31395);
nor U31743 (N_31743,N_31401,N_31358);
xor U31744 (N_31744,N_31332,N_31429);
xor U31745 (N_31745,N_31263,N_31333);
xnor U31746 (N_31746,N_31497,N_31451);
or U31747 (N_31747,N_31460,N_31347);
xnor U31748 (N_31748,N_31315,N_31328);
nor U31749 (N_31749,N_31473,N_31296);
xor U31750 (N_31750,N_31516,N_31748);
and U31751 (N_31751,N_31736,N_31569);
nor U31752 (N_31752,N_31591,N_31670);
and U31753 (N_31753,N_31587,N_31678);
and U31754 (N_31754,N_31721,N_31582);
xor U31755 (N_31755,N_31563,N_31652);
and U31756 (N_31756,N_31512,N_31541);
nand U31757 (N_31757,N_31644,N_31558);
or U31758 (N_31758,N_31654,N_31688);
or U31759 (N_31759,N_31610,N_31656);
and U31760 (N_31760,N_31514,N_31573);
or U31761 (N_31761,N_31566,N_31694);
nor U31762 (N_31762,N_31621,N_31584);
xor U31763 (N_31763,N_31513,N_31509);
or U31764 (N_31764,N_31506,N_31537);
and U31765 (N_31765,N_31615,N_31575);
and U31766 (N_31766,N_31552,N_31618);
nand U31767 (N_31767,N_31551,N_31627);
nor U31768 (N_31768,N_31714,N_31613);
nand U31769 (N_31769,N_31745,N_31539);
and U31770 (N_31770,N_31735,N_31704);
nand U31771 (N_31771,N_31668,N_31616);
xnor U31772 (N_31772,N_31528,N_31665);
xnor U31773 (N_31773,N_31550,N_31592);
and U31774 (N_31774,N_31548,N_31699);
nor U31775 (N_31775,N_31549,N_31589);
or U31776 (N_31776,N_31614,N_31635);
or U31777 (N_31777,N_31527,N_31701);
or U31778 (N_31778,N_31504,N_31674);
nand U31779 (N_31779,N_31706,N_31502);
nor U31780 (N_31780,N_31728,N_31588);
and U31781 (N_31781,N_31742,N_31727);
or U31782 (N_31782,N_31565,N_31529);
and U31783 (N_31783,N_31542,N_31581);
nand U31784 (N_31784,N_31687,N_31544);
or U31785 (N_31785,N_31645,N_31505);
nor U31786 (N_31786,N_31695,N_31692);
xnor U31787 (N_31787,N_31746,N_31737);
nor U31788 (N_31788,N_31586,N_31561);
or U31789 (N_31789,N_31572,N_31696);
nor U31790 (N_31790,N_31601,N_31686);
xnor U31791 (N_31791,N_31647,N_31590);
or U31792 (N_31792,N_31700,N_31612);
nor U31793 (N_31793,N_31648,N_31522);
and U31794 (N_31794,N_31500,N_31626);
xor U31795 (N_31795,N_31739,N_31707);
and U31796 (N_31796,N_31653,N_31507);
nand U31797 (N_31797,N_31603,N_31719);
and U31798 (N_31798,N_31718,N_31609);
nand U31799 (N_31799,N_31503,N_31651);
or U31800 (N_31800,N_31526,N_31743);
xor U31801 (N_31801,N_31725,N_31625);
xnor U31802 (N_31802,N_31667,N_31661);
and U31803 (N_31803,N_31734,N_31593);
or U31804 (N_31804,N_31532,N_31630);
and U31805 (N_31805,N_31567,N_31628);
nor U31806 (N_31806,N_31594,N_31732);
or U31807 (N_31807,N_31681,N_31657);
nand U31808 (N_31808,N_31679,N_31634);
or U31809 (N_31809,N_31556,N_31623);
nor U31810 (N_31810,N_31711,N_31713);
xor U31811 (N_31811,N_31517,N_31741);
or U31812 (N_31812,N_31545,N_31726);
nand U31813 (N_31813,N_31622,N_31632);
or U31814 (N_31814,N_31747,N_31724);
or U31815 (N_31815,N_31697,N_31641);
nand U31816 (N_31816,N_31619,N_31749);
and U31817 (N_31817,N_31599,N_31702);
and U31818 (N_31818,N_31511,N_31585);
or U31819 (N_31819,N_31631,N_31658);
nand U31820 (N_31820,N_31521,N_31597);
xnor U31821 (N_31821,N_31698,N_31543);
nand U31822 (N_31822,N_31524,N_31534);
xor U31823 (N_31823,N_31620,N_31717);
nor U31824 (N_31824,N_31571,N_31662);
nor U31825 (N_31825,N_31629,N_31643);
and U31826 (N_31826,N_31716,N_31682);
nand U31827 (N_31827,N_31579,N_31501);
and U31828 (N_31828,N_31650,N_31546);
nor U31829 (N_31829,N_31595,N_31538);
and U31830 (N_31830,N_31608,N_31530);
nor U31831 (N_31831,N_31605,N_31562);
nor U31832 (N_31832,N_31740,N_31576);
nor U31833 (N_31833,N_31515,N_31663);
xor U31834 (N_31834,N_31708,N_31518);
nor U31835 (N_31835,N_31535,N_31671);
and U31836 (N_31836,N_31690,N_31570);
nor U31837 (N_31837,N_31633,N_31577);
nand U31838 (N_31838,N_31683,N_31685);
or U31839 (N_31839,N_31606,N_31720);
nor U31840 (N_31840,N_31519,N_31723);
or U31841 (N_31841,N_31540,N_31693);
or U31842 (N_31842,N_31646,N_31624);
nor U31843 (N_31843,N_31596,N_31604);
nand U31844 (N_31844,N_31744,N_31637);
nand U31845 (N_31845,N_31611,N_31730);
nor U31846 (N_31846,N_31709,N_31639);
nand U31847 (N_31847,N_31520,N_31553);
and U31848 (N_31848,N_31600,N_31676);
xor U31849 (N_31849,N_31684,N_31508);
or U31850 (N_31850,N_31703,N_31525);
or U31851 (N_31851,N_31666,N_31705);
nand U31852 (N_31852,N_31554,N_31536);
nor U31853 (N_31853,N_31640,N_31729);
nand U31854 (N_31854,N_31580,N_31715);
or U31855 (N_31855,N_31677,N_31675);
or U31856 (N_31856,N_31607,N_31638);
and U31857 (N_31857,N_31673,N_31583);
nand U31858 (N_31858,N_31557,N_31533);
or U31859 (N_31859,N_31531,N_31691);
nor U31860 (N_31860,N_31602,N_31710);
nand U31861 (N_31861,N_31564,N_31560);
nor U31862 (N_31862,N_31642,N_31574);
xor U31863 (N_31863,N_31649,N_31731);
or U31864 (N_31864,N_31568,N_31617);
nand U31865 (N_31865,N_31722,N_31669);
xor U31866 (N_31866,N_31555,N_31712);
xnor U31867 (N_31867,N_31510,N_31689);
nor U31868 (N_31868,N_31660,N_31733);
or U31869 (N_31869,N_31672,N_31559);
or U31870 (N_31870,N_31680,N_31738);
and U31871 (N_31871,N_31598,N_31659);
and U31872 (N_31872,N_31523,N_31636);
xor U31873 (N_31873,N_31664,N_31578);
nor U31874 (N_31874,N_31655,N_31547);
nand U31875 (N_31875,N_31529,N_31590);
nor U31876 (N_31876,N_31638,N_31690);
xor U31877 (N_31877,N_31597,N_31741);
and U31878 (N_31878,N_31542,N_31710);
nand U31879 (N_31879,N_31625,N_31663);
nor U31880 (N_31880,N_31507,N_31717);
xor U31881 (N_31881,N_31569,N_31661);
nand U31882 (N_31882,N_31675,N_31545);
nand U31883 (N_31883,N_31553,N_31732);
and U31884 (N_31884,N_31662,N_31594);
and U31885 (N_31885,N_31550,N_31606);
nand U31886 (N_31886,N_31602,N_31740);
or U31887 (N_31887,N_31680,N_31608);
nand U31888 (N_31888,N_31621,N_31656);
and U31889 (N_31889,N_31544,N_31693);
nor U31890 (N_31890,N_31628,N_31631);
and U31891 (N_31891,N_31506,N_31733);
nand U31892 (N_31892,N_31702,N_31556);
xor U31893 (N_31893,N_31742,N_31575);
nand U31894 (N_31894,N_31531,N_31663);
and U31895 (N_31895,N_31544,N_31654);
nand U31896 (N_31896,N_31655,N_31624);
and U31897 (N_31897,N_31651,N_31592);
xnor U31898 (N_31898,N_31693,N_31531);
nand U31899 (N_31899,N_31631,N_31510);
and U31900 (N_31900,N_31615,N_31608);
nor U31901 (N_31901,N_31719,N_31673);
xor U31902 (N_31902,N_31524,N_31636);
or U31903 (N_31903,N_31661,N_31508);
or U31904 (N_31904,N_31568,N_31563);
nor U31905 (N_31905,N_31665,N_31738);
xnor U31906 (N_31906,N_31691,N_31524);
and U31907 (N_31907,N_31714,N_31679);
or U31908 (N_31908,N_31598,N_31727);
nor U31909 (N_31909,N_31622,N_31535);
nand U31910 (N_31910,N_31503,N_31522);
xor U31911 (N_31911,N_31553,N_31522);
xnor U31912 (N_31912,N_31501,N_31626);
nor U31913 (N_31913,N_31672,N_31700);
nor U31914 (N_31914,N_31629,N_31700);
xor U31915 (N_31915,N_31594,N_31695);
xnor U31916 (N_31916,N_31736,N_31663);
or U31917 (N_31917,N_31544,N_31519);
or U31918 (N_31918,N_31505,N_31581);
xor U31919 (N_31919,N_31606,N_31601);
nor U31920 (N_31920,N_31670,N_31620);
or U31921 (N_31921,N_31668,N_31701);
xnor U31922 (N_31922,N_31717,N_31730);
or U31923 (N_31923,N_31586,N_31659);
nand U31924 (N_31924,N_31592,N_31660);
xnor U31925 (N_31925,N_31507,N_31638);
nor U31926 (N_31926,N_31691,N_31603);
or U31927 (N_31927,N_31538,N_31738);
and U31928 (N_31928,N_31595,N_31542);
or U31929 (N_31929,N_31746,N_31638);
or U31930 (N_31930,N_31504,N_31664);
or U31931 (N_31931,N_31648,N_31523);
nor U31932 (N_31932,N_31582,N_31695);
nand U31933 (N_31933,N_31670,N_31692);
nor U31934 (N_31934,N_31656,N_31521);
and U31935 (N_31935,N_31517,N_31708);
nor U31936 (N_31936,N_31638,N_31686);
nor U31937 (N_31937,N_31548,N_31628);
nor U31938 (N_31938,N_31681,N_31545);
nand U31939 (N_31939,N_31607,N_31749);
nand U31940 (N_31940,N_31535,N_31506);
xor U31941 (N_31941,N_31585,N_31630);
and U31942 (N_31942,N_31696,N_31540);
or U31943 (N_31943,N_31601,N_31592);
and U31944 (N_31944,N_31564,N_31580);
nand U31945 (N_31945,N_31596,N_31657);
xnor U31946 (N_31946,N_31601,N_31530);
and U31947 (N_31947,N_31522,N_31582);
and U31948 (N_31948,N_31514,N_31550);
nand U31949 (N_31949,N_31666,N_31645);
nor U31950 (N_31950,N_31687,N_31644);
xnor U31951 (N_31951,N_31720,N_31725);
xor U31952 (N_31952,N_31719,N_31623);
xor U31953 (N_31953,N_31722,N_31622);
nor U31954 (N_31954,N_31554,N_31730);
nor U31955 (N_31955,N_31555,N_31502);
nor U31956 (N_31956,N_31731,N_31734);
nand U31957 (N_31957,N_31708,N_31639);
or U31958 (N_31958,N_31564,N_31745);
and U31959 (N_31959,N_31575,N_31573);
nor U31960 (N_31960,N_31677,N_31571);
xnor U31961 (N_31961,N_31599,N_31616);
and U31962 (N_31962,N_31550,N_31716);
xnor U31963 (N_31963,N_31716,N_31551);
xnor U31964 (N_31964,N_31748,N_31581);
or U31965 (N_31965,N_31740,N_31606);
or U31966 (N_31966,N_31527,N_31637);
xnor U31967 (N_31967,N_31565,N_31523);
nor U31968 (N_31968,N_31567,N_31633);
or U31969 (N_31969,N_31550,N_31553);
and U31970 (N_31970,N_31690,N_31696);
or U31971 (N_31971,N_31500,N_31635);
and U31972 (N_31972,N_31600,N_31572);
or U31973 (N_31973,N_31654,N_31709);
and U31974 (N_31974,N_31656,N_31590);
nand U31975 (N_31975,N_31697,N_31594);
nor U31976 (N_31976,N_31688,N_31588);
xor U31977 (N_31977,N_31612,N_31640);
or U31978 (N_31978,N_31598,N_31685);
or U31979 (N_31979,N_31725,N_31606);
or U31980 (N_31980,N_31726,N_31639);
and U31981 (N_31981,N_31545,N_31654);
xor U31982 (N_31982,N_31641,N_31672);
or U31983 (N_31983,N_31600,N_31725);
nand U31984 (N_31984,N_31748,N_31575);
xnor U31985 (N_31985,N_31556,N_31598);
and U31986 (N_31986,N_31545,N_31524);
nand U31987 (N_31987,N_31662,N_31577);
nor U31988 (N_31988,N_31518,N_31575);
or U31989 (N_31989,N_31698,N_31736);
nand U31990 (N_31990,N_31719,N_31652);
xnor U31991 (N_31991,N_31591,N_31706);
or U31992 (N_31992,N_31555,N_31666);
or U31993 (N_31993,N_31607,N_31718);
and U31994 (N_31994,N_31726,N_31745);
xor U31995 (N_31995,N_31557,N_31717);
or U31996 (N_31996,N_31514,N_31629);
or U31997 (N_31997,N_31503,N_31637);
nand U31998 (N_31998,N_31726,N_31684);
and U31999 (N_31999,N_31565,N_31725);
xnor U32000 (N_32000,N_31872,N_31884);
xor U32001 (N_32001,N_31886,N_31802);
nand U32002 (N_32002,N_31855,N_31757);
nor U32003 (N_32003,N_31946,N_31860);
or U32004 (N_32004,N_31966,N_31774);
and U32005 (N_32005,N_31851,N_31789);
and U32006 (N_32006,N_31873,N_31815);
and U32007 (N_32007,N_31791,N_31818);
nor U32008 (N_32008,N_31786,N_31954);
nor U32009 (N_32009,N_31928,N_31793);
and U32010 (N_32010,N_31974,N_31810);
nor U32011 (N_32011,N_31994,N_31890);
or U32012 (N_32012,N_31879,N_31907);
and U32013 (N_32013,N_31779,N_31836);
nand U32014 (N_32014,N_31854,N_31978);
nand U32015 (N_32015,N_31768,N_31766);
or U32016 (N_32016,N_31861,N_31877);
nand U32017 (N_32017,N_31900,N_31969);
or U32018 (N_32018,N_31807,N_31931);
xor U32019 (N_32019,N_31968,N_31770);
nand U32020 (N_32020,N_31845,N_31816);
nor U32021 (N_32021,N_31865,N_31924);
nor U32022 (N_32022,N_31891,N_31881);
nand U32023 (N_32023,N_31976,N_31763);
xor U32024 (N_32024,N_31787,N_31918);
and U32025 (N_32025,N_31961,N_31869);
xnor U32026 (N_32026,N_31795,N_31948);
nand U32027 (N_32027,N_31932,N_31822);
nand U32028 (N_32028,N_31936,N_31947);
and U32029 (N_32029,N_31964,N_31940);
xor U32030 (N_32030,N_31903,N_31844);
or U32031 (N_32031,N_31847,N_31980);
xor U32032 (N_32032,N_31797,N_31967);
nor U32033 (N_32033,N_31849,N_31832);
and U32034 (N_32034,N_31913,N_31819);
nor U32035 (N_32035,N_31899,N_31767);
nor U32036 (N_32036,N_31977,N_31916);
xnor U32037 (N_32037,N_31929,N_31755);
nor U32038 (N_32038,N_31826,N_31777);
nor U32039 (N_32039,N_31911,N_31963);
or U32040 (N_32040,N_31962,N_31781);
nand U32041 (N_32041,N_31874,N_31896);
nor U32042 (N_32042,N_31846,N_31842);
nand U32043 (N_32043,N_31857,N_31895);
nand U32044 (N_32044,N_31804,N_31956);
and U32045 (N_32045,N_31758,N_31983);
nand U32046 (N_32046,N_31971,N_31988);
or U32047 (N_32047,N_31871,N_31825);
nor U32048 (N_32048,N_31959,N_31973);
nand U32049 (N_32049,N_31848,N_31866);
and U32050 (N_32050,N_31939,N_31750);
nand U32051 (N_32051,N_31984,N_31934);
or U32052 (N_32052,N_31785,N_31904);
or U32053 (N_32053,N_31813,N_31981);
and U32054 (N_32054,N_31778,N_31835);
or U32055 (N_32055,N_31843,N_31965);
or U32056 (N_32056,N_31930,N_31852);
or U32057 (N_32057,N_31780,N_31937);
or U32058 (N_32058,N_31756,N_31831);
and U32059 (N_32059,N_31754,N_31839);
nand U32060 (N_32060,N_31878,N_31834);
nor U32061 (N_32061,N_31943,N_31970);
xor U32062 (N_32062,N_31838,N_31782);
and U32063 (N_32063,N_31910,N_31806);
or U32064 (N_32064,N_31771,N_31960);
nor U32065 (N_32065,N_31915,N_31908);
nor U32066 (N_32066,N_31985,N_31883);
and U32067 (N_32067,N_31803,N_31752);
and U32068 (N_32068,N_31761,N_31920);
or U32069 (N_32069,N_31993,N_31783);
and U32070 (N_32070,N_31811,N_31919);
nand U32071 (N_32071,N_31897,N_31769);
xor U32072 (N_32072,N_31944,N_31801);
nor U32073 (N_32073,N_31817,N_31868);
nor U32074 (N_32074,N_31906,N_31824);
or U32075 (N_32075,N_31827,N_31952);
nand U32076 (N_32076,N_31853,N_31975);
nand U32077 (N_32077,N_31773,N_31837);
and U32078 (N_32078,N_31850,N_31945);
and U32079 (N_32079,N_31859,N_31941);
xor U32080 (N_32080,N_31805,N_31829);
or U32081 (N_32081,N_31800,N_31989);
and U32082 (N_32082,N_31927,N_31885);
and U32083 (N_32083,N_31830,N_31799);
nor U32084 (N_32084,N_31856,N_31808);
and U32085 (N_32085,N_31902,N_31921);
nand U32086 (N_32086,N_31862,N_31759);
nor U32087 (N_32087,N_31958,N_31926);
or U32088 (N_32088,N_31905,N_31889);
xor U32089 (N_32089,N_31950,N_31955);
nand U32090 (N_32090,N_31898,N_31840);
nand U32091 (N_32091,N_31772,N_31991);
nor U32092 (N_32092,N_31938,N_31949);
and U32093 (N_32093,N_31760,N_31925);
and U32094 (N_32094,N_31870,N_31828);
nand U32095 (N_32095,N_31986,N_31796);
nand U32096 (N_32096,N_31979,N_31821);
nand U32097 (N_32097,N_31882,N_31792);
nor U32098 (N_32098,N_31923,N_31917);
nor U32099 (N_32099,N_31823,N_31775);
nor U32100 (N_32100,N_31909,N_31957);
xnor U32101 (N_32101,N_31982,N_31875);
xor U32102 (N_32102,N_31765,N_31809);
xnor U32103 (N_32103,N_31880,N_31751);
or U32104 (N_32104,N_31784,N_31992);
nor U32105 (N_32105,N_31753,N_31820);
nand U32106 (N_32106,N_31892,N_31841);
nor U32107 (N_32107,N_31833,N_31995);
nor U32108 (N_32108,N_31942,N_31998);
nor U32109 (N_32109,N_31933,N_31935);
nor U32110 (N_32110,N_31762,N_31790);
xnor U32111 (N_32111,N_31887,N_31999);
xnor U32112 (N_32112,N_31893,N_31814);
or U32113 (N_32113,N_31888,N_31864);
xnor U32114 (N_32114,N_31990,N_31798);
and U32115 (N_32115,N_31867,N_31953);
or U32116 (N_32116,N_31987,N_31764);
and U32117 (N_32117,N_31876,N_31858);
nor U32118 (N_32118,N_31997,N_31912);
nand U32119 (N_32119,N_31972,N_31901);
xor U32120 (N_32120,N_31914,N_31794);
and U32121 (N_32121,N_31788,N_31894);
nor U32122 (N_32122,N_31812,N_31776);
nor U32123 (N_32123,N_31996,N_31922);
nor U32124 (N_32124,N_31863,N_31951);
xnor U32125 (N_32125,N_31813,N_31886);
or U32126 (N_32126,N_31775,N_31838);
nand U32127 (N_32127,N_31820,N_31848);
and U32128 (N_32128,N_31914,N_31884);
xor U32129 (N_32129,N_31843,N_31925);
and U32130 (N_32130,N_31932,N_31910);
xor U32131 (N_32131,N_31891,N_31934);
and U32132 (N_32132,N_31856,N_31764);
or U32133 (N_32133,N_31856,N_31803);
and U32134 (N_32134,N_31765,N_31897);
or U32135 (N_32135,N_31902,N_31949);
or U32136 (N_32136,N_31830,N_31914);
or U32137 (N_32137,N_31884,N_31859);
nand U32138 (N_32138,N_31971,N_31790);
and U32139 (N_32139,N_31816,N_31787);
and U32140 (N_32140,N_31919,N_31804);
and U32141 (N_32141,N_31832,N_31866);
nand U32142 (N_32142,N_31851,N_31824);
or U32143 (N_32143,N_31860,N_31890);
nand U32144 (N_32144,N_31857,N_31852);
nand U32145 (N_32145,N_31957,N_31894);
xor U32146 (N_32146,N_31995,N_31808);
xnor U32147 (N_32147,N_31967,N_31832);
nor U32148 (N_32148,N_31968,N_31793);
nand U32149 (N_32149,N_31773,N_31841);
or U32150 (N_32150,N_31806,N_31785);
and U32151 (N_32151,N_31828,N_31853);
or U32152 (N_32152,N_31909,N_31846);
nand U32153 (N_32153,N_31963,N_31998);
xor U32154 (N_32154,N_31752,N_31816);
xor U32155 (N_32155,N_31876,N_31824);
and U32156 (N_32156,N_31858,N_31961);
xnor U32157 (N_32157,N_31916,N_31753);
nand U32158 (N_32158,N_31763,N_31954);
nand U32159 (N_32159,N_31840,N_31957);
nor U32160 (N_32160,N_31806,N_31798);
and U32161 (N_32161,N_31920,N_31972);
nor U32162 (N_32162,N_31819,N_31937);
nand U32163 (N_32163,N_31910,N_31999);
and U32164 (N_32164,N_31966,N_31996);
xnor U32165 (N_32165,N_31902,N_31755);
nor U32166 (N_32166,N_31847,N_31909);
or U32167 (N_32167,N_31955,N_31910);
nand U32168 (N_32168,N_31828,N_31919);
nor U32169 (N_32169,N_31957,N_31931);
and U32170 (N_32170,N_31888,N_31783);
nand U32171 (N_32171,N_31834,N_31981);
nor U32172 (N_32172,N_31937,N_31813);
nand U32173 (N_32173,N_31996,N_31899);
nor U32174 (N_32174,N_31751,N_31966);
and U32175 (N_32175,N_31820,N_31824);
xnor U32176 (N_32176,N_31989,N_31906);
nor U32177 (N_32177,N_31946,N_31868);
nor U32178 (N_32178,N_31942,N_31862);
and U32179 (N_32179,N_31954,N_31816);
nand U32180 (N_32180,N_31774,N_31840);
nand U32181 (N_32181,N_31910,N_31755);
and U32182 (N_32182,N_31818,N_31922);
nand U32183 (N_32183,N_31943,N_31758);
nor U32184 (N_32184,N_31906,N_31909);
and U32185 (N_32185,N_31940,N_31903);
and U32186 (N_32186,N_31916,N_31953);
and U32187 (N_32187,N_31970,N_31876);
xnor U32188 (N_32188,N_31867,N_31893);
nand U32189 (N_32189,N_31987,N_31981);
xnor U32190 (N_32190,N_31959,N_31965);
xor U32191 (N_32191,N_31767,N_31925);
nor U32192 (N_32192,N_31942,N_31902);
xnor U32193 (N_32193,N_31963,N_31944);
xnor U32194 (N_32194,N_31979,N_31773);
or U32195 (N_32195,N_31978,N_31763);
or U32196 (N_32196,N_31959,N_31896);
or U32197 (N_32197,N_31959,N_31850);
nand U32198 (N_32198,N_31751,N_31854);
nor U32199 (N_32199,N_31975,N_31915);
nor U32200 (N_32200,N_31885,N_31919);
xnor U32201 (N_32201,N_31870,N_31991);
nor U32202 (N_32202,N_31931,N_31777);
nand U32203 (N_32203,N_31752,N_31934);
nand U32204 (N_32204,N_31808,N_31974);
and U32205 (N_32205,N_31944,N_31883);
xor U32206 (N_32206,N_31816,N_31997);
nor U32207 (N_32207,N_31964,N_31898);
nand U32208 (N_32208,N_31980,N_31810);
or U32209 (N_32209,N_31853,N_31928);
xor U32210 (N_32210,N_31840,N_31899);
nand U32211 (N_32211,N_31927,N_31905);
xor U32212 (N_32212,N_31960,N_31979);
nand U32213 (N_32213,N_31939,N_31913);
or U32214 (N_32214,N_31882,N_31908);
nor U32215 (N_32215,N_31868,N_31750);
and U32216 (N_32216,N_31790,N_31954);
nand U32217 (N_32217,N_31958,N_31884);
and U32218 (N_32218,N_31901,N_31861);
nor U32219 (N_32219,N_31804,N_31911);
xor U32220 (N_32220,N_31782,N_31958);
nor U32221 (N_32221,N_31881,N_31773);
or U32222 (N_32222,N_31917,N_31824);
nor U32223 (N_32223,N_31896,N_31987);
xnor U32224 (N_32224,N_31971,N_31829);
xor U32225 (N_32225,N_31982,N_31935);
nor U32226 (N_32226,N_31903,N_31963);
xnor U32227 (N_32227,N_31848,N_31989);
nor U32228 (N_32228,N_31804,N_31854);
nand U32229 (N_32229,N_31968,N_31847);
or U32230 (N_32230,N_31885,N_31830);
or U32231 (N_32231,N_31855,N_31839);
xnor U32232 (N_32232,N_31968,N_31935);
xnor U32233 (N_32233,N_31791,N_31794);
nand U32234 (N_32234,N_31926,N_31778);
nand U32235 (N_32235,N_31841,N_31835);
and U32236 (N_32236,N_31950,N_31824);
nor U32237 (N_32237,N_31872,N_31831);
nor U32238 (N_32238,N_31982,N_31984);
nor U32239 (N_32239,N_31990,N_31899);
and U32240 (N_32240,N_31860,N_31829);
nor U32241 (N_32241,N_31867,N_31983);
and U32242 (N_32242,N_31963,N_31864);
and U32243 (N_32243,N_31774,N_31792);
nand U32244 (N_32244,N_31969,N_31857);
and U32245 (N_32245,N_31893,N_31859);
or U32246 (N_32246,N_31824,N_31763);
xor U32247 (N_32247,N_31955,N_31997);
nor U32248 (N_32248,N_31991,N_31963);
and U32249 (N_32249,N_31831,N_31944);
or U32250 (N_32250,N_32152,N_32196);
or U32251 (N_32251,N_32070,N_32123);
or U32252 (N_32252,N_32239,N_32090);
or U32253 (N_32253,N_32187,N_32171);
xnor U32254 (N_32254,N_32034,N_32100);
and U32255 (N_32255,N_32011,N_32247);
nor U32256 (N_32256,N_32053,N_32111);
xnor U32257 (N_32257,N_32003,N_32054);
xnor U32258 (N_32258,N_32118,N_32023);
and U32259 (N_32259,N_32197,N_32047);
nor U32260 (N_32260,N_32213,N_32240);
nor U32261 (N_32261,N_32243,N_32170);
and U32262 (N_32262,N_32065,N_32236);
and U32263 (N_32263,N_32201,N_32045);
xnor U32264 (N_32264,N_32177,N_32101);
xor U32265 (N_32265,N_32228,N_32126);
or U32266 (N_32266,N_32020,N_32218);
nor U32267 (N_32267,N_32216,N_32061);
nor U32268 (N_32268,N_32199,N_32175);
and U32269 (N_32269,N_32149,N_32233);
nand U32270 (N_32270,N_32106,N_32028);
or U32271 (N_32271,N_32227,N_32229);
nand U32272 (N_32272,N_32182,N_32242);
and U32273 (N_32273,N_32099,N_32159);
and U32274 (N_32274,N_32029,N_32209);
nor U32275 (N_32275,N_32220,N_32142);
xnor U32276 (N_32276,N_32075,N_32160);
nand U32277 (N_32277,N_32188,N_32109);
nor U32278 (N_32278,N_32022,N_32107);
and U32279 (N_32279,N_32163,N_32134);
xor U32280 (N_32280,N_32231,N_32012);
and U32281 (N_32281,N_32038,N_32004);
and U32282 (N_32282,N_32035,N_32194);
xnor U32283 (N_32283,N_32198,N_32108);
and U32284 (N_32284,N_32056,N_32086);
or U32285 (N_32285,N_32044,N_32122);
xnor U32286 (N_32286,N_32173,N_32165);
and U32287 (N_32287,N_32129,N_32195);
or U32288 (N_32288,N_32009,N_32151);
and U32289 (N_32289,N_32246,N_32205);
xor U32290 (N_32290,N_32076,N_32096);
and U32291 (N_32291,N_32016,N_32208);
nand U32292 (N_32292,N_32057,N_32148);
or U32293 (N_32293,N_32059,N_32221);
nand U32294 (N_32294,N_32131,N_32157);
nor U32295 (N_32295,N_32230,N_32013);
nor U32296 (N_32296,N_32002,N_32125);
nor U32297 (N_32297,N_32007,N_32060);
and U32298 (N_32298,N_32071,N_32183);
or U32299 (N_32299,N_32062,N_32133);
nor U32300 (N_32300,N_32166,N_32167);
xnor U32301 (N_32301,N_32006,N_32024);
xnor U32302 (N_32302,N_32051,N_32048);
nor U32303 (N_32303,N_32219,N_32223);
nor U32304 (N_32304,N_32036,N_32235);
nand U32305 (N_32305,N_32095,N_32128);
nand U32306 (N_32306,N_32110,N_32169);
and U32307 (N_32307,N_32077,N_32005);
nor U32308 (N_32308,N_32114,N_32244);
or U32309 (N_32309,N_32088,N_32084);
nor U32310 (N_32310,N_32092,N_32001);
nand U32311 (N_32311,N_32140,N_32185);
and U32312 (N_32312,N_32127,N_32189);
nand U32313 (N_32313,N_32224,N_32033);
xor U32314 (N_32314,N_32222,N_32050);
and U32315 (N_32315,N_32069,N_32079);
nor U32316 (N_32316,N_32237,N_32204);
or U32317 (N_32317,N_32226,N_32202);
and U32318 (N_32318,N_32078,N_32018);
xor U32319 (N_32319,N_32238,N_32105);
and U32320 (N_32320,N_32087,N_32217);
or U32321 (N_32321,N_32074,N_32066);
nand U32322 (N_32322,N_32156,N_32184);
or U32323 (N_32323,N_32207,N_32010);
xor U32324 (N_32324,N_32132,N_32147);
and U32325 (N_32325,N_32245,N_32161);
nand U32326 (N_32326,N_32141,N_32203);
or U32327 (N_32327,N_32021,N_32154);
xor U32328 (N_32328,N_32150,N_32072);
and U32329 (N_32329,N_32031,N_32039);
nand U32330 (N_32330,N_32081,N_32193);
nand U32331 (N_32331,N_32200,N_32052);
nor U32332 (N_32332,N_32211,N_32136);
nand U32333 (N_32333,N_32186,N_32063);
and U32334 (N_32334,N_32094,N_32085);
or U32335 (N_32335,N_32174,N_32168);
or U32336 (N_32336,N_32115,N_32046);
or U32337 (N_32337,N_32097,N_32093);
nor U32338 (N_32338,N_32146,N_32083);
nor U32339 (N_32339,N_32191,N_32055);
xor U32340 (N_32340,N_32089,N_32027);
and U32341 (N_32341,N_32014,N_32119);
nand U32342 (N_32342,N_32068,N_32120);
nand U32343 (N_32343,N_32135,N_32015);
xor U32344 (N_32344,N_32117,N_32190);
xnor U32345 (N_32345,N_32082,N_32113);
or U32346 (N_32346,N_32000,N_32025);
or U32347 (N_32347,N_32019,N_32249);
xnor U32348 (N_32348,N_32178,N_32241);
xor U32349 (N_32349,N_32121,N_32073);
nand U32350 (N_32350,N_32234,N_32064);
and U32351 (N_32351,N_32102,N_32037);
nand U32352 (N_32352,N_32130,N_32030);
nor U32353 (N_32353,N_32144,N_32192);
nor U32354 (N_32354,N_32098,N_32225);
and U32355 (N_32355,N_32176,N_32058);
or U32356 (N_32356,N_32206,N_32181);
or U32357 (N_32357,N_32138,N_32040);
or U32358 (N_32358,N_32026,N_32041);
and U32359 (N_32359,N_32210,N_32043);
or U32360 (N_32360,N_32032,N_32080);
or U32361 (N_32361,N_32008,N_32049);
or U32362 (N_32362,N_32232,N_32214);
and U32363 (N_32363,N_32158,N_32179);
xor U32364 (N_32364,N_32215,N_32017);
or U32365 (N_32365,N_32104,N_32124);
nand U32366 (N_32366,N_32103,N_32116);
and U32367 (N_32367,N_32091,N_32212);
nor U32368 (N_32368,N_32145,N_32164);
or U32369 (N_32369,N_32248,N_32067);
xor U32370 (N_32370,N_32139,N_32112);
and U32371 (N_32371,N_32162,N_32172);
nor U32372 (N_32372,N_32180,N_32153);
or U32373 (N_32373,N_32042,N_32143);
nand U32374 (N_32374,N_32155,N_32137);
or U32375 (N_32375,N_32019,N_32024);
or U32376 (N_32376,N_32027,N_32094);
nand U32377 (N_32377,N_32142,N_32078);
and U32378 (N_32378,N_32057,N_32203);
xnor U32379 (N_32379,N_32004,N_32093);
nand U32380 (N_32380,N_32004,N_32236);
and U32381 (N_32381,N_32099,N_32035);
or U32382 (N_32382,N_32237,N_32198);
and U32383 (N_32383,N_32224,N_32055);
nor U32384 (N_32384,N_32088,N_32201);
nor U32385 (N_32385,N_32137,N_32167);
and U32386 (N_32386,N_32083,N_32242);
nand U32387 (N_32387,N_32078,N_32162);
nand U32388 (N_32388,N_32181,N_32215);
or U32389 (N_32389,N_32110,N_32116);
and U32390 (N_32390,N_32199,N_32183);
nand U32391 (N_32391,N_32114,N_32153);
nand U32392 (N_32392,N_32008,N_32141);
nand U32393 (N_32393,N_32058,N_32059);
nand U32394 (N_32394,N_32145,N_32036);
nor U32395 (N_32395,N_32215,N_32011);
xnor U32396 (N_32396,N_32211,N_32106);
xnor U32397 (N_32397,N_32050,N_32235);
nand U32398 (N_32398,N_32109,N_32128);
and U32399 (N_32399,N_32022,N_32071);
or U32400 (N_32400,N_32019,N_32015);
and U32401 (N_32401,N_32170,N_32204);
xor U32402 (N_32402,N_32199,N_32040);
or U32403 (N_32403,N_32132,N_32009);
or U32404 (N_32404,N_32083,N_32189);
or U32405 (N_32405,N_32028,N_32141);
and U32406 (N_32406,N_32164,N_32143);
nor U32407 (N_32407,N_32080,N_32156);
xor U32408 (N_32408,N_32034,N_32098);
and U32409 (N_32409,N_32020,N_32016);
nor U32410 (N_32410,N_32147,N_32153);
and U32411 (N_32411,N_32238,N_32229);
xor U32412 (N_32412,N_32178,N_32201);
xnor U32413 (N_32413,N_32183,N_32062);
and U32414 (N_32414,N_32018,N_32058);
xnor U32415 (N_32415,N_32082,N_32222);
nand U32416 (N_32416,N_32242,N_32075);
xnor U32417 (N_32417,N_32185,N_32209);
and U32418 (N_32418,N_32216,N_32236);
xor U32419 (N_32419,N_32120,N_32218);
nand U32420 (N_32420,N_32193,N_32142);
nand U32421 (N_32421,N_32199,N_32001);
and U32422 (N_32422,N_32174,N_32073);
nand U32423 (N_32423,N_32022,N_32086);
xor U32424 (N_32424,N_32083,N_32092);
nand U32425 (N_32425,N_32130,N_32170);
and U32426 (N_32426,N_32164,N_32155);
xor U32427 (N_32427,N_32202,N_32051);
nor U32428 (N_32428,N_32241,N_32067);
and U32429 (N_32429,N_32094,N_32107);
or U32430 (N_32430,N_32187,N_32215);
nor U32431 (N_32431,N_32136,N_32015);
or U32432 (N_32432,N_32237,N_32105);
nor U32433 (N_32433,N_32247,N_32184);
or U32434 (N_32434,N_32239,N_32167);
nor U32435 (N_32435,N_32240,N_32234);
xnor U32436 (N_32436,N_32147,N_32063);
or U32437 (N_32437,N_32228,N_32171);
and U32438 (N_32438,N_32036,N_32080);
and U32439 (N_32439,N_32206,N_32003);
and U32440 (N_32440,N_32002,N_32146);
and U32441 (N_32441,N_32130,N_32023);
and U32442 (N_32442,N_32217,N_32073);
and U32443 (N_32443,N_32178,N_32031);
or U32444 (N_32444,N_32057,N_32137);
nor U32445 (N_32445,N_32132,N_32077);
nor U32446 (N_32446,N_32208,N_32144);
and U32447 (N_32447,N_32064,N_32235);
and U32448 (N_32448,N_32033,N_32019);
nor U32449 (N_32449,N_32066,N_32132);
or U32450 (N_32450,N_32093,N_32233);
and U32451 (N_32451,N_32197,N_32210);
nand U32452 (N_32452,N_32143,N_32102);
nor U32453 (N_32453,N_32223,N_32208);
or U32454 (N_32454,N_32242,N_32166);
or U32455 (N_32455,N_32180,N_32188);
nor U32456 (N_32456,N_32088,N_32143);
xnor U32457 (N_32457,N_32047,N_32182);
xnor U32458 (N_32458,N_32124,N_32005);
nor U32459 (N_32459,N_32170,N_32119);
and U32460 (N_32460,N_32069,N_32000);
xor U32461 (N_32461,N_32231,N_32219);
or U32462 (N_32462,N_32128,N_32004);
nand U32463 (N_32463,N_32072,N_32247);
xor U32464 (N_32464,N_32135,N_32103);
or U32465 (N_32465,N_32195,N_32077);
and U32466 (N_32466,N_32219,N_32008);
or U32467 (N_32467,N_32241,N_32087);
and U32468 (N_32468,N_32135,N_32221);
nor U32469 (N_32469,N_32058,N_32027);
nand U32470 (N_32470,N_32170,N_32184);
xor U32471 (N_32471,N_32181,N_32065);
xor U32472 (N_32472,N_32199,N_32082);
nor U32473 (N_32473,N_32038,N_32151);
nor U32474 (N_32474,N_32152,N_32170);
nand U32475 (N_32475,N_32155,N_32161);
nand U32476 (N_32476,N_32183,N_32113);
and U32477 (N_32477,N_32209,N_32100);
nand U32478 (N_32478,N_32239,N_32151);
nand U32479 (N_32479,N_32161,N_32232);
and U32480 (N_32480,N_32061,N_32245);
and U32481 (N_32481,N_32001,N_32162);
or U32482 (N_32482,N_32161,N_32008);
and U32483 (N_32483,N_32037,N_32201);
nand U32484 (N_32484,N_32147,N_32020);
nor U32485 (N_32485,N_32142,N_32211);
nor U32486 (N_32486,N_32222,N_32023);
nor U32487 (N_32487,N_32208,N_32068);
and U32488 (N_32488,N_32050,N_32037);
nand U32489 (N_32489,N_32130,N_32200);
and U32490 (N_32490,N_32233,N_32001);
nand U32491 (N_32491,N_32035,N_32225);
nand U32492 (N_32492,N_32246,N_32074);
or U32493 (N_32493,N_32145,N_32047);
nand U32494 (N_32494,N_32089,N_32131);
nor U32495 (N_32495,N_32203,N_32155);
or U32496 (N_32496,N_32049,N_32127);
or U32497 (N_32497,N_32029,N_32108);
and U32498 (N_32498,N_32171,N_32225);
and U32499 (N_32499,N_32228,N_32188);
xnor U32500 (N_32500,N_32288,N_32299);
nand U32501 (N_32501,N_32375,N_32310);
or U32502 (N_32502,N_32318,N_32270);
or U32503 (N_32503,N_32250,N_32448);
and U32504 (N_32504,N_32280,N_32394);
xor U32505 (N_32505,N_32285,N_32482);
xor U32506 (N_32506,N_32414,N_32301);
nand U32507 (N_32507,N_32272,N_32290);
and U32508 (N_32508,N_32460,N_32315);
or U32509 (N_32509,N_32372,N_32439);
or U32510 (N_32510,N_32387,N_32305);
nand U32511 (N_32511,N_32298,N_32327);
and U32512 (N_32512,N_32354,N_32342);
nand U32513 (N_32513,N_32287,N_32268);
nand U32514 (N_32514,N_32396,N_32263);
nor U32515 (N_32515,N_32476,N_32412);
and U32516 (N_32516,N_32421,N_32473);
or U32517 (N_32517,N_32488,N_32345);
or U32518 (N_32518,N_32450,N_32480);
and U32519 (N_32519,N_32340,N_32269);
or U32520 (N_32520,N_32359,N_32498);
or U32521 (N_32521,N_32432,N_32368);
nor U32522 (N_32522,N_32419,N_32471);
and U32523 (N_32523,N_32465,N_32462);
nor U32524 (N_32524,N_32437,N_32378);
or U32525 (N_32525,N_32281,N_32398);
nor U32526 (N_32526,N_32442,N_32477);
or U32527 (N_32527,N_32322,N_32324);
or U32528 (N_32528,N_32400,N_32466);
nor U32529 (N_32529,N_32409,N_32426);
or U32530 (N_32530,N_32313,N_32251);
nand U32531 (N_32531,N_32258,N_32303);
and U32532 (N_32532,N_32297,N_32289);
nand U32533 (N_32533,N_32389,N_32353);
nor U32534 (N_32534,N_32267,N_32443);
or U32535 (N_32535,N_32373,N_32374);
and U32536 (N_32536,N_32347,N_32323);
nor U32537 (N_32537,N_32311,N_32433);
nand U32538 (N_32538,N_32320,N_32326);
and U32539 (N_32539,N_32346,N_32475);
nor U32540 (N_32540,N_32492,N_32335);
nand U32541 (N_32541,N_32431,N_32478);
nand U32542 (N_32542,N_32390,N_32434);
nand U32543 (N_32543,N_32415,N_32422);
or U32544 (N_32544,N_32350,N_32486);
and U32545 (N_32545,N_32464,N_32380);
xnor U32546 (N_32546,N_32472,N_32276);
nor U32547 (N_32547,N_32312,N_32447);
nor U32548 (N_32548,N_32469,N_32406);
nand U32549 (N_32549,N_32252,N_32328);
xor U32550 (N_32550,N_32423,N_32444);
or U32551 (N_32551,N_32254,N_32411);
nor U32552 (N_32552,N_32352,N_32484);
and U32553 (N_32553,N_32256,N_32356);
or U32554 (N_32554,N_32336,N_32275);
nor U32555 (N_32555,N_32458,N_32489);
nand U32556 (N_32556,N_32262,N_32319);
or U32557 (N_32557,N_32457,N_32337);
nor U32558 (N_32558,N_32467,N_32377);
and U32559 (N_32559,N_32397,N_32405);
nand U32560 (N_32560,N_32391,N_32283);
and U32561 (N_32561,N_32449,N_32363);
or U32562 (N_32562,N_32470,N_32474);
and U32563 (N_32563,N_32325,N_32441);
nor U32564 (N_32564,N_32274,N_32461);
and U32565 (N_32565,N_32261,N_32392);
and U32566 (N_32566,N_32420,N_32402);
and U32567 (N_32567,N_32333,N_32381);
or U32568 (N_32568,N_32399,N_32279);
nor U32569 (N_32569,N_32459,N_32479);
nand U32570 (N_32570,N_32369,N_32408);
nor U32571 (N_32571,N_32413,N_32278);
and U32572 (N_32572,N_32349,N_32334);
and U32573 (N_32573,N_32296,N_32384);
or U32574 (N_32574,N_32355,N_32494);
xnor U32575 (N_32575,N_32253,N_32317);
or U32576 (N_32576,N_32401,N_32348);
nand U32577 (N_32577,N_32357,N_32371);
xnor U32578 (N_32578,N_32362,N_32496);
xnor U32579 (N_32579,N_32424,N_32383);
and U32580 (N_32580,N_32273,N_32367);
xnor U32581 (N_32581,N_32455,N_32435);
and U32582 (N_32582,N_32495,N_32264);
nand U32583 (N_32583,N_32440,N_32379);
nand U32584 (N_32584,N_32445,N_32497);
nand U32585 (N_32585,N_32265,N_32376);
nand U32586 (N_32586,N_32366,N_32385);
xnor U32587 (N_32587,N_32304,N_32308);
nor U32588 (N_32588,N_32292,N_32257);
xor U32589 (N_32589,N_32407,N_32314);
or U32590 (N_32590,N_32360,N_32452);
or U32591 (N_32591,N_32393,N_32271);
or U32592 (N_32592,N_32485,N_32259);
and U32593 (N_32593,N_32417,N_32425);
or U32594 (N_32594,N_32487,N_32351);
and U32595 (N_32595,N_32293,N_32302);
and U32596 (N_32596,N_32463,N_32404);
nand U32597 (N_32597,N_32429,N_32410);
nor U32598 (N_32598,N_32341,N_32343);
and U32599 (N_32599,N_32358,N_32266);
or U32600 (N_32600,N_32395,N_32329);
nand U32601 (N_32601,N_32446,N_32260);
or U32602 (N_32602,N_32416,N_32388);
nand U32603 (N_32603,N_32309,N_32306);
and U32604 (N_32604,N_32483,N_32330);
nor U32605 (N_32605,N_32316,N_32370);
nor U32606 (N_32606,N_32451,N_32291);
xnor U32607 (N_32607,N_32339,N_32454);
and U32608 (N_32608,N_32493,N_32300);
nor U32609 (N_32609,N_32338,N_32428);
nand U32610 (N_32610,N_32453,N_32403);
nand U32611 (N_32611,N_32436,N_32321);
nor U32612 (N_32612,N_32430,N_32331);
nor U32613 (N_32613,N_32307,N_32427);
nor U32614 (N_32614,N_32255,N_32481);
nor U32615 (N_32615,N_32277,N_32294);
nand U32616 (N_32616,N_32295,N_32344);
xor U32617 (N_32617,N_32386,N_32499);
xor U32618 (N_32618,N_32286,N_32491);
and U32619 (N_32619,N_32364,N_32284);
and U32620 (N_32620,N_32490,N_32438);
or U32621 (N_32621,N_32456,N_32468);
or U32622 (N_32622,N_32365,N_32332);
or U32623 (N_32623,N_32382,N_32418);
xnor U32624 (N_32624,N_32282,N_32361);
nand U32625 (N_32625,N_32308,N_32278);
nor U32626 (N_32626,N_32337,N_32437);
nor U32627 (N_32627,N_32486,N_32365);
or U32628 (N_32628,N_32411,N_32347);
or U32629 (N_32629,N_32251,N_32408);
xnor U32630 (N_32630,N_32440,N_32325);
or U32631 (N_32631,N_32270,N_32441);
nand U32632 (N_32632,N_32416,N_32264);
nand U32633 (N_32633,N_32435,N_32467);
nor U32634 (N_32634,N_32310,N_32358);
nand U32635 (N_32635,N_32370,N_32313);
or U32636 (N_32636,N_32293,N_32255);
xnor U32637 (N_32637,N_32366,N_32420);
or U32638 (N_32638,N_32253,N_32268);
and U32639 (N_32639,N_32430,N_32494);
or U32640 (N_32640,N_32466,N_32404);
nor U32641 (N_32641,N_32434,N_32258);
nand U32642 (N_32642,N_32427,N_32272);
nor U32643 (N_32643,N_32365,N_32443);
nor U32644 (N_32644,N_32396,N_32260);
or U32645 (N_32645,N_32479,N_32296);
and U32646 (N_32646,N_32438,N_32423);
xor U32647 (N_32647,N_32417,N_32277);
xnor U32648 (N_32648,N_32363,N_32289);
nand U32649 (N_32649,N_32473,N_32466);
and U32650 (N_32650,N_32288,N_32279);
nand U32651 (N_32651,N_32310,N_32318);
nor U32652 (N_32652,N_32496,N_32263);
or U32653 (N_32653,N_32380,N_32296);
nor U32654 (N_32654,N_32289,N_32412);
or U32655 (N_32655,N_32413,N_32425);
xnor U32656 (N_32656,N_32448,N_32310);
and U32657 (N_32657,N_32393,N_32454);
or U32658 (N_32658,N_32337,N_32297);
nor U32659 (N_32659,N_32497,N_32255);
nor U32660 (N_32660,N_32382,N_32484);
nor U32661 (N_32661,N_32300,N_32344);
xnor U32662 (N_32662,N_32465,N_32307);
nor U32663 (N_32663,N_32321,N_32302);
or U32664 (N_32664,N_32414,N_32380);
nor U32665 (N_32665,N_32270,N_32387);
and U32666 (N_32666,N_32491,N_32296);
nor U32667 (N_32667,N_32306,N_32410);
nand U32668 (N_32668,N_32251,N_32307);
nor U32669 (N_32669,N_32468,N_32440);
nand U32670 (N_32670,N_32298,N_32262);
nor U32671 (N_32671,N_32337,N_32412);
or U32672 (N_32672,N_32465,N_32375);
xor U32673 (N_32673,N_32251,N_32346);
and U32674 (N_32674,N_32455,N_32343);
or U32675 (N_32675,N_32411,N_32323);
nand U32676 (N_32676,N_32296,N_32270);
nor U32677 (N_32677,N_32491,N_32485);
or U32678 (N_32678,N_32395,N_32388);
and U32679 (N_32679,N_32476,N_32314);
xnor U32680 (N_32680,N_32415,N_32297);
or U32681 (N_32681,N_32380,N_32259);
xnor U32682 (N_32682,N_32441,N_32386);
xnor U32683 (N_32683,N_32371,N_32273);
nand U32684 (N_32684,N_32411,N_32271);
nand U32685 (N_32685,N_32302,N_32421);
nor U32686 (N_32686,N_32372,N_32271);
and U32687 (N_32687,N_32446,N_32298);
and U32688 (N_32688,N_32263,N_32460);
xnor U32689 (N_32689,N_32262,N_32455);
nor U32690 (N_32690,N_32420,N_32416);
and U32691 (N_32691,N_32497,N_32459);
xor U32692 (N_32692,N_32317,N_32498);
nand U32693 (N_32693,N_32384,N_32459);
and U32694 (N_32694,N_32305,N_32401);
nand U32695 (N_32695,N_32469,N_32276);
nor U32696 (N_32696,N_32310,N_32407);
nor U32697 (N_32697,N_32330,N_32413);
nor U32698 (N_32698,N_32422,N_32314);
nand U32699 (N_32699,N_32297,N_32433);
or U32700 (N_32700,N_32258,N_32255);
xor U32701 (N_32701,N_32380,N_32418);
or U32702 (N_32702,N_32421,N_32366);
and U32703 (N_32703,N_32427,N_32275);
nand U32704 (N_32704,N_32437,N_32389);
nand U32705 (N_32705,N_32439,N_32445);
and U32706 (N_32706,N_32342,N_32312);
or U32707 (N_32707,N_32336,N_32279);
nor U32708 (N_32708,N_32368,N_32388);
nor U32709 (N_32709,N_32348,N_32399);
or U32710 (N_32710,N_32299,N_32481);
xor U32711 (N_32711,N_32377,N_32264);
xnor U32712 (N_32712,N_32352,N_32435);
nor U32713 (N_32713,N_32323,N_32368);
xor U32714 (N_32714,N_32402,N_32251);
nand U32715 (N_32715,N_32480,N_32281);
nor U32716 (N_32716,N_32293,N_32306);
xnor U32717 (N_32717,N_32382,N_32427);
or U32718 (N_32718,N_32432,N_32471);
nor U32719 (N_32719,N_32423,N_32250);
nor U32720 (N_32720,N_32393,N_32474);
nand U32721 (N_32721,N_32383,N_32373);
nand U32722 (N_32722,N_32471,N_32307);
xnor U32723 (N_32723,N_32274,N_32433);
and U32724 (N_32724,N_32344,N_32481);
and U32725 (N_32725,N_32411,N_32438);
xor U32726 (N_32726,N_32328,N_32482);
xnor U32727 (N_32727,N_32418,N_32494);
nor U32728 (N_32728,N_32438,N_32450);
or U32729 (N_32729,N_32292,N_32288);
and U32730 (N_32730,N_32308,N_32317);
xor U32731 (N_32731,N_32332,N_32404);
or U32732 (N_32732,N_32277,N_32379);
nor U32733 (N_32733,N_32277,N_32288);
xor U32734 (N_32734,N_32489,N_32417);
and U32735 (N_32735,N_32404,N_32356);
xor U32736 (N_32736,N_32260,N_32357);
nand U32737 (N_32737,N_32467,N_32434);
nand U32738 (N_32738,N_32260,N_32386);
nand U32739 (N_32739,N_32290,N_32493);
xor U32740 (N_32740,N_32282,N_32374);
nand U32741 (N_32741,N_32397,N_32258);
and U32742 (N_32742,N_32321,N_32488);
nand U32743 (N_32743,N_32493,N_32274);
and U32744 (N_32744,N_32329,N_32357);
nor U32745 (N_32745,N_32415,N_32333);
nand U32746 (N_32746,N_32344,N_32296);
xnor U32747 (N_32747,N_32389,N_32282);
and U32748 (N_32748,N_32395,N_32332);
nor U32749 (N_32749,N_32375,N_32379);
or U32750 (N_32750,N_32518,N_32657);
and U32751 (N_32751,N_32739,N_32506);
xnor U32752 (N_32752,N_32643,N_32707);
nand U32753 (N_32753,N_32537,N_32538);
xnor U32754 (N_32754,N_32549,N_32604);
nand U32755 (N_32755,N_32599,N_32530);
or U32756 (N_32756,N_32561,N_32511);
nor U32757 (N_32757,N_32730,N_32658);
xor U32758 (N_32758,N_32503,N_32689);
and U32759 (N_32759,N_32570,N_32512);
nor U32760 (N_32760,N_32524,N_32714);
nor U32761 (N_32761,N_32558,N_32545);
nand U32762 (N_32762,N_32647,N_32559);
or U32763 (N_32763,N_32728,N_32605);
nor U32764 (N_32764,N_32639,N_32514);
xor U32765 (N_32765,N_32625,N_32653);
nor U32766 (N_32766,N_32567,N_32615);
nor U32767 (N_32767,N_32609,N_32645);
or U32768 (N_32768,N_32515,N_32541);
xnor U32769 (N_32769,N_32710,N_32579);
nand U32770 (N_32770,N_32576,N_32660);
and U32771 (N_32771,N_32581,N_32577);
nand U32772 (N_32772,N_32575,N_32742);
nand U32773 (N_32773,N_32664,N_32517);
xnor U32774 (N_32774,N_32614,N_32743);
or U32775 (N_32775,N_32641,N_32540);
and U32776 (N_32776,N_32523,N_32726);
nor U32777 (N_32777,N_32686,N_32556);
or U32778 (N_32778,N_32513,N_32594);
or U32779 (N_32779,N_32674,N_32626);
nand U32780 (N_32780,N_32613,N_32547);
and U32781 (N_32781,N_32569,N_32505);
xor U32782 (N_32782,N_32676,N_32695);
nand U32783 (N_32783,N_32555,N_32718);
and U32784 (N_32784,N_32670,N_32677);
or U32785 (N_32785,N_32691,N_32712);
nor U32786 (N_32786,N_32627,N_32732);
nand U32787 (N_32787,N_32528,N_32682);
nand U32788 (N_32788,N_32648,N_32701);
nor U32789 (N_32789,N_32694,N_32671);
and U32790 (N_32790,N_32562,N_32738);
or U32791 (N_32791,N_32659,N_32683);
and U32792 (N_32792,N_32527,N_32717);
xor U32793 (N_32793,N_32516,N_32650);
or U32794 (N_32794,N_32546,N_32551);
and U32795 (N_32795,N_32636,N_32709);
nor U32796 (N_32796,N_32640,N_32631);
and U32797 (N_32797,N_32571,N_32746);
xnor U32798 (N_32798,N_32704,N_32661);
or U32799 (N_32799,N_32603,N_32591);
xnor U32800 (N_32800,N_32584,N_32679);
and U32801 (N_32801,N_32520,N_32593);
and U32802 (N_32802,N_32667,N_32668);
nor U32803 (N_32803,N_32550,N_32544);
xnor U32804 (N_32804,N_32654,N_32587);
nand U32805 (N_32805,N_32629,N_32580);
xnor U32806 (N_32806,N_32500,N_32651);
nor U32807 (N_32807,N_32705,N_32669);
or U32808 (N_32808,N_32736,N_32568);
xnor U32809 (N_32809,N_32655,N_32735);
nor U32810 (N_32810,N_32716,N_32534);
nor U32811 (N_32811,N_32565,N_32554);
xor U32812 (N_32812,N_32632,N_32543);
nand U32813 (N_32813,N_32582,N_32630);
nand U32814 (N_32814,N_32733,N_32608);
and U32815 (N_32815,N_32521,N_32692);
nand U32816 (N_32816,N_32662,N_32620);
and U32817 (N_32817,N_32678,N_32573);
xnor U32818 (N_32818,N_32633,N_32532);
nor U32819 (N_32819,N_32720,N_32708);
and U32820 (N_32820,N_32646,N_32722);
and U32821 (N_32821,N_32607,N_32610);
nor U32822 (N_32822,N_32536,N_32697);
or U32823 (N_32823,N_32711,N_32699);
and U32824 (N_32824,N_32684,N_32602);
xnor U32825 (N_32825,N_32680,N_32749);
nand U32826 (N_32826,N_32618,N_32715);
nand U32827 (N_32827,N_32634,N_32729);
xnor U32828 (N_32828,N_32589,N_32535);
nor U32829 (N_32829,N_32504,N_32696);
and U32830 (N_32830,N_32566,N_32724);
nor U32831 (N_32831,N_32745,N_32588);
xor U32832 (N_32832,N_32578,N_32635);
and U32833 (N_32833,N_32507,N_32700);
and U32834 (N_32834,N_32687,N_32526);
nor U32835 (N_32835,N_32713,N_32508);
or U32836 (N_32836,N_32666,N_32598);
nor U32837 (N_32837,N_32590,N_32519);
xnor U32838 (N_32838,N_32552,N_32672);
nand U32839 (N_32839,N_32557,N_32531);
nor U32840 (N_32840,N_32611,N_32586);
nand U32841 (N_32841,N_32737,N_32731);
nor U32842 (N_32842,N_32595,N_32542);
nor U32843 (N_32843,N_32574,N_32606);
nor U32844 (N_32844,N_32688,N_32624);
or U32845 (N_32845,N_32601,N_32560);
or U32846 (N_32846,N_32741,N_32721);
nand U32847 (N_32847,N_32681,N_32690);
nand U32848 (N_32848,N_32525,N_32612);
and U32849 (N_32849,N_32501,N_32548);
nor U32850 (N_32850,N_32706,N_32748);
nand U32851 (N_32851,N_32665,N_32597);
nand U32852 (N_32852,N_32623,N_32649);
nand U32853 (N_32853,N_32727,N_32596);
nand U32854 (N_32854,N_32622,N_32734);
or U32855 (N_32855,N_32600,N_32572);
nand U32856 (N_32856,N_32656,N_32725);
nor U32857 (N_32857,N_32533,N_32663);
nor U32858 (N_32858,N_32522,N_32693);
xnor U32859 (N_32859,N_32644,N_32502);
xnor U32860 (N_32860,N_32621,N_32642);
or U32861 (N_32861,N_32616,N_32638);
nand U32862 (N_32862,N_32592,N_32744);
nor U32863 (N_32863,N_32509,N_32617);
nand U32864 (N_32864,N_32703,N_32553);
nand U32865 (N_32865,N_32510,N_32740);
nor U32866 (N_32866,N_32652,N_32564);
nor U32867 (N_32867,N_32637,N_32685);
and U32868 (N_32868,N_32698,N_32563);
nand U32869 (N_32869,N_32539,N_32673);
nor U32870 (N_32870,N_32747,N_32675);
and U32871 (N_32871,N_32583,N_32628);
nand U32872 (N_32872,N_32529,N_32723);
or U32873 (N_32873,N_32702,N_32719);
nor U32874 (N_32874,N_32585,N_32619);
and U32875 (N_32875,N_32594,N_32556);
xor U32876 (N_32876,N_32604,N_32541);
xnor U32877 (N_32877,N_32579,N_32541);
xnor U32878 (N_32878,N_32634,N_32690);
nor U32879 (N_32879,N_32647,N_32623);
nor U32880 (N_32880,N_32631,N_32726);
and U32881 (N_32881,N_32721,N_32641);
nor U32882 (N_32882,N_32557,N_32551);
xor U32883 (N_32883,N_32716,N_32598);
nand U32884 (N_32884,N_32677,N_32504);
and U32885 (N_32885,N_32718,N_32567);
nor U32886 (N_32886,N_32670,N_32686);
nor U32887 (N_32887,N_32675,N_32556);
nor U32888 (N_32888,N_32716,N_32518);
nor U32889 (N_32889,N_32539,N_32516);
nand U32890 (N_32890,N_32690,N_32691);
xor U32891 (N_32891,N_32695,N_32685);
or U32892 (N_32892,N_32624,N_32687);
xor U32893 (N_32893,N_32516,N_32540);
or U32894 (N_32894,N_32670,N_32681);
nand U32895 (N_32895,N_32580,N_32709);
and U32896 (N_32896,N_32703,N_32691);
nand U32897 (N_32897,N_32511,N_32687);
nand U32898 (N_32898,N_32660,N_32700);
or U32899 (N_32899,N_32550,N_32722);
and U32900 (N_32900,N_32675,N_32719);
or U32901 (N_32901,N_32541,N_32591);
xor U32902 (N_32902,N_32695,N_32675);
or U32903 (N_32903,N_32533,N_32520);
and U32904 (N_32904,N_32521,N_32705);
xor U32905 (N_32905,N_32589,N_32623);
nand U32906 (N_32906,N_32704,N_32601);
nand U32907 (N_32907,N_32685,N_32576);
and U32908 (N_32908,N_32723,N_32702);
nand U32909 (N_32909,N_32700,N_32561);
or U32910 (N_32910,N_32546,N_32734);
or U32911 (N_32911,N_32576,N_32516);
nand U32912 (N_32912,N_32665,N_32502);
or U32913 (N_32913,N_32731,N_32679);
nor U32914 (N_32914,N_32572,N_32668);
nor U32915 (N_32915,N_32576,N_32550);
nor U32916 (N_32916,N_32648,N_32570);
and U32917 (N_32917,N_32535,N_32678);
nand U32918 (N_32918,N_32628,N_32701);
nand U32919 (N_32919,N_32744,N_32666);
nand U32920 (N_32920,N_32738,N_32714);
or U32921 (N_32921,N_32542,N_32546);
or U32922 (N_32922,N_32641,N_32684);
or U32923 (N_32923,N_32626,N_32747);
nor U32924 (N_32924,N_32535,N_32598);
xnor U32925 (N_32925,N_32615,N_32547);
nand U32926 (N_32926,N_32540,N_32713);
nand U32927 (N_32927,N_32666,N_32749);
and U32928 (N_32928,N_32571,N_32658);
nand U32929 (N_32929,N_32677,N_32632);
nand U32930 (N_32930,N_32730,N_32625);
or U32931 (N_32931,N_32710,N_32581);
nand U32932 (N_32932,N_32724,N_32726);
or U32933 (N_32933,N_32628,N_32651);
nand U32934 (N_32934,N_32719,N_32743);
and U32935 (N_32935,N_32611,N_32702);
or U32936 (N_32936,N_32629,N_32624);
and U32937 (N_32937,N_32695,N_32740);
nand U32938 (N_32938,N_32605,N_32709);
nand U32939 (N_32939,N_32523,N_32745);
xor U32940 (N_32940,N_32644,N_32699);
and U32941 (N_32941,N_32624,N_32716);
and U32942 (N_32942,N_32568,N_32700);
nor U32943 (N_32943,N_32747,N_32571);
nand U32944 (N_32944,N_32742,N_32585);
nand U32945 (N_32945,N_32644,N_32689);
xnor U32946 (N_32946,N_32596,N_32544);
nor U32947 (N_32947,N_32698,N_32555);
nor U32948 (N_32948,N_32651,N_32692);
and U32949 (N_32949,N_32526,N_32553);
or U32950 (N_32950,N_32663,N_32638);
nor U32951 (N_32951,N_32501,N_32526);
or U32952 (N_32952,N_32581,N_32749);
nand U32953 (N_32953,N_32636,N_32535);
nor U32954 (N_32954,N_32664,N_32548);
or U32955 (N_32955,N_32687,N_32676);
xor U32956 (N_32956,N_32506,N_32529);
or U32957 (N_32957,N_32723,N_32524);
and U32958 (N_32958,N_32736,N_32620);
nand U32959 (N_32959,N_32599,N_32634);
xor U32960 (N_32960,N_32725,N_32558);
xnor U32961 (N_32961,N_32687,N_32677);
and U32962 (N_32962,N_32626,N_32636);
and U32963 (N_32963,N_32518,N_32558);
and U32964 (N_32964,N_32563,N_32534);
nand U32965 (N_32965,N_32507,N_32539);
xor U32966 (N_32966,N_32717,N_32519);
nand U32967 (N_32967,N_32539,N_32679);
xor U32968 (N_32968,N_32522,N_32543);
xnor U32969 (N_32969,N_32534,N_32633);
or U32970 (N_32970,N_32618,N_32684);
or U32971 (N_32971,N_32546,N_32638);
and U32972 (N_32972,N_32713,N_32562);
and U32973 (N_32973,N_32677,N_32719);
and U32974 (N_32974,N_32583,N_32504);
nor U32975 (N_32975,N_32624,N_32601);
nand U32976 (N_32976,N_32544,N_32654);
nor U32977 (N_32977,N_32618,N_32571);
nand U32978 (N_32978,N_32634,N_32548);
nand U32979 (N_32979,N_32656,N_32683);
and U32980 (N_32980,N_32531,N_32617);
nand U32981 (N_32981,N_32537,N_32743);
nor U32982 (N_32982,N_32624,N_32680);
and U32983 (N_32983,N_32716,N_32749);
nand U32984 (N_32984,N_32731,N_32586);
nand U32985 (N_32985,N_32743,N_32566);
nand U32986 (N_32986,N_32699,N_32685);
and U32987 (N_32987,N_32705,N_32656);
nand U32988 (N_32988,N_32587,N_32532);
and U32989 (N_32989,N_32735,N_32687);
or U32990 (N_32990,N_32573,N_32703);
nand U32991 (N_32991,N_32599,N_32728);
xor U32992 (N_32992,N_32644,N_32524);
nand U32993 (N_32993,N_32579,N_32530);
nor U32994 (N_32994,N_32595,N_32733);
nor U32995 (N_32995,N_32545,N_32573);
nand U32996 (N_32996,N_32727,N_32651);
xnor U32997 (N_32997,N_32568,N_32615);
xnor U32998 (N_32998,N_32508,N_32504);
and U32999 (N_32999,N_32726,N_32642);
and U33000 (N_33000,N_32956,N_32790);
or U33001 (N_33001,N_32752,N_32918);
or U33002 (N_33002,N_32810,N_32973);
and U33003 (N_33003,N_32875,N_32769);
and U33004 (N_33004,N_32835,N_32798);
xor U33005 (N_33005,N_32987,N_32914);
nor U33006 (N_33006,N_32885,N_32819);
nand U33007 (N_33007,N_32771,N_32799);
or U33008 (N_33008,N_32961,N_32755);
nor U33009 (N_33009,N_32944,N_32992);
and U33010 (N_33010,N_32809,N_32784);
xor U33011 (N_33011,N_32876,N_32990);
xnor U33012 (N_33012,N_32848,N_32903);
nor U33013 (N_33013,N_32985,N_32757);
nor U33014 (N_33014,N_32965,N_32861);
xor U33015 (N_33015,N_32772,N_32837);
and U33016 (N_33016,N_32860,N_32959);
and U33017 (N_33017,N_32920,N_32866);
xnor U33018 (N_33018,N_32847,N_32865);
nor U33019 (N_33019,N_32764,N_32917);
xor U33020 (N_33020,N_32887,N_32964);
nor U33021 (N_33021,N_32941,N_32932);
nand U33022 (N_33022,N_32983,N_32834);
nand U33023 (N_33023,N_32986,N_32766);
xor U33024 (N_33024,N_32765,N_32948);
or U33025 (N_33025,N_32921,N_32905);
or U33026 (N_33026,N_32972,N_32908);
and U33027 (N_33027,N_32853,N_32900);
nor U33028 (N_33028,N_32879,N_32770);
nor U33029 (N_33029,N_32786,N_32888);
or U33030 (N_33030,N_32803,N_32759);
nor U33031 (N_33031,N_32843,N_32906);
nor U33032 (N_33032,N_32813,N_32785);
or U33033 (N_33033,N_32831,N_32934);
nand U33034 (N_33034,N_32977,N_32807);
xnor U33035 (N_33035,N_32851,N_32890);
and U33036 (N_33036,N_32919,N_32871);
and U33037 (N_33037,N_32751,N_32780);
and U33038 (N_33038,N_32966,N_32911);
or U33039 (N_33039,N_32940,N_32946);
nor U33040 (N_33040,N_32818,N_32993);
nor U33041 (N_33041,N_32976,N_32870);
xnor U33042 (N_33042,N_32859,N_32849);
or U33043 (N_33043,N_32753,N_32894);
or U33044 (N_33044,N_32923,N_32945);
nor U33045 (N_33045,N_32823,N_32904);
xor U33046 (N_33046,N_32855,N_32762);
xor U33047 (N_33047,N_32916,N_32931);
and U33048 (N_33048,N_32816,N_32979);
xor U33049 (N_33049,N_32954,N_32867);
xor U33050 (N_33050,N_32792,N_32962);
nand U33051 (N_33051,N_32836,N_32938);
xnor U33052 (N_33052,N_32793,N_32841);
nor U33053 (N_33053,N_32833,N_32830);
xnor U33054 (N_33054,N_32984,N_32943);
or U33055 (N_33055,N_32891,N_32832);
nor U33056 (N_33056,N_32788,N_32768);
and U33057 (N_33057,N_32883,N_32936);
nand U33058 (N_33058,N_32902,N_32963);
nor U33059 (N_33059,N_32995,N_32817);
xor U33060 (N_33060,N_32774,N_32858);
and U33061 (N_33061,N_32930,N_32787);
and U33062 (N_33062,N_32822,N_32797);
or U33063 (N_33063,N_32750,N_32857);
or U33064 (N_33064,N_32981,N_32844);
or U33065 (N_33065,N_32850,N_32988);
nand U33066 (N_33066,N_32820,N_32852);
nor U33067 (N_33067,N_32805,N_32869);
nand U33068 (N_33068,N_32912,N_32808);
nor U33069 (N_33069,N_32892,N_32782);
or U33070 (N_33070,N_32991,N_32895);
xnor U33071 (N_33071,N_32969,N_32978);
xor U33072 (N_33072,N_32779,N_32804);
and U33073 (N_33073,N_32874,N_32922);
or U33074 (N_33074,N_32828,N_32846);
xnor U33075 (N_33075,N_32997,N_32928);
nand U33076 (N_33076,N_32913,N_32856);
xor U33077 (N_33077,N_32862,N_32795);
and U33078 (N_33078,N_32909,N_32781);
and U33079 (N_33079,N_32889,N_32796);
or U33080 (N_33080,N_32812,N_32801);
nand U33081 (N_33081,N_32821,N_32952);
xor U33082 (N_33082,N_32994,N_32957);
or U33083 (N_33083,N_32873,N_32975);
xor U33084 (N_33084,N_32926,N_32829);
nand U33085 (N_33085,N_32863,N_32935);
nor U33086 (N_33086,N_32947,N_32910);
and U33087 (N_33087,N_32791,N_32794);
or U33088 (N_33088,N_32838,N_32968);
nor U33089 (N_33089,N_32980,N_32842);
xnor U33090 (N_33090,N_32827,N_32896);
xor U33091 (N_33091,N_32802,N_32933);
or U33092 (N_33092,N_32880,N_32898);
nor U33093 (N_33093,N_32767,N_32881);
nor U33094 (N_33094,N_32815,N_32872);
and U33095 (N_33095,N_32942,N_32868);
and U33096 (N_33096,N_32925,N_32778);
nand U33097 (N_33097,N_32758,N_32998);
xnor U33098 (N_33098,N_32775,N_32877);
xor U33099 (N_33099,N_32949,N_32814);
and U33100 (N_33100,N_32996,N_32776);
or U33101 (N_33101,N_32806,N_32789);
and U33102 (N_33102,N_32878,N_32924);
nor U33103 (N_33103,N_32754,N_32929);
or U33104 (N_33104,N_32974,N_32886);
or U33105 (N_33105,N_32967,N_32955);
xnor U33106 (N_33106,N_32989,N_32839);
nand U33107 (N_33107,N_32761,N_32907);
nor U33108 (N_33108,N_32970,N_32777);
xor U33109 (N_33109,N_32864,N_32783);
and U33110 (N_33110,N_32826,N_32854);
nand U33111 (N_33111,N_32901,N_32760);
nand U33112 (N_33112,N_32950,N_32773);
nor U33113 (N_33113,N_32927,N_32756);
xor U33114 (N_33114,N_32845,N_32824);
and U33115 (N_33115,N_32899,N_32825);
or U33116 (N_33116,N_32884,N_32937);
xnor U33117 (N_33117,N_32811,N_32960);
and U33118 (N_33118,N_32763,N_32971);
or U33119 (N_33119,N_32915,N_32800);
nor U33120 (N_33120,N_32897,N_32840);
nor U33121 (N_33121,N_32893,N_32953);
and U33122 (N_33122,N_32882,N_32982);
nor U33123 (N_33123,N_32958,N_32999);
or U33124 (N_33124,N_32939,N_32951);
nand U33125 (N_33125,N_32869,N_32987);
nor U33126 (N_33126,N_32761,N_32894);
or U33127 (N_33127,N_32977,N_32883);
nor U33128 (N_33128,N_32913,N_32887);
nor U33129 (N_33129,N_32906,N_32862);
nand U33130 (N_33130,N_32819,N_32774);
and U33131 (N_33131,N_32792,N_32933);
nor U33132 (N_33132,N_32980,N_32968);
nand U33133 (N_33133,N_32856,N_32973);
xnor U33134 (N_33134,N_32918,N_32976);
or U33135 (N_33135,N_32888,N_32995);
and U33136 (N_33136,N_32812,N_32926);
nand U33137 (N_33137,N_32750,N_32938);
and U33138 (N_33138,N_32840,N_32775);
xnor U33139 (N_33139,N_32799,N_32939);
xnor U33140 (N_33140,N_32991,N_32939);
xor U33141 (N_33141,N_32770,N_32823);
nand U33142 (N_33142,N_32897,N_32817);
nor U33143 (N_33143,N_32957,N_32866);
or U33144 (N_33144,N_32786,N_32766);
and U33145 (N_33145,N_32960,N_32956);
xnor U33146 (N_33146,N_32910,N_32929);
xor U33147 (N_33147,N_32758,N_32924);
nand U33148 (N_33148,N_32750,N_32778);
and U33149 (N_33149,N_32753,N_32945);
or U33150 (N_33150,N_32797,N_32879);
nand U33151 (N_33151,N_32806,N_32954);
nand U33152 (N_33152,N_32792,N_32970);
and U33153 (N_33153,N_32818,N_32798);
nor U33154 (N_33154,N_32861,N_32983);
or U33155 (N_33155,N_32784,N_32957);
nor U33156 (N_33156,N_32837,N_32880);
xnor U33157 (N_33157,N_32877,N_32790);
and U33158 (N_33158,N_32983,N_32979);
or U33159 (N_33159,N_32794,N_32998);
or U33160 (N_33160,N_32841,N_32921);
or U33161 (N_33161,N_32829,N_32892);
xnor U33162 (N_33162,N_32762,N_32838);
nand U33163 (N_33163,N_32932,N_32985);
nand U33164 (N_33164,N_32930,N_32750);
xor U33165 (N_33165,N_32929,N_32773);
or U33166 (N_33166,N_32934,N_32852);
nand U33167 (N_33167,N_32967,N_32796);
xor U33168 (N_33168,N_32920,N_32860);
xnor U33169 (N_33169,N_32765,N_32768);
nor U33170 (N_33170,N_32978,N_32986);
xnor U33171 (N_33171,N_32758,N_32875);
and U33172 (N_33172,N_32760,N_32982);
nor U33173 (N_33173,N_32989,N_32937);
nor U33174 (N_33174,N_32947,N_32808);
nand U33175 (N_33175,N_32881,N_32945);
and U33176 (N_33176,N_32781,N_32988);
or U33177 (N_33177,N_32781,N_32857);
xor U33178 (N_33178,N_32963,N_32896);
or U33179 (N_33179,N_32926,N_32899);
or U33180 (N_33180,N_32768,N_32944);
nand U33181 (N_33181,N_32921,N_32874);
xnor U33182 (N_33182,N_32918,N_32764);
nor U33183 (N_33183,N_32806,N_32761);
nand U33184 (N_33184,N_32783,N_32866);
and U33185 (N_33185,N_32750,N_32797);
nand U33186 (N_33186,N_32767,N_32864);
or U33187 (N_33187,N_32825,N_32905);
xor U33188 (N_33188,N_32763,N_32905);
nand U33189 (N_33189,N_32957,N_32913);
nand U33190 (N_33190,N_32824,N_32968);
nand U33191 (N_33191,N_32836,N_32834);
and U33192 (N_33192,N_32926,N_32982);
and U33193 (N_33193,N_32974,N_32933);
nand U33194 (N_33194,N_32858,N_32903);
xor U33195 (N_33195,N_32852,N_32788);
xor U33196 (N_33196,N_32879,N_32882);
nand U33197 (N_33197,N_32925,N_32755);
nor U33198 (N_33198,N_32997,N_32824);
or U33199 (N_33199,N_32831,N_32836);
nand U33200 (N_33200,N_32830,N_32777);
xnor U33201 (N_33201,N_32865,N_32829);
nor U33202 (N_33202,N_32907,N_32775);
nor U33203 (N_33203,N_32877,N_32797);
nor U33204 (N_33204,N_32959,N_32962);
nand U33205 (N_33205,N_32978,N_32811);
xor U33206 (N_33206,N_32791,N_32998);
nor U33207 (N_33207,N_32839,N_32917);
nand U33208 (N_33208,N_32880,N_32968);
nand U33209 (N_33209,N_32853,N_32856);
xor U33210 (N_33210,N_32922,N_32783);
xnor U33211 (N_33211,N_32847,N_32758);
xor U33212 (N_33212,N_32882,N_32784);
and U33213 (N_33213,N_32755,N_32953);
xnor U33214 (N_33214,N_32956,N_32813);
xor U33215 (N_33215,N_32971,N_32892);
nand U33216 (N_33216,N_32750,N_32998);
and U33217 (N_33217,N_32851,N_32757);
nand U33218 (N_33218,N_32944,N_32972);
nor U33219 (N_33219,N_32868,N_32768);
nor U33220 (N_33220,N_32890,N_32887);
or U33221 (N_33221,N_32759,N_32931);
or U33222 (N_33222,N_32850,N_32896);
nand U33223 (N_33223,N_32836,N_32835);
xnor U33224 (N_33224,N_32902,N_32865);
nor U33225 (N_33225,N_32990,N_32863);
nand U33226 (N_33226,N_32806,N_32896);
xnor U33227 (N_33227,N_32761,N_32919);
or U33228 (N_33228,N_32807,N_32838);
and U33229 (N_33229,N_32958,N_32855);
nor U33230 (N_33230,N_32784,N_32815);
nor U33231 (N_33231,N_32778,N_32936);
xor U33232 (N_33232,N_32891,N_32750);
xor U33233 (N_33233,N_32801,N_32883);
or U33234 (N_33234,N_32839,N_32976);
xnor U33235 (N_33235,N_32874,N_32754);
nor U33236 (N_33236,N_32860,N_32984);
or U33237 (N_33237,N_32975,N_32901);
nand U33238 (N_33238,N_32904,N_32866);
or U33239 (N_33239,N_32877,N_32823);
or U33240 (N_33240,N_32906,N_32751);
and U33241 (N_33241,N_32824,N_32791);
or U33242 (N_33242,N_32864,N_32903);
nand U33243 (N_33243,N_32914,N_32859);
nand U33244 (N_33244,N_32921,N_32991);
xnor U33245 (N_33245,N_32786,N_32867);
and U33246 (N_33246,N_32755,N_32962);
nand U33247 (N_33247,N_32761,N_32778);
xor U33248 (N_33248,N_32896,N_32834);
nand U33249 (N_33249,N_32888,N_32802);
nor U33250 (N_33250,N_33063,N_33126);
nor U33251 (N_33251,N_33206,N_33168);
nor U33252 (N_33252,N_33127,N_33147);
nand U33253 (N_33253,N_33042,N_33078);
xor U33254 (N_33254,N_33227,N_33052);
nor U33255 (N_33255,N_33004,N_33069);
nand U33256 (N_33256,N_33019,N_33248);
or U33257 (N_33257,N_33010,N_33220);
nand U33258 (N_33258,N_33028,N_33232);
nand U33259 (N_33259,N_33136,N_33221);
or U33260 (N_33260,N_33102,N_33149);
or U33261 (N_33261,N_33035,N_33109);
xor U33262 (N_33262,N_33038,N_33225);
xnor U33263 (N_33263,N_33008,N_33119);
xnor U33264 (N_33264,N_33107,N_33047);
or U33265 (N_33265,N_33247,N_33021);
nand U33266 (N_33266,N_33110,N_33144);
xnor U33267 (N_33267,N_33186,N_33013);
nand U33268 (N_33268,N_33087,N_33002);
or U33269 (N_33269,N_33180,N_33000);
nor U33270 (N_33270,N_33037,N_33104);
nand U33271 (N_33271,N_33092,N_33018);
or U33272 (N_33272,N_33089,N_33123);
xnor U33273 (N_33273,N_33217,N_33094);
xnor U33274 (N_33274,N_33208,N_33080);
and U33275 (N_33275,N_33166,N_33143);
nand U33276 (N_33276,N_33154,N_33061);
nand U33277 (N_33277,N_33011,N_33121);
nand U33278 (N_33278,N_33233,N_33213);
nand U33279 (N_33279,N_33016,N_33029);
nand U33280 (N_33280,N_33053,N_33197);
or U33281 (N_33281,N_33098,N_33049);
and U33282 (N_33282,N_33193,N_33231);
nor U33283 (N_33283,N_33235,N_33006);
and U33284 (N_33284,N_33071,N_33074);
xor U33285 (N_33285,N_33161,N_33204);
or U33286 (N_33286,N_33160,N_33118);
or U33287 (N_33287,N_33129,N_33237);
xnor U33288 (N_33288,N_33088,N_33022);
xnor U33289 (N_33289,N_33108,N_33146);
and U33290 (N_33290,N_33044,N_33174);
nand U33291 (N_33291,N_33239,N_33077);
nor U33292 (N_33292,N_33076,N_33111);
or U33293 (N_33293,N_33219,N_33084);
xor U33294 (N_33294,N_33134,N_33142);
or U33295 (N_33295,N_33167,N_33106);
and U33296 (N_33296,N_33055,N_33086);
nand U33297 (N_33297,N_33113,N_33209);
and U33298 (N_33298,N_33195,N_33244);
nor U33299 (N_33299,N_33009,N_33015);
or U33300 (N_33300,N_33128,N_33056);
nor U33301 (N_33301,N_33179,N_33155);
nor U33302 (N_33302,N_33207,N_33159);
or U33303 (N_33303,N_33025,N_33068);
nand U33304 (N_33304,N_33041,N_33176);
nor U33305 (N_33305,N_33043,N_33026);
and U33306 (N_33306,N_33171,N_33040);
and U33307 (N_33307,N_33218,N_33045);
nor U33308 (N_33308,N_33082,N_33152);
nand U33309 (N_33309,N_33050,N_33188);
nand U33310 (N_33310,N_33222,N_33058);
nand U33311 (N_33311,N_33099,N_33183);
and U33312 (N_33312,N_33139,N_33132);
xor U33313 (N_33313,N_33242,N_33185);
and U33314 (N_33314,N_33115,N_33187);
or U33315 (N_33315,N_33212,N_33103);
and U33316 (N_33316,N_33205,N_33057);
nor U33317 (N_33317,N_33036,N_33177);
or U33318 (N_33318,N_33243,N_33158);
and U33319 (N_33319,N_33200,N_33059);
nor U33320 (N_33320,N_33001,N_33012);
and U33321 (N_33321,N_33031,N_33048);
xnor U33322 (N_33322,N_33075,N_33184);
nand U33323 (N_33323,N_33169,N_33032);
and U33324 (N_33324,N_33034,N_33162);
xnor U33325 (N_33325,N_33140,N_33112);
and U33326 (N_33326,N_33191,N_33051);
nor U33327 (N_33327,N_33100,N_33246);
nor U33328 (N_33328,N_33194,N_33124);
and U33329 (N_33329,N_33240,N_33066);
nand U33330 (N_33330,N_33137,N_33070);
xor U33331 (N_33331,N_33241,N_33223);
nand U33332 (N_33332,N_33173,N_33064);
and U33333 (N_33333,N_33216,N_33131);
xnor U33334 (N_33334,N_33007,N_33062);
nor U33335 (N_33335,N_33085,N_33153);
nor U33336 (N_33336,N_33083,N_33120);
xor U33337 (N_33337,N_33157,N_33067);
nand U33338 (N_33338,N_33156,N_33114);
xnor U33339 (N_33339,N_33125,N_33046);
nand U33340 (N_33340,N_33192,N_33150);
xnor U33341 (N_33341,N_33020,N_33095);
and U33342 (N_33342,N_33236,N_33033);
nand U33343 (N_33343,N_33017,N_33202);
xnor U33344 (N_33344,N_33163,N_33081);
xnor U33345 (N_33345,N_33190,N_33230);
xnor U33346 (N_33346,N_33172,N_33023);
nor U33347 (N_33347,N_33101,N_33229);
nor U33348 (N_33348,N_33234,N_33096);
or U33349 (N_33349,N_33214,N_33203);
or U33350 (N_33350,N_33079,N_33170);
nor U33351 (N_33351,N_33215,N_33226);
xor U33352 (N_33352,N_33141,N_33039);
nor U33353 (N_33353,N_33024,N_33189);
and U33354 (N_33354,N_33093,N_33003);
and U33355 (N_33355,N_33175,N_33138);
nand U33356 (N_33356,N_33164,N_33224);
or U33357 (N_33357,N_33145,N_33181);
and U33358 (N_33358,N_33060,N_33073);
xor U33359 (N_33359,N_33133,N_33249);
nand U33360 (N_33360,N_33211,N_33178);
nand U33361 (N_33361,N_33091,N_33030);
or U33362 (N_33362,N_33238,N_33148);
nand U33363 (N_33363,N_33210,N_33201);
nor U33364 (N_33364,N_33182,N_33065);
xnor U33365 (N_33365,N_33196,N_33097);
nor U33366 (N_33366,N_33198,N_33151);
xnor U33367 (N_33367,N_33122,N_33054);
and U33368 (N_33368,N_33005,N_33105);
nor U33369 (N_33369,N_33199,N_33245);
nand U33370 (N_33370,N_33116,N_33135);
or U33371 (N_33371,N_33117,N_33072);
nand U33372 (N_33372,N_33090,N_33165);
or U33373 (N_33373,N_33228,N_33130);
and U33374 (N_33374,N_33014,N_33027);
nor U33375 (N_33375,N_33136,N_33049);
and U33376 (N_33376,N_33095,N_33023);
or U33377 (N_33377,N_33248,N_33185);
xnor U33378 (N_33378,N_33132,N_33092);
nor U33379 (N_33379,N_33121,N_33229);
xnor U33380 (N_33380,N_33233,N_33149);
nand U33381 (N_33381,N_33089,N_33227);
and U33382 (N_33382,N_33249,N_33152);
nand U33383 (N_33383,N_33081,N_33036);
or U33384 (N_33384,N_33192,N_33086);
and U33385 (N_33385,N_33116,N_33176);
xor U33386 (N_33386,N_33007,N_33079);
or U33387 (N_33387,N_33129,N_33102);
and U33388 (N_33388,N_33210,N_33207);
nor U33389 (N_33389,N_33243,N_33015);
and U33390 (N_33390,N_33175,N_33198);
and U33391 (N_33391,N_33110,N_33129);
or U33392 (N_33392,N_33081,N_33001);
xnor U33393 (N_33393,N_33038,N_33051);
and U33394 (N_33394,N_33227,N_33211);
and U33395 (N_33395,N_33078,N_33228);
and U33396 (N_33396,N_33113,N_33023);
and U33397 (N_33397,N_33160,N_33197);
and U33398 (N_33398,N_33101,N_33202);
nand U33399 (N_33399,N_33098,N_33093);
nor U33400 (N_33400,N_33118,N_33088);
xor U33401 (N_33401,N_33160,N_33155);
or U33402 (N_33402,N_33125,N_33052);
nor U33403 (N_33403,N_33194,N_33240);
nor U33404 (N_33404,N_33080,N_33207);
nand U33405 (N_33405,N_33062,N_33032);
nand U33406 (N_33406,N_33045,N_33014);
nor U33407 (N_33407,N_33148,N_33056);
nor U33408 (N_33408,N_33149,N_33230);
and U33409 (N_33409,N_33038,N_33108);
or U33410 (N_33410,N_33187,N_33048);
and U33411 (N_33411,N_33220,N_33112);
nor U33412 (N_33412,N_33173,N_33144);
nor U33413 (N_33413,N_33167,N_33235);
xnor U33414 (N_33414,N_33080,N_33225);
nand U33415 (N_33415,N_33205,N_33132);
nand U33416 (N_33416,N_33041,N_33175);
nand U33417 (N_33417,N_33193,N_33077);
nor U33418 (N_33418,N_33165,N_33120);
xor U33419 (N_33419,N_33063,N_33201);
or U33420 (N_33420,N_33118,N_33180);
and U33421 (N_33421,N_33029,N_33192);
nand U33422 (N_33422,N_33112,N_33114);
nand U33423 (N_33423,N_33213,N_33112);
and U33424 (N_33424,N_33099,N_33038);
xnor U33425 (N_33425,N_33115,N_33008);
or U33426 (N_33426,N_33010,N_33078);
nand U33427 (N_33427,N_33232,N_33035);
nand U33428 (N_33428,N_33172,N_33008);
and U33429 (N_33429,N_33160,N_33081);
nor U33430 (N_33430,N_33036,N_33015);
and U33431 (N_33431,N_33021,N_33062);
xnor U33432 (N_33432,N_33196,N_33067);
and U33433 (N_33433,N_33212,N_33239);
nor U33434 (N_33434,N_33004,N_33079);
nor U33435 (N_33435,N_33026,N_33238);
xor U33436 (N_33436,N_33161,N_33228);
and U33437 (N_33437,N_33063,N_33067);
and U33438 (N_33438,N_33204,N_33206);
xor U33439 (N_33439,N_33112,N_33225);
nand U33440 (N_33440,N_33124,N_33183);
nand U33441 (N_33441,N_33040,N_33208);
and U33442 (N_33442,N_33041,N_33237);
and U33443 (N_33443,N_33157,N_33220);
or U33444 (N_33444,N_33212,N_33024);
nor U33445 (N_33445,N_33243,N_33038);
nor U33446 (N_33446,N_33101,N_33022);
nand U33447 (N_33447,N_33007,N_33169);
nand U33448 (N_33448,N_33050,N_33054);
or U33449 (N_33449,N_33002,N_33028);
nand U33450 (N_33450,N_33088,N_33161);
nor U33451 (N_33451,N_33235,N_33027);
xnor U33452 (N_33452,N_33241,N_33137);
or U33453 (N_33453,N_33071,N_33004);
xor U33454 (N_33454,N_33223,N_33048);
or U33455 (N_33455,N_33060,N_33132);
or U33456 (N_33456,N_33104,N_33164);
nor U33457 (N_33457,N_33158,N_33077);
nor U33458 (N_33458,N_33239,N_33228);
xnor U33459 (N_33459,N_33131,N_33000);
nand U33460 (N_33460,N_33239,N_33223);
nand U33461 (N_33461,N_33181,N_33063);
or U33462 (N_33462,N_33093,N_33193);
nand U33463 (N_33463,N_33243,N_33159);
xor U33464 (N_33464,N_33206,N_33105);
nand U33465 (N_33465,N_33085,N_33017);
nand U33466 (N_33466,N_33097,N_33003);
xor U33467 (N_33467,N_33042,N_33205);
nand U33468 (N_33468,N_33066,N_33181);
nand U33469 (N_33469,N_33188,N_33207);
and U33470 (N_33470,N_33117,N_33052);
and U33471 (N_33471,N_33212,N_33241);
nor U33472 (N_33472,N_33032,N_33031);
xor U33473 (N_33473,N_33219,N_33169);
xnor U33474 (N_33474,N_33046,N_33071);
nand U33475 (N_33475,N_33106,N_33200);
xnor U33476 (N_33476,N_33112,N_33128);
nor U33477 (N_33477,N_33113,N_33110);
xnor U33478 (N_33478,N_33118,N_33089);
nor U33479 (N_33479,N_33134,N_33242);
nand U33480 (N_33480,N_33009,N_33077);
and U33481 (N_33481,N_33246,N_33208);
nor U33482 (N_33482,N_33050,N_33032);
or U33483 (N_33483,N_33070,N_33240);
and U33484 (N_33484,N_33216,N_33060);
xor U33485 (N_33485,N_33013,N_33147);
nor U33486 (N_33486,N_33211,N_33079);
and U33487 (N_33487,N_33062,N_33108);
nor U33488 (N_33488,N_33033,N_33035);
or U33489 (N_33489,N_33213,N_33174);
xor U33490 (N_33490,N_33010,N_33216);
nand U33491 (N_33491,N_33123,N_33133);
nor U33492 (N_33492,N_33018,N_33217);
nor U33493 (N_33493,N_33074,N_33009);
xnor U33494 (N_33494,N_33053,N_33184);
nor U33495 (N_33495,N_33080,N_33083);
or U33496 (N_33496,N_33192,N_33016);
or U33497 (N_33497,N_33038,N_33071);
nor U33498 (N_33498,N_33032,N_33040);
and U33499 (N_33499,N_33210,N_33175);
xnor U33500 (N_33500,N_33276,N_33456);
xnor U33501 (N_33501,N_33462,N_33358);
nand U33502 (N_33502,N_33329,N_33430);
or U33503 (N_33503,N_33277,N_33493);
xnor U33504 (N_33504,N_33410,N_33280);
xnor U33505 (N_33505,N_33353,N_33408);
and U33506 (N_33506,N_33259,N_33427);
and U33507 (N_33507,N_33452,N_33285);
or U33508 (N_33508,N_33386,N_33472);
nor U33509 (N_33509,N_33346,N_33269);
xnor U33510 (N_33510,N_33378,N_33282);
and U33511 (N_33511,N_33313,N_33416);
nor U33512 (N_33512,N_33350,N_33455);
or U33513 (N_33513,N_33268,N_33398);
or U33514 (N_33514,N_33320,N_33314);
xnor U33515 (N_33515,N_33435,N_33360);
or U33516 (N_33516,N_33414,N_33404);
and U33517 (N_33517,N_33373,N_33470);
nand U33518 (N_33518,N_33279,N_33281);
nor U33519 (N_33519,N_33465,N_33389);
nand U33520 (N_33520,N_33262,N_33374);
nand U33521 (N_33521,N_33444,N_33383);
nor U33522 (N_33522,N_33365,N_33300);
nand U33523 (N_33523,N_33484,N_33490);
nor U33524 (N_33524,N_33468,N_33293);
nor U33525 (N_33525,N_33434,N_33390);
nor U33526 (N_33526,N_33460,N_33301);
nor U33527 (N_33527,N_33334,N_33442);
and U33528 (N_33528,N_33298,N_33466);
nand U33529 (N_33529,N_33479,N_33306);
xor U33530 (N_33530,N_33296,N_33337);
nor U33531 (N_33531,N_33445,N_33420);
or U33532 (N_33532,N_33255,N_33324);
nand U33533 (N_33533,N_33387,N_33368);
or U33534 (N_33534,N_33370,N_33403);
nor U33535 (N_33535,N_33292,N_33307);
nand U33536 (N_33536,N_33429,N_33270);
xor U33537 (N_33537,N_33357,N_33424);
or U33538 (N_33538,N_33375,N_33492);
xor U33539 (N_33539,N_33485,N_33401);
nand U33540 (N_33540,N_33464,N_33304);
xor U33541 (N_33541,N_33379,N_33459);
and U33542 (N_33542,N_33463,N_33339);
nand U33543 (N_33543,N_33412,N_33335);
xnor U33544 (N_33544,N_33362,N_33392);
xnor U33545 (N_33545,N_33415,N_33341);
xnor U33546 (N_33546,N_33473,N_33330);
nor U33547 (N_33547,N_33446,N_33297);
nand U33548 (N_33548,N_33467,N_33400);
nand U33549 (N_33549,N_33338,N_33257);
xnor U33550 (N_33550,N_33274,N_33331);
or U33551 (N_33551,N_33396,N_33278);
and U33552 (N_33552,N_33294,N_33482);
nor U33553 (N_33553,N_33326,N_33458);
nand U33554 (N_33554,N_33436,N_33423);
nand U33555 (N_33555,N_33433,N_33454);
and U33556 (N_33556,N_33265,N_33417);
xor U33557 (N_33557,N_33469,N_33431);
nor U33558 (N_33558,N_33305,N_33397);
or U33559 (N_33559,N_33289,N_33418);
nor U33560 (N_33560,N_33380,N_33391);
nand U33561 (N_33561,N_33325,N_33286);
nor U33562 (N_33562,N_33318,N_33352);
or U33563 (N_33563,N_33449,N_33252);
or U33564 (N_33564,N_33309,N_33495);
nor U33565 (N_33565,N_33336,N_33450);
nor U33566 (N_33566,N_33295,N_33290);
nor U33567 (N_33567,N_33475,N_33347);
nand U33568 (N_33568,N_33315,N_33369);
and U33569 (N_33569,N_33413,N_33310);
or U33570 (N_33570,N_33388,N_33421);
nor U33571 (N_33571,N_33251,N_33263);
nor U33572 (N_33572,N_33422,N_33394);
or U33573 (N_33573,N_33441,N_33471);
xnor U33574 (N_33574,N_33342,N_33481);
nand U33575 (N_33575,N_33399,N_33264);
xor U33576 (N_33576,N_33322,N_33409);
xor U33577 (N_33577,N_33443,N_33428);
xor U33578 (N_33578,N_33372,N_33411);
nor U33579 (N_33579,N_33425,N_33321);
nand U33580 (N_33580,N_33483,N_33432);
nor U33581 (N_33581,N_33451,N_33332);
and U33582 (N_33582,N_33317,N_33476);
or U33583 (N_33583,N_33377,N_33381);
or U33584 (N_33584,N_33497,N_33266);
or U33585 (N_33585,N_33393,N_33351);
nand U33586 (N_33586,N_33355,N_33498);
xor U33587 (N_33587,N_33384,N_33349);
nor U33588 (N_33588,N_33376,N_33478);
xnor U33589 (N_33589,N_33488,N_33486);
and U33590 (N_33590,N_33480,N_33323);
xnor U33591 (N_33591,N_33367,N_33440);
xnor U33592 (N_33592,N_33402,N_33288);
nand U33593 (N_33593,N_33494,N_33267);
or U33594 (N_33594,N_33489,N_33302);
nor U33595 (N_33595,N_33273,N_33345);
nor U33596 (N_33596,N_33354,N_33287);
or U33597 (N_33597,N_33438,N_33453);
and U33598 (N_33598,N_33256,N_33344);
or U33599 (N_33599,N_33271,N_33366);
or U33600 (N_33600,N_33406,N_33340);
nand U33601 (N_33601,N_33250,N_33343);
and U33602 (N_33602,N_33487,N_33364);
or U33603 (N_33603,N_33275,N_33437);
nand U33604 (N_33604,N_33272,N_33499);
xor U33605 (N_33605,N_33477,N_33308);
and U33606 (N_33606,N_33382,N_33407);
and U33607 (N_33607,N_33328,N_33311);
or U33608 (N_33608,N_33448,N_33426);
xnor U33609 (N_33609,N_33457,N_33348);
and U33610 (N_33610,N_33319,N_33356);
xor U33611 (N_33611,N_33405,N_33291);
nor U33612 (N_33612,N_33461,N_33258);
xor U33613 (N_33613,N_33283,N_33496);
nor U33614 (N_33614,N_33260,N_33419);
nor U33615 (N_33615,N_33371,N_33254);
nand U33616 (N_33616,N_33474,N_33333);
nand U33617 (N_33617,N_33395,N_33359);
nor U33618 (N_33618,N_33327,N_33312);
nor U33619 (N_33619,N_33316,N_33303);
and U33620 (N_33620,N_33363,N_33447);
and U33621 (N_33621,N_33439,N_33253);
and U33622 (N_33622,N_33284,N_33361);
or U33623 (N_33623,N_33491,N_33261);
xor U33624 (N_33624,N_33299,N_33385);
and U33625 (N_33625,N_33297,N_33426);
nor U33626 (N_33626,N_33322,N_33395);
nand U33627 (N_33627,N_33331,N_33273);
nand U33628 (N_33628,N_33326,N_33471);
nor U33629 (N_33629,N_33330,N_33468);
xor U33630 (N_33630,N_33462,N_33286);
nor U33631 (N_33631,N_33423,N_33496);
nor U33632 (N_33632,N_33490,N_33486);
nor U33633 (N_33633,N_33409,N_33358);
or U33634 (N_33634,N_33483,N_33412);
or U33635 (N_33635,N_33265,N_33346);
nor U33636 (N_33636,N_33412,N_33454);
or U33637 (N_33637,N_33279,N_33320);
nand U33638 (N_33638,N_33484,N_33389);
and U33639 (N_33639,N_33334,N_33274);
or U33640 (N_33640,N_33320,N_33484);
and U33641 (N_33641,N_33301,N_33467);
nor U33642 (N_33642,N_33364,N_33414);
or U33643 (N_33643,N_33424,N_33468);
or U33644 (N_33644,N_33482,N_33348);
and U33645 (N_33645,N_33324,N_33320);
nor U33646 (N_33646,N_33430,N_33352);
or U33647 (N_33647,N_33306,N_33430);
nor U33648 (N_33648,N_33378,N_33400);
nor U33649 (N_33649,N_33382,N_33302);
xnor U33650 (N_33650,N_33321,N_33414);
and U33651 (N_33651,N_33339,N_33337);
and U33652 (N_33652,N_33350,N_33497);
and U33653 (N_33653,N_33409,N_33331);
nor U33654 (N_33654,N_33300,N_33401);
nor U33655 (N_33655,N_33393,N_33406);
or U33656 (N_33656,N_33269,N_33343);
or U33657 (N_33657,N_33346,N_33481);
nand U33658 (N_33658,N_33275,N_33263);
or U33659 (N_33659,N_33424,N_33309);
xnor U33660 (N_33660,N_33264,N_33356);
or U33661 (N_33661,N_33385,N_33288);
nor U33662 (N_33662,N_33453,N_33301);
or U33663 (N_33663,N_33450,N_33357);
xor U33664 (N_33664,N_33374,N_33422);
and U33665 (N_33665,N_33336,N_33315);
xor U33666 (N_33666,N_33259,N_33377);
nor U33667 (N_33667,N_33356,N_33368);
or U33668 (N_33668,N_33379,N_33408);
and U33669 (N_33669,N_33380,N_33489);
and U33670 (N_33670,N_33269,N_33410);
nand U33671 (N_33671,N_33445,N_33258);
xnor U33672 (N_33672,N_33470,N_33355);
xor U33673 (N_33673,N_33391,N_33350);
or U33674 (N_33674,N_33450,N_33409);
and U33675 (N_33675,N_33288,N_33365);
or U33676 (N_33676,N_33413,N_33342);
and U33677 (N_33677,N_33466,N_33485);
and U33678 (N_33678,N_33441,N_33345);
and U33679 (N_33679,N_33348,N_33303);
nand U33680 (N_33680,N_33397,N_33353);
xnor U33681 (N_33681,N_33341,N_33303);
xor U33682 (N_33682,N_33336,N_33372);
xor U33683 (N_33683,N_33373,N_33370);
nand U33684 (N_33684,N_33312,N_33321);
nand U33685 (N_33685,N_33358,N_33333);
xnor U33686 (N_33686,N_33376,N_33267);
nand U33687 (N_33687,N_33465,N_33358);
and U33688 (N_33688,N_33448,N_33257);
or U33689 (N_33689,N_33407,N_33384);
nor U33690 (N_33690,N_33360,N_33304);
and U33691 (N_33691,N_33283,N_33268);
or U33692 (N_33692,N_33290,N_33459);
or U33693 (N_33693,N_33322,N_33424);
nor U33694 (N_33694,N_33354,N_33444);
and U33695 (N_33695,N_33479,N_33281);
nor U33696 (N_33696,N_33427,N_33460);
or U33697 (N_33697,N_33343,N_33465);
or U33698 (N_33698,N_33453,N_33355);
nand U33699 (N_33699,N_33469,N_33263);
xor U33700 (N_33700,N_33310,N_33374);
nand U33701 (N_33701,N_33382,N_33338);
nor U33702 (N_33702,N_33429,N_33494);
nand U33703 (N_33703,N_33430,N_33488);
nor U33704 (N_33704,N_33317,N_33456);
nor U33705 (N_33705,N_33346,N_33429);
or U33706 (N_33706,N_33392,N_33254);
nor U33707 (N_33707,N_33298,N_33307);
nand U33708 (N_33708,N_33397,N_33374);
xor U33709 (N_33709,N_33397,N_33432);
nand U33710 (N_33710,N_33381,N_33379);
and U33711 (N_33711,N_33442,N_33378);
nand U33712 (N_33712,N_33343,N_33394);
nor U33713 (N_33713,N_33459,N_33301);
or U33714 (N_33714,N_33328,N_33464);
or U33715 (N_33715,N_33257,N_33485);
and U33716 (N_33716,N_33299,N_33253);
and U33717 (N_33717,N_33325,N_33341);
xor U33718 (N_33718,N_33474,N_33297);
or U33719 (N_33719,N_33292,N_33431);
and U33720 (N_33720,N_33471,N_33478);
or U33721 (N_33721,N_33259,N_33324);
or U33722 (N_33722,N_33300,N_33302);
nor U33723 (N_33723,N_33307,N_33428);
or U33724 (N_33724,N_33462,N_33449);
nand U33725 (N_33725,N_33405,N_33440);
or U33726 (N_33726,N_33329,N_33424);
nor U33727 (N_33727,N_33449,N_33335);
nor U33728 (N_33728,N_33443,N_33317);
nand U33729 (N_33729,N_33314,N_33364);
and U33730 (N_33730,N_33472,N_33398);
and U33731 (N_33731,N_33312,N_33322);
and U33732 (N_33732,N_33337,N_33271);
nor U33733 (N_33733,N_33270,N_33333);
nor U33734 (N_33734,N_33415,N_33388);
or U33735 (N_33735,N_33361,N_33312);
xnor U33736 (N_33736,N_33283,N_33463);
nand U33737 (N_33737,N_33461,N_33371);
nand U33738 (N_33738,N_33307,N_33466);
or U33739 (N_33739,N_33281,N_33481);
nor U33740 (N_33740,N_33379,N_33417);
nor U33741 (N_33741,N_33280,N_33284);
or U33742 (N_33742,N_33331,N_33478);
nand U33743 (N_33743,N_33453,N_33315);
nand U33744 (N_33744,N_33465,N_33265);
nor U33745 (N_33745,N_33310,N_33458);
and U33746 (N_33746,N_33283,N_33418);
nor U33747 (N_33747,N_33477,N_33350);
nand U33748 (N_33748,N_33278,N_33296);
or U33749 (N_33749,N_33390,N_33488);
nor U33750 (N_33750,N_33505,N_33516);
nand U33751 (N_33751,N_33711,N_33695);
or U33752 (N_33752,N_33612,N_33598);
nand U33753 (N_33753,N_33506,N_33591);
nand U33754 (N_33754,N_33705,N_33699);
and U33755 (N_33755,N_33543,N_33640);
nand U33756 (N_33756,N_33568,N_33529);
or U33757 (N_33757,N_33658,N_33571);
nor U33758 (N_33758,N_33698,N_33637);
nor U33759 (N_33759,N_33703,N_33531);
or U33760 (N_33760,N_33585,N_33731);
xor U33761 (N_33761,N_33638,N_33580);
nand U33762 (N_33762,N_33670,N_33660);
nand U33763 (N_33763,N_33718,N_33737);
xnor U33764 (N_33764,N_33576,N_33667);
nand U33765 (N_33765,N_33528,N_33740);
nand U33766 (N_33766,N_33526,N_33558);
nor U33767 (N_33767,N_33641,N_33726);
xnor U33768 (N_33768,N_33566,N_33678);
nand U33769 (N_33769,N_33646,N_33693);
xnor U33770 (N_33770,N_33509,N_33501);
and U33771 (N_33771,N_33709,N_33743);
and U33772 (N_33772,N_33519,N_33672);
and U33773 (N_33773,N_33690,N_33653);
or U33774 (N_33774,N_33683,N_33630);
and U33775 (N_33775,N_33665,N_33602);
nand U33776 (N_33776,N_33560,N_33682);
nor U33777 (N_33777,N_33625,N_33574);
nand U33778 (N_33778,N_33639,N_33623);
and U33779 (N_33779,N_33621,N_33627);
nor U33780 (N_33780,N_33570,N_33680);
and U33781 (N_33781,N_33557,N_33618);
xnor U33782 (N_33782,N_33575,N_33527);
and U33783 (N_33783,N_33694,N_33596);
nor U33784 (N_33784,N_33707,N_33719);
and U33785 (N_33785,N_33628,N_33600);
xnor U33786 (N_33786,N_33684,N_33616);
or U33787 (N_33787,N_33545,N_33583);
nand U33788 (N_33788,N_33607,N_33524);
nor U33789 (N_33789,N_33689,N_33727);
or U33790 (N_33790,N_33702,N_33520);
nand U33791 (N_33791,N_33654,N_33721);
and U33792 (N_33792,N_33535,N_33569);
and U33793 (N_33793,N_33663,N_33552);
or U33794 (N_33794,N_33661,N_33581);
and U33795 (N_33795,N_33636,N_33554);
nor U33796 (N_33796,N_33746,N_33582);
or U33797 (N_33797,N_33687,N_33510);
xnor U33798 (N_33798,N_33530,N_33536);
or U33799 (N_33799,N_33652,N_33631);
or U33800 (N_33800,N_33634,N_33513);
nand U33801 (N_33801,N_33525,N_33728);
nor U33802 (N_33802,N_33723,N_33534);
xor U33803 (N_33803,N_33669,N_33700);
xnor U33804 (N_33804,N_33633,N_33714);
xnor U33805 (N_33805,N_33594,N_33502);
nand U33806 (N_33806,N_33503,N_33604);
and U33807 (N_33807,N_33565,N_33595);
or U33808 (N_33808,N_33567,N_33744);
and U33809 (N_33809,N_33648,N_33589);
nand U33810 (N_33810,N_33608,N_33725);
nor U33811 (N_33811,N_33708,N_33666);
xor U33812 (N_33812,N_33550,N_33624);
nor U33813 (N_33813,N_33538,N_33590);
and U33814 (N_33814,N_33650,N_33511);
nand U33815 (N_33815,N_33584,N_33617);
nand U33816 (N_33816,N_33720,N_33561);
nand U33817 (N_33817,N_33685,N_33573);
xor U33818 (N_33818,N_33671,N_33713);
and U33819 (N_33819,N_33729,N_33688);
or U33820 (N_33820,N_33610,N_33697);
xnor U33821 (N_33821,N_33504,N_33741);
and U33822 (N_33822,N_33717,N_33696);
xor U33823 (N_33823,N_33662,N_33605);
or U33824 (N_33824,N_33613,N_33572);
xor U33825 (N_33825,N_33715,N_33742);
xor U33826 (N_33826,N_33673,N_33619);
nor U33827 (N_33827,N_33593,N_33603);
nand U33828 (N_33828,N_33681,N_33562);
or U33829 (N_33829,N_33563,N_33588);
nor U33830 (N_33830,N_33732,N_33691);
and U33831 (N_33831,N_33547,N_33508);
and U33832 (N_33832,N_33692,N_33701);
xor U33833 (N_33833,N_33514,N_33577);
and U33834 (N_33834,N_33745,N_33674);
or U33835 (N_33835,N_33515,N_33614);
and U33836 (N_33836,N_33676,N_33645);
nand U33837 (N_33837,N_33643,N_33609);
and U33838 (N_33838,N_33539,N_33656);
and U33839 (N_33839,N_33749,N_33517);
xor U33840 (N_33840,N_33626,N_33512);
or U33841 (N_33841,N_33544,N_33710);
nor U33842 (N_33842,N_33522,N_33500);
and U33843 (N_33843,N_33601,N_33553);
or U33844 (N_33844,N_33651,N_33549);
xnor U33845 (N_33845,N_33537,N_33551);
or U33846 (N_33846,N_33541,N_33556);
and U33847 (N_33847,N_33716,N_33704);
xnor U33848 (N_33848,N_33735,N_33578);
xnor U33849 (N_33849,N_33712,N_33615);
nor U33850 (N_33850,N_33686,N_33657);
or U33851 (N_33851,N_33747,N_33722);
nand U33852 (N_33852,N_33597,N_33564);
or U33853 (N_33853,N_33655,N_33523);
and U33854 (N_33854,N_33668,N_33739);
nor U33855 (N_33855,N_33649,N_33606);
nand U33856 (N_33856,N_33706,N_33592);
and U33857 (N_33857,N_33748,N_33622);
xnor U33858 (N_33858,N_33738,N_33632);
or U33859 (N_33859,N_33677,N_33620);
xor U33860 (N_33860,N_33659,N_33579);
or U33861 (N_33861,N_33533,N_33644);
and U33862 (N_33862,N_33733,N_33540);
nand U33863 (N_33863,N_33664,N_33548);
nand U33864 (N_33864,N_33546,N_33507);
nand U33865 (N_33865,N_33559,N_33629);
nand U33866 (N_33866,N_33724,N_33555);
nor U33867 (N_33867,N_33587,N_33734);
and U33868 (N_33868,N_33642,N_33730);
nor U33869 (N_33869,N_33532,N_33635);
and U33870 (N_33870,N_33736,N_33599);
and U33871 (N_33871,N_33521,N_33542);
and U33872 (N_33872,N_33611,N_33679);
or U33873 (N_33873,N_33586,N_33647);
and U33874 (N_33874,N_33675,N_33518);
or U33875 (N_33875,N_33602,N_33538);
nor U33876 (N_33876,N_33511,N_33726);
xor U33877 (N_33877,N_33653,N_33600);
and U33878 (N_33878,N_33524,N_33643);
nor U33879 (N_33879,N_33574,N_33623);
and U33880 (N_33880,N_33655,N_33672);
xor U33881 (N_33881,N_33612,N_33729);
nand U33882 (N_33882,N_33627,N_33654);
or U33883 (N_33883,N_33520,N_33698);
or U33884 (N_33884,N_33679,N_33594);
nor U33885 (N_33885,N_33708,N_33624);
or U33886 (N_33886,N_33559,N_33529);
xnor U33887 (N_33887,N_33685,N_33589);
nand U33888 (N_33888,N_33606,N_33590);
or U33889 (N_33889,N_33677,N_33640);
nor U33890 (N_33890,N_33517,N_33628);
and U33891 (N_33891,N_33627,N_33677);
and U33892 (N_33892,N_33646,N_33647);
nor U33893 (N_33893,N_33711,N_33653);
nor U33894 (N_33894,N_33574,N_33604);
or U33895 (N_33895,N_33640,N_33658);
or U33896 (N_33896,N_33689,N_33621);
or U33897 (N_33897,N_33578,N_33539);
or U33898 (N_33898,N_33692,N_33693);
nor U33899 (N_33899,N_33678,N_33648);
nor U33900 (N_33900,N_33549,N_33539);
and U33901 (N_33901,N_33614,N_33720);
and U33902 (N_33902,N_33563,N_33624);
nor U33903 (N_33903,N_33611,N_33628);
nor U33904 (N_33904,N_33571,N_33680);
xnor U33905 (N_33905,N_33741,N_33587);
nand U33906 (N_33906,N_33591,N_33574);
or U33907 (N_33907,N_33722,N_33526);
or U33908 (N_33908,N_33528,N_33749);
xnor U33909 (N_33909,N_33550,N_33571);
and U33910 (N_33910,N_33509,N_33587);
nand U33911 (N_33911,N_33569,N_33548);
and U33912 (N_33912,N_33610,N_33629);
nand U33913 (N_33913,N_33506,N_33735);
nor U33914 (N_33914,N_33654,N_33502);
nand U33915 (N_33915,N_33512,N_33548);
nor U33916 (N_33916,N_33599,N_33524);
and U33917 (N_33917,N_33729,N_33740);
xnor U33918 (N_33918,N_33684,N_33609);
or U33919 (N_33919,N_33555,N_33606);
xnor U33920 (N_33920,N_33654,N_33541);
or U33921 (N_33921,N_33744,N_33590);
nor U33922 (N_33922,N_33707,N_33611);
and U33923 (N_33923,N_33720,N_33550);
xor U33924 (N_33924,N_33593,N_33634);
or U33925 (N_33925,N_33732,N_33552);
nand U33926 (N_33926,N_33515,N_33571);
and U33927 (N_33927,N_33715,N_33731);
or U33928 (N_33928,N_33520,N_33544);
and U33929 (N_33929,N_33744,N_33618);
or U33930 (N_33930,N_33644,N_33675);
xnor U33931 (N_33931,N_33708,N_33646);
nand U33932 (N_33932,N_33620,N_33511);
or U33933 (N_33933,N_33685,N_33594);
and U33934 (N_33934,N_33524,N_33624);
nor U33935 (N_33935,N_33502,N_33601);
nor U33936 (N_33936,N_33552,N_33647);
and U33937 (N_33937,N_33506,N_33637);
and U33938 (N_33938,N_33641,N_33514);
or U33939 (N_33939,N_33731,N_33699);
nand U33940 (N_33940,N_33641,N_33626);
xor U33941 (N_33941,N_33722,N_33585);
nor U33942 (N_33942,N_33600,N_33545);
nor U33943 (N_33943,N_33592,N_33611);
nand U33944 (N_33944,N_33598,N_33548);
or U33945 (N_33945,N_33507,N_33621);
and U33946 (N_33946,N_33636,N_33559);
nand U33947 (N_33947,N_33566,N_33741);
nand U33948 (N_33948,N_33725,N_33738);
nor U33949 (N_33949,N_33500,N_33542);
or U33950 (N_33950,N_33516,N_33536);
xor U33951 (N_33951,N_33671,N_33640);
nor U33952 (N_33952,N_33572,N_33629);
nor U33953 (N_33953,N_33738,N_33648);
xor U33954 (N_33954,N_33575,N_33668);
nand U33955 (N_33955,N_33534,N_33692);
xor U33956 (N_33956,N_33711,N_33561);
or U33957 (N_33957,N_33709,N_33697);
and U33958 (N_33958,N_33625,N_33646);
or U33959 (N_33959,N_33588,N_33598);
xor U33960 (N_33960,N_33693,N_33558);
nand U33961 (N_33961,N_33669,N_33698);
xor U33962 (N_33962,N_33660,N_33520);
or U33963 (N_33963,N_33523,N_33595);
xor U33964 (N_33964,N_33670,N_33553);
and U33965 (N_33965,N_33508,N_33577);
and U33966 (N_33966,N_33684,N_33570);
nand U33967 (N_33967,N_33580,N_33516);
or U33968 (N_33968,N_33695,N_33725);
and U33969 (N_33969,N_33680,N_33712);
xor U33970 (N_33970,N_33689,N_33582);
nor U33971 (N_33971,N_33582,N_33736);
or U33972 (N_33972,N_33627,N_33520);
nor U33973 (N_33973,N_33727,N_33683);
nor U33974 (N_33974,N_33525,N_33610);
xor U33975 (N_33975,N_33543,N_33713);
nand U33976 (N_33976,N_33553,N_33644);
nor U33977 (N_33977,N_33616,N_33728);
xnor U33978 (N_33978,N_33713,N_33608);
or U33979 (N_33979,N_33630,N_33596);
nor U33980 (N_33980,N_33526,N_33531);
xor U33981 (N_33981,N_33679,N_33559);
or U33982 (N_33982,N_33667,N_33749);
xnor U33983 (N_33983,N_33525,N_33548);
nor U33984 (N_33984,N_33606,N_33574);
nand U33985 (N_33985,N_33577,N_33611);
xnor U33986 (N_33986,N_33719,N_33657);
or U33987 (N_33987,N_33549,N_33684);
xor U33988 (N_33988,N_33719,N_33648);
or U33989 (N_33989,N_33511,N_33537);
nor U33990 (N_33990,N_33648,N_33657);
nand U33991 (N_33991,N_33684,N_33702);
nor U33992 (N_33992,N_33685,N_33742);
nand U33993 (N_33993,N_33635,N_33680);
xor U33994 (N_33994,N_33610,N_33645);
nor U33995 (N_33995,N_33605,N_33522);
xor U33996 (N_33996,N_33584,N_33600);
or U33997 (N_33997,N_33642,N_33558);
nand U33998 (N_33998,N_33617,N_33675);
or U33999 (N_33999,N_33670,N_33615);
nor U34000 (N_34000,N_33819,N_33985);
or U34001 (N_34001,N_33990,N_33908);
nand U34002 (N_34002,N_33842,N_33788);
and U34003 (N_34003,N_33952,N_33827);
or U34004 (N_34004,N_33978,N_33998);
xnor U34005 (N_34005,N_33996,N_33863);
nand U34006 (N_34006,N_33854,N_33942);
nor U34007 (N_34007,N_33866,N_33930);
nand U34008 (N_34008,N_33816,N_33888);
or U34009 (N_34009,N_33799,N_33922);
and U34010 (N_34010,N_33815,N_33931);
nor U34011 (N_34011,N_33977,N_33832);
or U34012 (N_34012,N_33783,N_33843);
and U34013 (N_34013,N_33806,N_33862);
nor U34014 (N_34014,N_33918,N_33754);
xor U34015 (N_34015,N_33982,N_33861);
nand U34016 (N_34016,N_33953,N_33856);
or U34017 (N_34017,N_33965,N_33786);
xnor U34018 (N_34018,N_33929,N_33813);
nand U34019 (N_34019,N_33988,N_33928);
nand U34020 (N_34020,N_33881,N_33831);
nand U34021 (N_34021,N_33959,N_33869);
xnor U34022 (N_34022,N_33895,N_33906);
or U34023 (N_34023,N_33807,N_33966);
nor U34024 (N_34024,N_33949,N_33987);
and U34025 (N_34025,N_33913,N_33890);
or U34026 (N_34026,N_33775,N_33904);
nand U34027 (N_34027,N_33903,N_33935);
nor U34028 (N_34028,N_33969,N_33814);
nand U34029 (N_34029,N_33844,N_33972);
nor U34030 (N_34030,N_33752,N_33980);
or U34031 (N_34031,N_33921,N_33841);
and U34032 (N_34032,N_33871,N_33757);
and U34033 (N_34033,N_33923,N_33766);
or U34034 (N_34034,N_33758,N_33967);
and U34035 (N_34035,N_33789,N_33857);
nor U34036 (N_34036,N_33771,N_33898);
nand U34037 (N_34037,N_33826,N_33925);
nor U34038 (N_34038,N_33920,N_33938);
and U34039 (N_34039,N_33941,N_33781);
or U34040 (N_34040,N_33860,N_33828);
nor U34041 (N_34041,N_33825,N_33932);
and U34042 (N_34042,N_33957,N_33896);
and U34043 (N_34043,N_33765,N_33894);
xor U34044 (N_34044,N_33847,N_33933);
xor U34045 (N_34045,N_33859,N_33776);
nor U34046 (N_34046,N_33790,N_33794);
xor U34047 (N_34047,N_33874,N_33811);
nor U34048 (N_34048,N_33915,N_33845);
nor U34049 (N_34049,N_33858,N_33808);
nand U34050 (N_34050,N_33768,N_33810);
nand U34051 (N_34051,N_33802,N_33839);
xor U34052 (N_34052,N_33779,N_33916);
xor U34053 (N_34053,N_33910,N_33917);
or U34054 (N_34054,N_33800,N_33974);
nand U34055 (N_34055,N_33855,N_33865);
or U34056 (N_34056,N_33804,N_33986);
xor U34057 (N_34057,N_33902,N_33853);
or U34058 (N_34058,N_33934,N_33885);
xnor U34059 (N_34059,N_33946,N_33911);
nand U34060 (N_34060,N_33919,N_33887);
nor U34061 (N_34061,N_33973,N_33840);
nor U34062 (N_34062,N_33963,N_33880);
nor U34063 (N_34063,N_33817,N_33835);
or U34064 (N_34064,N_33951,N_33899);
or U34065 (N_34065,N_33877,N_33867);
and U34066 (N_34066,N_33760,N_33883);
nor U34067 (N_34067,N_33753,N_33773);
and U34068 (N_34068,N_33927,N_33836);
nor U34069 (N_34069,N_33787,N_33884);
nor U34070 (N_34070,N_33780,N_33795);
nand U34071 (N_34071,N_33868,N_33995);
nor U34072 (N_34072,N_33848,N_33943);
xor U34073 (N_34073,N_33955,N_33960);
nor U34074 (N_34074,N_33846,N_33962);
and U34075 (N_34075,N_33886,N_33784);
or U34076 (N_34076,N_33999,N_33782);
nor U34077 (N_34077,N_33769,N_33979);
nand U34078 (N_34078,N_33756,N_33793);
nor U34079 (N_34079,N_33924,N_33777);
nand U34080 (N_34080,N_33778,N_33905);
or U34081 (N_34081,N_33803,N_33944);
xnor U34082 (N_34082,N_33961,N_33755);
or U34083 (N_34083,N_33770,N_33798);
nor U34084 (N_34084,N_33976,N_33812);
xor U34085 (N_34085,N_33889,N_33805);
nor U34086 (N_34086,N_33864,N_33914);
and U34087 (N_34087,N_33837,N_33975);
xor U34088 (N_34088,N_33993,N_33897);
nor U34089 (N_34089,N_33870,N_33852);
or U34090 (N_34090,N_33981,N_33833);
or U34091 (N_34091,N_33759,N_33948);
and U34092 (N_34092,N_33750,N_33909);
and U34093 (N_34093,N_33785,N_33772);
nand U34094 (N_34094,N_33774,N_33849);
nor U34095 (N_34095,N_33792,N_33876);
and U34096 (N_34096,N_33821,N_33971);
nor U34097 (N_34097,N_33926,N_33936);
nor U34098 (N_34098,N_33893,N_33997);
nor U34099 (N_34099,N_33947,N_33891);
or U34100 (N_34100,N_33940,N_33954);
nor U34101 (N_34101,N_33882,N_33791);
nor U34102 (N_34102,N_33992,N_33823);
xnor U34103 (N_34103,N_33838,N_33764);
or U34104 (N_34104,N_33989,N_33797);
nand U34105 (N_34105,N_33912,N_33875);
and U34106 (N_34106,N_33751,N_33850);
nor U34107 (N_34107,N_33984,N_33829);
nor U34108 (N_34108,N_33901,N_33822);
and U34109 (N_34109,N_33945,N_33956);
or U34110 (N_34110,N_33767,N_33879);
xor U34111 (N_34111,N_33818,N_33900);
nor U34112 (N_34112,N_33761,N_33801);
and U34113 (N_34113,N_33892,N_33950);
and U34114 (N_34114,N_33762,N_33970);
or U34115 (N_34115,N_33939,N_33983);
nor U34116 (N_34116,N_33796,N_33824);
and U34117 (N_34117,N_33873,N_33994);
xor U34118 (N_34118,N_33809,N_33872);
xnor U34119 (N_34119,N_33907,N_33878);
or U34120 (N_34120,N_33991,N_33763);
nand U34121 (N_34121,N_33834,N_33937);
nor U34122 (N_34122,N_33830,N_33820);
and U34123 (N_34123,N_33958,N_33964);
or U34124 (N_34124,N_33968,N_33851);
nor U34125 (N_34125,N_33815,N_33891);
or U34126 (N_34126,N_33823,N_33781);
xnor U34127 (N_34127,N_33812,N_33853);
xor U34128 (N_34128,N_33877,N_33963);
nand U34129 (N_34129,N_33804,N_33778);
xor U34130 (N_34130,N_33862,N_33891);
xnor U34131 (N_34131,N_33870,N_33908);
or U34132 (N_34132,N_33952,N_33820);
xor U34133 (N_34133,N_33869,N_33854);
nor U34134 (N_34134,N_33757,N_33929);
and U34135 (N_34135,N_33946,N_33886);
and U34136 (N_34136,N_33921,N_33992);
or U34137 (N_34137,N_33769,N_33951);
xnor U34138 (N_34138,N_33896,N_33826);
and U34139 (N_34139,N_33940,N_33840);
and U34140 (N_34140,N_33826,N_33988);
or U34141 (N_34141,N_33854,N_33868);
xnor U34142 (N_34142,N_33942,N_33974);
nand U34143 (N_34143,N_33939,N_33772);
xor U34144 (N_34144,N_33855,N_33804);
or U34145 (N_34145,N_33763,N_33805);
or U34146 (N_34146,N_33904,N_33945);
nand U34147 (N_34147,N_33992,N_33753);
or U34148 (N_34148,N_33972,N_33905);
nor U34149 (N_34149,N_33855,N_33901);
or U34150 (N_34150,N_33854,N_33788);
or U34151 (N_34151,N_33925,N_33995);
nand U34152 (N_34152,N_33938,N_33908);
and U34153 (N_34153,N_33797,N_33756);
nand U34154 (N_34154,N_33957,N_33915);
nand U34155 (N_34155,N_33832,N_33904);
xnor U34156 (N_34156,N_33907,N_33776);
nor U34157 (N_34157,N_33883,N_33908);
or U34158 (N_34158,N_33785,N_33813);
xnor U34159 (N_34159,N_33992,N_33938);
xor U34160 (N_34160,N_33861,N_33869);
or U34161 (N_34161,N_33991,N_33965);
nor U34162 (N_34162,N_33822,N_33872);
nor U34163 (N_34163,N_33999,N_33904);
nor U34164 (N_34164,N_33878,N_33811);
nor U34165 (N_34165,N_33802,N_33764);
nand U34166 (N_34166,N_33773,N_33814);
nand U34167 (N_34167,N_33898,N_33773);
nand U34168 (N_34168,N_33770,N_33972);
nor U34169 (N_34169,N_33811,N_33791);
nor U34170 (N_34170,N_33953,N_33988);
and U34171 (N_34171,N_33976,N_33978);
or U34172 (N_34172,N_33990,N_33781);
and U34173 (N_34173,N_33761,N_33959);
xnor U34174 (N_34174,N_33910,N_33890);
nor U34175 (N_34175,N_33800,N_33771);
or U34176 (N_34176,N_33921,N_33859);
or U34177 (N_34177,N_33919,N_33994);
nand U34178 (N_34178,N_33872,N_33860);
or U34179 (N_34179,N_33836,N_33912);
nand U34180 (N_34180,N_33972,N_33946);
nor U34181 (N_34181,N_33871,N_33920);
and U34182 (N_34182,N_33927,N_33847);
nor U34183 (N_34183,N_33984,N_33897);
xnor U34184 (N_34184,N_33890,N_33767);
nor U34185 (N_34185,N_33982,N_33810);
or U34186 (N_34186,N_33932,N_33751);
and U34187 (N_34187,N_33796,N_33998);
nor U34188 (N_34188,N_33905,N_33977);
nand U34189 (N_34189,N_33818,N_33841);
nand U34190 (N_34190,N_33974,N_33883);
or U34191 (N_34191,N_33768,N_33978);
xor U34192 (N_34192,N_33892,N_33962);
xor U34193 (N_34193,N_33830,N_33881);
nor U34194 (N_34194,N_33805,N_33932);
nor U34195 (N_34195,N_33931,N_33791);
and U34196 (N_34196,N_33936,N_33832);
and U34197 (N_34197,N_33884,N_33988);
nor U34198 (N_34198,N_33899,N_33758);
or U34199 (N_34199,N_33904,N_33872);
xnor U34200 (N_34200,N_33795,N_33931);
nor U34201 (N_34201,N_33924,N_33976);
nand U34202 (N_34202,N_33776,N_33951);
xor U34203 (N_34203,N_33839,N_33794);
nand U34204 (N_34204,N_33880,N_33884);
xnor U34205 (N_34205,N_33819,N_33932);
or U34206 (N_34206,N_33841,N_33909);
xor U34207 (N_34207,N_33883,N_33840);
nor U34208 (N_34208,N_33830,N_33852);
nand U34209 (N_34209,N_33846,N_33751);
nand U34210 (N_34210,N_33852,N_33913);
or U34211 (N_34211,N_33766,N_33791);
or U34212 (N_34212,N_33850,N_33968);
xnor U34213 (N_34213,N_33854,N_33768);
nor U34214 (N_34214,N_33968,N_33988);
nand U34215 (N_34215,N_33807,N_33903);
or U34216 (N_34216,N_33988,N_33998);
nand U34217 (N_34217,N_33848,N_33910);
or U34218 (N_34218,N_33820,N_33901);
or U34219 (N_34219,N_33932,N_33922);
and U34220 (N_34220,N_33865,N_33785);
and U34221 (N_34221,N_33841,N_33908);
and U34222 (N_34222,N_33760,N_33843);
xor U34223 (N_34223,N_33885,N_33896);
xor U34224 (N_34224,N_33815,N_33869);
and U34225 (N_34225,N_33982,N_33790);
or U34226 (N_34226,N_33847,N_33830);
nor U34227 (N_34227,N_33923,N_33868);
or U34228 (N_34228,N_33972,N_33859);
or U34229 (N_34229,N_33878,N_33877);
or U34230 (N_34230,N_33843,N_33805);
nand U34231 (N_34231,N_33809,N_33859);
xor U34232 (N_34232,N_33834,N_33981);
nand U34233 (N_34233,N_33838,N_33754);
nor U34234 (N_34234,N_33817,N_33937);
or U34235 (N_34235,N_33995,N_33794);
xor U34236 (N_34236,N_33902,N_33795);
nor U34237 (N_34237,N_33760,N_33891);
nor U34238 (N_34238,N_33929,N_33787);
and U34239 (N_34239,N_33825,N_33805);
nor U34240 (N_34240,N_33984,N_33801);
nand U34241 (N_34241,N_33786,N_33913);
and U34242 (N_34242,N_33917,N_33936);
nor U34243 (N_34243,N_33835,N_33872);
xnor U34244 (N_34244,N_33902,N_33962);
nand U34245 (N_34245,N_33944,N_33750);
xor U34246 (N_34246,N_33934,N_33780);
xnor U34247 (N_34247,N_33998,N_33807);
or U34248 (N_34248,N_33857,N_33947);
nand U34249 (N_34249,N_33907,N_33769);
xnor U34250 (N_34250,N_34178,N_34117);
xnor U34251 (N_34251,N_34130,N_34163);
and U34252 (N_34252,N_34046,N_34208);
and U34253 (N_34253,N_34247,N_34176);
or U34254 (N_34254,N_34233,N_34017);
xor U34255 (N_34255,N_34047,N_34169);
or U34256 (N_34256,N_34156,N_34166);
nor U34257 (N_34257,N_34001,N_34116);
nor U34258 (N_34258,N_34009,N_34063);
or U34259 (N_34259,N_34171,N_34081);
and U34260 (N_34260,N_34016,N_34077);
and U34261 (N_34261,N_34044,N_34232);
nand U34262 (N_34262,N_34099,N_34062);
or U34263 (N_34263,N_34150,N_34118);
or U34264 (N_34264,N_34058,N_34123);
nor U34265 (N_34265,N_34043,N_34033);
nor U34266 (N_34266,N_34141,N_34186);
nor U34267 (N_34267,N_34245,N_34144);
xor U34268 (N_34268,N_34216,N_34105);
xnor U34269 (N_34269,N_34097,N_34002);
or U34270 (N_34270,N_34050,N_34053);
xnor U34271 (N_34271,N_34126,N_34194);
nor U34272 (N_34272,N_34107,N_34101);
and U34273 (N_34273,N_34207,N_34157);
nand U34274 (N_34274,N_34195,N_34114);
xnor U34275 (N_34275,N_34168,N_34022);
or U34276 (N_34276,N_34012,N_34237);
or U34277 (N_34277,N_34206,N_34181);
and U34278 (N_34278,N_34080,N_34159);
xor U34279 (N_34279,N_34167,N_34111);
and U34280 (N_34280,N_34177,N_34246);
and U34281 (N_34281,N_34201,N_34148);
xor U34282 (N_34282,N_34010,N_34098);
and U34283 (N_34283,N_34106,N_34211);
nand U34284 (N_34284,N_34104,N_34125);
nor U34285 (N_34285,N_34205,N_34041);
and U34286 (N_34286,N_34242,N_34161);
nor U34287 (N_34287,N_34019,N_34028);
xnor U34288 (N_34288,N_34076,N_34225);
or U34289 (N_34289,N_34241,N_34122);
nand U34290 (N_34290,N_34222,N_34108);
nor U34291 (N_34291,N_34200,N_34187);
or U34292 (N_34292,N_34035,N_34224);
or U34293 (N_34293,N_34079,N_34221);
nand U34294 (N_34294,N_34090,N_34027);
or U34295 (N_34295,N_34109,N_34142);
nor U34296 (N_34296,N_34146,N_34103);
xnor U34297 (N_34297,N_34182,N_34093);
or U34298 (N_34298,N_34004,N_34049);
xnor U34299 (N_34299,N_34244,N_34005);
or U34300 (N_34300,N_34197,N_34214);
nand U34301 (N_34301,N_34191,N_34021);
nor U34302 (N_34302,N_34160,N_34149);
or U34303 (N_34303,N_34032,N_34204);
and U34304 (N_34304,N_34158,N_34086);
nor U34305 (N_34305,N_34089,N_34008);
nand U34306 (N_34306,N_34153,N_34115);
nor U34307 (N_34307,N_34219,N_34066);
nor U34308 (N_34308,N_34209,N_34154);
nand U34309 (N_34309,N_34075,N_34029);
xnor U34310 (N_34310,N_34034,N_34202);
nor U34311 (N_34311,N_34138,N_34213);
xnor U34312 (N_34312,N_34140,N_34120);
and U34313 (N_34313,N_34040,N_34127);
and U34314 (N_34314,N_34112,N_34220);
and U34315 (N_34315,N_34162,N_34070);
nor U34316 (N_34316,N_34087,N_34199);
or U34317 (N_34317,N_34180,N_34007);
and U34318 (N_34318,N_34018,N_34172);
nand U34319 (N_34319,N_34072,N_34051);
or U34320 (N_34320,N_34057,N_34184);
nand U34321 (N_34321,N_34023,N_34092);
xnor U34322 (N_34322,N_34226,N_34192);
xor U34323 (N_34323,N_34038,N_34006);
xor U34324 (N_34324,N_34152,N_34230);
and U34325 (N_34325,N_34024,N_34059);
nand U34326 (N_34326,N_34238,N_34031);
nor U34327 (N_34327,N_34030,N_34234);
or U34328 (N_34328,N_34131,N_34193);
and U34329 (N_34329,N_34048,N_34175);
or U34330 (N_34330,N_34203,N_34003);
xnor U34331 (N_34331,N_34217,N_34060);
or U34332 (N_34332,N_34143,N_34054);
nor U34333 (N_34333,N_34025,N_34134);
and U34334 (N_34334,N_34227,N_34095);
nor U34335 (N_34335,N_34198,N_34102);
nor U34336 (N_34336,N_34183,N_34243);
nor U34337 (N_34337,N_34085,N_34083);
nor U34338 (N_34338,N_34014,N_34067);
xnor U34339 (N_34339,N_34235,N_34020);
or U34340 (N_34340,N_34248,N_34124);
nand U34341 (N_34341,N_34042,N_34061);
xor U34342 (N_34342,N_34188,N_34133);
and U34343 (N_34343,N_34190,N_34147);
nor U34344 (N_34344,N_34056,N_34236);
nand U34345 (N_34345,N_34071,N_34039);
or U34346 (N_34346,N_34026,N_34229);
or U34347 (N_34347,N_34136,N_34151);
nand U34348 (N_34348,N_34055,N_34091);
and U34349 (N_34349,N_34174,N_34119);
or U34350 (N_34350,N_34084,N_34239);
xnor U34351 (N_34351,N_34170,N_34240);
nand U34352 (N_34352,N_34185,N_34082);
and U34353 (N_34353,N_34068,N_34015);
nand U34354 (N_34354,N_34189,N_34000);
or U34355 (N_34355,N_34132,N_34137);
nor U34356 (N_34356,N_34069,N_34165);
xnor U34357 (N_34357,N_34052,N_34218);
nor U34358 (N_34358,N_34212,N_34096);
xnor U34359 (N_34359,N_34228,N_34196);
or U34360 (N_34360,N_34100,N_34073);
nor U34361 (N_34361,N_34231,N_34179);
nor U34362 (N_34362,N_34128,N_34164);
and U34363 (N_34363,N_34088,N_34135);
and U34364 (N_34364,N_34065,N_34223);
or U34365 (N_34365,N_34094,N_34064);
and U34366 (N_34366,N_34074,N_34173);
xor U34367 (N_34367,N_34037,N_34249);
nor U34368 (N_34368,N_34121,N_34139);
nand U34369 (N_34369,N_34036,N_34129);
and U34370 (N_34370,N_34210,N_34113);
nor U34371 (N_34371,N_34145,N_34078);
nor U34372 (N_34372,N_34013,N_34155);
or U34373 (N_34373,N_34110,N_34011);
or U34374 (N_34374,N_34045,N_34215);
or U34375 (N_34375,N_34006,N_34229);
xor U34376 (N_34376,N_34051,N_34139);
and U34377 (N_34377,N_34171,N_34192);
or U34378 (N_34378,N_34096,N_34007);
nand U34379 (N_34379,N_34241,N_34202);
nand U34380 (N_34380,N_34127,N_34000);
and U34381 (N_34381,N_34193,N_34184);
and U34382 (N_34382,N_34104,N_34008);
or U34383 (N_34383,N_34218,N_34248);
xnor U34384 (N_34384,N_34236,N_34224);
nor U34385 (N_34385,N_34147,N_34189);
xnor U34386 (N_34386,N_34188,N_34081);
and U34387 (N_34387,N_34227,N_34023);
or U34388 (N_34388,N_34043,N_34150);
nand U34389 (N_34389,N_34170,N_34231);
and U34390 (N_34390,N_34069,N_34011);
or U34391 (N_34391,N_34164,N_34133);
nand U34392 (N_34392,N_34014,N_34195);
nor U34393 (N_34393,N_34197,N_34115);
nand U34394 (N_34394,N_34205,N_34152);
or U34395 (N_34395,N_34205,N_34168);
nor U34396 (N_34396,N_34135,N_34044);
nand U34397 (N_34397,N_34107,N_34088);
or U34398 (N_34398,N_34187,N_34127);
nand U34399 (N_34399,N_34034,N_34045);
nand U34400 (N_34400,N_34061,N_34157);
xor U34401 (N_34401,N_34196,N_34185);
nand U34402 (N_34402,N_34025,N_34149);
nand U34403 (N_34403,N_34239,N_34149);
nor U34404 (N_34404,N_34150,N_34053);
xnor U34405 (N_34405,N_34114,N_34179);
nor U34406 (N_34406,N_34138,N_34188);
nor U34407 (N_34407,N_34085,N_34102);
or U34408 (N_34408,N_34099,N_34059);
xnor U34409 (N_34409,N_34140,N_34221);
or U34410 (N_34410,N_34041,N_34084);
nand U34411 (N_34411,N_34211,N_34001);
or U34412 (N_34412,N_34180,N_34103);
or U34413 (N_34413,N_34140,N_34161);
and U34414 (N_34414,N_34220,N_34073);
nor U34415 (N_34415,N_34176,N_34089);
xnor U34416 (N_34416,N_34225,N_34106);
xnor U34417 (N_34417,N_34036,N_34194);
nor U34418 (N_34418,N_34226,N_34182);
nand U34419 (N_34419,N_34078,N_34098);
nor U34420 (N_34420,N_34109,N_34172);
or U34421 (N_34421,N_34035,N_34244);
nor U34422 (N_34422,N_34030,N_34071);
xor U34423 (N_34423,N_34178,N_34046);
nor U34424 (N_34424,N_34033,N_34244);
and U34425 (N_34425,N_34167,N_34145);
and U34426 (N_34426,N_34004,N_34243);
nor U34427 (N_34427,N_34055,N_34007);
or U34428 (N_34428,N_34111,N_34211);
nand U34429 (N_34429,N_34135,N_34190);
or U34430 (N_34430,N_34059,N_34141);
nand U34431 (N_34431,N_34015,N_34001);
or U34432 (N_34432,N_34058,N_34144);
nand U34433 (N_34433,N_34119,N_34139);
and U34434 (N_34434,N_34005,N_34029);
xor U34435 (N_34435,N_34080,N_34013);
xor U34436 (N_34436,N_34034,N_34057);
and U34437 (N_34437,N_34123,N_34067);
nor U34438 (N_34438,N_34138,N_34077);
nand U34439 (N_34439,N_34063,N_34228);
nand U34440 (N_34440,N_34026,N_34007);
nand U34441 (N_34441,N_34027,N_34053);
and U34442 (N_34442,N_34219,N_34083);
nor U34443 (N_34443,N_34246,N_34114);
nor U34444 (N_34444,N_34191,N_34178);
nand U34445 (N_34445,N_34098,N_34181);
and U34446 (N_34446,N_34068,N_34145);
nand U34447 (N_34447,N_34230,N_34079);
and U34448 (N_34448,N_34096,N_34150);
nor U34449 (N_34449,N_34036,N_34138);
and U34450 (N_34450,N_34080,N_34237);
xnor U34451 (N_34451,N_34018,N_34097);
and U34452 (N_34452,N_34221,N_34063);
or U34453 (N_34453,N_34097,N_34196);
xnor U34454 (N_34454,N_34150,N_34002);
nand U34455 (N_34455,N_34244,N_34089);
xor U34456 (N_34456,N_34083,N_34023);
and U34457 (N_34457,N_34217,N_34027);
or U34458 (N_34458,N_34236,N_34028);
and U34459 (N_34459,N_34057,N_34145);
or U34460 (N_34460,N_34172,N_34193);
xnor U34461 (N_34461,N_34041,N_34081);
nor U34462 (N_34462,N_34003,N_34074);
nand U34463 (N_34463,N_34114,N_34045);
nor U34464 (N_34464,N_34038,N_34184);
and U34465 (N_34465,N_34021,N_34236);
nand U34466 (N_34466,N_34047,N_34141);
xnor U34467 (N_34467,N_34100,N_34031);
and U34468 (N_34468,N_34023,N_34187);
nor U34469 (N_34469,N_34062,N_34050);
xnor U34470 (N_34470,N_34160,N_34057);
or U34471 (N_34471,N_34058,N_34206);
and U34472 (N_34472,N_34105,N_34074);
xor U34473 (N_34473,N_34158,N_34018);
xor U34474 (N_34474,N_34199,N_34013);
nor U34475 (N_34475,N_34122,N_34131);
and U34476 (N_34476,N_34032,N_34141);
and U34477 (N_34477,N_34099,N_34092);
xor U34478 (N_34478,N_34161,N_34027);
or U34479 (N_34479,N_34034,N_34090);
xor U34480 (N_34480,N_34034,N_34116);
nor U34481 (N_34481,N_34171,N_34161);
and U34482 (N_34482,N_34165,N_34148);
xor U34483 (N_34483,N_34216,N_34227);
and U34484 (N_34484,N_34079,N_34069);
or U34485 (N_34485,N_34200,N_34153);
nand U34486 (N_34486,N_34013,N_34169);
or U34487 (N_34487,N_34083,N_34069);
nor U34488 (N_34488,N_34181,N_34004);
and U34489 (N_34489,N_34115,N_34230);
nor U34490 (N_34490,N_34186,N_34241);
xor U34491 (N_34491,N_34115,N_34193);
and U34492 (N_34492,N_34031,N_34164);
nand U34493 (N_34493,N_34006,N_34105);
or U34494 (N_34494,N_34161,N_34120);
nand U34495 (N_34495,N_34156,N_34231);
xor U34496 (N_34496,N_34246,N_34193);
or U34497 (N_34497,N_34155,N_34032);
and U34498 (N_34498,N_34235,N_34091);
xor U34499 (N_34499,N_34196,N_34041);
nor U34500 (N_34500,N_34252,N_34445);
nand U34501 (N_34501,N_34286,N_34338);
nor U34502 (N_34502,N_34315,N_34327);
xnor U34503 (N_34503,N_34446,N_34494);
nand U34504 (N_34504,N_34326,N_34388);
nand U34505 (N_34505,N_34390,N_34425);
or U34506 (N_34506,N_34323,N_34284);
nor U34507 (N_34507,N_34322,N_34316);
or U34508 (N_34508,N_34357,N_34370);
nor U34509 (N_34509,N_34337,N_34373);
nand U34510 (N_34510,N_34410,N_34385);
and U34511 (N_34511,N_34438,N_34378);
and U34512 (N_34512,N_34401,N_34417);
or U34513 (N_34513,N_34333,N_34456);
xor U34514 (N_34514,N_34282,N_34273);
nand U34515 (N_34515,N_34490,N_34259);
and U34516 (N_34516,N_34383,N_34266);
and U34517 (N_34517,N_34355,N_34300);
nor U34518 (N_34518,N_34421,N_34442);
and U34519 (N_34519,N_34423,N_34405);
nor U34520 (N_34520,N_34270,N_34339);
nand U34521 (N_34521,N_34346,N_34400);
or U34522 (N_34522,N_34257,N_34368);
and U34523 (N_34523,N_34317,N_34308);
nor U34524 (N_34524,N_34439,N_34476);
and U34525 (N_34525,N_34447,N_34454);
nand U34526 (N_34526,N_34342,N_34499);
xor U34527 (N_34527,N_34485,N_34455);
nand U34528 (N_34528,N_34471,N_34440);
xor U34529 (N_34529,N_34379,N_34354);
nor U34530 (N_34530,N_34467,N_34486);
nor U34531 (N_34531,N_34459,N_34360);
nor U34532 (N_34532,N_34458,N_34324);
xor U34533 (N_34533,N_34399,N_34416);
and U34534 (N_34534,N_34328,N_34433);
and U34535 (N_34535,N_34392,N_34488);
or U34536 (N_34536,N_34406,N_34466);
nor U34537 (N_34537,N_34325,N_34281);
and U34538 (N_34538,N_34268,N_34428);
or U34539 (N_34539,N_34457,N_34278);
and U34540 (N_34540,N_34267,N_34441);
nor U34541 (N_34541,N_34253,N_34404);
or U34542 (N_34542,N_34381,N_34277);
nor U34543 (N_34543,N_34394,N_34351);
or U34544 (N_34544,N_34255,N_34396);
and U34545 (N_34545,N_34345,N_34483);
nand U34546 (N_34546,N_34313,N_34465);
nand U34547 (N_34547,N_34319,N_34302);
and U34548 (N_34548,N_34375,N_34290);
nand U34549 (N_34549,N_34418,N_34256);
nor U34550 (N_34550,N_34484,N_34434);
xnor U34551 (N_34551,N_34320,N_34479);
nor U34552 (N_34552,N_34402,N_34292);
and U34553 (N_34553,N_34336,N_34419);
nor U34554 (N_34554,N_34264,N_34389);
nand U34555 (N_34555,N_34321,N_34301);
and U34556 (N_34556,N_34332,N_34464);
nor U34557 (N_34557,N_34391,N_34344);
nand U34558 (N_34558,N_34353,N_34371);
nand U34559 (N_34559,N_34387,N_34409);
xnor U34560 (N_34560,N_34276,N_34450);
nand U34561 (N_34561,N_34411,N_34359);
and U34562 (N_34562,N_34312,N_34377);
or U34563 (N_34563,N_34343,N_34271);
nand U34564 (N_34564,N_34285,N_34334);
nand U34565 (N_34565,N_34463,N_34384);
and U34566 (N_34566,N_34374,N_34427);
xnor U34567 (N_34567,N_34356,N_34453);
or U34568 (N_34568,N_34426,N_34489);
nor U34569 (N_34569,N_34364,N_34497);
or U34570 (N_34570,N_34251,N_34296);
and U34571 (N_34571,N_34358,N_34480);
nand U34572 (N_34572,N_34376,N_34291);
nand U34573 (N_34573,N_34297,N_34261);
nor U34574 (N_34574,N_34275,N_34289);
nand U34575 (N_34575,N_34495,N_34303);
or U34576 (N_34576,N_34491,N_34469);
nand U34577 (N_34577,N_34340,N_34318);
nand U34578 (N_34578,N_34395,N_34386);
or U34579 (N_34579,N_34420,N_34350);
xnor U34580 (N_34580,N_34260,N_34330);
and U34581 (N_34581,N_34444,N_34413);
xnor U34582 (N_34582,N_34470,N_34430);
xor U34583 (N_34583,N_34362,N_34424);
xor U34584 (N_34584,N_34279,N_34380);
and U34585 (N_34585,N_34492,N_34365);
nand U34586 (N_34586,N_34493,N_34452);
nand U34587 (N_34587,N_34478,N_34403);
xor U34588 (N_34588,N_34487,N_34397);
or U34589 (N_34589,N_34462,N_34481);
and U34590 (N_34590,N_34472,N_34361);
nand U34591 (N_34591,N_34460,N_34262);
or U34592 (N_34592,N_34432,N_34451);
nand U34593 (N_34593,N_34429,N_34306);
nor U34594 (N_34594,N_34274,N_34448);
or U34595 (N_34595,N_34367,N_34415);
nor U34596 (N_34596,N_34348,N_34349);
or U34597 (N_34597,N_34283,N_34422);
nor U34598 (N_34598,N_34294,N_34254);
or U34599 (N_34599,N_34449,N_34498);
and U34600 (N_34600,N_34372,N_34258);
nand U34601 (N_34601,N_34263,N_34461);
xor U34602 (N_34602,N_34496,N_34482);
xnor U34603 (N_34603,N_34443,N_34398);
xor U34604 (N_34604,N_34280,N_34287);
nand U34605 (N_34605,N_34293,N_34414);
nand U34606 (N_34606,N_34269,N_34369);
nor U34607 (N_34607,N_34437,N_34335);
or U34608 (N_34608,N_34295,N_34304);
and U34609 (N_34609,N_34298,N_34407);
nand U34610 (N_34610,N_34329,N_34477);
and U34611 (N_34611,N_34311,N_34265);
or U34612 (N_34612,N_34366,N_34436);
xnor U34613 (N_34613,N_34310,N_34314);
nor U34614 (N_34614,N_34288,N_34307);
xnor U34615 (N_34615,N_34431,N_34408);
or U34616 (N_34616,N_34468,N_34382);
nor U34617 (N_34617,N_34473,N_34474);
nand U34618 (N_34618,N_34250,N_34347);
nand U34619 (N_34619,N_34412,N_34475);
xnor U34620 (N_34620,N_34309,N_34393);
and U34621 (N_34621,N_34363,N_34305);
xor U34622 (N_34622,N_34435,N_34352);
and U34623 (N_34623,N_34272,N_34331);
and U34624 (N_34624,N_34299,N_34341);
or U34625 (N_34625,N_34409,N_34355);
nand U34626 (N_34626,N_34371,N_34254);
xnor U34627 (N_34627,N_34291,N_34266);
nor U34628 (N_34628,N_34294,N_34261);
xnor U34629 (N_34629,N_34333,N_34338);
and U34630 (N_34630,N_34407,N_34361);
nor U34631 (N_34631,N_34290,N_34433);
nand U34632 (N_34632,N_34364,N_34400);
nor U34633 (N_34633,N_34445,N_34461);
xnor U34634 (N_34634,N_34430,N_34386);
and U34635 (N_34635,N_34275,N_34324);
xor U34636 (N_34636,N_34430,N_34342);
and U34637 (N_34637,N_34327,N_34405);
nor U34638 (N_34638,N_34397,N_34267);
and U34639 (N_34639,N_34452,N_34433);
and U34640 (N_34640,N_34408,N_34498);
nor U34641 (N_34641,N_34284,N_34296);
nor U34642 (N_34642,N_34442,N_34478);
nand U34643 (N_34643,N_34416,N_34310);
xnor U34644 (N_34644,N_34423,N_34479);
and U34645 (N_34645,N_34341,N_34324);
or U34646 (N_34646,N_34254,N_34435);
nand U34647 (N_34647,N_34318,N_34349);
nand U34648 (N_34648,N_34400,N_34413);
and U34649 (N_34649,N_34465,N_34381);
nor U34650 (N_34650,N_34459,N_34422);
and U34651 (N_34651,N_34359,N_34320);
and U34652 (N_34652,N_34405,N_34471);
nor U34653 (N_34653,N_34365,N_34291);
or U34654 (N_34654,N_34402,N_34327);
or U34655 (N_34655,N_34298,N_34374);
or U34656 (N_34656,N_34462,N_34373);
nand U34657 (N_34657,N_34355,N_34317);
nor U34658 (N_34658,N_34402,N_34496);
and U34659 (N_34659,N_34417,N_34352);
nor U34660 (N_34660,N_34470,N_34398);
xnor U34661 (N_34661,N_34339,N_34315);
and U34662 (N_34662,N_34269,N_34457);
nand U34663 (N_34663,N_34272,N_34364);
xnor U34664 (N_34664,N_34250,N_34483);
and U34665 (N_34665,N_34406,N_34495);
nor U34666 (N_34666,N_34482,N_34417);
nand U34667 (N_34667,N_34272,N_34273);
nor U34668 (N_34668,N_34361,N_34496);
or U34669 (N_34669,N_34393,N_34275);
nand U34670 (N_34670,N_34294,N_34390);
or U34671 (N_34671,N_34257,N_34307);
or U34672 (N_34672,N_34292,N_34351);
xnor U34673 (N_34673,N_34352,N_34408);
and U34674 (N_34674,N_34294,N_34385);
or U34675 (N_34675,N_34301,N_34390);
or U34676 (N_34676,N_34429,N_34255);
xnor U34677 (N_34677,N_34330,N_34347);
xor U34678 (N_34678,N_34437,N_34491);
nor U34679 (N_34679,N_34430,N_34395);
and U34680 (N_34680,N_34488,N_34254);
nand U34681 (N_34681,N_34344,N_34342);
or U34682 (N_34682,N_34365,N_34310);
nor U34683 (N_34683,N_34432,N_34360);
and U34684 (N_34684,N_34317,N_34469);
xnor U34685 (N_34685,N_34452,N_34375);
or U34686 (N_34686,N_34257,N_34286);
or U34687 (N_34687,N_34314,N_34493);
nor U34688 (N_34688,N_34302,N_34481);
nand U34689 (N_34689,N_34393,N_34353);
or U34690 (N_34690,N_34309,N_34361);
nand U34691 (N_34691,N_34266,N_34459);
or U34692 (N_34692,N_34314,N_34346);
nor U34693 (N_34693,N_34307,N_34469);
xnor U34694 (N_34694,N_34407,N_34275);
nand U34695 (N_34695,N_34456,N_34438);
or U34696 (N_34696,N_34422,N_34423);
xnor U34697 (N_34697,N_34397,N_34439);
and U34698 (N_34698,N_34251,N_34276);
xor U34699 (N_34699,N_34437,N_34383);
nand U34700 (N_34700,N_34281,N_34363);
and U34701 (N_34701,N_34433,N_34439);
nor U34702 (N_34702,N_34292,N_34344);
and U34703 (N_34703,N_34455,N_34263);
xor U34704 (N_34704,N_34318,N_34416);
nand U34705 (N_34705,N_34440,N_34456);
xnor U34706 (N_34706,N_34388,N_34479);
nand U34707 (N_34707,N_34350,N_34336);
nor U34708 (N_34708,N_34365,N_34333);
and U34709 (N_34709,N_34471,N_34304);
and U34710 (N_34710,N_34397,N_34466);
nor U34711 (N_34711,N_34433,N_34368);
xor U34712 (N_34712,N_34393,N_34290);
nand U34713 (N_34713,N_34461,N_34380);
or U34714 (N_34714,N_34434,N_34350);
nand U34715 (N_34715,N_34286,N_34392);
xor U34716 (N_34716,N_34331,N_34325);
nor U34717 (N_34717,N_34347,N_34276);
or U34718 (N_34718,N_34339,N_34395);
xnor U34719 (N_34719,N_34393,N_34366);
nand U34720 (N_34720,N_34385,N_34362);
or U34721 (N_34721,N_34335,N_34370);
nor U34722 (N_34722,N_34400,N_34398);
xor U34723 (N_34723,N_34451,N_34271);
xnor U34724 (N_34724,N_34302,N_34401);
xor U34725 (N_34725,N_34315,N_34392);
nand U34726 (N_34726,N_34381,N_34261);
xnor U34727 (N_34727,N_34257,N_34476);
xnor U34728 (N_34728,N_34292,N_34404);
and U34729 (N_34729,N_34289,N_34292);
nor U34730 (N_34730,N_34479,N_34285);
nand U34731 (N_34731,N_34392,N_34319);
or U34732 (N_34732,N_34299,N_34429);
or U34733 (N_34733,N_34310,N_34418);
or U34734 (N_34734,N_34438,N_34411);
nor U34735 (N_34735,N_34433,N_34362);
xnor U34736 (N_34736,N_34259,N_34418);
or U34737 (N_34737,N_34261,N_34416);
and U34738 (N_34738,N_34338,N_34375);
nor U34739 (N_34739,N_34406,N_34304);
or U34740 (N_34740,N_34345,N_34330);
or U34741 (N_34741,N_34384,N_34440);
nor U34742 (N_34742,N_34379,N_34314);
xnor U34743 (N_34743,N_34321,N_34470);
or U34744 (N_34744,N_34398,N_34410);
and U34745 (N_34745,N_34432,N_34404);
nor U34746 (N_34746,N_34400,N_34463);
or U34747 (N_34747,N_34276,N_34368);
nand U34748 (N_34748,N_34373,N_34285);
or U34749 (N_34749,N_34423,N_34317);
xor U34750 (N_34750,N_34657,N_34649);
nor U34751 (N_34751,N_34640,N_34598);
nor U34752 (N_34752,N_34638,N_34578);
nor U34753 (N_34753,N_34517,N_34548);
xnor U34754 (N_34754,N_34702,N_34632);
and U34755 (N_34755,N_34519,N_34642);
nand U34756 (N_34756,N_34583,N_34749);
nor U34757 (N_34757,N_34585,N_34500);
nand U34758 (N_34758,N_34626,N_34668);
xnor U34759 (N_34759,N_34603,N_34740);
or U34760 (N_34760,N_34606,N_34656);
xor U34761 (N_34761,N_34712,N_34727);
nor U34762 (N_34762,N_34644,N_34741);
or U34763 (N_34763,N_34501,N_34611);
or U34764 (N_34764,N_34739,N_34667);
xor U34765 (N_34765,N_34573,N_34680);
or U34766 (N_34766,N_34716,N_34708);
xor U34767 (N_34767,N_34562,N_34694);
xor U34768 (N_34768,N_34736,N_34744);
nand U34769 (N_34769,N_34648,N_34567);
and U34770 (N_34770,N_34590,N_34745);
or U34771 (N_34771,N_34618,N_34600);
nand U34772 (N_34772,N_34747,N_34614);
xnor U34773 (N_34773,N_34730,N_34544);
or U34774 (N_34774,N_34524,N_34564);
and U34775 (N_34775,N_34700,N_34530);
nor U34776 (N_34776,N_34684,N_34738);
nand U34777 (N_34777,N_34654,N_34610);
or U34778 (N_34778,N_34577,N_34613);
or U34779 (N_34779,N_34525,N_34677);
xor U34780 (N_34780,N_34529,N_34707);
or U34781 (N_34781,N_34591,N_34737);
xor U34782 (N_34782,N_34726,N_34629);
nor U34783 (N_34783,N_34622,N_34746);
xor U34784 (N_34784,N_34575,N_34572);
or U34785 (N_34785,N_34709,N_34602);
nor U34786 (N_34786,N_34513,N_34508);
and U34787 (N_34787,N_34701,N_34568);
nor U34788 (N_34788,N_34710,N_34691);
nor U34789 (N_34789,N_34672,N_34646);
or U34790 (N_34790,N_34506,N_34604);
or U34791 (N_34791,N_34621,N_34671);
or U34792 (N_34792,N_34687,N_34532);
xor U34793 (N_34793,N_34633,N_34725);
xnor U34794 (N_34794,N_34593,N_34509);
xnor U34795 (N_34795,N_34627,N_34516);
xor U34796 (N_34796,N_34503,N_34605);
nand U34797 (N_34797,N_34675,N_34673);
and U34798 (N_34798,N_34689,N_34540);
nor U34799 (N_34799,N_34734,N_34601);
and U34800 (N_34800,N_34713,N_34523);
xor U34801 (N_34801,N_34527,N_34594);
and U34802 (N_34802,N_34652,N_34696);
nand U34803 (N_34803,N_34674,N_34690);
nor U34804 (N_34804,N_34715,N_34528);
or U34805 (N_34805,N_34555,N_34685);
and U34806 (N_34806,N_34561,N_34559);
and U34807 (N_34807,N_34623,N_34514);
or U34808 (N_34808,N_34717,N_34520);
xor U34809 (N_34809,N_34609,N_34550);
or U34810 (N_34810,N_34661,N_34641);
nand U34811 (N_34811,N_34569,N_34551);
and U34812 (N_34812,N_34663,N_34732);
and U34813 (N_34813,N_34571,N_34616);
or U34814 (N_34814,N_34721,N_34659);
and U34815 (N_34815,N_34615,N_34580);
xor U34816 (N_34816,N_34536,N_34719);
xnor U34817 (N_34817,N_34537,N_34546);
and U34818 (N_34818,N_34669,N_34660);
or U34819 (N_34819,N_34699,N_34693);
or U34820 (N_34820,N_34556,N_34733);
nor U34821 (N_34821,N_34705,N_34552);
and U34822 (N_34822,N_34724,N_34534);
or U34823 (N_34823,N_34542,N_34698);
and U34824 (N_34824,N_34570,N_34630);
xor U34825 (N_34825,N_34612,N_34723);
nand U34826 (N_34826,N_34547,N_34579);
xor U34827 (N_34827,N_34566,N_34664);
nand U34828 (N_34828,N_34666,N_34505);
or U34829 (N_34829,N_34545,N_34620);
nor U34830 (N_34830,N_34617,N_34703);
or U34831 (N_34831,N_34718,N_34599);
xor U34832 (N_34832,N_34711,N_34643);
nand U34833 (N_34833,N_34565,N_34683);
and U34834 (N_34834,N_34742,N_34543);
nand U34835 (N_34835,N_34512,N_34589);
nor U34836 (N_34836,N_34706,N_34686);
nand U34837 (N_34837,N_34631,N_34697);
xor U34838 (N_34838,N_34587,N_34581);
nor U34839 (N_34839,N_34541,N_34533);
nor U34840 (N_34840,N_34679,N_34522);
xor U34841 (N_34841,N_34681,N_34607);
xor U34842 (N_34842,N_34743,N_34538);
nand U34843 (N_34843,N_34720,N_34658);
nand U34844 (N_34844,N_34692,N_34518);
or U34845 (N_34845,N_34504,N_34653);
and U34846 (N_34846,N_34704,N_34557);
or U34847 (N_34847,N_34507,N_34553);
and U34848 (N_34848,N_34574,N_34729);
nand U34849 (N_34849,N_34676,N_34558);
nor U34850 (N_34850,N_34526,N_34597);
xor U34851 (N_34851,N_34695,N_34624);
nor U34852 (N_34852,N_34678,N_34651);
nand U34853 (N_34853,N_34728,N_34735);
nand U34854 (N_34854,N_34628,N_34662);
nand U34855 (N_34855,N_34521,N_34655);
or U34856 (N_34856,N_34722,N_34634);
or U34857 (N_34857,N_34554,N_34665);
nand U34858 (N_34858,N_34586,N_34588);
xnor U34859 (N_34859,N_34637,N_34584);
or U34860 (N_34860,N_34502,N_34639);
and U34861 (N_34861,N_34647,N_34531);
nor U34862 (N_34862,N_34625,N_34682);
nand U34863 (N_34863,N_34619,N_34560);
xnor U34864 (N_34864,N_34635,N_34595);
and U34865 (N_34865,N_34539,N_34714);
nor U34866 (N_34866,N_34645,N_34688);
xnor U34867 (N_34867,N_34510,N_34511);
nand U34868 (N_34868,N_34748,N_34592);
nor U34869 (N_34869,N_34650,N_34670);
or U34870 (N_34870,N_34596,N_34576);
or U34871 (N_34871,N_34582,N_34636);
or U34872 (N_34872,N_34608,N_34515);
nand U34873 (N_34873,N_34535,N_34563);
nand U34874 (N_34874,N_34731,N_34549);
and U34875 (N_34875,N_34531,N_34512);
nand U34876 (N_34876,N_34509,N_34512);
and U34877 (N_34877,N_34712,N_34522);
nor U34878 (N_34878,N_34630,N_34679);
and U34879 (N_34879,N_34566,N_34667);
nor U34880 (N_34880,N_34637,N_34505);
nand U34881 (N_34881,N_34551,N_34528);
nor U34882 (N_34882,N_34507,N_34661);
nor U34883 (N_34883,N_34620,N_34578);
nand U34884 (N_34884,N_34603,N_34590);
nor U34885 (N_34885,N_34638,N_34676);
nor U34886 (N_34886,N_34533,N_34728);
or U34887 (N_34887,N_34619,N_34692);
nor U34888 (N_34888,N_34681,N_34648);
nor U34889 (N_34889,N_34621,N_34572);
xor U34890 (N_34890,N_34660,N_34623);
nand U34891 (N_34891,N_34706,N_34616);
nor U34892 (N_34892,N_34516,N_34508);
or U34893 (N_34893,N_34635,N_34567);
or U34894 (N_34894,N_34643,N_34585);
or U34895 (N_34895,N_34506,N_34726);
or U34896 (N_34896,N_34718,N_34503);
xor U34897 (N_34897,N_34546,N_34729);
or U34898 (N_34898,N_34616,N_34739);
or U34899 (N_34899,N_34664,N_34676);
or U34900 (N_34900,N_34521,N_34740);
nand U34901 (N_34901,N_34600,N_34682);
nor U34902 (N_34902,N_34547,N_34622);
nor U34903 (N_34903,N_34565,N_34604);
and U34904 (N_34904,N_34689,N_34622);
xnor U34905 (N_34905,N_34545,N_34532);
nor U34906 (N_34906,N_34701,N_34566);
nand U34907 (N_34907,N_34526,N_34660);
nand U34908 (N_34908,N_34563,N_34700);
nor U34909 (N_34909,N_34695,N_34736);
and U34910 (N_34910,N_34573,N_34719);
or U34911 (N_34911,N_34512,N_34533);
xor U34912 (N_34912,N_34704,N_34745);
nor U34913 (N_34913,N_34722,N_34637);
and U34914 (N_34914,N_34570,N_34647);
nor U34915 (N_34915,N_34615,N_34587);
nor U34916 (N_34916,N_34715,N_34570);
and U34917 (N_34917,N_34646,N_34559);
nor U34918 (N_34918,N_34669,N_34540);
or U34919 (N_34919,N_34592,N_34603);
xnor U34920 (N_34920,N_34741,N_34630);
or U34921 (N_34921,N_34548,N_34574);
nand U34922 (N_34922,N_34665,N_34699);
and U34923 (N_34923,N_34517,N_34716);
and U34924 (N_34924,N_34675,N_34605);
xor U34925 (N_34925,N_34580,N_34734);
and U34926 (N_34926,N_34689,N_34650);
or U34927 (N_34927,N_34556,N_34636);
or U34928 (N_34928,N_34581,N_34625);
and U34929 (N_34929,N_34590,N_34631);
and U34930 (N_34930,N_34528,N_34712);
nor U34931 (N_34931,N_34646,N_34520);
nor U34932 (N_34932,N_34668,N_34507);
xnor U34933 (N_34933,N_34700,N_34594);
or U34934 (N_34934,N_34630,N_34616);
nor U34935 (N_34935,N_34507,N_34550);
xnor U34936 (N_34936,N_34507,N_34555);
or U34937 (N_34937,N_34531,N_34635);
or U34938 (N_34938,N_34572,N_34576);
xnor U34939 (N_34939,N_34686,N_34684);
nand U34940 (N_34940,N_34501,N_34586);
or U34941 (N_34941,N_34548,N_34557);
and U34942 (N_34942,N_34728,N_34657);
xor U34943 (N_34943,N_34525,N_34712);
and U34944 (N_34944,N_34597,N_34574);
nor U34945 (N_34945,N_34553,N_34593);
xnor U34946 (N_34946,N_34555,N_34727);
and U34947 (N_34947,N_34628,N_34679);
xor U34948 (N_34948,N_34733,N_34537);
and U34949 (N_34949,N_34624,N_34609);
and U34950 (N_34950,N_34593,N_34526);
or U34951 (N_34951,N_34692,N_34655);
and U34952 (N_34952,N_34568,N_34524);
nand U34953 (N_34953,N_34529,N_34720);
nand U34954 (N_34954,N_34587,N_34569);
and U34955 (N_34955,N_34648,N_34619);
or U34956 (N_34956,N_34734,N_34648);
xor U34957 (N_34957,N_34613,N_34570);
xnor U34958 (N_34958,N_34522,N_34562);
nor U34959 (N_34959,N_34607,N_34585);
and U34960 (N_34960,N_34643,N_34570);
nor U34961 (N_34961,N_34504,N_34514);
and U34962 (N_34962,N_34678,N_34572);
and U34963 (N_34963,N_34680,N_34720);
xor U34964 (N_34964,N_34609,N_34589);
nand U34965 (N_34965,N_34682,N_34718);
xor U34966 (N_34966,N_34666,N_34642);
and U34967 (N_34967,N_34743,N_34679);
xor U34968 (N_34968,N_34594,N_34730);
nor U34969 (N_34969,N_34580,N_34710);
nor U34970 (N_34970,N_34723,N_34602);
xnor U34971 (N_34971,N_34556,N_34543);
nor U34972 (N_34972,N_34591,N_34588);
and U34973 (N_34973,N_34698,N_34529);
nor U34974 (N_34974,N_34527,N_34531);
nor U34975 (N_34975,N_34502,N_34688);
nor U34976 (N_34976,N_34633,N_34599);
nor U34977 (N_34977,N_34527,N_34671);
or U34978 (N_34978,N_34501,N_34509);
or U34979 (N_34979,N_34535,N_34736);
nor U34980 (N_34980,N_34587,N_34661);
and U34981 (N_34981,N_34518,N_34587);
nand U34982 (N_34982,N_34654,N_34591);
nand U34983 (N_34983,N_34561,N_34504);
nor U34984 (N_34984,N_34703,N_34520);
or U34985 (N_34985,N_34718,N_34656);
and U34986 (N_34986,N_34739,N_34642);
or U34987 (N_34987,N_34697,N_34736);
or U34988 (N_34988,N_34540,N_34501);
nor U34989 (N_34989,N_34515,N_34640);
and U34990 (N_34990,N_34706,N_34735);
or U34991 (N_34991,N_34721,N_34617);
and U34992 (N_34992,N_34530,N_34597);
xnor U34993 (N_34993,N_34622,N_34579);
nand U34994 (N_34994,N_34513,N_34641);
or U34995 (N_34995,N_34597,N_34664);
xor U34996 (N_34996,N_34588,N_34702);
xnor U34997 (N_34997,N_34592,N_34660);
or U34998 (N_34998,N_34602,N_34511);
nand U34999 (N_34999,N_34648,N_34548);
or U35000 (N_35000,N_34884,N_34880);
nand U35001 (N_35001,N_34864,N_34927);
xnor U35002 (N_35002,N_34854,N_34947);
xor U35003 (N_35003,N_34808,N_34761);
or U35004 (N_35004,N_34797,N_34815);
xnor U35005 (N_35005,N_34943,N_34857);
and U35006 (N_35006,N_34801,N_34922);
xor U35007 (N_35007,N_34931,N_34822);
nor U35008 (N_35008,N_34968,N_34982);
nor U35009 (N_35009,N_34755,N_34890);
nand U35010 (N_35010,N_34772,N_34987);
xnor U35011 (N_35011,N_34946,N_34830);
xor U35012 (N_35012,N_34877,N_34777);
and U35013 (N_35013,N_34984,N_34925);
or U35014 (N_35014,N_34969,N_34769);
nand U35015 (N_35015,N_34868,N_34846);
nand U35016 (N_35016,N_34985,N_34887);
nand U35017 (N_35017,N_34805,N_34926);
or U35018 (N_35018,N_34876,N_34756);
nor U35019 (N_35019,N_34998,N_34891);
and U35020 (N_35020,N_34763,N_34869);
nor U35021 (N_35021,N_34950,N_34765);
nand U35022 (N_35022,N_34752,N_34886);
nor U35023 (N_35023,N_34941,N_34767);
xnor U35024 (N_35024,N_34949,N_34849);
nand U35025 (N_35025,N_34821,N_34974);
nand U35026 (N_35026,N_34782,N_34972);
nor U35027 (N_35027,N_34806,N_34902);
nand U35028 (N_35028,N_34781,N_34938);
nor U35029 (N_35029,N_34778,N_34818);
xnor U35030 (N_35030,N_34910,N_34906);
nor U35031 (N_35031,N_34804,N_34836);
nor U35032 (N_35032,N_34934,N_34800);
xor U35033 (N_35033,N_34850,N_34856);
nor U35034 (N_35034,N_34990,N_34863);
nor U35035 (N_35035,N_34776,N_34954);
and U35036 (N_35036,N_34841,N_34758);
xnor U35037 (N_35037,N_34956,N_34770);
nor U35038 (N_35038,N_34789,N_34811);
or U35039 (N_35039,N_34795,N_34920);
and U35040 (N_35040,N_34895,N_34948);
or U35041 (N_35041,N_34855,N_34935);
and U35042 (N_35042,N_34843,N_34918);
and U35043 (N_35043,N_34989,N_34784);
xor U35044 (N_35044,N_34944,N_34757);
nor U35045 (N_35045,N_34996,N_34792);
and U35046 (N_35046,N_34958,N_34967);
and U35047 (N_35047,N_34865,N_34966);
or U35048 (N_35048,N_34889,N_34867);
nand U35049 (N_35049,N_34997,N_34764);
or U35050 (N_35050,N_34973,N_34881);
and U35051 (N_35051,N_34766,N_34909);
and U35052 (N_35052,N_34914,N_34845);
or U35053 (N_35053,N_34903,N_34754);
nor U35054 (N_35054,N_34970,N_34773);
nor U35055 (N_35055,N_34835,N_34838);
or U35056 (N_35056,N_34993,N_34809);
xnor U35057 (N_35057,N_34783,N_34951);
nor U35058 (N_35058,N_34957,N_34751);
xor U35059 (N_35059,N_34812,N_34753);
nand U35060 (N_35060,N_34768,N_34904);
and U35061 (N_35061,N_34759,N_34917);
or U35062 (N_35062,N_34991,N_34832);
nand U35063 (N_35063,N_34921,N_34977);
nor U35064 (N_35064,N_34813,N_34978);
nor U35065 (N_35065,N_34839,N_34919);
nand U35066 (N_35066,N_34882,N_34871);
and U35067 (N_35067,N_34858,N_34915);
nand U35068 (N_35068,N_34963,N_34840);
and U35069 (N_35069,N_34936,N_34851);
xor U35070 (N_35070,N_34897,N_34760);
or U35071 (N_35071,N_34975,N_34888);
and U35072 (N_35072,N_34861,N_34774);
xnor U35073 (N_35073,N_34872,N_34916);
or U35074 (N_35074,N_34962,N_34816);
xnor U35075 (N_35075,N_34896,N_34912);
and U35076 (N_35076,N_34873,N_34823);
xnor U35077 (N_35077,N_34893,N_34785);
nor U35078 (N_35078,N_34847,N_34908);
nand U35079 (N_35079,N_34810,N_34940);
nor U35080 (N_35080,N_34965,N_34961);
or U35081 (N_35081,N_34825,N_34979);
and U35082 (N_35082,N_34803,N_34786);
xnor U35083 (N_35083,N_34798,N_34999);
xor U35084 (N_35084,N_34976,N_34820);
nor U35085 (N_35085,N_34894,N_34953);
or U35086 (N_35086,N_34964,N_34874);
xnor U35087 (N_35087,N_34862,N_34992);
and U35088 (N_35088,N_34842,N_34794);
nand U35089 (N_35089,N_34980,N_34955);
nor U35090 (N_35090,N_34885,N_34945);
nor U35091 (N_35091,N_34911,N_34878);
xor U35092 (N_35092,N_34848,N_34762);
and U35093 (N_35093,N_34837,N_34929);
or U35094 (N_35094,N_34853,N_34779);
and U35095 (N_35095,N_34824,N_34807);
nor U35096 (N_35096,N_34960,N_34787);
nor U35097 (N_35097,N_34892,N_34870);
nand U35098 (N_35098,N_34826,N_34796);
nand U35099 (N_35099,N_34994,N_34900);
and U35100 (N_35100,N_34817,N_34750);
nor U35101 (N_35101,N_34829,N_34883);
and U35102 (N_35102,N_34937,N_34827);
and U35103 (N_35103,N_34942,N_34905);
and U35104 (N_35104,N_34860,N_34831);
nor U35105 (N_35105,N_34802,N_34907);
or U35106 (N_35106,N_34986,N_34952);
nand U35107 (N_35107,N_34866,N_34923);
xor U35108 (N_35108,N_34928,N_34988);
or U35109 (N_35109,N_34981,N_34859);
or U35110 (N_35110,N_34932,N_34793);
or U35111 (N_35111,N_34799,N_34775);
or U35112 (N_35112,N_34771,N_34833);
or U35113 (N_35113,N_34875,N_34995);
nor U35114 (N_35114,N_34780,N_34852);
or U35115 (N_35115,N_34844,N_34959);
nor U35116 (N_35116,N_34901,N_34924);
nand U35117 (N_35117,N_34814,N_34913);
nand U35118 (N_35118,N_34791,N_34971);
and U35119 (N_35119,N_34879,N_34788);
xor U35120 (N_35120,N_34828,N_34898);
or U35121 (N_35121,N_34790,N_34834);
xnor U35122 (N_35122,N_34933,N_34983);
xnor U35123 (N_35123,N_34899,N_34819);
or U35124 (N_35124,N_34930,N_34939);
and U35125 (N_35125,N_34858,N_34920);
or U35126 (N_35126,N_34765,N_34824);
xor U35127 (N_35127,N_34942,N_34860);
or U35128 (N_35128,N_34885,N_34790);
nor U35129 (N_35129,N_34941,N_34964);
nor U35130 (N_35130,N_34894,N_34984);
or U35131 (N_35131,N_34934,N_34858);
nor U35132 (N_35132,N_34993,N_34970);
nand U35133 (N_35133,N_34978,N_34931);
nand U35134 (N_35134,N_34840,N_34835);
and U35135 (N_35135,N_34879,N_34888);
or U35136 (N_35136,N_34790,N_34983);
or U35137 (N_35137,N_34884,N_34991);
nor U35138 (N_35138,N_34992,N_34809);
nand U35139 (N_35139,N_34933,N_34878);
nand U35140 (N_35140,N_34977,N_34816);
or U35141 (N_35141,N_34990,N_34950);
and U35142 (N_35142,N_34809,N_34751);
xor U35143 (N_35143,N_34950,N_34854);
nor U35144 (N_35144,N_34793,N_34766);
nor U35145 (N_35145,N_34961,N_34854);
xor U35146 (N_35146,N_34908,N_34964);
xor U35147 (N_35147,N_34815,N_34853);
xor U35148 (N_35148,N_34924,N_34931);
and U35149 (N_35149,N_34861,N_34941);
xor U35150 (N_35150,N_34821,N_34818);
and U35151 (N_35151,N_34950,N_34949);
nor U35152 (N_35152,N_34995,N_34963);
xnor U35153 (N_35153,N_34938,N_34857);
nor U35154 (N_35154,N_34940,N_34809);
and U35155 (N_35155,N_34886,N_34757);
or U35156 (N_35156,N_34877,N_34868);
xor U35157 (N_35157,N_34966,N_34883);
xor U35158 (N_35158,N_34822,N_34861);
nor U35159 (N_35159,N_34948,N_34768);
nand U35160 (N_35160,N_34784,N_34841);
and U35161 (N_35161,N_34794,N_34950);
or U35162 (N_35162,N_34802,N_34896);
nand U35163 (N_35163,N_34891,N_34973);
nor U35164 (N_35164,N_34863,N_34874);
nand U35165 (N_35165,N_34824,N_34897);
xnor U35166 (N_35166,N_34838,N_34887);
or U35167 (N_35167,N_34930,N_34957);
and U35168 (N_35168,N_34875,N_34834);
nor U35169 (N_35169,N_34826,N_34979);
nand U35170 (N_35170,N_34982,N_34971);
or U35171 (N_35171,N_34964,N_34871);
xor U35172 (N_35172,N_34954,N_34972);
or U35173 (N_35173,N_34974,N_34764);
or U35174 (N_35174,N_34921,N_34801);
or U35175 (N_35175,N_34824,N_34912);
nor U35176 (N_35176,N_34923,N_34841);
nor U35177 (N_35177,N_34960,N_34840);
nor U35178 (N_35178,N_34757,N_34965);
and U35179 (N_35179,N_34962,N_34846);
and U35180 (N_35180,N_34873,N_34834);
xor U35181 (N_35181,N_34961,N_34960);
nor U35182 (N_35182,N_34827,N_34907);
xor U35183 (N_35183,N_34891,N_34924);
nand U35184 (N_35184,N_34899,N_34825);
nand U35185 (N_35185,N_34817,N_34846);
or U35186 (N_35186,N_34825,N_34997);
xor U35187 (N_35187,N_34876,N_34775);
nor U35188 (N_35188,N_34883,N_34954);
nand U35189 (N_35189,N_34942,N_34890);
nor U35190 (N_35190,N_34994,N_34862);
nand U35191 (N_35191,N_34919,N_34976);
nand U35192 (N_35192,N_34985,N_34766);
and U35193 (N_35193,N_34986,N_34849);
xnor U35194 (N_35194,N_34906,N_34822);
nor U35195 (N_35195,N_34999,N_34856);
nand U35196 (N_35196,N_34958,N_34842);
nor U35197 (N_35197,N_34751,N_34767);
nand U35198 (N_35198,N_34981,N_34820);
nor U35199 (N_35199,N_34878,N_34941);
xnor U35200 (N_35200,N_34993,N_34829);
and U35201 (N_35201,N_34833,N_34854);
or U35202 (N_35202,N_34756,N_34911);
xor U35203 (N_35203,N_34768,N_34759);
or U35204 (N_35204,N_34760,N_34867);
or U35205 (N_35205,N_34760,N_34845);
and U35206 (N_35206,N_34874,N_34950);
xnor U35207 (N_35207,N_34841,N_34791);
nand U35208 (N_35208,N_34913,N_34861);
and U35209 (N_35209,N_34767,N_34844);
xor U35210 (N_35210,N_34879,N_34797);
and U35211 (N_35211,N_34915,N_34976);
xor U35212 (N_35212,N_34832,N_34771);
or U35213 (N_35213,N_34926,N_34828);
nor U35214 (N_35214,N_34957,N_34959);
nor U35215 (N_35215,N_34836,N_34822);
or U35216 (N_35216,N_34853,N_34929);
xor U35217 (N_35217,N_34810,N_34945);
or U35218 (N_35218,N_34991,N_34872);
nor U35219 (N_35219,N_34837,N_34877);
and U35220 (N_35220,N_34993,N_34827);
or U35221 (N_35221,N_34973,N_34779);
nand U35222 (N_35222,N_34796,N_34937);
nor U35223 (N_35223,N_34911,N_34785);
nor U35224 (N_35224,N_34899,N_34922);
nor U35225 (N_35225,N_34773,N_34807);
or U35226 (N_35226,N_34938,N_34831);
and U35227 (N_35227,N_34882,N_34839);
and U35228 (N_35228,N_34792,N_34797);
xnor U35229 (N_35229,N_34986,N_34866);
xnor U35230 (N_35230,N_34810,N_34799);
nor U35231 (N_35231,N_34910,N_34836);
or U35232 (N_35232,N_34820,N_34933);
xor U35233 (N_35233,N_34906,N_34928);
or U35234 (N_35234,N_34899,N_34913);
xor U35235 (N_35235,N_34930,N_34755);
nor U35236 (N_35236,N_34855,N_34802);
xor U35237 (N_35237,N_34888,N_34873);
nor U35238 (N_35238,N_34891,N_34954);
nand U35239 (N_35239,N_34818,N_34987);
xor U35240 (N_35240,N_34999,N_34773);
nor U35241 (N_35241,N_34990,N_34799);
or U35242 (N_35242,N_34969,N_34791);
xnor U35243 (N_35243,N_34993,N_34870);
or U35244 (N_35244,N_34940,N_34796);
nand U35245 (N_35245,N_34932,N_34758);
nor U35246 (N_35246,N_34962,N_34983);
or U35247 (N_35247,N_34767,N_34838);
or U35248 (N_35248,N_34978,N_34797);
xor U35249 (N_35249,N_34799,N_34757);
and U35250 (N_35250,N_35232,N_35219);
nand U35251 (N_35251,N_35248,N_35018);
nand U35252 (N_35252,N_35069,N_35187);
nor U35253 (N_35253,N_35234,N_35150);
nand U35254 (N_35254,N_35200,N_35146);
xnor U35255 (N_35255,N_35208,N_35129);
nand U35256 (N_35256,N_35089,N_35025);
xor U35257 (N_35257,N_35010,N_35065);
and U35258 (N_35258,N_35225,N_35206);
nand U35259 (N_35259,N_35212,N_35218);
or U35260 (N_35260,N_35107,N_35075);
xnor U35261 (N_35261,N_35229,N_35013);
and U35262 (N_35262,N_35245,N_35241);
or U35263 (N_35263,N_35246,N_35035);
nand U35264 (N_35264,N_35034,N_35004);
xor U35265 (N_35265,N_35233,N_35163);
nand U35266 (N_35266,N_35043,N_35153);
nor U35267 (N_35267,N_35030,N_35249);
nand U35268 (N_35268,N_35012,N_35160);
and U35269 (N_35269,N_35211,N_35120);
xor U35270 (N_35270,N_35175,N_35024);
xor U35271 (N_35271,N_35151,N_35164);
and U35272 (N_35272,N_35139,N_35056);
xnor U35273 (N_35273,N_35228,N_35230);
nand U35274 (N_35274,N_35115,N_35032);
nor U35275 (N_35275,N_35029,N_35008);
nand U35276 (N_35276,N_35040,N_35198);
nor U35277 (N_35277,N_35223,N_35201);
and U35278 (N_35278,N_35171,N_35240);
nor U35279 (N_35279,N_35048,N_35041);
nand U35280 (N_35280,N_35205,N_35042);
nand U35281 (N_35281,N_35131,N_35162);
nor U35282 (N_35282,N_35173,N_35085);
and U35283 (N_35283,N_35006,N_35105);
nand U35284 (N_35284,N_35189,N_35176);
xnor U35285 (N_35285,N_35074,N_35058);
and U35286 (N_35286,N_35028,N_35203);
nor U35287 (N_35287,N_35183,N_35033);
xnor U35288 (N_35288,N_35076,N_35073);
nand U35289 (N_35289,N_35207,N_35195);
and U35290 (N_35290,N_35098,N_35185);
and U35291 (N_35291,N_35236,N_35086);
or U35292 (N_35292,N_35093,N_35192);
nand U35293 (N_35293,N_35143,N_35050);
or U35294 (N_35294,N_35147,N_35216);
xor U35295 (N_35295,N_35044,N_35077);
xor U35296 (N_35296,N_35017,N_35156);
xor U35297 (N_35297,N_35088,N_35049);
or U35298 (N_35298,N_35174,N_35170);
or U35299 (N_35299,N_35047,N_35237);
nor U35300 (N_35300,N_35109,N_35190);
and U35301 (N_35301,N_35111,N_35217);
nor U35302 (N_35302,N_35031,N_35118);
and U35303 (N_35303,N_35071,N_35157);
and U35304 (N_35304,N_35178,N_35224);
xnor U35305 (N_35305,N_35130,N_35122);
nor U35306 (N_35306,N_35081,N_35113);
xnor U35307 (N_35307,N_35036,N_35072);
xnor U35308 (N_35308,N_35124,N_35084);
nor U35309 (N_35309,N_35144,N_35177);
or U35310 (N_35310,N_35083,N_35096);
or U35311 (N_35311,N_35213,N_35000);
and U35312 (N_35312,N_35057,N_35242);
or U35313 (N_35313,N_35243,N_35104);
or U35314 (N_35314,N_35142,N_35054);
nor U35315 (N_35315,N_35125,N_35166);
nor U35316 (N_35316,N_35014,N_35210);
nor U35317 (N_35317,N_35204,N_35051);
or U35318 (N_35318,N_35220,N_35094);
nor U35319 (N_35319,N_35019,N_35214);
or U35320 (N_35320,N_35001,N_35134);
xnor U35321 (N_35321,N_35137,N_35114);
nand U35322 (N_35322,N_35082,N_35168);
and U35323 (N_35323,N_35095,N_35064);
nand U35324 (N_35324,N_35127,N_35126);
or U35325 (N_35325,N_35103,N_35097);
and U35326 (N_35326,N_35116,N_35154);
nand U35327 (N_35327,N_35052,N_35101);
nor U35328 (N_35328,N_35016,N_35061);
and U35329 (N_35329,N_35179,N_35099);
xor U35330 (N_35330,N_35009,N_35112);
xnor U35331 (N_35331,N_35005,N_35021);
or U35332 (N_35332,N_35059,N_35138);
and U35333 (N_35333,N_35145,N_35123);
xor U35334 (N_35334,N_35169,N_35117);
nand U35335 (N_35335,N_35180,N_35038);
or U35336 (N_35336,N_35026,N_35020);
nand U35337 (N_35337,N_35110,N_35194);
xor U35338 (N_35338,N_35140,N_35108);
nor U35339 (N_35339,N_35239,N_35141);
and U35340 (N_35340,N_35102,N_35092);
xor U35341 (N_35341,N_35079,N_35002);
nor U35342 (N_35342,N_35159,N_35087);
xor U35343 (N_35343,N_35100,N_35136);
or U35344 (N_35344,N_35090,N_35149);
xnor U35345 (N_35345,N_35247,N_35161);
nand U35346 (N_35346,N_35148,N_35091);
or U35347 (N_35347,N_35011,N_35037);
and U35348 (N_35348,N_35045,N_35158);
nand U35349 (N_35349,N_35022,N_35231);
nand U35350 (N_35350,N_35066,N_35015);
xor U35351 (N_35351,N_35132,N_35106);
or U35352 (N_35352,N_35186,N_35023);
and U35353 (N_35353,N_35165,N_35226);
or U35354 (N_35354,N_35062,N_35182);
nand U35355 (N_35355,N_35039,N_35193);
nand U35356 (N_35356,N_35003,N_35070);
nand U35357 (N_35357,N_35181,N_35055);
xnor U35358 (N_35358,N_35191,N_35152);
and U35359 (N_35359,N_35080,N_35238);
nand U35360 (N_35360,N_35196,N_35063);
nor U35361 (N_35361,N_35184,N_35188);
xor U35362 (N_35362,N_35046,N_35133);
nor U35363 (N_35363,N_35197,N_35222);
nor U35364 (N_35364,N_35235,N_35172);
and U35365 (N_35365,N_35007,N_35215);
xor U35366 (N_35366,N_35078,N_35209);
nor U35367 (N_35367,N_35155,N_35068);
nor U35368 (N_35368,N_35128,N_35135);
nand U35369 (N_35369,N_35060,N_35167);
nor U35370 (N_35370,N_35221,N_35053);
or U35371 (N_35371,N_35027,N_35202);
nor U35372 (N_35372,N_35244,N_35227);
nand U35373 (N_35373,N_35199,N_35119);
nor U35374 (N_35374,N_35121,N_35067);
and U35375 (N_35375,N_35095,N_35102);
nor U35376 (N_35376,N_35217,N_35176);
xnor U35377 (N_35377,N_35062,N_35233);
nor U35378 (N_35378,N_35152,N_35160);
nand U35379 (N_35379,N_35022,N_35198);
or U35380 (N_35380,N_35012,N_35084);
nand U35381 (N_35381,N_35170,N_35239);
or U35382 (N_35382,N_35041,N_35093);
xor U35383 (N_35383,N_35119,N_35235);
nand U35384 (N_35384,N_35109,N_35247);
nand U35385 (N_35385,N_35210,N_35225);
or U35386 (N_35386,N_35095,N_35227);
or U35387 (N_35387,N_35218,N_35014);
nor U35388 (N_35388,N_35012,N_35188);
nand U35389 (N_35389,N_35061,N_35215);
nand U35390 (N_35390,N_35190,N_35010);
or U35391 (N_35391,N_35023,N_35199);
nand U35392 (N_35392,N_35083,N_35203);
nor U35393 (N_35393,N_35013,N_35126);
nand U35394 (N_35394,N_35104,N_35137);
and U35395 (N_35395,N_35187,N_35195);
nand U35396 (N_35396,N_35083,N_35163);
and U35397 (N_35397,N_35098,N_35163);
nand U35398 (N_35398,N_35148,N_35099);
nand U35399 (N_35399,N_35038,N_35133);
or U35400 (N_35400,N_35109,N_35229);
xor U35401 (N_35401,N_35174,N_35022);
nor U35402 (N_35402,N_35214,N_35096);
xor U35403 (N_35403,N_35052,N_35152);
nand U35404 (N_35404,N_35000,N_35102);
nand U35405 (N_35405,N_35126,N_35121);
nand U35406 (N_35406,N_35081,N_35156);
nand U35407 (N_35407,N_35173,N_35169);
and U35408 (N_35408,N_35224,N_35170);
xor U35409 (N_35409,N_35150,N_35051);
and U35410 (N_35410,N_35241,N_35225);
or U35411 (N_35411,N_35158,N_35153);
or U35412 (N_35412,N_35011,N_35133);
xnor U35413 (N_35413,N_35041,N_35092);
xor U35414 (N_35414,N_35206,N_35129);
or U35415 (N_35415,N_35143,N_35082);
xnor U35416 (N_35416,N_35218,N_35171);
nor U35417 (N_35417,N_35217,N_35040);
xnor U35418 (N_35418,N_35230,N_35065);
xnor U35419 (N_35419,N_35199,N_35203);
and U35420 (N_35420,N_35104,N_35028);
or U35421 (N_35421,N_35020,N_35063);
and U35422 (N_35422,N_35206,N_35014);
or U35423 (N_35423,N_35234,N_35183);
nor U35424 (N_35424,N_35095,N_35119);
and U35425 (N_35425,N_35000,N_35129);
or U35426 (N_35426,N_35037,N_35176);
xor U35427 (N_35427,N_35097,N_35028);
nand U35428 (N_35428,N_35030,N_35111);
nor U35429 (N_35429,N_35005,N_35163);
xnor U35430 (N_35430,N_35164,N_35226);
nor U35431 (N_35431,N_35022,N_35108);
or U35432 (N_35432,N_35181,N_35112);
or U35433 (N_35433,N_35177,N_35075);
nor U35434 (N_35434,N_35004,N_35235);
and U35435 (N_35435,N_35210,N_35169);
and U35436 (N_35436,N_35009,N_35054);
nor U35437 (N_35437,N_35226,N_35104);
nor U35438 (N_35438,N_35216,N_35229);
and U35439 (N_35439,N_35127,N_35072);
xnor U35440 (N_35440,N_35146,N_35121);
xnor U35441 (N_35441,N_35136,N_35202);
nand U35442 (N_35442,N_35166,N_35136);
or U35443 (N_35443,N_35086,N_35112);
nor U35444 (N_35444,N_35247,N_35004);
nand U35445 (N_35445,N_35043,N_35104);
and U35446 (N_35446,N_35208,N_35188);
xor U35447 (N_35447,N_35003,N_35249);
xnor U35448 (N_35448,N_35168,N_35031);
and U35449 (N_35449,N_35199,N_35214);
and U35450 (N_35450,N_35014,N_35011);
nand U35451 (N_35451,N_35007,N_35148);
xnor U35452 (N_35452,N_35102,N_35063);
nor U35453 (N_35453,N_35160,N_35229);
or U35454 (N_35454,N_35117,N_35165);
or U35455 (N_35455,N_35072,N_35000);
xnor U35456 (N_35456,N_35058,N_35120);
or U35457 (N_35457,N_35070,N_35012);
or U35458 (N_35458,N_35146,N_35168);
and U35459 (N_35459,N_35135,N_35010);
and U35460 (N_35460,N_35106,N_35183);
and U35461 (N_35461,N_35090,N_35088);
nand U35462 (N_35462,N_35245,N_35229);
xnor U35463 (N_35463,N_35089,N_35083);
nor U35464 (N_35464,N_35153,N_35247);
and U35465 (N_35465,N_35065,N_35160);
or U35466 (N_35466,N_35183,N_35016);
nor U35467 (N_35467,N_35201,N_35114);
and U35468 (N_35468,N_35120,N_35176);
nor U35469 (N_35469,N_35174,N_35057);
nor U35470 (N_35470,N_35078,N_35064);
xnor U35471 (N_35471,N_35124,N_35177);
and U35472 (N_35472,N_35028,N_35021);
nand U35473 (N_35473,N_35011,N_35111);
and U35474 (N_35474,N_35213,N_35120);
nor U35475 (N_35475,N_35006,N_35046);
nor U35476 (N_35476,N_35122,N_35108);
xnor U35477 (N_35477,N_35083,N_35187);
nand U35478 (N_35478,N_35049,N_35174);
xnor U35479 (N_35479,N_35012,N_35235);
nor U35480 (N_35480,N_35210,N_35131);
and U35481 (N_35481,N_35188,N_35193);
or U35482 (N_35482,N_35233,N_35236);
xnor U35483 (N_35483,N_35153,N_35146);
nand U35484 (N_35484,N_35055,N_35143);
nor U35485 (N_35485,N_35180,N_35064);
nand U35486 (N_35486,N_35109,N_35106);
nand U35487 (N_35487,N_35021,N_35247);
nor U35488 (N_35488,N_35200,N_35058);
nand U35489 (N_35489,N_35096,N_35221);
xnor U35490 (N_35490,N_35032,N_35047);
or U35491 (N_35491,N_35230,N_35037);
nor U35492 (N_35492,N_35062,N_35137);
or U35493 (N_35493,N_35038,N_35191);
or U35494 (N_35494,N_35246,N_35187);
and U35495 (N_35495,N_35222,N_35052);
nand U35496 (N_35496,N_35188,N_35132);
or U35497 (N_35497,N_35121,N_35108);
xor U35498 (N_35498,N_35118,N_35023);
xor U35499 (N_35499,N_35218,N_35118);
nor U35500 (N_35500,N_35348,N_35353);
or U35501 (N_35501,N_35349,N_35363);
nor U35502 (N_35502,N_35366,N_35458);
and U35503 (N_35503,N_35252,N_35296);
xor U35504 (N_35504,N_35358,N_35331);
or U35505 (N_35505,N_35310,N_35283);
or U35506 (N_35506,N_35309,N_35425);
or U35507 (N_35507,N_35317,N_35372);
xor U35508 (N_35508,N_35276,N_35327);
nor U35509 (N_35509,N_35350,N_35369);
nor U35510 (N_35510,N_35382,N_35298);
nor U35511 (N_35511,N_35470,N_35436);
nor U35512 (N_35512,N_35450,N_35263);
nor U35513 (N_35513,N_35275,N_35455);
or U35514 (N_35514,N_35356,N_35258);
and U35515 (N_35515,N_35497,N_35371);
nor U35516 (N_35516,N_35361,N_35341);
nand U35517 (N_35517,N_35365,N_35380);
xor U35518 (N_35518,N_35453,N_35291);
or U35519 (N_35519,N_35277,N_35415);
nor U35520 (N_35520,N_35411,N_35253);
or U35521 (N_35521,N_35280,N_35498);
and U35522 (N_35522,N_35461,N_35305);
nand U35523 (N_35523,N_35445,N_35447);
xnor U35524 (N_35524,N_35273,N_35367);
or U35525 (N_35525,N_35322,N_35430);
xnor U35526 (N_35526,N_35306,N_35478);
and U35527 (N_35527,N_35339,N_35389);
nand U35528 (N_35528,N_35408,N_35345);
or U35529 (N_35529,N_35499,N_35267);
and U35530 (N_35530,N_35364,N_35424);
nor U35531 (N_35531,N_35311,N_35293);
xnor U35532 (N_35532,N_35264,N_35347);
and U35533 (N_35533,N_35403,N_35261);
and U35534 (N_35534,N_35385,N_35495);
or U35535 (N_35535,N_35290,N_35270);
nor U35536 (N_35536,N_35302,N_35394);
nor U35537 (N_35537,N_35409,N_35457);
and U35538 (N_35538,N_35426,N_35360);
xor U35539 (N_35539,N_35390,N_35402);
nand U35540 (N_35540,N_35352,N_35320);
nand U35541 (N_35541,N_35384,N_35404);
and U35542 (N_35542,N_35449,N_35491);
xnor U35543 (N_35543,N_35300,N_35401);
and U35544 (N_35544,N_35286,N_35472);
and U35545 (N_35545,N_35395,N_35406);
xnor U35546 (N_35546,N_35255,N_35274);
nand U35547 (N_35547,N_35278,N_35440);
xnor U35548 (N_35548,N_35388,N_35407);
or U35549 (N_35549,N_35427,N_35464);
nor U35550 (N_35550,N_35379,N_35292);
xnor U35551 (N_35551,N_35471,N_35312);
or U35552 (N_35552,N_35257,N_35370);
and U35553 (N_35553,N_35304,N_35381);
xnor U35554 (N_35554,N_35465,N_35484);
or U35555 (N_35555,N_35467,N_35431);
and U35556 (N_35556,N_35333,N_35452);
or U35557 (N_35557,N_35256,N_35251);
or U35558 (N_35558,N_35490,N_35418);
nand U35559 (N_35559,N_35446,N_35285);
nand U35560 (N_35560,N_35271,N_35260);
nand U35561 (N_35561,N_35265,N_35414);
nor U35562 (N_35562,N_35315,N_35375);
nand U35563 (N_35563,N_35479,N_35288);
or U35564 (N_35564,N_35466,N_35337);
and U35565 (N_35565,N_35272,N_35405);
xnor U35566 (N_35566,N_35284,N_35432);
or U35567 (N_35567,N_35448,N_35462);
nor U35568 (N_35568,N_35357,N_35314);
xor U35569 (N_35569,N_35468,N_35480);
and U35570 (N_35570,N_35313,N_35266);
or U35571 (N_35571,N_35494,N_35281);
or U35572 (N_35572,N_35269,N_35477);
xor U35573 (N_35573,N_35412,N_35325);
nand U35574 (N_35574,N_35299,N_35469);
or U35575 (N_35575,N_35442,N_35307);
or U35576 (N_35576,N_35328,N_35376);
and U35577 (N_35577,N_35486,N_35485);
nor U35578 (N_35578,N_35393,N_35398);
xnor U35579 (N_35579,N_35294,N_35435);
nor U35580 (N_35580,N_35493,N_35437);
xor U35581 (N_35581,N_35316,N_35454);
and U35582 (N_35582,N_35259,N_35287);
xor U35583 (N_35583,N_35487,N_35308);
and U35584 (N_35584,N_35268,N_35362);
and U35585 (N_35585,N_35397,N_35489);
or U35586 (N_35586,N_35351,N_35250);
xor U35587 (N_35587,N_35496,N_35476);
nand U35588 (N_35588,N_35387,N_35355);
nor U35589 (N_35589,N_35340,N_35262);
and U35590 (N_35590,N_35399,N_35400);
or U35591 (N_35591,N_35475,N_35459);
nor U35592 (N_35592,N_35346,N_35460);
xnor U35593 (N_35593,N_35383,N_35413);
and U35594 (N_35594,N_35392,N_35279);
xnor U35595 (N_35595,N_35428,N_35441);
and U35596 (N_35596,N_35344,N_35378);
and U35597 (N_35597,N_35330,N_35359);
or U35598 (N_35598,N_35474,N_35396);
or U35599 (N_35599,N_35368,N_35438);
and U35600 (N_35600,N_35354,N_35318);
or U35601 (N_35601,N_35323,N_35332);
nand U35602 (N_35602,N_35433,N_35295);
xor U35603 (N_35603,N_35335,N_35334);
xor U35604 (N_35604,N_35421,N_35444);
xor U35605 (N_35605,N_35336,N_35492);
xnor U35606 (N_35606,N_35301,N_35488);
xor U35607 (N_35607,N_35319,N_35342);
or U35608 (N_35608,N_35420,N_35422);
nor U35609 (N_35609,N_35373,N_35324);
or U35610 (N_35610,N_35416,N_35410);
nand U35611 (N_35611,N_35451,N_35463);
nor U35612 (N_35612,N_35386,N_35326);
and U35613 (N_35613,N_35329,N_35439);
xnor U35614 (N_35614,N_35434,N_35443);
nor U35615 (N_35615,N_35423,N_35282);
and U35616 (N_35616,N_35482,N_35289);
or U35617 (N_35617,N_35297,N_35481);
nand U35618 (N_35618,N_35391,N_35303);
xnor U35619 (N_35619,N_35254,N_35456);
or U35620 (N_35620,N_35483,N_35429);
nand U35621 (N_35621,N_35417,N_35321);
nand U35622 (N_35622,N_35374,N_35338);
and U35623 (N_35623,N_35343,N_35377);
or U35624 (N_35624,N_35473,N_35419);
nand U35625 (N_35625,N_35380,N_35362);
or U35626 (N_35626,N_35360,N_35321);
or U35627 (N_35627,N_35453,N_35332);
nand U35628 (N_35628,N_35334,N_35371);
and U35629 (N_35629,N_35276,N_35478);
nand U35630 (N_35630,N_35297,N_35383);
xnor U35631 (N_35631,N_35442,N_35491);
and U35632 (N_35632,N_35432,N_35485);
or U35633 (N_35633,N_35491,N_35330);
nor U35634 (N_35634,N_35308,N_35254);
and U35635 (N_35635,N_35406,N_35402);
or U35636 (N_35636,N_35303,N_35376);
xor U35637 (N_35637,N_35339,N_35349);
xnor U35638 (N_35638,N_35419,N_35344);
nor U35639 (N_35639,N_35347,N_35323);
and U35640 (N_35640,N_35369,N_35431);
xor U35641 (N_35641,N_35274,N_35313);
and U35642 (N_35642,N_35337,N_35305);
and U35643 (N_35643,N_35403,N_35252);
or U35644 (N_35644,N_35386,N_35355);
xnor U35645 (N_35645,N_35496,N_35402);
xnor U35646 (N_35646,N_35390,N_35427);
and U35647 (N_35647,N_35320,N_35307);
nand U35648 (N_35648,N_35357,N_35325);
nand U35649 (N_35649,N_35310,N_35368);
nor U35650 (N_35650,N_35279,N_35410);
and U35651 (N_35651,N_35272,N_35327);
nand U35652 (N_35652,N_35401,N_35295);
and U35653 (N_35653,N_35315,N_35497);
and U35654 (N_35654,N_35256,N_35336);
xnor U35655 (N_35655,N_35350,N_35407);
and U35656 (N_35656,N_35374,N_35250);
nand U35657 (N_35657,N_35251,N_35291);
xor U35658 (N_35658,N_35486,N_35324);
nor U35659 (N_35659,N_35471,N_35324);
nor U35660 (N_35660,N_35416,N_35288);
and U35661 (N_35661,N_35439,N_35491);
or U35662 (N_35662,N_35458,N_35416);
xor U35663 (N_35663,N_35289,N_35366);
xor U35664 (N_35664,N_35454,N_35337);
nand U35665 (N_35665,N_35389,N_35366);
xnor U35666 (N_35666,N_35373,N_35480);
nor U35667 (N_35667,N_35369,N_35467);
nand U35668 (N_35668,N_35426,N_35345);
nor U35669 (N_35669,N_35387,N_35473);
and U35670 (N_35670,N_35343,N_35253);
and U35671 (N_35671,N_35498,N_35364);
and U35672 (N_35672,N_35323,N_35327);
and U35673 (N_35673,N_35255,N_35472);
xnor U35674 (N_35674,N_35365,N_35320);
xnor U35675 (N_35675,N_35379,N_35484);
nor U35676 (N_35676,N_35327,N_35291);
nor U35677 (N_35677,N_35312,N_35369);
xor U35678 (N_35678,N_35487,N_35261);
nand U35679 (N_35679,N_35321,N_35438);
nand U35680 (N_35680,N_35468,N_35279);
nor U35681 (N_35681,N_35330,N_35320);
xor U35682 (N_35682,N_35448,N_35449);
nor U35683 (N_35683,N_35479,N_35285);
xnor U35684 (N_35684,N_35458,N_35292);
or U35685 (N_35685,N_35477,N_35424);
nand U35686 (N_35686,N_35421,N_35332);
nor U35687 (N_35687,N_35410,N_35266);
xnor U35688 (N_35688,N_35386,N_35476);
nor U35689 (N_35689,N_35325,N_35305);
or U35690 (N_35690,N_35418,N_35337);
or U35691 (N_35691,N_35368,N_35329);
nand U35692 (N_35692,N_35374,N_35448);
xor U35693 (N_35693,N_35262,N_35254);
or U35694 (N_35694,N_35374,N_35430);
or U35695 (N_35695,N_35259,N_35285);
or U35696 (N_35696,N_35328,N_35295);
nand U35697 (N_35697,N_35286,N_35363);
nand U35698 (N_35698,N_35269,N_35316);
xor U35699 (N_35699,N_35268,N_35303);
xnor U35700 (N_35700,N_35320,N_35261);
nor U35701 (N_35701,N_35412,N_35486);
or U35702 (N_35702,N_35343,N_35497);
nor U35703 (N_35703,N_35266,N_35293);
nor U35704 (N_35704,N_35311,N_35414);
and U35705 (N_35705,N_35320,N_35303);
nor U35706 (N_35706,N_35255,N_35453);
and U35707 (N_35707,N_35396,N_35263);
and U35708 (N_35708,N_35305,N_35309);
and U35709 (N_35709,N_35484,N_35346);
and U35710 (N_35710,N_35405,N_35469);
and U35711 (N_35711,N_35330,N_35388);
and U35712 (N_35712,N_35311,N_35329);
nor U35713 (N_35713,N_35290,N_35363);
xor U35714 (N_35714,N_35269,N_35294);
nand U35715 (N_35715,N_35487,N_35265);
nand U35716 (N_35716,N_35385,N_35322);
nand U35717 (N_35717,N_35443,N_35295);
nand U35718 (N_35718,N_35291,N_35482);
xnor U35719 (N_35719,N_35479,N_35400);
nand U35720 (N_35720,N_35331,N_35430);
nand U35721 (N_35721,N_35420,N_35297);
nand U35722 (N_35722,N_35455,N_35324);
nand U35723 (N_35723,N_35422,N_35340);
nand U35724 (N_35724,N_35497,N_35265);
or U35725 (N_35725,N_35482,N_35334);
nor U35726 (N_35726,N_35373,N_35475);
nor U35727 (N_35727,N_35343,N_35470);
and U35728 (N_35728,N_35309,N_35432);
and U35729 (N_35729,N_35312,N_35496);
and U35730 (N_35730,N_35356,N_35335);
xor U35731 (N_35731,N_35435,N_35394);
and U35732 (N_35732,N_35297,N_35462);
nor U35733 (N_35733,N_35286,N_35496);
and U35734 (N_35734,N_35474,N_35408);
nand U35735 (N_35735,N_35387,N_35281);
xor U35736 (N_35736,N_35305,N_35329);
nor U35737 (N_35737,N_35432,N_35365);
nor U35738 (N_35738,N_35496,N_35381);
nand U35739 (N_35739,N_35250,N_35299);
nand U35740 (N_35740,N_35367,N_35499);
or U35741 (N_35741,N_35315,N_35453);
nor U35742 (N_35742,N_35287,N_35474);
nor U35743 (N_35743,N_35348,N_35433);
and U35744 (N_35744,N_35262,N_35315);
nand U35745 (N_35745,N_35273,N_35378);
nand U35746 (N_35746,N_35430,N_35401);
xnor U35747 (N_35747,N_35490,N_35327);
xnor U35748 (N_35748,N_35252,N_35372);
nor U35749 (N_35749,N_35483,N_35439);
or U35750 (N_35750,N_35623,N_35603);
nor U35751 (N_35751,N_35701,N_35551);
xor U35752 (N_35752,N_35631,N_35709);
nor U35753 (N_35753,N_35677,N_35669);
or U35754 (N_35754,N_35512,N_35724);
and U35755 (N_35755,N_35507,N_35736);
or U35756 (N_35756,N_35745,N_35649);
and U35757 (N_35757,N_35561,N_35719);
or U35758 (N_35758,N_35647,N_35521);
nand U35759 (N_35759,N_35590,N_35548);
or U35760 (N_35760,N_35661,N_35567);
and U35761 (N_35761,N_35565,N_35515);
nand U35762 (N_35762,N_35554,N_35558);
xor U35763 (N_35763,N_35697,N_35673);
nor U35764 (N_35764,N_35511,N_35714);
and U35765 (N_35765,N_35625,N_35648);
and U35766 (N_35766,N_35587,N_35718);
and U35767 (N_35767,N_35730,N_35549);
nand U35768 (N_35768,N_35675,N_35642);
nand U35769 (N_35769,N_35666,N_35566);
xor U35770 (N_35770,N_35505,N_35692);
nor U35771 (N_35771,N_35598,N_35615);
xnor U35772 (N_35772,N_35633,N_35576);
or U35773 (N_35773,N_35588,N_35572);
or U35774 (N_35774,N_35733,N_35609);
or U35775 (N_35775,N_35728,N_35513);
or U35776 (N_35776,N_35628,N_35651);
nor U35777 (N_35777,N_35681,N_35611);
nor U35778 (N_35778,N_35556,N_35531);
or U35779 (N_35779,N_35610,N_35746);
or U35780 (N_35780,N_35735,N_35620);
xor U35781 (N_35781,N_35510,N_35700);
xor U35782 (N_35782,N_35659,N_35656);
or U35783 (N_35783,N_35694,N_35635);
nor U35784 (N_35784,N_35687,N_35644);
or U35785 (N_35785,N_35641,N_35538);
or U35786 (N_35786,N_35508,N_35645);
xor U35787 (N_35787,N_35653,N_35529);
xnor U35788 (N_35788,N_35546,N_35643);
nand U35789 (N_35789,N_35721,N_35537);
and U35790 (N_35790,N_35679,N_35705);
and U35791 (N_35791,N_35711,N_35654);
and U35792 (N_35792,N_35589,N_35715);
nand U35793 (N_35793,N_35504,N_35562);
nor U35794 (N_35794,N_35703,N_35626);
nor U35795 (N_35795,N_35747,N_35748);
nand U35796 (N_35796,N_35682,N_35544);
nor U35797 (N_35797,N_35522,N_35665);
nand U35798 (N_35798,N_35591,N_35506);
nand U35799 (N_35799,N_35744,N_35691);
xnor U35800 (N_35800,N_35612,N_35698);
and U35801 (N_35801,N_35704,N_35624);
and U35802 (N_35802,N_35596,N_35541);
xor U35803 (N_35803,N_35637,N_35618);
nand U35804 (N_35804,N_35640,N_35743);
nand U35805 (N_35805,N_35706,N_35533);
nor U35806 (N_35806,N_35520,N_35502);
xor U35807 (N_35807,N_35571,N_35543);
nand U35808 (N_35808,N_35660,N_35713);
or U35809 (N_35809,N_35555,N_35634);
or U35810 (N_35810,N_35740,N_35619);
nand U35811 (N_35811,N_35726,N_35563);
nor U35812 (N_35812,N_35578,N_35509);
nor U35813 (N_35813,N_35530,N_35501);
nand U35814 (N_35814,N_35532,N_35630);
nor U35815 (N_35815,N_35584,N_35517);
or U35816 (N_35816,N_35586,N_35597);
or U35817 (N_35817,N_35707,N_35622);
or U35818 (N_35818,N_35749,N_35650);
and U35819 (N_35819,N_35632,N_35668);
nor U35820 (N_35820,N_35695,N_35674);
nor U35821 (N_35821,N_35734,N_35594);
nor U35822 (N_35822,N_35607,N_35540);
nand U35823 (N_35823,N_35592,N_35712);
nor U35824 (N_35824,N_35727,N_35720);
or U35825 (N_35825,N_35500,N_35729);
nand U35826 (N_35826,N_35608,N_35693);
nand U35827 (N_35827,N_35652,N_35577);
and U35828 (N_35828,N_35518,N_35685);
nand U35829 (N_35829,N_35629,N_35606);
xnor U35830 (N_35830,N_35680,N_35545);
nand U35831 (N_35831,N_35559,N_35684);
and U35832 (N_35832,N_35613,N_35683);
nand U35833 (N_35833,N_35573,N_35536);
nor U35834 (N_35834,N_35528,N_35671);
and U35835 (N_35835,N_35580,N_35604);
xor U35836 (N_35836,N_35568,N_35614);
and U35837 (N_35837,N_35579,N_35569);
nor U35838 (N_35838,N_35670,N_35737);
nor U35839 (N_35839,N_35723,N_35638);
nand U35840 (N_35840,N_35575,N_35672);
nand U35841 (N_35841,N_35526,N_35710);
xnor U35842 (N_35842,N_35539,N_35678);
or U35843 (N_35843,N_35655,N_35664);
xnor U35844 (N_35844,N_35617,N_35732);
nand U35845 (N_35845,N_35689,N_35658);
nand U35846 (N_35846,N_35534,N_35662);
and U35847 (N_35847,N_35605,N_35731);
xor U35848 (N_35848,N_35741,N_35593);
nand U35849 (N_35849,N_35702,N_35686);
nor U35850 (N_35850,N_35525,N_35742);
or U35851 (N_35851,N_35542,N_35583);
nor U35852 (N_35852,N_35547,N_35519);
and U35853 (N_35853,N_35722,N_35636);
nand U35854 (N_35854,N_35600,N_35535);
xor U35855 (N_35855,N_35708,N_35725);
xnor U35856 (N_35856,N_35516,N_35581);
xnor U35857 (N_35857,N_35688,N_35550);
or U35858 (N_35858,N_35599,N_35716);
or U35859 (N_35859,N_35663,N_35514);
and U35860 (N_35860,N_35739,N_35595);
nand U35861 (N_35861,N_35690,N_35657);
and U35862 (N_35862,N_35627,N_35602);
nor U35863 (N_35863,N_35553,N_35527);
or U35864 (N_35864,N_35574,N_35523);
nand U35865 (N_35865,N_35557,N_35738);
and U35866 (N_35866,N_35639,N_35552);
nand U35867 (N_35867,N_35570,N_35564);
nor U35868 (N_35868,N_35503,N_35621);
xor U35869 (N_35869,N_35524,N_35560);
or U35870 (N_35870,N_35582,N_35699);
or U35871 (N_35871,N_35646,N_35585);
and U35872 (N_35872,N_35601,N_35676);
or U35873 (N_35873,N_35717,N_35667);
xor U35874 (N_35874,N_35696,N_35616);
xor U35875 (N_35875,N_35625,N_35695);
nand U35876 (N_35876,N_35577,N_35683);
nand U35877 (N_35877,N_35528,N_35651);
nand U35878 (N_35878,N_35718,N_35555);
nor U35879 (N_35879,N_35734,N_35563);
xor U35880 (N_35880,N_35698,N_35579);
xor U35881 (N_35881,N_35546,N_35734);
and U35882 (N_35882,N_35650,N_35626);
or U35883 (N_35883,N_35504,N_35580);
or U35884 (N_35884,N_35688,N_35734);
nor U35885 (N_35885,N_35703,N_35618);
nor U35886 (N_35886,N_35516,N_35673);
or U35887 (N_35887,N_35663,N_35632);
xor U35888 (N_35888,N_35729,N_35579);
nand U35889 (N_35889,N_35737,N_35649);
and U35890 (N_35890,N_35580,N_35705);
nand U35891 (N_35891,N_35622,N_35727);
and U35892 (N_35892,N_35516,N_35579);
and U35893 (N_35893,N_35600,N_35681);
xor U35894 (N_35894,N_35677,N_35541);
and U35895 (N_35895,N_35500,N_35723);
nand U35896 (N_35896,N_35720,N_35565);
or U35897 (N_35897,N_35581,N_35603);
nand U35898 (N_35898,N_35741,N_35644);
nor U35899 (N_35899,N_35722,N_35681);
or U35900 (N_35900,N_35613,N_35580);
and U35901 (N_35901,N_35516,N_35546);
nand U35902 (N_35902,N_35743,N_35655);
nor U35903 (N_35903,N_35543,N_35590);
nor U35904 (N_35904,N_35697,N_35615);
or U35905 (N_35905,N_35620,N_35520);
nor U35906 (N_35906,N_35683,N_35518);
or U35907 (N_35907,N_35725,N_35614);
nand U35908 (N_35908,N_35646,N_35709);
nor U35909 (N_35909,N_35716,N_35690);
nand U35910 (N_35910,N_35547,N_35622);
nor U35911 (N_35911,N_35564,N_35522);
nor U35912 (N_35912,N_35661,N_35629);
xor U35913 (N_35913,N_35702,N_35512);
or U35914 (N_35914,N_35649,N_35522);
and U35915 (N_35915,N_35729,N_35690);
xor U35916 (N_35916,N_35629,N_35512);
nor U35917 (N_35917,N_35622,N_35665);
nand U35918 (N_35918,N_35735,N_35714);
nand U35919 (N_35919,N_35694,N_35608);
or U35920 (N_35920,N_35725,N_35742);
or U35921 (N_35921,N_35527,N_35714);
and U35922 (N_35922,N_35584,N_35736);
or U35923 (N_35923,N_35745,N_35533);
or U35924 (N_35924,N_35721,N_35615);
or U35925 (N_35925,N_35532,N_35733);
xnor U35926 (N_35926,N_35547,N_35692);
and U35927 (N_35927,N_35589,N_35584);
or U35928 (N_35928,N_35626,N_35744);
and U35929 (N_35929,N_35611,N_35577);
xnor U35930 (N_35930,N_35667,N_35624);
xor U35931 (N_35931,N_35516,N_35549);
and U35932 (N_35932,N_35694,N_35628);
nand U35933 (N_35933,N_35679,N_35598);
or U35934 (N_35934,N_35733,N_35647);
xor U35935 (N_35935,N_35524,N_35599);
or U35936 (N_35936,N_35711,N_35576);
nand U35937 (N_35937,N_35647,N_35617);
nor U35938 (N_35938,N_35624,N_35607);
nand U35939 (N_35939,N_35560,N_35671);
xnor U35940 (N_35940,N_35609,N_35544);
nand U35941 (N_35941,N_35706,N_35539);
and U35942 (N_35942,N_35624,N_35747);
nand U35943 (N_35943,N_35527,N_35660);
nor U35944 (N_35944,N_35718,N_35613);
or U35945 (N_35945,N_35749,N_35538);
nand U35946 (N_35946,N_35728,N_35726);
and U35947 (N_35947,N_35592,N_35743);
and U35948 (N_35948,N_35566,N_35658);
xor U35949 (N_35949,N_35516,N_35687);
xor U35950 (N_35950,N_35519,N_35655);
xnor U35951 (N_35951,N_35557,N_35533);
xnor U35952 (N_35952,N_35572,N_35644);
xor U35953 (N_35953,N_35675,N_35654);
or U35954 (N_35954,N_35749,N_35632);
or U35955 (N_35955,N_35723,N_35549);
or U35956 (N_35956,N_35675,N_35619);
or U35957 (N_35957,N_35576,N_35657);
nand U35958 (N_35958,N_35733,N_35690);
and U35959 (N_35959,N_35538,N_35732);
and U35960 (N_35960,N_35543,N_35540);
and U35961 (N_35961,N_35585,N_35676);
or U35962 (N_35962,N_35503,N_35566);
and U35963 (N_35963,N_35663,N_35558);
and U35964 (N_35964,N_35667,N_35634);
nor U35965 (N_35965,N_35730,N_35612);
nor U35966 (N_35966,N_35622,N_35605);
and U35967 (N_35967,N_35558,N_35685);
nand U35968 (N_35968,N_35504,N_35551);
xor U35969 (N_35969,N_35557,N_35563);
nor U35970 (N_35970,N_35668,N_35670);
xnor U35971 (N_35971,N_35588,N_35726);
and U35972 (N_35972,N_35602,N_35634);
and U35973 (N_35973,N_35597,N_35592);
xnor U35974 (N_35974,N_35540,N_35739);
nand U35975 (N_35975,N_35622,N_35692);
and U35976 (N_35976,N_35526,N_35516);
nand U35977 (N_35977,N_35675,N_35551);
nor U35978 (N_35978,N_35678,N_35629);
nor U35979 (N_35979,N_35749,N_35734);
nor U35980 (N_35980,N_35703,N_35690);
nand U35981 (N_35981,N_35715,N_35704);
and U35982 (N_35982,N_35574,N_35576);
or U35983 (N_35983,N_35611,N_35695);
nor U35984 (N_35984,N_35748,N_35536);
xnor U35985 (N_35985,N_35726,N_35574);
nand U35986 (N_35986,N_35553,N_35592);
xor U35987 (N_35987,N_35601,N_35619);
and U35988 (N_35988,N_35573,N_35575);
or U35989 (N_35989,N_35633,N_35652);
nor U35990 (N_35990,N_35618,N_35660);
nor U35991 (N_35991,N_35682,N_35602);
xnor U35992 (N_35992,N_35517,N_35501);
nor U35993 (N_35993,N_35654,N_35651);
and U35994 (N_35994,N_35547,N_35746);
nand U35995 (N_35995,N_35744,N_35720);
or U35996 (N_35996,N_35599,N_35637);
or U35997 (N_35997,N_35566,N_35659);
or U35998 (N_35998,N_35694,N_35682);
and U35999 (N_35999,N_35558,N_35591);
xor U36000 (N_36000,N_35921,N_35981);
or U36001 (N_36001,N_35914,N_35771);
and U36002 (N_36002,N_35823,N_35927);
nand U36003 (N_36003,N_35756,N_35901);
xnor U36004 (N_36004,N_35807,N_35933);
and U36005 (N_36005,N_35791,N_35881);
or U36006 (N_36006,N_35802,N_35822);
and U36007 (N_36007,N_35839,N_35836);
xnor U36008 (N_36008,N_35794,N_35997);
nor U36009 (N_36009,N_35887,N_35980);
or U36010 (N_36010,N_35984,N_35751);
and U36011 (N_36011,N_35967,N_35957);
or U36012 (N_36012,N_35994,N_35853);
nor U36013 (N_36013,N_35851,N_35828);
or U36014 (N_36014,N_35973,N_35963);
xnor U36015 (N_36015,N_35975,N_35867);
or U36016 (N_36016,N_35987,N_35805);
or U36017 (N_36017,N_35868,N_35934);
or U36018 (N_36018,N_35784,N_35939);
nand U36019 (N_36019,N_35972,N_35892);
xnor U36020 (N_36020,N_35782,N_35950);
nor U36021 (N_36021,N_35846,N_35837);
or U36022 (N_36022,N_35775,N_35960);
nor U36023 (N_36023,N_35962,N_35768);
nor U36024 (N_36024,N_35806,N_35835);
nor U36025 (N_36025,N_35863,N_35774);
nor U36026 (N_36026,N_35880,N_35964);
or U36027 (N_36027,N_35793,N_35841);
and U36028 (N_36028,N_35941,N_35917);
or U36029 (N_36029,N_35761,N_35808);
and U36030 (N_36030,N_35790,N_35924);
or U36031 (N_36031,N_35818,N_35845);
and U36032 (N_36032,N_35883,N_35843);
nand U36033 (N_36033,N_35780,N_35826);
and U36034 (N_36034,N_35936,N_35885);
or U36035 (N_36035,N_35849,N_35876);
nand U36036 (N_36036,N_35942,N_35872);
or U36037 (N_36037,N_35855,N_35988);
xnor U36038 (N_36038,N_35777,N_35852);
nor U36039 (N_36039,N_35860,N_35817);
xor U36040 (N_36040,N_35926,N_35765);
nor U36041 (N_36041,N_35955,N_35970);
nand U36042 (N_36042,N_35752,N_35976);
and U36043 (N_36043,N_35923,N_35781);
or U36044 (N_36044,N_35909,N_35848);
nand U36045 (N_36045,N_35918,N_35797);
nand U36046 (N_36046,N_35974,N_35778);
and U36047 (N_36047,N_35786,N_35940);
xor U36048 (N_36048,N_35903,N_35796);
or U36049 (N_36049,N_35882,N_35965);
nand U36050 (N_36050,N_35992,N_35819);
and U36051 (N_36051,N_35945,N_35913);
nand U36052 (N_36052,N_35821,N_35840);
and U36053 (N_36053,N_35888,N_35831);
or U36054 (N_36054,N_35857,N_35866);
and U36055 (N_36055,N_35847,N_35800);
or U36056 (N_36056,N_35982,N_35958);
nor U36057 (N_36057,N_35772,N_35906);
nand U36058 (N_36058,N_35759,N_35953);
and U36059 (N_36059,N_35971,N_35985);
or U36060 (N_36060,N_35877,N_35889);
or U36061 (N_36061,N_35993,N_35760);
and U36062 (N_36062,N_35838,N_35787);
nand U36063 (N_36063,N_35938,N_35832);
or U36064 (N_36064,N_35755,N_35912);
or U36065 (N_36065,N_35754,N_35978);
and U36066 (N_36066,N_35795,N_35825);
or U36067 (N_36067,N_35816,N_35799);
or U36068 (N_36068,N_35865,N_35925);
xnor U36069 (N_36069,N_35815,N_35900);
nand U36070 (N_36070,N_35859,N_35944);
nor U36071 (N_36071,N_35803,N_35928);
and U36072 (N_36072,N_35767,N_35873);
nand U36073 (N_36073,N_35813,N_35996);
xor U36074 (N_36074,N_35966,N_35779);
nand U36075 (N_36075,N_35809,N_35911);
nand U36076 (N_36076,N_35935,N_35764);
nand U36077 (N_36077,N_35879,N_35930);
nor U36078 (N_36078,N_35897,N_35789);
and U36079 (N_36079,N_35951,N_35814);
and U36080 (N_36080,N_35915,N_35827);
nand U36081 (N_36081,N_35758,N_35753);
nand U36082 (N_36082,N_35949,N_35968);
xnor U36083 (N_36083,N_35969,N_35861);
and U36084 (N_36084,N_35884,N_35983);
nand U36085 (N_36085,N_35820,N_35959);
and U36086 (N_36086,N_35919,N_35932);
and U36087 (N_36087,N_35812,N_35948);
nand U36088 (N_36088,N_35869,N_35990);
and U36089 (N_36089,N_35844,N_35995);
nor U36090 (N_36090,N_35874,N_35895);
and U36091 (N_36091,N_35770,N_35998);
nand U36092 (N_36092,N_35829,N_35878);
nor U36093 (N_36093,N_35893,N_35946);
xnor U36094 (N_36094,N_35858,N_35757);
and U36095 (N_36095,N_35811,N_35856);
and U36096 (N_36096,N_35750,N_35788);
nor U36097 (N_36097,N_35776,N_35999);
nand U36098 (N_36098,N_35952,N_35891);
and U36099 (N_36099,N_35850,N_35908);
nand U36100 (N_36100,N_35763,N_35766);
nor U36101 (N_36101,N_35896,N_35824);
nor U36102 (N_36102,N_35842,N_35870);
and U36103 (N_36103,N_35785,N_35986);
xnor U36104 (N_36104,N_35792,N_35905);
xor U36105 (N_36105,N_35894,N_35890);
or U36106 (N_36106,N_35991,N_35989);
nand U36107 (N_36107,N_35875,N_35956);
xnor U36108 (N_36108,N_35798,N_35910);
or U36109 (N_36109,N_35830,N_35834);
nand U36110 (N_36110,N_35916,N_35907);
nand U36111 (N_36111,N_35961,N_35954);
nor U36112 (N_36112,N_35801,N_35854);
or U36113 (N_36113,N_35810,N_35920);
or U36114 (N_36114,N_35902,N_35947);
and U36115 (N_36115,N_35864,N_35769);
nand U36116 (N_36116,N_35862,N_35886);
or U36117 (N_36117,N_35783,N_35871);
nand U36118 (N_36118,N_35899,N_35804);
xor U36119 (N_36119,N_35977,N_35904);
nor U36120 (N_36120,N_35943,N_35773);
and U36121 (N_36121,N_35833,N_35762);
xnor U36122 (N_36122,N_35931,N_35929);
and U36123 (N_36123,N_35937,N_35922);
nor U36124 (N_36124,N_35979,N_35898);
nor U36125 (N_36125,N_35834,N_35820);
and U36126 (N_36126,N_35979,N_35952);
xor U36127 (N_36127,N_35808,N_35813);
nor U36128 (N_36128,N_35896,N_35873);
nor U36129 (N_36129,N_35933,N_35819);
or U36130 (N_36130,N_35956,N_35877);
and U36131 (N_36131,N_35864,N_35819);
or U36132 (N_36132,N_35933,N_35974);
nand U36133 (N_36133,N_35813,N_35964);
nor U36134 (N_36134,N_35895,N_35793);
nor U36135 (N_36135,N_35891,N_35922);
nor U36136 (N_36136,N_35833,N_35975);
nor U36137 (N_36137,N_35944,N_35881);
xnor U36138 (N_36138,N_35924,N_35884);
or U36139 (N_36139,N_35968,N_35915);
and U36140 (N_36140,N_35995,N_35902);
nand U36141 (N_36141,N_35777,N_35912);
xor U36142 (N_36142,N_35812,N_35915);
or U36143 (N_36143,N_35875,N_35816);
and U36144 (N_36144,N_35898,N_35921);
nand U36145 (N_36145,N_35869,N_35880);
xor U36146 (N_36146,N_35985,N_35858);
or U36147 (N_36147,N_35859,N_35917);
nand U36148 (N_36148,N_35908,N_35894);
nor U36149 (N_36149,N_35837,N_35999);
and U36150 (N_36150,N_35870,N_35971);
xnor U36151 (N_36151,N_35778,N_35787);
xnor U36152 (N_36152,N_35751,N_35811);
or U36153 (N_36153,N_35843,N_35980);
and U36154 (N_36154,N_35952,N_35828);
and U36155 (N_36155,N_35952,N_35837);
or U36156 (N_36156,N_35766,N_35930);
nand U36157 (N_36157,N_35754,N_35788);
nand U36158 (N_36158,N_35751,N_35750);
and U36159 (N_36159,N_35829,N_35977);
xor U36160 (N_36160,N_35991,N_35882);
or U36161 (N_36161,N_35966,N_35875);
and U36162 (N_36162,N_35910,N_35773);
nor U36163 (N_36163,N_35935,N_35807);
nand U36164 (N_36164,N_35859,N_35985);
xor U36165 (N_36165,N_35760,N_35997);
nand U36166 (N_36166,N_35892,N_35968);
or U36167 (N_36167,N_35944,N_35817);
nor U36168 (N_36168,N_35868,N_35975);
or U36169 (N_36169,N_35750,N_35916);
nand U36170 (N_36170,N_35867,N_35820);
nand U36171 (N_36171,N_35852,N_35896);
xor U36172 (N_36172,N_35863,N_35891);
and U36173 (N_36173,N_35848,N_35904);
nor U36174 (N_36174,N_35851,N_35771);
xnor U36175 (N_36175,N_35762,N_35956);
xnor U36176 (N_36176,N_35836,N_35765);
nor U36177 (N_36177,N_35841,N_35811);
nor U36178 (N_36178,N_35894,N_35887);
nor U36179 (N_36179,N_35754,N_35917);
xor U36180 (N_36180,N_35988,N_35930);
xor U36181 (N_36181,N_35867,N_35753);
or U36182 (N_36182,N_35755,N_35770);
nor U36183 (N_36183,N_35862,N_35929);
nand U36184 (N_36184,N_35990,N_35799);
nor U36185 (N_36185,N_35779,N_35934);
xor U36186 (N_36186,N_35866,N_35783);
and U36187 (N_36187,N_35924,N_35839);
and U36188 (N_36188,N_35907,N_35812);
or U36189 (N_36189,N_35777,N_35856);
xnor U36190 (N_36190,N_35923,N_35884);
nand U36191 (N_36191,N_35961,N_35960);
nor U36192 (N_36192,N_35923,N_35937);
nor U36193 (N_36193,N_35793,N_35901);
nor U36194 (N_36194,N_35761,N_35840);
xnor U36195 (N_36195,N_35752,N_35998);
or U36196 (N_36196,N_35920,N_35949);
and U36197 (N_36197,N_35929,N_35944);
nand U36198 (N_36198,N_35864,N_35797);
and U36199 (N_36199,N_35780,N_35952);
xnor U36200 (N_36200,N_35884,N_35980);
xor U36201 (N_36201,N_35767,N_35816);
or U36202 (N_36202,N_35766,N_35875);
nor U36203 (N_36203,N_35785,N_35995);
or U36204 (N_36204,N_35999,N_35757);
xor U36205 (N_36205,N_35752,N_35977);
or U36206 (N_36206,N_35797,N_35863);
nor U36207 (N_36207,N_35801,N_35997);
or U36208 (N_36208,N_35821,N_35936);
xnor U36209 (N_36209,N_35884,N_35928);
nand U36210 (N_36210,N_35986,N_35853);
xor U36211 (N_36211,N_35892,N_35836);
nand U36212 (N_36212,N_35809,N_35990);
or U36213 (N_36213,N_35890,N_35958);
nor U36214 (N_36214,N_35908,N_35829);
xor U36215 (N_36215,N_35859,N_35897);
nand U36216 (N_36216,N_35960,N_35975);
and U36217 (N_36217,N_35768,N_35797);
xnor U36218 (N_36218,N_35790,N_35943);
xnor U36219 (N_36219,N_35853,N_35898);
nor U36220 (N_36220,N_35789,N_35985);
and U36221 (N_36221,N_35865,N_35884);
nor U36222 (N_36222,N_35976,N_35990);
xor U36223 (N_36223,N_35818,N_35914);
nor U36224 (N_36224,N_35800,N_35940);
xnor U36225 (N_36225,N_35901,N_35855);
nor U36226 (N_36226,N_35933,N_35751);
xor U36227 (N_36227,N_35881,N_35907);
xor U36228 (N_36228,N_35926,N_35799);
or U36229 (N_36229,N_35949,N_35753);
or U36230 (N_36230,N_35860,N_35982);
nand U36231 (N_36231,N_35934,N_35840);
nand U36232 (N_36232,N_35949,N_35983);
and U36233 (N_36233,N_35872,N_35821);
xor U36234 (N_36234,N_35895,N_35920);
and U36235 (N_36235,N_35771,N_35896);
nand U36236 (N_36236,N_35995,N_35885);
or U36237 (N_36237,N_35823,N_35863);
or U36238 (N_36238,N_35926,N_35885);
or U36239 (N_36239,N_35816,N_35963);
and U36240 (N_36240,N_35758,N_35848);
nor U36241 (N_36241,N_35928,N_35787);
or U36242 (N_36242,N_35927,N_35974);
xnor U36243 (N_36243,N_35849,N_35813);
nand U36244 (N_36244,N_35965,N_35847);
nor U36245 (N_36245,N_35851,N_35850);
nor U36246 (N_36246,N_35893,N_35921);
or U36247 (N_36247,N_35830,N_35885);
and U36248 (N_36248,N_35935,N_35781);
or U36249 (N_36249,N_35824,N_35847);
nand U36250 (N_36250,N_36232,N_36113);
nor U36251 (N_36251,N_36096,N_36198);
nor U36252 (N_36252,N_36147,N_36033);
nor U36253 (N_36253,N_36123,N_36202);
or U36254 (N_36254,N_36124,N_36017);
and U36255 (N_36255,N_36084,N_36183);
or U36256 (N_36256,N_36225,N_36083);
or U36257 (N_36257,N_36106,N_36093);
and U36258 (N_36258,N_36164,N_36039);
xnor U36259 (N_36259,N_36068,N_36026);
nand U36260 (N_36260,N_36206,N_36161);
xnor U36261 (N_36261,N_36234,N_36203);
nand U36262 (N_36262,N_36201,N_36244);
nor U36263 (N_36263,N_36142,N_36072);
nor U36264 (N_36264,N_36182,N_36020);
nand U36265 (N_36265,N_36197,N_36023);
xnor U36266 (N_36266,N_36220,N_36078);
xnor U36267 (N_36267,N_36181,N_36191);
xor U36268 (N_36268,N_36008,N_36235);
nand U36269 (N_36269,N_36100,N_36159);
xnor U36270 (N_36270,N_36111,N_36042);
nor U36271 (N_36271,N_36028,N_36097);
nand U36272 (N_36272,N_36036,N_36185);
and U36273 (N_36273,N_36057,N_36230);
nor U36274 (N_36274,N_36178,N_36085);
xnor U36275 (N_36275,N_36059,N_36027);
or U36276 (N_36276,N_36199,N_36200);
nand U36277 (N_36277,N_36153,N_36210);
or U36278 (N_36278,N_36025,N_36095);
or U36279 (N_36279,N_36247,N_36233);
nand U36280 (N_36280,N_36044,N_36052);
or U36281 (N_36281,N_36174,N_36176);
or U36282 (N_36282,N_36166,N_36104);
or U36283 (N_36283,N_36120,N_36040);
nand U36284 (N_36284,N_36238,N_36169);
and U36285 (N_36285,N_36126,N_36221);
and U36286 (N_36286,N_36156,N_36217);
and U36287 (N_36287,N_36158,N_36237);
nand U36288 (N_36288,N_36146,N_36196);
xnor U36289 (N_36289,N_36131,N_36157);
nand U36290 (N_36290,N_36140,N_36240);
or U36291 (N_36291,N_36089,N_36228);
or U36292 (N_36292,N_36035,N_36053);
nor U36293 (N_36293,N_36048,N_36115);
xnor U36294 (N_36294,N_36010,N_36070);
nor U36295 (N_36295,N_36179,N_36121);
and U36296 (N_36296,N_36170,N_36009);
or U36297 (N_36297,N_36007,N_36037);
or U36298 (N_36298,N_36049,N_36031);
nand U36299 (N_36299,N_36133,N_36110);
or U36300 (N_36300,N_36060,N_36224);
xnor U36301 (N_36301,N_36167,N_36154);
nor U36302 (N_36302,N_36137,N_36127);
and U36303 (N_36303,N_36103,N_36248);
nor U36304 (N_36304,N_36163,N_36148);
nor U36305 (N_36305,N_36223,N_36227);
xnor U36306 (N_36306,N_36135,N_36001);
nor U36307 (N_36307,N_36077,N_36193);
nand U36308 (N_36308,N_36136,N_36081);
nand U36309 (N_36309,N_36215,N_36139);
nand U36310 (N_36310,N_36018,N_36175);
nor U36311 (N_36311,N_36245,N_36216);
nor U36312 (N_36312,N_36029,N_36003);
or U36313 (N_36313,N_36032,N_36071);
nand U36314 (N_36314,N_36222,N_36122);
nor U36315 (N_36315,N_36046,N_36082);
or U36316 (N_36316,N_36192,N_36118);
or U36317 (N_36317,N_36030,N_36114);
nand U36318 (N_36318,N_36092,N_36058);
xor U36319 (N_36319,N_36173,N_36090);
or U36320 (N_36320,N_36226,N_36172);
or U36321 (N_36321,N_36079,N_36144);
nand U36322 (N_36322,N_36208,N_36205);
and U36323 (N_36323,N_36075,N_36239);
nor U36324 (N_36324,N_36125,N_36209);
nor U36325 (N_36325,N_36108,N_36102);
nor U36326 (N_36326,N_36012,N_36069);
and U36327 (N_36327,N_36129,N_36087);
xor U36328 (N_36328,N_36231,N_36246);
nor U36329 (N_36329,N_36051,N_36074);
or U36330 (N_36330,N_36004,N_36213);
and U36331 (N_36331,N_36091,N_36076);
nor U36332 (N_36332,N_36195,N_36150);
or U36333 (N_36333,N_36013,N_36015);
nand U36334 (N_36334,N_36065,N_36016);
nor U36335 (N_36335,N_36034,N_36101);
and U36336 (N_36336,N_36130,N_36080);
and U36337 (N_36337,N_36184,N_36038);
nor U36338 (N_36338,N_36119,N_36243);
or U36339 (N_36339,N_36180,N_36219);
and U36340 (N_36340,N_36000,N_36218);
and U36341 (N_36341,N_36006,N_36043);
xnor U36342 (N_36342,N_36128,N_36204);
or U36343 (N_36343,N_36152,N_36177);
nand U36344 (N_36344,N_36134,N_36056);
nand U36345 (N_36345,N_36050,N_36132);
or U36346 (N_36346,N_36073,N_36151);
nand U36347 (N_36347,N_36109,N_36117);
nor U36348 (N_36348,N_36187,N_36149);
xor U36349 (N_36349,N_36011,N_36145);
xnor U36350 (N_36350,N_36055,N_36047);
or U36351 (N_36351,N_36194,N_36054);
xor U36352 (N_36352,N_36189,N_36019);
nor U36353 (N_36353,N_36005,N_36155);
nand U36354 (N_36354,N_36105,N_36022);
nand U36355 (N_36355,N_36188,N_36063);
and U36356 (N_36356,N_36190,N_36229);
nor U36357 (N_36357,N_36211,N_36116);
and U36358 (N_36358,N_36168,N_36062);
or U36359 (N_36359,N_36061,N_36099);
nand U36360 (N_36360,N_36165,N_36094);
nand U36361 (N_36361,N_36041,N_36141);
or U36362 (N_36362,N_36242,N_36098);
nand U36363 (N_36363,N_36064,N_36066);
or U36364 (N_36364,N_36067,N_36045);
nand U36365 (N_36365,N_36088,N_36107);
and U36366 (N_36366,N_36002,N_36236);
or U36367 (N_36367,N_36112,N_36186);
or U36368 (N_36368,N_36143,N_36249);
xor U36369 (N_36369,N_36207,N_36160);
xnor U36370 (N_36370,N_36162,N_36138);
or U36371 (N_36371,N_36171,N_36214);
nand U36372 (N_36372,N_36212,N_36024);
and U36373 (N_36373,N_36086,N_36241);
nor U36374 (N_36374,N_36014,N_36021);
and U36375 (N_36375,N_36123,N_36185);
or U36376 (N_36376,N_36096,N_36053);
nand U36377 (N_36377,N_36157,N_36182);
nor U36378 (N_36378,N_36148,N_36218);
and U36379 (N_36379,N_36116,N_36136);
nand U36380 (N_36380,N_36233,N_36061);
and U36381 (N_36381,N_36089,N_36198);
or U36382 (N_36382,N_36184,N_36151);
and U36383 (N_36383,N_36110,N_36002);
xor U36384 (N_36384,N_36048,N_36192);
and U36385 (N_36385,N_36218,N_36204);
and U36386 (N_36386,N_36112,N_36102);
nand U36387 (N_36387,N_36042,N_36169);
nand U36388 (N_36388,N_36213,N_36169);
nand U36389 (N_36389,N_36223,N_36182);
nor U36390 (N_36390,N_36235,N_36068);
nand U36391 (N_36391,N_36107,N_36068);
and U36392 (N_36392,N_36097,N_36139);
or U36393 (N_36393,N_36012,N_36007);
nand U36394 (N_36394,N_36075,N_36161);
or U36395 (N_36395,N_36177,N_36121);
or U36396 (N_36396,N_36211,N_36088);
and U36397 (N_36397,N_36135,N_36167);
xor U36398 (N_36398,N_36016,N_36093);
xnor U36399 (N_36399,N_36111,N_36124);
or U36400 (N_36400,N_36142,N_36069);
nor U36401 (N_36401,N_36088,N_36210);
and U36402 (N_36402,N_36156,N_36167);
or U36403 (N_36403,N_36136,N_36027);
xnor U36404 (N_36404,N_36143,N_36119);
and U36405 (N_36405,N_36198,N_36041);
or U36406 (N_36406,N_36166,N_36236);
and U36407 (N_36407,N_36220,N_36207);
or U36408 (N_36408,N_36028,N_36219);
and U36409 (N_36409,N_36163,N_36242);
nor U36410 (N_36410,N_36040,N_36206);
xor U36411 (N_36411,N_36116,N_36229);
or U36412 (N_36412,N_36139,N_36020);
or U36413 (N_36413,N_36009,N_36182);
nand U36414 (N_36414,N_36145,N_36026);
or U36415 (N_36415,N_36018,N_36127);
xor U36416 (N_36416,N_36115,N_36133);
xor U36417 (N_36417,N_36208,N_36114);
or U36418 (N_36418,N_36068,N_36006);
nand U36419 (N_36419,N_36021,N_36246);
xnor U36420 (N_36420,N_36084,N_36234);
xnor U36421 (N_36421,N_36021,N_36139);
or U36422 (N_36422,N_36060,N_36158);
nor U36423 (N_36423,N_36223,N_36136);
and U36424 (N_36424,N_36069,N_36059);
nor U36425 (N_36425,N_36107,N_36085);
xnor U36426 (N_36426,N_36008,N_36075);
and U36427 (N_36427,N_36175,N_36110);
nor U36428 (N_36428,N_36176,N_36146);
xnor U36429 (N_36429,N_36221,N_36090);
xor U36430 (N_36430,N_36054,N_36191);
nand U36431 (N_36431,N_36087,N_36013);
nor U36432 (N_36432,N_36181,N_36116);
nor U36433 (N_36433,N_36045,N_36087);
and U36434 (N_36434,N_36242,N_36009);
xnor U36435 (N_36435,N_36248,N_36162);
nand U36436 (N_36436,N_36118,N_36209);
nor U36437 (N_36437,N_36099,N_36160);
and U36438 (N_36438,N_36098,N_36099);
nand U36439 (N_36439,N_36003,N_36191);
nor U36440 (N_36440,N_36124,N_36012);
or U36441 (N_36441,N_36107,N_36214);
or U36442 (N_36442,N_36186,N_36199);
xnor U36443 (N_36443,N_36179,N_36028);
and U36444 (N_36444,N_36060,N_36141);
and U36445 (N_36445,N_36067,N_36003);
and U36446 (N_36446,N_36115,N_36110);
nor U36447 (N_36447,N_36239,N_36086);
and U36448 (N_36448,N_36041,N_36162);
xnor U36449 (N_36449,N_36133,N_36123);
nor U36450 (N_36450,N_36159,N_36148);
nand U36451 (N_36451,N_36170,N_36053);
and U36452 (N_36452,N_36203,N_36064);
nor U36453 (N_36453,N_36011,N_36224);
and U36454 (N_36454,N_36124,N_36015);
nor U36455 (N_36455,N_36006,N_36149);
and U36456 (N_36456,N_36189,N_36177);
and U36457 (N_36457,N_36041,N_36173);
nand U36458 (N_36458,N_36147,N_36109);
nand U36459 (N_36459,N_36101,N_36115);
xnor U36460 (N_36460,N_36167,N_36111);
or U36461 (N_36461,N_36132,N_36053);
xnor U36462 (N_36462,N_36141,N_36134);
and U36463 (N_36463,N_36217,N_36102);
xnor U36464 (N_36464,N_36134,N_36091);
nand U36465 (N_36465,N_36224,N_36216);
and U36466 (N_36466,N_36129,N_36173);
nor U36467 (N_36467,N_36083,N_36241);
or U36468 (N_36468,N_36121,N_36051);
nor U36469 (N_36469,N_36020,N_36247);
xnor U36470 (N_36470,N_36013,N_36031);
nand U36471 (N_36471,N_36158,N_36235);
or U36472 (N_36472,N_36141,N_36121);
xor U36473 (N_36473,N_36072,N_36146);
nor U36474 (N_36474,N_36211,N_36067);
nor U36475 (N_36475,N_36030,N_36017);
nand U36476 (N_36476,N_36028,N_36200);
or U36477 (N_36477,N_36159,N_36015);
nand U36478 (N_36478,N_36068,N_36160);
or U36479 (N_36479,N_36057,N_36045);
xnor U36480 (N_36480,N_36030,N_36183);
nand U36481 (N_36481,N_36068,N_36119);
xor U36482 (N_36482,N_36167,N_36172);
or U36483 (N_36483,N_36034,N_36088);
xnor U36484 (N_36484,N_36072,N_36238);
nand U36485 (N_36485,N_36080,N_36145);
nor U36486 (N_36486,N_36189,N_36063);
xor U36487 (N_36487,N_36236,N_36006);
xor U36488 (N_36488,N_36007,N_36093);
nand U36489 (N_36489,N_36230,N_36025);
xor U36490 (N_36490,N_36197,N_36043);
or U36491 (N_36491,N_36069,N_36182);
xnor U36492 (N_36492,N_36042,N_36088);
nand U36493 (N_36493,N_36051,N_36227);
or U36494 (N_36494,N_36200,N_36149);
and U36495 (N_36495,N_36004,N_36210);
and U36496 (N_36496,N_36191,N_36217);
xnor U36497 (N_36497,N_36135,N_36047);
nand U36498 (N_36498,N_36173,N_36053);
or U36499 (N_36499,N_36024,N_36188);
and U36500 (N_36500,N_36271,N_36252);
and U36501 (N_36501,N_36447,N_36387);
nor U36502 (N_36502,N_36379,N_36299);
nor U36503 (N_36503,N_36439,N_36281);
xor U36504 (N_36504,N_36297,N_36315);
nand U36505 (N_36505,N_36260,N_36305);
nor U36506 (N_36506,N_36329,N_36463);
nor U36507 (N_36507,N_36441,N_36433);
or U36508 (N_36508,N_36264,N_36307);
nand U36509 (N_36509,N_36266,N_36255);
xor U36510 (N_36510,N_36282,N_36383);
nand U36511 (N_36511,N_36352,N_36429);
nor U36512 (N_36512,N_36341,N_36261);
xnor U36513 (N_36513,N_36391,N_36430);
nand U36514 (N_36514,N_36306,N_36423);
nor U36515 (N_36515,N_36374,N_36390);
xnor U36516 (N_36516,N_36464,N_36342);
nor U36517 (N_36517,N_36426,N_36365);
nand U36518 (N_36518,N_36411,N_36435);
nor U36519 (N_36519,N_36388,N_36358);
nand U36520 (N_36520,N_36437,N_36468);
and U36521 (N_36521,N_36256,N_36436);
or U36522 (N_36522,N_36325,N_36488);
and U36523 (N_36523,N_36336,N_36403);
nand U36524 (N_36524,N_36487,N_36348);
or U36525 (N_36525,N_36289,N_36253);
or U36526 (N_36526,N_36449,N_36398);
xor U36527 (N_36527,N_36312,N_36380);
or U36528 (N_36528,N_36457,N_36345);
and U36529 (N_36529,N_36385,N_36482);
xnor U36530 (N_36530,N_36273,N_36375);
nor U36531 (N_36531,N_36351,N_36421);
or U36532 (N_36532,N_36276,N_36400);
and U36533 (N_36533,N_36294,N_36443);
nor U36534 (N_36534,N_36369,N_36343);
or U36535 (N_36535,N_36347,N_36378);
nand U36536 (N_36536,N_36459,N_36491);
nor U36537 (N_36537,N_36458,N_36384);
nand U36538 (N_36538,N_36431,N_36417);
xnor U36539 (N_36539,N_36427,N_36267);
xnor U36540 (N_36540,N_36399,N_36333);
nor U36541 (N_36541,N_36259,N_36445);
nand U36542 (N_36542,N_36476,N_36360);
and U36543 (N_36543,N_36422,N_36469);
nand U36544 (N_36544,N_36442,N_36381);
nand U36545 (N_36545,N_36453,N_36461);
or U36546 (N_36546,N_36283,N_36250);
or U36547 (N_36547,N_36269,N_36415);
nor U36548 (N_36548,N_36328,N_36257);
xnor U36549 (N_36549,N_36414,N_36296);
nor U36550 (N_36550,N_36394,N_36489);
xor U36551 (N_36551,N_36478,N_36335);
nand U36552 (N_36552,N_36475,N_36485);
xnor U36553 (N_36553,N_36410,N_36324);
nor U36554 (N_36554,N_36496,N_36254);
nand U36555 (N_36555,N_36304,N_36474);
xor U36556 (N_36556,N_36331,N_36288);
nand U36557 (N_36557,N_36494,N_36327);
nand U36558 (N_36558,N_36302,N_36479);
nand U36559 (N_36559,N_36330,N_36280);
and U36560 (N_36560,N_36405,N_36492);
and U36561 (N_36561,N_36319,N_36397);
or U36562 (N_36562,N_36450,N_36285);
and U36563 (N_36563,N_36300,N_36301);
and U36564 (N_36564,N_36396,N_36310);
xor U36565 (N_36565,N_36408,N_36291);
nor U36566 (N_36566,N_36362,N_36371);
nand U36567 (N_36567,N_36434,N_36293);
nor U36568 (N_36568,N_36262,N_36286);
or U36569 (N_36569,N_36356,N_36424);
and U36570 (N_36570,N_36277,N_36298);
nor U36571 (N_36571,N_36361,N_36344);
nor U36572 (N_36572,N_36455,N_36389);
nand U36573 (N_36573,N_36416,N_36486);
and U36574 (N_36574,N_36418,N_36359);
nor U36575 (N_36575,N_36338,N_36373);
nor U36576 (N_36576,N_36406,N_36466);
xnor U36577 (N_36577,N_36386,N_36484);
or U36578 (N_36578,N_36263,N_36340);
xor U36579 (N_36579,N_36368,N_36446);
and U36580 (N_36580,N_36311,N_36448);
or U36581 (N_36581,N_36355,N_36275);
xor U36582 (N_36582,N_36470,N_36320);
nor U36583 (N_36583,N_36287,N_36454);
or U36584 (N_36584,N_36495,N_36308);
and U36585 (N_36585,N_36372,N_36357);
nor U36586 (N_36586,N_36465,N_36377);
nand U36587 (N_36587,N_36364,N_36425);
nor U36588 (N_36588,N_36498,N_36323);
and U36589 (N_36589,N_36317,N_36313);
nand U36590 (N_36590,N_36270,N_36303);
nand U36591 (N_36591,N_36451,N_36346);
and U36592 (N_36592,N_36392,N_36318);
nand U36593 (N_36593,N_36472,N_36265);
xnor U36594 (N_36594,N_36353,N_36395);
xor U36595 (N_36595,N_36409,N_36490);
xnor U36596 (N_36596,N_36493,N_36284);
nand U36597 (N_36597,N_36393,N_36258);
and U36598 (N_36598,N_36321,N_36367);
xor U36599 (N_36599,N_36272,N_36295);
xor U36600 (N_36600,N_36290,N_36322);
nor U36601 (N_36601,N_36382,N_36404);
nand U36602 (N_36602,N_36363,N_36477);
and U36603 (N_36603,N_36268,N_36292);
nand U36604 (N_36604,N_36462,N_36370);
and U36605 (N_36605,N_36420,N_36444);
and U36606 (N_36606,N_36402,N_36350);
and U36607 (N_36607,N_36376,N_36460);
or U36608 (N_36608,N_36334,N_36401);
or U36609 (N_36609,N_36497,N_36366);
nand U36610 (N_36610,N_36412,N_36279);
xor U36611 (N_36611,N_36432,N_36438);
xor U36612 (N_36612,N_36332,N_36499);
nand U36613 (N_36613,N_36483,N_36452);
nand U36614 (N_36614,N_36354,N_36339);
and U36615 (N_36615,N_36407,N_36428);
nand U36616 (N_36616,N_36471,N_36349);
and U36617 (N_36617,N_36419,N_36456);
and U36618 (N_36618,N_36413,N_36309);
or U36619 (N_36619,N_36467,N_36480);
nand U36620 (N_36620,N_36473,N_36481);
and U36621 (N_36621,N_36251,N_36440);
nand U36622 (N_36622,N_36314,N_36278);
and U36623 (N_36623,N_36274,N_36316);
or U36624 (N_36624,N_36326,N_36337);
and U36625 (N_36625,N_36394,N_36445);
nand U36626 (N_36626,N_36275,N_36331);
and U36627 (N_36627,N_36334,N_36391);
or U36628 (N_36628,N_36301,N_36278);
or U36629 (N_36629,N_36374,N_36312);
or U36630 (N_36630,N_36455,N_36313);
and U36631 (N_36631,N_36445,N_36497);
and U36632 (N_36632,N_36369,N_36330);
nor U36633 (N_36633,N_36398,N_36399);
and U36634 (N_36634,N_36262,N_36338);
nor U36635 (N_36635,N_36333,N_36286);
or U36636 (N_36636,N_36345,N_36409);
and U36637 (N_36637,N_36396,N_36294);
xor U36638 (N_36638,N_36337,N_36348);
nand U36639 (N_36639,N_36296,N_36402);
or U36640 (N_36640,N_36272,N_36466);
nand U36641 (N_36641,N_36381,N_36320);
xor U36642 (N_36642,N_36450,N_36458);
and U36643 (N_36643,N_36381,N_36394);
or U36644 (N_36644,N_36343,N_36399);
xor U36645 (N_36645,N_36438,N_36313);
xor U36646 (N_36646,N_36329,N_36405);
nand U36647 (N_36647,N_36329,N_36485);
xnor U36648 (N_36648,N_36364,N_36339);
nor U36649 (N_36649,N_36408,N_36255);
and U36650 (N_36650,N_36376,N_36350);
nand U36651 (N_36651,N_36380,N_36291);
nor U36652 (N_36652,N_36261,N_36256);
or U36653 (N_36653,N_36403,N_36457);
xnor U36654 (N_36654,N_36311,N_36276);
nor U36655 (N_36655,N_36263,N_36388);
or U36656 (N_36656,N_36366,N_36486);
or U36657 (N_36657,N_36309,N_36447);
and U36658 (N_36658,N_36372,N_36420);
xor U36659 (N_36659,N_36275,N_36335);
or U36660 (N_36660,N_36334,N_36317);
nor U36661 (N_36661,N_36263,N_36355);
nand U36662 (N_36662,N_36308,N_36477);
and U36663 (N_36663,N_36269,N_36318);
and U36664 (N_36664,N_36385,N_36337);
or U36665 (N_36665,N_36250,N_36481);
or U36666 (N_36666,N_36338,N_36423);
xnor U36667 (N_36667,N_36304,N_36312);
xnor U36668 (N_36668,N_36386,N_36492);
and U36669 (N_36669,N_36419,N_36368);
nand U36670 (N_36670,N_36414,N_36358);
nand U36671 (N_36671,N_36393,N_36284);
or U36672 (N_36672,N_36465,N_36353);
and U36673 (N_36673,N_36315,N_36488);
xor U36674 (N_36674,N_36418,N_36444);
or U36675 (N_36675,N_36296,N_36499);
and U36676 (N_36676,N_36465,N_36364);
nand U36677 (N_36677,N_36409,N_36405);
or U36678 (N_36678,N_36478,N_36294);
nor U36679 (N_36679,N_36437,N_36493);
and U36680 (N_36680,N_36292,N_36465);
or U36681 (N_36681,N_36458,N_36273);
nor U36682 (N_36682,N_36438,N_36378);
and U36683 (N_36683,N_36496,N_36469);
and U36684 (N_36684,N_36431,N_36254);
nor U36685 (N_36685,N_36406,N_36359);
nand U36686 (N_36686,N_36305,N_36320);
nor U36687 (N_36687,N_36316,N_36258);
and U36688 (N_36688,N_36271,N_36374);
and U36689 (N_36689,N_36454,N_36471);
nor U36690 (N_36690,N_36343,N_36497);
xnor U36691 (N_36691,N_36331,N_36342);
xnor U36692 (N_36692,N_36293,N_36416);
nand U36693 (N_36693,N_36458,N_36472);
xnor U36694 (N_36694,N_36387,N_36449);
xnor U36695 (N_36695,N_36291,N_36494);
nand U36696 (N_36696,N_36384,N_36362);
and U36697 (N_36697,N_36262,N_36408);
nor U36698 (N_36698,N_36486,N_36305);
and U36699 (N_36699,N_36465,N_36477);
nand U36700 (N_36700,N_36310,N_36319);
nor U36701 (N_36701,N_36291,N_36438);
or U36702 (N_36702,N_36396,N_36401);
or U36703 (N_36703,N_36356,N_36476);
or U36704 (N_36704,N_36402,N_36263);
nor U36705 (N_36705,N_36305,N_36322);
or U36706 (N_36706,N_36266,N_36318);
or U36707 (N_36707,N_36356,N_36265);
xnor U36708 (N_36708,N_36314,N_36274);
nor U36709 (N_36709,N_36355,N_36362);
xnor U36710 (N_36710,N_36356,N_36392);
and U36711 (N_36711,N_36452,N_36473);
or U36712 (N_36712,N_36343,N_36465);
nand U36713 (N_36713,N_36399,N_36410);
nor U36714 (N_36714,N_36296,N_36373);
nor U36715 (N_36715,N_36452,N_36272);
nor U36716 (N_36716,N_36456,N_36404);
nor U36717 (N_36717,N_36374,N_36303);
xnor U36718 (N_36718,N_36290,N_36396);
and U36719 (N_36719,N_36445,N_36427);
xor U36720 (N_36720,N_36317,N_36388);
and U36721 (N_36721,N_36324,N_36459);
or U36722 (N_36722,N_36275,N_36417);
nor U36723 (N_36723,N_36442,N_36479);
and U36724 (N_36724,N_36422,N_36391);
nand U36725 (N_36725,N_36265,N_36341);
nand U36726 (N_36726,N_36497,N_36393);
nand U36727 (N_36727,N_36324,N_36352);
nand U36728 (N_36728,N_36331,N_36464);
xor U36729 (N_36729,N_36287,N_36336);
nand U36730 (N_36730,N_36432,N_36266);
xnor U36731 (N_36731,N_36376,N_36259);
and U36732 (N_36732,N_36295,N_36325);
and U36733 (N_36733,N_36270,N_36299);
or U36734 (N_36734,N_36482,N_36273);
xnor U36735 (N_36735,N_36378,N_36450);
nand U36736 (N_36736,N_36398,N_36374);
nor U36737 (N_36737,N_36419,N_36350);
xnor U36738 (N_36738,N_36279,N_36313);
or U36739 (N_36739,N_36260,N_36442);
nor U36740 (N_36740,N_36266,N_36276);
xor U36741 (N_36741,N_36384,N_36486);
xor U36742 (N_36742,N_36342,N_36326);
and U36743 (N_36743,N_36418,N_36404);
xnor U36744 (N_36744,N_36387,N_36340);
and U36745 (N_36745,N_36278,N_36491);
or U36746 (N_36746,N_36304,N_36329);
nor U36747 (N_36747,N_36453,N_36281);
xnor U36748 (N_36748,N_36398,N_36263);
nor U36749 (N_36749,N_36497,N_36444);
nand U36750 (N_36750,N_36593,N_36532);
and U36751 (N_36751,N_36748,N_36542);
nor U36752 (N_36752,N_36676,N_36690);
nand U36753 (N_36753,N_36645,N_36728);
nor U36754 (N_36754,N_36683,N_36505);
and U36755 (N_36755,N_36732,N_36566);
or U36756 (N_36756,N_36692,N_36672);
and U36757 (N_36757,N_36580,N_36558);
xor U36758 (N_36758,N_36540,N_36638);
and U36759 (N_36759,N_36749,N_36565);
and U36760 (N_36760,N_36502,N_36698);
xnor U36761 (N_36761,N_36511,N_36605);
or U36762 (N_36762,N_36525,N_36710);
or U36763 (N_36763,N_36730,N_36648);
nand U36764 (N_36764,N_36569,N_36701);
nor U36765 (N_36765,N_36703,N_36723);
nand U36766 (N_36766,N_36623,N_36561);
and U36767 (N_36767,N_36545,N_36662);
xor U36768 (N_36768,N_36721,N_36613);
nand U36769 (N_36769,N_36520,N_36736);
and U36770 (N_36770,N_36513,N_36577);
or U36771 (N_36771,N_36504,N_36746);
or U36772 (N_36772,N_36568,N_36592);
xnor U36773 (N_36773,N_36589,N_36689);
and U36774 (N_36774,N_36691,N_36509);
or U36775 (N_36775,N_36702,N_36573);
nor U36776 (N_36776,N_36572,N_36633);
nand U36777 (N_36777,N_36590,N_36665);
nor U36778 (N_36778,N_36579,N_36621);
xnor U36779 (N_36779,N_36674,N_36680);
xor U36780 (N_36780,N_36678,N_36667);
nand U36781 (N_36781,N_36738,N_36506);
and U36782 (N_36782,N_36659,N_36503);
and U36783 (N_36783,N_36617,N_36669);
or U36784 (N_36784,N_36642,N_36534);
nor U36785 (N_36785,N_36584,N_36712);
nor U36786 (N_36786,N_36729,N_36528);
nand U36787 (N_36787,N_36629,N_36661);
and U36788 (N_36788,N_36630,N_36695);
nand U36789 (N_36789,N_36570,N_36601);
and U36790 (N_36790,N_36716,N_36640);
or U36791 (N_36791,N_36733,N_36608);
nand U36792 (N_36792,N_36521,N_36658);
xnor U36793 (N_36793,N_36596,N_36538);
nor U36794 (N_36794,N_36510,N_36527);
xor U36795 (N_36795,N_36576,N_36715);
nor U36796 (N_36796,N_36614,N_36734);
xor U36797 (N_36797,N_36536,N_36551);
and U36798 (N_36798,N_36663,N_36564);
nand U36799 (N_36799,N_36742,N_36556);
xor U36800 (N_36800,N_36516,N_36687);
xor U36801 (N_36801,N_36554,N_36660);
or U36802 (N_36802,N_36553,N_36581);
nor U36803 (N_36803,N_36681,N_36559);
nand U36804 (N_36804,N_36587,N_36644);
nand U36805 (N_36805,N_36624,N_36696);
and U36806 (N_36806,N_36620,N_36612);
or U36807 (N_36807,N_36602,N_36673);
and U36808 (N_36808,N_36567,N_36650);
nand U36809 (N_36809,N_36652,N_36731);
xor U36810 (N_36810,N_36529,N_36514);
xor U36811 (N_36811,N_36706,N_36643);
nand U36812 (N_36812,N_36607,N_36563);
nand U36813 (N_36813,N_36523,N_36726);
nor U36814 (N_36814,N_36657,N_36574);
nor U36815 (N_36815,N_36671,N_36519);
or U36816 (N_36816,N_36539,N_36699);
nand U36817 (N_36817,N_36641,N_36543);
or U36818 (N_36818,N_36526,N_36537);
xnor U36819 (N_36819,N_36597,N_36588);
nand U36820 (N_36820,N_36722,N_36595);
or U36821 (N_36821,N_36522,N_36653);
xnor U36822 (N_36822,N_36549,N_36707);
nand U36823 (N_36823,N_36560,N_36562);
nor U36824 (N_36824,N_36724,N_36649);
and U36825 (N_36825,N_36709,N_36626);
xor U36826 (N_36826,N_36725,N_36603);
or U36827 (N_36827,N_36670,N_36517);
and U36828 (N_36828,N_36741,N_36599);
xnor U36829 (N_36829,N_36524,N_36694);
nand U36830 (N_36830,N_36632,N_36664);
or U36831 (N_36831,N_36507,N_36578);
nand U36832 (N_36832,N_36541,N_36647);
and U36833 (N_36833,N_36646,N_36631);
or U36834 (N_36834,N_36708,N_36550);
nor U36835 (N_36835,N_36740,N_36591);
xor U36836 (N_36836,N_36594,N_36609);
or U36837 (N_36837,N_36552,N_36548);
and U36838 (N_36838,N_36697,N_36743);
nor U36839 (N_36839,N_36628,N_36622);
and U36840 (N_36840,N_36718,N_36693);
nand U36841 (N_36841,N_36747,N_36700);
or U36842 (N_36842,N_36704,N_36713);
and U36843 (N_36843,N_36583,N_36735);
nor U36844 (N_36844,N_36679,N_36615);
nor U36845 (N_36845,N_36546,N_36515);
and U36846 (N_36846,N_36688,N_36625);
xor U36847 (N_36847,N_36739,N_36600);
or U36848 (N_36848,N_36627,N_36727);
nand U36849 (N_36849,N_36639,N_36501);
and U36850 (N_36850,N_36705,N_36677);
nor U36851 (N_36851,N_36610,N_36711);
and U36852 (N_36852,N_36675,N_36531);
nor U36853 (N_36853,N_36655,N_36575);
nor U36854 (N_36854,N_36685,N_36555);
nor U36855 (N_36855,N_36737,N_36666);
xor U36856 (N_36856,N_36619,N_36616);
or U36857 (N_36857,N_36530,N_36618);
or U36858 (N_36858,N_36544,N_36719);
xnor U36859 (N_36859,N_36744,N_36634);
and U36860 (N_36860,N_36635,N_36557);
nor U36861 (N_36861,N_36637,N_36512);
xor U36862 (N_36862,N_36636,N_36586);
or U36863 (N_36863,N_36606,N_36656);
nor U36864 (N_36864,N_36533,N_36668);
or U36865 (N_36865,N_36714,N_36682);
nor U36866 (N_36866,N_36611,N_36720);
nor U36867 (N_36867,N_36571,N_36684);
xnor U36868 (N_36868,N_36500,N_36508);
nand U36869 (N_36869,N_36604,N_36535);
nor U36870 (N_36870,N_36717,N_36686);
and U36871 (N_36871,N_36654,N_36651);
nor U36872 (N_36872,N_36547,N_36598);
and U36873 (N_36873,N_36582,N_36585);
nand U36874 (N_36874,N_36745,N_36518);
nor U36875 (N_36875,N_36700,N_36715);
xor U36876 (N_36876,N_36694,N_36525);
and U36877 (N_36877,N_36535,N_36594);
nor U36878 (N_36878,N_36543,N_36563);
or U36879 (N_36879,N_36631,N_36721);
xnor U36880 (N_36880,N_36700,N_36606);
and U36881 (N_36881,N_36625,N_36636);
or U36882 (N_36882,N_36512,N_36580);
or U36883 (N_36883,N_36642,N_36528);
nor U36884 (N_36884,N_36687,N_36542);
nor U36885 (N_36885,N_36589,N_36517);
nand U36886 (N_36886,N_36539,N_36534);
nand U36887 (N_36887,N_36549,N_36700);
and U36888 (N_36888,N_36637,N_36740);
or U36889 (N_36889,N_36634,N_36591);
nor U36890 (N_36890,N_36544,N_36643);
or U36891 (N_36891,N_36551,N_36711);
nand U36892 (N_36892,N_36562,N_36632);
xnor U36893 (N_36893,N_36577,N_36503);
or U36894 (N_36894,N_36519,N_36574);
and U36895 (N_36895,N_36522,N_36529);
nor U36896 (N_36896,N_36718,N_36650);
nand U36897 (N_36897,N_36604,N_36658);
or U36898 (N_36898,N_36663,N_36705);
nor U36899 (N_36899,N_36590,N_36556);
xnor U36900 (N_36900,N_36706,N_36618);
nand U36901 (N_36901,N_36706,N_36686);
or U36902 (N_36902,N_36719,N_36737);
or U36903 (N_36903,N_36541,N_36716);
or U36904 (N_36904,N_36615,N_36501);
or U36905 (N_36905,N_36598,N_36625);
nand U36906 (N_36906,N_36587,N_36518);
nor U36907 (N_36907,N_36566,N_36576);
nand U36908 (N_36908,N_36642,N_36506);
nor U36909 (N_36909,N_36566,N_36575);
nand U36910 (N_36910,N_36742,N_36662);
xnor U36911 (N_36911,N_36724,N_36597);
and U36912 (N_36912,N_36721,N_36547);
or U36913 (N_36913,N_36600,N_36735);
or U36914 (N_36914,N_36613,N_36552);
and U36915 (N_36915,N_36704,N_36507);
xnor U36916 (N_36916,N_36545,N_36577);
nand U36917 (N_36917,N_36524,N_36661);
or U36918 (N_36918,N_36670,N_36525);
and U36919 (N_36919,N_36582,N_36724);
nor U36920 (N_36920,N_36660,N_36573);
or U36921 (N_36921,N_36674,N_36721);
nand U36922 (N_36922,N_36602,N_36622);
nand U36923 (N_36923,N_36699,N_36532);
xor U36924 (N_36924,N_36668,N_36727);
xor U36925 (N_36925,N_36509,N_36607);
and U36926 (N_36926,N_36585,N_36716);
or U36927 (N_36927,N_36695,N_36614);
nor U36928 (N_36928,N_36727,N_36620);
and U36929 (N_36929,N_36668,N_36525);
and U36930 (N_36930,N_36574,N_36648);
xnor U36931 (N_36931,N_36642,N_36661);
and U36932 (N_36932,N_36646,N_36744);
and U36933 (N_36933,N_36706,N_36683);
xnor U36934 (N_36934,N_36707,N_36717);
or U36935 (N_36935,N_36722,N_36507);
xor U36936 (N_36936,N_36544,N_36540);
and U36937 (N_36937,N_36692,N_36688);
and U36938 (N_36938,N_36715,N_36598);
nand U36939 (N_36939,N_36579,N_36652);
nand U36940 (N_36940,N_36586,N_36682);
nand U36941 (N_36941,N_36517,N_36685);
nand U36942 (N_36942,N_36607,N_36500);
nor U36943 (N_36943,N_36742,N_36741);
nand U36944 (N_36944,N_36585,N_36624);
or U36945 (N_36945,N_36530,N_36676);
or U36946 (N_36946,N_36569,N_36699);
and U36947 (N_36947,N_36719,N_36727);
and U36948 (N_36948,N_36654,N_36658);
nor U36949 (N_36949,N_36718,N_36555);
nor U36950 (N_36950,N_36503,N_36720);
and U36951 (N_36951,N_36691,N_36702);
and U36952 (N_36952,N_36517,N_36675);
nor U36953 (N_36953,N_36597,N_36570);
xor U36954 (N_36954,N_36529,N_36535);
nand U36955 (N_36955,N_36696,N_36671);
nor U36956 (N_36956,N_36625,N_36522);
nand U36957 (N_36957,N_36673,N_36628);
nand U36958 (N_36958,N_36747,N_36540);
or U36959 (N_36959,N_36668,N_36548);
xor U36960 (N_36960,N_36677,N_36607);
or U36961 (N_36961,N_36555,N_36683);
or U36962 (N_36962,N_36748,N_36519);
or U36963 (N_36963,N_36651,N_36599);
or U36964 (N_36964,N_36528,N_36618);
nor U36965 (N_36965,N_36565,N_36655);
and U36966 (N_36966,N_36693,N_36609);
or U36967 (N_36967,N_36678,N_36558);
nand U36968 (N_36968,N_36641,N_36617);
nor U36969 (N_36969,N_36702,N_36711);
or U36970 (N_36970,N_36559,N_36668);
or U36971 (N_36971,N_36644,N_36552);
nand U36972 (N_36972,N_36534,N_36740);
xor U36973 (N_36973,N_36607,N_36548);
and U36974 (N_36974,N_36629,N_36634);
nand U36975 (N_36975,N_36636,N_36717);
and U36976 (N_36976,N_36651,N_36658);
and U36977 (N_36977,N_36548,N_36608);
or U36978 (N_36978,N_36627,N_36671);
nor U36979 (N_36979,N_36539,N_36580);
and U36980 (N_36980,N_36687,N_36563);
or U36981 (N_36981,N_36650,N_36633);
nand U36982 (N_36982,N_36632,N_36607);
xor U36983 (N_36983,N_36733,N_36596);
xor U36984 (N_36984,N_36734,N_36716);
and U36985 (N_36985,N_36614,N_36636);
xnor U36986 (N_36986,N_36631,N_36642);
or U36987 (N_36987,N_36542,N_36569);
and U36988 (N_36988,N_36692,N_36641);
or U36989 (N_36989,N_36677,N_36597);
or U36990 (N_36990,N_36593,N_36730);
nor U36991 (N_36991,N_36647,N_36594);
nand U36992 (N_36992,N_36530,N_36721);
nor U36993 (N_36993,N_36745,N_36610);
nand U36994 (N_36994,N_36534,N_36744);
xor U36995 (N_36995,N_36736,N_36636);
nor U36996 (N_36996,N_36715,N_36741);
nand U36997 (N_36997,N_36608,N_36537);
nand U36998 (N_36998,N_36573,N_36683);
and U36999 (N_36999,N_36539,N_36569);
nand U37000 (N_37000,N_36783,N_36865);
nand U37001 (N_37001,N_36890,N_36806);
xor U37002 (N_37002,N_36915,N_36858);
or U37003 (N_37003,N_36784,N_36863);
nand U37004 (N_37004,N_36930,N_36847);
or U37005 (N_37005,N_36904,N_36959);
nand U37006 (N_37006,N_36960,N_36855);
and U37007 (N_37007,N_36899,N_36799);
nor U37008 (N_37008,N_36763,N_36813);
or U37009 (N_37009,N_36941,N_36795);
xnor U37010 (N_37010,N_36991,N_36800);
nor U37011 (N_37011,N_36946,N_36859);
nand U37012 (N_37012,N_36797,N_36810);
or U37013 (N_37013,N_36988,N_36777);
xor U37014 (N_37014,N_36823,N_36846);
nor U37015 (N_37015,N_36754,N_36868);
or U37016 (N_37016,N_36923,N_36866);
and U37017 (N_37017,N_36822,N_36985);
xor U37018 (N_37018,N_36876,N_36798);
nand U37019 (N_37019,N_36796,N_36818);
xnor U37020 (N_37020,N_36950,N_36966);
nor U37021 (N_37021,N_36885,N_36849);
nor U37022 (N_37022,N_36881,N_36967);
nor U37023 (N_37023,N_36907,N_36860);
and U37024 (N_37024,N_36828,N_36894);
or U37025 (N_37025,N_36751,N_36755);
or U37026 (N_37026,N_36870,N_36891);
nor U37027 (N_37027,N_36943,N_36952);
nor U37028 (N_37028,N_36989,N_36794);
nand U37029 (N_37029,N_36862,N_36958);
xnor U37030 (N_37030,N_36901,N_36767);
nand U37031 (N_37031,N_36786,N_36936);
or U37032 (N_37032,N_36949,N_36775);
xnor U37033 (N_37033,N_36955,N_36909);
and U37034 (N_37034,N_36987,N_36926);
and U37035 (N_37035,N_36999,N_36853);
nand U37036 (N_37036,N_36889,N_36875);
or U37037 (N_37037,N_36932,N_36805);
nand U37038 (N_37038,N_36954,N_36919);
xnor U37039 (N_37039,N_36925,N_36938);
xor U37040 (N_37040,N_36826,N_36906);
and U37041 (N_37041,N_36788,N_36856);
and U37042 (N_37042,N_36970,N_36912);
and U37043 (N_37043,N_36933,N_36836);
nand U37044 (N_37044,N_36778,N_36848);
xor U37045 (N_37045,N_36753,N_36845);
and U37046 (N_37046,N_36965,N_36927);
and U37047 (N_37047,N_36830,N_36759);
nand U37048 (N_37048,N_36896,N_36948);
nand U37049 (N_37049,N_36838,N_36825);
and U37050 (N_37050,N_36760,N_36893);
nor U37051 (N_37051,N_36764,N_36924);
nor U37052 (N_37052,N_36977,N_36976);
xnor U37053 (N_37053,N_36808,N_36821);
or U37054 (N_37054,N_36854,N_36843);
nor U37055 (N_37055,N_36766,N_36812);
nor U37056 (N_37056,N_36990,N_36884);
nor U37057 (N_37057,N_36779,N_36971);
nor U37058 (N_37058,N_36758,N_36892);
xnor U37059 (N_37059,N_36770,N_36809);
nor U37060 (N_37060,N_36895,N_36857);
xnor U37061 (N_37061,N_36968,N_36913);
xnor U37062 (N_37062,N_36833,N_36898);
nand U37063 (N_37063,N_36761,N_36835);
or U37064 (N_37064,N_36787,N_36922);
nor U37065 (N_37065,N_36842,N_36790);
or U37066 (N_37066,N_36935,N_36752);
nand U37067 (N_37067,N_36921,N_36867);
xor U37068 (N_37068,N_36888,N_36994);
nand U37069 (N_37069,N_36887,N_36993);
nor U37070 (N_37070,N_36911,N_36781);
xnor U37071 (N_37071,N_36757,N_36807);
nor U37072 (N_37072,N_36942,N_36956);
nor U37073 (N_37073,N_36947,N_36951);
and U37074 (N_37074,N_36829,N_36773);
nor U37075 (N_37075,N_36961,N_36872);
xor U37076 (N_37076,N_36834,N_36827);
nor U37077 (N_37077,N_36840,N_36819);
and U37078 (N_37078,N_36982,N_36992);
xnor U37079 (N_37079,N_36832,N_36883);
and U37080 (N_37080,N_36864,N_36981);
or U37081 (N_37081,N_36820,N_36851);
and U37082 (N_37082,N_36979,N_36918);
or U37083 (N_37083,N_36998,N_36953);
nand U37084 (N_37084,N_36869,N_36756);
xnor U37085 (N_37085,N_36916,N_36945);
xnor U37086 (N_37086,N_36877,N_36969);
nor U37087 (N_37087,N_36995,N_36815);
xnor U37088 (N_37088,N_36850,N_36780);
and U37089 (N_37089,N_36897,N_36874);
or U37090 (N_37090,N_36785,N_36974);
and U37091 (N_37091,N_36937,N_36983);
xnor U37092 (N_37092,N_36772,N_36886);
or U37093 (N_37093,N_36975,N_36944);
and U37094 (N_37094,N_36940,N_36978);
and U37095 (N_37095,N_36928,N_36917);
and U37096 (N_37096,N_36996,N_36931);
or U37097 (N_37097,N_36750,N_36771);
or U37098 (N_37098,N_36817,N_36803);
nor U37099 (N_37099,N_36934,N_36873);
nor U37100 (N_37100,N_36880,N_36816);
nand U37101 (N_37101,N_36984,N_36972);
and U37102 (N_37102,N_36882,N_36963);
nor U37103 (N_37103,N_36765,N_36811);
nor U37104 (N_37104,N_36878,N_36871);
nand U37105 (N_37105,N_36914,N_36939);
xor U37106 (N_37106,N_36839,N_36792);
and U37107 (N_37107,N_36910,N_36782);
or U37108 (N_37108,N_36903,N_36900);
xnor U37109 (N_37109,N_36997,N_36789);
xnor U37110 (N_37110,N_36908,N_36962);
nor U37111 (N_37111,N_36964,N_36791);
and U37112 (N_37112,N_36837,N_36920);
and U37113 (N_37113,N_36776,N_36986);
or U37114 (N_37114,N_36861,N_36902);
or U37115 (N_37115,N_36804,N_36929);
and U37116 (N_37116,N_36852,N_36802);
xor U37117 (N_37117,N_36801,N_36957);
and U37118 (N_37118,N_36973,N_36824);
and U37119 (N_37119,N_36905,N_36768);
nor U37120 (N_37120,N_36814,N_36774);
nand U37121 (N_37121,N_36844,N_36793);
nor U37122 (N_37122,N_36762,N_36980);
nand U37123 (N_37123,N_36841,N_36769);
or U37124 (N_37124,N_36879,N_36831);
nand U37125 (N_37125,N_36990,N_36917);
and U37126 (N_37126,N_36791,N_36797);
and U37127 (N_37127,N_36768,N_36765);
xor U37128 (N_37128,N_36833,N_36962);
xnor U37129 (N_37129,N_36930,N_36838);
nor U37130 (N_37130,N_36777,N_36948);
or U37131 (N_37131,N_36989,N_36944);
nand U37132 (N_37132,N_36853,N_36969);
nand U37133 (N_37133,N_36968,N_36940);
or U37134 (N_37134,N_36890,N_36965);
or U37135 (N_37135,N_36878,N_36981);
nand U37136 (N_37136,N_36776,N_36884);
nand U37137 (N_37137,N_36967,N_36788);
or U37138 (N_37138,N_36970,N_36765);
xnor U37139 (N_37139,N_36757,N_36784);
nand U37140 (N_37140,N_36970,N_36920);
nand U37141 (N_37141,N_36833,N_36965);
and U37142 (N_37142,N_36787,N_36939);
xnor U37143 (N_37143,N_36776,N_36795);
nand U37144 (N_37144,N_36948,N_36764);
nor U37145 (N_37145,N_36770,N_36802);
or U37146 (N_37146,N_36899,N_36939);
or U37147 (N_37147,N_36969,N_36762);
xor U37148 (N_37148,N_36921,N_36777);
nor U37149 (N_37149,N_36959,N_36923);
nor U37150 (N_37150,N_36832,N_36953);
or U37151 (N_37151,N_36833,N_36982);
nor U37152 (N_37152,N_36944,N_36757);
or U37153 (N_37153,N_36835,N_36823);
or U37154 (N_37154,N_36750,N_36797);
nor U37155 (N_37155,N_36770,N_36868);
and U37156 (N_37156,N_36761,N_36992);
or U37157 (N_37157,N_36803,N_36876);
xor U37158 (N_37158,N_36796,N_36803);
and U37159 (N_37159,N_36931,N_36750);
and U37160 (N_37160,N_36760,N_36889);
and U37161 (N_37161,N_36863,N_36995);
xnor U37162 (N_37162,N_36827,N_36823);
or U37163 (N_37163,N_36947,N_36977);
nand U37164 (N_37164,N_36987,N_36822);
xnor U37165 (N_37165,N_36986,N_36831);
and U37166 (N_37166,N_36897,N_36839);
and U37167 (N_37167,N_36813,N_36980);
and U37168 (N_37168,N_36928,N_36778);
nand U37169 (N_37169,N_36996,N_36824);
or U37170 (N_37170,N_36922,N_36762);
and U37171 (N_37171,N_36839,N_36834);
xor U37172 (N_37172,N_36920,N_36900);
nand U37173 (N_37173,N_36806,N_36924);
nand U37174 (N_37174,N_36855,N_36815);
nor U37175 (N_37175,N_36934,N_36923);
and U37176 (N_37176,N_36957,N_36950);
nand U37177 (N_37177,N_36846,N_36950);
nand U37178 (N_37178,N_36857,N_36821);
or U37179 (N_37179,N_36852,N_36862);
or U37180 (N_37180,N_36906,N_36894);
xor U37181 (N_37181,N_36755,N_36830);
and U37182 (N_37182,N_36872,N_36867);
nor U37183 (N_37183,N_36773,N_36828);
nor U37184 (N_37184,N_36771,N_36790);
nand U37185 (N_37185,N_36976,N_36958);
nand U37186 (N_37186,N_36884,N_36923);
xnor U37187 (N_37187,N_36773,N_36935);
or U37188 (N_37188,N_36850,N_36800);
xnor U37189 (N_37189,N_36903,N_36958);
or U37190 (N_37190,N_36833,N_36967);
or U37191 (N_37191,N_36976,N_36985);
nand U37192 (N_37192,N_36836,N_36852);
xnor U37193 (N_37193,N_36777,N_36971);
xnor U37194 (N_37194,N_36959,N_36965);
or U37195 (N_37195,N_36907,N_36967);
nor U37196 (N_37196,N_36784,N_36925);
or U37197 (N_37197,N_36986,N_36891);
xnor U37198 (N_37198,N_36872,N_36874);
or U37199 (N_37199,N_36944,N_36774);
xnor U37200 (N_37200,N_36984,N_36827);
xnor U37201 (N_37201,N_36992,N_36897);
nand U37202 (N_37202,N_36881,N_36827);
or U37203 (N_37203,N_36868,N_36926);
or U37204 (N_37204,N_36846,N_36932);
xnor U37205 (N_37205,N_36771,N_36850);
xnor U37206 (N_37206,N_36869,N_36955);
and U37207 (N_37207,N_36787,N_36836);
and U37208 (N_37208,N_36892,N_36787);
and U37209 (N_37209,N_36795,N_36888);
xor U37210 (N_37210,N_36834,N_36879);
nand U37211 (N_37211,N_36765,N_36909);
and U37212 (N_37212,N_36761,N_36942);
and U37213 (N_37213,N_36946,N_36803);
xor U37214 (N_37214,N_36918,N_36861);
xor U37215 (N_37215,N_36779,N_36794);
or U37216 (N_37216,N_36860,N_36891);
and U37217 (N_37217,N_36766,N_36897);
or U37218 (N_37218,N_36764,N_36879);
nand U37219 (N_37219,N_36792,N_36810);
nor U37220 (N_37220,N_36995,N_36784);
xnor U37221 (N_37221,N_36986,N_36871);
or U37222 (N_37222,N_36783,N_36921);
or U37223 (N_37223,N_36875,N_36870);
and U37224 (N_37224,N_36920,N_36923);
or U37225 (N_37225,N_36979,N_36909);
nand U37226 (N_37226,N_36826,N_36950);
and U37227 (N_37227,N_36851,N_36836);
nor U37228 (N_37228,N_36781,N_36941);
nor U37229 (N_37229,N_36774,N_36760);
xor U37230 (N_37230,N_36861,N_36831);
xnor U37231 (N_37231,N_36964,N_36858);
xor U37232 (N_37232,N_36838,N_36897);
and U37233 (N_37233,N_36970,N_36952);
and U37234 (N_37234,N_36990,N_36984);
nand U37235 (N_37235,N_36848,N_36929);
and U37236 (N_37236,N_36853,N_36785);
nor U37237 (N_37237,N_36953,N_36866);
xor U37238 (N_37238,N_36765,N_36875);
nor U37239 (N_37239,N_36900,N_36787);
and U37240 (N_37240,N_36946,N_36983);
nor U37241 (N_37241,N_36944,N_36968);
xnor U37242 (N_37242,N_36859,N_36954);
and U37243 (N_37243,N_36857,N_36776);
xnor U37244 (N_37244,N_36961,N_36853);
xnor U37245 (N_37245,N_36993,N_36975);
or U37246 (N_37246,N_36831,N_36779);
nand U37247 (N_37247,N_36937,N_36967);
nor U37248 (N_37248,N_36931,N_36896);
nor U37249 (N_37249,N_36796,N_36966);
xnor U37250 (N_37250,N_37018,N_37237);
nor U37251 (N_37251,N_37175,N_37130);
nor U37252 (N_37252,N_37203,N_37110);
xor U37253 (N_37253,N_37019,N_37092);
nand U37254 (N_37254,N_37173,N_37072);
and U37255 (N_37255,N_37049,N_37157);
xnor U37256 (N_37256,N_37042,N_37161);
xor U37257 (N_37257,N_37016,N_37166);
xor U37258 (N_37258,N_37176,N_37105);
and U37259 (N_37259,N_37025,N_37073);
and U37260 (N_37260,N_37233,N_37172);
and U37261 (N_37261,N_37099,N_37195);
nand U37262 (N_37262,N_37070,N_37201);
nor U37263 (N_37263,N_37200,N_37167);
nand U37264 (N_37264,N_37053,N_37026);
or U37265 (N_37265,N_37163,N_37035);
nand U37266 (N_37266,N_37226,N_37214);
or U37267 (N_37267,N_37224,N_37032);
nor U37268 (N_37268,N_37148,N_37075);
and U37269 (N_37269,N_37169,N_37074);
or U37270 (N_37270,N_37164,N_37118);
xor U37271 (N_37271,N_37139,N_37225);
or U37272 (N_37272,N_37242,N_37121);
and U37273 (N_37273,N_37227,N_37159);
nand U37274 (N_37274,N_37141,N_37085);
nor U37275 (N_37275,N_37089,N_37207);
nor U37276 (N_37276,N_37205,N_37097);
nand U37277 (N_37277,N_37014,N_37189);
xnor U37278 (N_37278,N_37088,N_37180);
xnor U37279 (N_37279,N_37082,N_37142);
or U37280 (N_37280,N_37048,N_37236);
nand U37281 (N_37281,N_37184,N_37125);
nand U37282 (N_37282,N_37179,N_37137);
or U37283 (N_37283,N_37196,N_37245);
nand U37284 (N_37284,N_37243,N_37024);
or U37285 (N_37285,N_37101,N_37168);
and U37286 (N_37286,N_37037,N_37104);
nor U37287 (N_37287,N_37140,N_37124);
nand U37288 (N_37288,N_37108,N_37079);
nand U37289 (N_37289,N_37011,N_37191);
nor U37290 (N_37290,N_37229,N_37199);
or U37291 (N_37291,N_37244,N_37246);
nand U37292 (N_37292,N_37057,N_37030);
xnor U37293 (N_37293,N_37007,N_37190);
and U37294 (N_37294,N_37083,N_37028);
and U37295 (N_37295,N_37249,N_37065);
nand U37296 (N_37296,N_37232,N_37036);
xnor U37297 (N_37297,N_37114,N_37020);
or U37298 (N_37298,N_37174,N_37235);
nand U37299 (N_37299,N_37132,N_37146);
or U37300 (N_37300,N_37153,N_37023);
or U37301 (N_37301,N_37033,N_37106);
xor U37302 (N_37302,N_37116,N_37077);
nand U37303 (N_37303,N_37021,N_37107);
or U37304 (N_37304,N_37050,N_37147);
nor U37305 (N_37305,N_37134,N_37046);
xnor U37306 (N_37306,N_37177,N_37160);
nand U37307 (N_37307,N_37061,N_37034);
nor U37308 (N_37308,N_37194,N_37043);
or U37309 (N_37309,N_37091,N_37223);
nand U37310 (N_37310,N_37062,N_37185);
nand U37311 (N_37311,N_37067,N_37170);
nand U37312 (N_37312,N_37239,N_37238);
xnor U37313 (N_37313,N_37133,N_37013);
nand U37314 (N_37314,N_37197,N_37060);
xnor U37315 (N_37315,N_37186,N_37071);
nor U37316 (N_37316,N_37211,N_37178);
nand U37317 (N_37317,N_37248,N_37206);
nor U37318 (N_37318,N_37158,N_37230);
nor U37319 (N_37319,N_37188,N_37216);
and U37320 (N_37320,N_37111,N_37187);
xor U37321 (N_37321,N_37241,N_37064);
nand U37322 (N_37322,N_37068,N_37156);
nor U37323 (N_37323,N_37222,N_37240);
or U37324 (N_37324,N_37117,N_37165);
or U37325 (N_37325,N_37144,N_37182);
nor U37326 (N_37326,N_37078,N_37202);
nor U37327 (N_37327,N_37131,N_37002);
nor U37328 (N_37328,N_37228,N_37076);
xnor U37329 (N_37329,N_37171,N_37152);
xor U37330 (N_37330,N_37059,N_37119);
nand U37331 (N_37331,N_37192,N_37154);
or U37332 (N_37332,N_37041,N_37127);
xor U37333 (N_37333,N_37098,N_37029);
or U37334 (N_37334,N_37058,N_37008);
nor U37335 (N_37335,N_37006,N_37220);
and U37336 (N_37336,N_37056,N_37090);
and U37337 (N_37337,N_37138,N_37219);
or U37338 (N_37338,N_37247,N_37069);
and U37339 (N_37339,N_37109,N_37151);
xor U37340 (N_37340,N_37123,N_37198);
or U37341 (N_37341,N_37149,N_37155);
or U37342 (N_37342,N_37093,N_37015);
and U37343 (N_37343,N_37055,N_37081);
nand U37344 (N_37344,N_37150,N_37003);
nand U37345 (N_37345,N_37215,N_37038);
or U37346 (N_37346,N_37066,N_37122);
xor U37347 (N_37347,N_37183,N_37017);
nor U37348 (N_37348,N_37095,N_37231);
or U37349 (N_37349,N_37045,N_37162);
and U37350 (N_37350,N_37126,N_37112);
or U37351 (N_37351,N_37009,N_37052);
nor U37352 (N_37352,N_37193,N_37102);
xnor U37353 (N_37353,N_37031,N_37209);
or U37354 (N_37354,N_37039,N_37000);
or U37355 (N_37355,N_37103,N_37136);
nand U37356 (N_37356,N_37218,N_37001);
nand U37357 (N_37357,N_37234,N_37084);
xnor U37358 (N_37358,N_37221,N_37120);
nor U37359 (N_37359,N_37094,N_37145);
or U37360 (N_37360,N_37113,N_37135);
nor U37361 (N_37361,N_37213,N_37063);
or U37362 (N_37362,N_37040,N_37010);
and U37363 (N_37363,N_37143,N_37210);
xor U37364 (N_37364,N_37212,N_37129);
xnor U37365 (N_37365,N_37051,N_37100);
nor U37366 (N_37366,N_37115,N_37004);
nor U37367 (N_37367,N_37087,N_37080);
or U37368 (N_37368,N_37217,N_37005);
and U37369 (N_37369,N_37208,N_37047);
nor U37370 (N_37370,N_37054,N_37204);
nand U37371 (N_37371,N_37086,N_37012);
xor U37372 (N_37372,N_37044,N_37128);
and U37373 (N_37373,N_37181,N_37096);
xnor U37374 (N_37374,N_37022,N_37027);
nor U37375 (N_37375,N_37085,N_37233);
nand U37376 (N_37376,N_37190,N_37235);
and U37377 (N_37377,N_37059,N_37037);
and U37378 (N_37378,N_37245,N_37035);
nor U37379 (N_37379,N_37125,N_37194);
or U37380 (N_37380,N_37073,N_37024);
and U37381 (N_37381,N_37122,N_37146);
nor U37382 (N_37382,N_37196,N_37059);
xor U37383 (N_37383,N_37205,N_37079);
nand U37384 (N_37384,N_37185,N_37105);
nor U37385 (N_37385,N_37164,N_37114);
nand U37386 (N_37386,N_37152,N_37231);
or U37387 (N_37387,N_37029,N_37069);
nand U37388 (N_37388,N_37075,N_37100);
and U37389 (N_37389,N_37236,N_37241);
nand U37390 (N_37390,N_37118,N_37241);
and U37391 (N_37391,N_37038,N_37200);
nor U37392 (N_37392,N_37099,N_37223);
and U37393 (N_37393,N_37128,N_37162);
or U37394 (N_37394,N_37097,N_37222);
and U37395 (N_37395,N_37186,N_37195);
nor U37396 (N_37396,N_37174,N_37017);
xnor U37397 (N_37397,N_37109,N_37106);
nand U37398 (N_37398,N_37087,N_37221);
nor U37399 (N_37399,N_37130,N_37014);
nand U37400 (N_37400,N_37035,N_37180);
or U37401 (N_37401,N_37052,N_37105);
xnor U37402 (N_37402,N_37111,N_37046);
or U37403 (N_37403,N_37160,N_37049);
nand U37404 (N_37404,N_37162,N_37008);
nand U37405 (N_37405,N_37025,N_37135);
or U37406 (N_37406,N_37146,N_37028);
and U37407 (N_37407,N_37146,N_37068);
and U37408 (N_37408,N_37127,N_37148);
nor U37409 (N_37409,N_37071,N_37087);
nand U37410 (N_37410,N_37141,N_37117);
xor U37411 (N_37411,N_37002,N_37186);
nor U37412 (N_37412,N_37075,N_37184);
xor U37413 (N_37413,N_37176,N_37182);
and U37414 (N_37414,N_37120,N_37127);
nor U37415 (N_37415,N_37129,N_37135);
and U37416 (N_37416,N_37020,N_37169);
and U37417 (N_37417,N_37192,N_37171);
and U37418 (N_37418,N_37246,N_37190);
nand U37419 (N_37419,N_37176,N_37169);
nor U37420 (N_37420,N_37112,N_37067);
and U37421 (N_37421,N_37101,N_37044);
and U37422 (N_37422,N_37065,N_37120);
nand U37423 (N_37423,N_37177,N_37234);
nand U37424 (N_37424,N_37151,N_37232);
and U37425 (N_37425,N_37080,N_37082);
and U37426 (N_37426,N_37171,N_37013);
nand U37427 (N_37427,N_37239,N_37058);
or U37428 (N_37428,N_37126,N_37111);
and U37429 (N_37429,N_37229,N_37071);
nand U37430 (N_37430,N_37172,N_37215);
xnor U37431 (N_37431,N_37053,N_37052);
xnor U37432 (N_37432,N_37246,N_37042);
nor U37433 (N_37433,N_37156,N_37029);
or U37434 (N_37434,N_37019,N_37178);
nor U37435 (N_37435,N_37047,N_37040);
xnor U37436 (N_37436,N_37237,N_37186);
or U37437 (N_37437,N_37045,N_37130);
nand U37438 (N_37438,N_37089,N_37200);
xor U37439 (N_37439,N_37081,N_37196);
xnor U37440 (N_37440,N_37104,N_37062);
nand U37441 (N_37441,N_37218,N_37098);
xnor U37442 (N_37442,N_37050,N_37201);
nor U37443 (N_37443,N_37117,N_37039);
xor U37444 (N_37444,N_37110,N_37023);
or U37445 (N_37445,N_37240,N_37001);
nor U37446 (N_37446,N_37087,N_37077);
xor U37447 (N_37447,N_37214,N_37113);
or U37448 (N_37448,N_37020,N_37102);
nor U37449 (N_37449,N_37229,N_37132);
nor U37450 (N_37450,N_37059,N_37111);
nor U37451 (N_37451,N_37234,N_37118);
xnor U37452 (N_37452,N_37039,N_37021);
nor U37453 (N_37453,N_37114,N_37092);
nor U37454 (N_37454,N_37029,N_37244);
nand U37455 (N_37455,N_37037,N_37127);
nor U37456 (N_37456,N_37247,N_37107);
and U37457 (N_37457,N_37199,N_37105);
or U37458 (N_37458,N_37003,N_37172);
or U37459 (N_37459,N_37107,N_37209);
nand U37460 (N_37460,N_37245,N_37027);
xor U37461 (N_37461,N_37001,N_37141);
nor U37462 (N_37462,N_37247,N_37214);
and U37463 (N_37463,N_37121,N_37222);
nand U37464 (N_37464,N_37152,N_37235);
nor U37465 (N_37465,N_37109,N_37017);
xor U37466 (N_37466,N_37179,N_37200);
and U37467 (N_37467,N_37028,N_37185);
and U37468 (N_37468,N_37132,N_37004);
and U37469 (N_37469,N_37179,N_37151);
xnor U37470 (N_37470,N_37041,N_37029);
xnor U37471 (N_37471,N_37041,N_37080);
and U37472 (N_37472,N_37095,N_37131);
nor U37473 (N_37473,N_37086,N_37165);
or U37474 (N_37474,N_37152,N_37167);
and U37475 (N_37475,N_37019,N_37168);
or U37476 (N_37476,N_37051,N_37001);
nor U37477 (N_37477,N_37015,N_37227);
and U37478 (N_37478,N_37127,N_37169);
nor U37479 (N_37479,N_37060,N_37237);
or U37480 (N_37480,N_37156,N_37047);
or U37481 (N_37481,N_37069,N_37059);
xnor U37482 (N_37482,N_37052,N_37029);
and U37483 (N_37483,N_37186,N_37190);
nand U37484 (N_37484,N_37152,N_37049);
or U37485 (N_37485,N_37103,N_37109);
and U37486 (N_37486,N_37237,N_37133);
xnor U37487 (N_37487,N_37241,N_37187);
nand U37488 (N_37488,N_37147,N_37174);
nor U37489 (N_37489,N_37041,N_37122);
nand U37490 (N_37490,N_37224,N_37165);
nand U37491 (N_37491,N_37047,N_37029);
xor U37492 (N_37492,N_37160,N_37013);
nand U37493 (N_37493,N_37133,N_37047);
xor U37494 (N_37494,N_37233,N_37193);
nor U37495 (N_37495,N_37223,N_37190);
xnor U37496 (N_37496,N_37035,N_37070);
nand U37497 (N_37497,N_37064,N_37097);
nor U37498 (N_37498,N_37004,N_37126);
and U37499 (N_37499,N_37216,N_37089);
and U37500 (N_37500,N_37399,N_37271);
nand U37501 (N_37501,N_37361,N_37485);
nor U37502 (N_37502,N_37265,N_37293);
or U37503 (N_37503,N_37490,N_37421);
or U37504 (N_37504,N_37251,N_37312);
or U37505 (N_37505,N_37376,N_37455);
xnor U37506 (N_37506,N_37306,N_37381);
xor U37507 (N_37507,N_37262,N_37428);
nand U37508 (N_37508,N_37266,N_37345);
nor U37509 (N_37509,N_37425,N_37420);
nor U37510 (N_37510,N_37462,N_37360);
or U37511 (N_37511,N_37260,N_37307);
xor U37512 (N_37512,N_37328,N_37364);
nand U37513 (N_37513,N_37458,N_37463);
or U37514 (N_37514,N_37253,N_37468);
nor U37515 (N_37515,N_37439,N_37349);
or U37516 (N_37516,N_37267,N_37337);
nor U37517 (N_37517,N_37286,N_37470);
nand U37518 (N_37518,N_37464,N_37344);
and U37519 (N_37519,N_37341,N_37448);
nor U37520 (N_37520,N_37302,N_37259);
and U37521 (N_37521,N_37409,N_37275);
nor U37522 (N_37522,N_37313,N_37291);
xnor U37523 (N_37523,N_37449,N_37352);
nand U37524 (N_37524,N_37412,N_37392);
nor U37525 (N_37525,N_37333,N_37445);
and U37526 (N_37526,N_37380,N_37467);
nand U37527 (N_37527,N_37287,N_37385);
nand U37528 (N_37528,N_37495,N_37438);
or U37529 (N_37529,N_37283,N_37367);
xnor U37530 (N_37530,N_37480,N_37303);
nor U37531 (N_37531,N_37358,N_37430);
nand U37532 (N_37532,N_37471,N_37432);
nand U37533 (N_37533,N_37365,N_37258);
nor U37534 (N_37534,N_37309,N_37459);
or U37535 (N_37535,N_37404,N_37279);
nand U37536 (N_37536,N_37378,N_37431);
or U37537 (N_37537,N_37408,N_37434);
xor U37538 (N_37538,N_37401,N_37478);
xnor U37539 (N_37539,N_37488,N_37387);
or U37540 (N_37540,N_37374,N_37450);
xor U37541 (N_37541,N_37294,N_37441);
nor U37542 (N_37542,N_37324,N_37362);
nand U37543 (N_37543,N_37422,N_37298);
nand U37544 (N_37544,N_37453,N_37405);
xor U37545 (N_37545,N_37496,N_37460);
nor U37546 (N_37546,N_37268,N_37413);
or U37547 (N_37547,N_37454,N_37386);
or U37548 (N_37548,N_37492,N_37284);
nor U37549 (N_37549,N_37280,N_37273);
nor U37550 (N_37550,N_37331,N_37311);
and U37551 (N_37551,N_37395,N_37411);
nand U37552 (N_37552,N_37288,N_37278);
or U37553 (N_37553,N_37444,N_37295);
nand U37554 (N_37554,N_37372,N_37274);
or U37555 (N_37555,N_37261,N_37406);
xor U37556 (N_37556,N_37499,N_37433);
xnor U37557 (N_37557,N_37343,N_37310);
xnor U37558 (N_37558,N_37415,N_37443);
and U37559 (N_37559,N_37410,N_37255);
nor U37560 (N_37560,N_37418,N_37263);
nor U37561 (N_37561,N_37322,N_37465);
nand U37562 (N_37562,N_37429,N_37289);
or U37563 (N_37563,N_37326,N_37327);
nand U37564 (N_37564,N_37350,N_37402);
or U37565 (N_37565,N_37250,N_37340);
nand U37566 (N_37566,N_37400,N_37417);
and U37567 (N_37567,N_37348,N_37325);
nand U37568 (N_37568,N_37272,N_37486);
nand U37569 (N_37569,N_37332,N_37476);
or U37570 (N_37570,N_37301,N_37384);
nor U37571 (N_37571,N_37423,N_37300);
and U37572 (N_37572,N_37456,N_37264);
and U37573 (N_37573,N_37317,N_37330);
or U37574 (N_37574,N_37357,N_37440);
nand U37575 (N_37575,N_37491,N_37282);
nand U37576 (N_37576,N_37403,N_37416);
nand U37577 (N_37577,N_37359,N_37355);
nor U37578 (N_37578,N_37369,N_37469);
xor U37579 (N_37579,N_37356,N_37335);
or U37580 (N_37580,N_37323,N_37479);
or U37581 (N_37581,N_37347,N_37393);
nand U37582 (N_37582,N_37474,N_37388);
xnor U37583 (N_37583,N_37375,N_37407);
nand U37584 (N_37584,N_37319,N_37320);
xor U37585 (N_37585,N_37382,N_37419);
or U37586 (N_37586,N_37316,N_37314);
nor U37587 (N_37587,N_37484,N_37397);
xor U37588 (N_37588,N_37398,N_37366);
nand U37589 (N_37589,N_37334,N_37477);
or U37590 (N_37590,N_37483,N_37472);
nand U37591 (N_37591,N_37368,N_37427);
xnor U37592 (N_37592,N_37497,N_37426);
xor U37593 (N_37593,N_37321,N_37457);
nand U37594 (N_37594,N_37481,N_37451);
and U37595 (N_37595,N_37493,N_37442);
nand U37596 (N_37596,N_37304,N_37342);
and U37597 (N_37597,N_37383,N_37329);
nor U37598 (N_37598,N_37414,N_37487);
or U37599 (N_37599,N_37257,N_37270);
xor U37600 (N_37600,N_37498,N_37363);
and U37601 (N_37601,N_37461,N_37285);
xor U37602 (N_37602,N_37276,N_37292);
or U37603 (N_37603,N_37308,N_37290);
nand U37604 (N_37604,N_37299,N_37339);
and U37605 (N_37605,N_37424,N_37338);
and U37606 (N_37606,N_37353,N_37254);
nor U37607 (N_37607,N_37305,N_37482);
and U37608 (N_37608,N_37394,N_37466);
and U37609 (N_37609,N_37281,N_37297);
nand U37610 (N_37610,N_37336,N_37315);
or U37611 (N_37611,N_37377,N_37447);
xor U37612 (N_37612,N_37277,N_37370);
and U37613 (N_37613,N_37446,N_37256);
nand U37614 (N_37614,N_37354,N_37473);
nor U37615 (N_37615,N_37346,N_37252);
and U37616 (N_37616,N_37452,N_37296);
or U37617 (N_37617,N_37373,N_37318);
nand U37618 (N_37618,N_37489,N_37475);
xnor U37619 (N_37619,N_37435,N_37269);
nand U37620 (N_37620,N_37391,N_37371);
and U37621 (N_37621,N_37436,N_37494);
or U37622 (N_37622,N_37437,N_37390);
nand U37623 (N_37623,N_37351,N_37379);
or U37624 (N_37624,N_37389,N_37396);
or U37625 (N_37625,N_37399,N_37329);
nor U37626 (N_37626,N_37386,N_37351);
or U37627 (N_37627,N_37470,N_37478);
nand U37628 (N_37628,N_37487,N_37444);
or U37629 (N_37629,N_37442,N_37285);
nor U37630 (N_37630,N_37287,N_37485);
xnor U37631 (N_37631,N_37438,N_37443);
nor U37632 (N_37632,N_37414,N_37266);
and U37633 (N_37633,N_37482,N_37326);
xnor U37634 (N_37634,N_37480,N_37420);
nand U37635 (N_37635,N_37290,N_37276);
and U37636 (N_37636,N_37437,N_37272);
xor U37637 (N_37637,N_37259,N_37497);
or U37638 (N_37638,N_37288,N_37355);
or U37639 (N_37639,N_37415,N_37399);
xor U37640 (N_37640,N_37277,N_37293);
xnor U37641 (N_37641,N_37267,N_37475);
xor U37642 (N_37642,N_37475,N_37304);
and U37643 (N_37643,N_37465,N_37319);
nand U37644 (N_37644,N_37293,N_37458);
xor U37645 (N_37645,N_37373,N_37456);
and U37646 (N_37646,N_37252,N_37364);
or U37647 (N_37647,N_37332,N_37326);
and U37648 (N_37648,N_37444,N_37310);
nand U37649 (N_37649,N_37268,N_37363);
xor U37650 (N_37650,N_37357,N_37310);
xnor U37651 (N_37651,N_37408,N_37460);
and U37652 (N_37652,N_37319,N_37334);
and U37653 (N_37653,N_37486,N_37433);
or U37654 (N_37654,N_37337,N_37288);
nand U37655 (N_37655,N_37369,N_37427);
nand U37656 (N_37656,N_37273,N_37481);
or U37657 (N_37657,N_37492,N_37384);
or U37658 (N_37658,N_37357,N_37400);
or U37659 (N_37659,N_37395,N_37254);
xor U37660 (N_37660,N_37255,N_37493);
and U37661 (N_37661,N_37474,N_37356);
nor U37662 (N_37662,N_37351,N_37262);
xor U37663 (N_37663,N_37398,N_37273);
nor U37664 (N_37664,N_37353,N_37460);
nand U37665 (N_37665,N_37284,N_37306);
or U37666 (N_37666,N_37261,N_37327);
or U37667 (N_37667,N_37334,N_37383);
nor U37668 (N_37668,N_37383,N_37361);
or U37669 (N_37669,N_37252,N_37390);
or U37670 (N_37670,N_37428,N_37342);
or U37671 (N_37671,N_37367,N_37454);
and U37672 (N_37672,N_37342,N_37459);
xnor U37673 (N_37673,N_37416,N_37324);
nand U37674 (N_37674,N_37351,N_37391);
nor U37675 (N_37675,N_37424,N_37400);
or U37676 (N_37676,N_37360,N_37322);
nand U37677 (N_37677,N_37294,N_37359);
and U37678 (N_37678,N_37416,N_37369);
or U37679 (N_37679,N_37473,N_37441);
xnor U37680 (N_37680,N_37481,N_37408);
and U37681 (N_37681,N_37336,N_37414);
xnor U37682 (N_37682,N_37255,N_37271);
nor U37683 (N_37683,N_37436,N_37382);
nand U37684 (N_37684,N_37319,N_37296);
or U37685 (N_37685,N_37282,N_37354);
or U37686 (N_37686,N_37434,N_37258);
xnor U37687 (N_37687,N_37409,N_37386);
nor U37688 (N_37688,N_37402,N_37428);
nor U37689 (N_37689,N_37434,N_37498);
nand U37690 (N_37690,N_37258,N_37426);
xor U37691 (N_37691,N_37353,N_37395);
nand U37692 (N_37692,N_37455,N_37280);
nor U37693 (N_37693,N_37421,N_37403);
nand U37694 (N_37694,N_37366,N_37474);
nor U37695 (N_37695,N_37278,N_37343);
or U37696 (N_37696,N_37458,N_37291);
nand U37697 (N_37697,N_37393,N_37472);
xor U37698 (N_37698,N_37398,N_37328);
xor U37699 (N_37699,N_37363,N_37467);
xnor U37700 (N_37700,N_37279,N_37497);
nand U37701 (N_37701,N_37262,N_37364);
nor U37702 (N_37702,N_37372,N_37436);
and U37703 (N_37703,N_37368,N_37439);
nor U37704 (N_37704,N_37478,N_37311);
or U37705 (N_37705,N_37339,N_37250);
or U37706 (N_37706,N_37476,N_37452);
or U37707 (N_37707,N_37400,N_37401);
nor U37708 (N_37708,N_37267,N_37278);
nand U37709 (N_37709,N_37313,N_37309);
or U37710 (N_37710,N_37314,N_37392);
nor U37711 (N_37711,N_37273,N_37456);
nand U37712 (N_37712,N_37372,N_37307);
nor U37713 (N_37713,N_37372,N_37269);
and U37714 (N_37714,N_37277,N_37416);
xnor U37715 (N_37715,N_37320,N_37400);
nor U37716 (N_37716,N_37299,N_37271);
nor U37717 (N_37717,N_37486,N_37449);
nand U37718 (N_37718,N_37281,N_37293);
nor U37719 (N_37719,N_37373,N_37262);
nor U37720 (N_37720,N_37429,N_37456);
nor U37721 (N_37721,N_37375,N_37452);
xnor U37722 (N_37722,N_37404,N_37485);
nand U37723 (N_37723,N_37482,N_37477);
or U37724 (N_37724,N_37459,N_37433);
xnor U37725 (N_37725,N_37281,N_37336);
and U37726 (N_37726,N_37488,N_37489);
and U37727 (N_37727,N_37320,N_37338);
or U37728 (N_37728,N_37383,N_37399);
nor U37729 (N_37729,N_37490,N_37492);
nor U37730 (N_37730,N_37479,N_37456);
or U37731 (N_37731,N_37342,N_37439);
nor U37732 (N_37732,N_37368,N_37261);
or U37733 (N_37733,N_37336,N_37438);
nand U37734 (N_37734,N_37454,N_37340);
xor U37735 (N_37735,N_37378,N_37408);
nand U37736 (N_37736,N_37385,N_37320);
xor U37737 (N_37737,N_37341,N_37483);
nor U37738 (N_37738,N_37363,N_37453);
and U37739 (N_37739,N_37366,N_37346);
xnor U37740 (N_37740,N_37300,N_37324);
nor U37741 (N_37741,N_37329,N_37303);
nand U37742 (N_37742,N_37324,N_37260);
and U37743 (N_37743,N_37398,N_37443);
or U37744 (N_37744,N_37336,N_37349);
or U37745 (N_37745,N_37459,N_37460);
nor U37746 (N_37746,N_37428,N_37258);
xnor U37747 (N_37747,N_37477,N_37496);
nand U37748 (N_37748,N_37472,N_37428);
and U37749 (N_37749,N_37370,N_37284);
nand U37750 (N_37750,N_37731,N_37590);
or U37751 (N_37751,N_37745,N_37527);
and U37752 (N_37752,N_37507,N_37649);
and U37753 (N_37753,N_37732,N_37515);
xnor U37754 (N_37754,N_37501,N_37603);
and U37755 (N_37755,N_37576,N_37529);
nor U37756 (N_37756,N_37674,N_37504);
nor U37757 (N_37757,N_37516,N_37610);
nand U37758 (N_37758,N_37729,N_37716);
and U37759 (N_37759,N_37690,N_37718);
and U37760 (N_37760,N_37606,N_37564);
or U37761 (N_37761,N_37531,N_37678);
xnor U37762 (N_37762,N_37633,N_37518);
and U37763 (N_37763,N_37626,N_37644);
and U37764 (N_37764,N_37503,N_37715);
or U37765 (N_37765,N_37701,N_37592);
nor U37766 (N_37766,N_37702,N_37523);
nand U37767 (N_37767,N_37589,N_37735);
or U37768 (N_37768,N_37643,N_37567);
nor U37769 (N_37769,N_37550,N_37645);
nor U37770 (N_37770,N_37709,N_37647);
xnor U37771 (N_37771,N_37585,N_37505);
xnor U37772 (N_37772,N_37604,N_37598);
nand U37773 (N_37773,N_37650,N_37570);
nor U37774 (N_37774,N_37584,N_37586);
nor U37775 (N_37775,N_37662,N_37736);
and U37776 (N_37776,N_37526,N_37713);
or U37777 (N_37777,N_37595,N_37582);
nand U37778 (N_37778,N_37688,N_37692);
xnor U37779 (N_37779,N_37656,N_37636);
nand U37780 (N_37780,N_37664,N_37661);
nand U37781 (N_37781,N_37545,N_37737);
xnor U37782 (N_37782,N_37700,N_37723);
nor U37783 (N_37783,N_37660,N_37691);
or U37784 (N_37784,N_37614,N_37539);
nor U37785 (N_37785,N_37743,N_37521);
and U37786 (N_37786,N_37547,N_37632);
nand U37787 (N_37787,N_37724,N_37608);
nand U37788 (N_37788,N_37548,N_37683);
nor U37789 (N_37789,N_37573,N_37609);
nand U37790 (N_37790,N_37658,N_37581);
nand U37791 (N_37791,N_37601,N_37525);
or U37792 (N_37792,N_37714,N_37634);
or U37793 (N_37793,N_37741,N_37607);
nand U37794 (N_37794,N_37568,N_37558);
and U37795 (N_37795,N_37559,N_37659);
xor U37796 (N_37796,N_37680,N_37617);
nand U37797 (N_37797,N_37642,N_37588);
nor U37798 (N_37798,N_37749,N_37596);
and U37799 (N_37799,N_37733,N_37562);
xnor U37800 (N_37800,N_37635,N_37599);
or U37801 (N_37801,N_37734,N_37639);
xor U37802 (N_37802,N_37679,N_37646);
and U37803 (N_37803,N_37566,N_37571);
and U37804 (N_37804,N_37513,N_37502);
and U37805 (N_37805,N_37542,N_37726);
or U37806 (N_37806,N_37528,N_37676);
and U37807 (N_37807,N_37675,N_37696);
xor U37808 (N_37808,N_37560,N_37579);
nand U37809 (N_37809,N_37623,N_37728);
xor U37810 (N_37810,N_37673,N_37685);
nand U37811 (N_37811,N_37651,N_37549);
nor U37812 (N_37812,N_37706,N_37552);
nand U37813 (N_37813,N_37511,N_37725);
or U37814 (N_37814,N_37671,N_37727);
nor U37815 (N_37815,N_37618,N_37537);
or U37816 (N_37816,N_37538,N_37575);
or U37817 (N_37817,N_37708,N_37668);
and U37818 (N_37818,N_37605,N_37583);
and U37819 (N_37819,N_37697,N_37682);
nor U37820 (N_37820,N_37543,N_37695);
nand U37821 (N_37821,N_37533,N_37517);
nand U37822 (N_37822,N_37613,N_37730);
or U37823 (N_37823,N_37594,N_37655);
nand U37824 (N_37824,N_37637,N_37654);
nand U37825 (N_37825,N_37554,N_37693);
and U37826 (N_37826,N_37593,N_37616);
or U37827 (N_37827,N_37711,N_37530);
or U37828 (N_37828,N_37563,N_37556);
and U37829 (N_37829,N_37565,N_37541);
nor U37830 (N_37830,N_37506,N_37689);
xor U37831 (N_37831,N_37739,N_37630);
and U37832 (N_37832,N_37519,N_37524);
nand U37833 (N_37833,N_37648,N_37686);
nor U37834 (N_37834,N_37687,N_37710);
or U37835 (N_37835,N_37699,N_37602);
nand U37836 (N_37836,N_37587,N_37705);
or U37837 (N_37837,N_37600,N_37667);
nand U37838 (N_37838,N_37712,N_37665);
nand U37839 (N_37839,N_37669,N_37744);
xnor U37840 (N_37840,N_37627,N_37572);
and U37841 (N_37841,N_37628,N_37738);
and U37842 (N_37842,N_37532,N_37622);
or U37843 (N_37843,N_37569,N_37707);
xor U37844 (N_37844,N_37694,N_37551);
xor U37845 (N_37845,N_37717,N_37631);
or U37846 (N_37846,N_37536,N_37722);
nand U37847 (N_37847,N_37684,N_37578);
or U37848 (N_37848,N_37509,N_37553);
nor U37849 (N_37849,N_37672,N_37640);
nor U37850 (N_37850,N_37580,N_37720);
or U37851 (N_37851,N_37619,N_37577);
nand U37852 (N_37852,N_37719,N_37520);
nand U37853 (N_37853,N_37522,N_37747);
and U37854 (N_37854,N_37611,N_37670);
nor U37855 (N_37855,N_37698,N_37663);
or U37856 (N_37856,N_37591,N_37508);
nor U37857 (N_37857,N_37677,N_37703);
or U37858 (N_37858,N_37657,N_37510);
or U37859 (N_37859,N_37561,N_37555);
or U37860 (N_37860,N_37641,N_37512);
or U37861 (N_37861,N_37625,N_37544);
xor U37862 (N_37862,N_37540,N_37534);
nor U37863 (N_37863,N_37704,N_37546);
nand U37864 (N_37864,N_37535,N_37621);
xnor U37865 (N_37865,N_37742,N_37721);
or U37866 (N_37866,N_37748,N_37615);
and U37867 (N_37867,N_37620,N_37597);
nand U37868 (N_37868,N_37653,N_37681);
nor U37869 (N_37869,N_37740,N_37612);
xor U37870 (N_37870,N_37666,N_37500);
and U37871 (N_37871,N_37652,N_37574);
xor U37872 (N_37872,N_37746,N_37624);
and U37873 (N_37873,N_37557,N_37638);
or U37874 (N_37874,N_37514,N_37629);
xor U37875 (N_37875,N_37533,N_37651);
and U37876 (N_37876,N_37673,N_37709);
and U37877 (N_37877,N_37590,N_37650);
nor U37878 (N_37878,N_37642,N_37592);
nor U37879 (N_37879,N_37520,N_37716);
and U37880 (N_37880,N_37542,N_37623);
or U37881 (N_37881,N_37701,N_37575);
xor U37882 (N_37882,N_37703,N_37506);
and U37883 (N_37883,N_37559,N_37670);
nand U37884 (N_37884,N_37643,N_37502);
xor U37885 (N_37885,N_37642,N_37614);
nor U37886 (N_37886,N_37644,N_37659);
nor U37887 (N_37887,N_37585,N_37521);
xor U37888 (N_37888,N_37690,N_37553);
nand U37889 (N_37889,N_37546,N_37621);
nand U37890 (N_37890,N_37575,N_37744);
nand U37891 (N_37891,N_37705,N_37744);
xor U37892 (N_37892,N_37626,N_37593);
xor U37893 (N_37893,N_37500,N_37630);
xor U37894 (N_37894,N_37562,N_37594);
and U37895 (N_37895,N_37586,N_37578);
nand U37896 (N_37896,N_37577,N_37546);
xnor U37897 (N_37897,N_37670,N_37570);
or U37898 (N_37898,N_37587,N_37547);
nand U37899 (N_37899,N_37540,N_37554);
nor U37900 (N_37900,N_37609,N_37713);
and U37901 (N_37901,N_37581,N_37537);
and U37902 (N_37902,N_37591,N_37659);
and U37903 (N_37903,N_37653,N_37537);
nor U37904 (N_37904,N_37637,N_37666);
and U37905 (N_37905,N_37650,N_37716);
nor U37906 (N_37906,N_37609,N_37508);
xnor U37907 (N_37907,N_37658,N_37615);
or U37908 (N_37908,N_37602,N_37704);
xor U37909 (N_37909,N_37673,N_37738);
and U37910 (N_37910,N_37629,N_37509);
or U37911 (N_37911,N_37555,N_37571);
and U37912 (N_37912,N_37646,N_37704);
nor U37913 (N_37913,N_37556,N_37626);
xnor U37914 (N_37914,N_37720,N_37503);
and U37915 (N_37915,N_37718,N_37647);
and U37916 (N_37916,N_37567,N_37610);
and U37917 (N_37917,N_37706,N_37610);
and U37918 (N_37918,N_37611,N_37505);
nand U37919 (N_37919,N_37724,N_37702);
nand U37920 (N_37920,N_37714,N_37669);
nand U37921 (N_37921,N_37679,N_37737);
and U37922 (N_37922,N_37664,N_37674);
or U37923 (N_37923,N_37729,N_37723);
or U37924 (N_37924,N_37682,N_37653);
and U37925 (N_37925,N_37677,N_37747);
or U37926 (N_37926,N_37540,N_37661);
and U37927 (N_37927,N_37602,N_37724);
nor U37928 (N_37928,N_37569,N_37719);
xnor U37929 (N_37929,N_37706,N_37646);
nor U37930 (N_37930,N_37732,N_37563);
nor U37931 (N_37931,N_37669,N_37538);
xnor U37932 (N_37932,N_37519,N_37670);
xor U37933 (N_37933,N_37725,N_37729);
nand U37934 (N_37934,N_37672,N_37737);
and U37935 (N_37935,N_37626,N_37611);
and U37936 (N_37936,N_37607,N_37551);
xnor U37937 (N_37937,N_37644,N_37708);
xor U37938 (N_37938,N_37704,N_37595);
or U37939 (N_37939,N_37664,N_37728);
nand U37940 (N_37940,N_37516,N_37604);
xnor U37941 (N_37941,N_37563,N_37539);
xnor U37942 (N_37942,N_37707,N_37691);
nand U37943 (N_37943,N_37539,N_37611);
nor U37944 (N_37944,N_37717,N_37508);
nor U37945 (N_37945,N_37731,N_37721);
and U37946 (N_37946,N_37599,N_37678);
nand U37947 (N_37947,N_37701,N_37742);
xnor U37948 (N_37948,N_37517,N_37512);
nor U37949 (N_37949,N_37698,N_37667);
or U37950 (N_37950,N_37673,N_37714);
nand U37951 (N_37951,N_37609,N_37720);
and U37952 (N_37952,N_37636,N_37540);
nand U37953 (N_37953,N_37533,N_37732);
nand U37954 (N_37954,N_37613,N_37573);
xor U37955 (N_37955,N_37683,N_37568);
or U37956 (N_37956,N_37619,N_37712);
nand U37957 (N_37957,N_37608,N_37557);
nor U37958 (N_37958,N_37562,N_37568);
and U37959 (N_37959,N_37663,N_37693);
nand U37960 (N_37960,N_37682,N_37597);
xor U37961 (N_37961,N_37736,N_37585);
nor U37962 (N_37962,N_37544,N_37602);
xnor U37963 (N_37963,N_37736,N_37722);
xor U37964 (N_37964,N_37703,N_37575);
or U37965 (N_37965,N_37580,N_37544);
nor U37966 (N_37966,N_37720,N_37585);
xor U37967 (N_37967,N_37673,N_37674);
or U37968 (N_37968,N_37575,N_37600);
xor U37969 (N_37969,N_37640,N_37511);
xor U37970 (N_37970,N_37500,N_37651);
or U37971 (N_37971,N_37514,N_37650);
or U37972 (N_37972,N_37531,N_37523);
or U37973 (N_37973,N_37606,N_37698);
nor U37974 (N_37974,N_37530,N_37695);
or U37975 (N_37975,N_37624,N_37562);
or U37976 (N_37976,N_37536,N_37539);
or U37977 (N_37977,N_37621,N_37612);
and U37978 (N_37978,N_37536,N_37746);
nand U37979 (N_37979,N_37616,N_37720);
nor U37980 (N_37980,N_37610,N_37561);
or U37981 (N_37981,N_37724,N_37607);
or U37982 (N_37982,N_37622,N_37726);
nand U37983 (N_37983,N_37574,N_37533);
nor U37984 (N_37984,N_37672,N_37517);
and U37985 (N_37985,N_37654,N_37687);
or U37986 (N_37986,N_37731,N_37598);
nor U37987 (N_37987,N_37580,N_37582);
nand U37988 (N_37988,N_37514,N_37533);
nor U37989 (N_37989,N_37630,N_37689);
nor U37990 (N_37990,N_37684,N_37727);
or U37991 (N_37991,N_37512,N_37652);
nand U37992 (N_37992,N_37684,N_37731);
xnor U37993 (N_37993,N_37594,N_37733);
xnor U37994 (N_37994,N_37569,N_37723);
nor U37995 (N_37995,N_37579,N_37702);
nor U37996 (N_37996,N_37502,N_37628);
xor U37997 (N_37997,N_37617,N_37519);
nor U37998 (N_37998,N_37614,N_37682);
or U37999 (N_37999,N_37572,N_37593);
xor U38000 (N_38000,N_37879,N_37789);
nor U38001 (N_38001,N_37781,N_37853);
nor U38002 (N_38002,N_37965,N_37855);
nand U38003 (N_38003,N_37783,N_37984);
nand U38004 (N_38004,N_37755,N_37894);
nand U38005 (N_38005,N_37768,N_37951);
nor U38006 (N_38006,N_37887,N_37839);
nand U38007 (N_38007,N_37901,N_37943);
nor U38008 (N_38008,N_37766,N_37751);
xnor U38009 (N_38009,N_37764,N_37888);
and U38010 (N_38010,N_37752,N_37865);
and U38011 (N_38011,N_37880,N_37905);
or U38012 (N_38012,N_37762,N_37979);
or U38013 (N_38013,N_37818,N_37904);
nand U38014 (N_38014,N_37833,N_37957);
xor U38015 (N_38015,N_37961,N_37930);
and U38016 (N_38016,N_37932,N_37948);
and U38017 (N_38017,N_37936,N_37843);
nand U38018 (N_38018,N_37829,N_37805);
and U38019 (N_38019,N_37836,N_37980);
nor U38020 (N_38020,N_37872,N_37852);
or U38021 (N_38021,N_37759,N_37810);
and U38022 (N_38022,N_37862,N_37777);
xnor U38023 (N_38023,N_37982,N_37999);
nand U38024 (N_38024,N_37858,N_37846);
nor U38025 (N_38025,N_37763,N_37920);
nand U38026 (N_38026,N_37840,N_37842);
nor U38027 (N_38027,N_37797,N_37791);
xnor U38028 (N_38028,N_37922,N_37754);
nand U38029 (N_38029,N_37778,N_37983);
xnor U38030 (N_38030,N_37807,N_37849);
and U38031 (N_38031,N_37854,N_37861);
and U38032 (N_38032,N_37919,N_37821);
nand U38033 (N_38033,N_37776,N_37947);
or U38034 (N_38034,N_37893,N_37954);
and U38035 (N_38035,N_37803,N_37851);
nor U38036 (N_38036,N_37952,N_37760);
nand U38037 (N_38037,N_37816,N_37761);
and U38038 (N_38038,N_37859,N_37820);
or U38039 (N_38039,N_37917,N_37796);
nand U38040 (N_38040,N_37799,N_37991);
nor U38041 (N_38041,N_37973,N_37966);
and U38042 (N_38042,N_37873,N_37771);
or U38043 (N_38043,N_37924,N_37918);
xnor U38044 (N_38044,N_37911,N_37995);
nor U38045 (N_38045,N_37906,N_37969);
or U38046 (N_38046,N_37756,N_37934);
or U38047 (N_38047,N_37875,N_37998);
and U38048 (N_38048,N_37750,N_37903);
nand U38049 (N_38049,N_37800,N_37925);
nand U38050 (N_38050,N_37914,N_37889);
or U38051 (N_38051,N_37856,N_37882);
xnor U38052 (N_38052,N_37886,N_37898);
and U38053 (N_38053,N_37775,N_37909);
nand U38054 (N_38054,N_37784,N_37967);
nand U38055 (N_38055,N_37923,N_37900);
nor U38056 (N_38056,N_37971,N_37990);
or U38057 (N_38057,N_37860,N_37790);
nand U38058 (N_38058,N_37956,N_37928);
nand U38059 (N_38059,N_37753,N_37835);
and U38060 (N_38060,N_37896,N_37832);
nand U38061 (N_38061,N_37828,N_37757);
or U38062 (N_38062,N_37804,N_37989);
xnor U38063 (N_38063,N_37985,N_37935);
xnor U38064 (N_38064,N_37826,N_37857);
xor U38065 (N_38065,N_37831,N_37892);
nand U38066 (N_38066,N_37782,N_37808);
nand U38067 (N_38067,N_37926,N_37823);
nand U38068 (N_38068,N_37822,N_37838);
or U38069 (N_38069,N_37815,N_37812);
or U38070 (N_38070,N_37830,N_37950);
nor U38071 (N_38071,N_37975,N_37787);
nand U38072 (N_38072,N_37793,N_37878);
xnor U38073 (N_38073,N_37987,N_37963);
and U38074 (N_38074,N_37848,N_37921);
nor U38075 (N_38075,N_37899,N_37931);
nand U38076 (N_38076,N_37976,N_37769);
nand U38077 (N_38077,N_37758,N_37780);
nand U38078 (N_38078,N_37994,N_37978);
xor U38079 (N_38079,N_37960,N_37847);
nand U38080 (N_38080,N_37958,N_37817);
nand U38081 (N_38081,N_37949,N_37874);
or U38082 (N_38082,N_37927,N_37915);
xnor U38083 (N_38083,N_37912,N_37794);
or U38084 (N_38084,N_37929,N_37814);
nand U38085 (N_38085,N_37850,N_37933);
xor U38086 (N_38086,N_37938,N_37902);
xor U38087 (N_38087,N_37767,N_37869);
nand U38088 (N_38088,N_37916,N_37992);
nor U38089 (N_38089,N_37786,N_37939);
xnor U38090 (N_38090,N_37942,N_37970);
or U38091 (N_38091,N_37773,N_37795);
xor U38092 (N_38092,N_37827,N_37981);
nor U38093 (N_38093,N_37968,N_37913);
xor U38094 (N_38094,N_37945,N_37964);
and U38095 (N_38095,N_37877,N_37774);
nand U38096 (N_38096,N_37824,N_37883);
nor U38097 (N_38097,N_37863,N_37955);
xor U38098 (N_38098,N_37798,N_37802);
or U38099 (N_38099,N_37772,N_37868);
nand U38100 (N_38100,N_37811,N_37834);
xor U38101 (N_38101,N_37876,N_37837);
nor U38102 (N_38102,N_37907,N_37908);
nor U38103 (N_38103,N_37910,N_37792);
xor U38104 (N_38104,N_37785,N_37940);
or U38105 (N_38105,N_37996,N_37825);
or U38106 (N_38106,N_37806,N_37809);
and U38107 (N_38107,N_37801,N_37977);
or U38108 (N_38108,N_37986,N_37770);
nand U38109 (N_38109,N_37988,N_37891);
or U38110 (N_38110,N_37813,N_37819);
nand U38111 (N_38111,N_37946,N_37867);
and U38112 (N_38112,N_37974,N_37890);
nor U38113 (N_38113,N_37884,N_37953);
xnor U38114 (N_38114,N_37871,N_37895);
or U38115 (N_38115,N_37962,N_37885);
or U38116 (N_38116,N_37937,N_37870);
xnor U38117 (N_38117,N_37944,N_37897);
and U38118 (N_38118,N_37972,N_37866);
xnor U38119 (N_38119,N_37765,N_37788);
xor U38120 (N_38120,N_37841,N_37993);
nor U38121 (N_38121,N_37881,N_37997);
nand U38122 (N_38122,N_37845,N_37779);
nand U38123 (N_38123,N_37941,N_37864);
nand U38124 (N_38124,N_37844,N_37959);
xor U38125 (N_38125,N_37987,N_37761);
nor U38126 (N_38126,N_37894,N_37774);
and U38127 (N_38127,N_37935,N_37955);
and U38128 (N_38128,N_37940,N_37863);
nand U38129 (N_38129,N_37862,N_37886);
xnor U38130 (N_38130,N_37861,N_37930);
or U38131 (N_38131,N_37780,N_37982);
nor U38132 (N_38132,N_37765,N_37953);
and U38133 (N_38133,N_37801,N_37966);
nand U38134 (N_38134,N_37949,N_37885);
nand U38135 (N_38135,N_37970,N_37901);
xnor U38136 (N_38136,N_37918,N_37942);
xnor U38137 (N_38137,N_37941,N_37937);
xnor U38138 (N_38138,N_37931,N_37813);
nor U38139 (N_38139,N_37897,N_37814);
xnor U38140 (N_38140,N_37849,N_37786);
nand U38141 (N_38141,N_37851,N_37891);
nor U38142 (N_38142,N_37946,N_37756);
or U38143 (N_38143,N_37757,N_37980);
nand U38144 (N_38144,N_37848,N_37813);
or U38145 (N_38145,N_37874,N_37758);
xnor U38146 (N_38146,N_37835,N_37907);
nor U38147 (N_38147,N_37777,N_37864);
nor U38148 (N_38148,N_37876,N_37890);
or U38149 (N_38149,N_37753,N_37829);
nor U38150 (N_38150,N_37819,N_37783);
or U38151 (N_38151,N_37929,N_37796);
nand U38152 (N_38152,N_37988,N_37975);
and U38153 (N_38153,N_37930,N_37791);
nand U38154 (N_38154,N_37859,N_37883);
and U38155 (N_38155,N_37993,N_37758);
and U38156 (N_38156,N_37883,N_37752);
xor U38157 (N_38157,N_37932,N_37772);
xnor U38158 (N_38158,N_37781,N_37838);
xor U38159 (N_38159,N_37945,N_37825);
nand U38160 (N_38160,N_37809,N_37852);
xnor U38161 (N_38161,N_37786,N_37913);
xnor U38162 (N_38162,N_37936,N_37878);
nor U38163 (N_38163,N_37897,N_37978);
nand U38164 (N_38164,N_37757,N_37764);
nor U38165 (N_38165,N_37975,N_37981);
and U38166 (N_38166,N_37965,N_37920);
nor U38167 (N_38167,N_37888,N_37825);
or U38168 (N_38168,N_37965,N_37882);
or U38169 (N_38169,N_37875,N_37957);
nand U38170 (N_38170,N_37968,N_37870);
nor U38171 (N_38171,N_37802,N_37838);
and U38172 (N_38172,N_37953,N_37986);
and U38173 (N_38173,N_37997,N_37782);
and U38174 (N_38174,N_37765,N_37858);
nand U38175 (N_38175,N_37765,N_37922);
nor U38176 (N_38176,N_37797,N_37960);
or U38177 (N_38177,N_37876,N_37946);
nor U38178 (N_38178,N_37861,N_37796);
nand U38179 (N_38179,N_37881,N_37873);
or U38180 (N_38180,N_37970,N_37991);
and U38181 (N_38181,N_37754,N_37988);
and U38182 (N_38182,N_37951,N_37935);
xor U38183 (N_38183,N_37935,N_37989);
and U38184 (N_38184,N_37946,N_37917);
or U38185 (N_38185,N_37940,N_37886);
nand U38186 (N_38186,N_37852,N_37991);
xnor U38187 (N_38187,N_37840,N_37847);
or U38188 (N_38188,N_37907,N_37803);
nor U38189 (N_38189,N_37920,N_37810);
and U38190 (N_38190,N_37805,N_37898);
nor U38191 (N_38191,N_37842,N_37789);
nor U38192 (N_38192,N_37829,N_37789);
xor U38193 (N_38193,N_37823,N_37800);
xor U38194 (N_38194,N_37874,N_37939);
and U38195 (N_38195,N_37873,N_37784);
nand U38196 (N_38196,N_37821,N_37932);
nand U38197 (N_38197,N_37964,N_37831);
and U38198 (N_38198,N_37786,N_37953);
nand U38199 (N_38199,N_37949,N_37944);
nor U38200 (N_38200,N_37945,N_37778);
nor U38201 (N_38201,N_37806,N_37838);
or U38202 (N_38202,N_37988,N_37893);
nand U38203 (N_38203,N_37883,N_37849);
or U38204 (N_38204,N_37895,N_37958);
xor U38205 (N_38205,N_37777,N_37916);
or U38206 (N_38206,N_37865,N_37789);
xor U38207 (N_38207,N_37792,N_37771);
nand U38208 (N_38208,N_37755,N_37939);
and U38209 (N_38209,N_37881,N_37796);
nor U38210 (N_38210,N_37981,N_37822);
nand U38211 (N_38211,N_37909,N_37965);
nand U38212 (N_38212,N_37750,N_37763);
or U38213 (N_38213,N_37787,N_37885);
nand U38214 (N_38214,N_37850,N_37895);
nand U38215 (N_38215,N_37799,N_37903);
xnor U38216 (N_38216,N_37775,N_37760);
and U38217 (N_38217,N_37904,N_37817);
and U38218 (N_38218,N_37900,N_37974);
nor U38219 (N_38219,N_37909,N_37830);
xnor U38220 (N_38220,N_37991,N_37905);
xor U38221 (N_38221,N_37765,N_37960);
and U38222 (N_38222,N_37923,N_37757);
xnor U38223 (N_38223,N_37966,N_37877);
nand U38224 (N_38224,N_37962,N_37961);
nor U38225 (N_38225,N_37772,N_37848);
nand U38226 (N_38226,N_37872,N_37767);
nor U38227 (N_38227,N_37769,N_37940);
nor U38228 (N_38228,N_37957,N_37819);
and U38229 (N_38229,N_37995,N_37993);
xnor U38230 (N_38230,N_37866,N_37872);
nor U38231 (N_38231,N_37971,N_37882);
or U38232 (N_38232,N_37767,N_37979);
nand U38233 (N_38233,N_37845,N_37905);
xnor U38234 (N_38234,N_37787,N_37921);
nor U38235 (N_38235,N_37768,N_37849);
nor U38236 (N_38236,N_37879,N_37934);
xor U38237 (N_38237,N_37798,N_37979);
nand U38238 (N_38238,N_37935,N_37798);
and U38239 (N_38239,N_37913,N_37932);
or U38240 (N_38240,N_37796,N_37914);
and U38241 (N_38241,N_37884,N_37830);
nor U38242 (N_38242,N_37964,N_37979);
or U38243 (N_38243,N_37997,N_37870);
and U38244 (N_38244,N_37865,N_37807);
nor U38245 (N_38245,N_37761,N_37829);
and U38246 (N_38246,N_37854,N_37843);
and U38247 (N_38247,N_37958,N_37778);
and U38248 (N_38248,N_37796,N_37916);
and U38249 (N_38249,N_37768,N_37883);
and U38250 (N_38250,N_38072,N_38002);
xor U38251 (N_38251,N_38070,N_38196);
xnor U38252 (N_38252,N_38159,N_38135);
or U38253 (N_38253,N_38049,N_38248);
and U38254 (N_38254,N_38079,N_38130);
nor U38255 (N_38255,N_38191,N_38077);
and U38256 (N_38256,N_38198,N_38028);
or U38257 (N_38257,N_38056,N_38004);
nand U38258 (N_38258,N_38085,N_38188);
and U38259 (N_38259,N_38060,N_38101);
or U38260 (N_38260,N_38010,N_38224);
or U38261 (N_38261,N_38216,N_38244);
nand U38262 (N_38262,N_38136,N_38182);
nand U38263 (N_38263,N_38051,N_38104);
xor U38264 (N_38264,N_38048,N_38126);
or U38265 (N_38265,N_38016,N_38213);
xnor U38266 (N_38266,N_38151,N_38155);
or U38267 (N_38267,N_38209,N_38128);
and U38268 (N_38268,N_38089,N_38084);
and U38269 (N_38269,N_38146,N_38121);
nand U38270 (N_38270,N_38001,N_38082);
nand U38271 (N_38271,N_38220,N_38117);
nand U38272 (N_38272,N_38204,N_38222);
or U38273 (N_38273,N_38205,N_38176);
or U38274 (N_38274,N_38074,N_38083);
nor U38275 (N_38275,N_38186,N_38158);
xor U38276 (N_38276,N_38228,N_38239);
nor U38277 (N_38277,N_38113,N_38131);
and U38278 (N_38278,N_38240,N_38147);
and U38279 (N_38279,N_38177,N_38125);
nor U38280 (N_38280,N_38039,N_38210);
nand U38281 (N_38281,N_38208,N_38179);
nor U38282 (N_38282,N_38093,N_38184);
or U38283 (N_38283,N_38118,N_38026);
xnor U38284 (N_38284,N_38092,N_38054);
xor U38285 (N_38285,N_38238,N_38171);
nand U38286 (N_38286,N_38031,N_38154);
and U38287 (N_38287,N_38116,N_38094);
nor U38288 (N_38288,N_38227,N_38180);
xnor U38289 (N_38289,N_38097,N_38133);
or U38290 (N_38290,N_38081,N_38067);
nor U38291 (N_38291,N_38021,N_38110);
xor U38292 (N_38292,N_38241,N_38107);
nor U38293 (N_38293,N_38119,N_38245);
nor U38294 (N_38294,N_38075,N_38024);
xnor U38295 (N_38295,N_38157,N_38071);
and U38296 (N_38296,N_38162,N_38078);
or U38297 (N_38297,N_38183,N_38005);
nor U38298 (N_38298,N_38129,N_38199);
nor U38299 (N_38299,N_38069,N_38042);
xnor U38300 (N_38300,N_38027,N_38018);
nor U38301 (N_38301,N_38038,N_38219);
or U38302 (N_38302,N_38233,N_38076);
nor U38303 (N_38303,N_38168,N_38006);
or U38304 (N_38304,N_38236,N_38058);
nand U38305 (N_38305,N_38211,N_38193);
and U38306 (N_38306,N_38178,N_38124);
xnor U38307 (N_38307,N_38195,N_38225);
xnor U38308 (N_38308,N_38014,N_38041);
nand U38309 (N_38309,N_38145,N_38165);
or U38310 (N_38310,N_38025,N_38142);
xor U38311 (N_38311,N_38098,N_38140);
and U38312 (N_38312,N_38230,N_38100);
xnor U38313 (N_38313,N_38111,N_38201);
nand U38314 (N_38314,N_38065,N_38115);
and U38315 (N_38315,N_38203,N_38009);
nand U38316 (N_38316,N_38008,N_38044);
nor U38317 (N_38317,N_38197,N_38175);
and U38318 (N_38318,N_38169,N_38217);
xor U38319 (N_38319,N_38234,N_38214);
and U38320 (N_38320,N_38189,N_38167);
nor U38321 (N_38321,N_38173,N_38045);
or U38322 (N_38322,N_38053,N_38020);
nor U38323 (N_38323,N_38139,N_38221);
and U38324 (N_38324,N_38088,N_38143);
and U38325 (N_38325,N_38108,N_38068);
nand U38326 (N_38326,N_38112,N_38181);
nand U38327 (N_38327,N_38091,N_38114);
nor U38328 (N_38328,N_38187,N_38012);
xnor U38329 (N_38329,N_38223,N_38153);
nor U38330 (N_38330,N_38023,N_38174);
nor U38331 (N_38331,N_38247,N_38161);
and U38332 (N_38332,N_38149,N_38017);
xnor U38333 (N_38333,N_38095,N_38015);
xor U38334 (N_38334,N_38096,N_38215);
xnor U38335 (N_38335,N_38192,N_38132);
nor U38336 (N_38336,N_38134,N_38099);
xnor U38337 (N_38337,N_38123,N_38090);
nand U38338 (N_38338,N_38235,N_38013);
nand U38339 (N_38339,N_38073,N_38127);
or U38340 (N_38340,N_38246,N_38226);
nand U38341 (N_38341,N_38034,N_38237);
nor U38342 (N_38342,N_38103,N_38029);
xnor U38343 (N_38343,N_38206,N_38106);
or U38344 (N_38344,N_38105,N_38064);
or U38345 (N_38345,N_38057,N_38249);
nand U38346 (N_38346,N_38122,N_38194);
nand U38347 (N_38347,N_38152,N_38086);
or U38348 (N_38348,N_38080,N_38207);
and U38349 (N_38349,N_38138,N_38137);
nand U38350 (N_38350,N_38166,N_38144);
xor U38351 (N_38351,N_38040,N_38200);
or U38352 (N_38352,N_38019,N_38170);
nand U38353 (N_38353,N_38059,N_38150);
nor U38354 (N_38354,N_38164,N_38109);
and U38355 (N_38355,N_38035,N_38063);
nor U38356 (N_38356,N_38032,N_38229);
nor U38357 (N_38357,N_38163,N_38011);
nand U38358 (N_38358,N_38037,N_38242);
and U38359 (N_38359,N_38000,N_38148);
xnor U38360 (N_38360,N_38050,N_38033);
and U38361 (N_38361,N_38087,N_38022);
xor U38362 (N_38362,N_38185,N_38003);
xor U38363 (N_38363,N_38030,N_38043);
or U38364 (N_38364,N_38102,N_38202);
and U38365 (N_38365,N_38066,N_38243);
xnor U38366 (N_38366,N_38172,N_38062);
nor U38367 (N_38367,N_38052,N_38047);
xor U38368 (N_38368,N_38046,N_38007);
or U38369 (N_38369,N_38156,N_38218);
nand U38370 (N_38370,N_38190,N_38036);
nand U38371 (N_38371,N_38231,N_38055);
xnor U38372 (N_38372,N_38061,N_38232);
or U38373 (N_38373,N_38120,N_38212);
nor U38374 (N_38374,N_38141,N_38160);
nor U38375 (N_38375,N_38108,N_38048);
nor U38376 (N_38376,N_38178,N_38240);
nand U38377 (N_38377,N_38112,N_38212);
or U38378 (N_38378,N_38005,N_38158);
nand U38379 (N_38379,N_38104,N_38039);
nor U38380 (N_38380,N_38049,N_38023);
nand U38381 (N_38381,N_38245,N_38031);
or U38382 (N_38382,N_38120,N_38200);
nor U38383 (N_38383,N_38114,N_38235);
or U38384 (N_38384,N_38200,N_38112);
and U38385 (N_38385,N_38020,N_38048);
and U38386 (N_38386,N_38161,N_38013);
nor U38387 (N_38387,N_38005,N_38166);
nand U38388 (N_38388,N_38035,N_38217);
or U38389 (N_38389,N_38121,N_38196);
and U38390 (N_38390,N_38241,N_38065);
nor U38391 (N_38391,N_38190,N_38215);
nor U38392 (N_38392,N_38107,N_38203);
nand U38393 (N_38393,N_38137,N_38151);
and U38394 (N_38394,N_38087,N_38075);
nor U38395 (N_38395,N_38085,N_38086);
xnor U38396 (N_38396,N_38163,N_38172);
xor U38397 (N_38397,N_38067,N_38235);
nor U38398 (N_38398,N_38233,N_38222);
nor U38399 (N_38399,N_38141,N_38202);
nor U38400 (N_38400,N_38249,N_38147);
or U38401 (N_38401,N_38182,N_38122);
nand U38402 (N_38402,N_38008,N_38199);
or U38403 (N_38403,N_38178,N_38027);
and U38404 (N_38404,N_38087,N_38154);
xnor U38405 (N_38405,N_38208,N_38152);
nor U38406 (N_38406,N_38088,N_38077);
nor U38407 (N_38407,N_38085,N_38069);
and U38408 (N_38408,N_38016,N_38246);
and U38409 (N_38409,N_38103,N_38027);
and U38410 (N_38410,N_38099,N_38118);
and U38411 (N_38411,N_38065,N_38057);
nor U38412 (N_38412,N_38234,N_38195);
and U38413 (N_38413,N_38117,N_38126);
nand U38414 (N_38414,N_38001,N_38186);
nor U38415 (N_38415,N_38110,N_38125);
and U38416 (N_38416,N_38093,N_38101);
or U38417 (N_38417,N_38112,N_38010);
nor U38418 (N_38418,N_38088,N_38013);
and U38419 (N_38419,N_38214,N_38199);
or U38420 (N_38420,N_38209,N_38208);
nand U38421 (N_38421,N_38117,N_38002);
xor U38422 (N_38422,N_38033,N_38091);
or U38423 (N_38423,N_38211,N_38180);
or U38424 (N_38424,N_38166,N_38101);
nand U38425 (N_38425,N_38103,N_38088);
or U38426 (N_38426,N_38085,N_38158);
nor U38427 (N_38427,N_38123,N_38233);
nand U38428 (N_38428,N_38213,N_38039);
nand U38429 (N_38429,N_38044,N_38191);
xnor U38430 (N_38430,N_38078,N_38177);
or U38431 (N_38431,N_38010,N_38183);
nor U38432 (N_38432,N_38144,N_38219);
and U38433 (N_38433,N_38187,N_38040);
xnor U38434 (N_38434,N_38152,N_38150);
or U38435 (N_38435,N_38013,N_38146);
nand U38436 (N_38436,N_38067,N_38148);
xor U38437 (N_38437,N_38227,N_38143);
and U38438 (N_38438,N_38165,N_38192);
and U38439 (N_38439,N_38040,N_38019);
or U38440 (N_38440,N_38000,N_38227);
or U38441 (N_38441,N_38004,N_38020);
nor U38442 (N_38442,N_38087,N_38191);
or U38443 (N_38443,N_38095,N_38025);
and U38444 (N_38444,N_38112,N_38006);
nand U38445 (N_38445,N_38226,N_38046);
nor U38446 (N_38446,N_38046,N_38225);
nor U38447 (N_38447,N_38184,N_38145);
or U38448 (N_38448,N_38091,N_38216);
nand U38449 (N_38449,N_38192,N_38154);
nor U38450 (N_38450,N_38114,N_38199);
nor U38451 (N_38451,N_38024,N_38036);
or U38452 (N_38452,N_38058,N_38099);
or U38453 (N_38453,N_38120,N_38039);
nand U38454 (N_38454,N_38097,N_38248);
xor U38455 (N_38455,N_38193,N_38081);
and U38456 (N_38456,N_38056,N_38206);
or U38457 (N_38457,N_38203,N_38118);
xnor U38458 (N_38458,N_38197,N_38007);
and U38459 (N_38459,N_38048,N_38167);
xnor U38460 (N_38460,N_38121,N_38037);
nor U38461 (N_38461,N_38064,N_38023);
xnor U38462 (N_38462,N_38156,N_38223);
xnor U38463 (N_38463,N_38058,N_38174);
nor U38464 (N_38464,N_38215,N_38133);
nor U38465 (N_38465,N_38233,N_38007);
nand U38466 (N_38466,N_38239,N_38001);
xnor U38467 (N_38467,N_38041,N_38202);
or U38468 (N_38468,N_38186,N_38203);
xnor U38469 (N_38469,N_38007,N_38006);
or U38470 (N_38470,N_38150,N_38239);
nor U38471 (N_38471,N_38244,N_38091);
xor U38472 (N_38472,N_38216,N_38181);
nand U38473 (N_38473,N_38090,N_38111);
xnor U38474 (N_38474,N_38183,N_38134);
nand U38475 (N_38475,N_38196,N_38130);
nand U38476 (N_38476,N_38046,N_38205);
and U38477 (N_38477,N_38230,N_38248);
or U38478 (N_38478,N_38044,N_38074);
or U38479 (N_38479,N_38055,N_38171);
xnor U38480 (N_38480,N_38059,N_38198);
nor U38481 (N_38481,N_38091,N_38167);
nand U38482 (N_38482,N_38099,N_38048);
xor U38483 (N_38483,N_38155,N_38046);
nor U38484 (N_38484,N_38188,N_38228);
nor U38485 (N_38485,N_38011,N_38075);
xor U38486 (N_38486,N_38033,N_38164);
nand U38487 (N_38487,N_38006,N_38053);
or U38488 (N_38488,N_38197,N_38107);
nor U38489 (N_38489,N_38183,N_38157);
nor U38490 (N_38490,N_38132,N_38168);
nor U38491 (N_38491,N_38064,N_38005);
nor U38492 (N_38492,N_38204,N_38033);
and U38493 (N_38493,N_38131,N_38171);
xor U38494 (N_38494,N_38208,N_38174);
nor U38495 (N_38495,N_38202,N_38170);
nand U38496 (N_38496,N_38084,N_38166);
or U38497 (N_38497,N_38062,N_38093);
and U38498 (N_38498,N_38123,N_38013);
nand U38499 (N_38499,N_38198,N_38184);
or U38500 (N_38500,N_38437,N_38351);
and U38501 (N_38501,N_38454,N_38383);
and U38502 (N_38502,N_38330,N_38285);
nor U38503 (N_38503,N_38290,N_38271);
and U38504 (N_38504,N_38413,N_38323);
nand U38505 (N_38505,N_38428,N_38334);
nor U38506 (N_38506,N_38306,N_38321);
and U38507 (N_38507,N_38436,N_38302);
nor U38508 (N_38508,N_38345,N_38344);
xnor U38509 (N_38509,N_38389,N_38253);
xor U38510 (N_38510,N_38269,N_38419);
or U38511 (N_38511,N_38267,N_38405);
or U38512 (N_38512,N_38422,N_38432);
nor U38513 (N_38513,N_38361,N_38494);
nand U38514 (N_38514,N_38399,N_38289);
nand U38515 (N_38515,N_38339,N_38411);
nand U38516 (N_38516,N_38470,N_38355);
nand U38517 (N_38517,N_38318,N_38426);
and U38518 (N_38518,N_38311,N_38486);
nand U38519 (N_38519,N_38392,N_38370);
nor U38520 (N_38520,N_38412,N_38309);
nand U38521 (N_38521,N_38319,N_38439);
and U38522 (N_38522,N_38406,N_38366);
and U38523 (N_38523,N_38433,N_38336);
nor U38524 (N_38524,N_38273,N_38372);
nand U38525 (N_38525,N_38382,N_38275);
and U38526 (N_38526,N_38260,N_38394);
and U38527 (N_38527,N_38281,N_38299);
nand U38528 (N_38528,N_38320,N_38356);
or U38529 (N_38529,N_38473,N_38430);
and U38530 (N_38530,N_38326,N_38386);
nand U38531 (N_38531,N_38313,N_38305);
and U38532 (N_38532,N_38468,N_38447);
nor U38533 (N_38533,N_38448,N_38373);
nand U38534 (N_38534,N_38272,N_38469);
and U38535 (N_38535,N_38300,N_38472);
and U38536 (N_38536,N_38446,N_38251);
and U38537 (N_38537,N_38458,N_38467);
or U38538 (N_38538,N_38292,N_38404);
xor U38539 (N_38539,N_38352,N_38354);
nand U38540 (N_38540,N_38474,N_38358);
nor U38541 (N_38541,N_38398,N_38315);
nand U38542 (N_38542,N_38441,N_38410);
nand U38543 (N_38543,N_38298,N_38431);
or U38544 (N_38544,N_38391,N_38387);
xnor U38545 (N_38545,N_38375,N_38371);
or U38546 (N_38546,N_38416,N_38477);
nand U38547 (N_38547,N_38396,N_38332);
nand U38548 (N_38548,N_38483,N_38489);
xor U38549 (N_38549,N_38350,N_38402);
xnor U38550 (N_38550,N_38367,N_38480);
xor U38551 (N_38551,N_38484,N_38445);
and U38552 (N_38552,N_38342,N_38481);
and U38553 (N_38553,N_38282,N_38308);
xnor U38554 (N_38554,N_38452,N_38459);
nand U38555 (N_38555,N_38393,N_38461);
or U38556 (N_38556,N_38429,N_38450);
xnor U38557 (N_38557,N_38363,N_38335);
or U38558 (N_38558,N_38485,N_38362);
xnor U38559 (N_38559,N_38258,N_38464);
nand U38560 (N_38560,N_38286,N_38257);
and U38561 (N_38561,N_38487,N_38284);
nand U38562 (N_38562,N_38353,N_38407);
nand U38563 (N_38563,N_38263,N_38415);
and U38564 (N_38564,N_38434,N_38337);
or U38565 (N_38565,N_38277,N_38423);
and U38566 (N_38566,N_38498,N_38291);
nor U38567 (N_38567,N_38368,N_38264);
nor U38568 (N_38568,N_38325,N_38380);
nand U38569 (N_38569,N_38471,N_38322);
nand U38570 (N_38570,N_38478,N_38384);
nor U38571 (N_38571,N_38314,N_38397);
nor U38572 (N_38572,N_38463,N_38347);
or U38573 (N_38573,N_38297,N_38390);
xor U38574 (N_38574,N_38421,N_38377);
nor U38575 (N_38575,N_38265,N_38427);
xnor U38576 (N_38576,N_38476,N_38466);
and U38577 (N_38577,N_38274,N_38425);
nand U38578 (N_38578,N_38493,N_38495);
nor U38579 (N_38579,N_38409,N_38346);
or U38580 (N_38580,N_38379,N_38418);
nor U38581 (N_38581,N_38499,N_38360);
nand U38582 (N_38582,N_38250,N_38435);
or U38583 (N_38583,N_38369,N_38276);
or U38584 (N_38584,N_38301,N_38288);
nor U38585 (N_38585,N_38252,N_38261);
or U38586 (N_38586,N_38255,N_38328);
or U38587 (N_38587,N_38293,N_38333);
nand U38588 (N_38588,N_38462,N_38482);
nand U38589 (N_38589,N_38451,N_38440);
and U38590 (N_38590,N_38400,N_38457);
or U38591 (N_38591,N_38338,N_38401);
nand U38592 (N_38592,N_38327,N_38294);
and U38593 (N_38593,N_38374,N_38388);
or U38594 (N_38594,N_38317,N_38341);
nor U38595 (N_38595,N_38455,N_38343);
nor U38596 (N_38596,N_38262,N_38312);
or U38597 (N_38597,N_38449,N_38340);
and U38598 (N_38598,N_38278,N_38438);
nor U38599 (N_38599,N_38479,N_38490);
nand U38600 (N_38600,N_38296,N_38408);
xor U38601 (N_38601,N_38492,N_38364);
or U38602 (N_38602,N_38417,N_38414);
or U38603 (N_38603,N_38270,N_38287);
xor U38604 (N_38604,N_38442,N_38376);
nor U38605 (N_38605,N_38349,N_38496);
xnor U38606 (N_38606,N_38395,N_38303);
or U38607 (N_38607,N_38488,N_38385);
nand U38608 (N_38608,N_38497,N_38465);
and U38609 (N_38609,N_38420,N_38357);
nor U38610 (N_38610,N_38348,N_38316);
nand U38611 (N_38611,N_38359,N_38266);
and U38612 (N_38612,N_38475,N_38256);
and U38613 (N_38613,N_38456,N_38444);
nand U38614 (N_38614,N_38460,N_38365);
xnor U38615 (N_38615,N_38381,N_38254);
and U38616 (N_38616,N_38324,N_38279);
or U38617 (N_38617,N_38268,N_38295);
nand U38618 (N_38618,N_38331,N_38307);
or U38619 (N_38619,N_38310,N_38304);
nor U38620 (N_38620,N_38378,N_38453);
nand U38621 (N_38621,N_38329,N_38283);
or U38622 (N_38622,N_38403,N_38424);
and U38623 (N_38623,N_38280,N_38491);
nand U38624 (N_38624,N_38259,N_38443);
and U38625 (N_38625,N_38415,N_38318);
xor U38626 (N_38626,N_38409,N_38255);
nand U38627 (N_38627,N_38446,N_38385);
nor U38628 (N_38628,N_38333,N_38311);
xnor U38629 (N_38629,N_38397,N_38267);
or U38630 (N_38630,N_38442,N_38294);
nor U38631 (N_38631,N_38297,N_38425);
nor U38632 (N_38632,N_38309,N_38292);
nor U38633 (N_38633,N_38467,N_38279);
and U38634 (N_38634,N_38366,N_38301);
nand U38635 (N_38635,N_38440,N_38488);
nor U38636 (N_38636,N_38272,N_38323);
and U38637 (N_38637,N_38471,N_38487);
and U38638 (N_38638,N_38292,N_38428);
and U38639 (N_38639,N_38284,N_38364);
or U38640 (N_38640,N_38399,N_38385);
xor U38641 (N_38641,N_38406,N_38376);
nor U38642 (N_38642,N_38372,N_38395);
nand U38643 (N_38643,N_38321,N_38358);
nor U38644 (N_38644,N_38384,N_38454);
nor U38645 (N_38645,N_38373,N_38475);
nand U38646 (N_38646,N_38260,N_38356);
nand U38647 (N_38647,N_38484,N_38279);
nor U38648 (N_38648,N_38414,N_38261);
nor U38649 (N_38649,N_38418,N_38450);
nand U38650 (N_38650,N_38492,N_38468);
nor U38651 (N_38651,N_38455,N_38282);
nand U38652 (N_38652,N_38407,N_38367);
nor U38653 (N_38653,N_38487,N_38320);
xor U38654 (N_38654,N_38384,N_38265);
or U38655 (N_38655,N_38353,N_38433);
nor U38656 (N_38656,N_38415,N_38402);
or U38657 (N_38657,N_38361,N_38328);
or U38658 (N_38658,N_38305,N_38472);
nand U38659 (N_38659,N_38378,N_38332);
nand U38660 (N_38660,N_38288,N_38479);
or U38661 (N_38661,N_38264,N_38314);
xor U38662 (N_38662,N_38370,N_38343);
xnor U38663 (N_38663,N_38366,N_38305);
nand U38664 (N_38664,N_38493,N_38359);
nor U38665 (N_38665,N_38264,N_38279);
or U38666 (N_38666,N_38360,N_38336);
xor U38667 (N_38667,N_38361,N_38438);
and U38668 (N_38668,N_38299,N_38398);
or U38669 (N_38669,N_38283,N_38361);
xor U38670 (N_38670,N_38398,N_38258);
xnor U38671 (N_38671,N_38366,N_38331);
or U38672 (N_38672,N_38337,N_38278);
and U38673 (N_38673,N_38279,N_38481);
xor U38674 (N_38674,N_38318,N_38497);
xor U38675 (N_38675,N_38381,N_38377);
or U38676 (N_38676,N_38266,N_38399);
xnor U38677 (N_38677,N_38288,N_38312);
xnor U38678 (N_38678,N_38477,N_38283);
and U38679 (N_38679,N_38447,N_38305);
or U38680 (N_38680,N_38456,N_38496);
nor U38681 (N_38681,N_38450,N_38495);
xnor U38682 (N_38682,N_38356,N_38365);
and U38683 (N_38683,N_38436,N_38414);
and U38684 (N_38684,N_38309,N_38326);
nand U38685 (N_38685,N_38260,N_38449);
nor U38686 (N_38686,N_38290,N_38378);
nand U38687 (N_38687,N_38378,N_38449);
nand U38688 (N_38688,N_38349,N_38298);
nor U38689 (N_38689,N_38269,N_38352);
and U38690 (N_38690,N_38251,N_38318);
nand U38691 (N_38691,N_38395,N_38383);
or U38692 (N_38692,N_38281,N_38353);
nor U38693 (N_38693,N_38307,N_38373);
or U38694 (N_38694,N_38462,N_38364);
and U38695 (N_38695,N_38335,N_38312);
or U38696 (N_38696,N_38274,N_38270);
xor U38697 (N_38697,N_38357,N_38290);
and U38698 (N_38698,N_38394,N_38286);
and U38699 (N_38699,N_38259,N_38258);
xor U38700 (N_38700,N_38408,N_38487);
nor U38701 (N_38701,N_38302,N_38311);
or U38702 (N_38702,N_38309,N_38323);
nor U38703 (N_38703,N_38262,N_38430);
nor U38704 (N_38704,N_38483,N_38382);
nand U38705 (N_38705,N_38264,N_38268);
xnor U38706 (N_38706,N_38470,N_38464);
or U38707 (N_38707,N_38445,N_38322);
nand U38708 (N_38708,N_38400,N_38264);
or U38709 (N_38709,N_38349,N_38312);
or U38710 (N_38710,N_38382,N_38306);
nand U38711 (N_38711,N_38253,N_38441);
nor U38712 (N_38712,N_38352,N_38418);
and U38713 (N_38713,N_38400,N_38374);
and U38714 (N_38714,N_38287,N_38492);
nor U38715 (N_38715,N_38255,N_38254);
and U38716 (N_38716,N_38422,N_38346);
nor U38717 (N_38717,N_38371,N_38271);
nand U38718 (N_38718,N_38489,N_38451);
and U38719 (N_38719,N_38408,N_38465);
nor U38720 (N_38720,N_38303,N_38408);
nor U38721 (N_38721,N_38313,N_38384);
or U38722 (N_38722,N_38454,N_38348);
nor U38723 (N_38723,N_38481,N_38488);
and U38724 (N_38724,N_38317,N_38417);
nand U38725 (N_38725,N_38330,N_38450);
nand U38726 (N_38726,N_38303,N_38455);
nor U38727 (N_38727,N_38267,N_38451);
nand U38728 (N_38728,N_38342,N_38306);
nor U38729 (N_38729,N_38395,N_38455);
or U38730 (N_38730,N_38364,N_38385);
nand U38731 (N_38731,N_38310,N_38464);
nand U38732 (N_38732,N_38332,N_38387);
and U38733 (N_38733,N_38342,N_38493);
nand U38734 (N_38734,N_38290,N_38393);
and U38735 (N_38735,N_38431,N_38339);
or U38736 (N_38736,N_38386,N_38324);
nand U38737 (N_38737,N_38351,N_38489);
or U38738 (N_38738,N_38305,N_38379);
or U38739 (N_38739,N_38271,N_38487);
nor U38740 (N_38740,N_38442,N_38256);
or U38741 (N_38741,N_38484,N_38332);
or U38742 (N_38742,N_38371,N_38404);
nand U38743 (N_38743,N_38374,N_38476);
nor U38744 (N_38744,N_38358,N_38445);
and U38745 (N_38745,N_38294,N_38453);
or U38746 (N_38746,N_38409,N_38430);
or U38747 (N_38747,N_38300,N_38461);
nand U38748 (N_38748,N_38381,N_38251);
nor U38749 (N_38749,N_38362,N_38493);
nand U38750 (N_38750,N_38733,N_38676);
nand U38751 (N_38751,N_38502,N_38720);
xor U38752 (N_38752,N_38659,N_38526);
nor U38753 (N_38753,N_38584,N_38637);
nand U38754 (N_38754,N_38599,N_38743);
and U38755 (N_38755,N_38678,N_38523);
or U38756 (N_38756,N_38545,N_38551);
or U38757 (N_38757,N_38604,N_38538);
nand U38758 (N_38758,N_38559,N_38650);
xor U38759 (N_38759,N_38593,N_38716);
and U38760 (N_38760,N_38556,N_38530);
xor U38761 (N_38761,N_38597,N_38671);
nand U38762 (N_38762,N_38610,N_38581);
or U38763 (N_38763,N_38702,N_38585);
nand U38764 (N_38764,N_38638,N_38516);
nand U38765 (N_38765,N_38669,N_38713);
or U38766 (N_38766,N_38614,N_38651);
nand U38767 (N_38767,N_38629,N_38700);
nor U38768 (N_38768,N_38693,N_38578);
and U38769 (N_38769,N_38665,N_38594);
and U38770 (N_38770,N_38505,N_38606);
xnor U38771 (N_38771,N_38673,N_38697);
xnor U38772 (N_38772,N_38736,N_38570);
nor U38773 (N_38773,N_38686,N_38692);
or U38774 (N_38774,N_38653,N_38684);
nand U38775 (N_38775,N_38520,N_38558);
or U38776 (N_38776,N_38740,N_38646);
or U38777 (N_38777,N_38577,N_38679);
and U38778 (N_38778,N_38633,N_38617);
xnor U38779 (N_38779,N_38544,N_38567);
nor U38780 (N_38780,N_38640,N_38627);
xor U38781 (N_38781,N_38726,N_38608);
nand U38782 (N_38782,N_38503,N_38722);
xnor U38783 (N_38783,N_38694,N_38601);
nand U38784 (N_38784,N_38623,N_38647);
and U38785 (N_38785,N_38712,N_38714);
nand U38786 (N_38786,N_38572,N_38685);
nor U38787 (N_38787,N_38718,N_38737);
xor U38788 (N_38788,N_38521,N_38555);
and U38789 (N_38789,N_38571,N_38724);
xnor U38790 (N_38790,N_38549,N_38660);
nand U38791 (N_38791,N_38500,N_38707);
nand U38792 (N_38792,N_38634,N_38546);
xor U38793 (N_38793,N_38698,N_38618);
or U38794 (N_38794,N_38525,N_38540);
and U38795 (N_38795,N_38613,N_38612);
or U38796 (N_38796,N_38598,N_38735);
and U38797 (N_38797,N_38732,N_38742);
xor U38798 (N_38798,N_38553,N_38682);
xnor U38799 (N_38799,N_38652,N_38605);
or U38800 (N_38800,N_38579,N_38699);
and U38801 (N_38801,N_38576,N_38519);
xor U38802 (N_38802,N_38518,N_38506);
or U38803 (N_38803,N_38661,N_38715);
and U38804 (N_38804,N_38644,N_38591);
xor U38805 (N_38805,N_38522,N_38547);
nand U38806 (N_38806,N_38690,N_38550);
nor U38807 (N_38807,N_38607,N_38619);
and U38808 (N_38808,N_38741,N_38729);
nor U38809 (N_38809,N_38527,N_38675);
nor U38810 (N_38810,N_38511,N_38536);
nor U38811 (N_38811,N_38552,N_38749);
nor U38812 (N_38812,N_38542,N_38711);
or U38813 (N_38813,N_38674,N_38664);
nor U38814 (N_38814,N_38744,N_38639);
nor U38815 (N_38815,N_38562,N_38709);
or U38816 (N_38816,N_38534,N_38717);
and U38817 (N_38817,N_38504,N_38509);
and U38818 (N_38818,N_38602,N_38573);
nor U38819 (N_38819,N_38668,N_38508);
xnor U38820 (N_38820,N_38636,N_38582);
nand U38821 (N_38821,N_38663,N_38658);
xor U38822 (N_38822,N_38512,N_38725);
and U38823 (N_38823,N_38730,N_38507);
xnor U38824 (N_38824,N_38710,N_38681);
nand U38825 (N_38825,N_38721,N_38734);
and U38826 (N_38826,N_38515,N_38603);
or U38827 (N_38827,N_38643,N_38696);
nor U38828 (N_38828,N_38514,N_38510);
nand U38829 (N_38829,N_38541,N_38641);
nand U38830 (N_38830,N_38532,N_38662);
and U38831 (N_38831,N_38738,N_38600);
nor U38832 (N_38832,N_38630,N_38667);
or U38833 (N_38833,N_38654,N_38719);
or U38834 (N_38834,N_38621,N_38628);
or U38835 (N_38835,N_38706,N_38580);
and U38836 (N_38836,N_38731,N_38746);
and U38837 (N_38837,N_38648,N_38535);
or U38838 (N_38838,N_38677,N_38590);
xnor U38839 (N_38839,N_38583,N_38561);
xnor U38840 (N_38840,N_38689,N_38595);
and U38841 (N_38841,N_38748,N_38632);
and U38842 (N_38842,N_38586,N_38529);
xnor U38843 (N_38843,N_38565,N_38539);
or U38844 (N_38844,N_38635,N_38655);
xor U38845 (N_38845,N_38611,N_38587);
xor U38846 (N_38846,N_38566,N_38588);
nor U38847 (N_38847,N_38703,N_38691);
nand U38848 (N_38848,N_38624,N_38657);
nor U38849 (N_38849,N_38688,N_38695);
nand U38850 (N_38850,N_38728,N_38723);
or U38851 (N_38851,N_38620,N_38528);
and U38852 (N_38852,N_38560,N_38642);
or U38853 (N_38853,N_38569,N_38649);
nor U38854 (N_38854,N_38574,N_38745);
nand U38855 (N_38855,N_38531,N_38513);
or U38856 (N_38856,N_38524,N_38656);
or U38857 (N_38857,N_38626,N_38589);
xor U38858 (N_38858,N_38687,N_38622);
xor U38859 (N_38859,N_38609,N_38616);
nor U38860 (N_38860,N_38537,N_38548);
and U38861 (N_38861,N_38704,N_38683);
and U38862 (N_38862,N_38564,N_38631);
nand U38863 (N_38863,N_38672,N_38533);
xnor U38864 (N_38864,N_38670,N_38680);
nand U38865 (N_38865,N_38727,N_38554);
and U38866 (N_38866,N_38563,N_38625);
nor U38867 (N_38867,N_38557,N_38708);
xnor U38868 (N_38868,N_38592,N_38705);
or U38869 (N_38869,N_38701,N_38543);
and U38870 (N_38870,N_38615,N_38645);
nand U38871 (N_38871,N_38501,N_38747);
and U38872 (N_38872,N_38517,N_38596);
xor U38873 (N_38873,N_38666,N_38575);
xnor U38874 (N_38874,N_38568,N_38739);
nor U38875 (N_38875,N_38554,N_38650);
nor U38876 (N_38876,N_38636,N_38685);
xor U38877 (N_38877,N_38565,N_38699);
and U38878 (N_38878,N_38719,N_38691);
and U38879 (N_38879,N_38704,N_38544);
and U38880 (N_38880,N_38504,N_38596);
nor U38881 (N_38881,N_38715,N_38727);
nor U38882 (N_38882,N_38631,N_38712);
and U38883 (N_38883,N_38565,N_38570);
nand U38884 (N_38884,N_38546,N_38707);
or U38885 (N_38885,N_38748,N_38505);
xnor U38886 (N_38886,N_38689,N_38578);
and U38887 (N_38887,N_38569,N_38634);
nor U38888 (N_38888,N_38684,N_38640);
nand U38889 (N_38889,N_38546,N_38725);
xor U38890 (N_38890,N_38668,N_38594);
nor U38891 (N_38891,N_38598,N_38573);
and U38892 (N_38892,N_38675,N_38678);
nor U38893 (N_38893,N_38537,N_38605);
or U38894 (N_38894,N_38530,N_38536);
or U38895 (N_38895,N_38517,N_38585);
nand U38896 (N_38896,N_38511,N_38605);
nand U38897 (N_38897,N_38697,N_38550);
xor U38898 (N_38898,N_38651,N_38507);
and U38899 (N_38899,N_38624,N_38532);
nor U38900 (N_38900,N_38672,N_38619);
and U38901 (N_38901,N_38667,N_38557);
and U38902 (N_38902,N_38591,N_38697);
or U38903 (N_38903,N_38725,N_38672);
xnor U38904 (N_38904,N_38700,N_38658);
nor U38905 (N_38905,N_38729,N_38669);
or U38906 (N_38906,N_38651,N_38677);
xnor U38907 (N_38907,N_38650,N_38522);
xnor U38908 (N_38908,N_38523,N_38568);
xnor U38909 (N_38909,N_38626,N_38623);
or U38910 (N_38910,N_38679,N_38554);
nor U38911 (N_38911,N_38580,N_38730);
nand U38912 (N_38912,N_38529,N_38627);
xor U38913 (N_38913,N_38744,N_38706);
and U38914 (N_38914,N_38703,N_38645);
nor U38915 (N_38915,N_38639,N_38512);
and U38916 (N_38916,N_38679,N_38659);
or U38917 (N_38917,N_38701,N_38559);
xnor U38918 (N_38918,N_38636,N_38593);
xor U38919 (N_38919,N_38730,N_38567);
nor U38920 (N_38920,N_38661,N_38519);
or U38921 (N_38921,N_38623,N_38703);
nor U38922 (N_38922,N_38535,N_38689);
xnor U38923 (N_38923,N_38711,N_38596);
nand U38924 (N_38924,N_38623,N_38660);
and U38925 (N_38925,N_38529,N_38654);
nor U38926 (N_38926,N_38710,N_38736);
nand U38927 (N_38927,N_38539,N_38519);
and U38928 (N_38928,N_38681,N_38673);
nand U38929 (N_38929,N_38729,N_38672);
and U38930 (N_38930,N_38741,N_38501);
xor U38931 (N_38931,N_38727,N_38571);
and U38932 (N_38932,N_38583,N_38578);
or U38933 (N_38933,N_38692,N_38624);
or U38934 (N_38934,N_38673,N_38509);
and U38935 (N_38935,N_38683,N_38570);
nand U38936 (N_38936,N_38534,N_38730);
nor U38937 (N_38937,N_38506,N_38523);
nand U38938 (N_38938,N_38614,N_38591);
xor U38939 (N_38939,N_38534,N_38708);
nor U38940 (N_38940,N_38508,N_38509);
and U38941 (N_38941,N_38649,N_38663);
xnor U38942 (N_38942,N_38639,N_38601);
nand U38943 (N_38943,N_38714,N_38672);
xor U38944 (N_38944,N_38556,N_38599);
nand U38945 (N_38945,N_38592,N_38602);
nand U38946 (N_38946,N_38592,N_38582);
xor U38947 (N_38947,N_38728,N_38630);
xnor U38948 (N_38948,N_38591,N_38616);
and U38949 (N_38949,N_38727,N_38541);
or U38950 (N_38950,N_38572,N_38627);
xnor U38951 (N_38951,N_38555,N_38736);
and U38952 (N_38952,N_38531,N_38527);
nand U38953 (N_38953,N_38594,N_38644);
nand U38954 (N_38954,N_38557,N_38565);
and U38955 (N_38955,N_38713,N_38708);
or U38956 (N_38956,N_38742,N_38525);
and U38957 (N_38957,N_38605,N_38530);
xnor U38958 (N_38958,N_38682,N_38726);
nor U38959 (N_38959,N_38644,N_38697);
nor U38960 (N_38960,N_38592,N_38529);
xnor U38961 (N_38961,N_38684,N_38581);
xor U38962 (N_38962,N_38645,N_38688);
nand U38963 (N_38963,N_38624,N_38749);
or U38964 (N_38964,N_38513,N_38743);
and U38965 (N_38965,N_38609,N_38684);
nor U38966 (N_38966,N_38580,N_38733);
nand U38967 (N_38967,N_38724,N_38681);
and U38968 (N_38968,N_38634,N_38622);
nor U38969 (N_38969,N_38699,N_38596);
nor U38970 (N_38970,N_38675,N_38744);
nand U38971 (N_38971,N_38579,N_38501);
nand U38972 (N_38972,N_38723,N_38668);
nor U38973 (N_38973,N_38547,N_38552);
nand U38974 (N_38974,N_38606,N_38502);
or U38975 (N_38975,N_38586,N_38523);
and U38976 (N_38976,N_38739,N_38641);
or U38977 (N_38977,N_38622,N_38552);
xnor U38978 (N_38978,N_38528,N_38624);
or U38979 (N_38979,N_38504,N_38512);
nand U38980 (N_38980,N_38746,N_38502);
or U38981 (N_38981,N_38564,N_38740);
and U38982 (N_38982,N_38739,N_38524);
or U38983 (N_38983,N_38684,N_38582);
and U38984 (N_38984,N_38581,N_38540);
and U38985 (N_38985,N_38713,N_38679);
or U38986 (N_38986,N_38519,N_38550);
nand U38987 (N_38987,N_38667,N_38681);
and U38988 (N_38988,N_38583,N_38702);
xor U38989 (N_38989,N_38653,N_38528);
xor U38990 (N_38990,N_38564,N_38625);
nand U38991 (N_38991,N_38591,N_38642);
nand U38992 (N_38992,N_38578,N_38674);
nand U38993 (N_38993,N_38734,N_38660);
nor U38994 (N_38994,N_38536,N_38729);
nand U38995 (N_38995,N_38564,N_38520);
xor U38996 (N_38996,N_38721,N_38702);
xor U38997 (N_38997,N_38578,N_38545);
or U38998 (N_38998,N_38734,N_38645);
xnor U38999 (N_38999,N_38743,N_38701);
and U39000 (N_39000,N_38782,N_38918);
or U39001 (N_39001,N_38949,N_38812);
nor U39002 (N_39002,N_38974,N_38943);
and U39003 (N_39003,N_38940,N_38937);
and U39004 (N_39004,N_38878,N_38787);
and U39005 (N_39005,N_38880,N_38972);
nand U39006 (N_39006,N_38927,N_38766);
nor U39007 (N_39007,N_38924,N_38803);
nand U39008 (N_39008,N_38768,N_38942);
and U39009 (N_39009,N_38896,N_38993);
nand U39010 (N_39010,N_38981,N_38914);
nor U39011 (N_39011,N_38967,N_38781);
nor U39012 (N_39012,N_38865,N_38952);
or U39013 (N_39013,N_38859,N_38917);
nor U39014 (N_39014,N_38759,N_38767);
and U39015 (N_39015,N_38854,N_38790);
and U39016 (N_39016,N_38794,N_38816);
nor U39017 (N_39017,N_38776,N_38826);
xor U39018 (N_39018,N_38801,N_38874);
nor U39019 (N_39019,N_38983,N_38906);
or U39020 (N_39020,N_38779,N_38910);
xnor U39021 (N_39021,N_38909,N_38979);
nand U39022 (N_39022,N_38875,N_38838);
nand U39023 (N_39023,N_38893,N_38948);
and U39024 (N_39024,N_38808,N_38793);
nor U39025 (N_39025,N_38856,N_38950);
and U39026 (N_39026,N_38897,N_38785);
xor U39027 (N_39027,N_38847,N_38822);
nor U39028 (N_39028,N_38925,N_38770);
nand U39029 (N_39029,N_38849,N_38971);
xor U39030 (N_39030,N_38962,N_38860);
or U39031 (N_39031,N_38858,N_38901);
or U39032 (N_39032,N_38944,N_38886);
nor U39033 (N_39033,N_38888,N_38818);
or U39034 (N_39034,N_38987,N_38795);
and U39035 (N_39035,N_38791,N_38800);
xnor U39036 (N_39036,N_38898,N_38783);
xnor U39037 (N_39037,N_38881,N_38923);
nor U39038 (N_39038,N_38955,N_38855);
xor U39039 (N_39039,N_38862,N_38991);
or U39040 (N_39040,N_38945,N_38934);
xnor U39041 (N_39041,N_38778,N_38756);
xor U39042 (N_39042,N_38840,N_38763);
xor U39043 (N_39043,N_38941,N_38866);
xnor U39044 (N_39044,N_38951,N_38879);
nor U39045 (N_39045,N_38830,N_38869);
nor U39046 (N_39046,N_38958,N_38841);
or U39047 (N_39047,N_38820,N_38931);
or U39048 (N_39048,N_38905,N_38761);
or U39049 (N_39049,N_38789,N_38873);
nand U39050 (N_39050,N_38960,N_38932);
and U39051 (N_39051,N_38844,N_38947);
nor U39052 (N_39052,N_38807,N_38842);
nor U39053 (N_39053,N_38902,N_38883);
xor U39054 (N_39054,N_38913,N_38821);
nor U39055 (N_39055,N_38895,N_38999);
nor U39056 (N_39056,N_38959,N_38775);
and U39057 (N_39057,N_38806,N_38824);
and U39058 (N_39058,N_38890,N_38996);
or U39059 (N_39059,N_38939,N_38760);
xnor U39060 (N_39060,N_38930,N_38980);
nor U39061 (N_39061,N_38815,N_38919);
nor U39062 (N_39062,N_38846,N_38753);
nand U39063 (N_39063,N_38839,N_38811);
nor U39064 (N_39064,N_38798,N_38894);
xnor U39065 (N_39065,N_38863,N_38965);
and U39066 (N_39066,N_38887,N_38836);
nand U39067 (N_39067,N_38900,N_38852);
xor U39068 (N_39068,N_38963,N_38825);
and U39069 (N_39069,N_38982,N_38904);
xor U39070 (N_39070,N_38764,N_38953);
xor U39071 (N_39071,N_38903,N_38968);
nor U39072 (N_39072,N_38851,N_38978);
or U39073 (N_39073,N_38975,N_38899);
nand U39074 (N_39074,N_38915,N_38845);
nor U39075 (N_39075,N_38837,N_38973);
and U39076 (N_39076,N_38833,N_38989);
and U39077 (N_39077,N_38802,N_38884);
nand U39078 (N_39078,N_38861,N_38867);
nand U39079 (N_39079,N_38929,N_38769);
or U39080 (N_39080,N_38977,N_38907);
nor U39081 (N_39081,N_38813,N_38876);
or U39082 (N_39082,N_38870,N_38857);
nand U39083 (N_39083,N_38786,N_38755);
or U39084 (N_39084,N_38889,N_38774);
nand U39085 (N_39085,N_38810,N_38936);
and U39086 (N_39086,N_38792,N_38938);
nand U39087 (N_39087,N_38809,N_38969);
or U39088 (N_39088,N_38750,N_38850);
nand U39089 (N_39089,N_38751,N_38788);
or U39090 (N_39090,N_38777,N_38926);
nor U39091 (N_39091,N_38928,N_38831);
nor U39092 (N_39092,N_38762,N_38864);
nand U39093 (N_39093,N_38920,N_38908);
nand U39094 (N_39094,N_38997,N_38758);
xor U39095 (N_39095,N_38805,N_38765);
or U39096 (N_39096,N_38985,N_38771);
or U39097 (N_39097,N_38922,N_38877);
and U39098 (N_39098,N_38804,N_38871);
xor U39099 (N_39099,N_38853,N_38957);
or U39100 (N_39100,N_38935,N_38998);
and U39101 (N_39101,N_38784,N_38892);
xnor U39102 (N_39102,N_38970,N_38992);
xor U39103 (N_39103,N_38921,N_38986);
or U39104 (N_39104,N_38994,N_38872);
or U39105 (N_39105,N_38946,N_38964);
or U39106 (N_39106,N_38772,N_38752);
nand U39107 (N_39107,N_38911,N_38754);
nand U39108 (N_39108,N_38796,N_38916);
xor U39109 (N_39109,N_38819,N_38933);
nor U39110 (N_39110,N_38988,N_38882);
xor U39111 (N_39111,N_38797,N_38868);
nand U39112 (N_39112,N_38832,N_38773);
and U39113 (N_39113,N_38956,N_38990);
or U39114 (N_39114,N_38799,N_38843);
nand U39115 (N_39115,N_38814,N_38891);
and U39116 (N_39116,N_38966,N_38828);
nor U39117 (N_39117,N_38984,N_38823);
nor U39118 (N_39118,N_38780,N_38757);
and U39119 (N_39119,N_38976,N_38885);
nand U39120 (N_39120,N_38829,N_38954);
and U39121 (N_39121,N_38995,N_38848);
and U39122 (N_39122,N_38834,N_38827);
or U39123 (N_39123,N_38817,N_38912);
nand U39124 (N_39124,N_38835,N_38961);
xor U39125 (N_39125,N_38821,N_38918);
xor U39126 (N_39126,N_38926,N_38845);
or U39127 (N_39127,N_38880,N_38831);
nand U39128 (N_39128,N_38987,N_38936);
or U39129 (N_39129,N_38870,N_38794);
xnor U39130 (N_39130,N_38931,N_38829);
or U39131 (N_39131,N_38787,N_38837);
or U39132 (N_39132,N_38941,N_38998);
or U39133 (N_39133,N_38991,N_38994);
nor U39134 (N_39134,N_38869,N_38862);
or U39135 (N_39135,N_38951,N_38787);
xor U39136 (N_39136,N_38760,N_38777);
and U39137 (N_39137,N_38971,N_38798);
nand U39138 (N_39138,N_38880,N_38877);
xor U39139 (N_39139,N_38959,N_38990);
nor U39140 (N_39140,N_38932,N_38974);
nor U39141 (N_39141,N_38953,N_38971);
or U39142 (N_39142,N_38848,N_38842);
nand U39143 (N_39143,N_38946,N_38759);
nand U39144 (N_39144,N_38963,N_38927);
and U39145 (N_39145,N_38954,N_38946);
and U39146 (N_39146,N_38897,N_38815);
nor U39147 (N_39147,N_38787,N_38851);
nand U39148 (N_39148,N_38960,N_38914);
or U39149 (N_39149,N_38821,N_38894);
or U39150 (N_39150,N_38876,N_38946);
and U39151 (N_39151,N_38840,N_38830);
nand U39152 (N_39152,N_38862,N_38912);
and U39153 (N_39153,N_38861,N_38966);
or U39154 (N_39154,N_38874,N_38836);
nor U39155 (N_39155,N_38974,N_38966);
and U39156 (N_39156,N_38915,N_38974);
and U39157 (N_39157,N_38863,N_38811);
nand U39158 (N_39158,N_38787,N_38899);
nor U39159 (N_39159,N_38900,N_38897);
nand U39160 (N_39160,N_38756,N_38903);
xnor U39161 (N_39161,N_38771,N_38994);
and U39162 (N_39162,N_38793,N_38881);
xor U39163 (N_39163,N_38819,N_38975);
and U39164 (N_39164,N_38885,N_38948);
or U39165 (N_39165,N_38833,N_38832);
nor U39166 (N_39166,N_38969,N_38799);
nand U39167 (N_39167,N_38917,N_38907);
or U39168 (N_39168,N_38849,N_38926);
and U39169 (N_39169,N_38932,N_38981);
or U39170 (N_39170,N_38964,N_38792);
xor U39171 (N_39171,N_38758,N_38944);
nor U39172 (N_39172,N_38801,N_38950);
xnor U39173 (N_39173,N_38784,N_38962);
xnor U39174 (N_39174,N_38860,N_38787);
xor U39175 (N_39175,N_38776,N_38771);
nand U39176 (N_39176,N_38926,N_38865);
xnor U39177 (N_39177,N_38781,N_38956);
and U39178 (N_39178,N_38815,N_38812);
and U39179 (N_39179,N_38882,N_38857);
and U39180 (N_39180,N_38865,N_38832);
xor U39181 (N_39181,N_38775,N_38911);
xor U39182 (N_39182,N_38972,N_38797);
and U39183 (N_39183,N_38820,N_38960);
xnor U39184 (N_39184,N_38812,N_38782);
xnor U39185 (N_39185,N_38815,N_38941);
nor U39186 (N_39186,N_38968,N_38762);
nand U39187 (N_39187,N_38940,N_38850);
nor U39188 (N_39188,N_38772,N_38978);
nand U39189 (N_39189,N_38891,N_38983);
or U39190 (N_39190,N_38817,N_38837);
nor U39191 (N_39191,N_38809,N_38833);
and U39192 (N_39192,N_38953,N_38773);
or U39193 (N_39193,N_38887,N_38844);
nand U39194 (N_39194,N_38805,N_38927);
nand U39195 (N_39195,N_38834,N_38986);
nor U39196 (N_39196,N_38952,N_38783);
nor U39197 (N_39197,N_38899,N_38818);
nor U39198 (N_39198,N_38869,N_38945);
and U39199 (N_39199,N_38879,N_38752);
nand U39200 (N_39200,N_38808,N_38879);
and U39201 (N_39201,N_38979,N_38965);
nand U39202 (N_39202,N_38997,N_38774);
nor U39203 (N_39203,N_38985,N_38975);
nand U39204 (N_39204,N_38901,N_38789);
and U39205 (N_39205,N_38884,N_38774);
xor U39206 (N_39206,N_38906,N_38808);
and U39207 (N_39207,N_38765,N_38797);
nand U39208 (N_39208,N_38798,N_38929);
nor U39209 (N_39209,N_38973,N_38799);
or U39210 (N_39210,N_38929,N_38946);
or U39211 (N_39211,N_38889,N_38942);
and U39212 (N_39212,N_38965,N_38964);
xor U39213 (N_39213,N_38846,N_38990);
nand U39214 (N_39214,N_38873,N_38869);
nand U39215 (N_39215,N_38969,N_38789);
nor U39216 (N_39216,N_38955,N_38789);
xnor U39217 (N_39217,N_38811,N_38945);
or U39218 (N_39218,N_38951,N_38805);
xnor U39219 (N_39219,N_38791,N_38752);
or U39220 (N_39220,N_38928,N_38890);
and U39221 (N_39221,N_38889,N_38946);
and U39222 (N_39222,N_38892,N_38796);
nand U39223 (N_39223,N_38895,N_38963);
xnor U39224 (N_39224,N_38845,N_38951);
xnor U39225 (N_39225,N_38790,N_38869);
or U39226 (N_39226,N_38929,N_38970);
and U39227 (N_39227,N_38924,N_38889);
nand U39228 (N_39228,N_38830,N_38979);
nor U39229 (N_39229,N_38765,N_38752);
nand U39230 (N_39230,N_38974,N_38965);
xnor U39231 (N_39231,N_38807,N_38812);
nand U39232 (N_39232,N_38987,N_38828);
nand U39233 (N_39233,N_38755,N_38944);
nand U39234 (N_39234,N_38844,N_38929);
or U39235 (N_39235,N_38933,N_38832);
nor U39236 (N_39236,N_38769,N_38801);
and U39237 (N_39237,N_38844,N_38779);
xor U39238 (N_39238,N_38840,N_38913);
xnor U39239 (N_39239,N_38758,N_38891);
or U39240 (N_39240,N_38944,N_38840);
and U39241 (N_39241,N_38974,N_38811);
and U39242 (N_39242,N_38974,N_38817);
xnor U39243 (N_39243,N_38980,N_38770);
and U39244 (N_39244,N_38962,N_38953);
xor U39245 (N_39245,N_38995,N_38868);
xnor U39246 (N_39246,N_38992,N_38842);
and U39247 (N_39247,N_38851,N_38801);
nor U39248 (N_39248,N_38957,N_38781);
xor U39249 (N_39249,N_38952,N_38960);
nor U39250 (N_39250,N_39012,N_39236);
nor U39251 (N_39251,N_39050,N_39185);
xnor U39252 (N_39252,N_39026,N_39029);
xor U39253 (N_39253,N_39062,N_39066);
and U39254 (N_39254,N_39244,N_39205);
or U39255 (N_39255,N_39229,N_39221);
or U39256 (N_39256,N_39051,N_39176);
or U39257 (N_39257,N_39111,N_39109);
nor U39258 (N_39258,N_39117,N_39160);
or U39259 (N_39259,N_39175,N_39241);
nand U39260 (N_39260,N_39195,N_39211);
and U39261 (N_39261,N_39219,N_39135);
xor U39262 (N_39262,N_39093,N_39094);
or U39263 (N_39263,N_39122,N_39120);
nand U39264 (N_39264,N_39082,N_39155);
and U39265 (N_39265,N_39202,N_39140);
or U39266 (N_39266,N_39225,N_39248);
xor U39267 (N_39267,N_39031,N_39194);
nand U39268 (N_39268,N_39000,N_39055);
xnor U39269 (N_39269,N_39075,N_39247);
or U39270 (N_39270,N_39243,N_39069);
nor U39271 (N_39271,N_39056,N_39071);
nand U39272 (N_39272,N_39072,N_39209);
nand U39273 (N_39273,N_39080,N_39037);
and U39274 (N_39274,N_39025,N_39108);
nand U39275 (N_39275,N_39131,N_39213);
xor U39276 (N_39276,N_39147,N_39145);
nand U39277 (N_39277,N_39114,N_39181);
nand U39278 (N_39278,N_39092,N_39127);
or U39279 (N_39279,N_39052,N_39138);
nand U39280 (N_39280,N_39076,N_39121);
xor U39281 (N_39281,N_39146,N_39234);
or U39282 (N_39282,N_39226,N_39227);
and U39283 (N_39283,N_39223,N_39218);
xor U39284 (N_39284,N_39063,N_39021);
nand U39285 (N_39285,N_39184,N_39079);
xnor U39286 (N_39286,N_39173,N_39210);
and U39287 (N_39287,N_39235,N_39123);
or U39288 (N_39288,N_39134,N_39097);
xnor U39289 (N_39289,N_39030,N_39095);
nor U39290 (N_39290,N_39084,N_39033);
nor U39291 (N_39291,N_39053,N_39070);
nor U39292 (N_39292,N_39208,N_39113);
or U39293 (N_39293,N_39083,N_39203);
or U39294 (N_39294,N_39158,N_39230);
nor U39295 (N_39295,N_39228,N_39174);
or U39296 (N_39296,N_39154,N_39179);
nor U39297 (N_39297,N_39129,N_39143);
nor U39298 (N_39298,N_39006,N_39172);
nor U39299 (N_39299,N_39077,N_39190);
nand U39300 (N_39300,N_39011,N_39239);
and U39301 (N_39301,N_39100,N_39180);
nor U39302 (N_39302,N_39197,N_39168);
nor U39303 (N_39303,N_39233,N_39152);
xor U39304 (N_39304,N_39048,N_39240);
nor U39305 (N_39305,N_39187,N_39073);
nand U39306 (N_39306,N_39047,N_39201);
or U39307 (N_39307,N_39137,N_39162);
nor U39308 (N_39308,N_39017,N_39101);
nor U39309 (N_39309,N_39098,N_39032);
or U39310 (N_39310,N_39115,N_39212);
nand U39311 (N_39311,N_39167,N_39039);
and U39312 (N_39312,N_39040,N_39242);
or U39313 (N_39313,N_39238,N_39118);
nand U39314 (N_39314,N_39088,N_39119);
and U39315 (N_39315,N_39237,N_39215);
nor U39316 (N_39316,N_39159,N_39018);
and U39317 (N_39317,N_39136,N_39177);
nand U39318 (N_39318,N_39058,N_39204);
nand U39319 (N_39319,N_39022,N_39103);
xor U39320 (N_39320,N_39151,N_39206);
xnor U39321 (N_39321,N_39186,N_39081);
and U39322 (N_39322,N_39045,N_39074);
xnor U39323 (N_39323,N_39170,N_39182);
or U39324 (N_39324,N_39112,N_39245);
nand U39325 (N_39325,N_39106,N_39096);
nor U39326 (N_39326,N_39016,N_39183);
or U39327 (N_39327,N_39041,N_39157);
xor U39328 (N_39328,N_39007,N_39141);
or U39329 (N_39329,N_39023,N_39156);
nand U39330 (N_39330,N_39102,N_39067);
nand U39331 (N_39331,N_39060,N_39091);
xor U39332 (N_39332,N_39133,N_39222);
nand U39333 (N_39333,N_39144,N_39036);
nor U39334 (N_39334,N_39089,N_39028);
and U39335 (N_39335,N_39005,N_39132);
nand U39336 (N_39336,N_39246,N_39224);
xnor U39337 (N_39337,N_39207,N_39216);
nand U39338 (N_39338,N_39249,N_39148);
xor U39339 (N_39339,N_39150,N_39139);
and U39340 (N_39340,N_39065,N_39166);
and U39341 (N_39341,N_39232,N_39200);
nand U39342 (N_39342,N_39003,N_39038);
or U39343 (N_39343,N_39042,N_39199);
nand U39344 (N_39344,N_39149,N_39068);
or U39345 (N_39345,N_39087,N_39214);
and U39346 (N_39346,N_39116,N_39002);
nor U39347 (N_39347,N_39078,N_39220);
nand U39348 (N_39348,N_39191,N_39164);
xnor U39349 (N_39349,N_39128,N_39196);
nor U39350 (N_39350,N_39217,N_39090);
nand U39351 (N_39351,N_39044,N_39193);
and U39352 (N_39352,N_39189,N_39231);
and U39353 (N_39353,N_39171,N_39099);
nand U39354 (N_39354,N_39125,N_39054);
nor U39355 (N_39355,N_39130,N_39027);
xor U39356 (N_39356,N_39015,N_39059);
or U39357 (N_39357,N_39014,N_39165);
or U39358 (N_39358,N_39019,N_39064);
or U39359 (N_39359,N_39046,N_39009);
nor U39360 (N_39360,N_39142,N_39035);
or U39361 (N_39361,N_39169,N_39008);
xor U39362 (N_39362,N_39124,N_39163);
nor U39363 (N_39363,N_39104,N_39105);
nor U39364 (N_39364,N_39013,N_39192);
nor U39365 (N_39365,N_39198,N_39085);
or U39366 (N_39366,N_39153,N_39107);
nand U39367 (N_39367,N_39188,N_39061);
or U39368 (N_39368,N_39001,N_39126);
nor U39369 (N_39369,N_39161,N_39010);
and U39370 (N_39370,N_39024,N_39086);
or U39371 (N_39371,N_39178,N_39057);
nand U39372 (N_39372,N_39020,N_39034);
xor U39373 (N_39373,N_39004,N_39110);
nand U39374 (N_39374,N_39043,N_39049);
and U39375 (N_39375,N_39185,N_39047);
or U39376 (N_39376,N_39101,N_39027);
nor U39377 (N_39377,N_39174,N_39062);
and U39378 (N_39378,N_39137,N_39178);
or U39379 (N_39379,N_39101,N_39152);
and U39380 (N_39380,N_39128,N_39069);
xor U39381 (N_39381,N_39065,N_39180);
or U39382 (N_39382,N_39187,N_39139);
or U39383 (N_39383,N_39187,N_39075);
nand U39384 (N_39384,N_39164,N_39186);
nand U39385 (N_39385,N_39085,N_39148);
nand U39386 (N_39386,N_39159,N_39183);
and U39387 (N_39387,N_39110,N_39241);
or U39388 (N_39388,N_39153,N_39008);
nor U39389 (N_39389,N_39044,N_39210);
and U39390 (N_39390,N_39132,N_39208);
or U39391 (N_39391,N_39211,N_39171);
or U39392 (N_39392,N_39193,N_39155);
or U39393 (N_39393,N_39162,N_39141);
and U39394 (N_39394,N_39128,N_39006);
and U39395 (N_39395,N_39031,N_39075);
xor U39396 (N_39396,N_39095,N_39018);
nor U39397 (N_39397,N_39008,N_39233);
xnor U39398 (N_39398,N_39049,N_39106);
or U39399 (N_39399,N_39127,N_39045);
nor U39400 (N_39400,N_39146,N_39199);
xnor U39401 (N_39401,N_39122,N_39196);
nor U39402 (N_39402,N_39151,N_39168);
or U39403 (N_39403,N_39215,N_39117);
nand U39404 (N_39404,N_39156,N_39151);
and U39405 (N_39405,N_39042,N_39031);
nor U39406 (N_39406,N_39128,N_39082);
xor U39407 (N_39407,N_39103,N_39192);
nor U39408 (N_39408,N_39057,N_39028);
nor U39409 (N_39409,N_39107,N_39160);
and U39410 (N_39410,N_39228,N_39108);
and U39411 (N_39411,N_39169,N_39088);
and U39412 (N_39412,N_39134,N_39026);
or U39413 (N_39413,N_39001,N_39232);
and U39414 (N_39414,N_39002,N_39140);
nor U39415 (N_39415,N_39120,N_39082);
nor U39416 (N_39416,N_39130,N_39104);
nand U39417 (N_39417,N_39015,N_39102);
or U39418 (N_39418,N_39090,N_39144);
nand U39419 (N_39419,N_39155,N_39100);
xnor U39420 (N_39420,N_39034,N_39244);
nor U39421 (N_39421,N_39015,N_39184);
or U39422 (N_39422,N_39095,N_39091);
xor U39423 (N_39423,N_39237,N_39050);
nand U39424 (N_39424,N_39012,N_39111);
and U39425 (N_39425,N_39121,N_39053);
nor U39426 (N_39426,N_39188,N_39242);
xnor U39427 (N_39427,N_39007,N_39023);
and U39428 (N_39428,N_39229,N_39114);
or U39429 (N_39429,N_39021,N_39180);
and U39430 (N_39430,N_39028,N_39030);
nand U39431 (N_39431,N_39060,N_39220);
and U39432 (N_39432,N_39133,N_39121);
nand U39433 (N_39433,N_39191,N_39206);
and U39434 (N_39434,N_39214,N_39089);
nand U39435 (N_39435,N_39123,N_39173);
nand U39436 (N_39436,N_39162,N_39146);
nand U39437 (N_39437,N_39134,N_39090);
or U39438 (N_39438,N_39151,N_39136);
nand U39439 (N_39439,N_39149,N_39041);
or U39440 (N_39440,N_39055,N_39095);
xnor U39441 (N_39441,N_39106,N_39229);
xor U39442 (N_39442,N_39205,N_39001);
xnor U39443 (N_39443,N_39146,N_39211);
and U39444 (N_39444,N_39193,N_39177);
or U39445 (N_39445,N_39237,N_39156);
and U39446 (N_39446,N_39047,N_39238);
xor U39447 (N_39447,N_39216,N_39201);
and U39448 (N_39448,N_39231,N_39205);
and U39449 (N_39449,N_39072,N_39056);
and U39450 (N_39450,N_39120,N_39077);
and U39451 (N_39451,N_39107,N_39084);
and U39452 (N_39452,N_39098,N_39013);
or U39453 (N_39453,N_39099,N_39247);
nor U39454 (N_39454,N_39056,N_39204);
xor U39455 (N_39455,N_39215,N_39207);
nor U39456 (N_39456,N_39195,N_39008);
or U39457 (N_39457,N_39232,N_39122);
and U39458 (N_39458,N_39193,N_39165);
nor U39459 (N_39459,N_39013,N_39217);
nor U39460 (N_39460,N_39191,N_39013);
and U39461 (N_39461,N_39045,N_39024);
nor U39462 (N_39462,N_39197,N_39056);
or U39463 (N_39463,N_39220,N_39174);
nand U39464 (N_39464,N_39166,N_39101);
xnor U39465 (N_39465,N_39038,N_39034);
nor U39466 (N_39466,N_39095,N_39207);
nor U39467 (N_39467,N_39102,N_39092);
or U39468 (N_39468,N_39057,N_39005);
or U39469 (N_39469,N_39230,N_39118);
xnor U39470 (N_39470,N_39076,N_39004);
xnor U39471 (N_39471,N_39095,N_39099);
or U39472 (N_39472,N_39228,N_39072);
nor U39473 (N_39473,N_39017,N_39024);
and U39474 (N_39474,N_39121,N_39018);
and U39475 (N_39475,N_39122,N_39123);
and U39476 (N_39476,N_39042,N_39038);
nand U39477 (N_39477,N_39230,N_39085);
and U39478 (N_39478,N_39164,N_39090);
nand U39479 (N_39479,N_39188,N_39031);
nor U39480 (N_39480,N_39150,N_39186);
xnor U39481 (N_39481,N_39240,N_39112);
nor U39482 (N_39482,N_39089,N_39213);
or U39483 (N_39483,N_39083,N_39031);
and U39484 (N_39484,N_39103,N_39002);
nand U39485 (N_39485,N_39213,N_39214);
nand U39486 (N_39486,N_39162,N_39055);
nor U39487 (N_39487,N_39085,N_39131);
and U39488 (N_39488,N_39024,N_39191);
xor U39489 (N_39489,N_39124,N_39032);
and U39490 (N_39490,N_39075,N_39060);
or U39491 (N_39491,N_39198,N_39142);
nand U39492 (N_39492,N_39118,N_39175);
or U39493 (N_39493,N_39016,N_39131);
nand U39494 (N_39494,N_39210,N_39095);
or U39495 (N_39495,N_39199,N_39020);
and U39496 (N_39496,N_39220,N_39092);
or U39497 (N_39497,N_39119,N_39125);
xor U39498 (N_39498,N_39059,N_39182);
and U39499 (N_39499,N_39243,N_39147);
xor U39500 (N_39500,N_39274,N_39486);
nand U39501 (N_39501,N_39277,N_39356);
or U39502 (N_39502,N_39372,N_39320);
and U39503 (N_39503,N_39445,N_39290);
and U39504 (N_39504,N_39266,N_39301);
and U39505 (N_39505,N_39463,N_39349);
xor U39506 (N_39506,N_39352,N_39473);
xnor U39507 (N_39507,N_39279,N_39407);
or U39508 (N_39508,N_39458,N_39385);
xnor U39509 (N_39509,N_39316,N_39427);
nand U39510 (N_39510,N_39269,N_39467);
nor U39511 (N_39511,N_39362,N_39480);
nand U39512 (N_39512,N_39478,N_39404);
nand U39513 (N_39513,N_39449,N_39283);
or U39514 (N_39514,N_39295,N_39298);
nor U39515 (N_39515,N_39296,N_39465);
or U39516 (N_39516,N_39475,N_39488);
nand U39517 (N_39517,N_39387,N_39335);
or U39518 (N_39518,N_39430,N_39423);
or U39519 (N_39519,N_39306,N_39280);
xnor U39520 (N_39520,N_39257,N_39273);
xnor U39521 (N_39521,N_39307,N_39343);
or U39522 (N_39522,N_39326,N_39336);
xnor U39523 (N_39523,N_39381,N_39328);
nor U39524 (N_39524,N_39254,N_39284);
xor U39525 (N_39525,N_39443,N_39383);
nand U39526 (N_39526,N_39384,N_39302);
xor U39527 (N_39527,N_39308,N_39304);
nand U39528 (N_39528,N_39278,N_39339);
xnor U39529 (N_39529,N_39377,N_39294);
nand U39530 (N_39530,N_39378,N_39347);
or U39531 (N_39531,N_39426,N_39435);
and U39532 (N_39532,N_39361,N_39312);
nor U39533 (N_39533,N_39322,N_39442);
xnor U39534 (N_39534,N_39440,N_39363);
nand U39535 (N_39535,N_39332,N_39472);
nor U39536 (N_39536,N_39432,N_39348);
xor U39537 (N_39537,N_39371,N_39360);
or U39538 (N_39538,N_39380,N_39439);
or U39539 (N_39539,N_39495,N_39469);
nand U39540 (N_39540,N_39450,N_39271);
xnor U39541 (N_39541,N_39350,N_39479);
xor U39542 (N_39542,N_39405,N_39419);
nor U39543 (N_39543,N_39499,N_39261);
or U39544 (N_39544,N_39461,N_39497);
or U39545 (N_39545,N_39428,N_39493);
or U39546 (N_39546,N_39297,N_39263);
xnor U39547 (N_39547,N_39264,N_39325);
nor U39548 (N_39548,N_39323,N_39342);
nor U39549 (N_39549,N_39414,N_39351);
nand U39550 (N_39550,N_39396,N_39267);
nor U39551 (N_39551,N_39253,N_39487);
and U39552 (N_39552,N_39317,N_39401);
xnor U39553 (N_39553,N_39410,N_39305);
xnor U39554 (N_39554,N_39376,N_39291);
or U39555 (N_39555,N_39303,N_39327);
xor U39556 (N_39556,N_39481,N_39437);
or U39557 (N_39557,N_39455,N_39345);
and U39558 (N_39558,N_39477,N_39412);
xor U39559 (N_39559,N_39260,N_39468);
or U39560 (N_39560,N_39397,N_39282);
xnor U39561 (N_39561,N_39448,N_39338);
nor U39562 (N_39562,N_39454,N_39402);
nand U39563 (N_39563,N_39334,N_39357);
xor U39564 (N_39564,N_39466,N_39258);
or U39565 (N_39565,N_39460,N_39311);
and U39566 (N_39566,N_39337,N_39386);
nand U39567 (N_39567,N_39299,N_39379);
or U39568 (N_39568,N_39392,N_39256);
xor U39569 (N_39569,N_39318,N_39436);
xor U39570 (N_39570,N_39496,N_39276);
and U39571 (N_39571,N_39359,N_39259);
and U39572 (N_39572,N_39418,N_39413);
nor U39573 (N_39573,N_39369,N_39319);
xor U39574 (N_39574,N_39484,N_39354);
xor U39575 (N_39575,N_39353,N_39330);
xor U39576 (N_39576,N_39394,N_39453);
and U39577 (N_39577,N_39390,N_39382);
or U39578 (N_39578,N_39288,N_39364);
nand U39579 (N_39579,N_39417,N_39375);
nand U39580 (N_39580,N_39331,N_39292);
xor U39581 (N_39581,N_39321,N_39441);
nand U39582 (N_39582,N_39491,N_39416);
xor U39583 (N_39583,N_39400,N_39374);
or U39584 (N_39584,N_39447,N_39251);
or U39585 (N_39585,N_39340,N_39399);
nor U39586 (N_39586,N_39265,N_39389);
xnor U39587 (N_39587,N_39252,N_39411);
and U39588 (N_39588,N_39434,N_39422);
and U39589 (N_39589,N_39398,N_39485);
xor U39590 (N_39590,N_39293,N_39365);
nor U39591 (N_39591,N_39367,N_39474);
and U39592 (N_39592,N_39344,N_39470);
nor U39593 (N_39593,N_39281,N_39346);
and U39594 (N_39594,N_39368,N_39272);
nand U39595 (N_39595,N_39433,N_39415);
or U39596 (N_39596,N_39255,N_39395);
or U39597 (N_39597,N_39483,N_39373);
or U39598 (N_39598,N_39444,N_39341);
xnor U39599 (N_39599,N_39355,N_39489);
nor U39600 (N_39600,N_39388,N_39451);
and U39601 (N_39601,N_39498,N_39464);
nor U39602 (N_39602,N_39425,N_39366);
and U39603 (N_39603,N_39314,N_39268);
and U39604 (N_39604,N_39421,N_39424);
and U39605 (N_39605,N_39309,N_39494);
and U39606 (N_39606,N_39250,N_39408);
and U39607 (N_39607,N_39286,N_39270);
nor U39608 (N_39608,N_39429,N_39313);
and U39609 (N_39609,N_39446,N_39329);
and U39610 (N_39610,N_39452,N_39370);
nand U39611 (N_39611,N_39409,N_39403);
xnor U39612 (N_39612,N_39406,N_39324);
or U39613 (N_39613,N_39310,N_39476);
nand U39614 (N_39614,N_39420,N_39287);
nor U39615 (N_39615,N_39431,N_39482);
xor U39616 (N_39616,N_39275,N_39333);
nor U39617 (N_39617,N_39456,N_39300);
or U39618 (N_39618,N_39462,N_39285);
xor U39619 (N_39619,N_39471,N_39490);
nor U39620 (N_39620,N_39457,N_39492);
nor U39621 (N_39621,N_39393,N_39391);
nor U39622 (N_39622,N_39438,N_39262);
nand U39623 (N_39623,N_39315,N_39459);
xor U39624 (N_39624,N_39358,N_39289);
nand U39625 (N_39625,N_39336,N_39293);
xor U39626 (N_39626,N_39443,N_39251);
nand U39627 (N_39627,N_39486,N_39291);
and U39628 (N_39628,N_39383,N_39371);
and U39629 (N_39629,N_39447,N_39470);
or U39630 (N_39630,N_39359,N_39448);
nor U39631 (N_39631,N_39495,N_39462);
or U39632 (N_39632,N_39494,N_39481);
and U39633 (N_39633,N_39270,N_39298);
nor U39634 (N_39634,N_39335,N_39407);
and U39635 (N_39635,N_39436,N_39355);
and U39636 (N_39636,N_39311,N_39426);
or U39637 (N_39637,N_39283,N_39450);
nor U39638 (N_39638,N_39434,N_39383);
or U39639 (N_39639,N_39369,N_39370);
nor U39640 (N_39640,N_39454,N_39447);
nand U39641 (N_39641,N_39325,N_39309);
xor U39642 (N_39642,N_39412,N_39328);
nor U39643 (N_39643,N_39277,N_39304);
xnor U39644 (N_39644,N_39390,N_39283);
nor U39645 (N_39645,N_39263,N_39468);
nand U39646 (N_39646,N_39411,N_39350);
or U39647 (N_39647,N_39394,N_39329);
xor U39648 (N_39648,N_39335,N_39494);
and U39649 (N_39649,N_39363,N_39279);
and U39650 (N_39650,N_39284,N_39373);
nor U39651 (N_39651,N_39399,N_39298);
xnor U39652 (N_39652,N_39389,N_39313);
or U39653 (N_39653,N_39487,N_39471);
and U39654 (N_39654,N_39320,N_39393);
xnor U39655 (N_39655,N_39405,N_39295);
or U39656 (N_39656,N_39301,N_39330);
or U39657 (N_39657,N_39266,N_39367);
nand U39658 (N_39658,N_39430,N_39491);
nor U39659 (N_39659,N_39295,N_39383);
nor U39660 (N_39660,N_39309,N_39331);
and U39661 (N_39661,N_39428,N_39374);
and U39662 (N_39662,N_39373,N_39302);
or U39663 (N_39663,N_39422,N_39376);
xor U39664 (N_39664,N_39326,N_39494);
nor U39665 (N_39665,N_39449,N_39267);
nand U39666 (N_39666,N_39413,N_39268);
xor U39667 (N_39667,N_39286,N_39488);
or U39668 (N_39668,N_39356,N_39483);
or U39669 (N_39669,N_39273,N_39295);
nor U39670 (N_39670,N_39269,N_39386);
or U39671 (N_39671,N_39461,N_39479);
and U39672 (N_39672,N_39354,N_39439);
xor U39673 (N_39673,N_39366,N_39348);
nand U39674 (N_39674,N_39323,N_39386);
nand U39675 (N_39675,N_39498,N_39409);
and U39676 (N_39676,N_39397,N_39413);
nor U39677 (N_39677,N_39498,N_39446);
xor U39678 (N_39678,N_39456,N_39338);
and U39679 (N_39679,N_39331,N_39328);
xor U39680 (N_39680,N_39363,N_39307);
nand U39681 (N_39681,N_39387,N_39478);
xnor U39682 (N_39682,N_39386,N_39484);
and U39683 (N_39683,N_39477,N_39341);
nand U39684 (N_39684,N_39277,N_39376);
or U39685 (N_39685,N_39263,N_39331);
nor U39686 (N_39686,N_39319,N_39489);
xor U39687 (N_39687,N_39430,N_39397);
xnor U39688 (N_39688,N_39462,N_39305);
nor U39689 (N_39689,N_39415,N_39302);
or U39690 (N_39690,N_39485,N_39486);
xnor U39691 (N_39691,N_39306,N_39348);
and U39692 (N_39692,N_39438,N_39303);
nor U39693 (N_39693,N_39472,N_39268);
or U39694 (N_39694,N_39301,N_39458);
xnor U39695 (N_39695,N_39469,N_39267);
or U39696 (N_39696,N_39383,N_39426);
and U39697 (N_39697,N_39393,N_39343);
nor U39698 (N_39698,N_39494,N_39304);
xor U39699 (N_39699,N_39368,N_39348);
xnor U39700 (N_39700,N_39370,N_39281);
nor U39701 (N_39701,N_39427,N_39390);
nor U39702 (N_39702,N_39250,N_39476);
nand U39703 (N_39703,N_39460,N_39431);
or U39704 (N_39704,N_39363,N_39284);
and U39705 (N_39705,N_39335,N_39386);
nor U39706 (N_39706,N_39285,N_39304);
nor U39707 (N_39707,N_39443,N_39390);
xnor U39708 (N_39708,N_39493,N_39469);
nor U39709 (N_39709,N_39474,N_39380);
nand U39710 (N_39710,N_39421,N_39407);
xnor U39711 (N_39711,N_39471,N_39375);
or U39712 (N_39712,N_39261,N_39403);
nand U39713 (N_39713,N_39299,N_39436);
and U39714 (N_39714,N_39304,N_39363);
nor U39715 (N_39715,N_39441,N_39275);
nand U39716 (N_39716,N_39282,N_39313);
or U39717 (N_39717,N_39453,N_39297);
nand U39718 (N_39718,N_39424,N_39450);
nor U39719 (N_39719,N_39397,N_39327);
and U39720 (N_39720,N_39469,N_39382);
and U39721 (N_39721,N_39439,N_39339);
and U39722 (N_39722,N_39255,N_39477);
or U39723 (N_39723,N_39411,N_39444);
xnor U39724 (N_39724,N_39340,N_39289);
nor U39725 (N_39725,N_39460,N_39418);
nand U39726 (N_39726,N_39339,N_39491);
or U39727 (N_39727,N_39296,N_39313);
xor U39728 (N_39728,N_39337,N_39353);
xnor U39729 (N_39729,N_39280,N_39384);
and U39730 (N_39730,N_39467,N_39314);
or U39731 (N_39731,N_39346,N_39282);
or U39732 (N_39732,N_39402,N_39472);
and U39733 (N_39733,N_39468,N_39267);
and U39734 (N_39734,N_39401,N_39481);
nand U39735 (N_39735,N_39471,N_39330);
xnor U39736 (N_39736,N_39273,N_39318);
and U39737 (N_39737,N_39486,N_39292);
nand U39738 (N_39738,N_39399,N_39331);
nand U39739 (N_39739,N_39328,N_39428);
xor U39740 (N_39740,N_39438,N_39415);
nand U39741 (N_39741,N_39348,N_39250);
and U39742 (N_39742,N_39283,N_39486);
or U39743 (N_39743,N_39373,N_39475);
nor U39744 (N_39744,N_39364,N_39418);
nor U39745 (N_39745,N_39266,N_39283);
xnor U39746 (N_39746,N_39307,N_39369);
xor U39747 (N_39747,N_39262,N_39496);
and U39748 (N_39748,N_39257,N_39398);
nand U39749 (N_39749,N_39498,N_39482);
xor U39750 (N_39750,N_39583,N_39568);
xor U39751 (N_39751,N_39520,N_39619);
xor U39752 (N_39752,N_39611,N_39692);
or U39753 (N_39753,N_39596,N_39645);
and U39754 (N_39754,N_39690,N_39601);
xnor U39755 (N_39755,N_39748,N_39639);
nand U39756 (N_39756,N_39537,N_39566);
or U39757 (N_39757,N_39512,N_39670);
and U39758 (N_39758,N_39637,N_39562);
xnor U39759 (N_39759,N_39703,N_39642);
or U39760 (N_39760,N_39713,N_39677);
xor U39761 (N_39761,N_39587,N_39501);
nand U39762 (N_39762,N_39660,N_39651);
nand U39763 (N_39763,N_39694,N_39631);
or U39764 (N_39764,N_39737,N_39648);
nor U39765 (N_39765,N_39618,N_39647);
or U39766 (N_39766,N_39653,N_39546);
nand U39767 (N_39767,N_39557,N_39600);
nand U39768 (N_39768,N_39593,N_39615);
nor U39769 (N_39769,N_39743,N_39712);
nand U39770 (N_39770,N_39742,N_39659);
nand U39771 (N_39771,N_39649,N_39612);
or U39772 (N_39772,N_39564,N_39630);
or U39773 (N_39773,N_39709,N_39716);
and U39774 (N_39774,N_39702,N_39578);
and U39775 (N_39775,N_39534,N_39706);
nand U39776 (N_39776,N_39538,N_39588);
and U39777 (N_39777,N_39582,N_39680);
nand U39778 (N_39778,N_39526,N_39589);
nor U39779 (N_39779,N_39700,N_39640);
or U39780 (N_39780,N_39745,N_39616);
nor U39781 (N_39781,N_39550,N_39540);
xor U39782 (N_39782,N_39511,N_39650);
or U39783 (N_39783,N_39524,N_39730);
or U39784 (N_39784,N_39559,N_39514);
or U39785 (N_39785,N_39608,N_39525);
nor U39786 (N_39786,N_39542,N_39580);
nand U39787 (N_39787,N_39641,N_39554);
nor U39788 (N_39788,N_39708,N_39747);
xnor U39789 (N_39789,N_39714,N_39543);
xor U39790 (N_39790,N_39688,N_39508);
xnor U39791 (N_39791,N_39729,N_39668);
nor U39792 (N_39792,N_39739,N_39719);
nor U39793 (N_39793,N_39691,N_39678);
and U39794 (N_39794,N_39516,N_39527);
xnor U39795 (N_39795,N_39685,N_39581);
nor U39796 (N_39796,N_39598,N_39698);
xor U39797 (N_39797,N_39635,N_39597);
and U39798 (N_39798,N_39561,N_39725);
nor U39799 (N_39799,N_39711,N_39614);
xor U39800 (N_39800,N_39654,N_39606);
nor U39801 (N_39801,N_39661,N_39515);
nor U39802 (N_39802,N_39664,N_39724);
nand U39803 (N_39803,N_39579,N_39658);
nand U39804 (N_39804,N_39662,N_39741);
or U39805 (N_39805,N_39684,N_39721);
xnor U39806 (N_39806,N_39699,N_39683);
nor U39807 (N_39807,N_39740,N_39715);
and U39808 (N_39808,N_39548,N_39536);
nor U39809 (N_39809,N_39657,N_39591);
nand U39810 (N_39810,N_39617,N_39517);
nor U39811 (N_39811,N_39652,N_39555);
xor U39812 (N_39812,N_39710,N_39529);
nor U39813 (N_39813,N_39633,N_39717);
nor U39814 (N_39814,N_39693,N_39528);
nand U39815 (N_39815,N_39585,N_39673);
and U39816 (N_39816,N_39560,N_39530);
nor U39817 (N_39817,N_39666,N_39682);
xnor U39818 (N_39818,N_39558,N_39569);
nand U39819 (N_39819,N_39502,N_39575);
and U39820 (N_39820,N_39628,N_39687);
xor U39821 (N_39821,N_39574,N_39704);
nor U39822 (N_39822,N_39571,N_39553);
nor U39823 (N_39823,N_39513,N_39733);
xnor U39824 (N_39824,N_39732,N_39636);
xnor U39825 (N_39825,N_39707,N_39663);
xnor U39826 (N_39826,N_39599,N_39720);
nand U39827 (N_39827,N_39624,N_39696);
xnor U39828 (N_39828,N_39686,N_39541);
nor U39829 (N_39829,N_39573,N_39665);
xor U39830 (N_39830,N_39738,N_39533);
xor U39831 (N_39831,N_39518,N_39552);
or U39832 (N_39832,N_39500,N_39504);
or U39833 (N_39833,N_39674,N_39605);
or U39834 (N_39834,N_39551,N_39695);
nor U39835 (N_39835,N_39697,N_39644);
or U39836 (N_39836,N_39655,N_39731);
nand U39837 (N_39837,N_39620,N_39531);
nand U39838 (N_39838,N_39602,N_39726);
xor U39839 (N_39839,N_39507,N_39592);
nor U39840 (N_39840,N_39625,N_39577);
nor U39841 (N_39841,N_39669,N_39643);
xor U39842 (N_39842,N_39728,N_39681);
xnor U39843 (N_39843,N_39632,N_39746);
nand U39844 (N_39844,N_39689,N_39595);
and U39845 (N_39845,N_39521,N_39638);
xnor U39846 (N_39846,N_39506,N_39672);
and U39847 (N_39847,N_39629,N_39532);
nand U39848 (N_39848,N_39545,N_39563);
or U39849 (N_39849,N_39572,N_39671);
and U39850 (N_39850,N_39609,N_39607);
nor U39851 (N_39851,N_39590,N_39544);
or U39852 (N_39852,N_39705,N_39621);
and U39853 (N_39853,N_39503,N_39679);
xor U39854 (N_39854,N_39567,N_39622);
and U39855 (N_39855,N_39556,N_39734);
nor U39856 (N_39856,N_39736,N_39610);
and U39857 (N_39857,N_39547,N_39667);
xnor U39858 (N_39858,N_39675,N_39509);
and U39859 (N_39859,N_39718,N_39701);
nor U39860 (N_39860,N_39505,N_39576);
and U39861 (N_39861,N_39510,N_39594);
and U39862 (N_39862,N_39570,N_39623);
and U39863 (N_39863,N_39519,N_39539);
nor U39864 (N_39864,N_39722,N_39646);
or U39865 (N_39865,N_39627,N_39603);
xor U39866 (N_39866,N_39735,N_39656);
xnor U39867 (N_39867,N_39613,N_39549);
nor U39868 (N_39868,N_39634,N_39523);
nand U39869 (N_39869,N_39744,N_39586);
nor U39870 (N_39870,N_39676,N_39727);
and U39871 (N_39871,N_39626,N_39723);
xnor U39872 (N_39872,N_39565,N_39522);
nor U39873 (N_39873,N_39535,N_39749);
nand U39874 (N_39874,N_39604,N_39584);
xor U39875 (N_39875,N_39562,N_39520);
and U39876 (N_39876,N_39674,N_39619);
and U39877 (N_39877,N_39743,N_39570);
or U39878 (N_39878,N_39513,N_39657);
nor U39879 (N_39879,N_39683,N_39703);
nor U39880 (N_39880,N_39606,N_39517);
nor U39881 (N_39881,N_39676,N_39586);
nand U39882 (N_39882,N_39717,N_39668);
nand U39883 (N_39883,N_39504,N_39694);
xor U39884 (N_39884,N_39615,N_39643);
and U39885 (N_39885,N_39532,N_39749);
or U39886 (N_39886,N_39502,N_39680);
xnor U39887 (N_39887,N_39632,N_39600);
nor U39888 (N_39888,N_39736,N_39716);
xor U39889 (N_39889,N_39703,N_39698);
nand U39890 (N_39890,N_39600,N_39563);
or U39891 (N_39891,N_39568,N_39632);
xor U39892 (N_39892,N_39500,N_39576);
and U39893 (N_39893,N_39701,N_39641);
and U39894 (N_39894,N_39716,N_39546);
and U39895 (N_39895,N_39683,N_39727);
nand U39896 (N_39896,N_39728,N_39651);
xor U39897 (N_39897,N_39743,N_39631);
or U39898 (N_39898,N_39577,N_39508);
or U39899 (N_39899,N_39556,N_39684);
xor U39900 (N_39900,N_39676,N_39592);
nand U39901 (N_39901,N_39596,N_39610);
nor U39902 (N_39902,N_39725,N_39522);
and U39903 (N_39903,N_39678,N_39739);
xnor U39904 (N_39904,N_39574,N_39741);
xor U39905 (N_39905,N_39567,N_39667);
nor U39906 (N_39906,N_39708,N_39605);
and U39907 (N_39907,N_39550,N_39514);
nand U39908 (N_39908,N_39666,N_39517);
or U39909 (N_39909,N_39543,N_39633);
nand U39910 (N_39910,N_39695,N_39562);
or U39911 (N_39911,N_39740,N_39612);
or U39912 (N_39912,N_39540,N_39697);
nand U39913 (N_39913,N_39690,N_39584);
and U39914 (N_39914,N_39500,N_39518);
xor U39915 (N_39915,N_39569,N_39617);
or U39916 (N_39916,N_39655,N_39537);
nand U39917 (N_39917,N_39682,N_39571);
xnor U39918 (N_39918,N_39732,N_39629);
or U39919 (N_39919,N_39513,N_39609);
or U39920 (N_39920,N_39646,N_39693);
or U39921 (N_39921,N_39686,N_39691);
nand U39922 (N_39922,N_39747,N_39501);
xor U39923 (N_39923,N_39677,N_39665);
and U39924 (N_39924,N_39541,N_39512);
xnor U39925 (N_39925,N_39591,N_39654);
and U39926 (N_39926,N_39728,N_39654);
xor U39927 (N_39927,N_39540,N_39533);
xor U39928 (N_39928,N_39508,N_39726);
or U39929 (N_39929,N_39614,N_39728);
nand U39930 (N_39930,N_39596,N_39733);
nor U39931 (N_39931,N_39541,N_39648);
nor U39932 (N_39932,N_39600,N_39514);
or U39933 (N_39933,N_39559,N_39616);
nand U39934 (N_39934,N_39541,N_39721);
xnor U39935 (N_39935,N_39527,N_39608);
nand U39936 (N_39936,N_39604,N_39653);
and U39937 (N_39937,N_39723,N_39596);
and U39938 (N_39938,N_39661,N_39574);
nor U39939 (N_39939,N_39651,N_39521);
and U39940 (N_39940,N_39565,N_39529);
or U39941 (N_39941,N_39658,N_39551);
nor U39942 (N_39942,N_39597,N_39560);
and U39943 (N_39943,N_39663,N_39617);
or U39944 (N_39944,N_39625,N_39736);
and U39945 (N_39945,N_39678,N_39567);
nand U39946 (N_39946,N_39739,N_39560);
xnor U39947 (N_39947,N_39565,N_39630);
nor U39948 (N_39948,N_39518,N_39557);
and U39949 (N_39949,N_39623,N_39739);
nor U39950 (N_39950,N_39581,N_39573);
or U39951 (N_39951,N_39539,N_39664);
nand U39952 (N_39952,N_39723,N_39528);
or U39953 (N_39953,N_39545,N_39590);
nor U39954 (N_39954,N_39545,N_39740);
xnor U39955 (N_39955,N_39616,N_39589);
or U39956 (N_39956,N_39554,N_39513);
and U39957 (N_39957,N_39693,N_39588);
and U39958 (N_39958,N_39640,N_39644);
xor U39959 (N_39959,N_39580,N_39521);
xnor U39960 (N_39960,N_39524,N_39621);
xor U39961 (N_39961,N_39685,N_39607);
nor U39962 (N_39962,N_39503,N_39586);
xnor U39963 (N_39963,N_39516,N_39709);
or U39964 (N_39964,N_39660,N_39511);
nand U39965 (N_39965,N_39655,N_39585);
xnor U39966 (N_39966,N_39551,N_39721);
nand U39967 (N_39967,N_39628,N_39643);
nor U39968 (N_39968,N_39602,N_39740);
nand U39969 (N_39969,N_39595,N_39545);
xor U39970 (N_39970,N_39651,N_39530);
and U39971 (N_39971,N_39665,N_39655);
nor U39972 (N_39972,N_39595,N_39588);
and U39973 (N_39973,N_39689,N_39698);
xnor U39974 (N_39974,N_39732,N_39549);
nor U39975 (N_39975,N_39733,N_39517);
nor U39976 (N_39976,N_39675,N_39528);
xnor U39977 (N_39977,N_39721,N_39574);
or U39978 (N_39978,N_39600,N_39671);
xor U39979 (N_39979,N_39726,N_39565);
or U39980 (N_39980,N_39662,N_39510);
or U39981 (N_39981,N_39743,N_39602);
nor U39982 (N_39982,N_39732,N_39628);
nor U39983 (N_39983,N_39692,N_39736);
nor U39984 (N_39984,N_39556,N_39736);
nand U39985 (N_39985,N_39749,N_39670);
or U39986 (N_39986,N_39575,N_39659);
or U39987 (N_39987,N_39690,N_39642);
nand U39988 (N_39988,N_39744,N_39515);
and U39989 (N_39989,N_39625,N_39678);
xor U39990 (N_39990,N_39721,N_39653);
or U39991 (N_39991,N_39658,N_39582);
and U39992 (N_39992,N_39701,N_39619);
nor U39993 (N_39993,N_39702,N_39539);
nor U39994 (N_39994,N_39652,N_39614);
xor U39995 (N_39995,N_39599,N_39688);
nor U39996 (N_39996,N_39709,N_39526);
nand U39997 (N_39997,N_39630,N_39663);
and U39998 (N_39998,N_39683,N_39720);
and U39999 (N_39999,N_39606,N_39551);
nor U40000 (N_40000,N_39831,N_39881);
nor U40001 (N_40001,N_39862,N_39990);
xnor U40002 (N_40002,N_39786,N_39766);
and U40003 (N_40003,N_39836,N_39888);
nand U40004 (N_40004,N_39972,N_39994);
or U40005 (N_40005,N_39984,N_39875);
xnor U40006 (N_40006,N_39856,N_39802);
and U40007 (N_40007,N_39872,N_39928);
nand U40008 (N_40008,N_39957,N_39828);
or U40009 (N_40009,N_39806,N_39937);
and U40010 (N_40010,N_39978,N_39807);
xnor U40011 (N_40011,N_39909,N_39868);
nand U40012 (N_40012,N_39827,N_39936);
and U40013 (N_40013,N_39846,N_39832);
or U40014 (N_40014,N_39764,N_39889);
nand U40015 (N_40015,N_39925,N_39753);
nand U40016 (N_40016,N_39910,N_39837);
or U40017 (N_40017,N_39991,N_39815);
nor U40018 (N_40018,N_39826,N_39800);
xor U40019 (N_40019,N_39897,N_39809);
xnor U40020 (N_40020,N_39901,N_39908);
nand U40021 (N_40021,N_39820,N_39964);
nand U40022 (N_40022,N_39911,N_39979);
xnor U40023 (N_40023,N_39933,N_39817);
xnor U40024 (N_40024,N_39920,N_39750);
and U40025 (N_40025,N_39969,N_39848);
nand U40026 (N_40026,N_39759,N_39976);
nand U40027 (N_40027,N_39918,N_39767);
nand U40028 (N_40028,N_39962,N_39842);
nand U40029 (N_40029,N_39961,N_39829);
and U40030 (N_40030,N_39801,N_39763);
nand U40031 (N_40031,N_39867,N_39954);
nand U40032 (N_40032,N_39851,N_39966);
xor U40033 (N_40033,N_39835,N_39812);
and U40034 (N_40034,N_39959,N_39768);
or U40035 (N_40035,N_39849,N_39886);
xor U40036 (N_40036,N_39915,N_39838);
or U40037 (N_40037,N_39900,N_39895);
xor U40038 (N_40038,N_39956,N_39960);
nor U40039 (N_40039,N_39791,N_39923);
and U40040 (N_40040,N_39771,N_39951);
nand U40041 (N_40041,N_39993,N_39916);
xnor U40042 (N_40042,N_39885,N_39874);
or U40043 (N_40043,N_39789,N_39762);
or U40044 (N_40044,N_39898,N_39891);
nor U40045 (N_40045,N_39782,N_39852);
nor U40046 (N_40046,N_39864,N_39769);
and U40047 (N_40047,N_39927,N_39830);
xnor U40048 (N_40048,N_39779,N_39955);
xor U40049 (N_40049,N_39825,N_39887);
and U40050 (N_40050,N_39879,N_39840);
xor U40051 (N_40051,N_39892,N_39822);
xnor U40052 (N_40052,N_39792,N_39989);
xnor U40053 (N_40053,N_39847,N_39761);
and U40054 (N_40054,N_39932,N_39788);
nand U40055 (N_40055,N_39783,N_39965);
nor U40056 (N_40056,N_39941,N_39947);
and U40057 (N_40057,N_39754,N_39811);
nand U40058 (N_40058,N_39839,N_39985);
or U40059 (N_40059,N_39902,N_39940);
xor U40060 (N_40060,N_39906,N_39859);
xnor U40061 (N_40061,N_39998,N_39796);
or U40062 (N_40062,N_39944,N_39958);
or U40063 (N_40063,N_39996,N_39913);
nand U40064 (N_40064,N_39883,N_39776);
nor U40065 (N_40065,N_39798,N_39905);
nand U40066 (N_40066,N_39751,N_39865);
and U40067 (N_40067,N_39884,N_39999);
nand U40068 (N_40068,N_39757,N_39890);
nand U40069 (N_40069,N_39992,N_39986);
and U40070 (N_40070,N_39995,N_39756);
xnor U40071 (N_40071,N_39950,N_39752);
or U40072 (N_40072,N_39912,N_39784);
nand U40073 (N_40073,N_39946,N_39758);
nor U40074 (N_40074,N_39870,N_39853);
nand U40075 (N_40075,N_39843,N_39882);
nand U40076 (N_40076,N_39949,N_39988);
or U40077 (N_40077,N_39975,N_39833);
xor U40078 (N_40078,N_39816,N_39777);
nor U40079 (N_40079,N_39795,N_39893);
and U40080 (N_40080,N_39952,N_39793);
and U40081 (N_40081,N_39805,N_39818);
or U40082 (N_40082,N_39931,N_39770);
nand U40083 (N_40083,N_39871,N_39861);
nand U40084 (N_40084,N_39904,N_39819);
or U40085 (N_40085,N_39866,N_39878);
or U40086 (N_40086,N_39930,N_39973);
and U40087 (N_40087,N_39857,N_39797);
xor U40088 (N_40088,N_39787,N_39813);
nand U40089 (N_40089,N_39987,N_39967);
and U40090 (N_40090,N_39997,N_39873);
and U40091 (N_40091,N_39983,N_39963);
and U40092 (N_40092,N_39773,N_39860);
nand U40093 (N_40093,N_39845,N_39760);
xor U40094 (N_40094,N_39968,N_39834);
nand U40095 (N_40095,N_39880,N_39917);
nor U40096 (N_40096,N_39799,N_39903);
nor U40097 (N_40097,N_39977,N_39844);
nor U40098 (N_40098,N_39877,N_39755);
nand U40099 (N_40099,N_39794,N_39803);
and U40100 (N_40100,N_39945,N_39971);
or U40101 (N_40101,N_39938,N_39953);
or U40102 (N_40102,N_39921,N_39785);
xor U40103 (N_40103,N_39778,N_39981);
nor U40104 (N_40104,N_39772,N_39854);
and U40105 (N_40105,N_39814,N_39922);
nor U40106 (N_40106,N_39855,N_39970);
nor U40107 (N_40107,N_39929,N_39980);
xnor U40108 (N_40108,N_39823,N_39924);
or U40109 (N_40109,N_39982,N_39943);
xnor U40110 (N_40110,N_39926,N_39869);
nand U40111 (N_40111,N_39858,N_39808);
nor U40112 (N_40112,N_39894,N_39781);
nor U40113 (N_40113,N_39935,N_39841);
or U40114 (N_40114,N_39765,N_39899);
and U40115 (N_40115,N_39790,N_39974);
or U40116 (N_40116,N_39780,N_39850);
xor U40117 (N_40117,N_39810,N_39804);
nor U40118 (N_40118,N_39896,N_39824);
xnor U40119 (N_40119,N_39919,N_39774);
nand U40120 (N_40120,N_39876,N_39863);
xor U40121 (N_40121,N_39907,N_39821);
and U40122 (N_40122,N_39939,N_39948);
nor U40123 (N_40123,N_39775,N_39942);
nor U40124 (N_40124,N_39934,N_39914);
nor U40125 (N_40125,N_39990,N_39936);
xnor U40126 (N_40126,N_39892,N_39888);
and U40127 (N_40127,N_39856,N_39903);
xor U40128 (N_40128,N_39788,N_39799);
nand U40129 (N_40129,N_39994,N_39921);
nor U40130 (N_40130,N_39979,N_39966);
or U40131 (N_40131,N_39979,N_39976);
xor U40132 (N_40132,N_39938,N_39811);
and U40133 (N_40133,N_39772,N_39984);
nor U40134 (N_40134,N_39975,N_39801);
nor U40135 (N_40135,N_39789,N_39787);
or U40136 (N_40136,N_39939,N_39917);
nand U40137 (N_40137,N_39944,N_39875);
xor U40138 (N_40138,N_39894,N_39836);
nor U40139 (N_40139,N_39993,N_39981);
xnor U40140 (N_40140,N_39944,N_39978);
and U40141 (N_40141,N_39885,N_39755);
or U40142 (N_40142,N_39781,N_39871);
or U40143 (N_40143,N_39867,N_39907);
and U40144 (N_40144,N_39753,N_39982);
nor U40145 (N_40145,N_39963,N_39938);
xor U40146 (N_40146,N_39924,N_39855);
or U40147 (N_40147,N_39855,N_39817);
and U40148 (N_40148,N_39784,N_39897);
and U40149 (N_40149,N_39938,N_39842);
nand U40150 (N_40150,N_39908,N_39999);
nand U40151 (N_40151,N_39800,N_39813);
xnor U40152 (N_40152,N_39859,N_39828);
nand U40153 (N_40153,N_39829,N_39967);
nor U40154 (N_40154,N_39827,N_39791);
and U40155 (N_40155,N_39984,N_39970);
xor U40156 (N_40156,N_39758,N_39816);
nor U40157 (N_40157,N_39875,N_39782);
xnor U40158 (N_40158,N_39996,N_39813);
and U40159 (N_40159,N_39901,N_39968);
and U40160 (N_40160,N_39877,N_39906);
nand U40161 (N_40161,N_39794,N_39828);
or U40162 (N_40162,N_39853,N_39829);
or U40163 (N_40163,N_39832,N_39977);
xor U40164 (N_40164,N_39940,N_39926);
and U40165 (N_40165,N_39760,N_39960);
or U40166 (N_40166,N_39995,N_39912);
nor U40167 (N_40167,N_39928,N_39788);
nand U40168 (N_40168,N_39921,N_39797);
xor U40169 (N_40169,N_39942,N_39869);
xnor U40170 (N_40170,N_39846,N_39813);
nor U40171 (N_40171,N_39841,N_39837);
nand U40172 (N_40172,N_39924,N_39893);
xnor U40173 (N_40173,N_39846,N_39988);
and U40174 (N_40174,N_39824,N_39987);
nand U40175 (N_40175,N_39941,N_39991);
nor U40176 (N_40176,N_39926,N_39909);
or U40177 (N_40177,N_39791,N_39759);
and U40178 (N_40178,N_39966,N_39985);
or U40179 (N_40179,N_39839,N_39794);
and U40180 (N_40180,N_39813,N_39878);
or U40181 (N_40181,N_39879,N_39850);
nor U40182 (N_40182,N_39924,N_39828);
nand U40183 (N_40183,N_39775,N_39861);
xor U40184 (N_40184,N_39957,N_39959);
nand U40185 (N_40185,N_39962,N_39816);
nand U40186 (N_40186,N_39894,N_39803);
and U40187 (N_40187,N_39843,N_39836);
or U40188 (N_40188,N_39822,N_39979);
or U40189 (N_40189,N_39956,N_39839);
and U40190 (N_40190,N_39905,N_39878);
and U40191 (N_40191,N_39978,N_39885);
or U40192 (N_40192,N_39965,N_39921);
xnor U40193 (N_40193,N_39760,N_39962);
nand U40194 (N_40194,N_39967,N_39953);
xor U40195 (N_40195,N_39993,N_39989);
nor U40196 (N_40196,N_39865,N_39821);
and U40197 (N_40197,N_39818,N_39769);
or U40198 (N_40198,N_39781,N_39788);
nand U40199 (N_40199,N_39811,N_39996);
and U40200 (N_40200,N_39769,N_39985);
nand U40201 (N_40201,N_39770,N_39951);
or U40202 (N_40202,N_39857,N_39784);
nand U40203 (N_40203,N_39898,N_39928);
xnor U40204 (N_40204,N_39910,N_39789);
nor U40205 (N_40205,N_39799,N_39900);
nor U40206 (N_40206,N_39937,N_39992);
nand U40207 (N_40207,N_39786,N_39894);
or U40208 (N_40208,N_39937,N_39826);
or U40209 (N_40209,N_39762,N_39770);
nand U40210 (N_40210,N_39776,N_39938);
nand U40211 (N_40211,N_39759,N_39963);
nand U40212 (N_40212,N_39895,N_39976);
nor U40213 (N_40213,N_39997,N_39805);
nor U40214 (N_40214,N_39762,N_39899);
nand U40215 (N_40215,N_39762,N_39869);
or U40216 (N_40216,N_39754,N_39910);
nand U40217 (N_40217,N_39758,N_39783);
or U40218 (N_40218,N_39868,N_39871);
or U40219 (N_40219,N_39756,N_39994);
xnor U40220 (N_40220,N_39962,N_39858);
or U40221 (N_40221,N_39881,N_39782);
nand U40222 (N_40222,N_39821,N_39804);
xor U40223 (N_40223,N_39905,N_39853);
nor U40224 (N_40224,N_39889,N_39755);
or U40225 (N_40225,N_39962,N_39825);
nand U40226 (N_40226,N_39958,N_39987);
or U40227 (N_40227,N_39751,N_39894);
xnor U40228 (N_40228,N_39763,N_39933);
nand U40229 (N_40229,N_39830,N_39793);
or U40230 (N_40230,N_39836,N_39778);
nand U40231 (N_40231,N_39982,N_39969);
xnor U40232 (N_40232,N_39857,N_39887);
xnor U40233 (N_40233,N_39784,N_39898);
or U40234 (N_40234,N_39951,N_39806);
nand U40235 (N_40235,N_39876,N_39799);
or U40236 (N_40236,N_39753,N_39957);
nand U40237 (N_40237,N_39916,N_39792);
nor U40238 (N_40238,N_39765,N_39799);
or U40239 (N_40239,N_39951,N_39970);
nand U40240 (N_40240,N_39961,N_39962);
xnor U40241 (N_40241,N_39975,N_39852);
nand U40242 (N_40242,N_39885,N_39768);
xnor U40243 (N_40243,N_39815,N_39859);
nor U40244 (N_40244,N_39914,N_39779);
nor U40245 (N_40245,N_39990,N_39901);
nand U40246 (N_40246,N_39938,N_39851);
or U40247 (N_40247,N_39859,N_39998);
nor U40248 (N_40248,N_39938,N_39861);
or U40249 (N_40249,N_39755,N_39855);
xor U40250 (N_40250,N_40042,N_40143);
xnor U40251 (N_40251,N_40191,N_40081);
and U40252 (N_40252,N_40128,N_40225);
and U40253 (N_40253,N_40233,N_40246);
nor U40254 (N_40254,N_40073,N_40004);
and U40255 (N_40255,N_40072,N_40240);
xor U40256 (N_40256,N_40175,N_40034);
nor U40257 (N_40257,N_40053,N_40141);
and U40258 (N_40258,N_40119,N_40161);
nor U40259 (N_40259,N_40186,N_40005);
nand U40260 (N_40260,N_40193,N_40060);
and U40261 (N_40261,N_40015,N_40234);
nand U40262 (N_40262,N_40007,N_40102);
or U40263 (N_40263,N_40242,N_40174);
or U40264 (N_40264,N_40021,N_40192);
and U40265 (N_40265,N_40054,N_40245);
xnor U40266 (N_40266,N_40076,N_40033);
or U40267 (N_40267,N_40224,N_40115);
nand U40268 (N_40268,N_40069,N_40010);
xnor U40269 (N_40269,N_40217,N_40228);
nand U40270 (N_40270,N_40249,N_40159);
nor U40271 (N_40271,N_40212,N_40024);
xnor U40272 (N_40272,N_40083,N_40110);
nand U40273 (N_40273,N_40014,N_40122);
xnor U40274 (N_40274,N_40170,N_40205);
and U40275 (N_40275,N_40220,N_40094);
nor U40276 (N_40276,N_40079,N_40109);
nand U40277 (N_40277,N_40199,N_40000);
or U40278 (N_40278,N_40086,N_40112);
and U40279 (N_40279,N_40055,N_40006);
nor U40280 (N_40280,N_40058,N_40023);
xor U40281 (N_40281,N_40099,N_40230);
and U40282 (N_40282,N_40198,N_40158);
or U40283 (N_40283,N_40195,N_40064);
nor U40284 (N_40284,N_40134,N_40100);
nor U40285 (N_40285,N_40116,N_40168);
and U40286 (N_40286,N_40190,N_40239);
or U40287 (N_40287,N_40038,N_40120);
or U40288 (N_40288,N_40148,N_40088);
nor U40289 (N_40289,N_40160,N_40065);
and U40290 (N_40290,N_40129,N_40169);
or U40291 (N_40291,N_40171,N_40046);
xor U40292 (N_40292,N_40057,N_40176);
xor U40293 (N_40293,N_40203,N_40036);
xor U40294 (N_40294,N_40179,N_40236);
xnor U40295 (N_40295,N_40151,N_40130);
or U40296 (N_40296,N_40216,N_40178);
xnor U40297 (N_40297,N_40135,N_40196);
or U40298 (N_40298,N_40009,N_40067);
and U40299 (N_40299,N_40043,N_40020);
nor U40300 (N_40300,N_40243,N_40184);
nor U40301 (N_40301,N_40204,N_40104);
nor U40302 (N_40302,N_40238,N_40050);
nor U40303 (N_40303,N_40044,N_40103);
or U40304 (N_40304,N_40030,N_40101);
nor U40305 (N_40305,N_40145,N_40215);
nand U40306 (N_40306,N_40183,N_40019);
and U40307 (N_40307,N_40098,N_40227);
nand U40308 (N_40308,N_40062,N_40095);
and U40309 (N_40309,N_40127,N_40206);
and U40310 (N_40310,N_40146,N_40113);
and U40311 (N_40311,N_40092,N_40096);
nand U40312 (N_40312,N_40185,N_40026);
and U40313 (N_40313,N_40084,N_40002);
or U40314 (N_40314,N_40016,N_40142);
nand U40315 (N_40315,N_40022,N_40211);
xnor U40316 (N_40316,N_40068,N_40149);
or U40317 (N_40317,N_40025,N_40125);
nand U40318 (N_40318,N_40162,N_40197);
xor U40319 (N_40319,N_40231,N_40241);
or U40320 (N_40320,N_40049,N_40153);
nor U40321 (N_40321,N_40133,N_40139);
or U40322 (N_40322,N_40035,N_40126);
nand U40323 (N_40323,N_40087,N_40173);
nand U40324 (N_40324,N_40226,N_40163);
or U40325 (N_40325,N_40031,N_40167);
and U40326 (N_40326,N_40201,N_40182);
nor U40327 (N_40327,N_40027,N_40066);
nor U40328 (N_40328,N_40123,N_40117);
nor U40329 (N_40329,N_40164,N_40091);
or U40330 (N_40330,N_40180,N_40047);
nand U40331 (N_40331,N_40029,N_40032);
and U40332 (N_40332,N_40045,N_40028);
xnor U40333 (N_40333,N_40235,N_40166);
or U40334 (N_40334,N_40012,N_40085);
xnor U40335 (N_40335,N_40209,N_40082);
nand U40336 (N_40336,N_40165,N_40075);
nor U40337 (N_40337,N_40107,N_40132);
xnor U40338 (N_40338,N_40189,N_40208);
xor U40339 (N_40339,N_40063,N_40070);
nor U40340 (N_40340,N_40061,N_40210);
xnor U40341 (N_40341,N_40011,N_40071);
or U40342 (N_40342,N_40108,N_40156);
and U40343 (N_40343,N_40232,N_40001);
nor U40344 (N_40344,N_40188,N_40200);
or U40345 (N_40345,N_40118,N_40137);
and U40346 (N_40346,N_40114,N_40041);
nor U40347 (N_40347,N_40213,N_40140);
xor U40348 (N_40348,N_40147,N_40177);
xor U40349 (N_40349,N_40039,N_40124);
and U40350 (N_40350,N_40152,N_40078);
nand U40351 (N_40351,N_40157,N_40051);
nor U40352 (N_40352,N_40222,N_40077);
nor U40353 (N_40353,N_40121,N_40154);
xnor U40354 (N_40354,N_40187,N_40052);
xor U40355 (N_40355,N_40181,N_40089);
nand U40356 (N_40356,N_40138,N_40248);
and U40357 (N_40357,N_40144,N_40194);
and U40358 (N_40358,N_40093,N_40008);
nand U40359 (N_40359,N_40247,N_40131);
nand U40360 (N_40360,N_40090,N_40003);
xor U40361 (N_40361,N_40056,N_40223);
and U40362 (N_40362,N_40105,N_40037);
or U40363 (N_40363,N_40111,N_40155);
or U40364 (N_40364,N_40136,N_40244);
xor U40365 (N_40365,N_40080,N_40218);
and U40366 (N_40366,N_40207,N_40214);
xnor U40367 (N_40367,N_40040,N_40202);
nand U40368 (N_40368,N_40172,N_40018);
and U40369 (N_40369,N_40074,N_40150);
or U40370 (N_40370,N_40017,N_40097);
nand U40371 (N_40371,N_40219,N_40237);
or U40372 (N_40372,N_40013,N_40048);
and U40373 (N_40373,N_40221,N_40059);
nor U40374 (N_40374,N_40106,N_40229);
or U40375 (N_40375,N_40207,N_40151);
nand U40376 (N_40376,N_40192,N_40042);
xor U40377 (N_40377,N_40083,N_40202);
or U40378 (N_40378,N_40206,N_40018);
and U40379 (N_40379,N_40180,N_40088);
and U40380 (N_40380,N_40237,N_40194);
nand U40381 (N_40381,N_40236,N_40079);
nand U40382 (N_40382,N_40158,N_40149);
or U40383 (N_40383,N_40230,N_40175);
nand U40384 (N_40384,N_40071,N_40155);
nand U40385 (N_40385,N_40118,N_40114);
nor U40386 (N_40386,N_40001,N_40220);
or U40387 (N_40387,N_40215,N_40225);
nor U40388 (N_40388,N_40037,N_40117);
xor U40389 (N_40389,N_40198,N_40107);
and U40390 (N_40390,N_40024,N_40242);
xnor U40391 (N_40391,N_40218,N_40060);
nand U40392 (N_40392,N_40208,N_40183);
nor U40393 (N_40393,N_40202,N_40041);
nor U40394 (N_40394,N_40033,N_40168);
xor U40395 (N_40395,N_40110,N_40167);
and U40396 (N_40396,N_40063,N_40036);
or U40397 (N_40397,N_40087,N_40032);
xnor U40398 (N_40398,N_40181,N_40108);
nor U40399 (N_40399,N_40233,N_40048);
nor U40400 (N_40400,N_40060,N_40189);
nand U40401 (N_40401,N_40106,N_40020);
xor U40402 (N_40402,N_40150,N_40089);
xor U40403 (N_40403,N_40042,N_40141);
xnor U40404 (N_40404,N_40167,N_40125);
and U40405 (N_40405,N_40003,N_40014);
nand U40406 (N_40406,N_40128,N_40141);
nand U40407 (N_40407,N_40184,N_40131);
nor U40408 (N_40408,N_40159,N_40106);
nand U40409 (N_40409,N_40076,N_40082);
nor U40410 (N_40410,N_40141,N_40107);
or U40411 (N_40411,N_40170,N_40174);
nand U40412 (N_40412,N_40237,N_40066);
nor U40413 (N_40413,N_40165,N_40017);
or U40414 (N_40414,N_40097,N_40015);
nand U40415 (N_40415,N_40060,N_40207);
and U40416 (N_40416,N_40238,N_40152);
or U40417 (N_40417,N_40204,N_40116);
and U40418 (N_40418,N_40009,N_40106);
and U40419 (N_40419,N_40034,N_40193);
or U40420 (N_40420,N_40212,N_40136);
or U40421 (N_40421,N_40121,N_40026);
nor U40422 (N_40422,N_40037,N_40120);
nor U40423 (N_40423,N_40060,N_40127);
or U40424 (N_40424,N_40011,N_40109);
nand U40425 (N_40425,N_40020,N_40014);
xnor U40426 (N_40426,N_40202,N_40197);
nand U40427 (N_40427,N_40244,N_40236);
and U40428 (N_40428,N_40062,N_40217);
xnor U40429 (N_40429,N_40011,N_40199);
nor U40430 (N_40430,N_40199,N_40248);
nand U40431 (N_40431,N_40014,N_40202);
or U40432 (N_40432,N_40194,N_40136);
and U40433 (N_40433,N_40028,N_40061);
nor U40434 (N_40434,N_40245,N_40065);
xnor U40435 (N_40435,N_40222,N_40133);
and U40436 (N_40436,N_40033,N_40165);
nand U40437 (N_40437,N_40138,N_40219);
and U40438 (N_40438,N_40063,N_40003);
and U40439 (N_40439,N_40007,N_40103);
nor U40440 (N_40440,N_40046,N_40123);
and U40441 (N_40441,N_40109,N_40144);
nor U40442 (N_40442,N_40231,N_40074);
nor U40443 (N_40443,N_40031,N_40084);
nor U40444 (N_40444,N_40098,N_40044);
and U40445 (N_40445,N_40235,N_40121);
xnor U40446 (N_40446,N_40125,N_40185);
or U40447 (N_40447,N_40147,N_40098);
xor U40448 (N_40448,N_40244,N_40086);
nand U40449 (N_40449,N_40222,N_40042);
or U40450 (N_40450,N_40005,N_40077);
xor U40451 (N_40451,N_40110,N_40128);
nand U40452 (N_40452,N_40058,N_40224);
nand U40453 (N_40453,N_40205,N_40228);
nand U40454 (N_40454,N_40006,N_40010);
or U40455 (N_40455,N_40217,N_40097);
and U40456 (N_40456,N_40000,N_40070);
nor U40457 (N_40457,N_40044,N_40231);
xor U40458 (N_40458,N_40082,N_40112);
xor U40459 (N_40459,N_40244,N_40150);
and U40460 (N_40460,N_40170,N_40046);
nor U40461 (N_40461,N_40103,N_40150);
nand U40462 (N_40462,N_40223,N_40049);
or U40463 (N_40463,N_40038,N_40128);
xor U40464 (N_40464,N_40244,N_40212);
or U40465 (N_40465,N_40147,N_40236);
nand U40466 (N_40466,N_40213,N_40235);
xnor U40467 (N_40467,N_40122,N_40189);
nor U40468 (N_40468,N_40142,N_40080);
xnor U40469 (N_40469,N_40077,N_40217);
nand U40470 (N_40470,N_40000,N_40187);
nand U40471 (N_40471,N_40041,N_40185);
nor U40472 (N_40472,N_40158,N_40058);
xnor U40473 (N_40473,N_40049,N_40245);
xnor U40474 (N_40474,N_40209,N_40031);
and U40475 (N_40475,N_40018,N_40061);
nand U40476 (N_40476,N_40224,N_40178);
xor U40477 (N_40477,N_40026,N_40113);
xor U40478 (N_40478,N_40018,N_40193);
xnor U40479 (N_40479,N_40212,N_40016);
and U40480 (N_40480,N_40130,N_40144);
nor U40481 (N_40481,N_40033,N_40010);
nor U40482 (N_40482,N_40092,N_40128);
or U40483 (N_40483,N_40007,N_40061);
nand U40484 (N_40484,N_40123,N_40016);
and U40485 (N_40485,N_40100,N_40212);
nor U40486 (N_40486,N_40179,N_40147);
xor U40487 (N_40487,N_40137,N_40195);
or U40488 (N_40488,N_40237,N_40013);
xor U40489 (N_40489,N_40152,N_40043);
xnor U40490 (N_40490,N_40194,N_40106);
or U40491 (N_40491,N_40209,N_40221);
or U40492 (N_40492,N_40150,N_40064);
and U40493 (N_40493,N_40056,N_40236);
nand U40494 (N_40494,N_40223,N_40245);
nand U40495 (N_40495,N_40030,N_40043);
and U40496 (N_40496,N_40177,N_40204);
or U40497 (N_40497,N_40069,N_40021);
or U40498 (N_40498,N_40240,N_40053);
nand U40499 (N_40499,N_40011,N_40038);
nor U40500 (N_40500,N_40387,N_40379);
or U40501 (N_40501,N_40269,N_40428);
and U40502 (N_40502,N_40346,N_40381);
or U40503 (N_40503,N_40455,N_40252);
and U40504 (N_40504,N_40450,N_40304);
nand U40505 (N_40505,N_40293,N_40330);
nor U40506 (N_40506,N_40266,N_40311);
nand U40507 (N_40507,N_40426,N_40321);
and U40508 (N_40508,N_40490,N_40338);
and U40509 (N_40509,N_40340,N_40421);
or U40510 (N_40510,N_40474,N_40345);
nand U40511 (N_40511,N_40283,N_40301);
and U40512 (N_40512,N_40414,N_40363);
xor U40513 (N_40513,N_40393,N_40373);
and U40514 (N_40514,N_40388,N_40313);
and U40515 (N_40515,N_40280,N_40361);
and U40516 (N_40516,N_40440,N_40480);
xor U40517 (N_40517,N_40377,N_40397);
and U40518 (N_40518,N_40425,N_40454);
and U40519 (N_40519,N_40289,N_40385);
nor U40520 (N_40520,N_40386,N_40374);
and U40521 (N_40521,N_40489,N_40306);
nor U40522 (N_40522,N_40255,N_40410);
and U40523 (N_40523,N_40453,N_40367);
xor U40524 (N_40524,N_40261,N_40403);
xor U40525 (N_40525,N_40407,N_40469);
or U40526 (N_40526,N_40436,N_40467);
nand U40527 (N_40527,N_40378,N_40282);
and U40528 (N_40528,N_40401,N_40492);
xnor U40529 (N_40529,N_40483,N_40427);
or U40530 (N_40530,N_40431,N_40267);
nor U40531 (N_40531,N_40417,N_40400);
and U40532 (N_40532,N_40302,N_40292);
xor U40533 (N_40533,N_40456,N_40333);
xnor U40534 (N_40534,N_40419,N_40380);
nand U40535 (N_40535,N_40351,N_40310);
nand U40536 (N_40536,N_40478,N_40487);
or U40537 (N_40537,N_40352,N_40299);
or U40538 (N_40538,N_40257,N_40498);
or U40539 (N_40539,N_40461,N_40260);
nand U40540 (N_40540,N_40324,N_40392);
and U40541 (N_40541,N_40491,N_40424);
and U40542 (N_40542,N_40368,N_40458);
nor U40543 (N_40543,N_40357,N_40296);
xnor U40544 (N_40544,N_40268,N_40308);
nand U40545 (N_40545,N_40452,N_40354);
nor U40546 (N_40546,N_40481,N_40300);
or U40547 (N_40547,N_40418,N_40320);
or U40548 (N_40548,N_40430,N_40499);
or U40549 (N_40549,N_40286,N_40375);
and U40550 (N_40550,N_40413,N_40332);
nor U40551 (N_40551,N_40314,N_40391);
nor U40552 (N_40552,N_40468,N_40295);
and U40553 (N_40553,N_40347,N_40274);
nor U40554 (N_40554,N_40256,N_40482);
nand U40555 (N_40555,N_40325,N_40285);
nor U40556 (N_40556,N_40350,N_40326);
xnor U40557 (N_40557,N_40359,N_40497);
xor U40558 (N_40558,N_40416,N_40264);
or U40559 (N_40559,N_40476,N_40429);
and U40560 (N_40560,N_40402,N_40395);
and U40561 (N_40561,N_40415,N_40254);
nor U40562 (N_40562,N_40370,N_40449);
nor U40563 (N_40563,N_40448,N_40464);
nand U40564 (N_40564,N_40253,N_40439);
xnor U40565 (N_40565,N_40488,N_40250);
or U40566 (N_40566,N_40327,N_40298);
xor U40567 (N_40567,N_40451,N_40466);
or U40568 (N_40568,N_40494,N_40420);
nand U40569 (N_40569,N_40463,N_40348);
nand U40570 (N_40570,N_40265,N_40344);
nand U40571 (N_40571,N_40318,N_40366);
nor U40572 (N_40572,N_40312,N_40287);
and U40573 (N_40573,N_40472,N_40339);
nor U40574 (N_40574,N_40406,N_40272);
xnor U40575 (N_40575,N_40276,N_40331);
or U40576 (N_40576,N_40432,N_40398);
nand U40577 (N_40577,N_40315,N_40273);
or U40578 (N_40578,N_40275,N_40382);
nor U40579 (N_40579,N_40495,N_40435);
or U40580 (N_40580,N_40364,N_40319);
and U40581 (N_40581,N_40307,N_40323);
and U40582 (N_40582,N_40437,N_40496);
or U40583 (N_40583,N_40457,N_40485);
and U40584 (N_40584,N_40342,N_40328);
nor U40585 (N_40585,N_40258,N_40404);
xor U40586 (N_40586,N_40390,N_40316);
nor U40587 (N_40587,N_40389,N_40423);
nand U40588 (N_40588,N_40441,N_40438);
or U40589 (N_40589,N_40278,N_40349);
nand U40590 (N_40590,N_40270,N_40465);
and U40591 (N_40591,N_40294,N_40411);
nor U40592 (N_40592,N_40251,N_40277);
nor U40593 (N_40593,N_40263,N_40412);
nand U40594 (N_40594,N_40262,N_40446);
or U40595 (N_40595,N_40281,N_40309);
nand U40596 (N_40596,N_40405,N_40334);
or U40597 (N_40597,N_40356,N_40443);
xnor U40598 (N_40598,N_40479,N_40445);
and U40599 (N_40599,N_40493,N_40409);
or U40600 (N_40600,N_40473,N_40329);
and U40601 (N_40601,N_40399,N_40297);
and U40602 (N_40602,N_40317,N_40394);
xnor U40603 (N_40603,N_40322,N_40470);
or U40604 (N_40604,N_40365,N_40279);
nand U40605 (N_40605,N_40372,N_40288);
and U40606 (N_40606,N_40336,N_40335);
and U40607 (N_40607,N_40362,N_40305);
or U40608 (N_40608,N_40290,N_40447);
nor U40609 (N_40609,N_40369,N_40442);
or U40610 (N_40610,N_40486,N_40355);
xor U40611 (N_40611,N_40337,N_40343);
nand U40612 (N_40612,N_40422,N_40303);
nand U40613 (N_40613,N_40384,N_40271);
nor U40614 (N_40614,N_40358,N_40408);
nor U40615 (N_40615,N_40396,N_40383);
or U40616 (N_40616,N_40353,N_40475);
xor U40617 (N_40617,N_40471,N_40477);
nor U40618 (N_40618,N_40371,N_40341);
xnor U40619 (N_40619,N_40434,N_40460);
nor U40620 (N_40620,N_40459,N_40484);
and U40621 (N_40621,N_40462,N_40376);
xnor U40622 (N_40622,N_40259,N_40291);
or U40623 (N_40623,N_40444,N_40433);
nor U40624 (N_40624,N_40360,N_40284);
nor U40625 (N_40625,N_40325,N_40415);
or U40626 (N_40626,N_40335,N_40479);
nor U40627 (N_40627,N_40477,N_40271);
and U40628 (N_40628,N_40468,N_40294);
nand U40629 (N_40629,N_40370,N_40290);
nand U40630 (N_40630,N_40442,N_40359);
and U40631 (N_40631,N_40295,N_40406);
xor U40632 (N_40632,N_40304,N_40322);
and U40633 (N_40633,N_40289,N_40316);
or U40634 (N_40634,N_40361,N_40356);
or U40635 (N_40635,N_40290,N_40466);
xnor U40636 (N_40636,N_40429,N_40498);
xnor U40637 (N_40637,N_40340,N_40487);
and U40638 (N_40638,N_40256,N_40307);
or U40639 (N_40639,N_40403,N_40253);
xnor U40640 (N_40640,N_40446,N_40450);
nand U40641 (N_40641,N_40459,N_40260);
nor U40642 (N_40642,N_40477,N_40345);
xor U40643 (N_40643,N_40294,N_40438);
or U40644 (N_40644,N_40345,N_40470);
and U40645 (N_40645,N_40424,N_40328);
and U40646 (N_40646,N_40283,N_40453);
or U40647 (N_40647,N_40264,N_40280);
or U40648 (N_40648,N_40340,N_40465);
nand U40649 (N_40649,N_40310,N_40303);
nand U40650 (N_40650,N_40437,N_40332);
and U40651 (N_40651,N_40300,N_40282);
xor U40652 (N_40652,N_40313,N_40379);
or U40653 (N_40653,N_40347,N_40404);
or U40654 (N_40654,N_40312,N_40440);
xnor U40655 (N_40655,N_40350,N_40275);
nor U40656 (N_40656,N_40396,N_40252);
xor U40657 (N_40657,N_40342,N_40488);
and U40658 (N_40658,N_40482,N_40411);
and U40659 (N_40659,N_40340,N_40276);
or U40660 (N_40660,N_40372,N_40333);
xnor U40661 (N_40661,N_40404,N_40406);
nor U40662 (N_40662,N_40356,N_40497);
or U40663 (N_40663,N_40280,N_40282);
nand U40664 (N_40664,N_40488,N_40309);
or U40665 (N_40665,N_40378,N_40268);
and U40666 (N_40666,N_40448,N_40479);
nand U40667 (N_40667,N_40444,N_40388);
nor U40668 (N_40668,N_40453,N_40446);
or U40669 (N_40669,N_40330,N_40335);
or U40670 (N_40670,N_40489,N_40309);
nand U40671 (N_40671,N_40336,N_40253);
nand U40672 (N_40672,N_40288,N_40385);
and U40673 (N_40673,N_40324,N_40334);
or U40674 (N_40674,N_40269,N_40284);
or U40675 (N_40675,N_40479,N_40288);
xnor U40676 (N_40676,N_40287,N_40333);
xor U40677 (N_40677,N_40418,N_40331);
or U40678 (N_40678,N_40391,N_40352);
nor U40679 (N_40679,N_40299,N_40322);
nand U40680 (N_40680,N_40439,N_40331);
nand U40681 (N_40681,N_40301,N_40323);
or U40682 (N_40682,N_40337,N_40414);
nor U40683 (N_40683,N_40322,N_40265);
and U40684 (N_40684,N_40302,N_40494);
or U40685 (N_40685,N_40336,N_40413);
nand U40686 (N_40686,N_40258,N_40474);
xnor U40687 (N_40687,N_40326,N_40411);
and U40688 (N_40688,N_40252,N_40496);
nor U40689 (N_40689,N_40276,N_40416);
nor U40690 (N_40690,N_40327,N_40289);
and U40691 (N_40691,N_40306,N_40408);
xor U40692 (N_40692,N_40341,N_40462);
and U40693 (N_40693,N_40439,N_40414);
or U40694 (N_40694,N_40301,N_40314);
nor U40695 (N_40695,N_40397,N_40371);
or U40696 (N_40696,N_40343,N_40383);
nand U40697 (N_40697,N_40364,N_40266);
xnor U40698 (N_40698,N_40266,N_40360);
nor U40699 (N_40699,N_40454,N_40391);
and U40700 (N_40700,N_40437,N_40319);
nor U40701 (N_40701,N_40264,N_40455);
nand U40702 (N_40702,N_40413,N_40277);
and U40703 (N_40703,N_40292,N_40484);
or U40704 (N_40704,N_40446,N_40251);
xor U40705 (N_40705,N_40303,N_40425);
nor U40706 (N_40706,N_40354,N_40343);
and U40707 (N_40707,N_40260,N_40361);
nand U40708 (N_40708,N_40275,N_40283);
nand U40709 (N_40709,N_40339,N_40445);
nand U40710 (N_40710,N_40429,N_40495);
xor U40711 (N_40711,N_40347,N_40301);
and U40712 (N_40712,N_40261,N_40389);
or U40713 (N_40713,N_40395,N_40494);
or U40714 (N_40714,N_40469,N_40446);
nand U40715 (N_40715,N_40462,N_40429);
xor U40716 (N_40716,N_40321,N_40404);
nand U40717 (N_40717,N_40296,N_40402);
or U40718 (N_40718,N_40367,N_40430);
xor U40719 (N_40719,N_40446,N_40421);
nor U40720 (N_40720,N_40251,N_40326);
nor U40721 (N_40721,N_40258,N_40478);
xnor U40722 (N_40722,N_40441,N_40253);
and U40723 (N_40723,N_40328,N_40391);
and U40724 (N_40724,N_40307,N_40406);
nor U40725 (N_40725,N_40339,N_40275);
nand U40726 (N_40726,N_40266,N_40298);
nand U40727 (N_40727,N_40288,N_40376);
and U40728 (N_40728,N_40325,N_40369);
xor U40729 (N_40729,N_40470,N_40440);
or U40730 (N_40730,N_40372,N_40427);
nor U40731 (N_40731,N_40470,N_40463);
xnor U40732 (N_40732,N_40424,N_40259);
nand U40733 (N_40733,N_40487,N_40291);
and U40734 (N_40734,N_40348,N_40432);
xor U40735 (N_40735,N_40326,N_40315);
and U40736 (N_40736,N_40466,N_40468);
and U40737 (N_40737,N_40363,N_40419);
xnor U40738 (N_40738,N_40492,N_40386);
xnor U40739 (N_40739,N_40413,N_40464);
and U40740 (N_40740,N_40321,N_40467);
or U40741 (N_40741,N_40306,N_40328);
nor U40742 (N_40742,N_40320,N_40494);
xnor U40743 (N_40743,N_40455,N_40303);
nand U40744 (N_40744,N_40440,N_40296);
xor U40745 (N_40745,N_40381,N_40258);
nand U40746 (N_40746,N_40480,N_40467);
nand U40747 (N_40747,N_40415,N_40450);
nor U40748 (N_40748,N_40487,N_40275);
and U40749 (N_40749,N_40377,N_40408);
nor U40750 (N_40750,N_40569,N_40536);
and U40751 (N_40751,N_40543,N_40529);
xor U40752 (N_40752,N_40650,N_40613);
or U40753 (N_40753,N_40680,N_40584);
or U40754 (N_40754,N_40702,N_40512);
and U40755 (N_40755,N_40735,N_40530);
or U40756 (N_40756,N_40544,N_40582);
or U40757 (N_40757,N_40557,N_40502);
or U40758 (N_40758,N_40696,N_40534);
nor U40759 (N_40759,N_40678,N_40733);
xnor U40760 (N_40760,N_40576,N_40659);
nor U40761 (N_40761,N_40522,N_40681);
nand U40762 (N_40762,N_40667,N_40662);
xnor U40763 (N_40763,N_40690,N_40615);
and U40764 (N_40764,N_40649,N_40636);
nand U40765 (N_40765,N_40596,N_40742);
and U40766 (N_40766,N_40575,N_40525);
nor U40767 (N_40767,N_40614,N_40588);
and U40768 (N_40768,N_40521,N_40602);
or U40769 (N_40769,N_40558,N_40703);
nor U40770 (N_40770,N_40620,N_40617);
xnor U40771 (N_40771,N_40689,N_40728);
and U40772 (N_40772,N_40545,N_40622);
and U40773 (N_40773,N_40727,N_40568);
and U40774 (N_40774,N_40510,N_40657);
nor U40775 (N_40775,N_40717,N_40719);
xor U40776 (N_40776,N_40720,N_40671);
xnor U40777 (N_40777,N_40586,N_40705);
xnor U40778 (N_40778,N_40523,N_40538);
and U40779 (N_40779,N_40707,N_40646);
nor U40780 (N_40780,N_40553,N_40716);
xor U40781 (N_40781,N_40692,N_40741);
or U40782 (N_40782,N_40583,N_40730);
xor U40783 (N_40783,N_40591,N_40592);
and U40784 (N_40784,N_40744,N_40748);
nor U40785 (N_40785,N_40539,N_40688);
nand U40786 (N_40786,N_40599,N_40611);
nor U40787 (N_40787,N_40648,N_40693);
nor U40788 (N_40788,N_40504,N_40736);
or U40789 (N_40789,N_40710,N_40652);
and U40790 (N_40790,N_40527,N_40714);
or U40791 (N_40791,N_40686,N_40628);
xnor U40792 (N_40792,N_40559,N_40640);
xnor U40793 (N_40793,N_40675,N_40605);
nand U40794 (N_40794,N_40713,N_40516);
nand U40795 (N_40795,N_40551,N_40724);
nand U40796 (N_40796,N_40734,N_40745);
nand U40797 (N_40797,N_40597,N_40743);
nand U40798 (N_40798,N_40631,N_40556);
nand U40799 (N_40799,N_40600,N_40718);
or U40800 (N_40800,N_40555,N_40587);
or U40801 (N_40801,N_40548,N_40700);
or U40802 (N_40802,N_40633,N_40601);
or U40803 (N_40803,N_40749,N_40715);
and U40804 (N_40804,N_40632,N_40624);
or U40805 (N_40805,N_40609,N_40722);
nor U40806 (N_40806,N_40658,N_40571);
xnor U40807 (N_40807,N_40520,N_40738);
nand U40808 (N_40808,N_40511,N_40500);
and U40809 (N_40809,N_40732,N_40721);
and U40810 (N_40810,N_40708,N_40656);
and U40811 (N_40811,N_40687,N_40607);
and U40812 (N_40812,N_40506,N_40517);
nor U40813 (N_40813,N_40641,N_40507);
nand U40814 (N_40814,N_40532,N_40739);
and U40815 (N_40815,N_40673,N_40616);
nor U40816 (N_40816,N_40729,N_40573);
and U40817 (N_40817,N_40590,N_40661);
nor U40818 (N_40818,N_40561,N_40644);
xnor U40819 (N_40819,N_40679,N_40654);
nand U40820 (N_40820,N_40503,N_40666);
or U40821 (N_40821,N_40547,N_40626);
or U40822 (N_40822,N_40706,N_40595);
xor U40823 (N_40823,N_40638,N_40723);
or U40824 (N_40824,N_40508,N_40540);
or U40825 (N_40825,N_40552,N_40712);
xnor U40826 (N_40826,N_40621,N_40672);
xnor U40827 (N_40827,N_40549,N_40637);
nand U40828 (N_40828,N_40580,N_40563);
and U40829 (N_40829,N_40655,N_40560);
and U40830 (N_40830,N_40585,N_40515);
and U40831 (N_40831,N_40701,N_40537);
and U40832 (N_40832,N_40726,N_40604);
nor U40833 (N_40833,N_40684,N_40629);
xnor U40834 (N_40834,N_40565,N_40518);
xnor U40835 (N_40835,N_40594,N_40564);
nand U40836 (N_40836,N_40685,N_40663);
nor U40837 (N_40837,N_40660,N_40669);
xnor U40838 (N_40838,N_40699,N_40501);
nand U40839 (N_40839,N_40581,N_40574);
or U40840 (N_40840,N_40567,N_40589);
and U40841 (N_40841,N_40608,N_40627);
or U40842 (N_40842,N_40695,N_40630);
nand U40843 (N_40843,N_40505,N_40531);
and U40844 (N_40844,N_40610,N_40546);
xnor U40845 (N_40845,N_40664,N_40645);
and U40846 (N_40846,N_40623,N_40677);
nand U40847 (N_40847,N_40528,N_40550);
nand U40848 (N_40848,N_40647,N_40704);
nand U40849 (N_40849,N_40603,N_40541);
nor U40850 (N_40850,N_40642,N_40566);
xor U40851 (N_40851,N_40577,N_40740);
nand U40852 (N_40852,N_40513,N_40542);
nand U40853 (N_40853,N_40634,N_40737);
xor U40854 (N_40854,N_40570,N_40682);
xnor U40855 (N_40855,N_40635,N_40731);
xnor U40856 (N_40856,N_40554,N_40578);
or U40857 (N_40857,N_40683,N_40618);
nor U40858 (N_40858,N_40691,N_40711);
xor U40859 (N_40859,N_40697,N_40606);
or U40860 (N_40860,N_40670,N_40562);
nor U40861 (N_40861,N_40535,N_40579);
nand U40862 (N_40862,N_40524,N_40725);
or U40863 (N_40863,N_40639,N_40619);
nor U40864 (N_40864,N_40509,N_40643);
or U40865 (N_40865,N_40526,N_40746);
xor U40866 (N_40866,N_40676,N_40598);
nand U40867 (N_40867,N_40625,N_40694);
and U40868 (N_40868,N_40612,N_40709);
nand U40869 (N_40869,N_40593,N_40519);
or U40870 (N_40870,N_40665,N_40668);
nand U40871 (N_40871,N_40747,N_40572);
and U40872 (N_40872,N_40674,N_40514);
xnor U40873 (N_40873,N_40651,N_40698);
nand U40874 (N_40874,N_40533,N_40653);
or U40875 (N_40875,N_40612,N_40679);
and U40876 (N_40876,N_40621,N_40575);
nor U40877 (N_40877,N_40517,N_40682);
nand U40878 (N_40878,N_40571,N_40547);
and U40879 (N_40879,N_40649,N_40511);
xnor U40880 (N_40880,N_40629,N_40513);
nand U40881 (N_40881,N_40716,N_40537);
xnor U40882 (N_40882,N_40548,N_40707);
and U40883 (N_40883,N_40683,N_40595);
nor U40884 (N_40884,N_40546,N_40557);
nor U40885 (N_40885,N_40690,N_40692);
xnor U40886 (N_40886,N_40585,N_40553);
nor U40887 (N_40887,N_40642,N_40720);
nand U40888 (N_40888,N_40552,N_40697);
or U40889 (N_40889,N_40631,N_40587);
and U40890 (N_40890,N_40655,N_40727);
or U40891 (N_40891,N_40681,N_40662);
nand U40892 (N_40892,N_40532,N_40630);
and U40893 (N_40893,N_40594,N_40610);
or U40894 (N_40894,N_40556,N_40542);
nor U40895 (N_40895,N_40618,N_40741);
nand U40896 (N_40896,N_40623,N_40699);
and U40897 (N_40897,N_40694,N_40733);
or U40898 (N_40898,N_40667,N_40604);
xnor U40899 (N_40899,N_40544,N_40629);
xor U40900 (N_40900,N_40694,N_40672);
or U40901 (N_40901,N_40545,N_40595);
nor U40902 (N_40902,N_40678,N_40706);
and U40903 (N_40903,N_40599,N_40560);
nor U40904 (N_40904,N_40718,N_40698);
xor U40905 (N_40905,N_40535,N_40547);
nor U40906 (N_40906,N_40706,N_40563);
nor U40907 (N_40907,N_40669,N_40521);
nand U40908 (N_40908,N_40548,N_40603);
xor U40909 (N_40909,N_40692,N_40589);
nor U40910 (N_40910,N_40643,N_40603);
nand U40911 (N_40911,N_40726,N_40605);
or U40912 (N_40912,N_40589,N_40701);
xor U40913 (N_40913,N_40688,N_40623);
xnor U40914 (N_40914,N_40619,N_40707);
nand U40915 (N_40915,N_40539,N_40698);
xor U40916 (N_40916,N_40704,N_40627);
and U40917 (N_40917,N_40514,N_40669);
xnor U40918 (N_40918,N_40705,N_40542);
and U40919 (N_40919,N_40651,N_40641);
nor U40920 (N_40920,N_40645,N_40513);
nor U40921 (N_40921,N_40543,N_40643);
and U40922 (N_40922,N_40558,N_40652);
nand U40923 (N_40923,N_40541,N_40506);
and U40924 (N_40924,N_40597,N_40744);
nor U40925 (N_40925,N_40576,N_40740);
and U40926 (N_40926,N_40618,N_40659);
and U40927 (N_40927,N_40604,N_40744);
or U40928 (N_40928,N_40747,N_40599);
and U40929 (N_40929,N_40531,N_40516);
and U40930 (N_40930,N_40629,N_40511);
nand U40931 (N_40931,N_40520,N_40661);
or U40932 (N_40932,N_40572,N_40557);
nand U40933 (N_40933,N_40616,N_40602);
or U40934 (N_40934,N_40692,N_40633);
nor U40935 (N_40935,N_40556,N_40627);
or U40936 (N_40936,N_40533,N_40744);
and U40937 (N_40937,N_40548,N_40510);
or U40938 (N_40938,N_40660,N_40588);
and U40939 (N_40939,N_40734,N_40518);
or U40940 (N_40940,N_40505,N_40669);
nand U40941 (N_40941,N_40541,N_40621);
nor U40942 (N_40942,N_40542,N_40601);
and U40943 (N_40943,N_40681,N_40698);
nor U40944 (N_40944,N_40742,N_40601);
nand U40945 (N_40945,N_40685,N_40588);
or U40946 (N_40946,N_40691,N_40527);
nor U40947 (N_40947,N_40658,N_40560);
nor U40948 (N_40948,N_40533,N_40630);
nand U40949 (N_40949,N_40621,N_40624);
or U40950 (N_40950,N_40512,N_40635);
and U40951 (N_40951,N_40611,N_40553);
nor U40952 (N_40952,N_40611,N_40632);
nand U40953 (N_40953,N_40723,N_40687);
and U40954 (N_40954,N_40685,N_40534);
or U40955 (N_40955,N_40692,N_40645);
nor U40956 (N_40956,N_40512,N_40746);
or U40957 (N_40957,N_40615,N_40677);
and U40958 (N_40958,N_40749,N_40633);
xnor U40959 (N_40959,N_40725,N_40565);
or U40960 (N_40960,N_40607,N_40649);
xnor U40961 (N_40961,N_40668,N_40509);
nand U40962 (N_40962,N_40717,N_40671);
nand U40963 (N_40963,N_40713,N_40627);
or U40964 (N_40964,N_40605,N_40659);
and U40965 (N_40965,N_40575,N_40545);
nor U40966 (N_40966,N_40585,N_40659);
and U40967 (N_40967,N_40743,N_40553);
and U40968 (N_40968,N_40527,N_40747);
xnor U40969 (N_40969,N_40706,N_40593);
nor U40970 (N_40970,N_40707,N_40669);
xor U40971 (N_40971,N_40607,N_40686);
nor U40972 (N_40972,N_40596,N_40697);
xor U40973 (N_40973,N_40604,N_40634);
nor U40974 (N_40974,N_40661,N_40725);
nor U40975 (N_40975,N_40649,N_40621);
nand U40976 (N_40976,N_40691,N_40607);
nand U40977 (N_40977,N_40640,N_40586);
xnor U40978 (N_40978,N_40596,N_40730);
xnor U40979 (N_40979,N_40720,N_40669);
xnor U40980 (N_40980,N_40570,N_40593);
xnor U40981 (N_40981,N_40594,N_40506);
nor U40982 (N_40982,N_40556,N_40643);
xnor U40983 (N_40983,N_40661,N_40612);
xnor U40984 (N_40984,N_40615,N_40678);
xnor U40985 (N_40985,N_40586,N_40663);
nand U40986 (N_40986,N_40707,N_40687);
xor U40987 (N_40987,N_40593,N_40564);
and U40988 (N_40988,N_40690,N_40664);
nand U40989 (N_40989,N_40597,N_40572);
xnor U40990 (N_40990,N_40630,N_40726);
nand U40991 (N_40991,N_40727,N_40633);
and U40992 (N_40992,N_40663,N_40544);
xnor U40993 (N_40993,N_40640,N_40615);
nand U40994 (N_40994,N_40621,N_40632);
or U40995 (N_40995,N_40663,N_40666);
nor U40996 (N_40996,N_40740,N_40720);
nor U40997 (N_40997,N_40586,N_40555);
nor U40998 (N_40998,N_40538,N_40637);
nand U40999 (N_40999,N_40704,N_40653);
xnor U41000 (N_41000,N_40772,N_40938);
and U41001 (N_41001,N_40916,N_40835);
nand U41002 (N_41002,N_40862,N_40834);
or U41003 (N_41003,N_40962,N_40908);
nor U41004 (N_41004,N_40879,N_40960);
and U41005 (N_41005,N_40993,N_40930);
xor U41006 (N_41006,N_40891,N_40795);
and U41007 (N_41007,N_40926,N_40771);
and U41008 (N_41008,N_40814,N_40924);
nor U41009 (N_41009,N_40756,N_40825);
or U41010 (N_41010,N_40997,N_40757);
or U41011 (N_41011,N_40932,N_40815);
or U41012 (N_41012,N_40858,N_40765);
nand U41013 (N_41013,N_40880,N_40863);
and U41014 (N_41014,N_40803,N_40837);
and U41015 (N_41015,N_40783,N_40827);
nand U41016 (N_41016,N_40994,N_40802);
xnor U41017 (N_41017,N_40974,N_40760);
and U41018 (N_41018,N_40910,N_40807);
and U41019 (N_41019,N_40884,N_40774);
or U41020 (N_41020,N_40770,N_40831);
nand U41021 (N_41021,N_40841,N_40819);
or U41022 (N_41022,N_40791,N_40763);
xor U41023 (N_41023,N_40887,N_40792);
or U41024 (N_41024,N_40768,N_40923);
nor U41025 (N_41025,N_40842,N_40868);
or U41026 (N_41026,N_40758,N_40816);
nor U41027 (N_41027,N_40843,N_40913);
xor U41028 (N_41028,N_40999,N_40904);
or U41029 (N_41029,N_40817,N_40839);
or U41030 (N_41030,N_40810,N_40821);
nand U41031 (N_41031,N_40988,N_40861);
or U41032 (N_41032,N_40968,N_40992);
xor U41033 (N_41033,N_40766,N_40948);
nor U41034 (N_41034,N_40995,N_40976);
or U41035 (N_41035,N_40941,N_40900);
and U41036 (N_41036,N_40801,N_40942);
nand U41037 (N_41037,N_40920,N_40922);
and U41038 (N_41038,N_40973,N_40873);
and U41039 (N_41039,N_40865,N_40851);
and U41040 (N_41040,N_40852,N_40806);
nor U41041 (N_41041,N_40944,N_40977);
and U41042 (N_41042,N_40940,N_40951);
nor U41043 (N_41043,N_40979,N_40934);
nor U41044 (N_41044,N_40897,N_40848);
nand U41045 (N_41045,N_40780,N_40845);
xor U41046 (N_41046,N_40933,N_40808);
or U41047 (N_41047,N_40833,N_40964);
and U41048 (N_41048,N_40917,N_40939);
and U41049 (N_41049,N_40869,N_40946);
or U41050 (N_41050,N_40824,N_40987);
nand U41051 (N_41051,N_40877,N_40965);
nand U41052 (N_41052,N_40996,N_40889);
and U41053 (N_41053,N_40892,N_40871);
and U41054 (N_41054,N_40844,N_40778);
and U41055 (N_41055,N_40828,N_40779);
xnor U41056 (N_41056,N_40928,N_40882);
nor U41057 (N_41057,N_40867,N_40752);
or U41058 (N_41058,N_40947,N_40911);
and U41059 (N_41059,N_40853,N_40901);
or U41060 (N_41060,N_40769,N_40898);
xnor U41061 (N_41061,N_40755,N_40903);
nand U41062 (N_41062,N_40982,N_40893);
or U41063 (N_41063,N_40966,N_40796);
or U41064 (N_41064,N_40914,N_40784);
or U41065 (N_41065,N_40986,N_40823);
nor U41066 (N_41066,N_40909,N_40886);
xor U41067 (N_41067,N_40989,N_40870);
nand U41068 (N_41068,N_40800,N_40754);
nor U41069 (N_41069,N_40972,N_40876);
nor U41070 (N_41070,N_40902,N_40840);
and U41071 (N_41071,N_40927,N_40912);
or U41072 (N_41072,N_40753,N_40856);
xor U41073 (N_41073,N_40885,N_40907);
and U41074 (N_41074,N_40931,N_40943);
nor U41075 (N_41075,N_40751,N_40915);
and U41076 (N_41076,N_40957,N_40854);
nand U41077 (N_41077,N_40857,N_40820);
nand U41078 (N_41078,N_40764,N_40929);
or U41079 (N_41079,N_40991,N_40855);
nor U41080 (N_41080,N_40955,N_40785);
and U41081 (N_41081,N_40925,N_40949);
nor U41082 (N_41082,N_40826,N_40937);
or U41083 (N_41083,N_40990,N_40789);
xor U41084 (N_41084,N_40775,N_40804);
nor U41085 (N_41085,N_40818,N_40980);
and U41086 (N_41086,N_40954,N_40809);
xor U41087 (N_41087,N_40847,N_40793);
nor U41088 (N_41088,N_40759,N_40894);
nor U41089 (N_41089,N_40899,N_40978);
nor U41090 (N_41090,N_40984,N_40935);
nand U41091 (N_41091,N_40822,N_40881);
or U41092 (N_41092,N_40945,N_40794);
xor U41093 (N_41093,N_40975,N_40866);
nor U41094 (N_41094,N_40788,N_40829);
and U41095 (N_41095,N_40776,N_40782);
nand U41096 (N_41096,N_40878,N_40919);
xor U41097 (N_41097,N_40985,N_40872);
and U41098 (N_41098,N_40781,N_40798);
xor U41099 (N_41099,N_40959,N_40761);
or U41100 (N_41100,N_40875,N_40936);
nand U41101 (N_41101,N_40864,N_40811);
and U41102 (N_41102,N_40918,N_40921);
and U41103 (N_41103,N_40983,N_40998);
nand U41104 (N_41104,N_40846,N_40956);
or U41105 (N_41105,N_40888,N_40836);
or U41106 (N_41106,N_40967,N_40952);
and U41107 (N_41107,N_40859,N_40860);
nor U41108 (N_41108,N_40797,N_40787);
and U41109 (N_41109,N_40958,N_40961);
and U41110 (N_41110,N_40838,N_40971);
nor U41111 (N_41111,N_40906,N_40762);
xnor U41112 (N_41112,N_40963,N_40812);
xnor U41113 (N_41113,N_40750,N_40786);
nor U41114 (N_41114,N_40777,N_40981);
nand U41115 (N_41115,N_40832,N_40830);
or U41116 (N_41116,N_40805,N_40883);
nor U41117 (N_41117,N_40896,N_40895);
nand U41118 (N_41118,N_40799,N_40969);
and U41119 (N_41119,N_40905,N_40890);
nor U41120 (N_41120,N_40874,N_40773);
and U41121 (N_41121,N_40813,N_40850);
xor U41122 (N_41122,N_40849,N_40767);
nand U41123 (N_41123,N_40790,N_40950);
xnor U41124 (N_41124,N_40970,N_40953);
nor U41125 (N_41125,N_40868,N_40928);
nor U41126 (N_41126,N_40871,N_40966);
or U41127 (N_41127,N_40990,N_40950);
xor U41128 (N_41128,N_40931,N_40876);
nor U41129 (N_41129,N_40961,N_40927);
or U41130 (N_41130,N_40794,N_40927);
xor U41131 (N_41131,N_40993,N_40903);
nor U41132 (N_41132,N_40859,N_40831);
xor U41133 (N_41133,N_40936,N_40758);
nor U41134 (N_41134,N_40884,N_40806);
nand U41135 (N_41135,N_40927,N_40944);
nor U41136 (N_41136,N_40872,N_40776);
or U41137 (N_41137,N_40897,N_40983);
and U41138 (N_41138,N_40928,N_40909);
xnor U41139 (N_41139,N_40912,N_40925);
nand U41140 (N_41140,N_40834,N_40800);
or U41141 (N_41141,N_40911,N_40962);
or U41142 (N_41142,N_40868,N_40845);
nor U41143 (N_41143,N_40753,N_40989);
nor U41144 (N_41144,N_40953,N_40851);
and U41145 (N_41145,N_40870,N_40756);
nand U41146 (N_41146,N_40961,N_40944);
xor U41147 (N_41147,N_40841,N_40778);
and U41148 (N_41148,N_40929,N_40935);
nand U41149 (N_41149,N_40958,N_40949);
and U41150 (N_41150,N_40877,N_40937);
or U41151 (N_41151,N_40807,N_40896);
or U41152 (N_41152,N_40791,N_40750);
or U41153 (N_41153,N_40996,N_40812);
or U41154 (N_41154,N_40840,N_40916);
nor U41155 (N_41155,N_40916,N_40952);
nor U41156 (N_41156,N_40983,N_40775);
and U41157 (N_41157,N_40799,N_40857);
nor U41158 (N_41158,N_40946,N_40773);
xnor U41159 (N_41159,N_40905,N_40949);
nand U41160 (N_41160,N_40997,N_40970);
and U41161 (N_41161,N_40877,N_40978);
nor U41162 (N_41162,N_40821,N_40901);
xnor U41163 (N_41163,N_40836,N_40881);
and U41164 (N_41164,N_40987,N_40852);
xor U41165 (N_41165,N_40889,N_40988);
and U41166 (N_41166,N_40937,N_40991);
nand U41167 (N_41167,N_40890,N_40946);
nand U41168 (N_41168,N_40966,N_40851);
or U41169 (N_41169,N_40899,N_40927);
xor U41170 (N_41170,N_40818,N_40955);
and U41171 (N_41171,N_40833,N_40916);
nand U41172 (N_41172,N_40864,N_40880);
or U41173 (N_41173,N_40793,N_40826);
nand U41174 (N_41174,N_40919,N_40858);
nand U41175 (N_41175,N_40769,N_40781);
nor U41176 (N_41176,N_40845,N_40917);
and U41177 (N_41177,N_40972,N_40771);
nor U41178 (N_41178,N_40811,N_40786);
nand U41179 (N_41179,N_40830,N_40881);
and U41180 (N_41180,N_40916,N_40869);
nor U41181 (N_41181,N_40934,N_40904);
nand U41182 (N_41182,N_40771,N_40937);
nand U41183 (N_41183,N_40913,N_40854);
or U41184 (N_41184,N_40854,N_40855);
nand U41185 (N_41185,N_40781,N_40818);
xor U41186 (N_41186,N_40887,N_40852);
nor U41187 (N_41187,N_40784,N_40794);
or U41188 (N_41188,N_40985,N_40958);
nor U41189 (N_41189,N_40794,N_40850);
or U41190 (N_41190,N_40922,N_40915);
or U41191 (N_41191,N_40846,N_40832);
or U41192 (N_41192,N_40988,N_40841);
nand U41193 (N_41193,N_40807,N_40956);
nand U41194 (N_41194,N_40877,N_40800);
nor U41195 (N_41195,N_40934,N_40750);
and U41196 (N_41196,N_40906,N_40831);
and U41197 (N_41197,N_40988,N_40919);
or U41198 (N_41198,N_40887,N_40831);
or U41199 (N_41199,N_40845,N_40970);
and U41200 (N_41200,N_40944,N_40976);
nor U41201 (N_41201,N_40988,N_40778);
nor U41202 (N_41202,N_40910,N_40771);
or U41203 (N_41203,N_40928,N_40770);
or U41204 (N_41204,N_40968,N_40927);
nand U41205 (N_41205,N_40837,N_40870);
xor U41206 (N_41206,N_40945,N_40913);
xor U41207 (N_41207,N_40995,N_40764);
xor U41208 (N_41208,N_40993,N_40875);
and U41209 (N_41209,N_40859,N_40804);
nand U41210 (N_41210,N_40765,N_40811);
and U41211 (N_41211,N_40937,N_40982);
or U41212 (N_41212,N_40853,N_40754);
nand U41213 (N_41213,N_40918,N_40850);
and U41214 (N_41214,N_40823,N_40871);
and U41215 (N_41215,N_40772,N_40924);
or U41216 (N_41216,N_40761,N_40844);
xnor U41217 (N_41217,N_40785,N_40840);
and U41218 (N_41218,N_40792,N_40882);
or U41219 (N_41219,N_40940,N_40784);
nand U41220 (N_41220,N_40984,N_40903);
and U41221 (N_41221,N_40894,N_40783);
nor U41222 (N_41222,N_40930,N_40989);
xor U41223 (N_41223,N_40985,N_40772);
xor U41224 (N_41224,N_40775,N_40791);
xor U41225 (N_41225,N_40778,N_40905);
and U41226 (N_41226,N_40854,N_40775);
and U41227 (N_41227,N_40774,N_40795);
xnor U41228 (N_41228,N_40806,N_40880);
xnor U41229 (N_41229,N_40939,N_40844);
and U41230 (N_41230,N_40808,N_40974);
nand U41231 (N_41231,N_40866,N_40762);
or U41232 (N_41232,N_40808,N_40998);
nor U41233 (N_41233,N_40849,N_40817);
or U41234 (N_41234,N_40756,N_40986);
or U41235 (N_41235,N_40904,N_40979);
or U41236 (N_41236,N_40862,N_40795);
xnor U41237 (N_41237,N_40988,N_40905);
nor U41238 (N_41238,N_40896,N_40760);
xor U41239 (N_41239,N_40918,N_40764);
or U41240 (N_41240,N_40863,N_40889);
and U41241 (N_41241,N_40780,N_40926);
and U41242 (N_41242,N_40770,N_40833);
or U41243 (N_41243,N_40805,N_40770);
and U41244 (N_41244,N_40783,N_40921);
and U41245 (N_41245,N_40985,N_40924);
xnor U41246 (N_41246,N_40977,N_40911);
xnor U41247 (N_41247,N_40752,N_40899);
xor U41248 (N_41248,N_40755,N_40859);
nand U41249 (N_41249,N_40905,N_40967);
or U41250 (N_41250,N_41077,N_41197);
nor U41251 (N_41251,N_41118,N_41199);
nor U41252 (N_41252,N_41101,N_41117);
and U41253 (N_41253,N_41207,N_41193);
nand U41254 (N_41254,N_41029,N_41106);
nor U41255 (N_41255,N_41176,N_41010);
and U41256 (N_41256,N_41088,N_41071);
nor U41257 (N_41257,N_41219,N_41189);
or U41258 (N_41258,N_41167,N_41142);
xnor U41259 (N_41259,N_41196,N_41217);
and U41260 (N_41260,N_41124,N_41178);
nand U41261 (N_41261,N_41125,N_41127);
nand U41262 (N_41262,N_41240,N_41113);
or U41263 (N_41263,N_41063,N_41062);
and U41264 (N_41264,N_41170,N_41021);
xor U41265 (N_41265,N_41109,N_41094);
and U41266 (N_41266,N_41216,N_41049);
or U41267 (N_41267,N_41036,N_41209);
nand U41268 (N_41268,N_41005,N_41091);
and U41269 (N_41269,N_41007,N_41107);
nor U41270 (N_41270,N_41237,N_41031);
nand U41271 (N_41271,N_41056,N_41030);
nor U41272 (N_41272,N_41085,N_41114);
nand U41273 (N_41273,N_41139,N_41152);
and U41274 (N_41274,N_41111,N_41080);
or U41275 (N_41275,N_41009,N_41149);
or U41276 (N_41276,N_41055,N_41132);
xor U41277 (N_41277,N_41203,N_41163);
nor U41278 (N_41278,N_41000,N_41110);
and U41279 (N_41279,N_41181,N_41060);
nor U41280 (N_41280,N_41228,N_41034);
or U41281 (N_41281,N_41025,N_41160);
and U41282 (N_41282,N_41001,N_41061);
nand U41283 (N_41283,N_41024,N_41246);
and U41284 (N_41284,N_41221,N_41171);
or U41285 (N_41285,N_41225,N_41116);
or U41286 (N_41286,N_41090,N_41128);
xnor U41287 (N_41287,N_41235,N_41115);
xor U41288 (N_41288,N_41184,N_41173);
or U41289 (N_41289,N_41103,N_41039);
xnor U41290 (N_41290,N_41230,N_41206);
xnor U41291 (N_41291,N_41015,N_41019);
and U41292 (N_41292,N_41134,N_41003);
xnor U41293 (N_41293,N_41122,N_41131);
or U41294 (N_41294,N_41180,N_41070);
or U41295 (N_41295,N_41017,N_41161);
xor U41296 (N_41296,N_41157,N_41130);
nor U41297 (N_41297,N_41084,N_41037);
or U41298 (N_41298,N_41166,N_41148);
nor U41299 (N_41299,N_41226,N_41045);
xnor U41300 (N_41300,N_41231,N_41182);
nor U41301 (N_41301,N_41175,N_41075);
nor U41302 (N_41302,N_41040,N_41201);
nor U41303 (N_41303,N_41057,N_41119);
nand U41304 (N_41304,N_41082,N_41096);
xnor U41305 (N_41305,N_41092,N_41027);
and U41306 (N_41306,N_41081,N_41086);
xnor U41307 (N_41307,N_41046,N_41064);
nor U41308 (N_41308,N_41105,N_41174);
and U41309 (N_41309,N_41162,N_41242);
and U41310 (N_41310,N_41195,N_41141);
nor U41311 (N_41311,N_41241,N_41190);
nor U41312 (N_41312,N_41013,N_41018);
or U41313 (N_41313,N_41028,N_41200);
nor U41314 (N_41314,N_41047,N_41043);
nand U41315 (N_41315,N_41194,N_41095);
xnor U41316 (N_41316,N_41068,N_41067);
nor U41317 (N_41317,N_41041,N_41243);
nor U41318 (N_41318,N_41072,N_41227);
nor U41319 (N_41319,N_41249,N_41098);
nand U41320 (N_41320,N_41198,N_41008);
and U41321 (N_41321,N_41129,N_41137);
and U41322 (N_41322,N_41154,N_41168);
nand U41323 (N_41323,N_41052,N_41074);
and U41324 (N_41324,N_41229,N_41026);
nor U41325 (N_41325,N_41053,N_41069);
and U41326 (N_41326,N_41022,N_41020);
nor U41327 (N_41327,N_41215,N_41108);
nor U41328 (N_41328,N_41218,N_41099);
nor U41329 (N_41329,N_41223,N_41136);
and U41330 (N_41330,N_41205,N_41126);
nand U41331 (N_41331,N_41054,N_41151);
nand U41332 (N_41332,N_41002,N_41222);
and U41333 (N_41333,N_41066,N_41204);
or U41334 (N_41334,N_41011,N_41073);
nand U41335 (N_41335,N_41112,N_41211);
xnor U41336 (N_41336,N_41210,N_41093);
and U41337 (N_41337,N_41038,N_41236);
xor U41338 (N_41338,N_41183,N_41089);
and U41339 (N_41339,N_41032,N_41083);
nand U41340 (N_41340,N_41239,N_41233);
xor U41341 (N_41341,N_41133,N_41153);
or U41342 (N_41342,N_41244,N_41042);
and U41343 (N_41343,N_41076,N_41104);
xnor U41344 (N_41344,N_41248,N_41065);
nor U41345 (N_41345,N_41012,N_41192);
nand U41346 (N_41346,N_41247,N_41006);
nand U41347 (N_41347,N_41033,N_41138);
xnor U41348 (N_41348,N_41156,N_41238);
xor U41349 (N_41349,N_41213,N_41147);
xnor U41350 (N_41350,N_41102,N_41035);
nor U41351 (N_41351,N_41078,N_41058);
nand U41352 (N_41352,N_41186,N_41191);
nand U41353 (N_41353,N_41120,N_41059);
and U41354 (N_41354,N_41208,N_41050);
xor U41355 (N_41355,N_41004,N_41179);
or U41356 (N_41356,N_41016,N_41158);
or U41357 (N_41357,N_41145,N_41135);
or U41358 (N_41358,N_41220,N_41097);
nand U41359 (N_41359,N_41143,N_41185);
xnor U41360 (N_41360,N_41165,N_41224);
and U41361 (N_41361,N_41023,N_41150);
nor U41362 (N_41362,N_41048,N_41155);
nand U41363 (N_41363,N_41140,N_41014);
nor U41364 (N_41364,N_41144,N_41159);
nand U41365 (N_41365,N_41172,N_41212);
nor U41366 (N_41366,N_41177,N_41214);
and U41367 (N_41367,N_41087,N_41164);
and U41368 (N_41368,N_41079,N_41123);
and U41369 (N_41369,N_41051,N_41044);
or U41370 (N_41370,N_41146,N_41234);
nand U41371 (N_41371,N_41187,N_41245);
nand U41372 (N_41372,N_41100,N_41188);
or U41373 (N_41373,N_41169,N_41121);
xor U41374 (N_41374,N_41232,N_41202);
nand U41375 (N_41375,N_41242,N_41173);
nor U41376 (N_41376,N_41209,N_41130);
xor U41377 (N_41377,N_41180,N_41111);
nand U41378 (N_41378,N_41044,N_41027);
nand U41379 (N_41379,N_41248,N_41237);
nor U41380 (N_41380,N_41039,N_41210);
and U41381 (N_41381,N_41043,N_41116);
xnor U41382 (N_41382,N_41095,N_41180);
nor U41383 (N_41383,N_41127,N_41159);
xor U41384 (N_41384,N_41007,N_41117);
nand U41385 (N_41385,N_41024,N_41089);
xor U41386 (N_41386,N_41184,N_41095);
xnor U41387 (N_41387,N_41096,N_41063);
and U41388 (N_41388,N_41070,N_41068);
and U41389 (N_41389,N_41082,N_41189);
or U41390 (N_41390,N_41089,N_41094);
and U41391 (N_41391,N_41101,N_41110);
and U41392 (N_41392,N_41192,N_41067);
or U41393 (N_41393,N_41108,N_41205);
and U41394 (N_41394,N_41142,N_41015);
nor U41395 (N_41395,N_41182,N_41047);
and U41396 (N_41396,N_41074,N_41006);
or U41397 (N_41397,N_41187,N_41036);
or U41398 (N_41398,N_41249,N_41169);
or U41399 (N_41399,N_41175,N_41222);
nor U41400 (N_41400,N_41215,N_41232);
or U41401 (N_41401,N_41023,N_41191);
xnor U41402 (N_41402,N_41080,N_41220);
nor U41403 (N_41403,N_41091,N_41006);
or U41404 (N_41404,N_41222,N_41193);
and U41405 (N_41405,N_41095,N_41143);
xor U41406 (N_41406,N_41036,N_41200);
and U41407 (N_41407,N_41133,N_41194);
nor U41408 (N_41408,N_41034,N_41020);
nand U41409 (N_41409,N_41177,N_41056);
and U41410 (N_41410,N_41224,N_41129);
xor U41411 (N_41411,N_41029,N_41050);
or U41412 (N_41412,N_41186,N_41052);
or U41413 (N_41413,N_41245,N_41138);
nand U41414 (N_41414,N_41008,N_41126);
and U41415 (N_41415,N_41069,N_41000);
nor U41416 (N_41416,N_41124,N_41025);
xnor U41417 (N_41417,N_41135,N_41148);
nor U41418 (N_41418,N_41211,N_41105);
or U41419 (N_41419,N_41077,N_41016);
xor U41420 (N_41420,N_41011,N_41070);
xor U41421 (N_41421,N_41201,N_41023);
nor U41422 (N_41422,N_41137,N_41015);
nand U41423 (N_41423,N_41083,N_41121);
nand U41424 (N_41424,N_41014,N_41042);
nor U41425 (N_41425,N_41225,N_41039);
or U41426 (N_41426,N_41200,N_41065);
or U41427 (N_41427,N_41186,N_41045);
or U41428 (N_41428,N_41200,N_41016);
nor U41429 (N_41429,N_41197,N_41037);
xnor U41430 (N_41430,N_41187,N_41226);
nand U41431 (N_41431,N_41119,N_41239);
nand U41432 (N_41432,N_41207,N_41087);
nand U41433 (N_41433,N_41058,N_41221);
xor U41434 (N_41434,N_41017,N_41131);
nand U41435 (N_41435,N_41152,N_41057);
xnor U41436 (N_41436,N_41188,N_41049);
or U41437 (N_41437,N_41238,N_41208);
nand U41438 (N_41438,N_41213,N_41133);
nand U41439 (N_41439,N_41171,N_41230);
and U41440 (N_41440,N_41009,N_41011);
xor U41441 (N_41441,N_41121,N_41109);
xnor U41442 (N_41442,N_41148,N_41091);
or U41443 (N_41443,N_41009,N_41091);
nand U41444 (N_41444,N_41050,N_41225);
and U41445 (N_41445,N_41148,N_41196);
xor U41446 (N_41446,N_41160,N_41093);
nor U41447 (N_41447,N_41116,N_41069);
nand U41448 (N_41448,N_41100,N_41051);
and U41449 (N_41449,N_41241,N_41192);
nand U41450 (N_41450,N_41135,N_41249);
or U41451 (N_41451,N_41020,N_41035);
and U41452 (N_41452,N_41153,N_41053);
and U41453 (N_41453,N_41007,N_41161);
or U41454 (N_41454,N_41072,N_41099);
or U41455 (N_41455,N_41181,N_41099);
nor U41456 (N_41456,N_41197,N_41055);
or U41457 (N_41457,N_41191,N_41033);
xnor U41458 (N_41458,N_41236,N_41167);
xor U41459 (N_41459,N_41070,N_41127);
nor U41460 (N_41460,N_41229,N_41093);
nor U41461 (N_41461,N_41200,N_41184);
and U41462 (N_41462,N_41075,N_41172);
nand U41463 (N_41463,N_41244,N_41084);
xnor U41464 (N_41464,N_41244,N_41234);
or U41465 (N_41465,N_41159,N_41156);
or U41466 (N_41466,N_41199,N_41080);
xor U41467 (N_41467,N_41226,N_41136);
xnor U41468 (N_41468,N_41029,N_41074);
and U41469 (N_41469,N_41109,N_41027);
xnor U41470 (N_41470,N_41115,N_41168);
and U41471 (N_41471,N_41101,N_41025);
xor U41472 (N_41472,N_41113,N_41043);
xnor U41473 (N_41473,N_41019,N_41095);
or U41474 (N_41474,N_41053,N_41176);
xnor U41475 (N_41475,N_41004,N_41075);
nor U41476 (N_41476,N_41170,N_41057);
or U41477 (N_41477,N_41046,N_41140);
nand U41478 (N_41478,N_41237,N_41148);
nor U41479 (N_41479,N_41164,N_41074);
and U41480 (N_41480,N_41176,N_41124);
nor U41481 (N_41481,N_41130,N_41185);
and U41482 (N_41482,N_41105,N_41169);
and U41483 (N_41483,N_41099,N_41192);
nor U41484 (N_41484,N_41064,N_41067);
nor U41485 (N_41485,N_41224,N_41013);
or U41486 (N_41486,N_41225,N_41112);
nand U41487 (N_41487,N_41016,N_41136);
xnor U41488 (N_41488,N_41192,N_41100);
and U41489 (N_41489,N_41050,N_41005);
or U41490 (N_41490,N_41211,N_41196);
nor U41491 (N_41491,N_41104,N_41022);
xnor U41492 (N_41492,N_41127,N_41240);
nor U41493 (N_41493,N_41236,N_41201);
nor U41494 (N_41494,N_41079,N_41049);
xnor U41495 (N_41495,N_41034,N_41155);
nand U41496 (N_41496,N_41101,N_41247);
nor U41497 (N_41497,N_41231,N_41235);
nand U41498 (N_41498,N_41158,N_41128);
nand U41499 (N_41499,N_41094,N_41165);
nand U41500 (N_41500,N_41272,N_41430);
or U41501 (N_41501,N_41390,N_41377);
nor U41502 (N_41502,N_41496,N_41270);
nand U41503 (N_41503,N_41266,N_41352);
xor U41504 (N_41504,N_41354,N_41326);
nor U41505 (N_41505,N_41321,N_41252);
xnor U41506 (N_41506,N_41314,N_41358);
nor U41507 (N_41507,N_41482,N_41269);
nor U41508 (N_41508,N_41435,N_41459);
and U41509 (N_41509,N_41399,N_41389);
and U41510 (N_41510,N_41294,N_41476);
or U41511 (N_41511,N_41264,N_41422);
xnor U41512 (N_41512,N_41299,N_41285);
or U41513 (N_41513,N_41401,N_41451);
xor U41514 (N_41514,N_41295,N_41356);
nor U41515 (N_41515,N_41472,N_41473);
xor U41516 (N_41516,N_41478,N_41268);
nor U41517 (N_41517,N_41336,N_41379);
nor U41518 (N_41518,N_41380,N_41384);
or U41519 (N_41519,N_41406,N_41421);
xor U41520 (N_41520,N_41329,N_41488);
and U41521 (N_41521,N_41259,N_41411);
or U41522 (N_41522,N_41431,N_41405);
nand U41523 (N_41523,N_41307,N_41479);
nand U41524 (N_41524,N_41491,N_41480);
nand U41525 (N_41525,N_41368,N_41466);
or U41526 (N_41526,N_41310,N_41357);
nor U41527 (N_41527,N_41391,N_41267);
xor U41528 (N_41528,N_41484,N_41322);
nand U41529 (N_41529,N_41372,N_41386);
nand U41530 (N_41530,N_41395,N_41412);
nand U41531 (N_41531,N_41427,N_41457);
nor U41532 (N_41532,N_41425,N_41424);
nor U41533 (N_41533,N_41319,N_41438);
xnor U41534 (N_41534,N_41261,N_41385);
or U41535 (N_41535,N_41446,N_41359);
nand U41536 (N_41536,N_41463,N_41419);
nand U41537 (N_41537,N_41392,N_41366);
xor U41538 (N_41538,N_41256,N_41464);
nor U41539 (N_41539,N_41426,N_41330);
xnor U41540 (N_41540,N_41339,N_41481);
or U41541 (N_41541,N_41304,N_41263);
or U41542 (N_41542,N_41404,N_41400);
or U41543 (N_41543,N_41346,N_41495);
and U41544 (N_41544,N_41283,N_41323);
nand U41545 (N_41545,N_41290,N_41287);
nor U41546 (N_41546,N_41442,N_41475);
nor U41547 (N_41547,N_41292,N_41331);
and U41548 (N_41548,N_41301,N_41351);
nand U41549 (N_41549,N_41432,N_41350);
nand U41550 (N_41550,N_41394,N_41460);
nor U41551 (N_41551,N_41362,N_41369);
nor U41552 (N_41552,N_41461,N_41393);
nor U41553 (N_41553,N_41361,N_41276);
and U41554 (N_41554,N_41251,N_41387);
nand U41555 (N_41555,N_41467,N_41429);
xor U41556 (N_41556,N_41250,N_41289);
xnor U41557 (N_41557,N_41277,N_41309);
nor U41558 (N_41558,N_41347,N_41338);
or U41559 (N_41559,N_41373,N_41408);
or U41560 (N_41560,N_41293,N_41410);
nand U41561 (N_41561,N_41344,N_41443);
nor U41562 (N_41562,N_41273,N_41317);
xor U41563 (N_41563,N_41282,N_41334);
and U41564 (N_41564,N_41291,N_41493);
and U41565 (N_41565,N_41341,N_41271);
and U41566 (N_41566,N_41397,N_41448);
nor U41567 (N_41567,N_41388,N_41367);
nand U41568 (N_41568,N_41279,N_41418);
nand U41569 (N_41569,N_41376,N_41409);
and U41570 (N_41570,N_41364,N_41474);
and U41571 (N_41571,N_41305,N_41253);
and U41572 (N_41572,N_41349,N_41313);
and U41573 (N_41573,N_41477,N_41320);
and U41574 (N_41574,N_41437,N_41257);
nor U41575 (N_41575,N_41444,N_41274);
and U41576 (N_41576,N_41449,N_41306);
or U41577 (N_41577,N_41447,N_41492);
or U41578 (N_41578,N_41468,N_41343);
or U41579 (N_41579,N_41450,N_41497);
xnor U41580 (N_41580,N_41433,N_41355);
nand U41581 (N_41581,N_41316,N_41416);
and U41582 (N_41582,N_41284,N_41265);
nand U41583 (N_41583,N_41396,N_41436);
nand U41584 (N_41584,N_41494,N_41469);
nor U41585 (N_41585,N_41365,N_41445);
xor U41586 (N_41586,N_41363,N_41303);
or U41587 (N_41587,N_41428,N_41337);
and U41588 (N_41588,N_41381,N_41402);
nor U41589 (N_41589,N_41378,N_41453);
or U41590 (N_41590,N_41286,N_41383);
nand U41591 (N_41591,N_41483,N_41403);
xor U41592 (N_41592,N_41420,N_41258);
or U41593 (N_41593,N_41324,N_41455);
nor U41594 (N_41594,N_41281,N_41414);
nand U41595 (N_41595,N_41333,N_41439);
xor U41596 (N_41596,N_41486,N_41327);
or U41597 (N_41597,N_41452,N_41441);
nor U41598 (N_41598,N_41311,N_41255);
nor U41599 (N_41599,N_41318,N_41315);
nor U41600 (N_41600,N_41465,N_41296);
and U41601 (N_41601,N_41454,N_41360);
xnor U41602 (N_41602,N_41374,N_41417);
nor U41603 (N_41603,N_41325,N_41288);
or U41604 (N_41604,N_41485,N_41382);
nand U41605 (N_41605,N_41300,N_41302);
or U41606 (N_41606,N_41348,N_41275);
or U41607 (N_41607,N_41370,N_41470);
nor U41608 (N_41608,N_41280,N_41345);
xnor U41609 (N_41609,N_41456,N_41413);
or U41610 (N_41610,N_41462,N_41340);
or U41611 (N_41611,N_41332,N_41254);
and U41612 (N_41612,N_41499,N_41407);
or U41613 (N_41613,N_41440,N_41375);
and U41614 (N_41614,N_41498,N_41260);
nand U41615 (N_41615,N_41353,N_41415);
xor U41616 (N_41616,N_41423,N_41371);
nand U41617 (N_41617,N_41490,N_41312);
nand U41618 (N_41618,N_41458,N_41298);
and U41619 (N_41619,N_41297,N_41328);
or U41620 (N_41620,N_41398,N_41335);
xnor U41621 (N_41621,N_41342,N_41471);
nand U41622 (N_41622,N_41434,N_41278);
xor U41623 (N_41623,N_41489,N_41262);
nor U41624 (N_41624,N_41308,N_41487);
nor U41625 (N_41625,N_41327,N_41416);
nor U41626 (N_41626,N_41498,N_41487);
nor U41627 (N_41627,N_41305,N_41429);
or U41628 (N_41628,N_41412,N_41465);
or U41629 (N_41629,N_41449,N_41432);
nor U41630 (N_41630,N_41338,N_41375);
and U41631 (N_41631,N_41440,N_41258);
nor U41632 (N_41632,N_41477,N_41316);
nor U41633 (N_41633,N_41262,N_41305);
or U41634 (N_41634,N_41464,N_41283);
and U41635 (N_41635,N_41344,N_41270);
xnor U41636 (N_41636,N_41415,N_41465);
xnor U41637 (N_41637,N_41479,N_41257);
nand U41638 (N_41638,N_41420,N_41484);
nand U41639 (N_41639,N_41481,N_41423);
or U41640 (N_41640,N_41487,N_41439);
nor U41641 (N_41641,N_41493,N_41283);
and U41642 (N_41642,N_41270,N_41323);
or U41643 (N_41643,N_41447,N_41348);
and U41644 (N_41644,N_41270,N_41299);
xor U41645 (N_41645,N_41277,N_41326);
or U41646 (N_41646,N_41458,N_41423);
and U41647 (N_41647,N_41269,N_41499);
nor U41648 (N_41648,N_41333,N_41470);
and U41649 (N_41649,N_41489,N_41334);
nor U41650 (N_41650,N_41475,N_41280);
or U41651 (N_41651,N_41437,N_41259);
nor U41652 (N_41652,N_41463,N_41302);
nand U41653 (N_41653,N_41485,N_41333);
and U41654 (N_41654,N_41397,N_41336);
or U41655 (N_41655,N_41482,N_41456);
nor U41656 (N_41656,N_41429,N_41339);
xnor U41657 (N_41657,N_41315,N_41266);
nand U41658 (N_41658,N_41428,N_41446);
nor U41659 (N_41659,N_41374,N_41307);
and U41660 (N_41660,N_41420,N_41401);
or U41661 (N_41661,N_41413,N_41304);
nand U41662 (N_41662,N_41338,N_41414);
nand U41663 (N_41663,N_41342,N_41460);
nor U41664 (N_41664,N_41474,N_41352);
or U41665 (N_41665,N_41439,N_41465);
nand U41666 (N_41666,N_41293,N_41475);
nand U41667 (N_41667,N_41493,N_41254);
xor U41668 (N_41668,N_41455,N_41292);
nor U41669 (N_41669,N_41333,N_41440);
and U41670 (N_41670,N_41252,N_41296);
nor U41671 (N_41671,N_41486,N_41458);
nand U41672 (N_41672,N_41471,N_41367);
or U41673 (N_41673,N_41327,N_41274);
nor U41674 (N_41674,N_41369,N_41399);
nor U41675 (N_41675,N_41382,N_41311);
or U41676 (N_41676,N_41423,N_41392);
and U41677 (N_41677,N_41358,N_41300);
nor U41678 (N_41678,N_41459,N_41451);
nor U41679 (N_41679,N_41357,N_41382);
nor U41680 (N_41680,N_41289,N_41357);
nand U41681 (N_41681,N_41437,N_41302);
nor U41682 (N_41682,N_41342,N_41275);
or U41683 (N_41683,N_41400,N_41405);
and U41684 (N_41684,N_41285,N_41338);
and U41685 (N_41685,N_41446,N_41385);
or U41686 (N_41686,N_41427,N_41323);
or U41687 (N_41687,N_41295,N_41405);
xor U41688 (N_41688,N_41435,N_41306);
and U41689 (N_41689,N_41408,N_41276);
nor U41690 (N_41690,N_41357,N_41323);
xnor U41691 (N_41691,N_41443,N_41490);
or U41692 (N_41692,N_41490,N_41410);
nand U41693 (N_41693,N_41362,N_41456);
or U41694 (N_41694,N_41271,N_41472);
nor U41695 (N_41695,N_41330,N_41349);
or U41696 (N_41696,N_41421,N_41432);
or U41697 (N_41697,N_41388,N_41273);
and U41698 (N_41698,N_41462,N_41369);
and U41699 (N_41699,N_41361,N_41409);
nor U41700 (N_41700,N_41351,N_41287);
nand U41701 (N_41701,N_41302,N_41416);
nor U41702 (N_41702,N_41398,N_41261);
or U41703 (N_41703,N_41339,N_41257);
nand U41704 (N_41704,N_41474,N_41399);
or U41705 (N_41705,N_41308,N_41419);
or U41706 (N_41706,N_41491,N_41300);
xor U41707 (N_41707,N_41302,N_41460);
or U41708 (N_41708,N_41361,N_41330);
and U41709 (N_41709,N_41342,N_41440);
xor U41710 (N_41710,N_41497,N_41496);
nor U41711 (N_41711,N_41401,N_41380);
xnor U41712 (N_41712,N_41295,N_41421);
nor U41713 (N_41713,N_41480,N_41401);
or U41714 (N_41714,N_41347,N_41361);
nand U41715 (N_41715,N_41250,N_41309);
nor U41716 (N_41716,N_41485,N_41330);
or U41717 (N_41717,N_41465,N_41485);
nor U41718 (N_41718,N_41305,N_41414);
and U41719 (N_41719,N_41256,N_41373);
or U41720 (N_41720,N_41262,N_41389);
nor U41721 (N_41721,N_41353,N_41387);
or U41722 (N_41722,N_41429,N_41259);
nand U41723 (N_41723,N_41321,N_41434);
and U41724 (N_41724,N_41329,N_41362);
nor U41725 (N_41725,N_41447,N_41459);
and U41726 (N_41726,N_41255,N_41375);
nand U41727 (N_41727,N_41346,N_41338);
or U41728 (N_41728,N_41298,N_41495);
or U41729 (N_41729,N_41337,N_41341);
nand U41730 (N_41730,N_41318,N_41474);
xnor U41731 (N_41731,N_41426,N_41457);
nand U41732 (N_41732,N_41290,N_41406);
nand U41733 (N_41733,N_41317,N_41406);
nor U41734 (N_41734,N_41318,N_41468);
nand U41735 (N_41735,N_41254,N_41305);
xnor U41736 (N_41736,N_41333,N_41357);
or U41737 (N_41737,N_41498,N_41332);
or U41738 (N_41738,N_41419,N_41251);
or U41739 (N_41739,N_41493,N_41297);
and U41740 (N_41740,N_41353,N_41354);
or U41741 (N_41741,N_41443,N_41432);
or U41742 (N_41742,N_41423,N_41289);
nand U41743 (N_41743,N_41439,N_41365);
xnor U41744 (N_41744,N_41291,N_41392);
and U41745 (N_41745,N_41489,N_41282);
nor U41746 (N_41746,N_41343,N_41293);
nor U41747 (N_41747,N_41332,N_41370);
nand U41748 (N_41748,N_41480,N_41355);
nor U41749 (N_41749,N_41421,N_41262);
or U41750 (N_41750,N_41704,N_41621);
or U41751 (N_41751,N_41510,N_41720);
or U41752 (N_41752,N_41663,N_41569);
nand U41753 (N_41753,N_41733,N_41718);
nand U41754 (N_41754,N_41624,N_41698);
and U41755 (N_41755,N_41532,N_41725);
or U41756 (N_41756,N_41578,N_41668);
and U41757 (N_41757,N_41575,N_41700);
nand U41758 (N_41758,N_41584,N_41640);
or U41759 (N_41759,N_41596,N_41722);
nand U41760 (N_41760,N_41664,N_41531);
and U41761 (N_41761,N_41709,N_41526);
xor U41762 (N_41762,N_41561,N_41748);
and U41763 (N_41763,N_41636,N_41551);
or U41764 (N_41764,N_41630,N_41628);
nand U41765 (N_41765,N_41649,N_41742);
nand U41766 (N_41766,N_41544,N_41588);
and U41767 (N_41767,N_41604,N_41629);
xor U41768 (N_41768,N_41595,N_41602);
xnor U41769 (N_41769,N_41574,N_41728);
nand U41770 (N_41770,N_41708,N_41688);
or U41771 (N_41771,N_41659,N_41502);
or U41772 (N_41772,N_41557,N_41723);
and U41773 (N_41773,N_41714,N_41665);
nand U41774 (N_41774,N_41740,N_41650);
nand U41775 (N_41775,N_41599,N_41731);
nor U41776 (N_41776,N_41506,N_41730);
or U41777 (N_41777,N_41517,N_41616);
nand U41778 (N_41778,N_41519,N_41556);
and U41779 (N_41779,N_41552,N_41514);
nor U41780 (N_41780,N_41530,N_41535);
xor U41781 (N_41781,N_41673,N_41712);
or U41782 (N_41782,N_41686,N_41738);
nor U41783 (N_41783,N_41706,N_41583);
or U41784 (N_41784,N_41560,N_41625);
and U41785 (N_41785,N_41694,N_41641);
nor U41786 (N_41786,N_41626,N_41562);
nand U41787 (N_41787,N_41726,N_41633);
nor U41788 (N_41788,N_41540,N_41503);
nand U41789 (N_41789,N_41538,N_41555);
or U41790 (N_41790,N_41716,N_41702);
nand U41791 (N_41791,N_41658,N_41548);
and U41792 (N_41792,N_41594,N_41539);
xnor U41793 (N_41793,N_41682,N_41642);
xnor U41794 (N_41794,N_41715,N_41719);
xor U41795 (N_41795,N_41666,N_41500);
or U41796 (N_41796,N_41597,N_41568);
and U41797 (N_41797,N_41573,N_41746);
nand U41798 (N_41798,N_41680,N_41611);
nor U41799 (N_41799,N_41581,N_41735);
nor U41800 (N_41800,N_41684,N_41580);
and U41801 (N_41801,N_41515,N_41732);
and U41802 (N_41802,N_41657,N_41729);
and U41803 (N_41803,N_41533,N_41632);
nand U41804 (N_41804,N_41634,N_41612);
or U41805 (N_41805,N_41577,N_41504);
xor U41806 (N_41806,N_41525,N_41727);
nor U41807 (N_41807,N_41615,N_41691);
and U41808 (N_41808,N_41619,N_41745);
and U41809 (N_41809,N_41547,N_41687);
or U41810 (N_41810,N_41553,N_41541);
xnor U41811 (N_41811,N_41603,N_41695);
and U41812 (N_41812,N_41737,N_41608);
nand U41813 (N_41813,N_41674,N_41651);
and U41814 (N_41814,N_41661,N_41711);
or U41815 (N_41815,N_41549,N_41647);
or U41816 (N_41816,N_41516,N_41672);
xnor U41817 (N_41817,N_41703,N_41523);
xor U41818 (N_41818,N_41618,N_41554);
or U41819 (N_41819,N_41724,N_41635);
xor U41820 (N_41820,N_41509,N_41550);
and U41821 (N_41821,N_41536,N_41566);
xnor U41822 (N_41822,N_41582,N_41613);
nand U41823 (N_41823,N_41591,N_41522);
xor U41824 (N_41824,N_41590,N_41736);
or U41825 (N_41825,N_41571,N_41690);
xnor U41826 (N_41826,N_41570,N_41652);
nor U41827 (N_41827,N_41564,N_41558);
nand U41828 (N_41828,N_41653,N_41643);
nand U41829 (N_41829,N_41678,N_41559);
nor U41830 (N_41830,N_41697,N_41639);
nor U41831 (N_41831,N_41614,N_41617);
xnor U41832 (N_41832,N_41671,N_41610);
xor U41833 (N_41833,N_41592,N_41622);
nand U41834 (N_41834,N_41741,N_41524);
and U41835 (N_41835,N_41676,N_41521);
nor U41836 (N_41836,N_41681,N_41601);
nor U41837 (N_41837,N_41670,N_41572);
or U41838 (N_41838,N_41696,N_41699);
xor U41839 (N_41839,N_41627,N_41623);
nor U41840 (N_41840,N_41645,N_41511);
xnor U41841 (N_41841,N_41537,N_41638);
and U41842 (N_41842,N_41543,N_41508);
xnor U41843 (N_41843,N_41589,N_41631);
xnor U41844 (N_41844,N_41646,N_41528);
xor U41845 (N_41845,N_41563,N_41520);
and U41846 (N_41846,N_41529,N_41744);
and U41847 (N_41847,N_41576,N_41606);
or U41848 (N_41848,N_41586,N_41689);
nand U41849 (N_41849,N_41713,N_41701);
and U41850 (N_41850,N_41734,N_41542);
nand U41851 (N_41851,N_41598,N_41512);
or U41852 (N_41852,N_41743,N_41667);
or U41853 (N_41853,N_41747,N_41721);
and U41854 (N_41854,N_41505,N_41707);
or U41855 (N_41855,N_41644,N_41705);
or U41856 (N_41856,N_41565,N_41679);
nand U41857 (N_41857,N_41749,N_41546);
nand U41858 (N_41858,N_41677,N_41654);
nand U41859 (N_41859,N_41739,N_41501);
xor U41860 (N_41860,N_41620,N_41710);
nand U41861 (N_41861,N_41579,N_41593);
xnor U41862 (N_41862,N_41567,N_41655);
xor U41863 (N_41863,N_41692,N_41669);
or U41864 (N_41864,N_41637,N_41587);
and U41865 (N_41865,N_41609,N_41607);
and U41866 (N_41866,N_41717,N_41648);
nor U41867 (N_41867,N_41600,N_41685);
nor U41868 (N_41868,N_41534,N_41683);
and U41869 (N_41869,N_41662,N_41527);
or U41870 (N_41870,N_41675,N_41518);
and U41871 (N_41871,N_41660,N_41693);
nand U41872 (N_41872,N_41605,N_41545);
nand U41873 (N_41873,N_41585,N_41507);
nor U41874 (N_41874,N_41513,N_41656);
nand U41875 (N_41875,N_41513,N_41643);
nand U41876 (N_41876,N_41567,N_41709);
or U41877 (N_41877,N_41508,N_41542);
nand U41878 (N_41878,N_41543,N_41688);
nor U41879 (N_41879,N_41613,N_41599);
and U41880 (N_41880,N_41571,N_41505);
nand U41881 (N_41881,N_41671,N_41528);
nand U41882 (N_41882,N_41648,N_41632);
and U41883 (N_41883,N_41696,N_41509);
xnor U41884 (N_41884,N_41604,N_41594);
nand U41885 (N_41885,N_41613,N_41606);
nor U41886 (N_41886,N_41607,N_41635);
and U41887 (N_41887,N_41564,N_41723);
and U41888 (N_41888,N_41700,N_41688);
nor U41889 (N_41889,N_41573,N_41555);
xor U41890 (N_41890,N_41731,N_41566);
nor U41891 (N_41891,N_41590,N_41720);
xor U41892 (N_41892,N_41686,N_41635);
or U41893 (N_41893,N_41694,N_41540);
nor U41894 (N_41894,N_41591,N_41679);
and U41895 (N_41895,N_41625,N_41681);
xor U41896 (N_41896,N_41674,N_41596);
and U41897 (N_41897,N_41529,N_41675);
or U41898 (N_41898,N_41667,N_41685);
or U41899 (N_41899,N_41654,N_41544);
or U41900 (N_41900,N_41666,N_41692);
nor U41901 (N_41901,N_41692,N_41564);
nor U41902 (N_41902,N_41520,N_41602);
nor U41903 (N_41903,N_41558,N_41694);
xor U41904 (N_41904,N_41636,N_41594);
and U41905 (N_41905,N_41638,N_41644);
nand U41906 (N_41906,N_41720,N_41619);
nor U41907 (N_41907,N_41676,N_41505);
and U41908 (N_41908,N_41506,N_41594);
nand U41909 (N_41909,N_41603,N_41719);
nand U41910 (N_41910,N_41728,N_41528);
or U41911 (N_41911,N_41721,N_41677);
nand U41912 (N_41912,N_41697,N_41660);
or U41913 (N_41913,N_41602,N_41509);
or U41914 (N_41914,N_41577,N_41697);
or U41915 (N_41915,N_41580,N_41602);
nand U41916 (N_41916,N_41699,N_41705);
nand U41917 (N_41917,N_41642,N_41541);
nand U41918 (N_41918,N_41708,N_41594);
and U41919 (N_41919,N_41596,N_41671);
xnor U41920 (N_41920,N_41555,N_41687);
nor U41921 (N_41921,N_41591,N_41613);
nor U41922 (N_41922,N_41649,N_41625);
xor U41923 (N_41923,N_41571,N_41692);
nor U41924 (N_41924,N_41589,N_41703);
or U41925 (N_41925,N_41656,N_41569);
or U41926 (N_41926,N_41609,N_41635);
xnor U41927 (N_41927,N_41655,N_41536);
nand U41928 (N_41928,N_41653,N_41667);
nand U41929 (N_41929,N_41704,N_41638);
nand U41930 (N_41930,N_41693,N_41641);
nor U41931 (N_41931,N_41707,N_41574);
and U41932 (N_41932,N_41565,N_41579);
and U41933 (N_41933,N_41517,N_41509);
and U41934 (N_41934,N_41529,N_41686);
nor U41935 (N_41935,N_41552,N_41550);
nand U41936 (N_41936,N_41510,N_41664);
nand U41937 (N_41937,N_41581,N_41644);
xor U41938 (N_41938,N_41658,N_41743);
nor U41939 (N_41939,N_41714,N_41716);
xnor U41940 (N_41940,N_41520,N_41638);
xor U41941 (N_41941,N_41651,N_41745);
nand U41942 (N_41942,N_41548,N_41674);
nand U41943 (N_41943,N_41677,N_41515);
xnor U41944 (N_41944,N_41566,N_41703);
nor U41945 (N_41945,N_41740,N_41658);
and U41946 (N_41946,N_41748,N_41721);
or U41947 (N_41947,N_41685,N_41714);
or U41948 (N_41948,N_41545,N_41716);
nand U41949 (N_41949,N_41612,N_41501);
xnor U41950 (N_41950,N_41555,N_41698);
and U41951 (N_41951,N_41591,N_41620);
nor U41952 (N_41952,N_41590,N_41730);
xor U41953 (N_41953,N_41566,N_41591);
nor U41954 (N_41954,N_41566,N_41556);
and U41955 (N_41955,N_41506,N_41623);
nor U41956 (N_41956,N_41667,N_41529);
nor U41957 (N_41957,N_41516,N_41619);
xor U41958 (N_41958,N_41724,N_41632);
or U41959 (N_41959,N_41690,N_41574);
nand U41960 (N_41960,N_41629,N_41623);
nor U41961 (N_41961,N_41686,N_41570);
nor U41962 (N_41962,N_41607,N_41739);
or U41963 (N_41963,N_41544,N_41690);
xnor U41964 (N_41964,N_41658,N_41566);
or U41965 (N_41965,N_41678,N_41683);
and U41966 (N_41966,N_41703,N_41697);
or U41967 (N_41967,N_41747,N_41695);
nor U41968 (N_41968,N_41542,N_41715);
or U41969 (N_41969,N_41629,N_41620);
or U41970 (N_41970,N_41729,N_41519);
nor U41971 (N_41971,N_41560,N_41572);
or U41972 (N_41972,N_41633,N_41745);
xor U41973 (N_41973,N_41699,N_41647);
and U41974 (N_41974,N_41519,N_41561);
and U41975 (N_41975,N_41744,N_41691);
xor U41976 (N_41976,N_41690,N_41678);
nand U41977 (N_41977,N_41580,N_41605);
nor U41978 (N_41978,N_41645,N_41600);
and U41979 (N_41979,N_41652,N_41589);
xnor U41980 (N_41980,N_41722,N_41646);
nand U41981 (N_41981,N_41557,N_41653);
nor U41982 (N_41982,N_41513,N_41683);
nor U41983 (N_41983,N_41526,N_41664);
and U41984 (N_41984,N_41741,N_41588);
or U41985 (N_41985,N_41743,N_41674);
or U41986 (N_41986,N_41530,N_41539);
xor U41987 (N_41987,N_41706,N_41516);
or U41988 (N_41988,N_41742,N_41703);
xnor U41989 (N_41989,N_41569,N_41592);
nand U41990 (N_41990,N_41561,N_41679);
and U41991 (N_41991,N_41512,N_41677);
nand U41992 (N_41992,N_41501,N_41500);
xor U41993 (N_41993,N_41693,N_41705);
and U41994 (N_41994,N_41623,N_41651);
nor U41995 (N_41995,N_41694,N_41667);
xnor U41996 (N_41996,N_41500,N_41627);
xnor U41997 (N_41997,N_41743,N_41702);
or U41998 (N_41998,N_41558,N_41603);
nor U41999 (N_41999,N_41717,N_41746);
or U42000 (N_42000,N_41868,N_41875);
nor U42001 (N_42001,N_41908,N_41975);
nor U42002 (N_42002,N_41825,N_41951);
or U42003 (N_42003,N_41824,N_41981);
nand U42004 (N_42004,N_41986,N_41897);
and U42005 (N_42005,N_41842,N_41906);
or U42006 (N_42006,N_41967,N_41899);
nor U42007 (N_42007,N_41773,N_41921);
xnor U42008 (N_42008,N_41954,N_41856);
or U42009 (N_42009,N_41940,N_41785);
or U42010 (N_42010,N_41929,N_41833);
or U42011 (N_42011,N_41896,N_41926);
xor U42012 (N_42012,N_41984,N_41861);
or U42013 (N_42013,N_41871,N_41881);
and U42014 (N_42014,N_41779,N_41783);
nor U42015 (N_42015,N_41752,N_41907);
xor U42016 (N_42016,N_41969,N_41877);
and U42017 (N_42017,N_41958,N_41862);
xor U42018 (N_42018,N_41972,N_41786);
xor U42019 (N_42019,N_41965,N_41860);
xor U42020 (N_42020,N_41953,N_41803);
or U42021 (N_42021,N_41855,N_41777);
nor U42022 (N_42022,N_41794,N_41928);
nand U42023 (N_42023,N_41775,N_41971);
xnor U42024 (N_42024,N_41863,N_41959);
xor U42025 (N_42025,N_41835,N_41859);
nand U42026 (N_42026,N_41991,N_41962);
nand U42027 (N_42027,N_41822,N_41820);
nand U42028 (N_42028,N_41780,N_41903);
and U42029 (N_42029,N_41900,N_41823);
nor U42030 (N_42030,N_41884,N_41767);
nand U42031 (N_42031,N_41916,N_41927);
xor U42032 (N_42032,N_41790,N_41996);
nor U42033 (N_42033,N_41994,N_41932);
or U42034 (N_42034,N_41924,N_41836);
and U42035 (N_42035,N_41768,N_41826);
and U42036 (N_42036,N_41944,N_41804);
nor U42037 (N_42037,N_41778,N_41821);
nor U42038 (N_42038,N_41960,N_41891);
and U42039 (N_42039,N_41978,N_41901);
nor U42040 (N_42040,N_41809,N_41925);
nor U42041 (N_42041,N_41890,N_41867);
nand U42042 (N_42042,N_41769,N_41930);
and U42043 (N_42043,N_41755,N_41808);
nor U42044 (N_42044,N_41968,N_41934);
nand U42045 (N_42045,N_41964,N_41914);
or U42046 (N_42046,N_41915,N_41760);
xnor U42047 (N_42047,N_41771,N_41963);
nor U42048 (N_42048,N_41789,N_41936);
and U42049 (N_42049,N_41750,N_41910);
and U42050 (N_42050,N_41883,N_41923);
or U42051 (N_42051,N_41957,N_41933);
xnor U42052 (N_42052,N_41788,N_41818);
nor U42053 (N_42053,N_41852,N_41799);
and U42054 (N_42054,N_41947,N_41840);
xnor U42055 (N_42055,N_41844,N_41917);
nand U42056 (N_42056,N_41931,N_41970);
xor U42057 (N_42057,N_41829,N_41977);
or U42058 (N_42058,N_41797,N_41961);
nor U42059 (N_42059,N_41943,N_41816);
nand U42060 (N_42060,N_41843,N_41999);
nor U42061 (N_42061,N_41873,N_41879);
nor U42062 (N_42062,N_41810,N_41819);
xor U42063 (N_42063,N_41827,N_41812);
nand U42064 (N_42064,N_41913,N_41832);
xor U42065 (N_42065,N_41898,N_41857);
nand U42066 (N_42066,N_41973,N_41802);
and U42067 (N_42067,N_41938,N_41974);
and U42068 (N_42068,N_41893,N_41949);
and U42069 (N_42069,N_41866,N_41865);
xnor U42070 (N_42070,N_41922,N_41800);
nor U42071 (N_42071,N_41992,N_41987);
nand U42072 (N_42072,N_41830,N_41754);
nor U42073 (N_42073,N_41990,N_41945);
or U42074 (N_42074,N_41904,N_41853);
or U42075 (N_42075,N_41806,N_41811);
xor U42076 (N_42076,N_41870,N_41849);
nand U42077 (N_42077,N_41985,N_41782);
or U42078 (N_42078,N_41937,N_41766);
xnor U42079 (N_42079,N_41791,N_41885);
nor U42080 (N_42080,N_41846,N_41792);
nor U42081 (N_42081,N_41787,N_41774);
nand U42082 (N_42082,N_41765,N_41858);
nor U42083 (N_42083,N_41876,N_41854);
or U42084 (N_42084,N_41874,N_41770);
xor U42085 (N_42085,N_41993,N_41887);
nand U42086 (N_42086,N_41894,N_41864);
and U42087 (N_42087,N_41998,N_41839);
and U42088 (N_42088,N_41761,N_41828);
nand U42089 (N_42089,N_41989,N_41946);
xor U42090 (N_42090,N_41912,N_41805);
or U42091 (N_42091,N_41952,N_41848);
nand U42092 (N_42092,N_41942,N_41880);
or U42093 (N_42093,N_41831,N_41872);
xnor U42094 (N_42094,N_41988,N_41888);
nand U42095 (N_42095,N_41753,N_41756);
and U42096 (N_42096,N_41918,N_41841);
and U42097 (N_42097,N_41758,N_41776);
nor U42098 (N_42098,N_41966,N_41911);
nand U42099 (N_42099,N_41935,N_41997);
nand U42100 (N_42100,N_41847,N_41793);
nor U42101 (N_42101,N_41878,N_41781);
or U42102 (N_42102,N_41834,N_41905);
nor U42103 (N_42103,N_41851,N_41979);
nor U42104 (N_42104,N_41995,N_41882);
or U42105 (N_42105,N_41950,N_41801);
and U42106 (N_42106,N_41902,N_41895);
nor U42107 (N_42107,N_41807,N_41980);
or U42108 (N_42108,N_41798,N_41976);
nand U42109 (N_42109,N_41762,N_41757);
or U42110 (N_42110,N_41815,N_41814);
xnor U42111 (N_42111,N_41796,N_41982);
or U42112 (N_42112,N_41919,N_41941);
or U42113 (N_42113,N_41948,N_41751);
nor U42114 (N_42114,N_41784,N_41763);
xor U42115 (N_42115,N_41772,N_41909);
and U42116 (N_42116,N_41813,N_41759);
nor U42117 (N_42117,N_41886,N_41817);
nor U42118 (N_42118,N_41850,N_41983);
nor U42119 (N_42119,N_41869,N_41955);
or U42120 (N_42120,N_41795,N_41939);
or U42121 (N_42121,N_41956,N_41838);
or U42122 (N_42122,N_41889,N_41764);
nand U42123 (N_42123,N_41837,N_41892);
or U42124 (N_42124,N_41845,N_41920);
xor U42125 (N_42125,N_41780,N_41910);
xor U42126 (N_42126,N_41912,N_41967);
xor U42127 (N_42127,N_41858,N_41951);
or U42128 (N_42128,N_41832,N_41863);
xnor U42129 (N_42129,N_41985,N_41805);
xnor U42130 (N_42130,N_41966,N_41753);
xnor U42131 (N_42131,N_41823,N_41846);
and U42132 (N_42132,N_41885,N_41905);
xor U42133 (N_42133,N_41774,N_41864);
and U42134 (N_42134,N_41866,N_41901);
xnor U42135 (N_42135,N_41755,N_41788);
and U42136 (N_42136,N_41955,N_41782);
or U42137 (N_42137,N_41900,N_41847);
nand U42138 (N_42138,N_41999,N_41830);
nor U42139 (N_42139,N_41872,N_41848);
xnor U42140 (N_42140,N_41963,N_41899);
or U42141 (N_42141,N_41783,N_41842);
and U42142 (N_42142,N_41788,N_41784);
nand U42143 (N_42143,N_41868,N_41918);
and U42144 (N_42144,N_41782,N_41874);
nor U42145 (N_42145,N_41860,N_41974);
or U42146 (N_42146,N_41988,N_41931);
and U42147 (N_42147,N_41887,N_41995);
nand U42148 (N_42148,N_41885,N_41952);
nand U42149 (N_42149,N_41866,N_41779);
nor U42150 (N_42150,N_41969,N_41788);
xor U42151 (N_42151,N_41798,N_41810);
xnor U42152 (N_42152,N_41951,N_41980);
and U42153 (N_42153,N_41822,N_41990);
xor U42154 (N_42154,N_41984,N_41953);
xnor U42155 (N_42155,N_41758,N_41988);
xnor U42156 (N_42156,N_41823,N_41770);
and U42157 (N_42157,N_41965,N_41878);
or U42158 (N_42158,N_41881,N_41978);
nor U42159 (N_42159,N_41959,N_41875);
xor U42160 (N_42160,N_41778,N_41957);
or U42161 (N_42161,N_41859,N_41962);
or U42162 (N_42162,N_41887,N_41800);
or U42163 (N_42163,N_41951,N_41927);
nor U42164 (N_42164,N_41899,N_41856);
nand U42165 (N_42165,N_41872,N_41826);
xnor U42166 (N_42166,N_41789,N_41888);
or U42167 (N_42167,N_41941,N_41897);
and U42168 (N_42168,N_41777,N_41841);
and U42169 (N_42169,N_41815,N_41829);
nand U42170 (N_42170,N_41793,N_41764);
nor U42171 (N_42171,N_41817,N_41835);
xnor U42172 (N_42172,N_41995,N_41774);
nor U42173 (N_42173,N_41996,N_41795);
or U42174 (N_42174,N_41777,N_41994);
or U42175 (N_42175,N_41937,N_41841);
nor U42176 (N_42176,N_41783,N_41825);
nor U42177 (N_42177,N_41999,N_41896);
nand U42178 (N_42178,N_41947,N_41807);
xnor U42179 (N_42179,N_41876,N_41886);
nor U42180 (N_42180,N_41983,N_41944);
nand U42181 (N_42181,N_41757,N_41846);
xnor U42182 (N_42182,N_41854,N_41889);
xor U42183 (N_42183,N_41772,N_41962);
and U42184 (N_42184,N_41945,N_41877);
nand U42185 (N_42185,N_41850,N_41852);
or U42186 (N_42186,N_41750,N_41922);
nor U42187 (N_42187,N_41922,N_41894);
nand U42188 (N_42188,N_41796,N_41817);
and U42189 (N_42189,N_41837,N_41855);
or U42190 (N_42190,N_41844,N_41756);
or U42191 (N_42191,N_41779,N_41880);
nor U42192 (N_42192,N_41752,N_41859);
and U42193 (N_42193,N_41903,N_41793);
xor U42194 (N_42194,N_41820,N_41981);
or U42195 (N_42195,N_41802,N_41764);
xnor U42196 (N_42196,N_41948,N_41762);
or U42197 (N_42197,N_41864,N_41965);
and U42198 (N_42198,N_41808,N_41910);
nand U42199 (N_42199,N_41830,N_41757);
and U42200 (N_42200,N_41926,N_41796);
xnor U42201 (N_42201,N_41927,N_41965);
nand U42202 (N_42202,N_41799,N_41905);
xor U42203 (N_42203,N_41885,N_41765);
xnor U42204 (N_42204,N_41832,N_41941);
nor U42205 (N_42205,N_41803,N_41787);
nand U42206 (N_42206,N_41756,N_41953);
and U42207 (N_42207,N_41890,N_41889);
nor U42208 (N_42208,N_41777,N_41853);
or U42209 (N_42209,N_41989,N_41910);
nand U42210 (N_42210,N_41987,N_41902);
nand U42211 (N_42211,N_41849,N_41880);
or U42212 (N_42212,N_41765,N_41842);
nor U42213 (N_42213,N_41814,N_41917);
nand U42214 (N_42214,N_41966,N_41830);
xor U42215 (N_42215,N_41790,N_41997);
nor U42216 (N_42216,N_41903,N_41756);
and U42217 (N_42217,N_41982,N_41893);
and U42218 (N_42218,N_41772,N_41902);
and U42219 (N_42219,N_41995,N_41959);
nand U42220 (N_42220,N_41941,N_41782);
or U42221 (N_42221,N_41784,N_41978);
and U42222 (N_42222,N_41806,N_41755);
nand U42223 (N_42223,N_41930,N_41915);
xor U42224 (N_42224,N_41803,N_41944);
nor U42225 (N_42225,N_41930,N_41880);
nor U42226 (N_42226,N_41875,N_41825);
and U42227 (N_42227,N_41931,N_41844);
nand U42228 (N_42228,N_41758,N_41860);
or U42229 (N_42229,N_41884,N_41949);
or U42230 (N_42230,N_41948,N_41878);
nand U42231 (N_42231,N_41805,N_41928);
or U42232 (N_42232,N_41886,N_41903);
nor U42233 (N_42233,N_41767,N_41811);
nor U42234 (N_42234,N_41963,N_41952);
xor U42235 (N_42235,N_41908,N_41803);
or U42236 (N_42236,N_41945,N_41935);
nor U42237 (N_42237,N_41901,N_41854);
xor U42238 (N_42238,N_41966,N_41824);
or U42239 (N_42239,N_41781,N_41844);
xnor U42240 (N_42240,N_41799,N_41966);
and U42241 (N_42241,N_41751,N_41964);
nor U42242 (N_42242,N_41837,N_41923);
or U42243 (N_42243,N_41950,N_41798);
and U42244 (N_42244,N_41853,N_41831);
and U42245 (N_42245,N_41962,N_41780);
nand U42246 (N_42246,N_41883,N_41880);
nand U42247 (N_42247,N_41927,N_41966);
nor U42248 (N_42248,N_41904,N_41970);
and U42249 (N_42249,N_41780,N_41774);
and U42250 (N_42250,N_42076,N_42039);
or U42251 (N_42251,N_42138,N_42149);
nor U42252 (N_42252,N_42112,N_42164);
xor U42253 (N_42253,N_42163,N_42187);
xor U42254 (N_42254,N_42158,N_42245);
nor U42255 (N_42255,N_42198,N_42231);
nand U42256 (N_42256,N_42229,N_42239);
nand U42257 (N_42257,N_42046,N_42101);
or U42258 (N_42258,N_42055,N_42027);
nand U42259 (N_42259,N_42157,N_42107);
or U42260 (N_42260,N_42233,N_42059);
nand U42261 (N_42261,N_42135,N_42012);
nor U42262 (N_42262,N_42122,N_42143);
and U42263 (N_42263,N_42038,N_42214);
nand U42264 (N_42264,N_42008,N_42051);
and U42265 (N_42265,N_42000,N_42177);
or U42266 (N_42266,N_42095,N_42146);
nor U42267 (N_42267,N_42193,N_42179);
nor U42268 (N_42268,N_42102,N_42105);
nor U42269 (N_42269,N_42232,N_42184);
nand U42270 (N_42270,N_42225,N_42220);
nor U42271 (N_42271,N_42137,N_42224);
and U42272 (N_42272,N_42018,N_42080);
nor U42273 (N_42273,N_42048,N_42007);
nor U42274 (N_42274,N_42026,N_42180);
xnor U42275 (N_42275,N_42049,N_42079);
and U42276 (N_42276,N_42111,N_42081);
or U42277 (N_42277,N_42246,N_42082);
xor U42278 (N_42278,N_42129,N_42170);
xor U42279 (N_42279,N_42036,N_42237);
nor U42280 (N_42280,N_42144,N_42070);
xor U42281 (N_42281,N_42185,N_42052);
or U42282 (N_42282,N_42011,N_42024);
nand U42283 (N_42283,N_42053,N_42096);
and U42284 (N_42284,N_42145,N_42009);
and U42285 (N_42285,N_42010,N_42086);
nand U42286 (N_42286,N_42132,N_42035);
nand U42287 (N_42287,N_42126,N_42114);
nand U42288 (N_42288,N_42094,N_42200);
or U42289 (N_42289,N_42241,N_42002);
or U42290 (N_42290,N_42209,N_42216);
xnor U42291 (N_42291,N_42085,N_42171);
nand U42292 (N_42292,N_42040,N_42175);
and U42293 (N_42293,N_42033,N_42037);
and U42294 (N_42294,N_42062,N_42226);
nor U42295 (N_42295,N_42196,N_42194);
or U42296 (N_42296,N_42019,N_42044);
xor U42297 (N_42297,N_42167,N_42159);
xnor U42298 (N_42298,N_42217,N_42067);
or U42299 (N_42299,N_42211,N_42188);
nand U42300 (N_42300,N_42092,N_42064);
and U42301 (N_42301,N_42191,N_42030);
nand U42302 (N_42302,N_42243,N_42091);
or U42303 (N_42303,N_42134,N_42029);
xor U42304 (N_42304,N_42069,N_42178);
or U42305 (N_42305,N_42238,N_42110);
and U42306 (N_42306,N_42127,N_42093);
or U42307 (N_42307,N_42058,N_42031);
nor U42308 (N_42308,N_42161,N_42025);
xor U42309 (N_42309,N_42150,N_42133);
and U42310 (N_42310,N_42203,N_42223);
xor U42311 (N_42311,N_42020,N_42090);
or U42312 (N_42312,N_42210,N_42130);
nor U42313 (N_42313,N_42097,N_42068);
or U42314 (N_42314,N_42087,N_42156);
nand U42315 (N_42315,N_42100,N_42140);
nand U42316 (N_42316,N_42227,N_42141);
nor U42317 (N_42317,N_42142,N_42181);
xnor U42318 (N_42318,N_42174,N_42098);
or U42319 (N_42319,N_42088,N_42074);
and U42320 (N_42320,N_42199,N_42023);
xor U42321 (N_42321,N_42128,N_42213);
and U42322 (N_42322,N_42115,N_42106);
nor U42323 (N_42323,N_42071,N_42244);
and U42324 (N_42324,N_42065,N_42057);
nand U42325 (N_42325,N_42108,N_42063);
nor U42326 (N_42326,N_42212,N_42022);
and U42327 (N_42327,N_42202,N_42197);
nand U42328 (N_42328,N_42124,N_42054);
and U42329 (N_42329,N_42016,N_42247);
xnor U42330 (N_42330,N_42207,N_42118);
and U42331 (N_42331,N_42152,N_42248);
nor U42332 (N_42332,N_42186,N_42240);
and U42333 (N_42333,N_42183,N_42201);
or U42334 (N_42334,N_42125,N_42249);
xnor U42335 (N_42335,N_42222,N_42168);
or U42336 (N_42336,N_42208,N_42117);
or U42337 (N_42337,N_42236,N_42103);
nand U42338 (N_42338,N_42041,N_42072);
nor U42339 (N_42339,N_42001,N_42113);
or U42340 (N_42340,N_42116,N_42083);
nand U42341 (N_42341,N_42136,N_42195);
nor U42342 (N_42342,N_42078,N_42189);
nor U42343 (N_42343,N_42089,N_42235);
nand U42344 (N_42344,N_42151,N_42148);
xnor U42345 (N_42345,N_42042,N_42034);
nand U42346 (N_42346,N_42073,N_42120);
or U42347 (N_42347,N_42190,N_42160);
nand U42348 (N_42348,N_42119,N_42066);
and U42349 (N_42349,N_42155,N_42215);
nor U42350 (N_42350,N_42099,N_42004);
nor U42351 (N_42351,N_42045,N_42221);
or U42352 (N_42352,N_42165,N_42205);
nor U42353 (N_42353,N_42121,N_42173);
nand U42354 (N_42354,N_42005,N_42003);
or U42355 (N_42355,N_42084,N_42228);
xor U42356 (N_42356,N_42242,N_42230);
and U42357 (N_42357,N_42014,N_42162);
nand U42358 (N_42358,N_42017,N_42050);
and U42359 (N_42359,N_42109,N_42056);
or U42360 (N_42360,N_42153,N_42234);
nor U42361 (N_42361,N_42028,N_42013);
or U42362 (N_42362,N_42032,N_42147);
xor U42363 (N_42363,N_42219,N_42104);
xor U42364 (N_42364,N_42166,N_42139);
xnor U42365 (N_42365,N_42043,N_42172);
or U42366 (N_42366,N_42021,N_42131);
nor U42367 (N_42367,N_42075,N_42060);
and U42368 (N_42368,N_42154,N_42204);
and U42369 (N_42369,N_42169,N_42182);
or U42370 (N_42370,N_42006,N_42077);
xor U42371 (N_42371,N_42176,N_42015);
nand U42372 (N_42372,N_42218,N_42206);
nor U42373 (N_42373,N_42047,N_42061);
nand U42374 (N_42374,N_42192,N_42123);
nand U42375 (N_42375,N_42029,N_42021);
and U42376 (N_42376,N_42013,N_42090);
nor U42377 (N_42377,N_42137,N_42043);
or U42378 (N_42378,N_42071,N_42143);
nor U42379 (N_42379,N_42142,N_42108);
nor U42380 (N_42380,N_42197,N_42237);
or U42381 (N_42381,N_42152,N_42020);
xnor U42382 (N_42382,N_42065,N_42051);
xnor U42383 (N_42383,N_42049,N_42208);
and U42384 (N_42384,N_42094,N_42172);
or U42385 (N_42385,N_42152,N_42071);
nand U42386 (N_42386,N_42022,N_42105);
xor U42387 (N_42387,N_42184,N_42040);
and U42388 (N_42388,N_42191,N_42118);
and U42389 (N_42389,N_42043,N_42023);
nand U42390 (N_42390,N_42137,N_42166);
nor U42391 (N_42391,N_42118,N_42063);
or U42392 (N_42392,N_42181,N_42057);
nand U42393 (N_42393,N_42045,N_42189);
or U42394 (N_42394,N_42079,N_42072);
or U42395 (N_42395,N_42075,N_42189);
xor U42396 (N_42396,N_42064,N_42036);
nor U42397 (N_42397,N_42170,N_42163);
nand U42398 (N_42398,N_42212,N_42248);
or U42399 (N_42399,N_42165,N_42070);
or U42400 (N_42400,N_42073,N_42050);
xor U42401 (N_42401,N_42159,N_42162);
xnor U42402 (N_42402,N_42064,N_42148);
xor U42403 (N_42403,N_42071,N_42183);
xor U42404 (N_42404,N_42062,N_42230);
xor U42405 (N_42405,N_42130,N_42018);
nand U42406 (N_42406,N_42022,N_42205);
xor U42407 (N_42407,N_42092,N_42094);
and U42408 (N_42408,N_42141,N_42043);
xnor U42409 (N_42409,N_42031,N_42217);
nand U42410 (N_42410,N_42201,N_42212);
or U42411 (N_42411,N_42062,N_42196);
and U42412 (N_42412,N_42185,N_42189);
nand U42413 (N_42413,N_42186,N_42203);
nor U42414 (N_42414,N_42198,N_42245);
and U42415 (N_42415,N_42132,N_42103);
and U42416 (N_42416,N_42162,N_42117);
nand U42417 (N_42417,N_42168,N_42050);
nand U42418 (N_42418,N_42087,N_42060);
nand U42419 (N_42419,N_42125,N_42037);
nand U42420 (N_42420,N_42248,N_42163);
or U42421 (N_42421,N_42140,N_42025);
xor U42422 (N_42422,N_42161,N_42121);
nand U42423 (N_42423,N_42121,N_42148);
or U42424 (N_42424,N_42166,N_42152);
nor U42425 (N_42425,N_42244,N_42236);
xor U42426 (N_42426,N_42005,N_42060);
nand U42427 (N_42427,N_42155,N_42082);
nor U42428 (N_42428,N_42097,N_42038);
nor U42429 (N_42429,N_42004,N_42137);
or U42430 (N_42430,N_42228,N_42186);
nor U42431 (N_42431,N_42081,N_42233);
and U42432 (N_42432,N_42025,N_42077);
and U42433 (N_42433,N_42000,N_42171);
xnor U42434 (N_42434,N_42022,N_42095);
and U42435 (N_42435,N_42134,N_42118);
or U42436 (N_42436,N_42135,N_42032);
nand U42437 (N_42437,N_42248,N_42087);
nor U42438 (N_42438,N_42010,N_42098);
or U42439 (N_42439,N_42056,N_42152);
or U42440 (N_42440,N_42018,N_42128);
xnor U42441 (N_42441,N_42046,N_42154);
or U42442 (N_42442,N_42041,N_42200);
nor U42443 (N_42443,N_42167,N_42161);
xor U42444 (N_42444,N_42127,N_42157);
nor U42445 (N_42445,N_42082,N_42106);
nand U42446 (N_42446,N_42070,N_42042);
nand U42447 (N_42447,N_42125,N_42063);
nor U42448 (N_42448,N_42161,N_42140);
or U42449 (N_42449,N_42217,N_42054);
xnor U42450 (N_42450,N_42232,N_42091);
or U42451 (N_42451,N_42000,N_42106);
and U42452 (N_42452,N_42203,N_42216);
and U42453 (N_42453,N_42047,N_42213);
nand U42454 (N_42454,N_42105,N_42043);
or U42455 (N_42455,N_42018,N_42022);
and U42456 (N_42456,N_42223,N_42225);
nor U42457 (N_42457,N_42181,N_42095);
or U42458 (N_42458,N_42119,N_42223);
nand U42459 (N_42459,N_42116,N_42110);
nand U42460 (N_42460,N_42177,N_42060);
or U42461 (N_42461,N_42032,N_42084);
nand U42462 (N_42462,N_42244,N_42029);
xnor U42463 (N_42463,N_42216,N_42014);
nand U42464 (N_42464,N_42179,N_42101);
or U42465 (N_42465,N_42227,N_42144);
xnor U42466 (N_42466,N_42203,N_42039);
and U42467 (N_42467,N_42242,N_42097);
nor U42468 (N_42468,N_42092,N_42199);
xor U42469 (N_42469,N_42063,N_42215);
nand U42470 (N_42470,N_42216,N_42011);
nand U42471 (N_42471,N_42173,N_42080);
xor U42472 (N_42472,N_42100,N_42119);
nor U42473 (N_42473,N_42134,N_42080);
and U42474 (N_42474,N_42049,N_42140);
nor U42475 (N_42475,N_42141,N_42000);
nor U42476 (N_42476,N_42026,N_42162);
nor U42477 (N_42477,N_42161,N_42242);
nand U42478 (N_42478,N_42132,N_42079);
nor U42479 (N_42479,N_42123,N_42221);
and U42480 (N_42480,N_42145,N_42052);
nand U42481 (N_42481,N_42180,N_42217);
nand U42482 (N_42482,N_42014,N_42238);
or U42483 (N_42483,N_42246,N_42172);
nor U42484 (N_42484,N_42192,N_42207);
and U42485 (N_42485,N_42088,N_42246);
or U42486 (N_42486,N_42117,N_42061);
xor U42487 (N_42487,N_42196,N_42026);
nor U42488 (N_42488,N_42161,N_42032);
or U42489 (N_42489,N_42227,N_42087);
or U42490 (N_42490,N_42228,N_42180);
nor U42491 (N_42491,N_42104,N_42137);
and U42492 (N_42492,N_42072,N_42024);
nand U42493 (N_42493,N_42182,N_42060);
and U42494 (N_42494,N_42168,N_42109);
nand U42495 (N_42495,N_42155,N_42114);
nor U42496 (N_42496,N_42090,N_42118);
xnor U42497 (N_42497,N_42085,N_42031);
nand U42498 (N_42498,N_42160,N_42001);
nor U42499 (N_42499,N_42118,N_42029);
xnor U42500 (N_42500,N_42477,N_42261);
and U42501 (N_42501,N_42475,N_42376);
or U42502 (N_42502,N_42322,N_42345);
and U42503 (N_42503,N_42339,N_42416);
xor U42504 (N_42504,N_42488,N_42495);
nand U42505 (N_42505,N_42410,N_42404);
nor U42506 (N_42506,N_42499,N_42281);
or U42507 (N_42507,N_42435,N_42434);
or U42508 (N_42508,N_42286,N_42327);
nand U42509 (N_42509,N_42310,N_42275);
and U42510 (N_42510,N_42268,N_42369);
or U42511 (N_42511,N_42332,N_42450);
or U42512 (N_42512,N_42315,N_42363);
or U42513 (N_42513,N_42287,N_42252);
xor U42514 (N_42514,N_42476,N_42259);
xnor U42515 (N_42515,N_42411,N_42457);
nor U42516 (N_42516,N_42378,N_42444);
or U42517 (N_42517,N_42452,N_42373);
xor U42518 (N_42518,N_42437,N_42489);
or U42519 (N_42519,N_42358,N_42302);
nand U42520 (N_42520,N_42494,N_42265);
nand U42521 (N_42521,N_42431,N_42372);
xor U42522 (N_42522,N_42405,N_42263);
and U42523 (N_42523,N_42468,N_42298);
nor U42524 (N_42524,N_42439,N_42390);
nor U42525 (N_42525,N_42326,N_42447);
nor U42526 (N_42526,N_42272,N_42423);
or U42527 (N_42527,N_42309,N_42473);
nor U42528 (N_42528,N_42253,N_42492);
and U42529 (N_42529,N_42328,N_42445);
xnor U42530 (N_42530,N_42269,N_42451);
and U42531 (N_42531,N_42481,N_42442);
and U42532 (N_42532,N_42375,N_42317);
or U42533 (N_42533,N_42251,N_42352);
xor U42534 (N_42534,N_42397,N_42365);
and U42535 (N_42535,N_42391,N_42325);
and U42536 (N_42536,N_42446,N_42455);
xor U42537 (N_42537,N_42316,N_42343);
or U42538 (N_42538,N_42408,N_42306);
or U42539 (N_42539,N_42285,N_42474);
xnor U42540 (N_42540,N_42467,N_42331);
xnor U42541 (N_42541,N_42333,N_42409);
and U42542 (N_42542,N_42480,N_42337);
xnor U42543 (N_42543,N_42303,N_42459);
nand U42544 (N_42544,N_42254,N_42496);
and U42545 (N_42545,N_42355,N_42460);
or U42546 (N_42546,N_42374,N_42371);
or U42547 (N_42547,N_42312,N_42277);
nand U42548 (N_42548,N_42466,N_42276);
xnor U42549 (N_42549,N_42314,N_42340);
nor U42550 (N_42550,N_42418,N_42427);
and U42551 (N_42551,N_42364,N_42382);
nor U42552 (N_42552,N_42484,N_42491);
nor U42553 (N_42553,N_42280,N_42386);
nand U42554 (N_42554,N_42320,N_42432);
nand U42555 (N_42555,N_42498,N_42262);
nand U42556 (N_42556,N_42255,N_42288);
nand U42557 (N_42557,N_42387,N_42299);
xnor U42558 (N_42558,N_42465,N_42295);
nor U42559 (N_42559,N_42300,N_42289);
xor U42560 (N_42560,N_42482,N_42313);
or U42561 (N_42561,N_42438,N_42385);
and U42562 (N_42562,N_42389,N_42301);
xor U42563 (N_42563,N_42440,N_42318);
nor U42564 (N_42564,N_42419,N_42461);
nand U42565 (N_42565,N_42384,N_42353);
nor U42566 (N_42566,N_42443,N_42449);
nor U42567 (N_42567,N_42383,N_42485);
or U42568 (N_42568,N_42270,N_42304);
and U42569 (N_42569,N_42324,N_42470);
nand U42570 (N_42570,N_42296,N_42273);
nor U42571 (N_42571,N_42278,N_42361);
and U42572 (N_42572,N_42456,N_42279);
xor U42573 (N_42573,N_42250,N_42330);
nor U42574 (N_42574,N_42347,N_42417);
nand U42575 (N_42575,N_42258,N_42349);
nor U42576 (N_42576,N_42308,N_42321);
and U42577 (N_42577,N_42424,N_42260);
nor U42578 (N_42578,N_42338,N_42307);
nand U42579 (N_42579,N_42336,N_42421);
xor U42580 (N_42580,N_42380,N_42462);
or U42581 (N_42581,N_42472,N_42478);
xnor U42582 (N_42582,N_42458,N_42311);
and U42583 (N_42583,N_42267,N_42399);
nand U42584 (N_42584,N_42290,N_42305);
and U42585 (N_42585,N_42362,N_42415);
xor U42586 (N_42586,N_42487,N_42256);
nand U42587 (N_42587,N_42403,N_42329);
nand U42588 (N_42588,N_42388,N_42264);
and U42589 (N_42589,N_42342,N_42422);
or U42590 (N_42590,N_42284,N_42335);
nor U42591 (N_42591,N_42293,N_42348);
or U42592 (N_42592,N_42395,N_42291);
nor U42593 (N_42593,N_42257,N_42346);
or U42594 (N_42594,N_42341,N_42282);
and U42595 (N_42595,N_42398,N_42370);
nand U42596 (N_42596,N_42266,N_42493);
nand U42597 (N_42597,N_42360,N_42426);
or U42598 (N_42598,N_42351,N_42486);
xor U42599 (N_42599,N_42441,N_42367);
and U42600 (N_42600,N_42497,N_42429);
or U42601 (N_42601,N_42377,N_42396);
xor U42602 (N_42602,N_42402,N_42464);
and U42603 (N_42603,N_42413,N_42368);
nand U42604 (N_42604,N_42294,N_42356);
nor U42605 (N_42605,N_42469,N_42490);
or U42606 (N_42606,N_42406,N_42425);
nand U42607 (N_42607,N_42344,N_42430);
nand U42608 (N_42608,N_42366,N_42271);
xnor U42609 (N_42609,N_42428,N_42463);
xor U42610 (N_42610,N_42392,N_42414);
and U42611 (N_42611,N_42407,N_42350);
nand U42612 (N_42612,N_42483,N_42453);
xnor U42613 (N_42613,N_42323,N_42479);
and U42614 (N_42614,N_42400,N_42381);
and U42615 (N_42615,N_42283,N_42274);
or U42616 (N_42616,N_42393,N_42354);
nand U42617 (N_42617,N_42454,N_42420);
and U42618 (N_42618,N_42359,N_42292);
xnor U42619 (N_42619,N_42297,N_42319);
nand U42620 (N_42620,N_42334,N_42436);
nor U42621 (N_42621,N_42448,N_42357);
nor U42622 (N_42622,N_42394,N_42471);
nand U42623 (N_42623,N_42433,N_42412);
xnor U42624 (N_42624,N_42379,N_42401);
nor U42625 (N_42625,N_42474,N_42287);
xor U42626 (N_42626,N_42386,N_42376);
or U42627 (N_42627,N_42448,N_42342);
and U42628 (N_42628,N_42396,N_42389);
nor U42629 (N_42629,N_42426,N_42432);
or U42630 (N_42630,N_42467,N_42454);
or U42631 (N_42631,N_42267,N_42407);
or U42632 (N_42632,N_42334,N_42372);
or U42633 (N_42633,N_42291,N_42471);
and U42634 (N_42634,N_42434,N_42479);
nand U42635 (N_42635,N_42470,N_42398);
or U42636 (N_42636,N_42417,N_42488);
nor U42637 (N_42637,N_42471,N_42434);
and U42638 (N_42638,N_42265,N_42296);
or U42639 (N_42639,N_42405,N_42311);
xor U42640 (N_42640,N_42429,N_42435);
or U42641 (N_42641,N_42322,N_42253);
nor U42642 (N_42642,N_42281,N_42430);
nand U42643 (N_42643,N_42258,N_42375);
and U42644 (N_42644,N_42389,N_42417);
xor U42645 (N_42645,N_42370,N_42389);
xnor U42646 (N_42646,N_42440,N_42314);
xor U42647 (N_42647,N_42442,N_42499);
xor U42648 (N_42648,N_42492,N_42266);
nor U42649 (N_42649,N_42498,N_42358);
and U42650 (N_42650,N_42437,N_42417);
nor U42651 (N_42651,N_42483,N_42427);
and U42652 (N_42652,N_42336,N_42313);
xor U42653 (N_42653,N_42293,N_42499);
nor U42654 (N_42654,N_42394,N_42355);
nand U42655 (N_42655,N_42477,N_42497);
nand U42656 (N_42656,N_42290,N_42315);
nor U42657 (N_42657,N_42380,N_42258);
nor U42658 (N_42658,N_42403,N_42414);
nor U42659 (N_42659,N_42309,N_42305);
nor U42660 (N_42660,N_42273,N_42271);
or U42661 (N_42661,N_42302,N_42333);
and U42662 (N_42662,N_42436,N_42469);
and U42663 (N_42663,N_42369,N_42469);
xnor U42664 (N_42664,N_42479,N_42381);
nor U42665 (N_42665,N_42318,N_42331);
xor U42666 (N_42666,N_42492,N_42256);
xor U42667 (N_42667,N_42473,N_42467);
and U42668 (N_42668,N_42429,N_42380);
nor U42669 (N_42669,N_42407,N_42459);
xnor U42670 (N_42670,N_42454,N_42275);
and U42671 (N_42671,N_42273,N_42328);
xor U42672 (N_42672,N_42446,N_42444);
and U42673 (N_42673,N_42495,N_42267);
and U42674 (N_42674,N_42448,N_42296);
nand U42675 (N_42675,N_42473,N_42499);
nor U42676 (N_42676,N_42373,N_42272);
xor U42677 (N_42677,N_42298,N_42446);
or U42678 (N_42678,N_42281,N_42444);
xnor U42679 (N_42679,N_42408,N_42331);
nand U42680 (N_42680,N_42268,N_42285);
nor U42681 (N_42681,N_42362,N_42421);
xor U42682 (N_42682,N_42278,N_42403);
nand U42683 (N_42683,N_42330,N_42264);
and U42684 (N_42684,N_42459,N_42299);
xnor U42685 (N_42685,N_42406,N_42478);
and U42686 (N_42686,N_42484,N_42369);
xnor U42687 (N_42687,N_42442,N_42378);
or U42688 (N_42688,N_42339,N_42371);
or U42689 (N_42689,N_42499,N_42398);
nor U42690 (N_42690,N_42454,N_42433);
and U42691 (N_42691,N_42298,N_42253);
nor U42692 (N_42692,N_42271,N_42445);
nand U42693 (N_42693,N_42342,N_42392);
nand U42694 (N_42694,N_42262,N_42386);
or U42695 (N_42695,N_42340,N_42278);
nand U42696 (N_42696,N_42460,N_42406);
or U42697 (N_42697,N_42460,N_42428);
nand U42698 (N_42698,N_42356,N_42434);
or U42699 (N_42699,N_42348,N_42311);
or U42700 (N_42700,N_42367,N_42375);
and U42701 (N_42701,N_42410,N_42354);
or U42702 (N_42702,N_42272,N_42493);
or U42703 (N_42703,N_42391,N_42420);
nor U42704 (N_42704,N_42466,N_42322);
nand U42705 (N_42705,N_42274,N_42278);
nand U42706 (N_42706,N_42437,N_42267);
and U42707 (N_42707,N_42414,N_42343);
and U42708 (N_42708,N_42267,N_42381);
xnor U42709 (N_42709,N_42362,N_42268);
or U42710 (N_42710,N_42339,N_42255);
and U42711 (N_42711,N_42357,N_42420);
nand U42712 (N_42712,N_42436,N_42472);
and U42713 (N_42713,N_42459,N_42293);
nand U42714 (N_42714,N_42404,N_42331);
xnor U42715 (N_42715,N_42278,N_42352);
xor U42716 (N_42716,N_42395,N_42311);
or U42717 (N_42717,N_42315,N_42340);
or U42718 (N_42718,N_42380,N_42260);
nand U42719 (N_42719,N_42432,N_42491);
nand U42720 (N_42720,N_42499,N_42448);
nor U42721 (N_42721,N_42498,N_42328);
and U42722 (N_42722,N_42495,N_42434);
xor U42723 (N_42723,N_42494,N_42260);
xnor U42724 (N_42724,N_42369,N_42401);
nor U42725 (N_42725,N_42262,N_42490);
nand U42726 (N_42726,N_42265,N_42305);
or U42727 (N_42727,N_42288,N_42405);
or U42728 (N_42728,N_42411,N_42425);
nor U42729 (N_42729,N_42460,N_42354);
xor U42730 (N_42730,N_42492,N_42497);
xnor U42731 (N_42731,N_42341,N_42307);
nand U42732 (N_42732,N_42261,N_42453);
and U42733 (N_42733,N_42283,N_42492);
nor U42734 (N_42734,N_42371,N_42421);
xnor U42735 (N_42735,N_42283,N_42490);
and U42736 (N_42736,N_42487,N_42326);
or U42737 (N_42737,N_42327,N_42287);
xnor U42738 (N_42738,N_42496,N_42334);
or U42739 (N_42739,N_42353,N_42327);
and U42740 (N_42740,N_42439,N_42415);
and U42741 (N_42741,N_42252,N_42392);
nand U42742 (N_42742,N_42396,N_42380);
xor U42743 (N_42743,N_42324,N_42410);
nor U42744 (N_42744,N_42279,N_42344);
and U42745 (N_42745,N_42371,N_42493);
nor U42746 (N_42746,N_42350,N_42455);
nor U42747 (N_42747,N_42362,N_42436);
and U42748 (N_42748,N_42253,N_42362);
nor U42749 (N_42749,N_42391,N_42274);
nor U42750 (N_42750,N_42683,N_42515);
and U42751 (N_42751,N_42651,N_42614);
xnor U42752 (N_42752,N_42578,N_42732);
nor U42753 (N_42753,N_42593,N_42510);
nand U42754 (N_42754,N_42659,N_42692);
nor U42755 (N_42755,N_42574,N_42560);
xor U42756 (N_42756,N_42680,N_42537);
nor U42757 (N_42757,N_42577,N_42517);
and U42758 (N_42758,N_42655,N_42598);
or U42759 (N_42759,N_42671,N_42632);
or U42760 (N_42760,N_42658,N_42738);
xnor U42761 (N_42761,N_42588,N_42693);
xor U42762 (N_42762,N_42511,N_42661);
and U42763 (N_42763,N_42597,N_42523);
nand U42764 (N_42764,N_42535,N_42694);
nand U42765 (N_42765,N_42739,N_42566);
nor U42766 (N_42766,N_42709,N_42534);
nor U42767 (N_42767,N_42706,N_42715);
nand U42768 (N_42768,N_42635,N_42616);
nor U42769 (N_42769,N_42507,N_42691);
and U42770 (N_42770,N_42639,N_42696);
and U42771 (N_42771,N_42613,N_42708);
nor U42772 (N_42772,N_42713,N_42521);
xor U42773 (N_42773,N_42512,N_42663);
xor U42774 (N_42774,N_42500,N_42531);
and U42775 (N_42775,N_42522,N_42625);
nand U42776 (N_42776,N_42684,N_42650);
xor U42777 (N_42777,N_42688,N_42711);
or U42778 (N_42778,N_42594,N_42723);
and U42779 (N_42779,N_42573,N_42689);
nand U42780 (N_42780,N_42528,N_42662);
nand U42781 (N_42781,N_42538,N_42619);
nand U42782 (N_42782,N_42552,N_42668);
nand U42783 (N_42783,N_42519,N_42508);
and U42784 (N_42784,N_42627,N_42716);
and U42785 (N_42785,N_42637,N_42717);
nor U42786 (N_42786,N_42645,N_42612);
nor U42787 (N_42787,N_42638,N_42643);
nand U42788 (N_42788,N_42745,N_42687);
nand U42789 (N_42789,N_42599,N_42622);
or U42790 (N_42790,N_42742,N_42749);
and U42791 (N_42791,N_42553,N_42626);
xor U42792 (N_42792,N_42660,N_42697);
nor U42793 (N_42793,N_42664,N_42605);
nand U42794 (N_42794,N_42722,N_42609);
and U42795 (N_42795,N_42737,N_42724);
and U42796 (N_42796,N_42561,N_42648);
xnor U42797 (N_42797,N_42590,N_42569);
or U42798 (N_42798,N_42563,N_42685);
nand U42799 (N_42799,N_42721,N_42733);
nand U42800 (N_42800,N_42505,N_42631);
and U42801 (N_42801,N_42618,N_42589);
nor U42802 (N_42802,N_42610,N_42529);
nand U42803 (N_42803,N_42666,N_42550);
or U42804 (N_42804,N_42501,N_42656);
xor U42805 (N_42805,N_42514,N_42678);
and U42806 (N_42806,N_42516,N_42608);
xnor U42807 (N_42807,N_42699,N_42587);
xor U42808 (N_42808,N_42543,N_42703);
or U42809 (N_42809,N_42576,N_42642);
and U42810 (N_42810,N_42503,N_42532);
or U42811 (N_42811,N_42546,N_42581);
and U42812 (N_42812,N_42542,N_42628);
nor U42813 (N_42813,N_42630,N_42747);
xnor U42814 (N_42814,N_42714,N_42585);
nand U42815 (N_42815,N_42541,N_42653);
or U42816 (N_42816,N_42556,N_42539);
xor U42817 (N_42817,N_42729,N_42735);
and U42818 (N_42818,N_42572,N_42743);
and U42819 (N_42819,N_42670,N_42741);
xor U42820 (N_42820,N_42611,N_42702);
xor U42821 (N_42821,N_42682,N_42633);
nand U42822 (N_42822,N_42586,N_42710);
xnor U42823 (N_42823,N_42654,N_42575);
xor U42824 (N_42824,N_42652,N_42551);
nand U42825 (N_42825,N_42718,N_42509);
and U42826 (N_42826,N_42557,N_42647);
and U42827 (N_42827,N_42533,N_42690);
and U42828 (N_42828,N_42502,N_42530);
nand U42829 (N_42829,N_42559,N_42667);
nor U42830 (N_42830,N_42669,N_42624);
nand U42831 (N_42831,N_42524,N_42513);
or U42832 (N_42832,N_42571,N_42634);
and U42833 (N_42833,N_42602,N_42606);
xor U42834 (N_42834,N_42579,N_42704);
or U42835 (N_42835,N_42504,N_42580);
nand U42836 (N_42836,N_42621,N_42665);
or U42837 (N_42837,N_42701,N_42712);
nor U42838 (N_42838,N_42746,N_42707);
or U42839 (N_42839,N_42558,N_42615);
and U42840 (N_42840,N_42565,N_42679);
nand U42841 (N_42841,N_42596,N_42641);
xnor U42842 (N_42842,N_42549,N_42730);
nor U42843 (N_42843,N_42603,N_42744);
or U42844 (N_42844,N_42601,N_42698);
nor U42845 (N_42845,N_42520,N_42544);
or U42846 (N_42846,N_42736,N_42740);
xor U42847 (N_42847,N_42540,N_42695);
and U42848 (N_42848,N_42526,N_42554);
nor U42849 (N_42849,N_42725,N_42681);
or U42850 (N_42850,N_42592,N_42617);
nor U42851 (N_42851,N_42726,N_42582);
and U42852 (N_42852,N_42527,N_42555);
nor U42853 (N_42853,N_42640,N_42727);
xnor U42854 (N_42854,N_42623,N_42570);
nor U42855 (N_42855,N_42677,N_42731);
or U42856 (N_42856,N_42674,N_42584);
xor U42857 (N_42857,N_42536,N_42562);
or U42858 (N_42858,N_42506,N_42646);
and U42859 (N_42859,N_42604,N_42547);
or U42860 (N_42860,N_42568,N_42686);
xnor U42861 (N_42861,N_42705,N_42545);
or U42862 (N_42862,N_42675,N_42607);
nand U42863 (N_42863,N_42676,N_42564);
nand U42864 (N_42864,N_42644,N_42595);
xnor U42865 (N_42865,N_42720,N_42620);
nor U42866 (N_42866,N_42657,N_42728);
and U42867 (N_42867,N_42525,N_42600);
xor U42868 (N_42868,N_42672,N_42583);
or U42869 (N_42869,N_42673,N_42636);
nor U42870 (N_42870,N_42629,N_42518);
nor U42871 (N_42871,N_42649,N_42591);
and U42872 (N_42872,N_42567,N_42719);
xnor U42873 (N_42873,N_42700,N_42734);
xnor U42874 (N_42874,N_42548,N_42748);
nor U42875 (N_42875,N_42656,N_42704);
and U42876 (N_42876,N_42739,N_42660);
nand U42877 (N_42877,N_42627,N_42739);
or U42878 (N_42878,N_42569,N_42656);
and U42879 (N_42879,N_42650,N_42717);
and U42880 (N_42880,N_42602,N_42669);
and U42881 (N_42881,N_42527,N_42711);
or U42882 (N_42882,N_42694,N_42744);
and U42883 (N_42883,N_42738,N_42707);
and U42884 (N_42884,N_42637,N_42679);
nor U42885 (N_42885,N_42640,N_42591);
or U42886 (N_42886,N_42550,N_42587);
xnor U42887 (N_42887,N_42605,N_42519);
nand U42888 (N_42888,N_42608,N_42578);
or U42889 (N_42889,N_42624,N_42543);
nor U42890 (N_42890,N_42671,N_42732);
or U42891 (N_42891,N_42602,N_42640);
nor U42892 (N_42892,N_42674,N_42630);
and U42893 (N_42893,N_42593,N_42577);
and U42894 (N_42894,N_42583,N_42500);
xnor U42895 (N_42895,N_42697,N_42679);
xnor U42896 (N_42896,N_42582,N_42679);
and U42897 (N_42897,N_42714,N_42582);
xor U42898 (N_42898,N_42735,N_42518);
xnor U42899 (N_42899,N_42656,N_42696);
nor U42900 (N_42900,N_42723,N_42593);
and U42901 (N_42901,N_42682,N_42683);
nand U42902 (N_42902,N_42522,N_42660);
nand U42903 (N_42903,N_42637,N_42607);
xnor U42904 (N_42904,N_42581,N_42575);
nor U42905 (N_42905,N_42702,N_42538);
or U42906 (N_42906,N_42623,N_42661);
or U42907 (N_42907,N_42653,N_42669);
nand U42908 (N_42908,N_42695,N_42521);
nand U42909 (N_42909,N_42516,N_42668);
nor U42910 (N_42910,N_42684,N_42592);
nand U42911 (N_42911,N_42695,N_42642);
and U42912 (N_42912,N_42729,N_42669);
nand U42913 (N_42913,N_42617,N_42570);
or U42914 (N_42914,N_42628,N_42714);
nor U42915 (N_42915,N_42543,N_42680);
xnor U42916 (N_42916,N_42674,N_42742);
nor U42917 (N_42917,N_42682,N_42601);
nor U42918 (N_42918,N_42596,N_42652);
nor U42919 (N_42919,N_42713,N_42710);
nor U42920 (N_42920,N_42570,N_42593);
nor U42921 (N_42921,N_42655,N_42714);
nand U42922 (N_42922,N_42532,N_42560);
nor U42923 (N_42923,N_42688,N_42680);
xnor U42924 (N_42924,N_42557,N_42665);
xor U42925 (N_42925,N_42654,N_42632);
nand U42926 (N_42926,N_42518,N_42610);
or U42927 (N_42927,N_42501,N_42502);
or U42928 (N_42928,N_42676,N_42710);
and U42929 (N_42929,N_42646,N_42607);
nor U42930 (N_42930,N_42683,N_42615);
nor U42931 (N_42931,N_42510,N_42532);
or U42932 (N_42932,N_42509,N_42678);
nand U42933 (N_42933,N_42686,N_42531);
nand U42934 (N_42934,N_42531,N_42566);
nor U42935 (N_42935,N_42619,N_42620);
nand U42936 (N_42936,N_42737,N_42742);
xor U42937 (N_42937,N_42569,N_42665);
or U42938 (N_42938,N_42702,N_42677);
or U42939 (N_42939,N_42679,N_42570);
or U42940 (N_42940,N_42724,N_42738);
nand U42941 (N_42941,N_42525,N_42682);
and U42942 (N_42942,N_42570,N_42521);
nor U42943 (N_42943,N_42611,N_42675);
or U42944 (N_42944,N_42535,N_42591);
nand U42945 (N_42945,N_42511,N_42650);
xor U42946 (N_42946,N_42535,N_42646);
or U42947 (N_42947,N_42586,N_42665);
and U42948 (N_42948,N_42747,N_42657);
nor U42949 (N_42949,N_42617,N_42735);
nor U42950 (N_42950,N_42511,N_42731);
nand U42951 (N_42951,N_42609,N_42710);
or U42952 (N_42952,N_42514,N_42698);
xor U42953 (N_42953,N_42747,N_42522);
nor U42954 (N_42954,N_42566,N_42700);
xor U42955 (N_42955,N_42581,N_42541);
and U42956 (N_42956,N_42691,N_42636);
xnor U42957 (N_42957,N_42655,N_42575);
or U42958 (N_42958,N_42661,N_42749);
xor U42959 (N_42959,N_42537,N_42722);
nand U42960 (N_42960,N_42726,N_42657);
nand U42961 (N_42961,N_42637,N_42697);
nand U42962 (N_42962,N_42731,N_42620);
or U42963 (N_42963,N_42515,N_42692);
xor U42964 (N_42964,N_42560,N_42584);
xnor U42965 (N_42965,N_42699,N_42664);
or U42966 (N_42966,N_42723,N_42744);
nor U42967 (N_42967,N_42639,N_42553);
and U42968 (N_42968,N_42525,N_42720);
nand U42969 (N_42969,N_42660,N_42519);
xor U42970 (N_42970,N_42546,N_42544);
xnor U42971 (N_42971,N_42638,N_42546);
or U42972 (N_42972,N_42545,N_42726);
xor U42973 (N_42973,N_42680,N_42670);
and U42974 (N_42974,N_42516,N_42745);
nor U42975 (N_42975,N_42740,N_42651);
xnor U42976 (N_42976,N_42695,N_42683);
nor U42977 (N_42977,N_42612,N_42748);
or U42978 (N_42978,N_42511,N_42563);
nor U42979 (N_42979,N_42591,N_42646);
nor U42980 (N_42980,N_42609,N_42608);
or U42981 (N_42981,N_42581,N_42665);
nor U42982 (N_42982,N_42749,N_42543);
nand U42983 (N_42983,N_42688,N_42673);
or U42984 (N_42984,N_42560,N_42523);
nor U42985 (N_42985,N_42653,N_42558);
or U42986 (N_42986,N_42507,N_42725);
and U42987 (N_42987,N_42605,N_42735);
xnor U42988 (N_42988,N_42605,N_42523);
nor U42989 (N_42989,N_42729,N_42565);
or U42990 (N_42990,N_42609,N_42701);
or U42991 (N_42991,N_42568,N_42507);
xnor U42992 (N_42992,N_42638,N_42606);
or U42993 (N_42993,N_42652,N_42734);
xnor U42994 (N_42994,N_42571,N_42501);
nor U42995 (N_42995,N_42589,N_42552);
or U42996 (N_42996,N_42653,N_42564);
or U42997 (N_42997,N_42553,N_42688);
or U42998 (N_42998,N_42667,N_42725);
or U42999 (N_42999,N_42619,N_42722);
or U43000 (N_43000,N_42989,N_42792);
or U43001 (N_43001,N_42966,N_42871);
nor U43002 (N_43002,N_42914,N_42875);
and U43003 (N_43003,N_42827,N_42802);
or U43004 (N_43004,N_42976,N_42838);
and U43005 (N_43005,N_42945,N_42795);
and U43006 (N_43006,N_42804,N_42988);
xnor U43007 (N_43007,N_42953,N_42915);
and U43008 (N_43008,N_42927,N_42797);
or U43009 (N_43009,N_42779,N_42984);
nand U43010 (N_43010,N_42985,N_42995);
or U43011 (N_43011,N_42811,N_42766);
nand U43012 (N_43012,N_42829,N_42867);
and U43013 (N_43013,N_42775,N_42866);
nand U43014 (N_43014,N_42922,N_42819);
nor U43015 (N_43015,N_42760,N_42852);
or U43016 (N_43016,N_42847,N_42986);
xnor U43017 (N_43017,N_42774,N_42937);
xnor U43018 (N_43018,N_42853,N_42783);
or U43019 (N_43019,N_42841,N_42877);
and U43020 (N_43020,N_42850,N_42778);
nor U43021 (N_43021,N_42998,N_42761);
and U43022 (N_43022,N_42786,N_42785);
or U43023 (N_43023,N_42815,N_42952);
and U43024 (N_43024,N_42809,N_42794);
and U43025 (N_43025,N_42924,N_42753);
and U43026 (N_43026,N_42928,N_42870);
and U43027 (N_43027,N_42773,N_42782);
and U43028 (N_43028,N_42756,N_42895);
and U43029 (N_43029,N_42769,N_42874);
nand U43030 (N_43030,N_42892,N_42939);
and U43031 (N_43031,N_42757,N_42816);
nor U43032 (N_43032,N_42938,N_42970);
xor U43033 (N_43033,N_42996,N_42948);
or U43034 (N_43034,N_42803,N_42967);
xnor U43035 (N_43035,N_42767,N_42911);
or U43036 (N_43036,N_42902,N_42878);
nor U43037 (N_43037,N_42865,N_42856);
or U43038 (N_43038,N_42910,N_42840);
nand U43039 (N_43039,N_42750,N_42981);
or U43040 (N_43040,N_42858,N_42861);
nor U43041 (N_43041,N_42823,N_42896);
nor U43042 (N_43042,N_42955,N_42889);
and U43043 (N_43043,N_42980,N_42975);
xor U43044 (N_43044,N_42810,N_42935);
or U43045 (N_43045,N_42831,N_42974);
nand U43046 (N_43046,N_42936,N_42876);
or U43047 (N_43047,N_42789,N_42772);
and U43048 (N_43048,N_42834,N_42848);
nand U43049 (N_43049,N_42891,N_42825);
nor U43050 (N_43050,N_42954,N_42755);
nand U43051 (N_43051,N_42971,N_42946);
xnor U43052 (N_43052,N_42805,N_42963);
and U43053 (N_43053,N_42784,N_42821);
and U43054 (N_43054,N_42758,N_42898);
xnor U43055 (N_43055,N_42934,N_42776);
and U43056 (N_43056,N_42991,N_42839);
nand U43057 (N_43057,N_42893,N_42899);
nor U43058 (N_43058,N_42987,N_42880);
nand U43059 (N_43059,N_42968,N_42930);
or U43060 (N_43060,N_42947,N_42798);
and U43061 (N_43061,N_42793,N_42799);
and U43062 (N_43062,N_42957,N_42860);
nor U43063 (N_43063,N_42796,N_42851);
nand U43064 (N_43064,N_42762,N_42908);
nor U43065 (N_43065,N_42864,N_42906);
nand U43066 (N_43066,N_42973,N_42763);
nor U43067 (N_43067,N_42904,N_42873);
xnor U43068 (N_43068,N_42997,N_42917);
xor U43069 (N_43069,N_42859,N_42923);
xor U43070 (N_43070,N_42836,N_42846);
nand U43071 (N_43071,N_42913,N_42887);
nand U43072 (N_43072,N_42949,N_42909);
and U43073 (N_43073,N_42978,N_42820);
or U43074 (N_43074,N_42872,N_42842);
nand U43075 (N_43075,N_42905,N_42884);
nand U43076 (N_43076,N_42977,N_42857);
or U43077 (N_43077,N_42907,N_42770);
xor U43078 (N_43078,N_42894,N_42943);
and U43079 (N_43079,N_42929,N_42926);
and U43080 (N_43080,N_42951,N_42863);
or U43081 (N_43081,N_42969,N_42849);
nor U43082 (N_43082,N_42854,N_42900);
nand U43083 (N_43083,N_42868,N_42788);
or U43084 (N_43084,N_42837,N_42808);
nand U43085 (N_43085,N_42807,N_42814);
or U43086 (N_43086,N_42932,N_42835);
and U43087 (N_43087,N_42781,N_42982);
nor U43088 (N_43088,N_42990,N_42959);
xnor U43089 (N_43089,N_42890,N_42994);
nor U43090 (N_43090,N_42919,N_42777);
and U43091 (N_43091,N_42818,N_42933);
xnor U43092 (N_43092,N_42941,N_42883);
xor U43093 (N_43093,N_42964,N_42921);
nand U43094 (N_43094,N_42958,N_42791);
or U43095 (N_43095,N_42888,N_42833);
and U43096 (N_43096,N_42845,N_42824);
xnor U43097 (N_43097,N_42806,N_42886);
and U43098 (N_43098,N_42993,N_42965);
nor U43099 (N_43099,N_42879,N_42813);
and U43100 (N_43100,N_42790,N_42830);
and U43101 (N_43101,N_42751,N_42801);
nand U43102 (N_43102,N_42983,N_42828);
nand U43103 (N_43103,N_42844,N_42916);
and U43104 (N_43104,N_42903,N_42925);
nor U43105 (N_43105,N_42956,N_42885);
xnor U43106 (N_43106,N_42787,N_42862);
and U43107 (N_43107,N_42881,N_42780);
nand U43108 (N_43108,N_42817,N_42812);
or U43109 (N_43109,N_42754,N_42999);
nand U43110 (N_43110,N_42765,N_42768);
or U43111 (N_43111,N_42992,N_42882);
nor U43112 (N_43112,N_42759,N_42944);
nor U43113 (N_43113,N_42961,N_42920);
nor U43114 (N_43114,N_42979,N_42940);
nor U43115 (N_43115,N_42897,N_42960);
xnor U43116 (N_43116,N_42950,N_42962);
or U43117 (N_43117,N_42912,N_42972);
nor U43118 (N_43118,N_42752,N_42822);
nor U43119 (N_43119,N_42771,N_42843);
xnor U43120 (N_43120,N_42832,N_42942);
nor U43121 (N_43121,N_42855,N_42901);
xnor U43122 (N_43122,N_42869,N_42800);
or U43123 (N_43123,N_42826,N_42918);
nor U43124 (N_43124,N_42764,N_42931);
nor U43125 (N_43125,N_42822,N_42948);
or U43126 (N_43126,N_42830,N_42872);
nand U43127 (N_43127,N_42918,N_42950);
or U43128 (N_43128,N_42769,N_42930);
nand U43129 (N_43129,N_42957,N_42824);
or U43130 (N_43130,N_42818,N_42856);
nor U43131 (N_43131,N_42881,N_42988);
nor U43132 (N_43132,N_42847,N_42860);
nand U43133 (N_43133,N_42948,N_42816);
nand U43134 (N_43134,N_42839,N_42890);
xor U43135 (N_43135,N_42967,N_42859);
xnor U43136 (N_43136,N_42913,N_42989);
or U43137 (N_43137,N_42836,N_42810);
xnor U43138 (N_43138,N_42862,N_42868);
nand U43139 (N_43139,N_42764,N_42773);
nand U43140 (N_43140,N_42913,N_42896);
nand U43141 (N_43141,N_42780,N_42951);
xnor U43142 (N_43142,N_42802,N_42839);
and U43143 (N_43143,N_42805,N_42775);
nor U43144 (N_43144,N_42925,N_42911);
or U43145 (N_43145,N_42753,N_42844);
xnor U43146 (N_43146,N_42763,N_42872);
and U43147 (N_43147,N_42896,N_42779);
or U43148 (N_43148,N_42898,N_42964);
nand U43149 (N_43149,N_42759,N_42773);
nand U43150 (N_43150,N_42974,N_42933);
or U43151 (N_43151,N_42904,N_42981);
and U43152 (N_43152,N_42761,N_42828);
and U43153 (N_43153,N_42816,N_42864);
xor U43154 (N_43154,N_42941,N_42884);
xnor U43155 (N_43155,N_42778,N_42974);
or U43156 (N_43156,N_42834,N_42890);
nand U43157 (N_43157,N_42945,N_42866);
and U43158 (N_43158,N_42864,N_42775);
xnor U43159 (N_43159,N_42842,N_42856);
or U43160 (N_43160,N_42870,N_42927);
nor U43161 (N_43161,N_42806,N_42807);
and U43162 (N_43162,N_42761,N_42923);
nor U43163 (N_43163,N_42851,N_42928);
nor U43164 (N_43164,N_42900,N_42998);
nor U43165 (N_43165,N_42775,N_42761);
nand U43166 (N_43166,N_42933,N_42839);
or U43167 (N_43167,N_42808,N_42774);
nand U43168 (N_43168,N_42957,N_42775);
or U43169 (N_43169,N_42973,N_42839);
or U43170 (N_43170,N_42764,N_42922);
xor U43171 (N_43171,N_42939,N_42767);
xnor U43172 (N_43172,N_42801,N_42821);
and U43173 (N_43173,N_42808,N_42873);
nor U43174 (N_43174,N_42815,N_42980);
nor U43175 (N_43175,N_42899,N_42775);
and U43176 (N_43176,N_42848,N_42828);
nand U43177 (N_43177,N_42928,N_42804);
or U43178 (N_43178,N_42909,N_42760);
or U43179 (N_43179,N_42977,N_42818);
xnor U43180 (N_43180,N_42866,N_42765);
and U43181 (N_43181,N_42821,N_42805);
or U43182 (N_43182,N_42847,N_42835);
or U43183 (N_43183,N_42873,N_42943);
or U43184 (N_43184,N_42939,N_42751);
xor U43185 (N_43185,N_42866,N_42836);
or U43186 (N_43186,N_42932,N_42802);
xnor U43187 (N_43187,N_42975,N_42943);
xor U43188 (N_43188,N_42879,N_42876);
or U43189 (N_43189,N_42764,N_42787);
and U43190 (N_43190,N_42951,N_42953);
xnor U43191 (N_43191,N_42889,N_42900);
nand U43192 (N_43192,N_42911,N_42766);
nor U43193 (N_43193,N_42923,N_42967);
or U43194 (N_43194,N_42849,N_42787);
nor U43195 (N_43195,N_42877,N_42928);
xnor U43196 (N_43196,N_42751,N_42869);
and U43197 (N_43197,N_42888,N_42775);
nor U43198 (N_43198,N_42800,N_42940);
xnor U43199 (N_43199,N_42987,N_42767);
nand U43200 (N_43200,N_42838,N_42796);
and U43201 (N_43201,N_42778,N_42814);
and U43202 (N_43202,N_42914,N_42802);
nor U43203 (N_43203,N_42857,N_42753);
nand U43204 (N_43204,N_42918,N_42945);
and U43205 (N_43205,N_42993,N_42868);
xnor U43206 (N_43206,N_42883,N_42782);
xnor U43207 (N_43207,N_42886,N_42989);
or U43208 (N_43208,N_42812,N_42892);
nand U43209 (N_43209,N_42777,N_42890);
or U43210 (N_43210,N_42976,N_42881);
nand U43211 (N_43211,N_42932,N_42956);
nand U43212 (N_43212,N_42757,N_42766);
nor U43213 (N_43213,N_42770,N_42823);
xnor U43214 (N_43214,N_42920,N_42890);
nor U43215 (N_43215,N_42809,N_42945);
or U43216 (N_43216,N_42799,N_42958);
or U43217 (N_43217,N_42750,N_42994);
and U43218 (N_43218,N_42858,N_42805);
and U43219 (N_43219,N_42946,N_42981);
xnor U43220 (N_43220,N_42817,N_42932);
and U43221 (N_43221,N_42816,N_42886);
xnor U43222 (N_43222,N_42877,N_42975);
or U43223 (N_43223,N_42958,N_42959);
or U43224 (N_43224,N_42954,N_42813);
nor U43225 (N_43225,N_42840,N_42826);
nor U43226 (N_43226,N_42960,N_42989);
and U43227 (N_43227,N_42776,N_42951);
xnor U43228 (N_43228,N_42834,N_42766);
and U43229 (N_43229,N_42841,N_42970);
or U43230 (N_43230,N_42820,N_42765);
xnor U43231 (N_43231,N_42933,N_42804);
nand U43232 (N_43232,N_42843,N_42972);
nor U43233 (N_43233,N_42995,N_42931);
or U43234 (N_43234,N_42911,N_42857);
nand U43235 (N_43235,N_42786,N_42750);
nand U43236 (N_43236,N_42877,N_42991);
xor U43237 (N_43237,N_42809,N_42771);
or U43238 (N_43238,N_42913,N_42948);
nor U43239 (N_43239,N_42859,N_42820);
nor U43240 (N_43240,N_42980,N_42832);
nand U43241 (N_43241,N_42946,N_42918);
nor U43242 (N_43242,N_42770,N_42920);
xor U43243 (N_43243,N_42935,N_42874);
xor U43244 (N_43244,N_42867,N_42805);
xnor U43245 (N_43245,N_42813,N_42851);
or U43246 (N_43246,N_42751,N_42980);
and U43247 (N_43247,N_42872,N_42890);
nor U43248 (N_43248,N_42885,N_42876);
or U43249 (N_43249,N_42998,N_42770);
nor U43250 (N_43250,N_43213,N_43113);
or U43251 (N_43251,N_43189,N_43088);
nand U43252 (N_43252,N_43159,N_43244);
nand U43253 (N_43253,N_43199,N_43000);
nor U43254 (N_43254,N_43120,N_43231);
or U43255 (N_43255,N_43025,N_43106);
nand U43256 (N_43256,N_43237,N_43082);
or U43257 (N_43257,N_43238,N_43191);
or U43258 (N_43258,N_43022,N_43172);
and U43259 (N_43259,N_43154,N_43174);
nor U43260 (N_43260,N_43206,N_43036);
or U43261 (N_43261,N_43029,N_43086);
xor U43262 (N_43262,N_43186,N_43239);
nor U43263 (N_43263,N_43085,N_43046);
nand U43264 (N_43264,N_43019,N_43247);
nor U43265 (N_43265,N_43081,N_43127);
nand U43266 (N_43266,N_43075,N_43087);
xnor U43267 (N_43267,N_43230,N_43011);
or U43268 (N_43268,N_43183,N_43077);
nand U43269 (N_43269,N_43134,N_43116);
or U43270 (N_43270,N_43150,N_43180);
nor U43271 (N_43271,N_43068,N_43208);
nor U43272 (N_43272,N_43061,N_43100);
nor U43273 (N_43273,N_43161,N_43115);
nand U43274 (N_43274,N_43016,N_43094);
nand U43275 (N_43275,N_43035,N_43048);
and U43276 (N_43276,N_43060,N_43198);
xnor U43277 (N_43277,N_43090,N_43064);
nand U43278 (N_43278,N_43181,N_43063);
nor U43279 (N_43279,N_43062,N_43190);
and U43280 (N_43280,N_43249,N_43155);
or U43281 (N_43281,N_43021,N_43076);
nor U43282 (N_43282,N_43053,N_43059);
nor U43283 (N_43283,N_43223,N_43142);
and U43284 (N_43284,N_43004,N_43099);
or U43285 (N_43285,N_43092,N_43138);
and U43286 (N_43286,N_43222,N_43158);
or U43287 (N_43287,N_43111,N_43041);
xor U43288 (N_43288,N_43013,N_43096);
xor U43289 (N_43289,N_43006,N_43105);
nand U43290 (N_43290,N_43139,N_43031);
nor U43291 (N_43291,N_43132,N_43078);
or U43292 (N_43292,N_43066,N_43215);
nor U43293 (N_43293,N_43095,N_43165);
or U43294 (N_43294,N_43187,N_43185);
nor U43295 (N_43295,N_43101,N_43028);
and U43296 (N_43296,N_43196,N_43147);
or U43297 (N_43297,N_43212,N_43024);
xor U43298 (N_43298,N_43093,N_43234);
and U43299 (N_43299,N_43129,N_43097);
nor U43300 (N_43300,N_43005,N_43117);
nand U43301 (N_43301,N_43176,N_43017);
or U43302 (N_43302,N_43131,N_43056);
and U43303 (N_43303,N_43151,N_43124);
and U43304 (N_43304,N_43235,N_43098);
nor U43305 (N_43305,N_43052,N_43042);
and U43306 (N_43306,N_43050,N_43074);
nand U43307 (N_43307,N_43130,N_43055);
and U43308 (N_43308,N_43207,N_43047);
nor U43309 (N_43309,N_43119,N_43170);
xnor U43310 (N_43310,N_43108,N_43102);
nor U43311 (N_43311,N_43168,N_43089);
nor U43312 (N_43312,N_43232,N_43173);
and U43313 (N_43313,N_43084,N_43146);
nand U43314 (N_43314,N_43080,N_43014);
nor U43315 (N_43315,N_43192,N_43141);
and U43316 (N_43316,N_43003,N_43103);
xor U43317 (N_43317,N_43203,N_43169);
nand U43318 (N_43318,N_43209,N_43073);
nor U43319 (N_43319,N_43160,N_43104);
and U43320 (N_43320,N_43164,N_43023);
and U43321 (N_43321,N_43193,N_43020);
xor U43322 (N_43322,N_43118,N_43045);
or U43323 (N_43323,N_43140,N_43034);
nand U43324 (N_43324,N_43243,N_43240);
and U43325 (N_43325,N_43219,N_43202);
nor U43326 (N_43326,N_43137,N_43040);
nand U43327 (N_43327,N_43224,N_43122);
or U43328 (N_43328,N_43070,N_43125);
xnor U43329 (N_43329,N_43133,N_43148);
nand U43330 (N_43330,N_43051,N_43184);
xor U43331 (N_43331,N_43166,N_43163);
nand U43332 (N_43332,N_43157,N_43188);
xor U43333 (N_43333,N_43049,N_43114);
xnor U43334 (N_43334,N_43057,N_43197);
and U43335 (N_43335,N_43221,N_43205);
nand U43336 (N_43336,N_43216,N_43144);
nand U43337 (N_43337,N_43143,N_43162);
xnor U43338 (N_43338,N_43091,N_43218);
and U43339 (N_43339,N_43149,N_43121);
nand U43340 (N_43340,N_43015,N_43226);
and U43341 (N_43341,N_43177,N_43010);
or U43342 (N_43342,N_43039,N_43178);
and U43343 (N_43343,N_43027,N_43241);
and U43344 (N_43344,N_43038,N_43242);
nor U43345 (N_43345,N_43037,N_43167);
nand U43346 (N_43346,N_43012,N_43245);
nor U43347 (N_43347,N_43246,N_43214);
and U43348 (N_43348,N_43128,N_43135);
xor U43349 (N_43349,N_43008,N_43152);
nor U43350 (N_43350,N_43071,N_43001);
or U43351 (N_43351,N_43026,N_43126);
and U43352 (N_43352,N_43211,N_43065);
or U43353 (N_43353,N_43228,N_43136);
xor U43354 (N_43354,N_43072,N_43079);
or U43355 (N_43355,N_43153,N_43009);
nor U43356 (N_43356,N_43156,N_43200);
or U43357 (N_43357,N_43201,N_43195);
and U43358 (N_43358,N_43033,N_43044);
xnor U43359 (N_43359,N_43171,N_43058);
or U43360 (N_43360,N_43032,N_43236);
xnor U43361 (N_43361,N_43107,N_43069);
xnor U43362 (N_43362,N_43123,N_43145);
and U43363 (N_43363,N_43182,N_43217);
nand U43364 (N_43364,N_43204,N_43233);
and U43365 (N_43365,N_43175,N_43083);
xnor U43366 (N_43366,N_43109,N_43248);
and U43367 (N_43367,N_43179,N_43067);
nor U43368 (N_43368,N_43112,N_43002);
or U43369 (N_43369,N_43210,N_43220);
and U43370 (N_43370,N_43225,N_43229);
nor U43371 (N_43371,N_43030,N_43194);
nand U43372 (N_43372,N_43018,N_43043);
and U43373 (N_43373,N_43054,N_43007);
nand U43374 (N_43374,N_43110,N_43227);
and U43375 (N_43375,N_43171,N_43143);
xnor U43376 (N_43376,N_43236,N_43018);
nand U43377 (N_43377,N_43112,N_43135);
xor U43378 (N_43378,N_43067,N_43016);
or U43379 (N_43379,N_43149,N_43176);
or U43380 (N_43380,N_43221,N_43161);
and U43381 (N_43381,N_43185,N_43246);
xnor U43382 (N_43382,N_43165,N_43133);
nor U43383 (N_43383,N_43094,N_43230);
or U43384 (N_43384,N_43210,N_43008);
nand U43385 (N_43385,N_43073,N_43026);
nor U43386 (N_43386,N_43186,N_43063);
nand U43387 (N_43387,N_43040,N_43159);
and U43388 (N_43388,N_43183,N_43035);
and U43389 (N_43389,N_43057,N_43075);
nand U43390 (N_43390,N_43147,N_43198);
nor U43391 (N_43391,N_43008,N_43103);
nand U43392 (N_43392,N_43156,N_43119);
or U43393 (N_43393,N_43041,N_43173);
nand U43394 (N_43394,N_43249,N_43020);
xor U43395 (N_43395,N_43081,N_43162);
or U43396 (N_43396,N_43015,N_43166);
or U43397 (N_43397,N_43200,N_43164);
nand U43398 (N_43398,N_43245,N_43139);
nor U43399 (N_43399,N_43031,N_43249);
nor U43400 (N_43400,N_43239,N_43146);
nor U43401 (N_43401,N_43176,N_43239);
nor U43402 (N_43402,N_43122,N_43011);
xor U43403 (N_43403,N_43109,N_43069);
or U43404 (N_43404,N_43035,N_43133);
and U43405 (N_43405,N_43079,N_43026);
xnor U43406 (N_43406,N_43152,N_43083);
and U43407 (N_43407,N_43168,N_43040);
nor U43408 (N_43408,N_43083,N_43177);
and U43409 (N_43409,N_43041,N_43245);
xor U43410 (N_43410,N_43123,N_43198);
nand U43411 (N_43411,N_43248,N_43132);
and U43412 (N_43412,N_43014,N_43017);
xnor U43413 (N_43413,N_43073,N_43180);
or U43414 (N_43414,N_43037,N_43003);
nor U43415 (N_43415,N_43105,N_43209);
or U43416 (N_43416,N_43228,N_43110);
or U43417 (N_43417,N_43036,N_43074);
or U43418 (N_43418,N_43016,N_43209);
xor U43419 (N_43419,N_43056,N_43174);
nor U43420 (N_43420,N_43132,N_43233);
or U43421 (N_43421,N_43164,N_43007);
or U43422 (N_43422,N_43083,N_43140);
nor U43423 (N_43423,N_43113,N_43009);
and U43424 (N_43424,N_43202,N_43240);
xor U43425 (N_43425,N_43078,N_43013);
and U43426 (N_43426,N_43058,N_43050);
xnor U43427 (N_43427,N_43134,N_43124);
nor U43428 (N_43428,N_43234,N_43223);
nor U43429 (N_43429,N_43075,N_43237);
xnor U43430 (N_43430,N_43009,N_43065);
and U43431 (N_43431,N_43229,N_43089);
or U43432 (N_43432,N_43117,N_43056);
nand U43433 (N_43433,N_43135,N_43094);
xor U43434 (N_43434,N_43002,N_43187);
and U43435 (N_43435,N_43109,N_43118);
nor U43436 (N_43436,N_43085,N_43057);
nand U43437 (N_43437,N_43219,N_43068);
or U43438 (N_43438,N_43219,N_43216);
nor U43439 (N_43439,N_43007,N_43189);
nor U43440 (N_43440,N_43237,N_43162);
nor U43441 (N_43441,N_43059,N_43074);
xnor U43442 (N_43442,N_43165,N_43227);
and U43443 (N_43443,N_43007,N_43203);
or U43444 (N_43444,N_43051,N_43077);
or U43445 (N_43445,N_43029,N_43219);
and U43446 (N_43446,N_43122,N_43203);
or U43447 (N_43447,N_43169,N_43056);
nand U43448 (N_43448,N_43124,N_43054);
nand U43449 (N_43449,N_43032,N_43222);
nor U43450 (N_43450,N_43245,N_43064);
nand U43451 (N_43451,N_43035,N_43154);
nor U43452 (N_43452,N_43116,N_43024);
nor U43453 (N_43453,N_43231,N_43165);
nand U43454 (N_43454,N_43213,N_43132);
and U43455 (N_43455,N_43190,N_43158);
or U43456 (N_43456,N_43002,N_43162);
and U43457 (N_43457,N_43218,N_43099);
xnor U43458 (N_43458,N_43158,N_43017);
and U43459 (N_43459,N_43236,N_43218);
and U43460 (N_43460,N_43171,N_43138);
nor U43461 (N_43461,N_43167,N_43023);
and U43462 (N_43462,N_43053,N_43022);
and U43463 (N_43463,N_43058,N_43025);
xnor U43464 (N_43464,N_43244,N_43045);
or U43465 (N_43465,N_43142,N_43132);
or U43466 (N_43466,N_43034,N_43214);
xor U43467 (N_43467,N_43146,N_43008);
or U43468 (N_43468,N_43021,N_43057);
nand U43469 (N_43469,N_43167,N_43115);
and U43470 (N_43470,N_43161,N_43057);
nor U43471 (N_43471,N_43004,N_43022);
nand U43472 (N_43472,N_43017,N_43218);
xnor U43473 (N_43473,N_43235,N_43071);
or U43474 (N_43474,N_43125,N_43011);
and U43475 (N_43475,N_43054,N_43201);
nor U43476 (N_43476,N_43138,N_43207);
xor U43477 (N_43477,N_43211,N_43245);
nand U43478 (N_43478,N_43141,N_43079);
xor U43479 (N_43479,N_43021,N_43065);
and U43480 (N_43480,N_43082,N_43014);
or U43481 (N_43481,N_43138,N_43021);
or U43482 (N_43482,N_43248,N_43131);
or U43483 (N_43483,N_43192,N_43116);
xnor U43484 (N_43484,N_43051,N_43033);
or U43485 (N_43485,N_43201,N_43119);
nor U43486 (N_43486,N_43050,N_43057);
xnor U43487 (N_43487,N_43102,N_43186);
nor U43488 (N_43488,N_43171,N_43045);
and U43489 (N_43489,N_43059,N_43028);
and U43490 (N_43490,N_43046,N_43151);
or U43491 (N_43491,N_43223,N_43204);
and U43492 (N_43492,N_43183,N_43174);
xor U43493 (N_43493,N_43031,N_43074);
and U43494 (N_43494,N_43249,N_43176);
xor U43495 (N_43495,N_43013,N_43108);
nor U43496 (N_43496,N_43193,N_43141);
xnor U43497 (N_43497,N_43123,N_43117);
nor U43498 (N_43498,N_43081,N_43211);
xor U43499 (N_43499,N_43214,N_43163);
xnor U43500 (N_43500,N_43391,N_43339);
nand U43501 (N_43501,N_43440,N_43389);
and U43502 (N_43502,N_43438,N_43295);
xnor U43503 (N_43503,N_43334,N_43497);
or U43504 (N_43504,N_43360,N_43484);
nand U43505 (N_43505,N_43340,N_43353);
or U43506 (N_43506,N_43271,N_43475);
or U43507 (N_43507,N_43418,N_43373);
nor U43508 (N_43508,N_43363,N_43355);
xnor U43509 (N_43509,N_43432,N_43376);
nor U43510 (N_43510,N_43284,N_43402);
nor U43511 (N_43511,N_43384,N_43368);
nor U43512 (N_43512,N_43419,N_43439);
nand U43513 (N_43513,N_43275,N_43348);
nand U43514 (N_43514,N_43252,N_43278);
xor U43515 (N_43515,N_43277,N_43385);
nor U43516 (N_43516,N_43483,N_43336);
xor U43517 (N_43517,N_43356,N_43319);
or U43518 (N_43518,N_43361,N_43399);
or U43519 (N_43519,N_43480,N_43343);
or U43520 (N_43520,N_43487,N_43297);
nor U43521 (N_43521,N_43309,N_43426);
nand U43522 (N_43522,N_43474,N_43411);
nand U43523 (N_43523,N_43308,N_43272);
xnor U43524 (N_43524,N_43320,N_43362);
and U43525 (N_43525,N_43281,N_43397);
or U43526 (N_43526,N_43366,N_43407);
xnor U43527 (N_43527,N_43381,N_43299);
xor U43528 (N_43528,N_43455,N_43428);
xor U43529 (N_43529,N_43491,N_43494);
nand U43530 (N_43530,N_43372,N_43436);
nor U43531 (N_43531,N_43341,N_43321);
nand U43532 (N_43532,N_43256,N_43267);
nand U43533 (N_43533,N_43324,N_43425);
xor U43534 (N_43534,N_43304,N_43383);
or U43535 (N_43535,N_43456,N_43251);
or U43536 (N_43536,N_43414,N_43467);
and U43537 (N_43537,N_43260,N_43345);
or U43538 (N_43538,N_43280,N_43496);
or U43539 (N_43539,N_43279,N_43250);
nor U43540 (N_43540,N_43378,N_43292);
nor U43541 (N_43541,N_43452,N_43396);
nor U43542 (N_43542,N_43421,N_43283);
or U43543 (N_43543,N_43305,N_43274);
xnor U43544 (N_43544,N_43406,N_43377);
nand U43545 (N_43545,N_43294,N_43329);
and U43546 (N_43546,N_43314,N_43437);
and U43547 (N_43547,N_43315,N_43388);
or U43548 (N_43548,N_43349,N_43394);
nand U43549 (N_43549,N_43403,N_43492);
or U43550 (N_43550,N_43273,N_43479);
and U43551 (N_43551,N_43259,N_43326);
or U43552 (N_43552,N_43293,N_43451);
nand U43553 (N_43553,N_43457,N_43369);
nand U43554 (N_43554,N_43476,N_43422);
and U43555 (N_43555,N_43318,N_43332);
or U43556 (N_43556,N_43431,N_43395);
or U43557 (N_43557,N_43330,N_43257);
nor U43558 (N_43558,N_43380,N_43371);
nor U43559 (N_43559,N_43323,N_43429);
and U43560 (N_43560,N_43253,N_43448);
nand U43561 (N_43561,N_43424,N_43382);
or U43562 (N_43562,N_43453,N_43410);
xor U43563 (N_43563,N_43365,N_43374);
and U43564 (N_43564,N_43352,N_43287);
or U43565 (N_43565,N_43423,N_43450);
xnor U43566 (N_43566,N_43392,N_43490);
and U43567 (N_43567,N_43289,N_43337);
and U43568 (N_43568,N_43335,N_43386);
xnor U43569 (N_43569,N_43291,N_43358);
xor U43570 (N_43570,N_43485,N_43290);
and U43571 (N_43571,N_43357,N_43390);
xnor U43572 (N_43572,N_43322,N_43401);
nand U43573 (N_43573,N_43300,N_43298);
nand U43574 (N_43574,N_43346,N_43409);
nand U43575 (N_43575,N_43460,N_43417);
or U43576 (N_43576,N_43462,N_43364);
xnor U43577 (N_43577,N_43493,N_43351);
or U43578 (N_43578,N_43420,N_43317);
xnor U43579 (N_43579,N_43285,N_43276);
nor U43580 (N_43580,N_43472,N_43473);
nand U43581 (N_43581,N_43446,N_43311);
or U43582 (N_43582,N_43470,N_43435);
xor U43583 (N_43583,N_43254,N_43313);
nor U43584 (N_43584,N_43264,N_43310);
or U43585 (N_43585,N_43255,N_43302);
and U43586 (N_43586,N_43408,N_43413);
xor U43587 (N_43587,N_43328,N_43379);
nor U43588 (N_43588,N_43306,N_43464);
nor U43589 (N_43589,N_43375,N_43288);
nor U43590 (N_43590,N_43477,N_43282);
nor U43591 (N_43591,N_43301,N_43303);
or U43592 (N_43592,N_43478,N_43465);
and U43593 (N_43593,N_43441,N_43458);
xor U43594 (N_43594,N_43482,N_43404);
or U43595 (N_43595,N_43486,N_43489);
or U43596 (N_43596,N_43498,N_43427);
xor U43597 (N_43597,N_43443,N_43488);
or U43598 (N_43598,N_43263,N_43459);
nand U43599 (N_43599,N_43433,N_43481);
or U43600 (N_43600,N_43350,N_43359);
nand U43601 (N_43601,N_43387,N_43444);
nor U43602 (N_43602,N_43412,N_43461);
nand U43603 (N_43603,N_43415,N_43463);
xor U43604 (N_43604,N_43342,N_43331);
or U43605 (N_43605,N_43258,N_43434);
or U43606 (N_43606,N_43327,N_43499);
nor U43607 (N_43607,N_43445,N_43312);
nor U43608 (N_43608,N_43398,N_43393);
nand U43609 (N_43609,N_43454,N_43269);
nor U43610 (N_43610,N_43296,N_43370);
and U43611 (N_43611,N_43266,N_43367);
and U43612 (N_43612,N_43265,N_43286);
xor U43613 (N_43613,N_43316,N_43262);
or U43614 (N_43614,N_43354,N_43468);
nand U43615 (N_43615,N_43347,N_43268);
xor U43616 (N_43616,N_43344,N_43416);
nor U43617 (N_43617,N_43466,N_43333);
xnor U43618 (N_43618,N_43270,N_43469);
and U43619 (N_43619,N_43400,N_43325);
nand U43620 (N_43620,N_43307,N_43495);
or U43621 (N_43621,N_43447,N_43430);
xor U43622 (N_43622,N_43449,N_43261);
nor U43623 (N_43623,N_43405,N_43338);
xnor U43624 (N_43624,N_43471,N_43442);
and U43625 (N_43625,N_43395,N_43265);
or U43626 (N_43626,N_43411,N_43410);
xor U43627 (N_43627,N_43325,N_43442);
or U43628 (N_43628,N_43498,N_43465);
nor U43629 (N_43629,N_43495,N_43377);
nand U43630 (N_43630,N_43329,N_43403);
or U43631 (N_43631,N_43278,N_43379);
xor U43632 (N_43632,N_43368,N_43291);
nand U43633 (N_43633,N_43345,N_43378);
xor U43634 (N_43634,N_43354,N_43322);
and U43635 (N_43635,N_43375,N_43403);
nor U43636 (N_43636,N_43321,N_43423);
or U43637 (N_43637,N_43381,N_43444);
or U43638 (N_43638,N_43357,N_43329);
xor U43639 (N_43639,N_43328,N_43419);
and U43640 (N_43640,N_43432,N_43445);
nand U43641 (N_43641,N_43320,N_43466);
nand U43642 (N_43642,N_43259,N_43301);
or U43643 (N_43643,N_43310,N_43405);
nand U43644 (N_43644,N_43478,N_43429);
and U43645 (N_43645,N_43460,N_43256);
nand U43646 (N_43646,N_43285,N_43344);
xor U43647 (N_43647,N_43317,N_43305);
and U43648 (N_43648,N_43374,N_43306);
xnor U43649 (N_43649,N_43409,N_43276);
xnor U43650 (N_43650,N_43475,N_43283);
xor U43651 (N_43651,N_43265,N_43353);
nand U43652 (N_43652,N_43422,N_43390);
nor U43653 (N_43653,N_43479,N_43395);
and U43654 (N_43654,N_43331,N_43462);
and U43655 (N_43655,N_43302,N_43470);
xnor U43656 (N_43656,N_43312,N_43268);
nor U43657 (N_43657,N_43300,N_43451);
and U43658 (N_43658,N_43336,N_43356);
xor U43659 (N_43659,N_43256,N_43438);
or U43660 (N_43660,N_43438,N_43316);
nand U43661 (N_43661,N_43392,N_43331);
and U43662 (N_43662,N_43442,N_43397);
xnor U43663 (N_43663,N_43443,N_43316);
and U43664 (N_43664,N_43392,N_43279);
and U43665 (N_43665,N_43461,N_43449);
nand U43666 (N_43666,N_43407,N_43314);
and U43667 (N_43667,N_43410,N_43333);
and U43668 (N_43668,N_43335,N_43267);
or U43669 (N_43669,N_43438,N_43428);
nand U43670 (N_43670,N_43310,N_43257);
xnor U43671 (N_43671,N_43445,N_43458);
nor U43672 (N_43672,N_43478,N_43402);
xnor U43673 (N_43673,N_43323,N_43316);
and U43674 (N_43674,N_43364,N_43372);
nor U43675 (N_43675,N_43474,N_43423);
nand U43676 (N_43676,N_43319,N_43456);
nand U43677 (N_43677,N_43298,N_43493);
xor U43678 (N_43678,N_43427,N_43398);
nand U43679 (N_43679,N_43444,N_43418);
xor U43680 (N_43680,N_43365,N_43258);
nand U43681 (N_43681,N_43454,N_43442);
or U43682 (N_43682,N_43251,N_43398);
or U43683 (N_43683,N_43459,N_43417);
or U43684 (N_43684,N_43272,N_43410);
and U43685 (N_43685,N_43294,N_43325);
or U43686 (N_43686,N_43495,N_43315);
xnor U43687 (N_43687,N_43273,N_43284);
or U43688 (N_43688,N_43468,N_43274);
nor U43689 (N_43689,N_43370,N_43271);
or U43690 (N_43690,N_43472,N_43496);
nand U43691 (N_43691,N_43278,N_43436);
or U43692 (N_43692,N_43357,N_43331);
and U43693 (N_43693,N_43446,N_43326);
or U43694 (N_43694,N_43272,N_43393);
or U43695 (N_43695,N_43366,N_43257);
nor U43696 (N_43696,N_43436,N_43362);
nor U43697 (N_43697,N_43340,N_43438);
nor U43698 (N_43698,N_43366,N_43428);
nand U43699 (N_43699,N_43264,N_43371);
or U43700 (N_43700,N_43450,N_43276);
nand U43701 (N_43701,N_43462,N_43345);
nor U43702 (N_43702,N_43479,N_43478);
xor U43703 (N_43703,N_43301,N_43331);
nor U43704 (N_43704,N_43285,N_43257);
nand U43705 (N_43705,N_43464,N_43316);
nand U43706 (N_43706,N_43486,N_43307);
or U43707 (N_43707,N_43476,N_43408);
and U43708 (N_43708,N_43409,N_43456);
xor U43709 (N_43709,N_43402,N_43274);
nand U43710 (N_43710,N_43267,N_43323);
nor U43711 (N_43711,N_43345,N_43448);
or U43712 (N_43712,N_43346,N_43442);
nor U43713 (N_43713,N_43463,N_43483);
nand U43714 (N_43714,N_43330,N_43331);
nand U43715 (N_43715,N_43294,N_43376);
and U43716 (N_43716,N_43486,N_43425);
nand U43717 (N_43717,N_43418,N_43420);
and U43718 (N_43718,N_43254,N_43280);
or U43719 (N_43719,N_43378,N_43327);
nand U43720 (N_43720,N_43428,N_43453);
nor U43721 (N_43721,N_43483,N_43268);
or U43722 (N_43722,N_43396,N_43338);
and U43723 (N_43723,N_43478,N_43457);
nor U43724 (N_43724,N_43479,N_43426);
xor U43725 (N_43725,N_43437,N_43482);
and U43726 (N_43726,N_43354,N_43464);
nand U43727 (N_43727,N_43286,N_43453);
xor U43728 (N_43728,N_43291,N_43361);
nor U43729 (N_43729,N_43484,N_43413);
xor U43730 (N_43730,N_43420,N_43291);
xor U43731 (N_43731,N_43487,N_43468);
and U43732 (N_43732,N_43315,N_43471);
or U43733 (N_43733,N_43444,N_43271);
nor U43734 (N_43734,N_43473,N_43337);
nor U43735 (N_43735,N_43466,N_43337);
xor U43736 (N_43736,N_43490,N_43304);
or U43737 (N_43737,N_43329,N_43384);
nor U43738 (N_43738,N_43425,N_43285);
nand U43739 (N_43739,N_43268,N_43495);
xor U43740 (N_43740,N_43481,N_43266);
xnor U43741 (N_43741,N_43309,N_43468);
nand U43742 (N_43742,N_43424,N_43310);
or U43743 (N_43743,N_43402,N_43294);
or U43744 (N_43744,N_43320,N_43281);
nor U43745 (N_43745,N_43279,N_43467);
nand U43746 (N_43746,N_43311,N_43491);
or U43747 (N_43747,N_43306,N_43451);
xor U43748 (N_43748,N_43282,N_43399);
xnor U43749 (N_43749,N_43255,N_43329);
xnor U43750 (N_43750,N_43693,N_43543);
and U43751 (N_43751,N_43646,N_43506);
and U43752 (N_43752,N_43664,N_43630);
nand U43753 (N_43753,N_43603,N_43586);
and U43754 (N_43754,N_43544,N_43721);
xor U43755 (N_43755,N_43591,N_43580);
and U43756 (N_43756,N_43548,N_43515);
and U43757 (N_43757,N_43676,N_43529);
or U43758 (N_43758,N_43553,N_43554);
xnor U43759 (N_43759,N_43604,N_43648);
or U43760 (N_43760,N_43702,N_43717);
nand U43761 (N_43761,N_43679,N_43734);
xor U43762 (N_43762,N_43527,N_43537);
nor U43763 (N_43763,N_43590,N_43598);
nand U43764 (N_43764,N_43644,N_43657);
xor U43765 (N_43765,N_43671,N_43565);
nand U43766 (N_43766,N_43577,N_43612);
nand U43767 (N_43767,N_43561,N_43592);
xnor U43768 (N_43768,N_43621,N_43663);
or U43769 (N_43769,N_43535,N_43528);
and U43770 (N_43770,N_43669,N_43678);
xor U43771 (N_43771,N_43504,N_43729);
and U43772 (N_43772,N_43708,N_43516);
or U43773 (N_43773,N_43631,N_43731);
nand U43774 (N_43774,N_43625,N_43611);
xor U43775 (N_43775,N_43524,N_43705);
or U43776 (N_43776,N_43744,N_43655);
nand U43777 (N_43777,N_43651,N_43736);
or U43778 (N_43778,N_43560,N_43667);
and U43779 (N_43779,N_43526,N_43509);
or U43780 (N_43780,N_43519,N_43672);
nor U43781 (N_43781,N_43733,N_43722);
or U43782 (N_43782,N_43587,N_43732);
xor U43783 (N_43783,N_43562,N_43707);
or U43784 (N_43784,N_43510,N_43634);
or U43785 (N_43785,N_43617,N_43737);
or U43786 (N_43786,N_43596,N_43607);
nor U43787 (N_43787,N_43749,N_43579);
nand U43788 (N_43788,N_43665,N_43581);
and U43789 (N_43789,N_43572,N_43501);
xor U43790 (N_43790,N_43532,N_43718);
nor U43791 (N_43791,N_43706,N_43574);
or U43792 (N_43792,N_43658,N_43575);
nand U43793 (N_43793,N_43578,N_43525);
nand U43794 (N_43794,N_43719,N_43571);
nand U43795 (N_43795,N_43688,N_43601);
and U43796 (N_43796,N_43726,N_43549);
nand U43797 (N_43797,N_43654,N_43710);
and U43798 (N_43798,N_43689,N_43683);
nor U43799 (N_43799,N_43594,N_43584);
and U43800 (N_43800,N_43540,N_43521);
nor U43801 (N_43801,N_43716,N_43588);
or U43802 (N_43802,N_43724,N_43536);
or U43803 (N_43803,N_43551,N_43725);
and U43804 (N_43804,N_43545,N_43686);
and U43805 (N_43805,N_43660,N_43567);
nand U43806 (N_43806,N_43748,N_43712);
xnor U43807 (N_43807,N_43653,N_43699);
nor U43808 (N_43808,N_43739,N_43583);
or U43809 (N_43809,N_43659,N_43742);
nand U43810 (N_43810,N_43640,N_43512);
nand U43811 (N_43811,N_43517,N_43511);
or U43812 (N_43812,N_43636,N_43747);
xor U43813 (N_43813,N_43623,N_43627);
nor U43814 (N_43814,N_43703,N_43616);
nand U43815 (N_43815,N_43620,N_43690);
and U43816 (N_43816,N_43670,N_43643);
and U43817 (N_43817,N_43738,N_43728);
or U43818 (N_43818,N_43568,N_43605);
or U43819 (N_43819,N_43713,N_43589);
or U43820 (N_43820,N_43522,N_43505);
nand U43821 (N_43821,N_43635,N_43582);
nor U43822 (N_43822,N_43730,N_43557);
and U43823 (N_43823,N_43656,N_43714);
nor U43824 (N_43824,N_43639,N_43727);
nand U43825 (N_43825,N_43685,N_43559);
nor U43826 (N_43826,N_43619,N_43741);
or U43827 (N_43827,N_43652,N_43618);
nand U43828 (N_43828,N_43723,N_43662);
nor U43829 (N_43829,N_43704,N_43602);
or U43830 (N_43830,N_43573,N_43599);
nand U43831 (N_43831,N_43502,N_43694);
nand U43832 (N_43832,N_43523,N_43614);
nor U43833 (N_43833,N_43638,N_43508);
xor U43834 (N_43834,N_43666,N_43696);
and U43835 (N_43835,N_43606,N_43675);
xnor U43836 (N_43836,N_43609,N_43624);
nand U43837 (N_43837,N_43746,N_43740);
or U43838 (N_43838,N_43674,N_43701);
nor U43839 (N_43839,N_43682,N_43613);
nor U43840 (N_43840,N_43745,N_43628);
nor U43841 (N_43841,N_43680,N_43534);
nor U43842 (N_43842,N_43615,N_43673);
nor U43843 (N_43843,N_43700,N_43556);
nand U43844 (N_43844,N_43697,N_43610);
nor U43845 (N_43845,N_43570,N_43743);
nand U43846 (N_43846,N_43563,N_43661);
xor U43847 (N_43847,N_43569,N_43629);
or U43848 (N_43848,N_43691,N_43626);
and U43849 (N_43849,N_43695,N_43715);
nand U43850 (N_43850,N_43711,N_43542);
nor U43851 (N_43851,N_43514,N_43552);
nand U43852 (N_43852,N_43555,N_43550);
and U43853 (N_43853,N_43507,N_43709);
nor U43854 (N_43854,N_43720,N_43649);
xor U43855 (N_43855,N_43642,N_43595);
nand U43856 (N_43856,N_43645,N_43593);
xnor U43857 (N_43857,N_43632,N_43564);
and U43858 (N_43858,N_43668,N_43531);
xor U43859 (N_43859,N_43558,N_43513);
xor U43860 (N_43860,N_43541,N_43547);
nand U43861 (N_43861,N_43647,N_43698);
nand U43862 (N_43862,N_43684,N_43566);
and U43863 (N_43863,N_43597,N_43622);
nor U43864 (N_43864,N_43503,N_43518);
xor U43865 (N_43865,N_43520,N_43608);
nor U43866 (N_43866,N_43500,N_43539);
nand U43867 (N_43867,N_43633,N_43538);
xnor U43868 (N_43868,N_43687,N_43585);
or U43869 (N_43869,N_43681,N_43576);
nand U43870 (N_43870,N_43692,N_43677);
and U43871 (N_43871,N_43546,N_43650);
nor U43872 (N_43872,N_43600,N_43530);
xor U43873 (N_43873,N_43735,N_43533);
xor U43874 (N_43874,N_43637,N_43641);
xor U43875 (N_43875,N_43593,N_43693);
xnor U43876 (N_43876,N_43548,N_43722);
and U43877 (N_43877,N_43730,N_43746);
nand U43878 (N_43878,N_43739,N_43533);
nand U43879 (N_43879,N_43515,N_43724);
xor U43880 (N_43880,N_43586,N_43724);
xnor U43881 (N_43881,N_43628,N_43608);
or U43882 (N_43882,N_43709,N_43676);
nand U43883 (N_43883,N_43509,N_43539);
and U43884 (N_43884,N_43693,N_43619);
xor U43885 (N_43885,N_43525,N_43694);
nor U43886 (N_43886,N_43518,N_43730);
nor U43887 (N_43887,N_43589,N_43569);
xnor U43888 (N_43888,N_43530,N_43575);
nor U43889 (N_43889,N_43588,N_43734);
nor U43890 (N_43890,N_43542,N_43577);
nor U43891 (N_43891,N_43591,N_43541);
nor U43892 (N_43892,N_43526,N_43669);
and U43893 (N_43893,N_43676,N_43637);
nor U43894 (N_43894,N_43702,N_43565);
or U43895 (N_43895,N_43560,N_43538);
or U43896 (N_43896,N_43534,N_43565);
xor U43897 (N_43897,N_43580,N_43593);
and U43898 (N_43898,N_43534,N_43543);
xor U43899 (N_43899,N_43732,N_43747);
nor U43900 (N_43900,N_43502,N_43683);
nand U43901 (N_43901,N_43677,N_43672);
or U43902 (N_43902,N_43630,N_43643);
xor U43903 (N_43903,N_43739,N_43661);
nor U43904 (N_43904,N_43535,N_43582);
and U43905 (N_43905,N_43632,N_43665);
xnor U43906 (N_43906,N_43532,N_43508);
xnor U43907 (N_43907,N_43707,N_43667);
nand U43908 (N_43908,N_43662,N_43554);
nand U43909 (N_43909,N_43510,N_43722);
nand U43910 (N_43910,N_43525,N_43703);
and U43911 (N_43911,N_43706,N_43539);
xnor U43912 (N_43912,N_43578,N_43509);
nand U43913 (N_43913,N_43703,N_43560);
and U43914 (N_43914,N_43677,N_43614);
nor U43915 (N_43915,N_43554,N_43748);
and U43916 (N_43916,N_43524,N_43545);
or U43917 (N_43917,N_43566,N_43688);
nand U43918 (N_43918,N_43672,N_43615);
nand U43919 (N_43919,N_43673,N_43608);
or U43920 (N_43920,N_43738,N_43721);
nor U43921 (N_43921,N_43554,N_43556);
or U43922 (N_43922,N_43670,N_43651);
or U43923 (N_43923,N_43702,N_43525);
xor U43924 (N_43924,N_43591,N_43588);
and U43925 (N_43925,N_43546,N_43648);
and U43926 (N_43926,N_43500,N_43731);
nor U43927 (N_43927,N_43658,N_43586);
and U43928 (N_43928,N_43518,N_43704);
nor U43929 (N_43929,N_43621,N_43649);
xor U43930 (N_43930,N_43649,N_43622);
and U43931 (N_43931,N_43572,N_43621);
nand U43932 (N_43932,N_43712,N_43669);
nor U43933 (N_43933,N_43746,N_43585);
nor U43934 (N_43934,N_43600,N_43595);
xor U43935 (N_43935,N_43580,N_43627);
nand U43936 (N_43936,N_43656,N_43580);
nand U43937 (N_43937,N_43515,N_43735);
xor U43938 (N_43938,N_43537,N_43708);
or U43939 (N_43939,N_43541,N_43668);
nand U43940 (N_43940,N_43591,N_43535);
and U43941 (N_43941,N_43638,N_43575);
nor U43942 (N_43942,N_43734,N_43652);
nand U43943 (N_43943,N_43679,N_43675);
xnor U43944 (N_43944,N_43644,N_43662);
nand U43945 (N_43945,N_43735,N_43728);
nand U43946 (N_43946,N_43700,N_43553);
xor U43947 (N_43947,N_43559,N_43633);
xnor U43948 (N_43948,N_43624,N_43617);
and U43949 (N_43949,N_43729,N_43683);
nor U43950 (N_43950,N_43730,N_43614);
or U43951 (N_43951,N_43656,N_43569);
nor U43952 (N_43952,N_43610,N_43525);
nand U43953 (N_43953,N_43693,N_43606);
or U43954 (N_43954,N_43630,N_43568);
or U43955 (N_43955,N_43748,N_43555);
or U43956 (N_43956,N_43651,N_43693);
nor U43957 (N_43957,N_43647,N_43676);
or U43958 (N_43958,N_43715,N_43541);
nand U43959 (N_43959,N_43556,N_43710);
or U43960 (N_43960,N_43549,N_43625);
and U43961 (N_43961,N_43598,N_43576);
nor U43962 (N_43962,N_43660,N_43513);
nor U43963 (N_43963,N_43669,N_43507);
nor U43964 (N_43964,N_43665,N_43508);
nand U43965 (N_43965,N_43739,N_43721);
xnor U43966 (N_43966,N_43700,N_43662);
nor U43967 (N_43967,N_43693,N_43682);
xor U43968 (N_43968,N_43576,N_43608);
and U43969 (N_43969,N_43590,N_43583);
nand U43970 (N_43970,N_43591,N_43694);
xnor U43971 (N_43971,N_43687,N_43570);
xnor U43972 (N_43972,N_43585,N_43506);
xor U43973 (N_43973,N_43620,N_43747);
nand U43974 (N_43974,N_43687,N_43600);
and U43975 (N_43975,N_43507,N_43646);
and U43976 (N_43976,N_43746,N_43511);
nand U43977 (N_43977,N_43580,N_43734);
and U43978 (N_43978,N_43712,N_43639);
nand U43979 (N_43979,N_43653,N_43718);
nor U43980 (N_43980,N_43500,N_43522);
or U43981 (N_43981,N_43684,N_43712);
nand U43982 (N_43982,N_43708,N_43745);
nand U43983 (N_43983,N_43683,N_43548);
or U43984 (N_43984,N_43618,N_43722);
or U43985 (N_43985,N_43698,N_43718);
nor U43986 (N_43986,N_43518,N_43514);
and U43987 (N_43987,N_43695,N_43617);
xnor U43988 (N_43988,N_43629,N_43665);
and U43989 (N_43989,N_43534,N_43617);
and U43990 (N_43990,N_43524,N_43560);
and U43991 (N_43991,N_43655,N_43505);
nor U43992 (N_43992,N_43512,N_43709);
nor U43993 (N_43993,N_43597,N_43534);
nor U43994 (N_43994,N_43608,N_43516);
nor U43995 (N_43995,N_43515,N_43608);
xnor U43996 (N_43996,N_43644,N_43659);
xor U43997 (N_43997,N_43501,N_43578);
nor U43998 (N_43998,N_43589,N_43739);
xor U43999 (N_43999,N_43527,N_43521);
nand U44000 (N_44000,N_43927,N_43940);
xor U44001 (N_44001,N_43791,N_43951);
or U44002 (N_44002,N_43928,N_43878);
xnor U44003 (N_44003,N_43916,N_43958);
or U44004 (N_44004,N_43873,N_43967);
nor U44005 (N_44005,N_43972,N_43908);
or U44006 (N_44006,N_43917,N_43897);
and U44007 (N_44007,N_43919,N_43805);
nor U44008 (N_44008,N_43876,N_43865);
xnor U44009 (N_44009,N_43808,N_43848);
and U44010 (N_44010,N_43936,N_43816);
nand U44011 (N_44011,N_43771,N_43831);
nor U44012 (N_44012,N_43989,N_43993);
and U44013 (N_44013,N_43773,N_43900);
and U44014 (N_44014,N_43861,N_43923);
and U44015 (N_44015,N_43815,N_43851);
nand U44016 (N_44016,N_43870,N_43864);
or U44017 (N_44017,N_43968,N_43941);
nand U44018 (N_44018,N_43899,N_43948);
nand U44019 (N_44019,N_43889,N_43838);
nor U44020 (N_44020,N_43798,N_43888);
nor U44021 (N_44021,N_43860,N_43754);
xor U44022 (N_44022,N_43772,N_43759);
xor U44023 (N_44023,N_43783,N_43953);
or U44024 (N_44024,N_43938,N_43866);
nor U44025 (N_44025,N_43875,N_43949);
or U44026 (N_44026,N_43843,N_43869);
nor U44027 (N_44027,N_43756,N_43966);
nand U44028 (N_44028,N_43884,N_43987);
and U44029 (N_44029,N_43804,N_43852);
and U44030 (N_44030,N_43982,N_43867);
xor U44031 (N_44031,N_43956,N_43925);
xor U44032 (N_44032,N_43767,N_43763);
nand U44033 (N_44033,N_43766,N_43817);
nor U44034 (N_44034,N_43818,N_43887);
and U44035 (N_44035,N_43809,N_43904);
xnor U44036 (N_44036,N_43957,N_43932);
nand U44037 (N_44037,N_43833,N_43994);
xnor U44038 (N_44038,N_43862,N_43942);
xnor U44039 (N_44039,N_43820,N_43929);
nor U44040 (N_44040,N_43837,N_43910);
or U44041 (N_44041,N_43827,N_43841);
or U44042 (N_44042,N_43881,N_43825);
nor U44043 (N_44043,N_43947,N_43757);
nand U44044 (N_44044,N_43935,N_43988);
and U44045 (N_44045,N_43853,N_43937);
nor U44046 (N_44046,N_43981,N_43903);
or U44047 (N_44047,N_43905,N_43964);
nand U44048 (N_44048,N_43859,N_43915);
and U44049 (N_44049,N_43943,N_43777);
and U44050 (N_44050,N_43890,N_43883);
nand U44051 (N_44051,N_43855,N_43984);
xnor U44052 (N_44052,N_43781,N_43785);
xnor U44053 (N_44053,N_43946,N_43882);
nor U44054 (N_44054,N_43811,N_43802);
nand U44055 (N_44055,N_43832,N_43793);
nand U44056 (N_44056,N_43921,N_43834);
and U44057 (N_44057,N_43877,N_43758);
nor U44058 (N_44058,N_43858,N_43906);
nand U44059 (N_44059,N_43800,N_43991);
and U44060 (N_44060,N_43914,N_43891);
or U44061 (N_44061,N_43918,N_43770);
xor U44062 (N_44062,N_43954,N_43774);
nand U44063 (N_44063,N_43750,N_43846);
nand U44064 (N_44064,N_43874,N_43795);
and U44065 (N_44065,N_43896,N_43835);
or U44066 (N_44066,N_43769,N_43751);
nor U44067 (N_44067,N_43924,N_43965);
nand U44068 (N_44068,N_43780,N_43779);
or U44069 (N_44069,N_43911,N_43907);
or U44070 (N_44070,N_43952,N_43782);
nor U44071 (N_44071,N_43973,N_43999);
nor U44072 (N_44072,N_43950,N_43930);
nand U44073 (N_44073,N_43912,N_43845);
xnor U44074 (N_44074,N_43819,N_43979);
or U44075 (N_44075,N_43892,N_43787);
or U44076 (N_44076,N_43898,N_43776);
nand U44077 (N_44077,N_43985,N_43944);
or U44078 (N_44078,N_43803,N_43926);
and U44079 (N_44079,N_43960,N_43807);
or U44080 (N_44080,N_43920,N_43857);
xor U44081 (N_44081,N_43792,N_43755);
nor U44082 (N_44082,N_43856,N_43998);
xnor U44083 (N_44083,N_43871,N_43799);
or U44084 (N_44084,N_43959,N_43922);
nor U44085 (N_44085,N_43901,N_43753);
nand U44086 (N_44086,N_43879,N_43868);
nor U44087 (N_44087,N_43830,N_43761);
and U44088 (N_44088,N_43764,N_43933);
nand U44089 (N_44089,N_43854,N_43885);
nand U44090 (N_44090,N_43978,N_43789);
or U44091 (N_44091,N_43801,N_43863);
and U44092 (N_44092,N_43934,N_43939);
or U44093 (N_44093,N_43963,N_43806);
and U44094 (N_44094,N_43955,N_43880);
xnor U44095 (N_44095,N_43823,N_43962);
nand U44096 (N_44096,N_43977,N_43992);
xor U44097 (N_44097,N_43849,N_43828);
and U44098 (N_44098,N_43821,N_43762);
xor U44099 (N_44099,N_43990,N_43765);
or U44100 (N_44100,N_43796,N_43894);
and U44101 (N_44101,N_43840,N_43931);
or U44102 (N_44102,N_43760,N_43961);
nand U44103 (N_44103,N_43822,N_43986);
xor U44104 (N_44104,N_43970,N_43975);
nor U44105 (N_44105,N_43974,N_43893);
xor U44106 (N_44106,N_43797,N_43829);
nor U44107 (N_44107,N_43997,N_43980);
xnor U44108 (N_44108,N_43788,N_43886);
or U44109 (N_44109,N_43786,N_43971);
and U44110 (N_44110,N_43895,N_43768);
nor U44111 (N_44111,N_43812,N_43969);
or U44112 (N_44112,N_43995,N_43842);
or U44113 (N_44113,N_43752,N_43839);
or U44114 (N_44114,N_43850,N_43983);
nor U44115 (N_44115,N_43824,N_43913);
xnor U44116 (N_44116,N_43847,N_43810);
nand U44117 (N_44117,N_43976,N_43813);
and U44118 (N_44118,N_43945,N_43872);
and U44119 (N_44119,N_43775,N_43826);
nor U44120 (N_44120,N_43902,N_43784);
nand U44121 (N_44121,N_43814,N_43836);
and U44122 (N_44122,N_43790,N_43996);
nand U44123 (N_44123,N_43909,N_43844);
xor U44124 (N_44124,N_43794,N_43778);
and U44125 (N_44125,N_43823,N_43790);
and U44126 (N_44126,N_43824,N_43955);
and U44127 (N_44127,N_43861,N_43806);
xnor U44128 (N_44128,N_43770,N_43795);
or U44129 (N_44129,N_43880,N_43875);
and U44130 (N_44130,N_43774,N_43765);
nand U44131 (N_44131,N_43826,N_43841);
nor U44132 (N_44132,N_43841,N_43797);
nand U44133 (N_44133,N_43757,N_43986);
or U44134 (N_44134,N_43851,N_43965);
nand U44135 (N_44135,N_43923,N_43866);
nor U44136 (N_44136,N_43916,N_43953);
nor U44137 (N_44137,N_43920,N_43872);
xor U44138 (N_44138,N_43910,N_43887);
or U44139 (N_44139,N_43814,N_43880);
or U44140 (N_44140,N_43786,N_43915);
or U44141 (N_44141,N_43965,N_43927);
or U44142 (N_44142,N_43924,N_43934);
nor U44143 (N_44143,N_43823,N_43855);
nand U44144 (N_44144,N_43939,N_43959);
nand U44145 (N_44145,N_43816,N_43801);
or U44146 (N_44146,N_43909,N_43822);
and U44147 (N_44147,N_43814,N_43952);
or U44148 (N_44148,N_43967,N_43843);
or U44149 (N_44149,N_43768,N_43901);
nor U44150 (N_44150,N_43936,N_43841);
and U44151 (N_44151,N_43934,N_43770);
nand U44152 (N_44152,N_43999,N_43834);
xor U44153 (N_44153,N_43755,N_43851);
xor U44154 (N_44154,N_43976,N_43949);
nand U44155 (N_44155,N_43942,N_43946);
xnor U44156 (N_44156,N_43934,N_43919);
and U44157 (N_44157,N_43888,N_43958);
and U44158 (N_44158,N_43861,N_43813);
nor U44159 (N_44159,N_43789,N_43835);
nand U44160 (N_44160,N_43949,N_43954);
xor U44161 (N_44161,N_43883,N_43928);
or U44162 (N_44162,N_43823,N_43909);
or U44163 (N_44163,N_43991,N_43782);
nor U44164 (N_44164,N_43783,N_43903);
nor U44165 (N_44165,N_43822,N_43870);
and U44166 (N_44166,N_43859,N_43923);
and U44167 (N_44167,N_43976,N_43893);
xor U44168 (N_44168,N_43781,N_43818);
nand U44169 (N_44169,N_43812,N_43852);
xor U44170 (N_44170,N_43794,N_43951);
or U44171 (N_44171,N_43883,N_43750);
nor U44172 (N_44172,N_43961,N_43852);
nor U44173 (N_44173,N_43771,N_43978);
or U44174 (N_44174,N_43861,N_43777);
xnor U44175 (N_44175,N_43924,N_43911);
xnor U44176 (N_44176,N_43824,N_43795);
xnor U44177 (N_44177,N_43910,N_43771);
or U44178 (N_44178,N_43979,N_43949);
nand U44179 (N_44179,N_43996,N_43977);
nand U44180 (N_44180,N_43820,N_43971);
and U44181 (N_44181,N_43773,N_43934);
nand U44182 (N_44182,N_43872,N_43826);
or U44183 (N_44183,N_43789,N_43788);
xnor U44184 (N_44184,N_43980,N_43919);
and U44185 (N_44185,N_43771,N_43785);
nor U44186 (N_44186,N_43790,N_43863);
nand U44187 (N_44187,N_43803,N_43901);
nand U44188 (N_44188,N_43754,N_43802);
nor U44189 (N_44189,N_43925,N_43917);
nor U44190 (N_44190,N_43970,N_43750);
xor U44191 (N_44191,N_43860,N_43904);
nor U44192 (N_44192,N_43797,N_43843);
or U44193 (N_44193,N_43755,N_43886);
nand U44194 (N_44194,N_43858,N_43809);
nand U44195 (N_44195,N_43950,N_43999);
and U44196 (N_44196,N_43888,N_43821);
and U44197 (N_44197,N_43864,N_43857);
or U44198 (N_44198,N_43793,N_43788);
nand U44199 (N_44199,N_43827,N_43850);
xor U44200 (N_44200,N_43881,N_43821);
or U44201 (N_44201,N_43904,N_43784);
xor U44202 (N_44202,N_43811,N_43902);
or U44203 (N_44203,N_43881,N_43909);
nor U44204 (N_44204,N_43885,N_43821);
and U44205 (N_44205,N_43961,N_43977);
xnor U44206 (N_44206,N_43780,N_43893);
or U44207 (N_44207,N_43893,N_43940);
xnor U44208 (N_44208,N_43867,N_43914);
nand U44209 (N_44209,N_43785,N_43871);
or U44210 (N_44210,N_43846,N_43959);
or U44211 (N_44211,N_43793,N_43951);
and U44212 (N_44212,N_43927,N_43960);
xnor U44213 (N_44213,N_43803,N_43912);
nor U44214 (N_44214,N_43964,N_43883);
nor U44215 (N_44215,N_43815,N_43790);
xor U44216 (N_44216,N_43880,N_43877);
or U44217 (N_44217,N_43928,N_43811);
and U44218 (N_44218,N_43890,N_43865);
nor U44219 (N_44219,N_43894,N_43957);
nand U44220 (N_44220,N_43825,N_43786);
nor U44221 (N_44221,N_43767,N_43995);
xor U44222 (N_44222,N_43981,N_43770);
or U44223 (N_44223,N_43791,N_43849);
nor U44224 (N_44224,N_43791,N_43952);
nand U44225 (N_44225,N_43981,N_43938);
or U44226 (N_44226,N_43938,N_43909);
or U44227 (N_44227,N_43795,N_43994);
nor U44228 (N_44228,N_43963,N_43798);
and U44229 (N_44229,N_43933,N_43803);
nor U44230 (N_44230,N_43761,N_43835);
xor U44231 (N_44231,N_43876,N_43921);
xnor U44232 (N_44232,N_43862,N_43767);
and U44233 (N_44233,N_43860,N_43768);
and U44234 (N_44234,N_43875,N_43928);
and U44235 (N_44235,N_43881,N_43925);
and U44236 (N_44236,N_43959,N_43941);
nand U44237 (N_44237,N_43774,N_43936);
nor U44238 (N_44238,N_43864,N_43770);
nand U44239 (N_44239,N_43792,N_43969);
or U44240 (N_44240,N_43948,N_43906);
or U44241 (N_44241,N_43887,N_43978);
or U44242 (N_44242,N_43941,N_43892);
and U44243 (N_44243,N_43856,N_43832);
and U44244 (N_44244,N_43977,N_43910);
nand U44245 (N_44245,N_43884,N_43758);
nor U44246 (N_44246,N_43990,N_43973);
nor U44247 (N_44247,N_43932,N_43813);
nor U44248 (N_44248,N_43961,N_43950);
nor U44249 (N_44249,N_43751,N_43898);
xnor U44250 (N_44250,N_44106,N_44172);
nor U44251 (N_44251,N_44022,N_44230);
nor U44252 (N_44252,N_44203,N_44048);
or U44253 (N_44253,N_44213,N_44136);
and U44254 (N_44254,N_44241,N_44159);
nand U44255 (N_44255,N_44229,N_44085);
and U44256 (N_44256,N_44031,N_44070);
xnor U44257 (N_44257,N_44118,N_44166);
nor U44258 (N_44258,N_44157,N_44043);
nor U44259 (N_44259,N_44158,N_44001);
nor U44260 (N_44260,N_44000,N_44104);
and U44261 (N_44261,N_44169,N_44093);
or U44262 (N_44262,N_44117,N_44021);
nand U44263 (N_44263,N_44096,N_44201);
or U44264 (N_44264,N_44202,N_44235);
nand U44265 (N_44265,N_44216,N_44236);
nor U44266 (N_44266,N_44206,N_44121);
xor U44267 (N_44267,N_44137,N_44223);
nor U44268 (N_44268,N_44039,N_44146);
and U44269 (N_44269,N_44155,N_44029);
nor U44270 (N_44270,N_44242,N_44176);
or U44271 (N_44271,N_44164,N_44220);
nor U44272 (N_44272,N_44006,N_44145);
xor U44273 (N_44273,N_44171,N_44204);
nor U44274 (N_44274,N_44081,N_44094);
nand U44275 (N_44275,N_44091,N_44027);
nor U44276 (N_44276,N_44234,N_44161);
xor U44277 (N_44277,N_44101,N_44073);
or U44278 (N_44278,N_44011,N_44240);
nand U44279 (N_44279,N_44126,N_44141);
xnor U44280 (N_44280,N_44009,N_44153);
xor U44281 (N_44281,N_44113,N_44030);
nor U44282 (N_44282,N_44135,N_44130);
and U44283 (N_44283,N_44023,N_44092);
nor U44284 (N_44284,N_44119,N_44087);
nand U44285 (N_44285,N_44187,N_44124);
xor U44286 (N_44286,N_44175,N_44185);
or U44287 (N_44287,N_44148,N_44042);
nand U44288 (N_44288,N_44076,N_44177);
or U44289 (N_44289,N_44154,N_44014);
and U44290 (N_44290,N_44125,N_44238);
or U44291 (N_44291,N_44064,N_44061);
nand U44292 (N_44292,N_44032,N_44035);
nor U44293 (N_44293,N_44019,N_44059);
xnor U44294 (N_44294,N_44150,N_44116);
xor U44295 (N_44295,N_44215,N_44008);
xor U44296 (N_44296,N_44170,N_44017);
and U44297 (N_44297,N_44003,N_44013);
or U44298 (N_44298,N_44162,N_44114);
xnor U44299 (N_44299,N_44034,N_44134);
nand U44300 (N_44300,N_44189,N_44036);
xor U44301 (N_44301,N_44111,N_44005);
and U44302 (N_44302,N_44247,N_44103);
nand U44303 (N_44303,N_44211,N_44195);
xnor U44304 (N_44304,N_44098,N_44115);
nor U44305 (N_44305,N_44004,N_44208);
or U44306 (N_44306,N_44192,N_44142);
or U44307 (N_44307,N_44075,N_44167);
nand U44308 (N_44308,N_44231,N_44173);
and U44309 (N_44309,N_44198,N_44024);
nor U44310 (N_44310,N_44178,N_44056);
nor U44311 (N_44311,N_44127,N_44156);
or U44312 (N_44312,N_44071,N_44160);
nand U44313 (N_44313,N_44168,N_44144);
and U44314 (N_44314,N_44131,N_44110);
nor U44315 (N_44315,N_44239,N_44214);
xnor U44316 (N_44316,N_44140,N_44107);
nor U44317 (N_44317,N_44199,N_44217);
nand U44318 (N_44318,N_44020,N_44197);
nand U44319 (N_44319,N_44243,N_44180);
nand U44320 (N_44320,N_44225,N_44190);
xor U44321 (N_44321,N_44191,N_44016);
or U44322 (N_44322,N_44222,N_44049);
nand U44323 (N_44323,N_44086,N_44249);
and U44324 (N_44324,N_44041,N_44200);
or U44325 (N_44325,N_44149,N_44139);
nand U44326 (N_44326,N_44143,N_44037);
nand U44327 (N_44327,N_44083,N_44147);
and U44328 (N_44328,N_44188,N_44015);
and U44329 (N_44329,N_44212,N_44072);
nor U44330 (N_44330,N_44053,N_44219);
and U44331 (N_44331,N_44052,N_44120);
and U44332 (N_44332,N_44078,N_44095);
xor U44333 (N_44333,N_44038,N_44179);
or U44334 (N_44334,N_44066,N_44057);
nand U44335 (N_44335,N_44163,N_44068);
or U44336 (N_44336,N_44050,N_44062);
or U44337 (N_44337,N_44207,N_44184);
nor U44338 (N_44338,N_44209,N_44074);
or U44339 (N_44339,N_44221,N_44122);
and U44340 (N_44340,N_44181,N_44194);
nor U44341 (N_44341,N_44226,N_44100);
and U44342 (N_44342,N_44099,N_44065);
nand U44343 (N_44343,N_44077,N_44069);
xor U44344 (N_44344,N_44007,N_44105);
xnor U44345 (N_44345,N_44132,N_44228);
or U44346 (N_44346,N_44193,N_44112);
nand U44347 (N_44347,N_44128,N_44205);
xnor U44348 (N_44348,N_44089,N_44248);
and U44349 (N_44349,N_44010,N_44186);
nor U44350 (N_44350,N_44046,N_44060);
nor U44351 (N_44351,N_44088,N_44183);
or U44352 (N_44352,N_44097,N_44210);
and U44353 (N_44353,N_44109,N_44227);
or U44354 (N_44354,N_44084,N_44033);
and U44355 (N_44355,N_44026,N_44218);
xor U44356 (N_44356,N_44151,N_44080);
xor U44357 (N_44357,N_44123,N_44055);
nor U44358 (N_44358,N_44040,N_44067);
nor U44359 (N_44359,N_44045,N_44063);
nand U44360 (N_44360,N_44174,N_44044);
nor U44361 (N_44361,N_44233,N_44246);
nand U44362 (N_44362,N_44047,N_44012);
or U44363 (N_44363,N_44018,N_44051);
and U44364 (N_44364,N_44138,N_44090);
xnor U44365 (N_44365,N_44025,N_44182);
and U44366 (N_44366,N_44237,N_44129);
or U44367 (N_44367,N_44152,N_44002);
xnor U44368 (N_44368,N_44102,N_44028);
nor U44369 (N_44369,N_44054,N_44224);
nor U44370 (N_44370,N_44082,N_44058);
or U44371 (N_44371,N_44196,N_44133);
and U44372 (N_44372,N_44108,N_44232);
and U44373 (N_44373,N_44244,N_44165);
xor U44374 (N_44374,N_44079,N_44245);
nand U44375 (N_44375,N_44050,N_44055);
nor U44376 (N_44376,N_44187,N_44097);
nor U44377 (N_44377,N_44173,N_44051);
xor U44378 (N_44378,N_44126,N_44104);
xnor U44379 (N_44379,N_44194,N_44226);
nor U44380 (N_44380,N_44051,N_44125);
nand U44381 (N_44381,N_44040,N_44183);
or U44382 (N_44382,N_44210,N_44100);
or U44383 (N_44383,N_44232,N_44163);
xor U44384 (N_44384,N_44058,N_44028);
or U44385 (N_44385,N_44046,N_44094);
xor U44386 (N_44386,N_44212,N_44115);
xor U44387 (N_44387,N_44172,N_44022);
or U44388 (N_44388,N_44046,N_44176);
and U44389 (N_44389,N_44145,N_44061);
xnor U44390 (N_44390,N_44193,N_44002);
nand U44391 (N_44391,N_44072,N_44228);
nor U44392 (N_44392,N_44112,N_44084);
nor U44393 (N_44393,N_44035,N_44069);
nor U44394 (N_44394,N_44157,N_44067);
nand U44395 (N_44395,N_44217,N_44015);
or U44396 (N_44396,N_44099,N_44217);
nor U44397 (N_44397,N_44130,N_44173);
and U44398 (N_44398,N_44245,N_44095);
nor U44399 (N_44399,N_44178,N_44146);
or U44400 (N_44400,N_44141,N_44199);
nand U44401 (N_44401,N_44035,N_44023);
nor U44402 (N_44402,N_44153,N_44045);
nor U44403 (N_44403,N_44071,N_44222);
or U44404 (N_44404,N_44023,N_44008);
and U44405 (N_44405,N_44239,N_44111);
xnor U44406 (N_44406,N_44065,N_44061);
xnor U44407 (N_44407,N_44023,N_44209);
nor U44408 (N_44408,N_44153,N_44232);
nand U44409 (N_44409,N_44206,N_44150);
xor U44410 (N_44410,N_44064,N_44214);
and U44411 (N_44411,N_44050,N_44153);
or U44412 (N_44412,N_44056,N_44117);
nor U44413 (N_44413,N_44219,N_44133);
or U44414 (N_44414,N_44140,N_44165);
xnor U44415 (N_44415,N_44157,N_44148);
nor U44416 (N_44416,N_44217,N_44237);
nor U44417 (N_44417,N_44062,N_44111);
nor U44418 (N_44418,N_44170,N_44003);
and U44419 (N_44419,N_44042,N_44133);
nor U44420 (N_44420,N_44195,N_44204);
xor U44421 (N_44421,N_44207,N_44139);
nor U44422 (N_44422,N_44152,N_44043);
nand U44423 (N_44423,N_44046,N_44138);
xnor U44424 (N_44424,N_44211,N_44085);
or U44425 (N_44425,N_44245,N_44205);
nor U44426 (N_44426,N_44016,N_44107);
nand U44427 (N_44427,N_44087,N_44140);
and U44428 (N_44428,N_44017,N_44192);
and U44429 (N_44429,N_44177,N_44214);
nor U44430 (N_44430,N_44131,N_44133);
or U44431 (N_44431,N_44186,N_44181);
nand U44432 (N_44432,N_44231,N_44210);
xnor U44433 (N_44433,N_44036,N_44041);
nor U44434 (N_44434,N_44047,N_44203);
nor U44435 (N_44435,N_44145,N_44219);
and U44436 (N_44436,N_44014,N_44024);
or U44437 (N_44437,N_44072,N_44168);
and U44438 (N_44438,N_44202,N_44241);
or U44439 (N_44439,N_44244,N_44015);
or U44440 (N_44440,N_44100,N_44206);
xnor U44441 (N_44441,N_44171,N_44212);
and U44442 (N_44442,N_44085,N_44205);
nand U44443 (N_44443,N_44076,N_44005);
nor U44444 (N_44444,N_44102,N_44046);
nor U44445 (N_44445,N_44118,N_44063);
and U44446 (N_44446,N_44021,N_44191);
nand U44447 (N_44447,N_44047,N_44181);
and U44448 (N_44448,N_44005,N_44027);
or U44449 (N_44449,N_44068,N_44135);
nand U44450 (N_44450,N_44068,N_44248);
xnor U44451 (N_44451,N_44210,N_44078);
and U44452 (N_44452,N_44128,N_44139);
and U44453 (N_44453,N_44170,N_44167);
nor U44454 (N_44454,N_44223,N_44034);
or U44455 (N_44455,N_44182,N_44094);
nor U44456 (N_44456,N_44171,N_44198);
and U44457 (N_44457,N_44244,N_44238);
and U44458 (N_44458,N_44229,N_44038);
or U44459 (N_44459,N_44021,N_44024);
nor U44460 (N_44460,N_44039,N_44059);
or U44461 (N_44461,N_44081,N_44114);
or U44462 (N_44462,N_44058,N_44038);
nand U44463 (N_44463,N_44212,N_44167);
and U44464 (N_44464,N_44171,N_44044);
and U44465 (N_44465,N_44016,N_44165);
or U44466 (N_44466,N_44046,N_44066);
and U44467 (N_44467,N_44011,N_44012);
nand U44468 (N_44468,N_44081,N_44095);
or U44469 (N_44469,N_44220,N_44035);
and U44470 (N_44470,N_44218,N_44233);
xor U44471 (N_44471,N_44221,N_44124);
and U44472 (N_44472,N_44030,N_44010);
or U44473 (N_44473,N_44101,N_44107);
nor U44474 (N_44474,N_44194,N_44115);
and U44475 (N_44475,N_44132,N_44063);
xor U44476 (N_44476,N_44120,N_44053);
nor U44477 (N_44477,N_44187,N_44056);
and U44478 (N_44478,N_44091,N_44141);
or U44479 (N_44479,N_44073,N_44085);
xnor U44480 (N_44480,N_44138,N_44027);
nand U44481 (N_44481,N_44231,N_44136);
xnor U44482 (N_44482,N_44111,N_44034);
xor U44483 (N_44483,N_44243,N_44068);
or U44484 (N_44484,N_44187,N_44158);
or U44485 (N_44485,N_44052,N_44057);
xor U44486 (N_44486,N_44158,N_44201);
nand U44487 (N_44487,N_44136,N_44089);
xor U44488 (N_44488,N_44072,N_44068);
and U44489 (N_44489,N_44026,N_44161);
and U44490 (N_44490,N_44148,N_44150);
and U44491 (N_44491,N_44226,N_44007);
or U44492 (N_44492,N_44026,N_44168);
nor U44493 (N_44493,N_44127,N_44191);
xor U44494 (N_44494,N_44068,N_44176);
or U44495 (N_44495,N_44225,N_44200);
nor U44496 (N_44496,N_44162,N_44150);
nand U44497 (N_44497,N_44172,N_44086);
and U44498 (N_44498,N_44073,N_44127);
nor U44499 (N_44499,N_44075,N_44162);
nor U44500 (N_44500,N_44313,N_44256);
xnor U44501 (N_44501,N_44371,N_44448);
or U44502 (N_44502,N_44403,N_44336);
and U44503 (N_44503,N_44299,N_44285);
nand U44504 (N_44504,N_44374,N_44386);
xnor U44505 (N_44505,N_44387,N_44320);
nand U44506 (N_44506,N_44291,N_44308);
nor U44507 (N_44507,N_44491,N_44485);
nor U44508 (N_44508,N_44353,N_44437);
nor U44509 (N_44509,N_44406,N_44344);
nand U44510 (N_44510,N_44267,N_44447);
nor U44511 (N_44511,N_44394,N_44358);
and U44512 (N_44512,N_44278,N_44276);
xor U44513 (N_44513,N_44427,N_44468);
or U44514 (N_44514,N_44296,N_44472);
nand U44515 (N_44515,N_44456,N_44328);
nand U44516 (N_44516,N_44304,N_44423);
nor U44517 (N_44517,N_44426,N_44262);
or U44518 (N_44518,N_44381,N_44463);
nand U44519 (N_44519,N_44316,N_44382);
nand U44520 (N_44520,N_44415,N_44473);
nand U44521 (N_44521,N_44300,N_44494);
nor U44522 (N_44522,N_44481,N_44274);
or U44523 (N_44523,N_44462,N_44496);
nor U44524 (N_44524,N_44337,N_44297);
nand U44525 (N_44525,N_44453,N_44409);
xnor U44526 (N_44526,N_44432,N_44351);
nor U44527 (N_44527,N_44323,N_44352);
nor U44528 (N_44528,N_44376,N_44330);
nor U44529 (N_44529,N_44250,N_44377);
nand U44530 (N_44530,N_44417,N_44321);
nand U44531 (N_44531,N_44272,N_44478);
and U44532 (N_44532,N_44343,N_44266);
nand U44533 (N_44533,N_44441,N_44332);
xnor U44534 (N_44534,N_44399,N_44388);
nor U44535 (N_44535,N_44268,N_44355);
and U44536 (N_44536,N_44383,N_44412);
nand U44537 (N_44537,N_44322,N_44293);
xnor U44538 (N_44538,N_44260,N_44338);
nor U44539 (N_44539,N_44324,N_44252);
and U44540 (N_44540,N_44364,N_44436);
or U44541 (N_44541,N_44442,N_44366);
or U44542 (N_44542,N_44348,N_44258);
nor U44543 (N_44543,N_44269,N_44424);
and U44544 (N_44544,N_44411,N_44356);
or U44545 (N_44545,N_44452,N_44284);
or U44546 (N_44546,N_44295,N_44370);
xor U44547 (N_44547,N_44360,N_44404);
nor U44548 (N_44548,N_44407,N_44421);
nor U44549 (N_44549,N_44326,N_44401);
or U44550 (N_44550,N_44280,N_44471);
or U44551 (N_44551,N_44487,N_44331);
or U44552 (N_44552,N_44385,N_44484);
and U44553 (N_44553,N_44464,N_44251);
nor U44554 (N_44554,N_44342,N_44265);
and U44555 (N_44555,N_44290,N_44283);
or U44556 (N_44556,N_44460,N_44334);
nand U44557 (N_44557,N_44480,N_44439);
nor U44558 (N_44558,N_44461,N_44349);
nor U44559 (N_44559,N_44271,N_44482);
or U44560 (N_44560,N_44368,N_44493);
and U44561 (N_44561,N_44372,N_44489);
and U44562 (N_44562,N_44444,N_44302);
xnor U44563 (N_44563,N_44305,N_44257);
nand U44564 (N_44564,N_44475,N_44490);
xnor U44565 (N_44565,N_44255,N_44354);
or U44566 (N_44566,N_44390,N_44379);
or U44567 (N_44567,N_44314,N_44365);
or U44568 (N_44568,N_44497,N_44483);
nor U44569 (N_44569,N_44346,N_44395);
and U44570 (N_44570,N_44286,N_44428);
nand U44571 (N_44571,N_44451,N_44359);
nand U44572 (N_44572,N_44422,N_44357);
and U44573 (N_44573,N_44378,N_44495);
nor U44574 (N_44574,N_44420,N_44341);
xnor U44575 (N_44575,N_44446,N_44329);
nand U44576 (N_44576,N_44413,N_44339);
and U44577 (N_44577,N_44288,N_44465);
and U44578 (N_44578,N_44315,N_44384);
nand U44579 (N_44579,N_44367,N_44392);
nor U44580 (N_44580,N_44333,N_44369);
or U44581 (N_44581,N_44431,N_44325);
and U44582 (N_44582,N_44393,N_44294);
nand U44583 (N_44583,N_44459,N_44309);
nor U44584 (N_44584,N_44479,N_44474);
xor U44585 (N_44585,N_44466,N_44312);
and U44586 (N_44586,N_44467,N_44317);
or U44587 (N_44587,N_44318,N_44301);
or U44588 (N_44588,N_44273,N_44263);
and U44589 (N_44589,N_44414,N_44270);
nor U44590 (N_44590,N_44476,N_44259);
and U44591 (N_44591,N_44405,N_44418);
nand U44592 (N_44592,N_44430,N_44375);
nor U44593 (N_44593,N_44327,N_44498);
nor U44594 (N_44594,N_44350,N_44373);
or U44595 (N_44595,N_44402,N_44279);
or U44596 (N_44596,N_44287,N_44298);
nor U44597 (N_44597,N_44454,N_44281);
and U44598 (N_44598,N_44362,N_44419);
nor U44599 (N_44599,N_44282,N_44492);
and U44600 (N_44600,N_44398,N_44455);
or U44601 (N_44601,N_44261,N_44380);
or U44602 (N_44602,N_44307,N_44400);
or U44603 (N_44603,N_44486,N_44335);
nor U44604 (N_44604,N_44397,N_44303);
nand U44605 (N_44605,N_44429,N_44319);
nand U44606 (N_44606,N_44275,N_44340);
and U44607 (N_44607,N_44306,N_44408);
nand U44608 (N_44608,N_44443,N_44396);
nor U44609 (N_44609,N_44450,N_44347);
or U44610 (N_44610,N_44345,N_44445);
or U44611 (N_44611,N_44391,N_44361);
or U44612 (N_44612,N_44310,N_44253);
nor U44613 (N_44613,N_44477,N_44311);
xor U44614 (N_44614,N_44438,N_44289);
or U44615 (N_44615,N_44458,N_44277);
and U44616 (N_44616,N_44292,N_44457);
and U44617 (N_44617,N_44440,N_44363);
or U44618 (N_44618,N_44449,N_44434);
and U44619 (N_44619,N_44470,N_44410);
or U44620 (N_44620,N_44254,N_44469);
nor U44621 (N_44621,N_44499,N_44433);
or U44622 (N_44622,N_44488,N_44435);
nor U44623 (N_44623,N_44416,N_44264);
nand U44624 (N_44624,N_44389,N_44425);
or U44625 (N_44625,N_44424,N_44494);
and U44626 (N_44626,N_44303,N_44295);
and U44627 (N_44627,N_44290,N_44356);
or U44628 (N_44628,N_44312,N_44468);
and U44629 (N_44629,N_44260,N_44489);
nand U44630 (N_44630,N_44270,N_44302);
nor U44631 (N_44631,N_44362,N_44436);
or U44632 (N_44632,N_44379,N_44407);
and U44633 (N_44633,N_44292,N_44484);
or U44634 (N_44634,N_44363,N_44281);
or U44635 (N_44635,N_44357,N_44311);
and U44636 (N_44636,N_44315,N_44458);
nor U44637 (N_44637,N_44446,N_44429);
and U44638 (N_44638,N_44374,N_44482);
and U44639 (N_44639,N_44376,N_44279);
or U44640 (N_44640,N_44432,N_44325);
xnor U44641 (N_44641,N_44467,N_44267);
nand U44642 (N_44642,N_44389,N_44300);
and U44643 (N_44643,N_44324,N_44463);
nand U44644 (N_44644,N_44451,N_44408);
nor U44645 (N_44645,N_44474,N_44397);
xor U44646 (N_44646,N_44276,N_44454);
nand U44647 (N_44647,N_44367,N_44493);
or U44648 (N_44648,N_44493,N_44331);
or U44649 (N_44649,N_44252,N_44361);
nand U44650 (N_44650,N_44417,N_44428);
and U44651 (N_44651,N_44470,N_44370);
xnor U44652 (N_44652,N_44337,N_44394);
xor U44653 (N_44653,N_44477,N_44476);
or U44654 (N_44654,N_44397,N_44345);
or U44655 (N_44655,N_44278,N_44404);
nor U44656 (N_44656,N_44480,N_44484);
nor U44657 (N_44657,N_44273,N_44306);
nand U44658 (N_44658,N_44312,N_44321);
or U44659 (N_44659,N_44328,N_44465);
nand U44660 (N_44660,N_44490,N_44419);
and U44661 (N_44661,N_44454,N_44437);
nor U44662 (N_44662,N_44443,N_44352);
nand U44663 (N_44663,N_44273,N_44433);
nor U44664 (N_44664,N_44354,N_44413);
nor U44665 (N_44665,N_44388,N_44442);
or U44666 (N_44666,N_44397,N_44263);
nor U44667 (N_44667,N_44497,N_44347);
and U44668 (N_44668,N_44297,N_44316);
xnor U44669 (N_44669,N_44279,N_44396);
nand U44670 (N_44670,N_44414,N_44292);
nor U44671 (N_44671,N_44334,N_44383);
nand U44672 (N_44672,N_44313,N_44464);
or U44673 (N_44673,N_44263,N_44480);
nor U44674 (N_44674,N_44413,N_44369);
xnor U44675 (N_44675,N_44480,N_44282);
nand U44676 (N_44676,N_44431,N_44363);
nand U44677 (N_44677,N_44262,N_44464);
and U44678 (N_44678,N_44253,N_44367);
nor U44679 (N_44679,N_44255,N_44264);
nand U44680 (N_44680,N_44318,N_44270);
nand U44681 (N_44681,N_44312,N_44270);
or U44682 (N_44682,N_44387,N_44351);
xnor U44683 (N_44683,N_44319,N_44461);
or U44684 (N_44684,N_44484,N_44375);
xnor U44685 (N_44685,N_44422,N_44254);
and U44686 (N_44686,N_44325,N_44439);
nand U44687 (N_44687,N_44347,N_44484);
xor U44688 (N_44688,N_44411,N_44382);
and U44689 (N_44689,N_44270,N_44258);
xor U44690 (N_44690,N_44320,N_44375);
and U44691 (N_44691,N_44380,N_44384);
or U44692 (N_44692,N_44451,N_44491);
nor U44693 (N_44693,N_44319,N_44406);
xnor U44694 (N_44694,N_44496,N_44254);
xnor U44695 (N_44695,N_44443,N_44259);
or U44696 (N_44696,N_44379,N_44423);
xnor U44697 (N_44697,N_44484,N_44267);
or U44698 (N_44698,N_44429,N_44397);
xnor U44699 (N_44699,N_44400,N_44262);
or U44700 (N_44700,N_44492,N_44496);
nand U44701 (N_44701,N_44322,N_44487);
nor U44702 (N_44702,N_44433,N_44256);
nor U44703 (N_44703,N_44277,N_44262);
xnor U44704 (N_44704,N_44280,N_44475);
or U44705 (N_44705,N_44320,N_44346);
or U44706 (N_44706,N_44444,N_44473);
and U44707 (N_44707,N_44372,N_44282);
and U44708 (N_44708,N_44256,N_44332);
nand U44709 (N_44709,N_44417,N_44397);
xor U44710 (N_44710,N_44490,N_44496);
xnor U44711 (N_44711,N_44467,N_44336);
and U44712 (N_44712,N_44495,N_44380);
xnor U44713 (N_44713,N_44341,N_44360);
nor U44714 (N_44714,N_44336,N_44255);
nor U44715 (N_44715,N_44321,N_44440);
and U44716 (N_44716,N_44372,N_44429);
xnor U44717 (N_44717,N_44318,N_44350);
and U44718 (N_44718,N_44294,N_44420);
xnor U44719 (N_44719,N_44396,N_44310);
and U44720 (N_44720,N_44383,N_44347);
and U44721 (N_44721,N_44341,N_44343);
xnor U44722 (N_44722,N_44273,N_44435);
nand U44723 (N_44723,N_44477,N_44384);
xnor U44724 (N_44724,N_44354,N_44311);
xnor U44725 (N_44725,N_44404,N_44460);
or U44726 (N_44726,N_44450,N_44437);
or U44727 (N_44727,N_44444,N_44330);
xor U44728 (N_44728,N_44371,N_44314);
xor U44729 (N_44729,N_44436,N_44482);
or U44730 (N_44730,N_44349,N_44393);
and U44731 (N_44731,N_44458,N_44253);
or U44732 (N_44732,N_44286,N_44330);
nor U44733 (N_44733,N_44354,N_44397);
xor U44734 (N_44734,N_44379,N_44408);
xor U44735 (N_44735,N_44489,N_44270);
nand U44736 (N_44736,N_44372,N_44365);
nor U44737 (N_44737,N_44332,N_44470);
nor U44738 (N_44738,N_44446,N_44254);
xor U44739 (N_44739,N_44254,N_44324);
or U44740 (N_44740,N_44262,N_44415);
xor U44741 (N_44741,N_44347,N_44264);
nand U44742 (N_44742,N_44281,N_44441);
xnor U44743 (N_44743,N_44448,N_44460);
nand U44744 (N_44744,N_44399,N_44486);
or U44745 (N_44745,N_44357,N_44271);
or U44746 (N_44746,N_44399,N_44373);
and U44747 (N_44747,N_44292,N_44458);
nand U44748 (N_44748,N_44340,N_44312);
nand U44749 (N_44749,N_44333,N_44345);
nor U44750 (N_44750,N_44636,N_44508);
or U44751 (N_44751,N_44551,N_44665);
xnor U44752 (N_44752,N_44727,N_44711);
and U44753 (N_44753,N_44748,N_44658);
and U44754 (N_44754,N_44734,N_44697);
xor U44755 (N_44755,N_44714,N_44504);
xnor U44756 (N_44756,N_44547,N_44688);
xnor U44757 (N_44757,N_44732,N_44634);
nand U44758 (N_44758,N_44605,N_44707);
nand U44759 (N_44759,N_44570,N_44703);
nand U44760 (N_44760,N_44720,N_44516);
nor U44761 (N_44761,N_44611,N_44723);
nor U44762 (N_44762,N_44626,N_44582);
nor U44763 (N_44763,N_44594,N_44555);
nand U44764 (N_44764,N_44619,N_44671);
and U44765 (N_44765,N_44562,N_44637);
nor U44766 (N_44766,N_44689,N_44678);
or U44767 (N_44767,N_44602,N_44685);
xor U44768 (N_44768,N_44642,N_44625);
nor U44769 (N_44769,N_44735,N_44531);
and U44770 (N_44770,N_44561,N_44725);
and U44771 (N_44771,N_44526,N_44583);
and U44772 (N_44772,N_44541,N_44532);
and U44773 (N_44773,N_44533,N_44606);
nor U44774 (N_44774,N_44747,N_44717);
nor U44775 (N_44775,N_44715,N_44627);
xor U44776 (N_44776,N_44586,N_44608);
xor U44777 (N_44777,N_44505,N_44670);
or U44778 (N_44778,N_44668,N_44742);
and U44779 (N_44779,N_44568,N_44639);
nor U44780 (N_44780,N_44730,N_44556);
nor U44781 (N_44781,N_44716,N_44679);
nand U44782 (N_44782,N_44593,N_44614);
xnor U44783 (N_44783,N_44745,N_44540);
and U44784 (N_44784,N_44530,N_44575);
xnor U44785 (N_44785,N_44534,N_44560);
or U44786 (N_44786,N_44584,N_44643);
xnor U44787 (N_44787,N_44631,N_44513);
and U44788 (N_44788,N_44522,N_44527);
xor U44789 (N_44789,N_44511,N_44749);
nor U44790 (N_44790,N_44552,N_44563);
nand U44791 (N_44791,N_44687,N_44672);
and U44792 (N_44792,N_44739,N_44537);
xnor U44793 (N_44793,N_44663,N_44623);
nor U44794 (N_44794,N_44694,N_44598);
nor U44795 (N_44795,N_44573,N_44553);
nor U44796 (N_44796,N_44655,N_44743);
nand U44797 (N_44797,N_44656,N_44550);
xnor U44798 (N_44798,N_44510,N_44645);
xor U44799 (N_44799,N_44708,N_44684);
nand U44800 (N_44800,N_44673,N_44740);
nand U44801 (N_44801,N_44613,N_44503);
or U44802 (N_44802,N_44710,N_44667);
xor U44803 (N_44803,N_44520,N_44559);
or U44804 (N_44804,N_44622,N_44744);
or U44805 (N_44805,N_44557,N_44579);
and U44806 (N_44806,N_44741,N_44603);
or U44807 (N_44807,N_44549,N_44691);
xor U44808 (N_44808,N_44698,N_44506);
xnor U44809 (N_44809,N_44539,N_44523);
nor U44810 (N_44810,N_44578,N_44628);
and U44811 (N_44811,N_44538,N_44746);
and U44812 (N_44812,N_44607,N_44693);
xnor U44813 (N_44813,N_44692,N_44659);
nor U44814 (N_44814,N_44542,N_44721);
nor U44815 (N_44815,N_44638,N_44501);
and U44816 (N_44816,N_44737,N_44621);
xnor U44817 (N_44817,N_44565,N_44669);
and U44818 (N_44818,N_44596,N_44515);
and U44819 (N_44819,N_44731,N_44564);
or U44820 (N_44820,N_44571,N_44652);
nor U44821 (N_44821,N_44618,N_44657);
xnor U44822 (N_44822,N_44728,N_44686);
or U44823 (N_44823,N_44680,N_44690);
nor U44824 (N_44824,N_44558,N_44644);
nor U44825 (N_44825,N_44640,N_44566);
xor U44826 (N_44826,N_44543,N_44632);
nand U44827 (N_44827,N_44509,N_44733);
nor U44828 (N_44828,N_44514,N_44529);
nand U44829 (N_44829,N_44507,N_44599);
xnor U44830 (N_44830,N_44600,N_44719);
nor U44831 (N_44831,N_44718,N_44545);
or U44832 (N_44832,N_44726,N_44554);
xor U44833 (N_44833,N_44674,N_44683);
or U44834 (N_44834,N_44612,N_44661);
xnor U44835 (N_44835,N_44700,N_44620);
nand U44836 (N_44836,N_44701,N_44589);
nor U44837 (N_44837,N_44724,N_44712);
and U44838 (N_44838,N_44648,N_44597);
nor U44839 (N_44839,N_44702,N_44569);
or U44840 (N_44840,N_44524,N_44604);
or U44841 (N_44841,N_44706,N_44588);
or U44842 (N_44842,N_44546,N_44601);
nand U44843 (N_44843,N_44544,N_44617);
or U44844 (N_44844,N_44709,N_44535);
and U44845 (N_44845,N_44677,N_44654);
nand U44846 (N_44846,N_44641,N_44675);
xnor U44847 (N_44847,N_44681,N_44660);
nand U44848 (N_44848,N_44525,N_44517);
or U44849 (N_44849,N_44528,N_44649);
xor U44850 (N_44850,N_44647,N_44592);
nor U44851 (N_44851,N_44630,N_44574);
or U44852 (N_44852,N_44572,N_44666);
and U44853 (N_44853,N_44738,N_44610);
or U44854 (N_44854,N_44653,N_44502);
and U44855 (N_44855,N_44664,N_44696);
and U44856 (N_44856,N_44587,N_44595);
and U44857 (N_44857,N_44576,N_44695);
xnor U44858 (N_44858,N_44624,N_44650);
nand U44859 (N_44859,N_44577,N_44646);
or U44860 (N_44860,N_44635,N_44722);
nand U44861 (N_44861,N_44609,N_44633);
xnor U44862 (N_44862,N_44591,N_44651);
nor U44863 (N_44863,N_44682,N_44662);
xnor U44864 (N_44864,N_44512,N_44699);
xnor U44865 (N_44865,N_44705,N_44616);
nor U44866 (N_44866,N_44704,N_44676);
nand U44867 (N_44867,N_44585,N_44519);
xnor U44868 (N_44868,N_44500,N_44567);
nand U44869 (N_44869,N_44521,N_44629);
or U44870 (N_44870,N_44590,N_44713);
nand U44871 (N_44871,N_44729,N_44615);
nand U44872 (N_44872,N_44518,N_44736);
xnor U44873 (N_44873,N_44548,N_44580);
nand U44874 (N_44874,N_44536,N_44581);
nor U44875 (N_44875,N_44619,N_44745);
or U44876 (N_44876,N_44574,N_44546);
xor U44877 (N_44877,N_44638,N_44687);
nand U44878 (N_44878,N_44728,N_44500);
nand U44879 (N_44879,N_44725,N_44706);
or U44880 (N_44880,N_44616,N_44532);
nor U44881 (N_44881,N_44685,N_44601);
or U44882 (N_44882,N_44690,N_44616);
xnor U44883 (N_44883,N_44685,N_44616);
or U44884 (N_44884,N_44640,N_44591);
or U44885 (N_44885,N_44558,N_44571);
xnor U44886 (N_44886,N_44629,N_44724);
or U44887 (N_44887,N_44594,N_44727);
nand U44888 (N_44888,N_44584,N_44542);
xnor U44889 (N_44889,N_44710,N_44542);
and U44890 (N_44890,N_44558,N_44541);
nor U44891 (N_44891,N_44684,N_44623);
nand U44892 (N_44892,N_44627,N_44686);
nand U44893 (N_44893,N_44606,N_44508);
xnor U44894 (N_44894,N_44544,N_44572);
xnor U44895 (N_44895,N_44710,N_44609);
or U44896 (N_44896,N_44539,N_44660);
nand U44897 (N_44897,N_44688,N_44674);
and U44898 (N_44898,N_44534,N_44638);
or U44899 (N_44899,N_44745,N_44515);
nor U44900 (N_44900,N_44515,N_44651);
xnor U44901 (N_44901,N_44674,N_44573);
nand U44902 (N_44902,N_44706,N_44641);
nand U44903 (N_44903,N_44642,N_44629);
or U44904 (N_44904,N_44741,N_44666);
xor U44905 (N_44905,N_44642,N_44682);
or U44906 (N_44906,N_44674,N_44511);
nor U44907 (N_44907,N_44645,N_44527);
or U44908 (N_44908,N_44619,N_44746);
and U44909 (N_44909,N_44564,N_44607);
xor U44910 (N_44910,N_44732,N_44747);
or U44911 (N_44911,N_44707,N_44577);
or U44912 (N_44912,N_44623,N_44665);
nor U44913 (N_44913,N_44636,N_44745);
and U44914 (N_44914,N_44513,N_44733);
xnor U44915 (N_44915,N_44712,N_44644);
or U44916 (N_44916,N_44619,N_44638);
or U44917 (N_44917,N_44672,N_44686);
and U44918 (N_44918,N_44546,N_44560);
xnor U44919 (N_44919,N_44654,N_44556);
nor U44920 (N_44920,N_44634,N_44560);
and U44921 (N_44921,N_44671,N_44580);
xor U44922 (N_44922,N_44700,N_44526);
xor U44923 (N_44923,N_44576,N_44590);
xor U44924 (N_44924,N_44612,N_44540);
nor U44925 (N_44925,N_44660,N_44513);
nand U44926 (N_44926,N_44547,N_44662);
xor U44927 (N_44927,N_44595,N_44652);
nand U44928 (N_44928,N_44603,N_44629);
nand U44929 (N_44929,N_44609,N_44612);
or U44930 (N_44930,N_44708,N_44517);
or U44931 (N_44931,N_44697,N_44596);
xnor U44932 (N_44932,N_44552,N_44583);
nor U44933 (N_44933,N_44506,N_44592);
and U44934 (N_44934,N_44643,N_44541);
nand U44935 (N_44935,N_44649,N_44612);
nor U44936 (N_44936,N_44574,N_44745);
and U44937 (N_44937,N_44727,N_44613);
and U44938 (N_44938,N_44662,N_44572);
nor U44939 (N_44939,N_44692,N_44701);
nor U44940 (N_44940,N_44572,N_44686);
xor U44941 (N_44941,N_44702,N_44611);
or U44942 (N_44942,N_44544,N_44629);
or U44943 (N_44943,N_44642,N_44557);
nand U44944 (N_44944,N_44578,N_44584);
nor U44945 (N_44945,N_44603,N_44544);
and U44946 (N_44946,N_44600,N_44727);
nand U44947 (N_44947,N_44512,N_44516);
xnor U44948 (N_44948,N_44718,N_44692);
nand U44949 (N_44949,N_44548,N_44591);
nand U44950 (N_44950,N_44583,N_44573);
nand U44951 (N_44951,N_44740,N_44627);
and U44952 (N_44952,N_44737,N_44660);
or U44953 (N_44953,N_44592,N_44692);
or U44954 (N_44954,N_44746,N_44669);
nand U44955 (N_44955,N_44678,N_44609);
or U44956 (N_44956,N_44653,N_44567);
nand U44957 (N_44957,N_44736,N_44521);
and U44958 (N_44958,N_44560,N_44734);
and U44959 (N_44959,N_44740,N_44593);
and U44960 (N_44960,N_44710,N_44715);
xor U44961 (N_44961,N_44707,N_44579);
or U44962 (N_44962,N_44740,N_44618);
nand U44963 (N_44963,N_44665,N_44611);
nand U44964 (N_44964,N_44570,N_44542);
nor U44965 (N_44965,N_44545,N_44634);
nor U44966 (N_44966,N_44689,N_44603);
and U44967 (N_44967,N_44626,N_44635);
xnor U44968 (N_44968,N_44515,N_44584);
nand U44969 (N_44969,N_44652,N_44515);
xnor U44970 (N_44970,N_44555,N_44619);
nand U44971 (N_44971,N_44703,N_44629);
and U44972 (N_44972,N_44739,N_44728);
and U44973 (N_44973,N_44641,N_44582);
xnor U44974 (N_44974,N_44702,N_44517);
or U44975 (N_44975,N_44641,N_44536);
nand U44976 (N_44976,N_44699,N_44655);
or U44977 (N_44977,N_44688,N_44516);
or U44978 (N_44978,N_44719,N_44525);
and U44979 (N_44979,N_44609,N_44665);
and U44980 (N_44980,N_44674,N_44547);
and U44981 (N_44981,N_44641,N_44632);
nor U44982 (N_44982,N_44588,N_44512);
nand U44983 (N_44983,N_44573,N_44640);
and U44984 (N_44984,N_44650,N_44647);
or U44985 (N_44985,N_44636,N_44732);
nor U44986 (N_44986,N_44578,N_44718);
nand U44987 (N_44987,N_44639,N_44746);
and U44988 (N_44988,N_44715,N_44522);
or U44989 (N_44989,N_44748,N_44592);
nand U44990 (N_44990,N_44747,N_44635);
nand U44991 (N_44991,N_44541,N_44606);
and U44992 (N_44992,N_44739,N_44686);
nor U44993 (N_44993,N_44547,N_44513);
xnor U44994 (N_44994,N_44698,N_44747);
nand U44995 (N_44995,N_44547,N_44668);
and U44996 (N_44996,N_44560,N_44638);
or U44997 (N_44997,N_44655,N_44559);
or U44998 (N_44998,N_44520,N_44665);
nand U44999 (N_44999,N_44743,N_44669);
xor U45000 (N_45000,N_44829,N_44965);
xnor U45001 (N_45001,N_44928,N_44915);
nor U45002 (N_45002,N_44853,N_44873);
nor U45003 (N_45003,N_44983,N_44843);
nand U45004 (N_45004,N_44909,N_44916);
or U45005 (N_45005,N_44845,N_44976);
and U45006 (N_45006,N_44929,N_44819);
and U45007 (N_45007,N_44778,N_44856);
or U45008 (N_45008,N_44939,N_44973);
xnor U45009 (N_45009,N_44805,N_44954);
or U45010 (N_45010,N_44995,N_44807);
xnor U45011 (N_45011,N_44774,N_44849);
nand U45012 (N_45012,N_44957,N_44885);
xor U45013 (N_45013,N_44759,N_44974);
nand U45014 (N_45014,N_44935,N_44964);
or U45015 (N_45015,N_44967,N_44989);
or U45016 (N_45016,N_44852,N_44832);
xnor U45017 (N_45017,N_44810,N_44861);
xor U45018 (N_45018,N_44945,N_44898);
xnor U45019 (N_45019,N_44806,N_44753);
nor U45020 (N_45020,N_44760,N_44893);
nand U45021 (N_45021,N_44814,N_44970);
nor U45022 (N_45022,N_44889,N_44796);
xor U45023 (N_45023,N_44775,N_44878);
xnor U45024 (N_45024,N_44791,N_44867);
xnor U45025 (N_45025,N_44801,N_44818);
nor U45026 (N_45026,N_44783,N_44999);
or U45027 (N_45027,N_44834,N_44812);
nand U45028 (N_45028,N_44897,N_44790);
nand U45029 (N_45029,N_44811,N_44798);
xnor U45030 (N_45030,N_44837,N_44895);
xnor U45031 (N_45031,N_44793,N_44952);
xnor U45032 (N_45032,N_44802,N_44971);
nand U45033 (N_45033,N_44771,N_44824);
nand U45034 (N_45034,N_44857,N_44998);
or U45035 (N_45035,N_44922,N_44933);
or U45036 (N_45036,N_44904,N_44926);
nor U45037 (N_45037,N_44982,N_44890);
and U45038 (N_45038,N_44772,N_44899);
xnor U45039 (N_45039,N_44993,N_44960);
nand U45040 (N_45040,N_44820,N_44984);
nand U45041 (N_45041,N_44881,N_44794);
and U45042 (N_45042,N_44887,N_44862);
xor U45043 (N_45043,N_44836,N_44827);
nor U45044 (N_45044,N_44882,N_44940);
xnor U45045 (N_45045,N_44879,N_44786);
nor U45046 (N_45046,N_44846,N_44813);
or U45047 (N_45047,N_44808,N_44868);
nand U45048 (N_45048,N_44880,N_44961);
nand U45049 (N_45049,N_44752,N_44988);
nor U45050 (N_45050,N_44951,N_44850);
nor U45051 (N_45051,N_44833,N_44949);
or U45052 (N_45052,N_44839,N_44870);
nand U45053 (N_45053,N_44944,N_44844);
xnor U45054 (N_45054,N_44785,N_44804);
xnor U45055 (N_45055,N_44918,N_44923);
or U45056 (N_45056,N_44886,N_44750);
nand U45057 (N_45057,N_44979,N_44779);
nor U45058 (N_45058,N_44787,N_44828);
nor U45059 (N_45059,N_44821,N_44866);
or U45060 (N_45060,N_44859,N_44831);
nand U45061 (N_45061,N_44883,N_44816);
and U45062 (N_45062,N_44770,N_44950);
or U45063 (N_45063,N_44826,N_44830);
nor U45064 (N_45064,N_44815,N_44797);
nor U45065 (N_45065,N_44756,N_44766);
and U45066 (N_45066,N_44872,N_44884);
xor U45067 (N_45067,N_44972,N_44925);
nand U45068 (N_45068,N_44931,N_44914);
and U45069 (N_45069,N_44764,N_44767);
or U45070 (N_45070,N_44768,N_44854);
nand U45071 (N_45071,N_44875,N_44910);
or U45072 (N_45072,N_44865,N_44847);
and U45073 (N_45073,N_44871,N_44876);
nand U45074 (N_45074,N_44955,N_44874);
or U45075 (N_45075,N_44919,N_44788);
nand U45076 (N_45076,N_44855,N_44763);
nor U45077 (N_45077,N_44994,N_44927);
nor U45078 (N_45078,N_44948,N_44959);
nor U45079 (N_45079,N_44858,N_44755);
nor U45080 (N_45080,N_44992,N_44968);
and U45081 (N_45081,N_44758,N_44913);
nor U45082 (N_45082,N_44977,N_44908);
and U45083 (N_45083,N_44990,N_44907);
nand U45084 (N_45084,N_44917,N_44838);
nor U45085 (N_45085,N_44891,N_44869);
nand U45086 (N_45086,N_44911,N_44892);
nand U45087 (N_45087,N_44920,N_44888);
or U45088 (N_45088,N_44841,N_44803);
and U45089 (N_45089,N_44963,N_44943);
nand U45090 (N_45090,N_44900,N_44937);
nand U45091 (N_45091,N_44978,N_44936);
nand U45092 (N_45092,N_44924,N_44981);
nor U45093 (N_45093,N_44905,N_44921);
nand U45094 (N_45094,N_44780,N_44942);
nand U45095 (N_45095,N_44860,N_44840);
nand U45096 (N_45096,N_44941,N_44902);
nor U45097 (N_45097,N_44762,N_44835);
nor U45098 (N_45098,N_44784,N_44894);
or U45099 (N_45099,N_44958,N_44906);
and U45100 (N_45100,N_44754,N_44903);
xnor U45101 (N_45101,N_44848,N_44825);
nand U45102 (N_45102,N_44896,N_44946);
nor U45103 (N_45103,N_44863,N_44817);
xnor U45104 (N_45104,N_44877,N_44966);
or U45105 (N_45105,N_44947,N_44956);
xnor U45106 (N_45106,N_44757,N_44792);
and U45107 (N_45107,N_44795,N_44776);
and U45108 (N_45108,N_44962,N_44842);
or U45109 (N_45109,N_44751,N_44938);
or U45110 (N_45110,N_44822,N_44997);
nor U45111 (N_45111,N_44901,N_44934);
nor U45112 (N_45112,N_44823,N_44987);
nor U45113 (N_45113,N_44782,N_44969);
and U45114 (N_45114,N_44789,N_44975);
xor U45115 (N_45115,N_44930,N_44851);
nand U45116 (N_45116,N_44800,N_44809);
nand U45117 (N_45117,N_44985,N_44761);
nand U45118 (N_45118,N_44986,N_44912);
nand U45119 (N_45119,N_44781,N_44953);
nor U45120 (N_45120,N_44765,N_44799);
xor U45121 (N_45121,N_44773,N_44777);
nand U45122 (N_45122,N_44991,N_44932);
xor U45123 (N_45123,N_44769,N_44864);
nor U45124 (N_45124,N_44980,N_44996);
nor U45125 (N_45125,N_44824,N_44925);
or U45126 (N_45126,N_44987,N_44766);
xor U45127 (N_45127,N_44870,N_44983);
and U45128 (N_45128,N_44945,N_44892);
and U45129 (N_45129,N_44997,N_44843);
xor U45130 (N_45130,N_44922,N_44924);
nor U45131 (N_45131,N_44781,N_44963);
and U45132 (N_45132,N_44799,N_44885);
or U45133 (N_45133,N_44852,N_44930);
and U45134 (N_45134,N_44820,N_44858);
or U45135 (N_45135,N_44807,N_44914);
or U45136 (N_45136,N_44789,N_44933);
or U45137 (N_45137,N_44819,N_44935);
xnor U45138 (N_45138,N_44990,N_44937);
nand U45139 (N_45139,N_44861,N_44956);
nand U45140 (N_45140,N_44812,N_44915);
and U45141 (N_45141,N_44808,N_44899);
or U45142 (N_45142,N_44849,N_44986);
nor U45143 (N_45143,N_44901,N_44859);
and U45144 (N_45144,N_44800,N_44949);
nor U45145 (N_45145,N_44952,N_44805);
and U45146 (N_45146,N_44931,N_44758);
or U45147 (N_45147,N_44772,N_44942);
xnor U45148 (N_45148,N_44893,N_44828);
nor U45149 (N_45149,N_44801,N_44797);
nor U45150 (N_45150,N_44916,N_44789);
nor U45151 (N_45151,N_44855,N_44760);
nor U45152 (N_45152,N_44904,N_44765);
or U45153 (N_45153,N_44784,N_44976);
nor U45154 (N_45154,N_44806,N_44892);
or U45155 (N_45155,N_44790,N_44775);
and U45156 (N_45156,N_44898,N_44913);
and U45157 (N_45157,N_44858,N_44948);
and U45158 (N_45158,N_44824,N_44762);
and U45159 (N_45159,N_44985,N_44884);
and U45160 (N_45160,N_44781,N_44810);
or U45161 (N_45161,N_44928,N_44789);
and U45162 (N_45162,N_44778,N_44933);
nor U45163 (N_45163,N_44971,N_44878);
and U45164 (N_45164,N_44844,N_44904);
xnor U45165 (N_45165,N_44897,N_44871);
xnor U45166 (N_45166,N_44952,N_44839);
nor U45167 (N_45167,N_44766,N_44764);
nand U45168 (N_45168,N_44758,N_44898);
nor U45169 (N_45169,N_44997,N_44804);
and U45170 (N_45170,N_44813,N_44893);
and U45171 (N_45171,N_44943,N_44985);
nor U45172 (N_45172,N_44818,N_44952);
or U45173 (N_45173,N_44766,N_44838);
or U45174 (N_45174,N_44954,N_44849);
nor U45175 (N_45175,N_44865,N_44830);
nand U45176 (N_45176,N_44882,N_44792);
nor U45177 (N_45177,N_44999,N_44883);
nand U45178 (N_45178,N_44929,N_44763);
nand U45179 (N_45179,N_44824,N_44914);
and U45180 (N_45180,N_44835,N_44975);
nand U45181 (N_45181,N_44988,N_44972);
nand U45182 (N_45182,N_44950,N_44841);
xnor U45183 (N_45183,N_44922,N_44887);
xor U45184 (N_45184,N_44945,N_44750);
and U45185 (N_45185,N_44897,N_44830);
nand U45186 (N_45186,N_44995,N_44896);
nor U45187 (N_45187,N_44982,N_44781);
or U45188 (N_45188,N_44967,N_44769);
or U45189 (N_45189,N_44808,N_44788);
xor U45190 (N_45190,N_44796,N_44876);
xor U45191 (N_45191,N_44912,N_44816);
xor U45192 (N_45192,N_44908,N_44928);
or U45193 (N_45193,N_44794,N_44863);
and U45194 (N_45194,N_44883,N_44978);
nor U45195 (N_45195,N_44809,N_44775);
nand U45196 (N_45196,N_44993,N_44995);
or U45197 (N_45197,N_44819,N_44860);
nand U45198 (N_45198,N_44969,N_44948);
xnor U45199 (N_45199,N_44979,N_44834);
and U45200 (N_45200,N_44956,N_44874);
or U45201 (N_45201,N_44990,N_44985);
or U45202 (N_45202,N_44834,N_44813);
xor U45203 (N_45203,N_44940,N_44947);
nor U45204 (N_45204,N_44882,N_44868);
nand U45205 (N_45205,N_44965,N_44952);
xor U45206 (N_45206,N_44839,N_44803);
and U45207 (N_45207,N_44781,N_44827);
and U45208 (N_45208,N_44934,N_44775);
and U45209 (N_45209,N_44852,N_44800);
nor U45210 (N_45210,N_44942,N_44881);
nor U45211 (N_45211,N_44917,N_44853);
and U45212 (N_45212,N_44962,N_44869);
xor U45213 (N_45213,N_44865,N_44961);
nand U45214 (N_45214,N_44909,N_44796);
nand U45215 (N_45215,N_44855,N_44756);
xnor U45216 (N_45216,N_44883,N_44841);
nand U45217 (N_45217,N_44867,N_44945);
and U45218 (N_45218,N_44761,N_44784);
xnor U45219 (N_45219,N_44880,N_44850);
and U45220 (N_45220,N_44949,N_44856);
xnor U45221 (N_45221,N_44916,N_44976);
nor U45222 (N_45222,N_44875,N_44960);
nand U45223 (N_45223,N_44893,N_44871);
and U45224 (N_45224,N_44849,N_44988);
xnor U45225 (N_45225,N_44989,N_44929);
nor U45226 (N_45226,N_44813,N_44958);
and U45227 (N_45227,N_44931,N_44843);
nand U45228 (N_45228,N_44864,N_44830);
xor U45229 (N_45229,N_44921,N_44788);
nor U45230 (N_45230,N_44976,N_44988);
and U45231 (N_45231,N_44847,N_44769);
or U45232 (N_45232,N_44812,N_44912);
nand U45233 (N_45233,N_44940,N_44913);
or U45234 (N_45234,N_44856,N_44971);
nor U45235 (N_45235,N_44766,N_44820);
and U45236 (N_45236,N_44805,N_44756);
nand U45237 (N_45237,N_44778,N_44945);
or U45238 (N_45238,N_44970,N_44804);
xor U45239 (N_45239,N_44887,N_44978);
xor U45240 (N_45240,N_44853,N_44805);
or U45241 (N_45241,N_44763,N_44948);
and U45242 (N_45242,N_44880,N_44930);
xnor U45243 (N_45243,N_44908,N_44886);
or U45244 (N_45244,N_44875,N_44950);
or U45245 (N_45245,N_44963,N_44858);
nor U45246 (N_45246,N_44757,N_44923);
nand U45247 (N_45247,N_44811,N_44806);
xor U45248 (N_45248,N_44784,N_44815);
nor U45249 (N_45249,N_44890,N_44796);
and U45250 (N_45250,N_45046,N_45023);
or U45251 (N_45251,N_45246,N_45004);
or U45252 (N_45252,N_45062,N_45170);
and U45253 (N_45253,N_45152,N_45154);
nand U45254 (N_45254,N_45191,N_45225);
nand U45255 (N_45255,N_45197,N_45002);
and U45256 (N_45256,N_45175,N_45146);
and U45257 (N_45257,N_45035,N_45166);
and U45258 (N_45258,N_45027,N_45034);
nand U45259 (N_45259,N_45235,N_45082);
and U45260 (N_45260,N_45015,N_45118);
xnor U45261 (N_45261,N_45212,N_45112);
nor U45262 (N_45262,N_45202,N_45053);
or U45263 (N_45263,N_45177,N_45243);
nor U45264 (N_45264,N_45092,N_45199);
xor U45265 (N_45265,N_45041,N_45215);
nor U45266 (N_45266,N_45066,N_45061);
or U45267 (N_45267,N_45237,N_45240);
xnor U45268 (N_45268,N_45007,N_45226);
nand U45269 (N_45269,N_45142,N_45052);
and U45270 (N_45270,N_45141,N_45228);
nand U45271 (N_45271,N_45130,N_45070);
nand U45272 (N_45272,N_45072,N_45245);
or U45273 (N_45273,N_45242,N_45137);
or U45274 (N_45274,N_45074,N_45234);
or U45275 (N_45275,N_45117,N_45075);
nand U45276 (N_45276,N_45220,N_45045);
and U45277 (N_45277,N_45151,N_45203);
xnor U45278 (N_45278,N_45022,N_45110);
or U45279 (N_45279,N_45050,N_45216);
or U45280 (N_45280,N_45176,N_45206);
nor U45281 (N_45281,N_45005,N_45194);
or U45282 (N_45282,N_45103,N_45223);
and U45283 (N_45283,N_45094,N_45087);
or U45284 (N_45284,N_45059,N_45196);
nor U45285 (N_45285,N_45148,N_45195);
and U45286 (N_45286,N_45078,N_45042);
or U45287 (N_45287,N_45143,N_45001);
nand U45288 (N_45288,N_45158,N_45201);
nor U45289 (N_45289,N_45133,N_45207);
nor U45290 (N_45290,N_45003,N_45162);
or U45291 (N_45291,N_45138,N_45069);
nor U45292 (N_45292,N_45222,N_45032);
and U45293 (N_45293,N_45014,N_45244);
xor U45294 (N_45294,N_45021,N_45127);
nand U45295 (N_45295,N_45164,N_45036);
nor U45296 (N_45296,N_45178,N_45033);
nand U45297 (N_45297,N_45150,N_45120);
nand U45298 (N_45298,N_45031,N_45081);
nor U45299 (N_45299,N_45239,N_45089);
or U45300 (N_45300,N_45219,N_45085);
and U45301 (N_45301,N_45205,N_45067);
nand U45302 (N_45302,N_45048,N_45038);
and U45303 (N_45303,N_45088,N_45128);
nand U45304 (N_45304,N_45065,N_45121);
and U45305 (N_45305,N_45132,N_45054);
nand U45306 (N_45306,N_45084,N_45165);
and U45307 (N_45307,N_45044,N_45096);
nor U45308 (N_45308,N_45119,N_45068);
xnor U45309 (N_45309,N_45080,N_45125);
or U45310 (N_45310,N_45188,N_45129);
and U45311 (N_45311,N_45083,N_45018);
nand U45312 (N_45312,N_45009,N_45167);
xor U45313 (N_45313,N_45111,N_45173);
and U45314 (N_45314,N_45140,N_45122);
or U45315 (N_45315,N_45079,N_45183);
and U45316 (N_45316,N_45247,N_45218);
xor U45317 (N_45317,N_45017,N_45076);
nand U45318 (N_45318,N_45236,N_45116);
or U45319 (N_45319,N_45221,N_45213);
or U45320 (N_45320,N_45229,N_45248);
xnor U45321 (N_45321,N_45123,N_45064);
nand U45322 (N_45322,N_45055,N_45232);
or U45323 (N_45323,N_45159,N_45093);
nand U45324 (N_45324,N_45171,N_45058);
xor U45325 (N_45325,N_45105,N_45131);
xnor U45326 (N_45326,N_45114,N_45006);
or U45327 (N_45327,N_45185,N_45107);
xnor U45328 (N_45328,N_45249,N_45180);
nor U45329 (N_45329,N_45214,N_45182);
and U45330 (N_45330,N_45156,N_45153);
nor U45331 (N_45331,N_45211,N_45099);
xnor U45332 (N_45332,N_45139,N_45012);
xor U45333 (N_45333,N_45101,N_45086);
nand U45334 (N_45334,N_45172,N_45060);
or U45335 (N_45335,N_45056,N_45174);
nor U45336 (N_45336,N_45169,N_45010);
and U45337 (N_45337,N_45043,N_45011);
and U45338 (N_45338,N_45208,N_45217);
and U45339 (N_45339,N_45097,N_45233);
xnor U45340 (N_45340,N_45073,N_45184);
xnor U45341 (N_45341,N_45230,N_45108);
nor U45342 (N_45342,N_45057,N_45135);
or U45343 (N_45343,N_45019,N_45095);
and U45344 (N_45344,N_45100,N_45030);
nand U45345 (N_45345,N_45238,N_45026);
and U45346 (N_45346,N_45077,N_45209);
or U45347 (N_45347,N_45040,N_45104);
xnor U45348 (N_45348,N_45024,N_45210);
xnor U45349 (N_45349,N_45227,N_45028);
xnor U45350 (N_45350,N_45186,N_45109);
nor U45351 (N_45351,N_45071,N_45193);
and U45352 (N_45352,N_45091,N_45047);
nand U45353 (N_45353,N_45204,N_45157);
xnor U45354 (N_45354,N_45020,N_45013);
nor U45355 (N_45355,N_45163,N_45147);
nor U45356 (N_45356,N_45025,N_45098);
nand U45357 (N_45357,N_45008,N_45190);
and U45358 (N_45358,N_45160,N_45063);
xor U45359 (N_45359,N_45029,N_45049);
or U45360 (N_45360,N_45168,N_45189);
nor U45361 (N_45361,N_45016,N_45181);
nand U45362 (N_45362,N_45134,N_45149);
nor U45363 (N_45363,N_45115,N_45161);
or U45364 (N_45364,N_45102,N_45126);
xnor U45365 (N_45365,N_45000,N_45241);
nand U45366 (N_45366,N_45179,N_45198);
xor U45367 (N_45367,N_45231,N_45144);
and U45368 (N_45368,N_45200,N_45106);
and U45369 (N_45369,N_45224,N_45051);
and U45370 (N_45370,N_45187,N_45136);
xor U45371 (N_45371,N_45113,N_45090);
nand U45372 (N_45372,N_45037,N_45124);
nand U45373 (N_45373,N_45145,N_45192);
nand U45374 (N_45374,N_45039,N_45155);
nand U45375 (N_45375,N_45027,N_45038);
or U45376 (N_45376,N_45011,N_45031);
nand U45377 (N_45377,N_45068,N_45177);
nor U45378 (N_45378,N_45082,N_45061);
nand U45379 (N_45379,N_45031,N_45216);
xnor U45380 (N_45380,N_45139,N_45107);
nor U45381 (N_45381,N_45145,N_45097);
or U45382 (N_45382,N_45071,N_45131);
nand U45383 (N_45383,N_45019,N_45030);
or U45384 (N_45384,N_45209,N_45041);
xor U45385 (N_45385,N_45238,N_45226);
or U45386 (N_45386,N_45062,N_45221);
or U45387 (N_45387,N_45098,N_45071);
xor U45388 (N_45388,N_45179,N_45199);
nor U45389 (N_45389,N_45141,N_45244);
or U45390 (N_45390,N_45108,N_45217);
and U45391 (N_45391,N_45091,N_45117);
and U45392 (N_45392,N_45210,N_45208);
and U45393 (N_45393,N_45007,N_45055);
nor U45394 (N_45394,N_45052,N_45198);
and U45395 (N_45395,N_45168,N_45064);
nor U45396 (N_45396,N_45202,N_45030);
nor U45397 (N_45397,N_45155,N_45216);
and U45398 (N_45398,N_45158,N_45087);
and U45399 (N_45399,N_45194,N_45098);
and U45400 (N_45400,N_45173,N_45102);
or U45401 (N_45401,N_45122,N_45085);
and U45402 (N_45402,N_45176,N_45116);
and U45403 (N_45403,N_45043,N_45130);
or U45404 (N_45404,N_45150,N_45182);
nor U45405 (N_45405,N_45178,N_45235);
or U45406 (N_45406,N_45198,N_45246);
or U45407 (N_45407,N_45119,N_45137);
or U45408 (N_45408,N_45114,N_45118);
xnor U45409 (N_45409,N_45193,N_45010);
nor U45410 (N_45410,N_45188,N_45089);
xor U45411 (N_45411,N_45046,N_45233);
nor U45412 (N_45412,N_45100,N_45064);
nor U45413 (N_45413,N_45054,N_45197);
nand U45414 (N_45414,N_45120,N_45052);
and U45415 (N_45415,N_45126,N_45011);
xor U45416 (N_45416,N_45234,N_45210);
and U45417 (N_45417,N_45141,N_45099);
nand U45418 (N_45418,N_45211,N_45068);
nor U45419 (N_45419,N_45161,N_45207);
and U45420 (N_45420,N_45061,N_45040);
xnor U45421 (N_45421,N_45084,N_45135);
or U45422 (N_45422,N_45182,N_45188);
nor U45423 (N_45423,N_45027,N_45168);
nor U45424 (N_45424,N_45122,N_45166);
nand U45425 (N_45425,N_45008,N_45191);
nor U45426 (N_45426,N_45124,N_45033);
nand U45427 (N_45427,N_45140,N_45036);
nand U45428 (N_45428,N_45116,N_45106);
nand U45429 (N_45429,N_45025,N_45226);
nor U45430 (N_45430,N_45157,N_45223);
nand U45431 (N_45431,N_45145,N_45246);
and U45432 (N_45432,N_45209,N_45174);
nor U45433 (N_45433,N_45104,N_45192);
nor U45434 (N_45434,N_45117,N_45174);
and U45435 (N_45435,N_45093,N_45180);
nor U45436 (N_45436,N_45174,N_45094);
xnor U45437 (N_45437,N_45166,N_45059);
nor U45438 (N_45438,N_45096,N_45224);
nand U45439 (N_45439,N_45127,N_45124);
and U45440 (N_45440,N_45127,N_45106);
or U45441 (N_45441,N_45187,N_45121);
nand U45442 (N_45442,N_45233,N_45112);
or U45443 (N_45443,N_45063,N_45134);
nor U45444 (N_45444,N_45210,N_45051);
xnor U45445 (N_45445,N_45209,N_45049);
nor U45446 (N_45446,N_45144,N_45062);
or U45447 (N_45447,N_45243,N_45049);
and U45448 (N_45448,N_45047,N_45194);
nand U45449 (N_45449,N_45146,N_45109);
xnor U45450 (N_45450,N_45189,N_45108);
xor U45451 (N_45451,N_45045,N_45071);
nand U45452 (N_45452,N_45173,N_45166);
and U45453 (N_45453,N_45021,N_45161);
nor U45454 (N_45454,N_45071,N_45052);
xnor U45455 (N_45455,N_45246,N_45056);
and U45456 (N_45456,N_45127,N_45175);
nand U45457 (N_45457,N_45024,N_45080);
nand U45458 (N_45458,N_45138,N_45115);
nand U45459 (N_45459,N_45015,N_45051);
and U45460 (N_45460,N_45096,N_45083);
and U45461 (N_45461,N_45159,N_45231);
nand U45462 (N_45462,N_45231,N_45052);
nor U45463 (N_45463,N_45085,N_45238);
xnor U45464 (N_45464,N_45112,N_45031);
nand U45465 (N_45465,N_45028,N_45134);
nand U45466 (N_45466,N_45037,N_45033);
xnor U45467 (N_45467,N_45189,N_45159);
xnor U45468 (N_45468,N_45145,N_45122);
xor U45469 (N_45469,N_45197,N_45232);
or U45470 (N_45470,N_45082,N_45223);
xor U45471 (N_45471,N_45055,N_45198);
or U45472 (N_45472,N_45173,N_45080);
nor U45473 (N_45473,N_45236,N_45201);
nor U45474 (N_45474,N_45241,N_45120);
nand U45475 (N_45475,N_45182,N_45185);
or U45476 (N_45476,N_45033,N_45214);
nand U45477 (N_45477,N_45206,N_45204);
and U45478 (N_45478,N_45208,N_45190);
nand U45479 (N_45479,N_45230,N_45121);
nor U45480 (N_45480,N_45219,N_45247);
or U45481 (N_45481,N_45153,N_45070);
nor U45482 (N_45482,N_45154,N_45047);
nand U45483 (N_45483,N_45166,N_45121);
and U45484 (N_45484,N_45061,N_45249);
nand U45485 (N_45485,N_45011,N_45069);
nand U45486 (N_45486,N_45201,N_45109);
and U45487 (N_45487,N_45082,N_45016);
and U45488 (N_45488,N_45213,N_45043);
nand U45489 (N_45489,N_45176,N_45010);
or U45490 (N_45490,N_45021,N_45037);
nor U45491 (N_45491,N_45205,N_45148);
nand U45492 (N_45492,N_45224,N_45065);
xnor U45493 (N_45493,N_45234,N_45100);
nand U45494 (N_45494,N_45110,N_45030);
and U45495 (N_45495,N_45234,N_45093);
nor U45496 (N_45496,N_45083,N_45144);
nor U45497 (N_45497,N_45177,N_45124);
or U45498 (N_45498,N_45100,N_45208);
nor U45499 (N_45499,N_45237,N_45069);
nand U45500 (N_45500,N_45485,N_45399);
nand U45501 (N_45501,N_45374,N_45397);
or U45502 (N_45502,N_45305,N_45487);
and U45503 (N_45503,N_45271,N_45379);
nand U45504 (N_45504,N_45347,N_45328);
nor U45505 (N_45505,N_45279,N_45355);
and U45506 (N_45506,N_45484,N_45345);
nand U45507 (N_45507,N_45283,N_45474);
or U45508 (N_45508,N_45442,N_45260);
and U45509 (N_45509,N_45288,N_45480);
and U45510 (N_45510,N_45381,N_45323);
nand U45511 (N_45511,N_45286,N_45313);
or U45512 (N_45512,N_45359,N_45386);
xnor U45513 (N_45513,N_45327,N_45306);
and U45514 (N_45514,N_45486,N_45371);
and U45515 (N_45515,N_45380,N_45274);
or U45516 (N_45516,N_45264,N_45431);
xor U45517 (N_45517,N_45451,N_45301);
xnor U45518 (N_45518,N_45297,N_45463);
nand U45519 (N_45519,N_45389,N_45369);
and U45520 (N_45520,N_45496,N_45479);
nand U45521 (N_45521,N_45395,N_45449);
xnor U45522 (N_45522,N_45372,N_45481);
or U45523 (N_45523,N_45482,N_45307);
and U45524 (N_45524,N_45289,N_45438);
or U45525 (N_45525,N_45319,N_45278);
nor U45526 (N_45526,N_45346,N_45337);
nor U45527 (N_45527,N_45497,N_45348);
nor U45528 (N_45528,N_45317,N_45310);
nand U45529 (N_45529,N_45471,N_45312);
nand U45530 (N_45530,N_45304,N_45410);
and U45531 (N_45531,N_45360,N_45367);
and U45532 (N_45532,N_45258,N_45425);
and U45533 (N_45533,N_45423,N_45448);
or U45534 (N_45534,N_45309,N_45419);
nand U45535 (N_45535,N_45356,N_45368);
and U45536 (N_45536,N_45262,N_45466);
and U45537 (N_45537,N_45365,N_45458);
or U45538 (N_45538,N_45266,N_45468);
and U45539 (N_45539,N_45447,N_45461);
xor U45540 (N_45540,N_45424,N_45401);
xnor U45541 (N_45541,N_45455,N_45391);
nand U45542 (N_45542,N_45402,N_45341);
xor U45543 (N_45543,N_45364,N_45334);
or U45544 (N_45544,N_45352,N_45417);
xor U45545 (N_45545,N_45351,N_45429);
nor U45546 (N_45546,N_45490,N_45441);
or U45547 (N_45547,N_45287,N_45412);
and U45548 (N_45548,N_45376,N_45445);
nand U45549 (N_45549,N_45415,N_45488);
xor U45550 (N_45550,N_45370,N_45459);
nor U45551 (N_45551,N_45383,N_45489);
nor U45552 (N_45552,N_45392,N_45333);
and U45553 (N_45553,N_45433,N_45408);
or U45554 (N_45554,N_45465,N_45320);
nor U45555 (N_45555,N_45495,N_45450);
or U45556 (N_45556,N_45349,N_45403);
nand U45557 (N_45557,N_45361,N_45387);
nand U45558 (N_45558,N_45250,N_45270);
xor U45559 (N_45559,N_45322,N_45321);
or U45560 (N_45560,N_45358,N_45362);
xnor U45561 (N_45561,N_45453,N_45439);
xor U45562 (N_45562,N_45340,N_45492);
nor U45563 (N_45563,N_45342,N_45295);
xnor U45564 (N_45564,N_45284,N_45498);
nor U45565 (N_45565,N_45382,N_45343);
nor U45566 (N_45566,N_45363,N_45263);
and U45567 (N_45567,N_45261,N_45446);
nor U45568 (N_45568,N_45469,N_45409);
nor U45569 (N_45569,N_45332,N_45316);
nor U45570 (N_45570,N_45427,N_45375);
or U45571 (N_45571,N_45285,N_45338);
xnor U45572 (N_45572,N_45298,N_45475);
nand U45573 (N_45573,N_45434,N_45472);
xor U45574 (N_45574,N_45325,N_45331);
or U45575 (N_45575,N_45467,N_45291);
xor U45576 (N_45576,N_45357,N_45252);
xnor U45577 (N_45577,N_45437,N_45418);
or U45578 (N_45578,N_45335,N_45462);
or U45579 (N_45579,N_45253,N_45407);
nor U45580 (N_45580,N_45398,N_45470);
or U45581 (N_45581,N_45394,N_45454);
nor U45582 (N_45582,N_45413,N_45436);
and U45583 (N_45583,N_45339,N_45493);
and U45584 (N_45584,N_45483,N_45396);
nor U45585 (N_45585,N_45494,N_45254);
nand U45586 (N_45586,N_45390,N_45435);
and U45587 (N_45587,N_45315,N_45251);
nor U45588 (N_45588,N_45460,N_45299);
xor U45589 (N_45589,N_45336,N_45293);
and U45590 (N_45590,N_45416,N_45350);
xnor U45591 (N_45591,N_45272,N_45384);
nand U45592 (N_45592,N_45354,N_45378);
nor U45593 (N_45593,N_45268,N_45281);
nor U45594 (N_45594,N_45290,N_45473);
xor U45595 (N_45595,N_45256,N_45280);
xnor U45596 (N_45596,N_45428,N_45267);
nor U45597 (N_45597,N_45430,N_45276);
xor U45598 (N_45598,N_45314,N_45452);
and U45599 (N_45599,N_45464,N_45311);
or U45600 (N_45600,N_45443,N_45414);
nand U45601 (N_45601,N_45330,N_45294);
xor U45602 (N_45602,N_45302,N_45303);
nand U45603 (N_45603,N_45257,N_45326);
nor U45604 (N_45604,N_45476,N_45404);
nor U45605 (N_45605,N_45259,N_45478);
xor U45606 (N_45606,N_45292,N_45324);
nor U45607 (N_45607,N_45456,N_45318);
nand U45608 (N_45608,N_45411,N_45296);
nand U45609 (N_45609,N_45426,N_45300);
nor U45610 (N_45610,N_45432,N_45405);
xnor U45611 (N_45611,N_45269,N_45444);
nand U45612 (N_45612,N_45499,N_45440);
nand U45613 (N_45613,N_45377,N_45277);
or U45614 (N_45614,N_45308,N_45255);
and U45615 (N_45615,N_45393,N_45353);
xor U45616 (N_45616,N_45265,N_45457);
and U45617 (N_45617,N_45406,N_45422);
or U45618 (N_45618,N_45388,N_45344);
and U45619 (N_45619,N_45275,N_45329);
nand U45620 (N_45620,N_45273,N_45491);
nor U45621 (N_45621,N_45282,N_45421);
and U45622 (N_45622,N_45385,N_45420);
nor U45623 (N_45623,N_45477,N_45400);
nor U45624 (N_45624,N_45373,N_45366);
nor U45625 (N_45625,N_45287,N_45409);
nor U45626 (N_45626,N_45364,N_45264);
and U45627 (N_45627,N_45434,N_45274);
nand U45628 (N_45628,N_45362,N_45472);
nor U45629 (N_45629,N_45476,N_45383);
and U45630 (N_45630,N_45319,N_45256);
nand U45631 (N_45631,N_45489,N_45436);
and U45632 (N_45632,N_45426,N_45447);
nor U45633 (N_45633,N_45268,N_45364);
or U45634 (N_45634,N_45405,N_45392);
and U45635 (N_45635,N_45284,N_45300);
or U45636 (N_45636,N_45338,N_45486);
or U45637 (N_45637,N_45284,N_45417);
and U45638 (N_45638,N_45327,N_45362);
and U45639 (N_45639,N_45276,N_45469);
nand U45640 (N_45640,N_45330,N_45359);
xor U45641 (N_45641,N_45337,N_45451);
and U45642 (N_45642,N_45432,N_45433);
xnor U45643 (N_45643,N_45480,N_45314);
nand U45644 (N_45644,N_45495,N_45306);
xor U45645 (N_45645,N_45267,N_45407);
nand U45646 (N_45646,N_45332,N_45401);
xnor U45647 (N_45647,N_45409,N_45463);
nor U45648 (N_45648,N_45361,N_45389);
nand U45649 (N_45649,N_45392,N_45270);
nand U45650 (N_45650,N_45488,N_45394);
nand U45651 (N_45651,N_45323,N_45281);
xor U45652 (N_45652,N_45379,N_45448);
and U45653 (N_45653,N_45423,N_45252);
and U45654 (N_45654,N_45303,N_45361);
nor U45655 (N_45655,N_45412,N_45334);
and U45656 (N_45656,N_45264,N_45255);
nand U45657 (N_45657,N_45364,N_45333);
and U45658 (N_45658,N_45317,N_45265);
or U45659 (N_45659,N_45350,N_45294);
and U45660 (N_45660,N_45367,N_45425);
or U45661 (N_45661,N_45290,N_45489);
xnor U45662 (N_45662,N_45349,N_45399);
nand U45663 (N_45663,N_45466,N_45496);
nor U45664 (N_45664,N_45390,N_45410);
nand U45665 (N_45665,N_45312,N_45337);
or U45666 (N_45666,N_45322,N_45435);
xnor U45667 (N_45667,N_45434,N_45379);
or U45668 (N_45668,N_45339,N_45342);
nor U45669 (N_45669,N_45376,N_45462);
nand U45670 (N_45670,N_45372,N_45428);
and U45671 (N_45671,N_45478,N_45386);
xor U45672 (N_45672,N_45345,N_45487);
or U45673 (N_45673,N_45377,N_45324);
nand U45674 (N_45674,N_45333,N_45338);
or U45675 (N_45675,N_45453,N_45422);
xnor U45676 (N_45676,N_45364,N_45278);
nand U45677 (N_45677,N_45395,N_45322);
and U45678 (N_45678,N_45477,N_45393);
nand U45679 (N_45679,N_45455,N_45337);
or U45680 (N_45680,N_45345,N_45499);
or U45681 (N_45681,N_45291,N_45424);
nor U45682 (N_45682,N_45414,N_45423);
nor U45683 (N_45683,N_45380,N_45285);
or U45684 (N_45684,N_45421,N_45417);
xnor U45685 (N_45685,N_45488,N_45347);
xnor U45686 (N_45686,N_45295,N_45477);
xnor U45687 (N_45687,N_45481,N_45472);
nand U45688 (N_45688,N_45485,N_45290);
or U45689 (N_45689,N_45344,N_45339);
nand U45690 (N_45690,N_45489,N_45442);
or U45691 (N_45691,N_45472,N_45419);
or U45692 (N_45692,N_45466,N_45360);
or U45693 (N_45693,N_45454,N_45429);
nor U45694 (N_45694,N_45333,N_45382);
or U45695 (N_45695,N_45356,N_45456);
or U45696 (N_45696,N_45472,N_45324);
nor U45697 (N_45697,N_45297,N_45279);
or U45698 (N_45698,N_45434,N_45331);
nand U45699 (N_45699,N_45361,N_45324);
or U45700 (N_45700,N_45475,N_45323);
nor U45701 (N_45701,N_45294,N_45315);
xnor U45702 (N_45702,N_45454,N_45405);
or U45703 (N_45703,N_45316,N_45424);
xnor U45704 (N_45704,N_45345,N_45344);
and U45705 (N_45705,N_45355,N_45427);
nor U45706 (N_45706,N_45331,N_45405);
nand U45707 (N_45707,N_45479,N_45264);
or U45708 (N_45708,N_45344,N_45457);
nor U45709 (N_45709,N_45264,N_45336);
and U45710 (N_45710,N_45263,N_45428);
xor U45711 (N_45711,N_45287,N_45478);
xor U45712 (N_45712,N_45349,N_45412);
nand U45713 (N_45713,N_45309,N_45386);
and U45714 (N_45714,N_45381,N_45313);
and U45715 (N_45715,N_45369,N_45295);
or U45716 (N_45716,N_45387,N_45421);
nand U45717 (N_45717,N_45470,N_45294);
xnor U45718 (N_45718,N_45286,N_45266);
nand U45719 (N_45719,N_45394,N_45499);
nor U45720 (N_45720,N_45488,N_45335);
or U45721 (N_45721,N_45339,N_45417);
xnor U45722 (N_45722,N_45298,N_45499);
and U45723 (N_45723,N_45255,N_45465);
or U45724 (N_45724,N_45304,N_45417);
nand U45725 (N_45725,N_45305,N_45357);
xor U45726 (N_45726,N_45270,N_45320);
nor U45727 (N_45727,N_45419,N_45480);
or U45728 (N_45728,N_45325,N_45499);
nor U45729 (N_45729,N_45421,N_45453);
xor U45730 (N_45730,N_45344,N_45463);
nor U45731 (N_45731,N_45452,N_45261);
xor U45732 (N_45732,N_45465,N_45279);
nand U45733 (N_45733,N_45365,N_45251);
xor U45734 (N_45734,N_45434,N_45432);
nor U45735 (N_45735,N_45296,N_45454);
xor U45736 (N_45736,N_45482,N_45332);
and U45737 (N_45737,N_45487,N_45452);
and U45738 (N_45738,N_45282,N_45477);
nand U45739 (N_45739,N_45499,N_45443);
nand U45740 (N_45740,N_45260,N_45426);
nor U45741 (N_45741,N_45394,N_45268);
and U45742 (N_45742,N_45458,N_45499);
nor U45743 (N_45743,N_45483,N_45321);
and U45744 (N_45744,N_45269,N_45258);
or U45745 (N_45745,N_45428,N_45260);
and U45746 (N_45746,N_45317,N_45358);
and U45747 (N_45747,N_45406,N_45438);
or U45748 (N_45748,N_45383,N_45327);
nor U45749 (N_45749,N_45403,N_45308);
and U45750 (N_45750,N_45525,N_45648);
nor U45751 (N_45751,N_45651,N_45501);
nand U45752 (N_45752,N_45670,N_45715);
or U45753 (N_45753,N_45539,N_45674);
nor U45754 (N_45754,N_45581,N_45644);
and U45755 (N_45755,N_45510,N_45526);
nor U45756 (N_45756,N_45742,N_45589);
nor U45757 (N_45757,N_45628,N_45558);
or U45758 (N_45758,N_45575,N_45506);
and U45759 (N_45759,N_45641,N_45690);
nor U45760 (N_45760,N_45657,N_45730);
or U45761 (N_45761,N_45549,N_45547);
or U45762 (N_45762,N_45631,N_45602);
and U45763 (N_45763,N_45598,N_45746);
nor U45764 (N_45764,N_45633,N_45565);
or U45765 (N_45765,N_45551,N_45530);
or U45766 (N_45766,N_45745,N_45554);
xor U45767 (N_45767,N_45749,N_45584);
nand U45768 (N_45768,N_45500,N_45647);
nor U45769 (N_45769,N_45684,N_45531);
or U45770 (N_45770,N_45679,N_45614);
nand U45771 (N_45771,N_45702,N_45552);
nor U45772 (N_45772,N_45662,N_45603);
xor U45773 (N_45773,N_45509,N_45747);
nand U45774 (N_45774,N_45527,N_45518);
nand U45775 (N_45775,N_45536,N_45600);
and U45776 (N_45776,N_45706,N_45592);
nand U45777 (N_45777,N_45741,N_45704);
nand U45778 (N_45778,N_45634,N_45686);
and U45779 (N_45779,N_45635,N_45619);
or U45780 (N_45780,N_45541,N_45519);
or U45781 (N_45781,N_45587,N_45595);
and U45782 (N_45782,N_45740,N_45650);
and U45783 (N_45783,N_45543,N_45532);
and U45784 (N_45784,N_45523,N_45548);
xor U45785 (N_45785,N_45658,N_45724);
or U45786 (N_45786,N_45528,N_45620);
xnor U45787 (N_45787,N_45534,N_45728);
or U45788 (N_45788,N_45629,N_45639);
nor U45789 (N_45789,N_45712,N_45597);
and U45790 (N_45790,N_45569,N_45550);
and U45791 (N_45791,N_45721,N_45585);
nor U45792 (N_45792,N_45701,N_45748);
and U45793 (N_45793,N_45508,N_45642);
or U45794 (N_45794,N_45638,N_45676);
or U45795 (N_45795,N_45533,N_45599);
nor U45796 (N_45796,N_45618,N_45529);
and U45797 (N_45797,N_45653,N_45668);
and U45798 (N_45798,N_45563,N_45511);
or U45799 (N_45799,N_45683,N_45714);
or U45800 (N_45800,N_45744,N_45695);
nor U45801 (N_45801,N_45659,N_45698);
nand U45802 (N_45802,N_45694,N_45682);
nand U45803 (N_45803,N_45535,N_45718);
nand U45804 (N_45804,N_45703,N_45738);
nor U45805 (N_45805,N_45708,N_45732);
nand U45806 (N_45806,N_45725,N_45636);
or U45807 (N_45807,N_45666,N_45722);
nor U45808 (N_45808,N_45571,N_45665);
or U45809 (N_45809,N_45545,N_45719);
or U45810 (N_45810,N_45577,N_45556);
xor U45811 (N_45811,N_45664,N_45623);
xnor U45812 (N_45812,N_45553,N_45699);
and U45813 (N_45813,N_45546,N_45726);
and U45814 (N_45814,N_45669,N_45615);
nor U45815 (N_45815,N_45613,N_45542);
or U45816 (N_45816,N_45705,N_45608);
nand U45817 (N_45817,N_45514,N_45522);
and U45818 (N_45818,N_45579,N_45517);
xnor U45819 (N_45819,N_45538,N_45520);
nor U45820 (N_45820,N_45561,N_45649);
nand U45821 (N_45821,N_45559,N_45643);
or U45822 (N_45822,N_45504,N_45604);
xnor U45823 (N_45823,N_45612,N_45507);
xnor U45824 (N_45824,N_45734,N_45557);
xor U45825 (N_45825,N_45692,N_45717);
or U45826 (N_45826,N_45729,N_45564);
and U45827 (N_45827,N_45652,N_45617);
nand U45828 (N_45828,N_45691,N_45743);
or U45829 (N_45829,N_45663,N_45606);
and U45830 (N_45830,N_45630,N_45685);
and U45831 (N_45831,N_45582,N_45537);
and U45832 (N_45832,N_45656,N_45637);
nand U45833 (N_45833,N_45544,N_45601);
nand U45834 (N_45834,N_45687,N_45661);
and U45835 (N_45835,N_45524,N_45667);
nor U45836 (N_45836,N_45594,N_45503);
nand U45837 (N_45837,N_45671,N_45568);
xnor U45838 (N_45838,N_45591,N_45723);
nor U45839 (N_45839,N_45516,N_45632);
or U45840 (N_45840,N_45626,N_45609);
and U45841 (N_45841,N_45567,N_45576);
or U45842 (N_45842,N_45590,N_45583);
nand U45843 (N_45843,N_45621,N_45593);
nand U45844 (N_45844,N_45521,N_45570);
xor U45845 (N_45845,N_45515,N_45720);
xnor U45846 (N_45846,N_45512,N_45578);
nand U45847 (N_45847,N_45689,N_45605);
nand U45848 (N_45848,N_45560,N_45646);
or U45849 (N_45849,N_45513,N_45739);
and U45850 (N_45850,N_45680,N_45502);
nand U45851 (N_45851,N_45611,N_45627);
and U45852 (N_45852,N_45640,N_45700);
nor U45853 (N_45853,N_45711,N_45681);
and U45854 (N_45854,N_45673,N_45654);
or U45855 (N_45855,N_45622,N_45616);
and U45856 (N_45856,N_45716,N_45713);
nor U45857 (N_45857,N_45677,N_45586);
nand U45858 (N_45858,N_45709,N_45660);
xnor U45859 (N_45859,N_45625,N_45580);
and U45860 (N_45860,N_45624,N_45736);
xnor U45861 (N_45861,N_45555,N_45727);
xor U45862 (N_45862,N_45672,N_45573);
or U45863 (N_45863,N_45607,N_45610);
and U45864 (N_45864,N_45731,N_45697);
nor U45865 (N_45865,N_45707,N_45678);
xnor U45866 (N_45866,N_45688,N_45574);
nor U45867 (N_45867,N_45733,N_45572);
nor U45868 (N_45868,N_45696,N_45655);
or U45869 (N_45869,N_45588,N_45540);
or U45870 (N_45870,N_45735,N_45645);
or U45871 (N_45871,N_45596,N_45710);
nor U45872 (N_45872,N_45566,N_45505);
nor U45873 (N_45873,N_45737,N_45562);
and U45874 (N_45874,N_45693,N_45675);
and U45875 (N_45875,N_45548,N_45509);
xor U45876 (N_45876,N_45507,N_45676);
or U45877 (N_45877,N_45585,N_45595);
and U45878 (N_45878,N_45524,N_45506);
and U45879 (N_45879,N_45673,N_45574);
or U45880 (N_45880,N_45569,N_45564);
nand U45881 (N_45881,N_45640,N_45674);
and U45882 (N_45882,N_45650,N_45526);
xor U45883 (N_45883,N_45647,N_45608);
or U45884 (N_45884,N_45737,N_45607);
nor U45885 (N_45885,N_45630,N_45749);
xnor U45886 (N_45886,N_45677,N_45723);
nand U45887 (N_45887,N_45667,N_45638);
nor U45888 (N_45888,N_45627,N_45670);
or U45889 (N_45889,N_45722,N_45564);
xor U45890 (N_45890,N_45745,N_45689);
or U45891 (N_45891,N_45581,N_45523);
or U45892 (N_45892,N_45679,N_45567);
nand U45893 (N_45893,N_45595,N_45582);
or U45894 (N_45894,N_45699,N_45652);
nand U45895 (N_45895,N_45593,N_45540);
and U45896 (N_45896,N_45627,N_45531);
and U45897 (N_45897,N_45739,N_45602);
nand U45898 (N_45898,N_45504,N_45556);
nor U45899 (N_45899,N_45556,N_45619);
xor U45900 (N_45900,N_45518,N_45545);
xnor U45901 (N_45901,N_45635,N_45602);
xor U45902 (N_45902,N_45695,N_45619);
nor U45903 (N_45903,N_45693,N_45511);
nor U45904 (N_45904,N_45659,N_45568);
or U45905 (N_45905,N_45737,N_45668);
or U45906 (N_45906,N_45621,N_45501);
and U45907 (N_45907,N_45584,N_45629);
and U45908 (N_45908,N_45554,N_45645);
nand U45909 (N_45909,N_45590,N_45657);
or U45910 (N_45910,N_45544,N_45586);
and U45911 (N_45911,N_45519,N_45524);
and U45912 (N_45912,N_45512,N_45703);
xnor U45913 (N_45913,N_45504,N_45589);
xor U45914 (N_45914,N_45559,N_45744);
xnor U45915 (N_45915,N_45712,N_45505);
or U45916 (N_45916,N_45612,N_45747);
xnor U45917 (N_45917,N_45611,N_45646);
nor U45918 (N_45918,N_45674,N_45703);
or U45919 (N_45919,N_45531,N_45529);
or U45920 (N_45920,N_45637,N_45683);
nor U45921 (N_45921,N_45657,N_45613);
nor U45922 (N_45922,N_45731,N_45524);
or U45923 (N_45923,N_45722,N_45572);
and U45924 (N_45924,N_45501,N_45529);
and U45925 (N_45925,N_45700,N_45699);
and U45926 (N_45926,N_45583,N_45747);
xor U45927 (N_45927,N_45525,N_45538);
or U45928 (N_45928,N_45661,N_45673);
or U45929 (N_45929,N_45645,N_45727);
or U45930 (N_45930,N_45621,N_45560);
or U45931 (N_45931,N_45723,N_45668);
nor U45932 (N_45932,N_45654,N_45584);
xor U45933 (N_45933,N_45617,N_45573);
or U45934 (N_45934,N_45630,N_45621);
and U45935 (N_45935,N_45592,N_45586);
nand U45936 (N_45936,N_45629,N_45534);
and U45937 (N_45937,N_45614,N_45605);
xnor U45938 (N_45938,N_45646,N_45634);
xor U45939 (N_45939,N_45561,N_45667);
xor U45940 (N_45940,N_45559,N_45656);
xnor U45941 (N_45941,N_45606,N_45519);
nand U45942 (N_45942,N_45703,N_45618);
nor U45943 (N_45943,N_45582,N_45580);
or U45944 (N_45944,N_45603,N_45746);
or U45945 (N_45945,N_45594,N_45746);
or U45946 (N_45946,N_45688,N_45569);
nor U45947 (N_45947,N_45662,N_45648);
nand U45948 (N_45948,N_45684,N_45594);
and U45949 (N_45949,N_45575,N_45648);
and U45950 (N_45950,N_45585,N_45644);
and U45951 (N_45951,N_45691,N_45593);
xor U45952 (N_45952,N_45603,N_45502);
xor U45953 (N_45953,N_45694,N_45699);
xnor U45954 (N_45954,N_45683,N_45610);
xor U45955 (N_45955,N_45708,N_45701);
nand U45956 (N_45956,N_45689,N_45629);
xor U45957 (N_45957,N_45703,N_45682);
and U45958 (N_45958,N_45540,N_45666);
or U45959 (N_45959,N_45686,N_45737);
nor U45960 (N_45960,N_45632,N_45741);
or U45961 (N_45961,N_45558,N_45707);
and U45962 (N_45962,N_45654,N_45639);
nor U45963 (N_45963,N_45532,N_45594);
and U45964 (N_45964,N_45507,N_45689);
and U45965 (N_45965,N_45523,N_45738);
xnor U45966 (N_45966,N_45617,N_45555);
xor U45967 (N_45967,N_45652,N_45560);
nor U45968 (N_45968,N_45602,N_45523);
xor U45969 (N_45969,N_45564,N_45664);
nor U45970 (N_45970,N_45689,N_45737);
xnor U45971 (N_45971,N_45534,N_45532);
and U45972 (N_45972,N_45632,N_45729);
nand U45973 (N_45973,N_45599,N_45612);
and U45974 (N_45974,N_45650,N_45533);
nand U45975 (N_45975,N_45675,N_45651);
or U45976 (N_45976,N_45601,N_45673);
nand U45977 (N_45977,N_45616,N_45687);
nand U45978 (N_45978,N_45662,N_45744);
and U45979 (N_45979,N_45695,N_45528);
or U45980 (N_45980,N_45623,N_45609);
nor U45981 (N_45981,N_45550,N_45623);
nand U45982 (N_45982,N_45642,N_45727);
nand U45983 (N_45983,N_45511,N_45729);
xnor U45984 (N_45984,N_45536,N_45673);
xnor U45985 (N_45985,N_45515,N_45575);
nand U45986 (N_45986,N_45500,N_45534);
or U45987 (N_45987,N_45596,N_45538);
and U45988 (N_45988,N_45666,N_45526);
nor U45989 (N_45989,N_45628,N_45724);
nand U45990 (N_45990,N_45680,N_45586);
nand U45991 (N_45991,N_45582,N_45719);
xnor U45992 (N_45992,N_45567,N_45514);
and U45993 (N_45993,N_45644,N_45636);
and U45994 (N_45994,N_45660,N_45604);
nand U45995 (N_45995,N_45674,N_45563);
nand U45996 (N_45996,N_45731,N_45532);
nand U45997 (N_45997,N_45637,N_45747);
nor U45998 (N_45998,N_45670,N_45700);
nand U45999 (N_45999,N_45533,N_45652);
and U46000 (N_46000,N_45949,N_45764);
xor U46001 (N_46001,N_45817,N_45879);
xor U46002 (N_46002,N_45829,N_45998);
nor U46003 (N_46003,N_45915,N_45780);
and U46004 (N_46004,N_45835,N_45993);
nor U46005 (N_46005,N_45801,N_45920);
and U46006 (N_46006,N_45972,N_45784);
xnor U46007 (N_46007,N_45957,N_45753);
nand U46008 (N_46008,N_45927,N_45837);
nand U46009 (N_46009,N_45865,N_45904);
nand U46010 (N_46010,N_45838,N_45751);
or U46011 (N_46011,N_45875,N_45812);
and U46012 (N_46012,N_45975,N_45902);
nor U46013 (N_46013,N_45762,N_45997);
xnor U46014 (N_46014,N_45897,N_45776);
and U46015 (N_46015,N_45987,N_45825);
and U46016 (N_46016,N_45916,N_45851);
nand U46017 (N_46017,N_45775,N_45768);
nand U46018 (N_46018,N_45863,N_45956);
nor U46019 (N_46019,N_45900,N_45894);
or U46020 (N_46020,N_45983,N_45815);
nor U46021 (N_46021,N_45982,N_45771);
nand U46022 (N_46022,N_45866,N_45846);
and U46023 (N_46023,N_45928,N_45790);
and U46024 (N_46024,N_45887,N_45889);
and U46025 (N_46025,N_45994,N_45988);
nor U46026 (N_46026,N_45864,N_45845);
xor U46027 (N_46027,N_45999,N_45870);
xor U46028 (N_46028,N_45763,N_45770);
nor U46029 (N_46029,N_45824,N_45756);
and U46030 (N_46030,N_45926,N_45939);
xor U46031 (N_46031,N_45867,N_45818);
and U46032 (N_46032,N_45809,N_45974);
nand U46033 (N_46033,N_45929,N_45934);
and U46034 (N_46034,N_45789,N_45787);
or U46035 (N_46035,N_45954,N_45816);
xor U46036 (N_46036,N_45759,N_45944);
and U46037 (N_46037,N_45914,N_45839);
xor U46038 (N_46038,N_45858,N_45805);
nand U46039 (N_46039,N_45951,N_45912);
nand U46040 (N_46040,N_45862,N_45895);
nand U46041 (N_46041,N_45847,N_45832);
nor U46042 (N_46042,N_45883,N_45868);
xnor U46043 (N_46043,N_45891,N_45774);
xnor U46044 (N_46044,N_45853,N_45948);
or U46045 (N_46045,N_45917,N_45826);
nor U46046 (N_46046,N_45992,N_45821);
nand U46047 (N_46047,N_45856,N_45802);
nor U46048 (N_46048,N_45849,N_45943);
nand U46049 (N_46049,N_45785,N_45991);
nor U46050 (N_46050,N_45947,N_45886);
xor U46051 (N_46051,N_45871,N_45976);
xnor U46052 (N_46052,N_45986,N_45810);
or U46053 (N_46053,N_45936,N_45901);
nor U46054 (N_46054,N_45755,N_45781);
nor U46055 (N_46055,N_45841,N_45808);
nor U46056 (N_46056,N_45823,N_45857);
xnor U46057 (N_46057,N_45990,N_45799);
nor U46058 (N_46058,N_45783,N_45950);
xnor U46059 (N_46059,N_45923,N_45910);
xnor U46060 (N_46060,N_45820,N_45946);
or U46061 (N_46061,N_45859,N_45911);
nand U46062 (N_46062,N_45773,N_45968);
and U46063 (N_46063,N_45873,N_45814);
xnor U46064 (N_46064,N_45971,N_45788);
nor U46065 (N_46065,N_45919,N_45852);
nand U46066 (N_46066,N_45804,N_45767);
nor U46067 (N_46067,N_45938,N_45981);
or U46068 (N_46068,N_45973,N_45960);
or U46069 (N_46069,N_45791,N_45778);
nor U46070 (N_46070,N_45893,N_45888);
and U46071 (N_46071,N_45798,N_45874);
or U46072 (N_46072,N_45786,N_45962);
nand U46073 (N_46073,N_45933,N_45827);
xor U46074 (N_46074,N_45937,N_45909);
xor U46075 (N_46075,N_45931,N_45892);
and U46076 (N_46076,N_45842,N_45899);
or U46077 (N_46077,N_45766,N_45854);
or U46078 (N_46078,N_45978,N_45752);
xnor U46079 (N_46079,N_45796,N_45930);
nor U46080 (N_46080,N_45795,N_45807);
nor U46081 (N_46081,N_45833,N_45855);
or U46082 (N_46082,N_45964,N_45958);
nand U46083 (N_46083,N_45800,N_45906);
nand U46084 (N_46084,N_45794,N_45880);
nand U46085 (N_46085,N_45952,N_45877);
and U46086 (N_46086,N_45830,N_45924);
nor U46087 (N_46087,N_45872,N_45869);
and U46088 (N_46088,N_45876,N_45935);
xnor U46089 (N_46089,N_45861,N_45942);
or U46090 (N_46090,N_45761,N_45806);
nand U46091 (N_46091,N_45966,N_45757);
or U46092 (N_46092,N_45918,N_45977);
nand U46093 (N_46093,N_45922,N_45792);
xnor U46094 (N_46094,N_45836,N_45878);
nor U46095 (N_46095,N_45758,N_45813);
or U46096 (N_46096,N_45777,N_45995);
or U46097 (N_46097,N_45765,N_45925);
nor U46098 (N_46098,N_45908,N_45890);
nor U46099 (N_46099,N_45782,N_45996);
xnor U46100 (N_46100,N_45980,N_45811);
xnor U46101 (N_46101,N_45819,N_45769);
nor U46102 (N_46102,N_45989,N_45967);
nand U46103 (N_46103,N_45905,N_45860);
xnor U46104 (N_46104,N_45898,N_45896);
or U46105 (N_46105,N_45844,N_45961);
nor U46106 (N_46106,N_45955,N_45803);
or U46107 (N_46107,N_45760,N_45884);
nor U46108 (N_46108,N_45921,N_45848);
and U46109 (N_46109,N_45850,N_45941);
and U46110 (N_46110,N_45828,N_45882);
nor U46111 (N_46111,N_45831,N_45750);
nand U46112 (N_46112,N_45822,N_45969);
nand U46113 (N_46113,N_45772,N_45970);
and U46114 (N_46114,N_45834,N_45793);
xor U46115 (N_46115,N_45903,N_45779);
xor U46116 (N_46116,N_45959,N_45953);
nand U46117 (N_46117,N_45885,N_45913);
or U46118 (N_46118,N_45965,N_45881);
and U46119 (N_46119,N_45945,N_45843);
nand U46120 (N_46120,N_45940,N_45932);
or U46121 (N_46121,N_45979,N_45797);
and U46122 (N_46122,N_45963,N_45907);
or U46123 (N_46123,N_45754,N_45984);
or U46124 (N_46124,N_45985,N_45840);
nand U46125 (N_46125,N_45920,N_45982);
xor U46126 (N_46126,N_45966,N_45946);
or U46127 (N_46127,N_45904,N_45918);
nor U46128 (N_46128,N_45799,N_45901);
xor U46129 (N_46129,N_45771,N_45887);
or U46130 (N_46130,N_45844,N_45880);
nor U46131 (N_46131,N_45817,N_45975);
xnor U46132 (N_46132,N_45907,N_45842);
or U46133 (N_46133,N_45928,N_45806);
nor U46134 (N_46134,N_45965,N_45853);
nor U46135 (N_46135,N_45943,N_45833);
and U46136 (N_46136,N_45945,N_45937);
xor U46137 (N_46137,N_45783,N_45780);
xnor U46138 (N_46138,N_45858,N_45777);
or U46139 (N_46139,N_45905,N_45977);
or U46140 (N_46140,N_45768,N_45960);
and U46141 (N_46141,N_45930,N_45928);
nand U46142 (N_46142,N_45845,N_45981);
and U46143 (N_46143,N_45973,N_45935);
nand U46144 (N_46144,N_45808,N_45806);
xor U46145 (N_46145,N_45761,N_45927);
nand U46146 (N_46146,N_45866,N_45783);
or U46147 (N_46147,N_45846,N_45929);
or U46148 (N_46148,N_45849,N_45817);
nor U46149 (N_46149,N_45946,N_45782);
xnor U46150 (N_46150,N_45883,N_45943);
xnor U46151 (N_46151,N_45767,N_45934);
or U46152 (N_46152,N_45797,N_45761);
xor U46153 (N_46153,N_45870,N_45841);
nor U46154 (N_46154,N_45908,N_45984);
nor U46155 (N_46155,N_45886,N_45775);
xor U46156 (N_46156,N_45902,N_45916);
or U46157 (N_46157,N_45814,N_45848);
nand U46158 (N_46158,N_45963,N_45884);
nor U46159 (N_46159,N_45929,N_45886);
or U46160 (N_46160,N_45892,N_45944);
or U46161 (N_46161,N_45990,N_45875);
nor U46162 (N_46162,N_45835,N_45757);
or U46163 (N_46163,N_45867,N_45922);
nor U46164 (N_46164,N_45940,N_45936);
nor U46165 (N_46165,N_45785,N_45754);
and U46166 (N_46166,N_45915,N_45795);
xnor U46167 (N_46167,N_45910,N_45993);
xor U46168 (N_46168,N_45951,N_45858);
xnor U46169 (N_46169,N_45816,N_45984);
nand U46170 (N_46170,N_45757,N_45980);
nor U46171 (N_46171,N_45806,N_45805);
xor U46172 (N_46172,N_45933,N_45872);
and U46173 (N_46173,N_45844,N_45782);
or U46174 (N_46174,N_45791,N_45772);
nand U46175 (N_46175,N_45976,N_45959);
nor U46176 (N_46176,N_45757,N_45826);
xnor U46177 (N_46177,N_45761,N_45870);
xor U46178 (N_46178,N_45792,N_45949);
nor U46179 (N_46179,N_45969,N_45913);
and U46180 (N_46180,N_45799,N_45991);
and U46181 (N_46181,N_45768,N_45806);
nand U46182 (N_46182,N_45758,N_45823);
or U46183 (N_46183,N_45813,N_45992);
nor U46184 (N_46184,N_45838,N_45912);
nor U46185 (N_46185,N_45813,N_45863);
or U46186 (N_46186,N_45988,N_45945);
or U46187 (N_46187,N_45993,N_45800);
nor U46188 (N_46188,N_45919,N_45752);
and U46189 (N_46189,N_45773,N_45761);
nor U46190 (N_46190,N_45760,N_45854);
or U46191 (N_46191,N_45825,N_45812);
and U46192 (N_46192,N_45844,N_45965);
xor U46193 (N_46193,N_45902,N_45949);
xnor U46194 (N_46194,N_45798,N_45780);
xor U46195 (N_46195,N_45931,N_45797);
or U46196 (N_46196,N_45801,N_45969);
and U46197 (N_46197,N_45791,N_45780);
or U46198 (N_46198,N_45820,N_45895);
nor U46199 (N_46199,N_45947,N_45864);
and U46200 (N_46200,N_45962,N_45852);
nor U46201 (N_46201,N_45792,N_45867);
xnor U46202 (N_46202,N_45953,N_45806);
xor U46203 (N_46203,N_45961,N_45969);
or U46204 (N_46204,N_45964,N_45915);
or U46205 (N_46205,N_45897,N_45911);
nand U46206 (N_46206,N_45926,N_45868);
nor U46207 (N_46207,N_45904,N_45922);
xnor U46208 (N_46208,N_45970,N_45782);
xor U46209 (N_46209,N_45821,N_45996);
nor U46210 (N_46210,N_45905,N_45867);
xor U46211 (N_46211,N_45780,N_45853);
nor U46212 (N_46212,N_45804,N_45753);
and U46213 (N_46213,N_45752,N_45837);
or U46214 (N_46214,N_45968,N_45763);
nand U46215 (N_46215,N_45983,N_45933);
xor U46216 (N_46216,N_45764,N_45964);
or U46217 (N_46217,N_45937,N_45821);
or U46218 (N_46218,N_45984,N_45856);
xor U46219 (N_46219,N_45989,N_45810);
nand U46220 (N_46220,N_45815,N_45897);
nor U46221 (N_46221,N_45865,N_45972);
xor U46222 (N_46222,N_45996,N_45769);
nand U46223 (N_46223,N_45878,N_45899);
nor U46224 (N_46224,N_45789,N_45842);
and U46225 (N_46225,N_45810,N_45834);
nand U46226 (N_46226,N_45886,N_45888);
and U46227 (N_46227,N_45869,N_45768);
and U46228 (N_46228,N_45824,N_45874);
nor U46229 (N_46229,N_45771,N_45946);
and U46230 (N_46230,N_45839,N_45953);
and U46231 (N_46231,N_45970,N_45872);
or U46232 (N_46232,N_45852,N_45756);
nor U46233 (N_46233,N_45786,N_45989);
nor U46234 (N_46234,N_45819,N_45864);
and U46235 (N_46235,N_45780,N_45815);
nor U46236 (N_46236,N_45852,N_45904);
and U46237 (N_46237,N_45977,N_45875);
xnor U46238 (N_46238,N_45811,N_45751);
nor U46239 (N_46239,N_45816,N_45858);
xnor U46240 (N_46240,N_45928,N_45840);
xor U46241 (N_46241,N_45826,N_45773);
xnor U46242 (N_46242,N_45870,N_45757);
nor U46243 (N_46243,N_45880,N_45757);
and U46244 (N_46244,N_45903,N_45929);
nand U46245 (N_46245,N_45962,N_45854);
or U46246 (N_46246,N_45975,N_45852);
nand U46247 (N_46247,N_45997,N_45862);
and U46248 (N_46248,N_45905,N_45921);
and U46249 (N_46249,N_45932,N_45879);
and U46250 (N_46250,N_46007,N_46181);
and U46251 (N_46251,N_46241,N_46059);
xnor U46252 (N_46252,N_46021,N_46222);
or U46253 (N_46253,N_46178,N_46191);
or U46254 (N_46254,N_46030,N_46065);
nor U46255 (N_46255,N_46019,N_46011);
and U46256 (N_46256,N_46123,N_46046);
and U46257 (N_46257,N_46055,N_46047);
and U46258 (N_46258,N_46200,N_46010);
and U46259 (N_46259,N_46216,N_46048);
and U46260 (N_46260,N_46195,N_46056);
xnor U46261 (N_46261,N_46132,N_46185);
nand U46262 (N_46262,N_46208,N_46173);
xnor U46263 (N_46263,N_46001,N_46203);
or U46264 (N_46264,N_46229,N_46108);
xor U46265 (N_46265,N_46221,N_46008);
and U46266 (N_46266,N_46044,N_46149);
xnor U46267 (N_46267,N_46086,N_46169);
or U46268 (N_46268,N_46189,N_46163);
and U46269 (N_46269,N_46031,N_46128);
or U46270 (N_46270,N_46093,N_46207);
and U46271 (N_46271,N_46246,N_46198);
nand U46272 (N_46272,N_46182,N_46218);
and U46273 (N_46273,N_46150,N_46175);
nand U46274 (N_46274,N_46183,N_46227);
and U46275 (N_46275,N_46094,N_46244);
or U46276 (N_46276,N_46122,N_46170);
nand U46277 (N_46277,N_46049,N_46077);
nor U46278 (N_46278,N_46157,N_46014);
nor U46279 (N_46279,N_46211,N_46147);
or U46280 (N_46280,N_46034,N_46112);
nor U46281 (N_46281,N_46167,N_46103);
nor U46282 (N_46282,N_46239,N_46105);
or U46283 (N_46283,N_46206,N_46201);
nand U46284 (N_46284,N_46004,N_46113);
and U46285 (N_46285,N_46158,N_46151);
nor U46286 (N_46286,N_46025,N_46115);
xor U46287 (N_46287,N_46141,N_46002);
and U46288 (N_46288,N_46058,N_46243);
xor U46289 (N_46289,N_46231,N_46165);
xnor U46290 (N_46290,N_46172,N_46090);
or U46291 (N_46291,N_46040,N_46135);
and U46292 (N_46292,N_46152,N_46130);
nand U46293 (N_46293,N_46080,N_46045);
or U46294 (N_46294,N_46196,N_46085);
nand U46295 (N_46295,N_46136,N_46225);
nor U46296 (N_46296,N_46022,N_46199);
nand U46297 (N_46297,N_46162,N_46212);
and U46298 (N_46298,N_46076,N_46042);
xor U46299 (N_46299,N_46125,N_46133);
or U46300 (N_46300,N_46068,N_46037);
nor U46301 (N_46301,N_46180,N_46116);
or U46302 (N_46302,N_46064,N_46043);
and U46303 (N_46303,N_46102,N_46119);
and U46304 (N_46304,N_46186,N_46174);
nor U46305 (N_46305,N_46005,N_46168);
xnor U46306 (N_46306,N_46213,N_46033);
and U46307 (N_46307,N_46016,N_46220);
nand U46308 (N_46308,N_46024,N_46069);
and U46309 (N_46309,N_46171,N_46204);
nand U46310 (N_46310,N_46029,N_46015);
nor U46311 (N_46311,N_46249,N_46083);
and U46312 (N_46312,N_46032,N_46143);
and U46313 (N_46313,N_46230,N_46101);
nor U46314 (N_46314,N_46139,N_46228);
nand U46315 (N_46315,N_46134,N_46209);
or U46316 (N_46316,N_46138,N_46193);
xnor U46317 (N_46317,N_46248,N_46109);
xor U46318 (N_46318,N_46131,N_46236);
nor U46319 (N_46319,N_46197,N_46051);
or U46320 (N_46320,N_46041,N_46081);
nor U46321 (N_46321,N_46217,N_46145);
or U46322 (N_46322,N_46177,N_46053);
and U46323 (N_46323,N_46070,N_46137);
or U46324 (N_46324,N_46234,N_46121);
or U46325 (N_46325,N_46050,N_46091);
nand U46326 (N_46326,N_46194,N_46009);
or U46327 (N_46327,N_46071,N_46142);
nand U46328 (N_46328,N_46219,N_46214);
nor U46329 (N_46329,N_46066,N_46082);
or U46330 (N_46330,N_46052,N_46224);
or U46331 (N_46331,N_46003,N_46153);
or U46332 (N_46332,N_46054,N_46072);
nand U46333 (N_46333,N_46018,N_46144);
nor U46334 (N_46334,N_46060,N_46164);
and U46335 (N_46335,N_46089,N_46120);
nand U46336 (N_46336,N_46245,N_46006);
nor U46337 (N_46337,N_46099,N_46100);
nor U46338 (N_46338,N_46036,N_46154);
or U46339 (N_46339,N_46238,N_46097);
nor U46340 (N_46340,N_46190,N_46179);
and U46341 (N_46341,N_46156,N_46240);
xnor U46342 (N_46342,N_46184,N_46247);
or U46343 (N_46343,N_46104,N_46235);
nand U46344 (N_46344,N_46166,N_46129);
nor U46345 (N_46345,N_46148,N_46028);
nor U46346 (N_46346,N_46092,N_46242);
and U46347 (N_46347,N_46078,N_46017);
or U46348 (N_46348,N_46187,N_46000);
and U46349 (N_46349,N_46233,N_46107);
nor U46350 (N_46350,N_46188,N_46013);
xnor U46351 (N_46351,N_46075,N_46088);
or U46352 (N_46352,N_46226,N_46114);
nor U46353 (N_46353,N_46205,N_46126);
nor U46354 (N_46354,N_46232,N_46161);
nand U46355 (N_46355,N_46127,N_46095);
nor U46356 (N_46356,N_46012,N_46118);
nand U46357 (N_46357,N_46237,N_46146);
nor U46358 (N_46358,N_46038,N_46098);
or U46359 (N_46359,N_46210,N_46160);
nand U46360 (N_46360,N_46061,N_46035);
xor U46361 (N_46361,N_46087,N_46106);
nand U46362 (N_46362,N_46062,N_46084);
or U46363 (N_46363,N_46202,N_46026);
xnor U46364 (N_46364,N_46176,N_46020);
and U46365 (N_46365,N_46057,N_46039);
nor U46366 (N_46366,N_46140,N_46074);
and U46367 (N_46367,N_46063,N_46155);
and U46368 (N_46368,N_46159,N_46192);
nand U46369 (N_46369,N_46067,N_46110);
or U46370 (N_46370,N_46096,N_46079);
and U46371 (N_46371,N_46124,N_46215);
xor U46372 (N_46372,N_46117,N_46111);
xor U46373 (N_46373,N_46223,N_46023);
or U46374 (N_46374,N_46073,N_46027);
or U46375 (N_46375,N_46117,N_46198);
or U46376 (N_46376,N_46093,N_46136);
and U46377 (N_46377,N_46161,N_46101);
xor U46378 (N_46378,N_46173,N_46028);
or U46379 (N_46379,N_46078,N_46133);
and U46380 (N_46380,N_46014,N_46156);
nand U46381 (N_46381,N_46150,N_46133);
xnor U46382 (N_46382,N_46197,N_46055);
nor U46383 (N_46383,N_46247,N_46129);
or U46384 (N_46384,N_46009,N_46097);
xor U46385 (N_46385,N_46208,N_46046);
and U46386 (N_46386,N_46042,N_46173);
nand U46387 (N_46387,N_46111,N_46091);
nand U46388 (N_46388,N_46175,N_46165);
xnor U46389 (N_46389,N_46154,N_46225);
or U46390 (N_46390,N_46061,N_46023);
xnor U46391 (N_46391,N_46230,N_46146);
nand U46392 (N_46392,N_46138,N_46192);
nor U46393 (N_46393,N_46079,N_46214);
nor U46394 (N_46394,N_46063,N_46220);
nand U46395 (N_46395,N_46239,N_46108);
and U46396 (N_46396,N_46226,N_46230);
and U46397 (N_46397,N_46179,N_46175);
or U46398 (N_46398,N_46024,N_46090);
and U46399 (N_46399,N_46067,N_46061);
nor U46400 (N_46400,N_46236,N_46112);
and U46401 (N_46401,N_46098,N_46167);
and U46402 (N_46402,N_46243,N_46060);
nor U46403 (N_46403,N_46054,N_46145);
or U46404 (N_46404,N_46036,N_46176);
and U46405 (N_46405,N_46214,N_46228);
or U46406 (N_46406,N_46222,N_46199);
or U46407 (N_46407,N_46082,N_46177);
and U46408 (N_46408,N_46180,N_46050);
or U46409 (N_46409,N_46160,N_46244);
xor U46410 (N_46410,N_46026,N_46044);
xnor U46411 (N_46411,N_46103,N_46249);
xnor U46412 (N_46412,N_46084,N_46041);
nor U46413 (N_46413,N_46234,N_46095);
nand U46414 (N_46414,N_46009,N_46220);
or U46415 (N_46415,N_46167,N_46073);
nand U46416 (N_46416,N_46112,N_46168);
xor U46417 (N_46417,N_46204,N_46201);
nor U46418 (N_46418,N_46085,N_46106);
and U46419 (N_46419,N_46069,N_46195);
or U46420 (N_46420,N_46023,N_46097);
nand U46421 (N_46421,N_46204,N_46050);
or U46422 (N_46422,N_46162,N_46215);
nand U46423 (N_46423,N_46052,N_46101);
nor U46424 (N_46424,N_46064,N_46037);
xor U46425 (N_46425,N_46008,N_46224);
or U46426 (N_46426,N_46249,N_46183);
nand U46427 (N_46427,N_46008,N_46097);
nand U46428 (N_46428,N_46211,N_46184);
nor U46429 (N_46429,N_46185,N_46182);
nand U46430 (N_46430,N_46238,N_46189);
nor U46431 (N_46431,N_46027,N_46204);
xnor U46432 (N_46432,N_46140,N_46055);
and U46433 (N_46433,N_46136,N_46249);
or U46434 (N_46434,N_46190,N_46104);
and U46435 (N_46435,N_46235,N_46055);
nand U46436 (N_46436,N_46129,N_46215);
or U46437 (N_46437,N_46190,N_46133);
nand U46438 (N_46438,N_46040,N_46060);
or U46439 (N_46439,N_46132,N_46228);
nand U46440 (N_46440,N_46112,N_46160);
nand U46441 (N_46441,N_46119,N_46070);
nand U46442 (N_46442,N_46111,N_46153);
nand U46443 (N_46443,N_46122,N_46035);
nand U46444 (N_46444,N_46185,N_46079);
nand U46445 (N_46445,N_46081,N_46156);
nand U46446 (N_46446,N_46050,N_46174);
or U46447 (N_46447,N_46074,N_46070);
nor U46448 (N_46448,N_46194,N_46079);
and U46449 (N_46449,N_46076,N_46037);
or U46450 (N_46450,N_46236,N_46064);
nand U46451 (N_46451,N_46091,N_46044);
or U46452 (N_46452,N_46010,N_46099);
xor U46453 (N_46453,N_46015,N_46218);
or U46454 (N_46454,N_46194,N_46071);
nand U46455 (N_46455,N_46008,N_46124);
and U46456 (N_46456,N_46065,N_46191);
nand U46457 (N_46457,N_46183,N_46155);
or U46458 (N_46458,N_46047,N_46146);
and U46459 (N_46459,N_46222,N_46122);
or U46460 (N_46460,N_46135,N_46016);
or U46461 (N_46461,N_46111,N_46184);
or U46462 (N_46462,N_46014,N_46249);
nor U46463 (N_46463,N_46050,N_46085);
nor U46464 (N_46464,N_46121,N_46017);
nand U46465 (N_46465,N_46081,N_46057);
nand U46466 (N_46466,N_46115,N_46096);
xor U46467 (N_46467,N_46167,N_46130);
nand U46468 (N_46468,N_46103,N_46176);
xnor U46469 (N_46469,N_46246,N_46010);
and U46470 (N_46470,N_46125,N_46174);
and U46471 (N_46471,N_46136,N_46162);
nand U46472 (N_46472,N_46175,N_46109);
nor U46473 (N_46473,N_46166,N_46029);
xor U46474 (N_46474,N_46203,N_46123);
or U46475 (N_46475,N_46162,N_46121);
and U46476 (N_46476,N_46154,N_46174);
xnor U46477 (N_46477,N_46096,N_46223);
xnor U46478 (N_46478,N_46127,N_46184);
xnor U46479 (N_46479,N_46072,N_46181);
nand U46480 (N_46480,N_46070,N_46248);
or U46481 (N_46481,N_46170,N_46193);
xor U46482 (N_46482,N_46002,N_46061);
xor U46483 (N_46483,N_46191,N_46213);
or U46484 (N_46484,N_46051,N_46178);
nand U46485 (N_46485,N_46177,N_46225);
nand U46486 (N_46486,N_46249,N_46154);
and U46487 (N_46487,N_46234,N_46076);
and U46488 (N_46488,N_46175,N_46220);
nor U46489 (N_46489,N_46168,N_46192);
nand U46490 (N_46490,N_46130,N_46243);
and U46491 (N_46491,N_46142,N_46190);
nor U46492 (N_46492,N_46057,N_46040);
xor U46493 (N_46493,N_46145,N_46193);
nor U46494 (N_46494,N_46145,N_46122);
and U46495 (N_46495,N_46163,N_46090);
or U46496 (N_46496,N_46084,N_46111);
nand U46497 (N_46497,N_46214,N_46102);
xnor U46498 (N_46498,N_46018,N_46157);
or U46499 (N_46499,N_46247,N_46023);
xor U46500 (N_46500,N_46438,N_46278);
nand U46501 (N_46501,N_46307,N_46434);
or U46502 (N_46502,N_46300,N_46403);
nor U46503 (N_46503,N_46474,N_46364);
nand U46504 (N_46504,N_46436,N_46431);
xor U46505 (N_46505,N_46303,N_46387);
xnor U46506 (N_46506,N_46411,N_46425);
nand U46507 (N_46507,N_46294,N_46275);
and U46508 (N_46508,N_46476,N_46441);
nor U46509 (N_46509,N_46258,N_46333);
and U46510 (N_46510,N_46488,N_46435);
nand U46511 (N_46511,N_46397,N_46311);
and U46512 (N_46512,N_46326,N_46382);
or U46513 (N_46513,N_46454,N_46388);
or U46514 (N_46514,N_46408,N_46473);
or U46515 (N_46515,N_46396,N_46318);
xor U46516 (N_46516,N_46464,N_46290);
xnor U46517 (N_46517,N_46460,N_46301);
nand U46518 (N_46518,N_46412,N_46305);
nand U46519 (N_46519,N_46314,N_46283);
or U46520 (N_46520,N_46368,N_46274);
and U46521 (N_46521,N_46292,N_46400);
and U46522 (N_46522,N_46369,N_46445);
nand U46523 (N_46523,N_46362,N_46325);
xnor U46524 (N_46524,N_46321,N_46443);
and U46525 (N_46525,N_46337,N_46461);
nand U46526 (N_46526,N_46279,N_46291);
xor U46527 (N_46527,N_46486,N_46354);
nand U46528 (N_46528,N_46379,N_46330);
and U46529 (N_46529,N_46253,N_46478);
nor U46530 (N_46530,N_46350,N_46427);
xnor U46531 (N_46531,N_46293,N_46365);
nor U46532 (N_46532,N_46463,N_46410);
xnor U46533 (N_46533,N_46328,N_46252);
nor U46534 (N_46534,N_46334,N_46415);
and U46535 (N_46535,N_46457,N_46356);
and U46536 (N_46536,N_46261,N_46381);
nor U46537 (N_46537,N_46298,N_46455);
nand U46538 (N_46538,N_46484,N_46419);
and U46539 (N_46539,N_46270,N_46492);
and U46540 (N_46540,N_46495,N_46479);
and U46541 (N_46541,N_46348,N_46340);
nand U46542 (N_46542,N_46355,N_46416);
and U46543 (N_46543,N_46444,N_46341);
and U46544 (N_46544,N_46485,N_46272);
nand U46545 (N_46545,N_46332,N_46376);
or U46546 (N_46546,N_46377,N_46451);
or U46547 (N_46547,N_46498,N_46407);
nand U46548 (N_46548,N_46353,N_46256);
and U46549 (N_46549,N_46393,N_46289);
nor U46550 (N_46550,N_46367,N_46442);
nand U46551 (N_46551,N_46255,N_46342);
or U46552 (N_46552,N_46277,N_46259);
nor U46553 (N_46553,N_46312,N_46349);
nand U46554 (N_46554,N_46296,N_46361);
xnor U46555 (N_46555,N_46469,N_46446);
xnor U46556 (N_46556,N_46375,N_46497);
or U46557 (N_46557,N_46327,N_46264);
and U46558 (N_46558,N_46331,N_46316);
xnor U46559 (N_46559,N_46392,N_46406);
and U46560 (N_46560,N_46459,N_46266);
and U46561 (N_46561,N_46466,N_46384);
xor U46562 (N_46562,N_46339,N_46386);
and U46563 (N_46563,N_46372,N_46366);
nor U46564 (N_46564,N_46491,N_46271);
and U46565 (N_46565,N_46371,N_46468);
xor U46566 (N_46566,N_46329,N_46346);
or U46567 (N_46567,N_46475,N_46380);
nor U46568 (N_46568,N_46470,N_46399);
xor U46569 (N_46569,N_46324,N_46430);
or U46570 (N_46570,N_46398,N_46404);
or U46571 (N_46571,N_46286,N_46414);
xor U46572 (N_46572,N_46257,N_46458);
and U46573 (N_46573,N_46343,N_46347);
nand U46574 (N_46574,N_46378,N_46323);
or U46575 (N_46575,N_46302,N_46417);
or U46576 (N_46576,N_46453,N_46304);
and U46577 (N_46577,N_46281,N_46269);
xnor U46578 (N_46578,N_46424,N_46359);
xnor U46579 (N_46579,N_46482,N_46383);
nor U46580 (N_46580,N_46450,N_46260);
xnor U46581 (N_46581,N_46351,N_46370);
and U46582 (N_46582,N_46280,N_46481);
nor U46583 (N_46583,N_46336,N_46320);
and U46584 (N_46584,N_46447,N_46480);
nand U46585 (N_46585,N_46319,N_46405);
or U46586 (N_46586,N_46308,N_46490);
nor U46587 (N_46587,N_46487,N_46413);
or U46588 (N_46588,N_46306,N_46448);
and U46589 (N_46589,N_46250,N_46373);
xnor U46590 (N_46590,N_46428,N_46267);
and U46591 (N_46591,N_46284,N_46317);
nor U46592 (N_46592,N_46360,N_46254);
xnor U46593 (N_46593,N_46437,N_46322);
nand U46594 (N_46594,N_46456,N_46295);
xor U46595 (N_46595,N_46483,N_46477);
and U46596 (N_46596,N_46287,N_46313);
nand U46597 (N_46597,N_46345,N_46462);
and U46598 (N_46598,N_46489,N_46285);
xnor U46599 (N_46599,N_46315,N_46268);
nand U46600 (N_46600,N_46309,N_46374);
and U46601 (N_46601,N_46394,N_46265);
or U46602 (N_46602,N_46262,N_46297);
or U46603 (N_46603,N_46421,N_46494);
or U46604 (N_46604,N_46344,N_46429);
xor U46605 (N_46605,N_46439,N_46401);
nand U46606 (N_46606,N_46471,N_46465);
nand U46607 (N_46607,N_46472,N_46282);
xnor U46608 (N_46608,N_46288,N_46263);
nor U46609 (N_46609,N_46493,N_46389);
or U46610 (N_46610,N_46422,N_46335);
nor U46611 (N_46611,N_46385,N_46418);
nand U46612 (N_46612,N_46299,N_46440);
and U46613 (N_46613,N_46402,N_46467);
or U46614 (N_46614,N_46338,N_46452);
or U46615 (N_46615,N_46310,N_46449);
or U46616 (N_46616,N_46499,N_46273);
xor U46617 (N_46617,N_46426,N_46352);
or U46618 (N_46618,N_46358,N_46409);
nand U46619 (N_46619,N_46357,N_46390);
nand U46620 (N_46620,N_46433,N_46420);
and U46621 (N_46621,N_46395,N_46391);
or U46622 (N_46622,N_46432,N_46496);
nand U46623 (N_46623,N_46363,N_46251);
nand U46624 (N_46624,N_46423,N_46276);
xnor U46625 (N_46625,N_46413,N_46257);
xnor U46626 (N_46626,N_46327,N_46423);
nand U46627 (N_46627,N_46403,N_46408);
and U46628 (N_46628,N_46361,N_46396);
or U46629 (N_46629,N_46341,N_46460);
and U46630 (N_46630,N_46385,N_46376);
nor U46631 (N_46631,N_46425,N_46422);
and U46632 (N_46632,N_46331,N_46398);
nor U46633 (N_46633,N_46380,N_46498);
xnor U46634 (N_46634,N_46408,N_46325);
xor U46635 (N_46635,N_46436,N_46333);
nor U46636 (N_46636,N_46499,N_46319);
and U46637 (N_46637,N_46319,N_46318);
xnor U46638 (N_46638,N_46360,N_46273);
and U46639 (N_46639,N_46443,N_46308);
xor U46640 (N_46640,N_46274,N_46414);
nand U46641 (N_46641,N_46411,N_46368);
nand U46642 (N_46642,N_46391,N_46428);
and U46643 (N_46643,N_46354,N_46293);
nand U46644 (N_46644,N_46400,N_46419);
nand U46645 (N_46645,N_46393,N_46454);
nor U46646 (N_46646,N_46397,N_46341);
or U46647 (N_46647,N_46326,N_46489);
and U46648 (N_46648,N_46415,N_46351);
nand U46649 (N_46649,N_46271,N_46424);
xnor U46650 (N_46650,N_46396,N_46338);
nor U46651 (N_46651,N_46326,N_46288);
and U46652 (N_46652,N_46497,N_46431);
nand U46653 (N_46653,N_46459,N_46407);
xor U46654 (N_46654,N_46461,N_46279);
nor U46655 (N_46655,N_46466,N_46450);
nor U46656 (N_46656,N_46296,N_46450);
and U46657 (N_46657,N_46318,N_46373);
and U46658 (N_46658,N_46354,N_46341);
and U46659 (N_46659,N_46288,N_46439);
xor U46660 (N_46660,N_46267,N_46438);
or U46661 (N_46661,N_46493,N_46380);
and U46662 (N_46662,N_46366,N_46395);
or U46663 (N_46663,N_46285,N_46415);
or U46664 (N_46664,N_46443,N_46455);
and U46665 (N_46665,N_46485,N_46497);
and U46666 (N_46666,N_46387,N_46357);
or U46667 (N_46667,N_46379,N_46367);
or U46668 (N_46668,N_46378,N_46296);
and U46669 (N_46669,N_46320,N_46360);
xor U46670 (N_46670,N_46281,N_46407);
xor U46671 (N_46671,N_46257,N_46407);
or U46672 (N_46672,N_46310,N_46360);
xor U46673 (N_46673,N_46315,N_46456);
nor U46674 (N_46674,N_46299,N_46498);
xnor U46675 (N_46675,N_46325,N_46370);
nor U46676 (N_46676,N_46438,N_46286);
and U46677 (N_46677,N_46471,N_46399);
nand U46678 (N_46678,N_46485,N_46364);
and U46679 (N_46679,N_46348,N_46465);
or U46680 (N_46680,N_46470,N_46377);
xnor U46681 (N_46681,N_46260,N_46322);
xnor U46682 (N_46682,N_46477,N_46312);
or U46683 (N_46683,N_46349,N_46497);
and U46684 (N_46684,N_46252,N_46405);
nor U46685 (N_46685,N_46305,N_46473);
or U46686 (N_46686,N_46476,N_46483);
nor U46687 (N_46687,N_46469,N_46317);
xor U46688 (N_46688,N_46382,N_46417);
or U46689 (N_46689,N_46412,N_46485);
and U46690 (N_46690,N_46395,N_46294);
and U46691 (N_46691,N_46496,N_46423);
xor U46692 (N_46692,N_46448,N_46344);
nor U46693 (N_46693,N_46431,N_46493);
nor U46694 (N_46694,N_46326,N_46304);
nor U46695 (N_46695,N_46317,N_46392);
and U46696 (N_46696,N_46405,N_46285);
nor U46697 (N_46697,N_46331,N_46261);
xnor U46698 (N_46698,N_46287,N_46377);
nand U46699 (N_46699,N_46499,N_46425);
and U46700 (N_46700,N_46441,N_46253);
or U46701 (N_46701,N_46396,N_46289);
or U46702 (N_46702,N_46468,N_46476);
xnor U46703 (N_46703,N_46366,N_46392);
or U46704 (N_46704,N_46311,N_46498);
or U46705 (N_46705,N_46343,N_46393);
xnor U46706 (N_46706,N_46309,N_46440);
xnor U46707 (N_46707,N_46298,N_46313);
or U46708 (N_46708,N_46448,N_46351);
or U46709 (N_46709,N_46331,N_46442);
or U46710 (N_46710,N_46344,N_46360);
nor U46711 (N_46711,N_46391,N_46497);
nor U46712 (N_46712,N_46459,N_46467);
and U46713 (N_46713,N_46486,N_46393);
or U46714 (N_46714,N_46440,N_46277);
xor U46715 (N_46715,N_46369,N_46470);
nor U46716 (N_46716,N_46474,N_46414);
xnor U46717 (N_46717,N_46485,N_46311);
and U46718 (N_46718,N_46250,N_46444);
nand U46719 (N_46719,N_46346,N_46413);
xor U46720 (N_46720,N_46360,N_46332);
nor U46721 (N_46721,N_46303,N_46362);
and U46722 (N_46722,N_46326,N_46370);
nand U46723 (N_46723,N_46375,N_46255);
nor U46724 (N_46724,N_46385,N_46338);
or U46725 (N_46725,N_46260,N_46377);
and U46726 (N_46726,N_46453,N_46457);
nor U46727 (N_46727,N_46251,N_46491);
nand U46728 (N_46728,N_46466,N_46300);
xnor U46729 (N_46729,N_46486,N_46270);
and U46730 (N_46730,N_46308,N_46299);
and U46731 (N_46731,N_46450,N_46323);
or U46732 (N_46732,N_46289,N_46416);
or U46733 (N_46733,N_46331,N_46301);
and U46734 (N_46734,N_46469,N_46343);
or U46735 (N_46735,N_46258,N_46371);
nor U46736 (N_46736,N_46397,N_46361);
nor U46737 (N_46737,N_46377,N_46328);
and U46738 (N_46738,N_46356,N_46422);
or U46739 (N_46739,N_46252,N_46302);
or U46740 (N_46740,N_46441,N_46402);
xnor U46741 (N_46741,N_46442,N_46309);
nor U46742 (N_46742,N_46449,N_46440);
nor U46743 (N_46743,N_46270,N_46362);
and U46744 (N_46744,N_46436,N_46421);
and U46745 (N_46745,N_46255,N_46357);
and U46746 (N_46746,N_46481,N_46474);
xnor U46747 (N_46747,N_46489,N_46346);
nor U46748 (N_46748,N_46303,N_46318);
xnor U46749 (N_46749,N_46262,N_46468);
nand U46750 (N_46750,N_46661,N_46546);
nor U46751 (N_46751,N_46567,N_46624);
and U46752 (N_46752,N_46521,N_46692);
and U46753 (N_46753,N_46588,N_46647);
nor U46754 (N_46754,N_46620,N_46511);
xor U46755 (N_46755,N_46659,N_46633);
or U46756 (N_46756,N_46506,N_46741);
nor U46757 (N_46757,N_46686,N_46621);
nor U46758 (N_46758,N_46527,N_46535);
and U46759 (N_46759,N_46644,N_46690);
nand U46760 (N_46760,N_46580,N_46597);
or U46761 (N_46761,N_46502,N_46678);
nand U46762 (N_46762,N_46704,N_46524);
and U46763 (N_46763,N_46585,N_46572);
nor U46764 (N_46764,N_46691,N_46592);
or U46765 (N_46765,N_46587,N_46709);
or U46766 (N_46766,N_46549,N_46662);
xnor U46767 (N_46767,N_46573,N_46627);
nor U46768 (N_46768,N_46653,N_46618);
nand U46769 (N_46769,N_46687,N_46697);
and U46770 (N_46770,N_46566,N_46702);
or U46771 (N_46771,N_46735,N_46666);
nor U46772 (N_46772,N_46615,N_46715);
nor U46773 (N_46773,N_46552,N_46510);
nand U46774 (N_46774,N_46718,N_46614);
nor U46775 (N_46775,N_46571,N_46551);
or U46776 (N_46776,N_46579,N_46746);
nand U46777 (N_46777,N_46721,N_46658);
or U46778 (N_46778,N_46730,N_46663);
xor U46779 (N_46779,N_46557,N_46714);
or U46780 (N_46780,N_46544,N_46748);
xnor U46781 (N_46781,N_46637,N_46628);
xnor U46782 (N_46782,N_46708,N_46584);
nand U46783 (N_46783,N_46560,N_46516);
nand U46784 (N_46784,N_46734,N_46533);
or U46785 (N_46785,N_46643,N_46582);
nand U46786 (N_46786,N_46529,N_46558);
or U46787 (N_46787,N_46609,N_46564);
xnor U46788 (N_46788,N_46530,N_46668);
nand U46789 (N_46789,N_46747,N_46606);
or U46790 (N_46790,N_46684,N_46539);
nand U46791 (N_46791,N_46595,N_46739);
or U46792 (N_46792,N_46727,N_46639);
and U46793 (N_46793,N_46669,N_46542);
nor U46794 (N_46794,N_46737,N_46561);
and U46795 (N_46795,N_46505,N_46512);
and U46796 (N_46796,N_46645,N_46685);
or U46797 (N_46797,N_46673,N_46581);
and U46798 (N_46798,N_46519,N_46728);
and U46799 (N_46799,N_46532,N_46711);
xnor U46800 (N_46800,N_46553,N_46513);
xnor U46801 (N_46801,N_46696,N_46503);
and U46802 (N_46802,N_46742,N_46672);
nor U46803 (N_46803,N_46738,N_46689);
nor U46804 (N_46804,N_46607,N_46724);
and U46805 (N_46805,N_46594,N_46731);
or U46806 (N_46806,N_46586,N_46712);
or U46807 (N_46807,N_46682,N_46634);
nand U46808 (N_46808,N_46676,N_46719);
and U46809 (N_46809,N_46548,N_46547);
and U46810 (N_46810,N_46694,N_46660);
xnor U46811 (N_46811,N_46622,N_46670);
nor U46812 (N_46812,N_46514,N_46578);
xnor U46813 (N_46813,N_46574,N_46612);
nand U46814 (N_46814,N_46652,N_46657);
xor U46815 (N_46815,N_46635,N_46610);
nor U46816 (N_46816,N_46743,N_46613);
or U46817 (N_46817,N_46650,N_46568);
xnor U46818 (N_46818,N_46744,N_46555);
or U46819 (N_46819,N_46675,N_46641);
and U46820 (N_46820,N_46693,N_46733);
nand U46821 (N_46821,N_46536,N_46596);
nor U46822 (N_46822,N_46745,N_46648);
nor U46823 (N_46823,N_46570,N_46683);
and U46824 (N_46824,N_46525,N_46665);
nor U46825 (N_46825,N_46541,N_46608);
and U46826 (N_46826,N_46654,N_46729);
or U46827 (N_46827,N_46522,N_46664);
and U46828 (N_46828,N_46720,N_46629);
nor U46829 (N_46829,N_46563,N_46601);
and U46830 (N_46830,N_46501,N_46680);
nor U46831 (N_46831,N_46705,N_46545);
nand U46832 (N_46832,N_46713,N_46520);
and U46833 (N_46833,N_46651,N_46716);
xor U46834 (N_46834,N_46632,N_46554);
and U46835 (N_46835,N_46515,N_46626);
and U46836 (N_46836,N_46740,N_46577);
and U46837 (N_46837,N_46600,N_46543);
and U46838 (N_46838,N_46500,N_46504);
xor U46839 (N_46839,N_46698,N_46725);
nor U46840 (N_46840,N_46569,N_46593);
and U46841 (N_46841,N_46508,N_46736);
and U46842 (N_46842,N_46642,N_46617);
xnor U46843 (N_46843,N_46667,N_46625);
xor U46844 (N_46844,N_46540,N_46707);
nand U46845 (N_46845,N_46605,N_46559);
nor U46846 (N_46846,N_46699,N_46603);
nand U46847 (N_46847,N_46636,N_46732);
or U46848 (N_46848,N_46526,N_46726);
xnor U46849 (N_46849,N_46722,N_46590);
or U46850 (N_46850,N_46531,N_46674);
or U46851 (N_46851,N_46681,N_46583);
nor U46852 (N_46852,N_46523,N_46565);
or U46853 (N_46853,N_46591,N_46640);
nor U46854 (N_46854,N_46749,N_46517);
nor U46855 (N_46855,N_46695,N_46646);
xnor U46856 (N_46856,N_46710,N_46677);
xor U46857 (N_46857,N_46619,N_46671);
or U46858 (N_46858,N_46589,N_46616);
xnor U46859 (N_46859,N_46538,N_46550);
or U46860 (N_46860,N_46518,N_46700);
and U46861 (N_46861,N_46575,N_46534);
and U46862 (N_46862,N_46537,N_46528);
or U46863 (N_46863,N_46688,N_46602);
nor U46864 (N_46864,N_46723,N_46703);
or U46865 (N_46865,N_46556,N_46562);
nand U46866 (N_46866,N_46598,N_46623);
and U46867 (N_46867,N_46576,N_46656);
nor U46868 (N_46868,N_46638,N_46701);
and U46869 (N_46869,N_46611,N_46706);
and U46870 (N_46870,N_46679,N_46630);
and U46871 (N_46871,N_46717,N_46507);
and U46872 (N_46872,N_46599,N_46649);
or U46873 (N_46873,N_46631,N_46509);
xor U46874 (N_46874,N_46604,N_46655);
and U46875 (N_46875,N_46738,N_46581);
nand U46876 (N_46876,N_46701,N_46707);
xor U46877 (N_46877,N_46602,N_46511);
nand U46878 (N_46878,N_46704,N_46688);
or U46879 (N_46879,N_46628,N_46529);
and U46880 (N_46880,N_46690,N_46566);
or U46881 (N_46881,N_46685,N_46526);
xor U46882 (N_46882,N_46698,N_46630);
or U46883 (N_46883,N_46648,N_46684);
nand U46884 (N_46884,N_46529,N_46728);
nand U46885 (N_46885,N_46509,N_46596);
nor U46886 (N_46886,N_46563,N_46717);
and U46887 (N_46887,N_46505,N_46623);
and U46888 (N_46888,N_46652,N_46611);
xnor U46889 (N_46889,N_46612,N_46644);
nand U46890 (N_46890,N_46617,N_46585);
xnor U46891 (N_46891,N_46564,N_46526);
nor U46892 (N_46892,N_46648,N_46596);
xnor U46893 (N_46893,N_46695,N_46552);
or U46894 (N_46894,N_46655,N_46711);
and U46895 (N_46895,N_46515,N_46567);
nor U46896 (N_46896,N_46533,N_46521);
xor U46897 (N_46897,N_46682,N_46695);
nor U46898 (N_46898,N_46675,N_46599);
xnor U46899 (N_46899,N_46698,N_46672);
or U46900 (N_46900,N_46546,N_46597);
nand U46901 (N_46901,N_46692,N_46734);
nand U46902 (N_46902,N_46636,N_46509);
nand U46903 (N_46903,N_46525,N_46599);
and U46904 (N_46904,N_46527,N_46536);
nor U46905 (N_46905,N_46594,N_46562);
nor U46906 (N_46906,N_46650,N_46512);
nand U46907 (N_46907,N_46511,N_46627);
and U46908 (N_46908,N_46675,N_46749);
xnor U46909 (N_46909,N_46725,N_46567);
nor U46910 (N_46910,N_46514,N_46607);
and U46911 (N_46911,N_46510,N_46592);
xnor U46912 (N_46912,N_46716,N_46646);
nand U46913 (N_46913,N_46593,N_46510);
xor U46914 (N_46914,N_46626,N_46576);
nand U46915 (N_46915,N_46697,N_46663);
xnor U46916 (N_46916,N_46618,N_46655);
or U46917 (N_46917,N_46713,N_46651);
or U46918 (N_46918,N_46584,N_46501);
or U46919 (N_46919,N_46709,N_46546);
nand U46920 (N_46920,N_46672,N_46697);
xor U46921 (N_46921,N_46501,N_46726);
or U46922 (N_46922,N_46518,N_46620);
or U46923 (N_46923,N_46513,N_46602);
and U46924 (N_46924,N_46501,N_46601);
nor U46925 (N_46925,N_46520,N_46646);
or U46926 (N_46926,N_46626,N_46691);
or U46927 (N_46927,N_46645,N_46513);
nor U46928 (N_46928,N_46526,N_46513);
nor U46929 (N_46929,N_46712,N_46585);
nand U46930 (N_46930,N_46633,N_46562);
xor U46931 (N_46931,N_46654,N_46639);
nand U46932 (N_46932,N_46712,N_46504);
or U46933 (N_46933,N_46665,N_46551);
nor U46934 (N_46934,N_46573,N_46583);
nor U46935 (N_46935,N_46609,N_46533);
and U46936 (N_46936,N_46665,N_46663);
and U46937 (N_46937,N_46569,N_46654);
nand U46938 (N_46938,N_46596,N_46678);
or U46939 (N_46939,N_46516,N_46661);
xor U46940 (N_46940,N_46713,N_46529);
nor U46941 (N_46941,N_46580,N_46591);
nand U46942 (N_46942,N_46615,N_46554);
xnor U46943 (N_46943,N_46599,N_46645);
nor U46944 (N_46944,N_46695,N_46568);
or U46945 (N_46945,N_46619,N_46733);
xnor U46946 (N_46946,N_46708,N_46705);
nand U46947 (N_46947,N_46647,N_46685);
nor U46948 (N_46948,N_46737,N_46685);
or U46949 (N_46949,N_46724,N_46522);
nor U46950 (N_46950,N_46706,N_46677);
and U46951 (N_46951,N_46697,N_46595);
nor U46952 (N_46952,N_46737,N_46545);
or U46953 (N_46953,N_46533,N_46682);
nor U46954 (N_46954,N_46720,N_46732);
nor U46955 (N_46955,N_46576,N_46678);
xnor U46956 (N_46956,N_46626,N_46539);
or U46957 (N_46957,N_46654,N_46699);
nor U46958 (N_46958,N_46629,N_46525);
nor U46959 (N_46959,N_46653,N_46613);
or U46960 (N_46960,N_46527,N_46731);
and U46961 (N_46961,N_46505,N_46719);
xnor U46962 (N_46962,N_46661,N_46644);
xor U46963 (N_46963,N_46710,N_46655);
xor U46964 (N_46964,N_46697,N_46679);
and U46965 (N_46965,N_46628,N_46662);
or U46966 (N_46966,N_46687,N_46742);
and U46967 (N_46967,N_46703,N_46542);
and U46968 (N_46968,N_46710,N_46712);
or U46969 (N_46969,N_46593,N_46588);
xnor U46970 (N_46970,N_46585,N_46638);
or U46971 (N_46971,N_46693,N_46547);
xnor U46972 (N_46972,N_46702,N_46628);
xnor U46973 (N_46973,N_46649,N_46739);
or U46974 (N_46974,N_46513,N_46695);
nor U46975 (N_46975,N_46605,N_46689);
nand U46976 (N_46976,N_46726,N_46676);
and U46977 (N_46977,N_46714,N_46538);
and U46978 (N_46978,N_46523,N_46515);
and U46979 (N_46979,N_46624,N_46636);
or U46980 (N_46980,N_46532,N_46547);
and U46981 (N_46981,N_46560,N_46628);
and U46982 (N_46982,N_46743,N_46733);
xor U46983 (N_46983,N_46614,N_46717);
and U46984 (N_46984,N_46684,N_46680);
or U46985 (N_46985,N_46688,N_46540);
and U46986 (N_46986,N_46554,N_46737);
nor U46987 (N_46987,N_46648,N_46525);
or U46988 (N_46988,N_46546,N_46670);
or U46989 (N_46989,N_46717,N_46596);
and U46990 (N_46990,N_46551,N_46509);
and U46991 (N_46991,N_46589,N_46518);
and U46992 (N_46992,N_46654,N_46567);
or U46993 (N_46993,N_46506,N_46677);
xor U46994 (N_46994,N_46715,N_46667);
nor U46995 (N_46995,N_46549,N_46551);
and U46996 (N_46996,N_46518,N_46636);
nand U46997 (N_46997,N_46631,N_46694);
xor U46998 (N_46998,N_46682,N_46616);
nor U46999 (N_46999,N_46512,N_46682);
and U47000 (N_47000,N_46960,N_46761);
or U47001 (N_47001,N_46996,N_46959);
and U47002 (N_47002,N_46913,N_46887);
or U47003 (N_47003,N_46900,N_46822);
nor U47004 (N_47004,N_46999,N_46926);
nor U47005 (N_47005,N_46944,N_46813);
xor U47006 (N_47006,N_46973,N_46940);
xnor U47007 (N_47007,N_46980,N_46861);
or U47008 (N_47008,N_46930,N_46911);
or U47009 (N_47009,N_46833,N_46829);
nor U47010 (N_47010,N_46751,N_46789);
nor U47011 (N_47011,N_46947,N_46756);
xnor U47012 (N_47012,N_46938,N_46910);
nor U47013 (N_47013,N_46794,N_46948);
nor U47014 (N_47014,N_46962,N_46974);
xnor U47015 (N_47015,N_46847,N_46872);
nor U47016 (N_47016,N_46891,N_46839);
and U47017 (N_47017,N_46988,N_46969);
or U47018 (N_47018,N_46840,N_46846);
nor U47019 (N_47019,N_46752,N_46936);
or U47020 (N_47020,N_46904,N_46773);
or U47021 (N_47021,N_46848,N_46866);
or U47022 (N_47022,N_46803,N_46933);
nor U47023 (N_47023,N_46915,N_46986);
xor U47024 (N_47024,N_46838,N_46855);
or U47025 (N_47025,N_46992,N_46985);
and U47026 (N_47026,N_46819,N_46903);
nand U47027 (N_47027,N_46865,N_46876);
nor U47028 (N_47028,N_46957,N_46864);
and U47029 (N_47029,N_46852,N_46873);
nor U47030 (N_47030,N_46827,N_46856);
nor U47031 (N_47031,N_46899,N_46858);
nand U47032 (N_47032,N_46995,N_46878);
nor U47033 (N_47033,N_46853,N_46975);
nand U47034 (N_47034,N_46919,N_46890);
nor U47035 (N_47035,N_46954,N_46921);
nand U47036 (N_47036,N_46805,N_46800);
xor U47037 (N_47037,N_46791,N_46880);
nor U47038 (N_47038,N_46871,N_46877);
nor U47039 (N_47039,N_46835,N_46777);
and U47040 (N_47040,N_46909,N_46780);
nand U47041 (N_47041,N_46949,N_46997);
xnor U47042 (N_47042,N_46811,N_46793);
nand U47043 (N_47043,N_46883,N_46893);
xnor U47044 (N_47044,N_46993,N_46812);
nor U47045 (N_47045,N_46897,N_46758);
xor U47046 (N_47046,N_46932,N_46809);
or U47047 (N_47047,N_46970,N_46823);
nor U47048 (N_47048,N_46977,N_46831);
nand U47049 (N_47049,N_46929,N_46917);
and U47050 (N_47050,N_46796,N_46792);
and U47051 (N_47051,N_46895,N_46770);
nand U47052 (N_47052,N_46862,N_46854);
or U47053 (N_47053,N_46912,N_46801);
or U47054 (N_47054,N_46828,N_46968);
nand U47055 (N_47055,N_46928,N_46908);
and U47056 (N_47056,N_46953,N_46905);
or U47057 (N_47057,N_46884,N_46764);
nand U47058 (N_47058,N_46766,N_46989);
and U47059 (N_47059,N_46771,N_46788);
and U47060 (N_47060,N_46804,N_46981);
and U47061 (N_47061,N_46881,N_46907);
and U47062 (N_47062,N_46830,N_46857);
xor U47063 (N_47063,N_46863,N_46879);
xor U47064 (N_47064,N_46979,N_46841);
nor U47065 (N_47065,N_46760,N_46934);
or U47066 (N_47066,N_46869,N_46951);
or U47067 (N_47067,N_46935,N_46843);
or U47068 (N_47068,N_46785,N_46956);
nor U47069 (N_47069,N_46914,N_46783);
nand U47070 (N_47070,N_46987,N_46939);
or U47071 (N_47071,N_46781,N_46918);
or U47072 (N_47072,N_46983,N_46994);
nor U47073 (N_47073,N_46757,N_46927);
nor U47074 (N_47074,N_46937,N_46765);
nand U47075 (N_47075,N_46844,N_46799);
xor U47076 (N_47076,N_46920,N_46946);
or U47077 (N_47077,N_46806,N_46963);
nand U47078 (N_47078,N_46860,N_46961);
and U47079 (N_47079,N_46776,N_46754);
nand U47080 (N_47080,N_46824,N_46825);
or U47081 (N_47081,N_46851,N_46889);
or U47082 (N_47082,N_46849,N_46998);
nor U47083 (N_47083,N_46941,N_46759);
or U47084 (N_47084,N_46774,N_46964);
nor U47085 (N_47085,N_46815,N_46808);
xor U47086 (N_47086,N_46984,N_46894);
nand U47087 (N_47087,N_46882,N_46836);
nor U47088 (N_47088,N_46787,N_46931);
nor U47089 (N_47089,N_46779,N_46901);
xnor U47090 (N_47090,N_46845,N_46972);
or U47091 (N_47091,N_46784,N_46820);
nand U47092 (N_47092,N_46782,N_46795);
nand U47093 (N_47093,N_46924,N_46925);
or U47094 (N_47094,N_46753,N_46943);
or U47095 (N_47095,N_46775,N_46867);
nor U47096 (N_47096,N_46790,N_46875);
or U47097 (N_47097,N_46842,N_46902);
or U47098 (N_47098,N_46814,N_46991);
nand U47099 (N_47099,N_46955,N_46976);
nor U47100 (N_47100,N_46906,N_46898);
nor U47101 (N_47101,N_46817,N_46942);
nand U47102 (N_47102,N_46971,N_46923);
xor U47103 (N_47103,N_46945,N_46802);
nand U47104 (N_47104,N_46922,N_46834);
nor U47105 (N_47105,N_46952,N_46896);
nand U47106 (N_47106,N_46797,N_46885);
nor U47107 (N_47107,N_46762,N_46886);
xnor U47108 (N_47108,N_46786,N_46916);
nand U47109 (N_47109,N_46778,N_46850);
xnor U47110 (N_47110,N_46763,N_46816);
or U47111 (N_47111,N_46868,N_46958);
xnor U47112 (N_47112,N_46768,N_46888);
and U47113 (N_47113,N_46767,N_46837);
xnor U47114 (N_47114,N_46832,N_46950);
or U47115 (N_47115,N_46965,N_46978);
or U47116 (N_47116,N_46967,N_46798);
nor U47117 (N_47117,N_46892,N_46826);
nand U47118 (N_47118,N_46769,N_46750);
and U47119 (N_47119,N_46870,N_46990);
nand U47120 (N_47120,N_46982,N_46859);
and U47121 (N_47121,N_46807,N_46772);
or U47122 (N_47122,N_46818,N_46966);
and U47123 (N_47123,N_46810,N_46874);
nor U47124 (N_47124,N_46755,N_46821);
nand U47125 (N_47125,N_46853,N_46836);
or U47126 (N_47126,N_46973,N_46852);
xnor U47127 (N_47127,N_46971,N_46865);
nand U47128 (N_47128,N_46851,N_46976);
xor U47129 (N_47129,N_46999,N_46796);
nor U47130 (N_47130,N_46827,N_46924);
nor U47131 (N_47131,N_46997,N_46785);
nand U47132 (N_47132,N_46845,N_46842);
or U47133 (N_47133,N_46852,N_46813);
or U47134 (N_47134,N_46955,N_46759);
nor U47135 (N_47135,N_46975,N_46771);
nor U47136 (N_47136,N_46816,N_46776);
and U47137 (N_47137,N_46813,N_46916);
xnor U47138 (N_47138,N_46915,N_46851);
or U47139 (N_47139,N_46933,N_46799);
nand U47140 (N_47140,N_46838,N_46824);
or U47141 (N_47141,N_46857,N_46761);
or U47142 (N_47142,N_46824,N_46906);
xor U47143 (N_47143,N_46804,N_46777);
or U47144 (N_47144,N_46775,N_46786);
nand U47145 (N_47145,N_46760,N_46902);
xnor U47146 (N_47146,N_46832,N_46921);
nor U47147 (N_47147,N_46777,N_46755);
nor U47148 (N_47148,N_46809,N_46972);
nand U47149 (N_47149,N_46859,N_46983);
or U47150 (N_47150,N_46992,N_46955);
nor U47151 (N_47151,N_46775,N_46919);
and U47152 (N_47152,N_46930,N_46942);
xor U47153 (N_47153,N_46930,N_46953);
nand U47154 (N_47154,N_46831,N_46786);
xor U47155 (N_47155,N_46859,N_46804);
nor U47156 (N_47156,N_46870,N_46809);
nand U47157 (N_47157,N_46881,N_46942);
and U47158 (N_47158,N_46900,N_46852);
nand U47159 (N_47159,N_46956,N_46810);
and U47160 (N_47160,N_46934,N_46793);
nand U47161 (N_47161,N_46814,N_46809);
and U47162 (N_47162,N_46926,N_46942);
nor U47163 (N_47163,N_46945,N_46774);
or U47164 (N_47164,N_46897,N_46876);
nand U47165 (N_47165,N_46860,N_46883);
xor U47166 (N_47166,N_46991,N_46912);
nand U47167 (N_47167,N_46785,N_46895);
nand U47168 (N_47168,N_46998,N_46868);
nand U47169 (N_47169,N_46933,N_46946);
xnor U47170 (N_47170,N_46924,N_46794);
nand U47171 (N_47171,N_46806,N_46988);
and U47172 (N_47172,N_46811,N_46892);
nor U47173 (N_47173,N_46919,N_46805);
and U47174 (N_47174,N_46905,N_46892);
nor U47175 (N_47175,N_46848,N_46956);
nor U47176 (N_47176,N_46951,N_46768);
and U47177 (N_47177,N_46814,N_46836);
nand U47178 (N_47178,N_46846,N_46806);
and U47179 (N_47179,N_46854,N_46762);
or U47180 (N_47180,N_46932,N_46754);
xnor U47181 (N_47181,N_46799,N_46775);
or U47182 (N_47182,N_46783,N_46907);
xor U47183 (N_47183,N_46820,N_46791);
xnor U47184 (N_47184,N_46814,N_46798);
nor U47185 (N_47185,N_46910,N_46803);
nand U47186 (N_47186,N_46818,N_46938);
or U47187 (N_47187,N_46917,N_46989);
xor U47188 (N_47188,N_46824,N_46969);
nand U47189 (N_47189,N_46926,N_46970);
nor U47190 (N_47190,N_46998,N_46980);
nor U47191 (N_47191,N_46814,N_46859);
nand U47192 (N_47192,N_46754,N_46935);
or U47193 (N_47193,N_46949,N_46803);
nand U47194 (N_47194,N_46975,N_46887);
and U47195 (N_47195,N_46983,N_46842);
or U47196 (N_47196,N_46834,N_46848);
nand U47197 (N_47197,N_46905,N_46769);
and U47198 (N_47198,N_46884,N_46822);
nand U47199 (N_47199,N_46984,N_46815);
nand U47200 (N_47200,N_46770,N_46937);
xor U47201 (N_47201,N_46785,N_46942);
or U47202 (N_47202,N_46943,N_46975);
xnor U47203 (N_47203,N_46892,N_46962);
nand U47204 (N_47204,N_46813,N_46947);
and U47205 (N_47205,N_46936,N_46773);
and U47206 (N_47206,N_46867,N_46831);
nor U47207 (N_47207,N_46836,N_46751);
and U47208 (N_47208,N_46937,N_46794);
nand U47209 (N_47209,N_46887,N_46760);
or U47210 (N_47210,N_46898,N_46808);
or U47211 (N_47211,N_46829,N_46947);
or U47212 (N_47212,N_46768,N_46813);
nand U47213 (N_47213,N_46804,N_46755);
xor U47214 (N_47214,N_46963,N_46853);
and U47215 (N_47215,N_46932,N_46874);
nand U47216 (N_47216,N_46983,N_46891);
nor U47217 (N_47217,N_46820,N_46827);
or U47218 (N_47218,N_46834,N_46971);
xnor U47219 (N_47219,N_46895,N_46763);
or U47220 (N_47220,N_46779,N_46981);
xnor U47221 (N_47221,N_46791,N_46814);
or U47222 (N_47222,N_46776,N_46876);
nor U47223 (N_47223,N_46942,N_46939);
xor U47224 (N_47224,N_46755,N_46800);
and U47225 (N_47225,N_46823,N_46833);
nor U47226 (N_47226,N_46866,N_46936);
nand U47227 (N_47227,N_46758,N_46994);
nand U47228 (N_47228,N_46778,N_46896);
or U47229 (N_47229,N_46956,N_46885);
nor U47230 (N_47230,N_46942,N_46953);
xor U47231 (N_47231,N_46852,N_46770);
nor U47232 (N_47232,N_46815,N_46882);
and U47233 (N_47233,N_46797,N_46949);
and U47234 (N_47234,N_46996,N_46753);
xor U47235 (N_47235,N_46830,N_46751);
nor U47236 (N_47236,N_46834,N_46841);
and U47237 (N_47237,N_46991,N_46951);
or U47238 (N_47238,N_46766,N_46931);
and U47239 (N_47239,N_46872,N_46925);
xnor U47240 (N_47240,N_46789,N_46793);
nand U47241 (N_47241,N_46955,N_46893);
or U47242 (N_47242,N_46768,N_46759);
nor U47243 (N_47243,N_46816,N_46912);
nor U47244 (N_47244,N_46776,N_46805);
xnor U47245 (N_47245,N_46974,N_46782);
nand U47246 (N_47246,N_46981,N_46793);
xnor U47247 (N_47247,N_46980,N_46826);
and U47248 (N_47248,N_46952,N_46814);
or U47249 (N_47249,N_46896,N_46963);
nand U47250 (N_47250,N_47248,N_47006);
nor U47251 (N_47251,N_47180,N_47225);
and U47252 (N_47252,N_47005,N_47001);
and U47253 (N_47253,N_47109,N_47030);
and U47254 (N_47254,N_47198,N_47157);
nand U47255 (N_47255,N_47056,N_47012);
xor U47256 (N_47256,N_47127,N_47094);
and U47257 (N_47257,N_47239,N_47107);
nor U47258 (N_47258,N_47151,N_47085);
xor U47259 (N_47259,N_47045,N_47224);
nand U47260 (N_47260,N_47037,N_47172);
xnor U47261 (N_47261,N_47209,N_47115);
or U47262 (N_47262,N_47059,N_47153);
nand U47263 (N_47263,N_47245,N_47110);
xor U47264 (N_47264,N_47167,N_47144);
xor U47265 (N_47265,N_47104,N_47081);
nand U47266 (N_47266,N_47074,N_47228);
nand U47267 (N_47267,N_47114,N_47047);
xor U47268 (N_47268,N_47139,N_47206);
or U47269 (N_47269,N_47022,N_47116);
nor U47270 (N_47270,N_47219,N_47051);
and U47271 (N_47271,N_47147,N_47054);
nand U47272 (N_47272,N_47055,N_47076);
xor U47273 (N_47273,N_47191,N_47243);
and U47274 (N_47274,N_47154,N_47231);
nand U47275 (N_47275,N_47077,N_47038);
nor U47276 (N_47276,N_47003,N_47132);
and U47277 (N_47277,N_47176,N_47020);
nand U47278 (N_47278,N_47100,N_47237);
nor U47279 (N_47279,N_47185,N_47235);
xnor U47280 (N_47280,N_47016,N_47041);
nor U47281 (N_47281,N_47009,N_47194);
or U47282 (N_47282,N_47143,N_47192);
nand U47283 (N_47283,N_47044,N_47145);
nor U47284 (N_47284,N_47092,N_47230);
nand U47285 (N_47285,N_47199,N_47096);
xnor U47286 (N_47286,N_47025,N_47174);
nor U47287 (N_47287,N_47046,N_47148);
nor U47288 (N_47288,N_47029,N_47138);
nand U47289 (N_47289,N_47182,N_47200);
nor U47290 (N_47290,N_47010,N_47043);
nand U47291 (N_47291,N_47164,N_47117);
or U47292 (N_47292,N_47018,N_47213);
nor U47293 (N_47293,N_47238,N_47101);
and U47294 (N_47294,N_47063,N_47031);
and U47295 (N_47295,N_47080,N_47119);
and U47296 (N_47296,N_47024,N_47071);
and U47297 (N_47297,N_47236,N_47083);
and U47298 (N_47298,N_47052,N_47129);
or U47299 (N_47299,N_47134,N_47124);
nor U47300 (N_47300,N_47075,N_47082);
nor U47301 (N_47301,N_47093,N_47216);
and U47302 (N_47302,N_47165,N_47067);
and U47303 (N_47303,N_47208,N_47222);
nand U47304 (N_47304,N_47210,N_47155);
nand U47305 (N_47305,N_47215,N_47152);
and U47306 (N_47306,N_47162,N_47135);
or U47307 (N_47307,N_47220,N_47202);
or U47308 (N_47308,N_47106,N_47068);
or U47309 (N_47309,N_47179,N_47190);
xnor U47310 (N_47310,N_47084,N_47048);
nand U47311 (N_47311,N_47140,N_47049);
and U47312 (N_47312,N_47232,N_47072);
nor U47313 (N_47313,N_47234,N_47150);
nor U47314 (N_47314,N_47008,N_47111);
nand U47315 (N_47315,N_47073,N_47069);
xor U47316 (N_47316,N_47229,N_47189);
nor U47317 (N_47317,N_47136,N_47175);
xnor U47318 (N_47318,N_47122,N_47195);
xnor U47319 (N_47319,N_47181,N_47166);
nand U47320 (N_47320,N_47097,N_47098);
xor U47321 (N_47321,N_47207,N_47099);
nor U47322 (N_47322,N_47177,N_47034);
nand U47323 (N_47323,N_47014,N_47205);
and U47324 (N_47324,N_47214,N_47050);
xnor U47325 (N_47325,N_47168,N_47184);
or U47326 (N_47326,N_47078,N_47170);
nand U47327 (N_47327,N_47217,N_47169);
xnor U47328 (N_47328,N_47105,N_47211);
and U47329 (N_47329,N_47186,N_47171);
nand U47330 (N_47330,N_47201,N_47019);
and U47331 (N_47331,N_47137,N_47108);
or U47332 (N_47332,N_47090,N_47249);
nor U47333 (N_47333,N_47086,N_47026);
or U47334 (N_47334,N_47032,N_47218);
nand U47335 (N_47335,N_47203,N_47027);
xor U47336 (N_47336,N_47028,N_47088);
or U47337 (N_47337,N_47133,N_47146);
and U47338 (N_47338,N_47062,N_47233);
nand U47339 (N_47339,N_47002,N_47053);
or U47340 (N_47340,N_47011,N_47247);
nor U47341 (N_47341,N_47040,N_47130);
nor U47342 (N_47342,N_47188,N_47023);
xor U47343 (N_47343,N_47226,N_47042);
nand U47344 (N_47344,N_47193,N_47121);
and U47345 (N_47345,N_47013,N_47197);
xnor U47346 (N_47346,N_47187,N_47065);
nor U47347 (N_47347,N_47178,N_47033);
and U47348 (N_47348,N_47141,N_47173);
xor U47349 (N_47349,N_47064,N_47123);
nand U47350 (N_47350,N_47183,N_47240);
and U47351 (N_47351,N_47163,N_47125);
and U47352 (N_47352,N_47058,N_47103);
nand U47353 (N_47353,N_47212,N_47036);
nor U47354 (N_47354,N_47223,N_47204);
or U47355 (N_47355,N_47159,N_47087);
and U47356 (N_47356,N_47007,N_47039);
nand U47357 (N_47357,N_47089,N_47079);
nor U47358 (N_47358,N_47221,N_47102);
and U47359 (N_47359,N_47227,N_47149);
or U47360 (N_47360,N_47000,N_47061);
or U47361 (N_47361,N_47241,N_47126);
nor U47362 (N_47362,N_47095,N_47242);
or U47363 (N_47363,N_47196,N_47120);
xnor U47364 (N_47364,N_47244,N_47035);
or U47365 (N_47365,N_47004,N_47017);
xnor U47366 (N_47366,N_47246,N_47057);
xor U47367 (N_47367,N_47160,N_47015);
or U47368 (N_47368,N_47142,N_47066);
or U47369 (N_47369,N_47131,N_47112);
or U47370 (N_47370,N_47091,N_47156);
and U47371 (N_47371,N_47113,N_47118);
nor U47372 (N_47372,N_47158,N_47070);
or U47373 (N_47373,N_47161,N_47060);
or U47374 (N_47374,N_47021,N_47128);
nor U47375 (N_47375,N_47025,N_47149);
nor U47376 (N_47376,N_47107,N_47219);
nor U47377 (N_47377,N_47216,N_47085);
nor U47378 (N_47378,N_47164,N_47023);
and U47379 (N_47379,N_47101,N_47022);
xor U47380 (N_47380,N_47204,N_47149);
or U47381 (N_47381,N_47015,N_47065);
or U47382 (N_47382,N_47169,N_47133);
xor U47383 (N_47383,N_47029,N_47139);
xnor U47384 (N_47384,N_47151,N_47026);
and U47385 (N_47385,N_47191,N_47167);
xor U47386 (N_47386,N_47190,N_47188);
xnor U47387 (N_47387,N_47237,N_47051);
nor U47388 (N_47388,N_47162,N_47059);
nand U47389 (N_47389,N_47151,N_47113);
and U47390 (N_47390,N_47159,N_47038);
or U47391 (N_47391,N_47049,N_47056);
xnor U47392 (N_47392,N_47009,N_47198);
xor U47393 (N_47393,N_47078,N_47165);
nor U47394 (N_47394,N_47016,N_47196);
xnor U47395 (N_47395,N_47057,N_47063);
or U47396 (N_47396,N_47045,N_47098);
nor U47397 (N_47397,N_47021,N_47034);
or U47398 (N_47398,N_47196,N_47195);
xnor U47399 (N_47399,N_47093,N_47083);
nand U47400 (N_47400,N_47119,N_47117);
xor U47401 (N_47401,N_47178,N_47024);
nor U47402 (N_47402,N_47196,N_47249);
xnor U47403 (N_47403,N_47083,N_47151);
nor U47404 (N_47404,N_47172,N_47243);
xor U47405 (N_47405,N_47009,N_47093);
or U47406 (N_47406,N_47229,N_47047);
xnor U47407 (N_47407,N_47036,N_47051);
and U47408 (N_47408,N_47142,N_47063);
nor U47409 (N_47409,N_47128,N_47225);
or U47410 (N_47410,N_47133,N_47102);
nand U47411 (N_47411,N_47083,N_47002);
and U47412 (N_47412,N_47146,N_47194);
nor U47413 (N_47413,N_47053,N_47069);
xor U47414 (N_47414,N_47098,N_47070);
or U47415 (N_47415,N_47212,N_47002);
and U47416 (N_47416,N_47234,N_47223);
nor U47417 (N_47417,N_47019,N_47241);
nor U47418 (N_47418,N_47104,N_47054);
nor U47419 (N_47419,N_47110,N_47105);
xnor U47420 (N_47420,N_47012,N_47036);
or U47421 (N_47421,N_47112,N_47164);
and U47422 (N_47422,N_47101,N_47035);
or U47423 (N_47423,N_47097,N_47113);
nand U47424 (N_47424,N_47144,N_47064);
xor U47425 (N_47425,N_47151,N_47194);
or U47426 (N_47426,N_47083,N_47010);
and U47427 (N_47427,N_47217,N_47204);
nor U47428 (N_47428,N_47060,N_47000);
and U47429 (N_47429,N_47230,N_47125);
and U47430 (N_47430,N_47099,N_47136);
and U47431 (N_47431,N_47102,N_47162);
xnor U47432 (N_47432,N_47107,N_47176);
and U47433 (N_47433,N_47118,N_47112);
or U47434 (N_47434,N_47186,N_47178);
or U47435 (N_47435,N_47156,N_47246);
or U47436 (N_47436,N_47247,N_47228);
nor U47437 (N_47437,N_47053,N_47115);
nor U47438 (N_47438,N_47105,N_47237);
nor U47439 (N_47439,N_47230,N_47099);
nand U47440 (N_47440,N_47097,N_47002);
xor U47441 (N_47441,N_47067,N_47060);
nor U47442 (N_47442,N_47072,N_47067);
nand U47443 (N_47443,N_47132,N_47240);
nor U47444 (N_47444,N_47020,N_47041);
nor U47445 (N_47445,N_47154,N_47172);
and U47446 (N_47446,N_47205,N_47031);
and U47447 (N_47447,N_47111,N_47029);
nor U47448 (N_47448,N_47231,N_47236);
nand U47449 (N_47449,N_47230,N_47088);
nand U47450 (N_47450,N_47062,N_47065);
nand U47451 (N_47451,N_47169,N_47092);
or U47452 (N_47452,N_47200,N_47192);
and U47453 (N_47453,N_47149,N_47016);
or U47454 (N_47454,N_47098,N_47170);
xor U47455 (N_47455,N_47149,N_47100);
and U47456 (N_47456,N_47074,N_47055);
nand U47457 (N_47457,N_47211,N_47104);
and U47458 (N_47458,N_47165,N_47139);
and U47459 (N_47459,N_47089,N_47237);
and U47460 (N_47460,N_47001,N_47046);
nor U47461 (N_47461,N_47139,N_47083);
xnor U47462 (N_47462,N_47084,N_47180);
nor U47463 (N_47463,N_47071,N_47116);
nor U47464 (N_47464,N_47232,N_47115);
nor U47465 (N_47465,N_47158,N_47188);
and U47466 (N_47466,N_47103,N_47150);
nor U47467 (N_47467,N_47189,N_47051);
and U47468 (N_47468,N_47084,N_47230);
or U47469 (N_47469,N_47210,N_47227);
nor U47470 (N_47470,N_47137,N_47035);
or U47471 (N_47471,N_47087,N_47108);
nand U47472 (N_47472,N_47070,N_47009);
nor U47473 (N_47473,N_47054,N_47237);
nor U47474 (N_47474,N_47151,N_47139);
and U47475 (N_47475,N_47220,N_47033);
or U47476 (N_47476,N_47144,N_47171);
and U47477 (N_47477,N_47019,N_47088);
nor U47478 (N_47478,N_47046,N_47232);
or U47479 (N_47479,N_47106,N_47238);
nand U47480 (N_47480,N_47159,N_47221);
and U47481 (N_47481,N_47084,N_47003);
or U47482 (N_47482,N_47214,N_47144);
nor U47483 (N_47483,N_47072,N_47214);
nand U47484 (N_47484,N_47033,N_47051);
or U47485 (N_47485,N_47005,N_47026);
xnor U47486 (N_47486,N_47057,N_47182);
xor U47487 (N_47487,N_47080,N_47168);
nand U47488 (N_47488,N_47026,N_47176);
xnor U47489 (N_47489,N_47241,N_47101);
or U47490 (N_47490,N_47159,N_47203);
nand U47491 (N_47491,N_47179,N_47003);
nand U47492 (N_47492,N_47188,N_47124);
and U47493 (N_47493,N_47221,N_47076);
nand U47494 (N_47494,N_47157,N_47118);
or U47495 (N_47495,N_47076,N_47162);
nand U47496 (N_47496,N_47248,N_47117);
nor U47497 (N_47497,N_47176,N_47198);
or U47498 (N_47498,N_47098,N_47151);
nor U47499 (N_47499,N_47208,N_47233);
xor U47500 (N_47500,N_47262,N_47429);
nor U47501 (N_47501,N_47255,N_47287);
nor U47502 (N_47502,N_47407,N_47288);
nand U47503 (N_47503,N_47486,N_47479);
nor U47504 (N_47504,N_47430,N_47369);
or U47505 (N_47505,N_47379,N_47415);
nor U47506 (N_47506,N_47483,N_47421);
or U47507 (N_47507,N_47260,N_47375);
nor U47508 (N_47508,N_47391,N_47378);
nor U47509 (N_47509,N_47400,N_47303);
xor U47510 (N_47510,N_47385,N_47322);
nor U47511 (N_47511,N_47296,N_47371);
xor U47512 (N_47512,N_47336,N_47282);
and U47513 (N_47513,N_47317,N_47291);
and U47514 (N_47514,N_47398,N_47320);
xor U47515 (N_47515,N_47356,N_47332);
nand U47516 (N_47516,N_47498,N_47493);
nor U47517 (N_47517,N_47406,N_47267);
and U47518 (N_47518,N_47402,N_47269);
and U47519 (N_47519,N_47372,N_47456);
and U47520 (N_47520,N_47444,N_47339);
nor U47521 (N_47521,N_47341,N_47480);
and U47522 (N_47522,N_47422,N_47273);
or U47523 (N_47523,N_47284,N_47266);
nor U47524 (N_47524,N_47350,N_47495);
or U47525 (N_47525,N_47488,N_47411);
xor U47526 (N_47526,N_47366,N_47474);
or U47527 (N_47527,N_47481,N_47251);
and U47528 (N_47528,N_47397,N_47252);
xor U47529 (N_47529,N_47327,N_47263);
xnor U47530 (N_47530,N_47308,N_47264);
xor U47531 (N_47531,N_47404,N_47302);
nor U47532 (N_47532,N_47340,N_47329);
and U47533 (N_47533,N_47470,N_47399);
xor U47534 (N_47534,N_47275,N_47448);
nor U47535 (N_47535,N_47443,N_47394);
and U47536 (N_47536,N_47294,N_47360);
xnor U47537 (N_47537,N_47463,N_47405);
and U47538 (N_47538,N_47442,N_47484);
or U47539 (N_47539,N_47307,N_47491);
nor U47540 (N_47540,N_47281,N_47330);
xor U47541 (N_47541,N_47487,N_47439);
xor U47542 (N_47542,N_47344,N_47462);
nand U47543 (N_47543,N_47457,N_47349);
nand U47544 (N_47544,N_47318,N_47426);
nor U47545 (N_47545,N_47335,N_47297);
nand U47546 (N_47546,N_47300,N_47359);
xor U47547 (N_47547,N_47445,N_47496);
xnor U47548 (N_47548,N_47272,N_47253);
xnor U47549 (N_47549,N_47265,N_47433);
nand U47550 (N_47550,N_47290,N_47475);
nor U47551 (N_47551,N_47434,N_47295);
nor U47552 (N_47552,N_47388,N_47380);
nor U47553 (N_47553,N_47353,N_47467);
nand U47554 (N_47554,N_47293,N_47315);
or U47555 (N_47555,N_47271,N_47348);
nand U47556 (N_47556,N_47384,N_47321);
xor U47557 (N_47557,N_47280,N_47499);
or U47558 (N_47558,N_47468,N_47323);
or U47559 (N_47559,N_47314,N_47452);
xor U47560 (N_47560,N_47390,N_47345);
nor U47561 (N_47561,N_47497,N_47438);
nor U47562 (N_47562,N_47392,N_47283);
nand U47563 (N_47563,N_47424,N_47373);
or U47564 (N_47564,N_47403,N_47285);
and U47565 (N_47565,N_47432,N_47367);
and U47566 (N_47566,N_47370,N_47277);
nand U47567 (N_47567,N_47408,N_47358);
or U47568 (N_47568,N_47446,N_47286);
nor U47569 (N_47569,N_47450,N_47482);
nand U47570 (N_47570,N_47436,N_47449);
nand U47571 (N_47571,N_47361,N_47472);
xnor U47572 (N_47572,N_47417,N_47374);
or U47573 (N_47573,N_47478,N_47362);
nor U47574 (N_47574,N_47453,N_47250);
and U47575 (N_47575,N_47412,N_47469);
nand U47576 (N_47576,N_47276,N_47324);
xor U47577 (N_47577,N_47337,N_47334);
and U47578 (N_47578,N_47428,N_47455);
nand U47579 (N_47579,N_47427,N_47425);
and U47580 (N_47580,N_47414,N_47257);
and U47581 (N_47581,N_47325,N_47363);
xor U47582 (N_47582,N_47461,N_47313);
xor U47583 (N_47583,N_47351,N_47395);
xor U47584 (N_47584,N_47459,N_47460);
nand U47585 (N_47585,N_47458,N_47298);
and U47586 (N_47586,N_47376,N_47401);
xor U47587 (N_47587,N_47274,N_47454);
or U47588 (N_47588,N_47268,N_47471);
and U47589 (N_47589,N_47368,N_47310);
and U47590 (N_47590,N_47473,N_47346);
nor U47591 (N_47591,N_47355,N_47333);
nand U47592 (N_47592,N_47347,N_47387);
nor U47593 (N_47593,N_47466,N_47354);
or U47594 (N_47594,N_47309,N_47259);
nand U47595 (N_47595,N_47440,N_47338);
xor U47596 (N_47596,N_47447,N_47492);
and U47597 (N_47597,N_47476,N_47365);
nor U47598 (N_47598,N_47494,N_47256);
or U47599 (N_47599,N_47328,N_47410);
nor U47600 (N_47600,N_47301,N_47357);
nor U47601 (N_47601,N_47416,N_47396);
nor U47602 (N_47602,N_47413,N_47258);
xnor U47603 (N_47603,N_47254,N_47431);
xnor U47604 (N_47604,N_47312,N_47377);
or U47605 (N_47605,N_47299,N_47331);
nor U47606 (N_47606,N_47420,N_47465);
xnor U47607 (N_47607,N_47326,N_47489);
xnor U47608 (N_47608,N_47304,N_47393);
or U47609 (N_47609,N_47477,N_47279);
nand U47610 (N_47610,N_47386,N_47278);
nand U47611 (N_47611,N_47261,N_47451);
or U47612 (N_47612,N_47485,N_47437);
or U47613 (N_47613,N_47306,N_47409);
nor U47614 (N_47614,N_47441,N_47292);
nand U47615 (N_47615,N_47382,N_47342);
nor U47616 (N_47616,N_47364,N_47381);
xor U47617 (N_47617,N_47418,N_47316);
or U47618 (N_47618,N_47305,N_47389);
xnor U47619 (N_47619,N_47270,N_47343);
xnor U47620 (N_47620,N_47435,N_47352);
nor U47621 (N_47621,N_47383,N_47419);
nor U47622 (N_47622,N_47423,N_47319);
or U47623 (N_47623,N_47311,N_47490);
nand U47624 (N_47624,N_47289,N_47464);
and U47625 (N_47625,N_47404,N_47306);
or U47626 (N_47626,N_47414,N_47411);
and U47627 (N_47627,N_47478,N_47394);
nand U47628 (N_47628,N_47404,N_47304);
and U47629 (N_47629,N_47306,N_47471);
or U47630 (N_47630,N_47379,N_47307);
or U47631 (N_47631,N_47393,N_47441);
nand U47632 (N_47632,N_47445,N_47418);
or U47633 (N_47633,N_47267,N_47470);
xor U47634 (N_47634,N_47366,N_47450);
nor U47635 (N_47635,N_47374,N_47293);
or U47636 (N_47636,N_47437,N_47463);
xor U47637 (N_47637,N_47330,N_47416);
nor U47638 (N_47638,N_47252,N_47255);
nand U47639 (N_47639,N_47484,N_47370);
nand U47640 (N_47640,N_47456,N_47450);
and U47641 (N_47641,N_47407,N_47259);
nor U47642 (N_47642,N_47262,N_47482);
nor U47643 (N_47643,N_47317,N_47305);
or U47644 (N_47644,N_47331,N_47398);
xnor U47645 (N_47645,N_47317,N_47324);
or U47646 (N_47646,N_47378,N_47363);
nor U47647 (N_47647,N_47451,N_47443);
xor U47648 (N_47648,N_47446,N_47292);
nand U47649 (N_47649,N_47430,N_47441);
or U47650 (N_47650,N_47314,N_47360);
and U47651 (N_47651,N_47473,N_47421);
nor U47652 (N_47652,N_47264,N_47378);
nand U47653 (N_47653,N_47323,N_47273);
or U47654 (N_47654,N_47290,N_47319);
nor U47655 (N_47655,N_47371,N_47378);
or U47656 (N_47656,N_47376,N_47463);
nand U47657 (N_47657,N_47499,N_47362);
or U47658 (N_47658,N_47294,N_47270);
nor U47659 (N_47659,N_47265,N_47271);
and U47660 (N_47660,N_47337,N_47415);
or U47661 (N_47661,N_47476,N_47357);
and U47662 (N_47662,N_47412,N_47475);
and U47663 (N_47663,N_47264,N_47437);
or U47664 (N_47664,N_47394,N_47297);
and U47665 (N_47665,N_47339,N_47492);
xor U47666 (N_47666,N_47284,N_47352);
and U47667 (N_47667,N_47440,N_47299);
and U47668 (N_47668,N_47314,N_47286);
or U47669 (N_47669,N_47494,N_47363);
or U47670 (N_47670,N_47257,N_47405);
and U47671 (N_47671,N_47412,N_47396);
xnor U47672 (N_47672,N_47380,N_47492);
nand U47673 (N_47673,N_47251,N_47472);
and U47674 (N_47674,N_47328,N_47464);
nor U47675 (N_47675,N_47279,N_47397);
xnor U47676 (N_47676,N_47448,N_47407);
nand U47677 (N_47677,N_47251,N_47354);
nand U47678 (N_47678,N_47468,N_47311);
nand U47679 (N_47679,N_47321,N_47463);
or U47680 (N_47680,N_47300,N_47302);
xor U47681 (N_47681,N_47430,N_47498);
and U47682 (N_47682,N_47469,N_47377);
or U47683 (N_47683,N_47385,N_47374);
nand U47684 (N_47684,N_47372,N_47358);
and U47685 (N_47685,N_47359,N_47355);
xnor U47686 (N_47686,N_47289,N_47273);
nand U47687 (N_47687,N_47259,N_47276);
and U47688 (N_47688,N_47323,N_47471);
or U47689 (N_47689,N_47262,N_47264);
or U47690 (N_47690,N_47328,N_47330);
or U47691 (N_47691,N_47303,N_47263);
xnor U47692 (N_47692,N_47352,N_47318);
or U47693 (N_47693,N_47354,N_47323);
and U47694 (N_47694,N_47376,N_47406);
nand U47695 (N_47695,N_47438,N_47297);
and U47696 (N_47696,N_47289,N_47379);
and U47697 (N_47697,N_47296,N_47260);
and U47698 (N_47698,N_47362,N_47320);
and U47699 (N_47699,N_47472,N_47318);
nand U47700 (N_47700,N_47426,N_47413);
and U47701 (N_47701,N_47331,N_47316);
or U47702 (N_47702,N_47482,N_47471);
nor U47703 (N_47703,N_47305,N_47394);
or U47704 (N_47704,N_47440,N_47410);
nand U47705 (N_47705,N_47299,N_47492);
and U47706 (N_47706,N_47494,N_47394);
xnor U47707 (N_47707,N_47469,N_47259);
nor U47708 (N_47708,N_47366,N_47260);
and U47709 (N_47709,N_47343,N_47372);
xor U47710 (N_47710,N_47487,N_47288);
nor U47711 (N_47711,N_47258,N_47468);
nor U47712 (N_47712,N_47269,N_47274);
nor U47713 (N_47713,N_47371,N_47403);
and U47714 (N_47714,N_47291,N_47347);
and U47715 (N_47715,N_47326,N_47486);
or U47716 (N_47716,N_47376,N_47331);
nand U47717 (N_47717,N_47491,N_47250);
nand U47718 (N_47718,N_47423,N_47403);
or U47719 (N_47719,N_47456,N_47319);
nand U47720 (N_47720,N_47352,N_47386);
nor U47721 (N_47721,N_47417,N_47398);
and U47722 (N_47722,N_47358,N_47478);
and U47723 (N_47723,N_47317,N_47253);
nand U47724 (N_47724,N_47395,N_47274);
xnor U47725 (N_47725,N_47394,N_47401);
nor U47726 (N_47726,N_47424,N_47419);
nand U47727 (N_47727,N_47457,N_47490);
and U47728 (N_47728,N_47270,N_47325);
or U47729 (N_47729,N_47396,N_47299);
nor U47730 (N_47730,N_47379,N_47420);
nand U47731 (N_47731,N_47289,N_47311);
nor U47732 (N_47732,N_47292,N_47295);
xor U47733 (N_47733,N_47311,N_47432);
and U47734 (N_47734,N_47333,N_47278);
and U47735 (N_47735,N_47371,N_47458);
and U47736 (N_47736,N_47445,N_47477);
and U47737 (N_47737,N_47434,N_47269);
or U47738 (N_47738,N_47429,N_47316);
and U47739 (N_47739,N_47380,N_47478);
or U47740 (N_47740,N_47306,N_47377);
xor U47741 (N_47741,N_47355,N_47351);
nor U47742 (N_47742,N_47345,N_47365);
and U47743 (N_47743,N_47351,N_47309);
nor U47744 (N_47744,N_47440,N_47298);
or U47745 (N_47745,N_47266,N_47451);
and U47746 (N_47746,N_47466,N_47398);
or U47747 (N_47747,N_47288,N_47499);
nand U47748 (N_47748,N_47257,N_47358);
nand U47749 (N_47749,N_47277,N_47499);
or U47750 (N_47750,N_47589,N_47603);
or U47751 (N_47751,N_47745,N_47680);
and U47752 (N_47752,N_47531,N_47575);
or U47753 (N_47753,N_47585,N_47558);
or U47754 (N_47754,N_47631,N_47650);
xnor U47755 (N_47755,N_47696,N_47678);
or U47756 (N_47756,N_47547,N_47605);
xnor U47757 (N_47757,N_47746,N_47566);
xnor U47758 (N_47758,N_47526,N_47702);
or U47759 (N_47759,N_47685,N_47601);
or U47760 (N_47760,N_47712,N_47738);
nor U47761 (N_47761,N_47710,N_47659);
and U47762 (N_47762,N_47512,N_47607);
nand U47763 (N_47763,N_47509,N_47546);
nor U47764 (N_47764,N_47731,N_47513);
or U47765 (N_47765,N_47724,N_47540);
and U47766 (N_47766,N_47682,N_47639);
nor U47767 (N_47767,N_47728,N_47528);
or U47768 (N_47768,N_47611,N_47642);
xnor U47769 (N_47769,N_47576,N_47584);
nand U47770 (N_47770,N_47637,N_47583);
nand U47771 (N_47771,N_47523,N_47617);
nand U47772 (N_47772,N_47560,N_47687);
nor U47773 (N_47773,N_47552,N_47729);
nand U47774 (N_47774,N_47630,N_47638);
or U47775 (N_47775,N_47660,N_47532);
nor U47776 (N_47776,N_47634,N_47569);
xor U47777 (N_47777,N_47635,N_47608);
nor U47778 (N_47778,N_47591,N_47570);
xnor U47779 (N_47779,N_47725,N_47747);
and U47780 (N_47780,N_47507,N_47657);
xor U47781 (N_47781,N_47735,N_47707);
nor U47782 (N_47782,N_47694,N_47614);
xor U47783 (N_47783,N_47730,N_47538);
and U47784 (N_47784,N_47664,N_47711);
or U47785 (N_47785,N_47612,N_47633);
nand U47786 (N_47786,N_47697,N_47740);
and U47787 (N_47787,N_47718,N_47628);
nand U47788 (N_47788,N_47555,N_47717);
nand U47789 (N_47789,N_47535,N_47530);
nand U47790 (N_47790,N_47652,N_47503);
xnor U47791 (N_47791,N_47577,N_47520);
or U47792 (N_47792,N_47596,N_47534);
xnor U47793 (N_47793,N_47529,N_47599);
nand U47794 (N_47794,N_47699,N_47594);
or U47795 (N_47795,N_47705,N_47582);
or U47796 (N_47796,N_47501,N_47537);
nand U47797 (N_47797,N_47624,N_47713);
or U47798 (N_47798,N_47504,N_47675);
nand U47799 (N_47799,N_47654,N_47616);
or U47800 (N_47800,N_47506,N_47684);
and U47801 (N_47801,N_47500,N_47693);
or U47802 (N_47802,N_47743,N_47627);
or U47803 (N_47803,N_47598,N_47539);
nand U47804 (N_47804,N_47604,N_47622);
or U47805 (N_47805,N_47602,N_47597);
nor U47806 (N_47806,N_47579,N_47609);
xnor U47807 (N_47807,N_47514,N_47715);
nor U47808 (N_47808,N_47681,N_47714);
or U47809 (N_47809,N_47703,N_47700);
and U47810 (N_47810,N_47742,N_47571);
and U47811 (N_47811,N_47722,N_47510);
xor U47812 (N_47812,N_47556,N_47688);
xor U47813 (N_47813,N_47677,N_47647);
nand U47814 (N_47814,N_47665,N_47698);
nor U47815 (N_47815,N_47643,N_47648);
nor U47816 (N_47816,N_47661,N_47586);
or U47817 (N_47817,N_47541,N_47690);
nor U47818 (N_47818,N_47545,N_47610);
nor U47819 (N_47819,N_47587,N_47739);
or U47820 (N_47820,N_47533,N_47590);
xor U47821 (N_47821,N_47606,N_47691);
nor U47822 (N_47822,N_47559,N_47595);
and U47823 (N_47823,N_47625,N_47706);
nand U47824 (N_47824,N_47557,N_47658);
or U47825 (N_47825,N_47508,N_47679);
xnor U47826 (N_47826,N_47549,N_47502);
nand U47827 (N_47827,N_47709,N_47553);
and U47828 (N_47828,N_47588,N_47673);
and U47829 (N_47829,N_47593,N_47734);
nor U47830 (N_47830,N_47723,N_47686);
and U47831 (N_47831,N_47737,N_47720);
or U47832 (N_47832,N_47667,N_47732);
nand U47833 (N_47833,N_47581,N_47568);
nor U47834 (N_47834,N_47562,N_47613);
or U47835 (N_47835,N_47719,N_47561);
nand U47836 (N_47836,N_47662,N_47550);
and U47837 (N_47837,N_47736,N_47708);
nand U47838 (N_47838,N_47542,N_47640);
and U47839 (N_47839,N_47641,N_47521);
or U47840 (N_47840,N_47565,N_47692);
xor U47841 (N_47841,N_47656,N_47676);
and U47842 (N_47842,N_47668,N_47551);
or U47843 (N_47843,N_47563,N_47600);
or U47844 (N_47844,N_47518,N_47619);
and U47845 (N_47845,N_47716,N_47554);
or U47846 (N_47846,N_47623,N_47592);
and U47847 (N_47847,N_47567,N_47727);
or U47848 (N_47848,N_47525,N_47663);
and U47849 (N_47849,N_47516,N_47651);
nand U47850 (N_47850,N_47701,N_47536);
nand U47851 (N_47851,N_47683,N_47618);
or U47852 (N_47852,N_47519,N_47649);
nor U47853 (N_47853,N_47666,N_47749);
nor U47854 (N_47854,N_47741,N_47572);
xnor U47855 (N_47855,N_47669,N_47644);
nor U47856 (N_47856,N_47629,N_47524);
or U47857 (N_47857,N_47670,N_47653);
xor U47858 (N_47858,N_47674,N_47574);
nand U47859 (N_47859,N_47548,N_47748);
xor U47860 (N_47860,N_47626,N_47621);
nor U47861 (N_47861,N_47515,N_47580);
nor U47862 (N_47862,N_47511,N_47695);
nor U47863 (N_47863,N_47721,N_47544);
xor U47864 (N_47864,N_47505,N_47578);
nand U47865 (N_47865,N_47527,N_47615);
xor U47866 (N_47866,N_47645,N_47517);
nand U47867 (N_47867,N_47672,N_47620);
or U47868 (N_47868,N_47744,N_47655);
nand U47869 (N_47869,N_47704,N_47646);
or U47870 (N_47870,N_47733,N_47632);
and U47871 (N_47871,N_47689,N_47573);
or U47872 (N_47872,N_47636,N_47564);
and U47873 (N_47873,N_47543,N_47522);
nor U47874 (N_47874,N_47671,N_47726);
and U47875 (N_47875,N_47738,N_47507);
nand U47876 (N_47876,N_47596,N_47671);
nand U47877 (N_47877,N_47599,N_47631);
xnor U47878 (N_47878,N_47544,N_47531);
nand U47879 (N_47879,N_47528,N_47627);
nand U47880 (N_47880,N_47737,N_47517);
xnor U47881 (N_47881,N_47506,N_47569);
or U47882 (N_47882,N_47730,N_47592);
and U47883 (N_47883,N_47640,N_47661);
nand U47884 (N_47884,N_47545,N_47635);
nand U47885 (N_47885,N_47572,N_47612);
nor U47886 (N_47886,N_47706,N_47508);
xor U47887 (N_47887,N_47653,N_47700);
and U47888 (N_47888,N_47614,N_47737);
nand U47889 (N_47889,N_47691,N_47571);
nand U47890 (N_47890,N_47667,N_47614);
nor U47891 (N_47891,N_47589,N_47662);
nand U47892 (N_47892,N_47655,N_47687);
xor U47893 (N_47893,N_47743,N_47729);
nand U47894 (N_47894,N_47732,N_47639);
nor U47895 (N_47895,N_47577,N_47612);
and U47896 (N_47896,N_47711,N_47616);
or U47897 (N_47897,N_47663,N_47740);
or U47898 (N_47898,N_47571,N_47594);
and U47899 (N_47899,N_47551,N_47675);
or U47900 (N_47900,N_47618,N_47635);
nand U47901 (N_47901,N_47627,N_47554);
and U47902 (N_47902,N_47517,N_47709);
and U47903 (N_47903,N_47535,N_47511);
or U47904 (N_47904,N_47588,N_47708);
and U47905 (N_47905,N_47519,N_47563);
nor U47906 (N_47906,N_47630,N_47525);
nor U47907 (N_47907,N_47507,N_47649);
and U47908 (N_47908,N_47524,N_47627);
xor U47909 (N_47909,N_47713,N_47634);
and U47910 (N_47910,N_47585,N_47612);
xor U47911 (N_47911,N_47731,N_47559);
and U47912 (N_47912,N_47670,N_47512);
or U47913 (N_47913,N_47687,N_47624);
and U47914 (N_47914,N_47502,N_47629);
nor U47915 (N_47915,N_47712,N_47628);
xnor U47916 (N_47916,N_47622,N_47629);
and U47917 (N_47917,N_47682,N_47705);
xnor U47918 (N_47918,N_47645,N_47552);
xnor U47919 (N_47919,N_47564,N_47523);
nor U47920 (N_47920,N_47742,N_47659);
and U47921 (N_47921,N_47542,N_47732);
or U47922 (N_47922,N_47690,N_47688);
nand U47923 (N_47923,N_47581,N_47596);
nand U47924 (N_47924,N_47588,N_47580);
or U47925 (N_47925,N_47685,N_47513);
and U47926 (N_47926,N_47559,N_47509);
xnor U47927 (N_47927,N_47565,N_47725);
or U47928 (N_47928,N_47596,N_47625);
or U47929 (N_47929,N_47735,N_47507);
nor U47930 (N_47930,N_47719,N_47603);
nor U47931 (N_47931,N_47589,N_47687);
xor U47932 (N_47932,N_47574,N_47520);
xnor U47933 (N_47933,N_47533,N_47545);
xnor U47934 (N_47934,N_47622,N_47619);
and U47935 (N_47935,N_47566,N_47515);
nor U47936 (N_47936,N_47726,N_47738);
and U47937 (N_47937,N_47677,N_47603);
and U47938 (N_47938,N_47637,N_47709);
nand U47939 (N_47939,N_47661,N_47559);
and U47940 (N_47940,N_47740,N_47675);
or U47941 (N_47941,N_47730,N_47603);
nand U47942 (N_47942,N_47502,N_47737);
nand U47943 (N_47943,N_47687,N_47512);
and U47944 (N_47944,N_47697,N_47581);
or U47945 (N_47945,N_47743,N_47736);
and U47946 (N_47946,N_47681,N_47509);
nor U47947 (N_47947,N_47651,N_47553);
nor U47948 (N_47948,N_47538,N_47512);
nand U47949 (N_47949,N_47722,N_47690);
or U47950 (N_47950,N_47667,N_47549);
or U47951 (N_47951,N_47700,N_47685);
nand U47952 (N_47952,N_47619,N_47749);
or U47953 (N_47953,N_47513,N_47676);
and U47954 (N_47954,N_47645,N_47534);
or U47955 (N_47955,N_47690,N_47713);
nor U47956 (N_47956,N_47533,N_47517);
nor U47957 (N_47957,N_47617,N_47682);
or U47958 (N_47958,N_47720,N_47733);
nor U47959 (N_47959,N_47536,N_47719);
and U47960 (N_47960,N_47709,N_47621);
and U47961 (N_47961,N_47576,N_47648);
and U47962 (N_47962,N_47617,N_47637);
nand U47963 (N_47963,N_47710,N_47645);
xnor U47964 (N_47964,N_47589,N_47546);
nor U47965 (N_47965,N_47742,N_47654);
nor U47966 (N_47966,N_47579,N_47602);
xor U47967 (N_47967,N_47719,N_47569);
nor U47968 (N_47968,N_47706,N_47522);
and U47969 (N_47969,N_47666,N_47542);
and U47970 (N_47970,N_47514,N_47619);
or U47971 (N_47971,N_47538,N_47724);
nand U47972 (N_47972,N_47531,N_47628);
and U47973 (N_47973,N_47688,N_47739);
xnor U47974 (N_47974,N_47728,N_47658);
and U47975 (N_47975,N_47667,N_47711);
xnor U47976 (N_47976,N_47715,N_47524);
and U47977 (N_47977,N_47565,N_47594);
nor U47978 (N_47978,N_47523,N_47689);
and U47979 (N_47979,N_47514,N_47504);
nand U47980 (N_47980,N_47735,N_47684);
nor U47981 (N_47981,N_47679,N_47506);
nor U47982 (N_47982,N_47505,N_47695);
nand U47983 (N_47983,N_47713,N_47665);
or U47984 (N_47984,N_47533,N_47587);
nand U47985 (N_47985,N_47539,N_47604);
nand U47986 (N_47986,N_47743,N_47669);
xnor U47987 (N_47987,N_47747,N_47718);
or U47988 (N_47988,N_47542,N_47506);
xor U47989 (N_47989,N_47688,N_47543);
xor U47990 (N_47990,N_47722,N_47575);
and U47991 (N_47991,N_47680,N_47627);
nor U47992 (N_47992,N_47543,N_47735);
nor U47993 (N_47993,N_47622,N_47714);
nor U47994 (N_47994,N_47575,N_47671);
or U47995 (N_47995,N_47625,N_47684);
nor U47996 (N_47996,N_47650,N_47592);
or U47997 (N_47997,N_47725,N_47676);
and U47998 (N_47998,N_47681,N_47654);
and U47999 (N_47999,N_47584,N_47666);
and U48000 (N_48000,N_47842,N_47761);
and U48001 (N_48001,N_47918,N_47792);
nor U48002 (N_48002,N_47795,N_47836);
and U48003 (N_48003,N_47862,N_47932);
nor U48004 (N_48004,N_47951,N_47967);
xnor U48005 (N_48005,N_47944,N_47999);
nand U48006 (N_48006,N_47764,N_47930);
nor U48007 (N_48007,N_47876,N_47911);
nor U48008 (N_48008,N_47898,N_47858);
or U48009 (N_48009,N_47996,N_47960);
nand U48010 (N_48010,N_47859,N_47760);
xor U48011 (N_48011,N_47936,N_47756);
nand U48012 (N_48012,N_47916,N_47846);
and U48013 (N_48013,N_47841,N_47924);
xor U48014 (N_48014,N_47750,N_47907);
and U48015 (N_48015,N_47820,N_47892);
xor U48016 (N_48016,N_47801,N_47905);
xnor U48017 (N_48017,N_47782,N_47803);
nand U48018 (N_48018,N_47853,N_47894);
nor U48019 (N_48019,N_47783,N_47948);
nor U48020 (N_48020,N_47827,N_47775);
xor U48021 (N_48021,N_47947,N_47763);
or U48022 (N_48022,N_47772,N_47903);
or U48023 (N_48023,N_47909,N_47881);
and U48024 (N_48024,N_47840,N_47878);
or U48025 (N_48025,N_47856,N_47785);
nand U48026 (N_48026,N_47987,N_47794);
xnor U48027 (N_48027,N_47904,N_47824);
or U48028 (N_48028,N_47786,N_47755);
nor U48029 (N_48029,N_47979,N_47938);
and U48030 (N_48030,N_47995,N_47864);
xor U48031 (N_48031,N_47828,N_47754);
or U48032 (N_48032,N_47971,N_47757);
or U48033 (N_48033,N_47880,N_47810);
xnor U48034 (N_48034,N_47983,N_47867);
nor U48035 (N_48035,N_47869,N_47807);
or U48036 (N_48036,N_47788,N_47900);
nand U48037 (N_48037,N_47844,N_47787);
nand U48038 (N_48038,N_47839,N_47920);
xor U48039 (N_48039,N_47848,N_47861);
xor U48040 (N_48040,N_47774,N_47950);
or U48041 (N_48041,N_47789,N_47857);
nor U48042 (N_48042,N_47797,N_47809);
nand U48043 (N_48043,N_47834,N_47925);
or U48044 (N_48044,N_47891,N_47934);
xnor U48045 (N_48045,N_47994,N_47997);
nand U48046 (N_48046,N_47959,N_47890);
and U48047 (N_48047,N_47769,N_47850);
or U48048 (N_48048,N_47957,N_47854);
nor U48049 (N_48049,N_47865,N_47779);
nand U48050 (N_48050,N_47781,N_47833);
or U48051 (N_48051,N_47902,N_47768);
or U48052 (N_48052,N_47819,N_47991);
nor U48053 (N_48053,N_47816,N_47884);
nor U48054 (N_48054,N_47949,N_47956);
nor U48055 (N_48055,N_47993,N_47863);
nor U48056 (N_48056,N_47778,N_47897);
or U48057 (N_48057,N_47955,N_47855);
nand U48058 (N_48058,N_47968,N_47998);
or U48059 (N_48059,N_47912,N_47910);
and U48060 (N_48060,N_47838,N_47917);
or U48061 (N_48061,N_47899,N_47766);
xnor U48062 (N_48062,N_47817,N_47988);
or U48063 (N_48063,N_47751,N_47939);
nor U48064 (N_48064,N_47821,N_47847);
or U48065 (N_48065,N_47926,N_47978);
nand U48066 (N_48066,N_47874,N_47931);
nor U48067 (N_48067,N_47770,N_47826);
xor U48068 (N_48068,N_47776,N_47849);
or U48069 (N_48069,N_47753,N_47919);
nand U48070 (N_48070,N_47972,N_47800);
xnor U48071 (N_48071,N_47812,N_47954);
and U48072 (N_48072,N_47773,N_47831);
and U48073 (N_48073,N_47870,N_47806);
nor U48074 (N_48074,N_47829,N_47771);
or U48075 (N_48075,N_47875,N_47977);
or U48076 (N_48076,N_47990,N_47941);
or U48077 (N_48077,N_47958,N_47837);
and U48078 (N_48078,N_47922,N_47966);
nor U48079 (N_48079,N_47946,N_47992);
or U48080 (N_48080,N_47893,N_47798);
nor U48081 (N_48081,N_47935,N_47866);
nand U48082 (N_48082,N_47942,N_47943);
and U48083 (N_48083,N_47981,N_47835);
nand U48084 (N_48084,N_47882,N_47815);
xor U48085 (N_48085,N_47928,N_47762);
nor U48086 (N_48086,N_47872,N_47962);
xor U48087 (N_48087,N_47984,N_47982);
or U48088 (N_48088,N_47964,N_47906);
nor U48089 (N_48089,N_47752,N_47961);
or U48090 (N_48090,N_47963,N_47885);
nor U48091 (N_48091,N_47965,N_47860);
or U48092 (N_48092,N_47940,N_47868);
and U48093 (N_48093,N_47808,N_47901);
nand U48094 (N_48094,N_47818,N_47843);
or U48095 (N_48095,N_47896,N_47851);
and U48096 (N_48096,N_47871,N_47758);
or U48097 (N_48097,N_47780,N_47980);
nand U48098 (N_48098,N_47879,N_47927);
xnor U48099 (N_48099,N_47759,N_47790);
xnor U48100 (N_48100,N_47873,N_47793);
nor U48101 (N_48101,N_47945,N_47830);
nand U48102 (N_48102,N_47802,N_47814);
xnor U48103 (N_48103,N_47986,N_47952);
nor U48104 (N_48104,N_47832,N_47895);
xnor U48105 (N_48105,N_47813,N_47976);
xor U48106 (N_48106,N_47974,N_47908);
nand U48107 (N_48107,N_47929,N_47886);
and U48108 (N_48108,N_47985,N_47845);
or U48109 (N_48109,N_47888,N_47914);
or U48110 (N_48110,N_47953,N_47805);
and U48111 (N_48111,N_47825,N_47989);
nor U48112 (N_48112,N_47975,N_47765);
and U48113 (N_48113,N_47811,N_47877);
and U48114 (N_48114,N_47852,N_47889);
nor U48115 (N_48115,N_47767,N_47883);
xor U48116 (N_48116,N_47791,N_47784);
or U48117 (N_48117,N_47823,N_47887);
nand U48118 (N_48118,N_47915,N_47796);
xor U48119 (N_48119,N_47804,N_47933);
xor U48120 (N_48120,N_47970,N_47822);
nor U48121 (N_48121,N_47777,N_47921);
or U48122 (N_48122,N_47973,N_47969);
and U48123 (N_48123,N_47923,N_47799);
nor U48124 (N_48124,N_47913,N_47937);
xor U48125 (N_48125,N_47838,N_47980);
and U48126 (N_48126,N_47951,N_47921);
xor U48127 (N_48127,N_47880,N_47921);
xor U48128 (N_48128,N_47831,N_47895);
or U48129 (N_48129,N_47820,N_47985);
and U48130 (N_48130,N_47973,N_47904);
and U48131 (N_48131,N_47937,N_47895);
or U48132 (N_48132,N_47976,N_47824);
nor U48133 (N_48133,N_47862,N_47757);
and U48134 (N_48134,N_47963,N_47860);
nor U48135 (N_48135,N_47790,N_47773);
and U48136 (N_48136,N_47983,N_47871);
xnor U48137 (N_48137,N_47982,N_47888);
nor U48138 (N_48138,N_47894,N_47753);
or U48139 (N_48139,N_47869,N_47991);
xor U48140 (N_48140,N_47794,N_47773);
or U48141 (N_48141,N_47752,N_47884);
or U48142 (N_48142,N_47920,N_47791);
xor U48143 (N_48143,N_47813,N_47875);
nand U48144 (N_48144,N_47830,N_47871);
or U48145 (N_48145,N_47993,N_47788);
and U48146 (N_48146,N_47939,N_47827);
xor U48147 (N_48147,N_47912,N_47877);
nor U48148 (N_48148,N_47986,N_47990);
or U48149 (N_48149,N_47883,N_47836);
xor U48150 (N_48150,N_47813,N_47995);
nand U48151 (N_48151,N_47997,N_47765);
and U48152 (N_48152,N_47872,N_47824);
nor U48153 (N_48153,N_47848,N_47886);
xor U48154 (N_48154,N_47752,N_47872);
xnor U48155 (N_48155,N_47841,N_47979);
nor U48156 (N_48156,N_47960,N_47918);
or U48157 (N_48157,N_47793,N_47833);
and U48158 (N_48158,N_47920,N_47845);
or U48159 (N_48159,N_47769,N_47811);
nand U48160 (N_48160,N_47835,N_47775);
or U48161 (N_48161,N_47828,N_47960);
nor U48162 (N_48162,N_47834,N_47819);
and U48163 (N_48163,N_47912,N_47887);
xnor U48164 (N_48164,N_47933,N_47773);
or U48165 (N_48165,N_47989,N_47879);
nand U48166 (N_48166,N_47783,N_47942);
nand U48167 (N_48167,N_47788,N_47790);
and U48168 (N_48168,N_47797,N_47778);
xor U48169 (N_48169,N_47801,N_47897);
nand U48170 (N_48170,N_47767,N_47913);
or U48171 (N_48171,N_47793,N_47970);
nand U48172 (N_48172,N_47812,N_47785);
xor U48173 (N_48173,N_47903,N_47801);
and U48174 (N_48174,N_47922,N_47903);
xor U48175 (N_48175,N_47976,N_47841);
or U48176 (N_48176,N_47876,N_47884);
nor U48177 (N_48177,N_47926,N_47835);
or U48178 (N_48178,N_47756,N_47840);
or U48179 (N_48179,N_47810,N_47806);
or U48180 (N_48180,N_47794,N_47768);
or U48181 (N_48181,N_47862,N_47839);
nor U48182 (N_48182,N_47909,N_47938);
xor U48183 (N_48183,N_47782,N_47942);
or U48184 (N_48184,N_47764,N_47887);
xnor U48185 (N_48185,N_47964,N_47942);
nor U48186 (N_48186,N_47869,N_47979);
xor U48187 (N_48187,N_47997,N_47888);
nor U48188 (N_48188,N_47823,N_47980);
and U48189 (N_48189,N_47875,N_47863);
nand U48190 (N_48190,N_47783,N_47773);
nor U48191 (N_48191,N_47849,N_47799);
nor U48192 (N_48192,N_47874,N_47961);
or U48193 (N_48193,N_47807,N_47912);
xor U48194 (N_48194,N_47876,N_47987);
and U48195 (N_48195,N_47788,N_47922);
and U48196 (N_48196,N_47831,N_47890);
or U48197 (N_48197,N_47920,N_47874);
xnor U48198 (N_48198,N_47891,N_47983);
nand U48199 (N_48199,N_47784,N_47764);
nor U48200 (N_48200,N_47911,N_47804);
xnor U48201 (N_48201,N_47935,N_47936);
and U48202 (N_48202,N_47955,N_47980);
or U48203 (N_48203,N_47807,N_47802);
nor U48204 (N_48204,N_47908,N_47787);
xor U48205 (N_48205,N_47767,N_47805);
and U48206 (N_48206,N_47949,N_47839);
nand U48207 (N_48207,N_47957,N_47811);
nand U48208 (N_48208,N_47940,N_47862);
nand U48209 (N_48209,N_47799,N_47833);
nor U48210 (N_48210,N_47936,N_47990);
xor U48211 (N_48211,N_47825,N_47919);
nand U48212 (N_48212,N_47879,N_47919);
or U48213 (N_48213,N_47813,N_47882);
xor U48214 (N_48214,N_47944,N_47977);
nand U48215 (N_48215,N_47910,N_47781);
nand U48216 (N_48216,N_47978,N_47820);
or U48217 (N_48217,N_47787,N_47750);
and U48218 (N_48218,N_47873,N_47996);
nand U48219 (N_48219,N_47799,N_47933);
nand U48220 (N_48220,N_47955,N_47953);
nor U48221 (N_48221,N_47820,N_47852);
nand U48222 (N_48222,N_47807,N_47853);
or U48223 (N_48223,N_47982,N_47933);
nand U48224 (N_48224,N_47852,N_47952);
or U48225 (N_48225,N_47887,N_47991);
and U48226 (N_48226,N_47964,N_47916);
or U48227 (N_48227,N_47884,N_47833);
xnor U48228 (N_48228,N_47943,N_47894);
nor U48229 (N_48229,N_47920,N_47789);
xor U48230 (N_48230,N_47925,N_47909);
xor U48231 (N_48231,N_47863,N_47840);
and U48232 (N_48232,N_47847,N_47781);
nor U48233 (N_48233,N_47788,N_47770);
and U48234 (N_48234,N_47791,N_47865);
nor U48235 (N_48235,N_47985,N_47975);
and U48236 (N_48236,N_47965,N_47978);
or U48237 (N_48237,N_47900,N_47889);
or U48238 (N_48238,N_47806,N_47770);
and U48239 (N_48239,N_47836,N_47774);
nand U48240 (N_48240,N_47878,N_47819);
and U48241 (N_48241,N_47995,N_47915);
nand U48242 (N_48242,N_47969,N_47817);
nand U48243 (N_48243,N_47970,N_47760);
nand U48244 (N_48244,N_47999,N_47916);
xor U48245 (N_48245,N_47860,N_47957);
or U48246 (N_48246,N_47838,N_47778);
or U48247 (N_48247,N_47978,N_47765);
nand U48248 (N_48248,N_47867,N_47959);
nor U48249 (N_48249,N_47981,N_47867);
nor U48250 (N_48250,N_48078,N_48072);
xor U48251 (N_48251,N_48179,N_48089);
and U48252 (N_48252,N_48230,N_48035);
nand U48253 (N_48253,N_48170,N_48200);
nand U48254 (N_48254,N_48055,N_48049);
and U48255 (N_48255,N_48087,N_48084);
or U48256 (N_48256,N_48086,N_48067);
or U48257 (N_48257,N_48209,N_48199);
and U48258 (N_48258,N_48233,N_48020);
or U48259 (N_48259,N_48228,N_48081);
and U48260 (N_48260,N_48217,N_48010);
nor U48261 (N_48261,N_48120,N_48158);
and U48262 (N_48262,N_48042,N_48095);
nand U48263 (N_48263,N_48106,N_48163);
and U48264 (N_48264,N_48050,N_48039);
and U48265 (N_48265,N_48202,N_48156);
nand U48266 (N_48266,N_48136,N_48013);
and U48267 (N_48267,N_48249,N_48130);
or U48268 (N_48268,N_48237,N_48041);
and U48269 (N_48269,N_48167,N_48148);
nor U48270 (N_48270,N_48145,N_48248);
nor U48271 (N_48271,N_48162,N_48022);
and U48272 (N_48272,N_48026,N_48242);
xnor U48273 (N_48273,N_48169,N_48241);
nor U48274 (N_48274,N_48213,N_48168);
nand U48275 (N_48275,N_48238,N_48031);
or U48276 (N_48276,N_48066,N_48061);
and U48277 (N_48277,N_48060,N_48208);
nand U48278 (N_48278,N_48027,N_48194);
nor U48279 (N_48279,N_48048,N_48015);
nor U48280 (N_48280,N_48152,N_48117);
xnor U48281 (N_48281,N_48235,N_48108);
xnor U48282 (N_48282,N_48220,N_48150);
and U48283 (N_48283,N_48166,N_48184);
and U48284 (N_48284,N_48001,N_48044);
nor U48285 (N_48285,N_48180,N_48164);
nor U48286 (N_48286,N_48111,N_48149);
xnor U48287 (N_48287,N_48146,N_48033);
xnor U48288 (N_48288,N_48114,N_48131);
nor U48289 (N_48289,N_48183,N_48077);
nor U48290 (N_48290,N_48219,N_48009);
nor U48291 (N_48291,N_48211,N_48103);
nor U48292 (N_48292,N_48173,N_48215);
and U48293 (N_48293,N_48176,N_48017);
or U48294 (N_48294,N_48032,N_48038);
xnor U48295 (N_48295,N_48126,N_48040);
and U48296 (N_48296,N_48161,N_48094);
nand U48297 (N_48297,N_48037,N_48046);
and U48298 (N_48298,N_48189,N_48098);
nand U48299 (N_48299,N_48064,N_48122);
xnor U48300 (N_48300,N_48076,N_48236);
nand U48301 (N_48301,N_48141,N_48082);
and U48302 (N_48302,N_48139,N_48043);
nand U48303 (N_48303,N_48070,N_48204);
xnor U48304 (N_48304,N_48210,N_48196);
nor U48305 (N_48305,N_48011,N_48193);
or U48306 (N_48306,N_48069,N_48191);
xor U48307 (N_48307,N_48000,N_48028);
and U48308 (N_48308,N_48216,N_48102);
nor U48309 (N_48309,N_48109,N_48240);
xnor U48310 (N_48310,N_48008,N_48014);
xnor U48311 (N_48311,N_48195,N_48071);
or U48312 (N_48312,N_48115,N_48177);
xor U48313 (N_48313,N_48036,N_48100);
or U48314 (N_48314,N_48129,N_48187);
and U48315 (N_48315,N_48075,N_48097);
or U48316 (N_48316,N_48118,N_48052);
xor U48317 (N_48317,N_48218,N_48023);
or U48318 (N_48318,N_48239,N_48025);
and U48319 (N_48319,N_48154,N_48016);
xnor U48320 (N_48320,N_48155,N_48062);
xnor U48321 (N_48321,N_48172,N_48030);
nor U48322 (N_48322,N_48053,N_48201);
nand U48323 (N_48323,N_48143,N_48113);
nand U48324 (N_48324,N_48185,N_48175);
nand U48325 (N_48325,N_48214,N_48063);
and U48326 (N_48326,N_48018,N_48178);
xnor U48327 (N_48327,N_48153,N_48142);
and U48328 (N_48328,N_48006,N_48007);
nor U48329 (N_48329,N_48065,N_48144);
nand U48330 (N_48330,N_48083,N_48207);
xnor U48331 (N_48331,N_48192,N_48088);
xnor U48332 (N_48332,N_48073,N_48024);
or U48333 (N_48333,N_48138,N_48128);
xor U48334 (N_48334,N_48221,N_48079);
nor U48335 (N_48335,N_48080,N_48247);
and U48336 (N_48336,N_48159,N_48134);
and U48337 (N_48337,N_48234,N_48123);
or U48338 (N_48338,N_48151,N_48160);
nor U48339 (N_48339,N_48112,N_48034);
and U48340 (N_48340,N_48212,N_48054);
and U48341 (N_48341,N_48056,N_48232);
nand U48342 (N_48342,N_48188,N_48005);
xnor U48343 (N_48343,N_48205,N_48047);
or U48344 (N_48344,N_48225,N_48093);
nor U48345 (N_48345,N_48068,N_48229);
or U48346 (N_48346,N_48181,N_48002);
nand U48347 (N_48347,N_48245,N_48121);
nand U48348 (N_48348,N_48231,N_48099);
xor U48349 (N_48349,N_48105,N_48085);
and U48350 (N_48350,N_48182,N_48058);
or U48351 (N_48351,N_48174,N_48132);
or U48352 (N_48352,N_48092,N_48059);
or U48353 (N_48353,N_48222,N_48246);
nor U48354 (N_48354,N_48090,N_48012);
nor U48355 (N_48355,N_48110,N_48165);
and U48356 (N_48356,N_48157,N_48127);
or U48357 (N_48357,N_48171,N_48147);
or U48358 (N_48358,N_48116,N_48045);
xor U48359 (N_48359,N_48224,N_48227);
or U48360 (N_48360,N_48074,N_48135);
xnor U48361 (N_48361,N_48133,N_48107);
or U48362 (N_48362,N_48203,N_48124);
xor U48363 (N_48363,N_48119,N_48091);
nor U48364 (N_48364,N_48243,N_48198);
or U48365 (N_48365,N_48125,N_48137);
nand U48366 (N_48366,N_48140,N_48057);
or U48367 (N_48367,N_48051,N_48190);
xor U48368 (N_48368,N_48096,N_48021);
and U48369 (N_48369,N_48019,N_48004);
and U48370 (N_48370,N_48029,N_48226);
and U48371 (N_48371,N_48223,N_48197);
nor U48372 (N_48372,N_48101,N_48244);
nand U48373 (N_48373,N_48003,N_48186);
or U48374 (N_48374,N_48206,N_48104);
nor U48375 (N_48375,N_48011,N_48060);
nand U48376 (N_48376,N_48239,N_48117);
xor U48377 (N_48377,N_48186,N_48167);
nor U48378 (N_48378,N_48121,N_48044);
xor U48379 (N_48379,N_48059,N_48150);
xor U48380 (N_48380,N_48249,N_48216);
or U48381 (N_48381,N_48179,N_48019);
and U48382 (N_48382,N_48102,N_48184);
xor U48383 (N_48383,N_48096,N_48018);
nor U48384 (N_48384,N_48121,N_48013);
xor U48385 (N_48385,N_48060,N_48062);
nor U48386 (N_48386,N_48089,N_48209);
xor U48387 (N_48387,N_48140,N_48205);
nand U48388 (N_48388,N_48201,N_48045);
or U48389 (N_48389,N_48089,N_48103);
nand U48390 (N_48390,N_48174,N_48190);
and U48391 (N_48391,N_48058,N_48018);
nand U48392 (N_48392,N_48083,N_48148);
nand U48393 (N_48393,N_48055,N_48130);
or U48394 (N_48394,N_48221,N_48139);
and U48395 (N_48395,N_48005,N_48090);
xor U48396 (N_48396,N_48192,N_48180);
nor U48397 (N_48397,N_48150,N_48136);
or U48398 (N_48398,N_48211,N_48005);
or U48399 (N_48399,N_48072,N_48090);
nand U48400 (N_48400,N_48067,N_48209);
nor U48401 (N_48401,N_48055,N_48223);
or U48402 (N_48402,N_48017,N_48022);
or U48403 (N_48403,N_48200,N_48066);
nand U48404 (N_48404,N_48090,N_48195);
nand U48405 (N_48405,N_48087,N_48029);
or U48406 (N_48406,N_48182,N_48075);
or U48407 (N_48407,N_48192,N_48225);
or U48408 (N_48408,N_48020,N_48103);
nand U48409 (N_48409,N_48236,N_48104);
and U48410 (N_48410,N_48032,N_48177);
nor U48411 (N_48411,N_48035,N_48102);
nor U48412 (N_48412,N_48085,N_48219);
nand U48413 (N_48413,N_48066,N_48009);
and U48414 (N_48414,N_48083,N_48123);
nand U48415 (N_48415,N_48089,N_48238);
and U48416 (N_48416,N_48028,N_48016);
nor U48417 (N_48417,N_48001,N_48149);
and U48418 (N_48418,N_48056,N_48205);
or U48419 (N_48419,N_48128,N_48162);
nand U48420 (N_48420,N_48177,N_48056);
and U48421 (N_48421,N_48206,N_48130);
and U48422 (N_48422,N_48055,N_48186);
or U48423 (N_48423,N_48063,N_48171);
or U48424 (N_48424,N_48030,N_48020);
nor U48425 (N_48425,N_48225,N_48100);
and U48426 (N_48426,N_48246,N_48184);
and U48427 (N_48427,N_48226,N_48194);
or U48428 (N_48428,N_48116,N_48220);
and U48429 (N_48429,N_48099,N_48211);
nor U48430 (N_48430,N_48088,N_48037);
nand U48431 (N_48431,N_48063,N_48156);
nand U48432 (N_48432,N_48206,N_48173);
nand U48433 (N_48433,N_48151,N_48117);
nor U48434 (N_48434,N_48001,N_48198);
and U48435 (N_48435,N_48055,N_48085);
nand U48436 (N_48436,N_48184,N_48061);
nor U48437 (N_48437,N_48154,N_48168);
nor U48438 (N_48438,N_48249,N_48174);
nor U48439 (N_48439,N_48173,N_48058);
nor U48440 (N_48440,N_48136,N_48021);
nor U48441 (N_48441,N_48206,N_48124);
nor U48442 (N_48442,N_48098,N_48024);
nor U48443 (N_48443,N_48180,N_48042);
xnor U48444 (N_48444,N_48008,N_48111);
nand U48445 (N_48445,N_48126,N_48245);
and U48446 (N_48446,N_48012,N_48209);
nand U48447 (N_48447,N_48234,N_48047);
nand U48448 (N_48448,N_48164,N_48228);
xor U48449 (N_48449,N_48153,N_48005);
xor U48450 (N_48450,N_48138,N_48189);
or U48451 (N_48451,N_48227,N_48068);
nand U48452 (N_48452,N_48204,N_48202);
and U48453 (N_48453,N_48058,N_48046);
xor U48454 (N_48454,N_48207,N_48074);
nor U48455 (N_48455,N_48011,N_48002);
or U48456 (N_48456,N_48168,N_48192);
and U48457 (N_48457,N_48172,N_48173);
and U48458 (N_48458,N_48085,N_48024);
nand U48459 (N_48459,N_48018,N_48211);
and U48460 (N_48460,N_48004,N_48047);
xor U48461 (N_48461,N_48129,N_48054);
or U48462 (N_48462,N_48025,N_48189);
nand U48463 (N_48463,N_48002,N_48100);
or U48464 (N_48464,N_48191,N_48086);
or U48465 (N_48465,N_48211,N_48127);
nor U48466 (N_48466,N_48132,N_48000);
or U48467 (N_48467,N_48152,N_48011);
nor U48468 (N_48468,N_48226,N_48025);
and U48469 (N_48469,N_48127,N_48247);
nor U48470 (N_48470,N_48036,N_48238);
xnor U48471 (N_48471,N_48203,N_48181);
nand U48472 (N_48472,N_48202,N_48209);
xnor U48473 (N_48473,N_48100,N_48167);
nand U48474 (N_48474,N_48158,N_48188);
nor U48475 (N_48475,N_48180,N_48215);
and U48476 (N_48476,N_48106,N_48116);
nor U48477 (N_48477,N_48060,N_48136);
and U48478 (N_48478,N_48206,N_48099);
nand U48479 (N_48479,N_48050,N_48053);
nor U48480 (N_48480,N_48140,N_48011);
nor U48481 (N_48481,N_48018,N_48195);
nand U48482 (N_48482,N_48170,N_48039);
and U48483 (N_48483,N_48179,N_48205);
or U48484 (N_48484,N_48197,N_48056);
nor U48485 (N_48485,N_48122,N_48248);
nor U48486 (N_48486,N_48011,N_48197);
nand U48487 (N_48487,N_48160,N_48020);
xnor U48488 (N_48488,N_48141,N_48027);
and U48489 (N_48489,N_48235,N_48152);
and U48490 (N_48490,N_48236,N_48043);
nor U48491 (N_48491,N_48248,N_48157);
and U48492 (N_48492,N_48157,N_48106);
or U48493 (N_48493,N_48208,N_48220);
nor U48494 (N_48494,N_48206,N_48112);
nand U48495 (N_48495,N_48088,N_48039);
nor U48496 (N_48496,N_48066,N_48241);
and U48497 (N_48497,N_48173,N_48040);
or U48498 (N_48498,N_48107,N_48024);
nand U48499 (N_48499,N_48218,N_48108);
and U48500 (N_48500,N_48340,N_48422);
nand U48501 (N_48501,N_48485,N_48286);
nand U48502 (N_48502,N_48489,N_48398);
and U48503 (N_48503,N_48289,N_48278);
nand U48504 (N_48504,N_48363,N_48268);
nor U48505 (N_48505,N_48439,N_48322);
or U48506 (N_48506,N_48317,N_48281);
or U48507 (N_48507,N_48313,N_48396);
nor U48508 (N_48508,N_48464,N_48385);
nor U48509 (N_48509,N_48453,N_48465);
xor U48510 (N_48510,N_48351,N_48434);
nand U48511 (N_48511,N_48495,N_48306);
and U48512 (N_48512,N_48339,N_48491);
nand U48513 (N_48513,N_48372,N_48460);
nor U48514 (N_48514,N_48357,N_48315);
nand U48515 (N_48515,N_48471,N_48272);
nand U48516 (N_48516,N_48253,N_48438);
xor U48517 (N_48517,N_48492,N_48259);
nor U48518 (N_48518,N_48264,N_48271);
or U48519 (N_48519,N_48314,N_48276);
and U48520 (N_48520,N_48343,N_48328);
nand U48521 (N_48521,N_48404,N_48327);
nor U48522 (N_48522,N_48473,N_48494);
nand U48523 (N_48523,N_48361,N_48486);
xor U48524 (N_48524,N_48330,N_48291);
nor U48525 (N_48525,N_48305,N_48430);
nor U48526 (N_48526,N_48300,N_48381);
nor U48527 (N_48527,N_48456,N_48435);
nor U48528 (N_48528,N_48400,N_48394);
and U48529 (N_48529,N_48299,N_48304);
and U48530 (N_48530,N_48288,N_48302);
or U48531 (N_48531,N_48475,N_48362);
and U48532 (N_48532,N_48303,N_48251);
xnor U48533 (N_48533,N_48265,N_48364);
or U48534 (N_48534,N_48488,N_48321);
xor U48535 (N_48535,N_48297,N_48437);
nand U48536 (N_48536,N_48285,N_48451);
xnor U48537 (N_48537,N_48334,N_48454);
xnor U48538 (N_48538,N_48498,N_48267);
xor U48539 (N_48539,N_48405,N_48371);
or U48540 (N_48540,N_48425,N_48294);
nor U48541 (N_48541,N_48252,N_48255);
xnor U48542 (N_48542,N_48307,N_48256);
and U48543 (N_48543,N_48375,N_48496);
xnor U48544 (N_48544,N_48277,N_48308);
and U48545 (N_48545,N_48316,N_48369);
or U48546 (N_48546,N_48287,N_48312);
and U48547 (N_48547,N_48382,N_48335);
nor U48548 (N_48548,N_48254,N_48478);
and U48549 (N_48549,N_48349,N_48436);
nand U48550 (N_48550,N_48386,N_48426);
and U48551 (N_48551,N_48416,N_48499);
and U48552 (N_48552,N_48350,N_48470);
xor U48553 (N_48553,N_48411,N_48283);
nor U48554 (N_48554,N_48459,N_48332);
nand U48555 (N_48555,N_48387,N_48466);
or U48556 (N_48556,N_48427,N_48290);
xor U48557 (N_48557,N_48341,N_48417);
nand U48558 (N_48558,N_48452,N_48463);
or U48559 (N_48559,N_48458,N_48358);
xnor U48560 (N_48560,N_48389,N_48424);
and U48561 (N_48561,N_48445,N_48431);
xor U48562 (N_48562,N_48354,N_48298);
and U48563 (N_48563,N_48409,N_48432);
nand U48564 (N_48564,N_48338,N_48482);
nand U48565 (N_48565,N_48379,N_48457);
or U48566 (N_48566,N_48367,N_48266);
and U48567 (N_48567,N_48423,N_48447);
or U48568 (N_48568,N_48415,N_48376);
and U48569 (N_48569,N_48476,N_48433);
nand U48570 (N_48570,N_48260,N_48352);
or U48571 (N_48571,N_48270,N_48301);
and U48572 (N_48572,N_48257,N_48356);
or U48573 (N_48573,N_48323,N_48262);
xnor U48574 (N_48574,N_48269,N_48368);
nor U48575 (N_48575,N_48261,N_48383);
nand U48576 (N_48576,N_48370,N_48449);
xnor U48577 (N_48577,N_48331,N_48468);
or U48578 (N_48578,N_48472,N_48326);
and U48579 (N_48579,N_48414,N_48483);
or U48580 (N_48580,N_48420,N_48462);
or U48581 (N_48581,N_48295,N_48388);
xnor U48582 (N_48582,N_48380,N_48273);
nor U48583 (N_48583,N_48467,N_48408);
and U48584 (N_48584,N_48345,N_48441);
nor U48585 (N_48585,N_48481,N_48342);
nand U48586 (N_48586,N_48395,N_48347);
nand U48587 (N_48587,N_48353,N_48263);
nor U48588 (N_48588,N_48402,N_48250);
or U48589 (N_48589,N_48324,N_48365);
or U48590 (N_48590,N_48310,N_48325);
nor U48591 (N_48591,N_48329,N_48280);
xnor U48592 (N_48592,N_48344,N_48355);
nand U48593 (N_48593,N_48275,N_48455);
xnor U48594 (N_48594,N_48446,N_48418);
and U48595 (N_48595,N_48378,N_48443);
nand U48596 (N_48596,N_48480,N_48474);
or U48597 (N_48597,N_48279,N_48318);
and U48598 (N_48598,N_48390,N_48292);
and U48599 (N_48599,N_48377,N_48333);
or U48600 (N_48600,N_48442,N_48274);
and U48601 (N_48601,N_48497,N_48469);
xor U48602 (N_48602,N_48360,N_48319);
nand U48603 (N_48603,N_48419,N_48309);
and U48604 (N_48604,N_48413,N_48407);
and U48605 (N_48605,N_48258,N_48428);
nand U48606 (N_48606,N_48401,N_48448);
xnor U48607 (N_48607,N_48373,N_48348);
nor U48608 (N_48608,N_48337,N_48391);
or U48609 (N_48609,N_48421,N_48336);
or U48610 (N_48610,N_48403,N_48429);
and U48611 (N_48611,N_48282,N_48384);
or U48612 (N_48612,N_48487,N_48284);
and U48613 (N_48613,N_48374,N_48320);
nand U48614 (N_48614,N_48366,N_48444);
or U48615 (N_48615,N_48412,N_48490);
or U48616 (N_48616,N_48410,N_48296);
or U48617 (N_48617,N_48484,N_48311);
nand U48618 (N_48618,N_48293,N_48399);
or U48619 (N_48619,N_48479,N_48440);
nand U48620 (N_48620,N_48393,N_48359);
nor U48621 (N_48621,N_48346,N_48477);
and U48622 (N_48622,N_48450,N_48406);
or U48623 (N_48623,N_48461,N_48493);
xor U48624 (N_48624,N_48397,N_48392);
and U48625 (N_48625,N_48463,N_48259);
nor U48626 (N_48626,N_48470,N_48487);
or U48627 (N_48627,N_48386,N_48367);
nor U48628 (N_48628,N_48315,N_48490);
nand U48629 (N_48629,N_48463,N_48475);
nor U48630 (N_48630,N_48251,N_48283);
nor U48631 (N_48631,N_48356,N_48279);
or U48632 (N_48632,N_48418,N_48324);
nand U48633 (N_48633,N_48426,N_48267);
or U48634 (N_48634,N_48339,N_48458);
or U48635 (N_48635,N_48367,N_48376);
and U48636 (N_48636,N_48346,N_48378);
nand U48637 (N_48637,N_48487,N_48427);
nor U48638 (N_48638,N_48403,N_48325);
nor U48639 (N_48639,N_48332,N_48344);
nand U48640 (N_48640,N_48285,N_48286);
or U48641 (N_48641,N_48365,N_48404);
xor U48642 (N_48642,N_48282,N_48414);
xnor U48643 (N_48643,N_48256,N_48285);
nor U48644 (N_48644,N_48309,N_48487);
nor U48645 (N_48645,N_48421,N_48378);
xnor U48646 (N_48646,N_48385,N_48288);
xnor U48647 (N_48647,N_48420,N_48267);
nor U48648 (N_48648,N_48378,N_48286);
and U48649 (N_48649,N_48354,N_48456);
nor U48650 (N_48650,N_48404,N_48408);
or U48651 (N_48651,N_48313,N_48460);
or U48652 (N_48652,N_48368,N_48361);
xor U48653 (N_48653,N_48317,N_48448);
nor U48654 (N_48654,N_48417,N_48425);
nor U48655 (N_48655,N_48342,N_48359);
nor U48656 (N_48656,N_48285,N_48393);
or U48657 (N_48657,N_48390,N_48442);
nor U48658 (N_48658,N_48355,N_48321);
and U48659 (N_48659,N_48316,N_48324);
and U48660 (N_48660,N_48330,N_48445);
and U48661 (N_48661,N_48436,N_48261);
nor U48662 (N_48662,N_48291,N_48332);
and U48663 (N_48663,N_48421,N_48454);
xor U48664 (N_48664,N_48499,N_48320);
nor U48665 (N_48665,N_48360,N_48484);
and U48666 (N_48666,N_48385,N_48342);
and U48667 (N_48667,N_48306,N_48289);
nand U48668 (N_48668,N_48471,N_48485);
or U48669 (N_48669,N_48326,N_48323);
and U48670 (N_48670,N_48317,N_48461);
nor U48671 (N_48671,N_48445,N_48392);
xnor U48672 (N_48672,N_48444,N_48460);
nand U48673 (N_48673,N_48292,N_48251);
nand U48674 (N_48674,N_48472,N_48296);
nand U48675 (N_48675,N_48465,N_48377);
nand U48676 (N_48676,N_48267,N_48338);
or U48677 (N_48677,N_48297,N_48389);
nand U48678 (N_48678,N_48428,N_48322);
xnor U48679 (N_48679,N_48383,N_48411);
and U48680 (N_48680,N_48412,N_48345);
or U48681 (N_48681,N_48475,N_48361);
nor U48682 (N_48682,N_48257,N_48461);
and U48683 (N_48683,N_48356,N_48473);
xor U48684 (N_48684,N_48401,N_48409);
xnor U48685 (N_48685,N_48451,N_48379);
and U48686 (N_48686,N_48385,N_48302);
nor U48687 (N_48687,N_48285,N_48370);
xor U48688 (N_48688,N_48423,N_48437);
and U48689 (N_48689,N_48496,N_48454);
nor U48690 (N_48690,N_48275,N_48352);
xor U48691 (N_48691,N_48414,N_48435);
or U48692 (N_48692,N_48258,N_48313);
nor U48693 (N_48693,N_48405,N_48341);
nand U48694 (N_48694,N_48400,N_48302);
xor U48695 (N_48695,N_48383,N_48256);
and U48696 (N_48696,N_48268,N_48460);
and U48697 (N_48697,N_48283,N_48449);
nand U48698 (N_48698,N_48346,N_48299);
nor U48699 (N_48699,N_48488,N_48313);
or U48700 (N_48700,N_48468,N_48356);
or U48701 (N_48701,N_48320,N_48443);
and U48702 (N_48702,N_48406,N_48464);
or U48703 (N_48703,N_48282,N_48385);
and U48704 (N_48704,N_48279,N_48381);
nor U48705 (N_48705,N_48438,N_48313);
xnor U48706 (N_48706,N_48263,N_48483);
xor U48707 (N_48707,N_48388,N_48296);
nor U48708 (N_48708,N_48406,N_48295);
or U48709 (N_48709,N_48440,N_48263);
nor U48710 (N_48710,N_48307,N_48342);
nand U48711 (N_48711,N_48378,N_48403);
or U48712 (N_48712,N_48384,N_48492);
xnor U48713 (N_48713,N_48462,N_48449);
nand U48714 (N_48714,N_48494,N_48404);
or U48715 (N_48715,N_48337,N_48439);
nand U48716 (N_48716,N_48406,N_48498);
nor U48717 (N_48717,N_48358,N_48282);
xor U48718 (N_48718,N_48290,N_48422);
or U48719 (N_48719,N_48347,N_48287);
nor U48720 (N_48720,N_48396,N_48432);
nor U48721 (N_48721,N_48468,N_48426);
xnor U48722 (N_48722,N_48417,N_48283);
nor U48723 (N_48723,N_48264,N_48435);
and U48724 (N_48724,N_48279,N_48470);
nand U48725 (N_48725,N_48463,N_48466);
nor U48726 (N_48726,N_48472,N_48390);
nor U48727 (N_48727,N_48338,N_48284);
xnor U48728 (N_48728,N_48433,N_48361);
or U48729 (N_48729,N_48328,N_48449);
or U48730 (N_48730,N_48402,N_48456);
and U48731 (N_48731,N_48463,N_48444);
nor U48732 (N_48732,N_48270,N_48393);
and U48733 (N_48733,N_48325,N_48339);
xor U48734 (N_48734,N_48326,N_48385);
and U48735 (N_48735,N_48279,N_48348);
and U48736 (N_48736,N_48302,N_48348);
xnor U48737 (N_48737,N_48265,N_48430);
or U48738 (N_48738,N_48265,N_48369);
xor U48739 (N_48739,N_48454,N_48278);
or U48740 (N_48740,N_48335,N_48434);
xnor U48741 (N_48741,N_48321,N_48269);
nor U48742 (N_48742,N_48314,N_48476);
nand U48743 (N_48743,N_48346,N_48491);
nor U48744 (N_48744,N_48323,N_48437);
and U48745 (N_48745,N_48257,N_48494);
or U48746 (N_48746,N_48422,N_48394);
or U48747 (N_48747,N_48383,N_48287);
and U48748 (N_48748,N_48342,N_48444);
or U48749 (N_48749,N_48342,N_48303);
nand U48750 (N_48750,N_48738,N_48737);
and U48751 (N_48751,N_48660,N_48650);
or U48752 (N_48752,N_48619,N_48569);
nand U48753 (N_48753,N_48731,N_48587);
nand U48754 (N_48754,N_48654,N_48739);
or U48755 (N_48755,N_48642,N_48597);
nand U48756 (N_48756,N_48567,N_48518);
xor U48757 (N_48757,N_48524,N_48720);
xor U48758 (N_48758,N_48555,N_48529);
or U48759 (N_48759,N_48576,N_48583);
xnor U48760 (N_48760,N_48709,N_48584);
xor U48761 (N_48761,N_48546,N_48512);
nand U48762 (N_48762,N_48504,N_48548);
xnor U48763 (N_48763,N_48649,N_48532);
xor U48764 (N_48764,N_48594,N_48668);
and U48765 (N_48765,N_48600,N_48615);
or U48766 (N_48766,N_48684,N_48707);
xor U48767 (N_48767,N_48581,N_48562);
or U48768 (N_48768,N_48664,N_48685);
or U48769 (N_48769,N_48675,N_48509);
and U48770 (N_48770,N_48609,N_48634);
xnor U48771 (N_48771,N_48582,N_48696);
nand U48772 (N_48772,N_48551,N_48645);
or U48773 (N_48773,N_48710,N_48703);
or U48774 (N_48774,N_48687,N_48617);
xnor U48775 (N_48775,N_48718,N_48655);
and U48776 (N_48776,N_48560,N_48699);
or U48777 (N_48777,N_48653,N_48639);
nand U48778 (N_48778,N_48697,N_48537);
xor U48779 (N_48779,N_48622,N_48591);
and U48780 (N_48780,N_48605,N_48701);
and U48781 (N_48781,N_48662,N_48745);
nor U48782 (N_48782,N_48531,N_48572);
nand U48783 (N_48783,N_48514,N_48728);
nor U48784 (N_48784,N_48734,N_48667);
and U48785 (N_48785,N_48610,N_48693);
and U48786 (N_48786,N_48553,N_48636);
nor U48787 (N_48787,N_48680,N_48694);
nor U48788 (N_48788,N_48590,N_48652);
or U48789 (N_48789,N_48657,N_48723);
nand U48790 (N_48790,N_48640,N_48677);
nand U48791 (N_48791,N_48500,N_48742);
xnor U48792 (N_48792,N_48603,N_48700);
or U48793 (N_48793,N_48540,N_48674);
nand U48794 (N_48794,N_48580,N_48545);
xor U48795 (N_48795,N_48564,N_48632);
nor U48796 (N_48796,N_48690,N_48679);
or U48797 (N_48797,N_48596,N_48656);
or U48798 (N_48798,N_48698,N_48706);
and U48799 (N_48799,N_48541,N_48724);
nand U48800 (N_48800,N_48643,N_48683);
xnor U48801 (N_48801,N_48507,N_48542);
or U48802 (N_48802,N_48614,N_48549);
and U48803 (N_48803,N_48611,N_48501);
nor U48804 (N_48804,N_48601,N_48519);
nand U48805 (N_48805,N_48563,N_48565);
xnor U48806 (N_48806,N_48666,N_48641);
nand U48807 (N_48807,N_48744,N_48574);
and U48808 (N_48808,N_48613,N_48722);
and U48809 (N_48809,N_48628,N_48708);
xor U48810 (N_48810,N_48711,N_48535);
and U48811 (N_48811,N_48525,N_48612);
nor U48812 (N_48812,N_48559,N_48659);
nor U48813 (N_48813,N_48646,N_48616);
xnor U48814 (N_48814,N_48705,N_48658);
nand U48815 (N_48815,N_48624,N_48593);
nor U48816 (N_48816,N_48558,N_48681);
and U48817 (N_48817,N_48638,N_48536);
and U48818 (N_48818,N_48626,N_48644);
and U48819 (N_48819,N_48573,N_48550);
and U48820 (N_48820,N_48589,N_48586);
nand U48821 (N_48821,N_48665,N_48689);
or U48822 (N_48822,N_48741,N_48727);
and U48823 (N_48823,N_48682,N_48527);
xor U48824 (N_48824,N_48726,N_48577);
xnor U48825 (N_48825,N_48678,N_48733);
and U48826 (N_48826,N_48543,N_48714);
and U48827 (N_48827,N_48676,N_48716);
xnor U48828 (N_48828,N_48721,N_48595);
xnor U48829 (N_48829,N_48521,N_48719);
nand U48830 (N_48830,N_48604,N_48740);
nand U48831 (N_48831,N_48575,N_48561);
and U48832 (N_48832,N_48534,N_48633);
or U48833 (N_48833,N_48625,N_48637);
and U48834 (N_48834,N_48522,N_48673);
xor U48835 (N_48835,N_48506,N_48533);
and U48836 (N_48836,N_48648,N_48651);
and U48837 (N_48837,N_48544,N_48602);
or U48838 (N_48838,N_48528,N_48688);
nand U48839 (N_48839,N_48513,N_48630);
and U48840 (N_48840,N_48510,N_48515);
nand U48841 (N_48841,N_48557,N_48552);
and U48842 (N_48842,N_48671,N_48547);
xor U48843 (N_48843,N_48566,N_48505);
or U48844 (N_48844,N_48704,N_48517);
xnor U48845 (N_48845,N_48554,N_48618);
xor U48846 (N_48846,N_48599,N_48712);
nor U48847 (N_48847,N_48672,N_48730);
nand U48848 (N_48848,N_48691,N_48661);
or U48849 (N_48849,N_48556,N_48508);
nor U48850 (N_48850,N_48607,N_48732);
nand U48851 (N_48851,N_48623,N_48725);
xnor U48852 (N_48852,N_48627,N_48606);
nand U48853 (N_48853,N_48692,N_48598);
xor U48854 (N_48854,N_48539,N_48746);
or U48855 (N_48855,N_48511,N_48735);
or U48856 (N_48856,N_48747,N_48520);
xnor U48857 (N_48857,N_48663,N_48503);
nor U48858 (N_48858,N_48686,N_48749);
and U48859 (N_48859,N_48621,N_48713);
nand U48860 (N_48860,N_48635,N_48570);
nor U48861 (N_48861,N_48729,N_48629);
or U48862 (N_48862,N_48736,N_48578);
and U48863 (N_48863,N_48585,N_48670);
nor U48864 (N_48864,N_48717,N_48715);
and U48865 (N_48865,N_48695,N_48538);
or U48866 (N_48866,N_48502,N_48743);
xnor U48867 (N_48867,N_48608,N_48702);
nor U48868 (N_48868,N_48571,N_48620);
xnor U48869 (N_48869,N_48631,N_48748);
nand U48870 (N_48870,N_48579,N_48516);
nand U48871 (N_48871,N_48568,N_48530);
or U48872 (N_48872,N_48523,N_48526);
nor U48873 (N_48873,N_48588,N_48592);
and U48874 (N_48874,N_48669,N_48647);
and U48875 (N_48875,N_48560,N_48545);
nand U48876 (N_48876,N_48609,N_48511);
and U48877 (N_48877,N_48568,N_48676);
nor U48878 (N_48878,N_48563,N_48503);
nand U48879 (N_48879,N_48575,N_48710);
nor U48880 (N_48880,N_48739,N_48674);
or U48881 (N_48881,N_48511,N_48605);
and U48882 (N_48882,N_48522,N_48590);
nand U48883 (N_48883,N_48690,N_48611);
or U48884 (N_48884,N_48564,N_48689);
and U48885 (N_48885,N_48741,N_48515);
xor U48886 (N_48886,N_48637,N_48603);
nor U48887 (N_48887,N_48711,N_48665);
or U48888 (N_48888,N_48513,N_48606);
and U48889 (N_48889,N_48662,N_48664);
or U48890 (N_48890,N_48729,N_48728);
nor U48891 (N_48891,N_48582,N_48697);
or U48892 (N_48892,N_48703,N_48573);
xor U48893 (N_48893,N_48633,N_48619);
and U48894 (N_48894,N_48684,N_48734);
xnor U48895 (N_48895,N_48621,N_48647);
or U48896 (N_48896,N_48611,N_48596);
nand U48897 (N_48897,N_48590,N_48547);
and U48898 (N_48898,N_48682,N_48548);
nand U48899 (N_48899,N_48593,N_48570);
nor U48900 (N_48900,N_48681,N_48673);
nor U48901 (N_48901,N_48667,N_48558);
nand U48902 (N_48902,N_48548,N_48661);
nand U48903 (N_48903,N_48658,N_48569);
and U48904 (N_48904,N_48688,N_48566);
nor U48905 (N_48905,N_48546,N_48644);
and U48906 (N_48906,N_48590,N_48613);
nand U48907 (N_48907,N_48544,N_48626);
or U48908 (N_48908,N_48697,N_48514);
nor U48909 (N_48909,N_48565,N_48531);
nor U48910 (N_48910,N_48569,N_48629);
or U48911 (N_48911,N_48716,N_48516);
and U48912 (N_48912,N_48552,N_48735);
nand U48913 (N_48913,N_48698,N_48537);
xor U48914 (N_48914,N_48661,N_48743);
and U48915 (N_48915,N_48523,N_48721);
or U48916 (N_48916,N_48532,N_48604);
and U48917 (N_48917,N_48669,N_48562);
nand U48918 (N_48918,N_48600,N_48552);
and U48919 (N_48919,N_48635,N_48667);
nand U48920 (N_48920,N_48746,N_48663);
nor U48921 (N_48921,N_48570,N_48522);
nand U48922 (N_48922,N_48554,N_48551);
nand U48923 (N_48923,N_48692,N_48605);
xor U48924 (N_48924,N_48516,N_48683);
xnor U48925 (N_48925,N_48670,N_48573);
and U48926 (N_48926,N_48561,N_48533);
and U48927 (N_48927,N_48744,N_48709);
xor U48928 (N_48928,N_48599,N_48604);
or U48929 (N_48929,N_48746,N_48703);
nand U48930 (N_48930,N_48712,N_48622);
nor U48931 (N_48931,N_48715,N_48663);
nand U48932 (N_48932,N_48517,N_48547);
nand U48933 (N_48933,N_48688,N_48705);
or U48934 (N_48934,N_48535,N_48723);
xnor U48935 (N_48935,N_48506,N_48588);
or U48936 (N_48936,N_48503,N_48685);
nand U48937 (N_48937,N_48727,N_48564);
and U48938 (N_48938,N_48558,N_48592);
and U48939 (N_48939,N_48652,N_48684);
and U48940 (N_48940,N_48610,N_48511);
nor U48941 (N_48941,N_48717,N_48566);
or U48942 (N_48942,N_48624,N_48724);
nor U48943 (N_48943,N_48568,N_48644);
nor U48944 (N_48944,N_48576,N_48517);
or U48945 (N_48945,N_48586,N_48715);
xor U48946 (N_48946,N_48700,N_48505);
and U48947 (N_48947,N_48611,N_48732);
and U48948 (N_48948,N_48557,N_48509);
or U48949 (N_48949,N_48679,N_48677);
nand U48950 (N_48950,N_48700,N_48745);
xnor U48951 (N_48951,N_48507,N_48653);
nand U48952 (N_48952,N_48712,N_48570);
nand U48953 (N_48953,N_48587,N_48527);
or U48954 (N_48954,N_48504,N_48628);
or U48955 (N_48955,N_48516,N_48522);
xnor U48956 (N_48956,N_48731,N_48536);
and U48957 (N_48957,N_48596,N_48645);
or U48958 (N_48958,N_48557,N_48514);
and U48959 (N_48959,N_48694,N_48591);
and U48960 (N_48960,N_48605,N_48539);
nand U48961 (N_48961,N_48556,N_48538);
and U48962 (N_48962,N_48511,N_48528);
nor U48963 (N_48963,N_48728,N_48655);
and U48964 (N_48964,N_48664,N_48734);
nor U48965 (N_48965,N_48613,N_48662);
nand U48966 (N_48966,N_48559,N_48618);
or U48967 (N_48967,N_48689,N_48730);
nand U48968 (N_48968,N_48516,N_48611);
or U48969 (N_48969,N_48635,N_48579);
nor U48970 (N_48970,N_48664,N_48549);
or U48971 (N_48971,N_48551,N_48662);
and U48972 (N_48972,N_48662,N_48723);
nand U48973 (N_48973,N_48730,N_48581);
or U48974 (N_48974,N_48540,N_48574);
nor U48975 (N_48975,N_48622,N_48715);
and U48976 (N_48976,N_48666,N_48639);
nand U48977 (N_48977,N_48611,N_48503);
xnor U48978 (N_48978,N_48500,N_48549);
xor U48979 (N_48979,N_48508,N_48674);
or U48980 (N_48980,N_48505,N_48529);
nor U48981 (N_48981,N_48558,N_48695);
or U48982 (N_48982,N_48596,N_48599);
or U48983 (N_48983,N_48557,N_48695);
or U48984 (N_48984,N_48557,N_48601);
xnor U48985 (N_48985,N_48680,N_48596);
or U48986 (N_48986,N_48702,N_48538);
and U48987 (N_48987,N_48735,N_48585);
xor U48988 (N_48988,N_48684,N_48574);
nand U48989 (N_48989,N_48656,N_48741);
and U48990 (N_48990,N_48706,N_48687);
or U48991 (N_48991,N_48556,N_48544);
nor U48992 (N_48992,N_48571,N_48736);
and U48993 (N_48993,N_48719,N_48683);
or U48994 (N_48994,N_48726,N_48734);
and U48995 (N_48995,N_48660,N_48694);
or U48996 (N_48996,N_48630,N_48601);
xor U48997 (N_48997,N_48738,N_48696);
xor U48998 (N_48998,N_48529,N_48675);
nor U48999 (N_48999,N_48658,N_48575);
nor U49000 (N_49000,N_48959,N_48753);
xnor U49001 (N_49001,N_48992,N_48991);
nor U49002 (N_49002,N_48907,N_48935);
and U49003 (N_49003,N_48882,N_48864);
nor U49004 (N_49004,N_48853,N_48788);
nor U49005 (N_49005,N_48970,N_48912);
nand U49006 (N_49006,N_48986,N_48793);
or U49007 (N_49007,N_48758,N_48792);
nor U49008 (N_49008,N_48893,N_48760);
and U49009 (N_49009,N_48955,N_48862);
nor U49010 (N_49010,N_48763,N_48876);
nand U49011 (N_49011,N_48939,N_48757);
xor U49012 (N_49012,N_48999,N_48827);
nor U49013 (N_49013,N_48817,N_48985);
or U49014 (N_49014,N_48924,N_48868);
nand U49015 (N_49015,N_48797,N_48831);
nor U49016 (N_49016,N_48799,N_48766);
nor U49017 (N_49017,N_48805,N_48949);
and U49018 (N_49018,N_48937,N_48789);
nand U49019 (N_49019,N_48978,N_48928);
xor U49020 (N_49020,N_48989,N_48946);
nand U49021 (N_49021,N_48869,N_48752);
and U49022 (N_49022,N_48948,N_48809);
xor U49023 (N_49023,N_48993,N_48828);
xnor U49024 (N_49024,N_48759,N_48934);
nand U49025 (N_49025,N_48814,N_48865);
xnor U49026 (N_49026,N_48834,N_48932);
and U49027 (N_49027,N_48866,N_48765);
or U49028 (N_49028,N_48919,N_48899);
and U49029 (N_49029,N_48849,N_48963);
xor U49030 (N_49030,N_48777,N_48863);
nor U49031 (N_49031,N_48841,N_48943);
or U49032 (N_49032,N_48988,N_48861);
xor U49033 (N_49033,N_48826,N_48904);
nor U49034 (N_49034,N_48927,N_48780);
and U49035 (N_49035,N_48870,N_48901);
nor U49036 (N_49036,N_48878,N_48824);
xor U49037 (N_49037,N_48857,N_48855);
xnor U49038 (N_49038,N_48945,N_48917);
nor U49039 (N_49039,N_48965,N_48957);
and U49040 (N_49040,N_48930,N_48845);
and U49041 (N_49041,N_48852,N_48925);
or U49042 (N_49042,N_48967,N_48846);
nand U49043 (N_49043,N_48835,N_48860);
nor U49044 (N_49044,N_48848,N_48975);
and U49045 (N_49045,N_48931,N_48896);
and U49046 (N_49046,N_48764,N_48881);
nand U49047 (N_49047,N_48856,N_48898);
or U49048 (N_49048,N_48808,N_48905);
nor U49049 (N_49049,N_48964,N_48954);
nor U49050 (N_49050,N_48920,N_48794);
or U49051 (N_49051,N_48938,N_48921);
xnor U49052 (N_49052,N_48790,N_48810);
or U49053 (N_49053,N_48804,N_48781);
nor U49054 (N_49054,N_48908,N_48821);
or U49055 (N_49055,N_48941,N_48916);
or U49056 (N_49056,N_48983,N_48906);
or U49057 (N_49057,N_48889,N_48982);
or U49058 (N_49058,N_48940,N_48770);
nand U49059 (N_49059,N_48891,N_48858);
xor U49060 (N_49060,N_48971,N_48913);
or U49061 (N_49061,N_48922,N_48902);
nor U49062 (N_49062,N_48769,N_48969);
nor U49063 (N_49063,N_48953,N_48818);
nor U49064 (N_49064,N_48762,N_48888);
and U49065 (N_49065,N_48775,N_48806);
or U49066 (N_49066,N_48754,N_48859);
nand U49067 (N_49067,N_48977,N_48877);
xnor U49068 (N_49068,N_48773,N_48926);
nand U49069 (N_49069,N_48851,N_48874);
and U49070 (N_49070,N_48990,N_48783);
or U49071 (N_49071,N_48767,N_48812);
or U49072 (N_49072,N_48998,N_48784);
nor U49073 (N_49073,N_48825,N_48750);
nor U49074 (N_49074,N_48795,N_48802);
xor U49075 (N_49075,N_48847,N_48819);
nand U49076 (N_49076,N_48816,N_48867);
nand U49077 (N_49077,N_48997,N_48914);
or U49078 (N_49078,N_48800,N_48933);
and U49079 (N_49079,N_48952,N_48897);
or U49080 (N_49080,N_48838,N_48796);
nand U49081 (N_49081,N_48798,N_48961);
and U49082 (N_49082,N_48813,N_48942);
nor U49083 (N_49083,N_48911,N_48918);
nor U49084 (N_49084,N_48958,N_48972);
nor U49085 (N_49085,N_48785,N_48909);
xor U49086 (N_49086,N_48973,N_48976);
and U49087 (N_49087,N_48979,N_48923);
and U49088 (N_49088,N_48815,N_48832);
xnor U49089 (N_49089,N_48885,N_48968);
and U49090 (N_49090,N_48887,N_48974);
or U49091 (N_49091,N_48822,N_48837);
nor U49092 (N_49092,N_48761,N_48915);
nand U49093 (N_49093,N_48774,N_48883);
and U49094 (N_49094,N_48807,N_48950);
nor U49095 (N_49095,N_48879,N_48929);
xnor U49096 (N_49096,N_48768,N_48872);
nor U49097 (N_49097,N_48778,N_48829);
nor U49098 (N_49098,N_48786,N_48854);
xor U49099 (N_49099,N_48951,N_48886);
or U49100 (N_49100,N_48944,N_48894);
nand U49101 (N_49101,N_48987,N_48980);
xnor U49102 (N_49102,N_48772,N_48842);
and U49103 (N_49103,N_48830,N_48996);
xnor U49104 (N_49104,N_48803,N_48823);
or U49105 (N_49105,N_48984,N_48850);
or U49106 (N_49106,N_48836,N_48755);
nor U49107 (N_49107,N_48947,N_48956);
nor U49108 (N_49108,N_48995,N_48910);
nand U49109 (N_49109,N_48779,N_48962);
nand U49110 (N_49110,N_48776,N_48751);
xnor U49111 (N_49111,N_48801,N_48840);
nor U49112 (N_49112,N_48884,N_48756);
nand U49113 (N_49113,N_48839,N_48820);
xnor U49114 (N_49114,N_48875,N_48960);
nor U49115 (N_49115,N_48966,N_48936);
nor U49116 (N_49116,N_48873,N_48791);
nand U49117 (N_49117,N_48843,N_48895);
and U49118 (N_49118,N_48782,N_48892);
or U49119 (N_49119,N_48890,N_48787);
xor U49120 (N_49120,N_48811,N_48771);
nand U49121 (N_49121,N_48903,N_48871);
nor U49122 (N_49122,N_48900,N_48994);
xnor U49123 (N_49123,N_48844,N_48880);
xor U49124 (N_49124,N_48833,N_48981);
and U49125 (N_49125,N_48827,N_48822);
and U49126 (N_49126,N_48830,N_48990);
nand U49127 (N_49127,N_48863,N_48825);
xor U49128 (N_49128,N_48824,N_48924);
nand U49129 (N_49129,N_48770,N_48815);
nand U49130 (N_49130,N_48849,N_48793);
xnor U49131 (N_49131,N_48771,N_48916);
nor U49132 (N_49132,N_48760,N_48990);
and U49133 (N_49133,N_48989,N_48980);
nor U49134 (N_49134,N_48776,N_48884);
and U49135 (N_49135,N_48952,N_48762);
and U49136 (N_49136,N_48774,N_48816);
or U49137 (N_49137,N_48958,N_48902);
or U49138 (N_49138,N_48994,N_48831);
nor U49139 (N_49139,N_48793,N_48812);
nand U49140 (N_49140,N_48869,N_48892);
and U49141 (N_49141,N_48765,N_48783);
and U49142 (N_49142,N_48816,N_48920);
and U49143 (N_49143,N_48948,N_48785);
nand U49144 (N_49144,N_48955,N_48880);
xor U49145 (N_49145,N_48787,N_48816);
or U49146 (N_49146,N_48861,N_48839);
and U49147 (N_49147,N_48840,N_48837);
or U49148 (N_49148,N_48994,N_48979);
or U49149 (N_49149,N_48973,N_48754);
nand U49150 (N_49150,N_48780,N_48786);
and U49151 (N_49151,N_48912,N_48793);
or U49152 (N_49152,N_48953,N_48892);
nor U49153 (N_49153,N_48909,N_48825);
nor U49154 (N_49154,N_48913,N_48880);
nor U49155 (N_49155,N_48755,N_48900);
or U49156 (N_49156,N_48803,N_48838);
nand U49157 (N_49157,N_48963,N_48877);
xor U49158 (N_49158,N_48880,N_48982);
and U49159 (N_49159,N_48874,N_48967);
xnor U49160 (N_49160,N_48969,N_48968);
xnor U49161 (N_49161,N_48849,N_48870);
xor U49162 (N_49162,N_48751,N_48982);
or U49163 (N_49163,N_48912,N_48825);
xnor U49164 (N_49164,N_48750,N_48999);
xnor U49165 (N_49165,N_48920,N_48899);
nand U49166 (N_49166,N_48782,N_48963);
xor U49167 (N_49167,N_48832,N_48912);
nor U49168 (N_49168,N_48864,N_48819);
or U49169 (N_49169,N_48929,N_48837);
and U49170 (N_49170,N_48916,N_48822);
or U49171 (N_49171,N_48762,N_48914);
and U49172 (N_49172,N_48759,N_48805);
nand U49173 (N_49173,N_48854,N_48784);
nand U49174 (N_49174,N_48780,N_48993);
and U49175 (N_49175,N_48847,N_48770);
and U49176 (N_49176,N_48971,N_48881);
and U49177 (N_49177,N_48814,N_48888);
nand U49178 (N_49178,N_48797,N_48909);
or U49179 (N_49179,N_48861,N_48770);
xor U49180 (N_49180,N_48948,N_48987);
nand U49181 (N_49181,N_48996,N_48978);
or U49182 (N_49182,N_48777,N_48935);
nand U49183 (N_49183,N_48992,N_48842);
nor U49184 (N_49184,N_48956,N_48869);
nor U49185 (N_49185,N_48946,N_48857);
nand U49186 (N_49186,N_48944,N_48940);
nand U49187 (N_49187,N_48871,N_48802);
xnor U49188 (N_49188,N_48785,N_48996);
nand U49189 (N_49189,N_48933,N_48757);
nor U49190 (N_49190,N_48850,N_48950);
xnor U49191 (N_49191,N_48832,N_48822);
nor U49192 (N_49192,N_48867,N_48783);
or U49193 (N_49193,N_48757,N_48899);
xor U49194 (N_49194,N_48870,N_48763);
or U49195 (N_49195,N_48915,N_48776);
nor U49196 (N_49196,N_48815,N_48961);
xor U49197 (N_49197,N_48951,N_48916);
or U49198 (N_49198,N_48918,N_48775);
xor U49199 (N_49199,N_48801,N_48780);
nand U49200 (N_49200,N_48751,N_48787);
xor U49201 (N_49201,N_48812,N_48800);
or U49202 (N_49202,N_48927,N_48837);
or U49203 (N_49203,N_48778,N_48974);
or U49204 (N_49204,N_48780,N_48791);
or U49205 (N_49205,N_48907,N_48882);
or U49206 (N_49206,N_48968,N_48841);
or U49207 (N_49207,N_48773,N_48882);
xnor U49208 (N_49208,N_48804,N_48827);
and U49209 (N_49209,N_48987,N_48969);
nor U49210 (N_49210,N_48905,N_48964);
nand U49211 (N_49211,N_48997,N_48896);
or U49212 (N_49212,N_48806,N_48888);
nor U49213 (N_49213,N_48989,N_48824);
and U49214 (N_49214,N_48811,N_48997);
nand U49215 (N_49215,N_48934,N_48842);
xnor U49216 (N_49216,N_48794,N_48946);
or U49217 (N_49217,N_48800,N_48864);
nor U49218 (N_49218,N_48981,N_48831);
and U49219 (N_49219,N_48947,N_48831);
nand U49220 (N_49220,N_48865,N_48889);
xnor U49221 (N_49221,N_48751,N_48893);
and U49222 (N_49222,N_48863,N_48937);
xnor U49223 (N_49223,N_48939,N_48836);
nand U49224 (N_49224,N_48798,N_48979);
xnor U49225 (N_49225,N_48903,N_48752);
nand U49226 (N_49226,N_48813,N_48957);
nor U49227 (N_49227,N_48837,N_48793);
and U49228 (N_49228,N_48944,N_48996);
or U49229 (N_49229,N_48804,N_48873);
nand U49230 (N_49230,N_48783,N_48869);
nor U49231 (N_49231,N_48827,N_48903);
nand U49232 (N_49232,N_48966,N_48983);
xnor U49233 (N_49233,N_48865,N_48803);
nand U49234 (N_49234,N_48848,N_48821);
xnor U49235 (N_49235,N_48859,N_48922);
nand U49236 (N_49236,N_48751,N_48825);
and U49237 (N_49237,N_48919,N_48963);
or U49238 (N_49238,N_48851,N_48946);
nand U49239 (N_49239,N_48786,N_48810);
nor U49240 (N_49240,N_48810,N_48841);
nor U49241 (N_49241,N_48771,N_48951);
nor U49242 (N_49242,N_48949,N_48892);
and U49243 (N_49243,N_48866,N_48841);
xnor U49244 (N_49244,N_48867,N_48809);
xor U49245 (N_49245,N_48807,N_48831);
nor U49246 (N_49246,N_48954,N_48895);
nor U49247 (N_49247,N_48865,N_48769);
xnor U49248 (N_49248,N_48987,N_48872);
or U49249 (N_49249,N_48868,N_48971);
nand U49250 (N_49250,N_49096,N_49231);
and U49251 (N_49251,N_49072,N_49172);
nor U49252 (N_49252,N_49039,N_49109);
nand U49253 (N_49253,N_49153,N_49022);
nor U49254 (N_49254,N_49246,N_49228);
and U49255 (N_49255,N_49210,N_49043);
or U49256 (N_49256,N_49019,N_49040);
and U49257 (N_49257,N_49171,N_49107);
and U49258 (N_49258,N_49010,N_49012);
or U49259 (N_49259,N_49178,N_49220);
nand U49260 (N_49260,N_49011,N_49121);
and U49261 (N_49261,N_49078,N_49106);
xor U49262 (N_49262,N_49196,N_49021);
and U49263 (N_49263,N_49104,N_49057);
xor U49264 (N_49264,N_49023,N_49071);
nand U49265 (N_49265,N_49005,N_49180);
or U49266 (N_49266,N_49234,N_49076);
xor U49267 (N_49267,N_49144,N_49099);
nor U49268 (N_49268,N_49214,N_49129);
or U49269 (N_49269,N_49070,N_49111);
nor U49270 (N_49270,N_49035,N_49113);
or U49271 (N_49271,N_49055,N_49002);
and U49272 (N_49272,N_49068,N_49212);
xor U49273 (N_49273,N_49173,N_49056);
or U49274 (N_49274,N_49226,N_49175);
nor U49275 (N_49275,N_49095,N_49126);
nand U49276 (N_49276,N_49045,N_49247);
and U49277 (N_49277,N_49000,N_49191);
xor U49278 (N_49278,N_49058,N_49028);
and U49279 (N_49279,N_49177,N_49026);
xnor U49280 (N_49280,N_49052,N_49051);
and U49281 (N_49281,N_49073,N_49018);
nand U49282 (N_49282,N_49193,N_49119);
and U49283 (N_49283,N_49088,N_49053);
nor U49284 (N_49284,N_49075,N_49165);
nor U49285 (N_49285,N_49067,N_49184);
or U49286 (N_49286,N_49091,N_49114);
and U49287 (N_49287,N_49050,N_49224);
and U49288 (N_49288,N_49098,N_49062);
nand U49289 (N_49289,N_49235,N_49029);
and U49290 (N_49290,N_49036,N_49080);
nand U49291 (N_49291,N_49017,N_49030);
nand U49292 (N_49292,N_49089,N_49118);
or U49293 (N_49293,N_49083,N_49239);
nand U49294 (N_49294,N_49047,N_49154);
or U49295 (N_49295,N_49189,N_49065);
nor U49296 (N_49296,N_49122,N_49031);
and U49297 (N_49297,N_49117,N_49216);
and U49298 (N_49298,N_49008,N_49157);
and U49299 (N_49299,N_49128,N_49248);
nor U49300 (N_49300,N_49219,N_49186);
nand U49301 (N_49301,N_49194,N_49102);
xnor U49302 (N_49302,N_49044,N_49218);
and U49303 (N_49303,N_49124,N_49025);
nand U49304 (N_49304,N_49140,N_49203);
xor U49305 (N_49305,N_49230,N_49201);
xnor U49306 (N_49306,N_49169,N_49241);
nor U49307 (N_49307,N_49181,N_49245);
nand U49308 (N_49308,N_49211,N_49227);
xor U49309 (N_49309,N_49166,N_49127);
or U49310 (N_49310,N_49131,N_49027);
nand U49311 (N_49311,N_49134,N_49249);
or U49312 (N_49312,N_49199,N_49105);
or U49313 (N_49313,N_49158,N_49074);
or U49314 (N_49314,N_49229,N_49185);
nand U49315 (N_49315,N_49160,N_49207);
and U49316 (N_49316,N_49009,N_49132);
nand U49317 (N_49317,N_49142,N_49222);
nor U49318 (N_49318,N_49032,N_49146);
and U49319 (N_49319,N_49206,N_49110);
and U49320 (N_49320,N_49163,N_49174);
xnor U49321 (N_49321,N_49094,N_49108);
and U49322 (N_49322,N_49200,N_49188);
or U49323 (N_49323,N_49152,N_49197);
and U49324 (N_49324,N_49167,N_49164);
and U49325 (N_49325,N_49033,N_49014);
or U49326 (N_49326,N_49244,N_49112);
or U49327 (N_49327,N_49020,N_49084);
or U49328 (N_49328,N_49037,N_49209);
or U49329 (N_49329,N_49147,N_49069);
nor U49330 (N_49330,N_49048,N_49149);
and U49331 (N_49331,N_49046,N_49015);
and U49332 (N_49332,N_49064,N_49097);
xor U49333 (N_49333,N_49202,N_49170);
and U49334 (N_49334,N_49100,N_49049);
nand U49335 (N_49335,N_49139,N_49116);
nand U49336 (N_49336,N_49162,N_49133);
nor U49337 (N_49337,N_49238,N_49081);
nand U49338 (N_49338,N_49087,N_49183);
nor U49339 (N_49339,N_49063,N_49092);
and U49340 (N_49340,N_49198,N_49013);
and U49341 (N_49341,N_49115,N_49205);
nand U49342 (N_49342,N_49217,N_49120);
and U49343 (N_49343,N_49093,N_49077);
xnor U49344 (N_49344,N_49061,N_49066);
xor U49345 (N_49345,N_49060,N_49232);
nand U49346 (N_49346,N_49240,N_49101);
xnor U49347 (N_49347,N_49190,N_49042);
xnor U49348 (N_49348,N_49024,N_49242);
or U49349 (N_49349,N_49156,N_49138);
or U49350 (N_49350,N_49001,N_49213);
xnor U49351 (N_49351,N_49145,N_49237);
xnor U49352 (N_49352,N_49137,N_49192);
or U49353 (N_49353,N_49215,N_49155);
nand U49354 (N_49354,N_49243,N_49233);
xnor U49355 (N_49355,N_49176,N_49208);
nor U49356 (N_49356,N_49086,N_49016);
nand U49357 (N_49357,N_49143,N_49182);
nand U49358 (N_49358,N_49079,N_49225);
nor U49359 (N_49359,N_49161,N_49195);
nand U49360 (N_49360,N_49103,N_49003);
xnor U49361 (N_49361,N_49159,N_49136);
or U49362 (N_49362,N_49123,N_49151);
xnor U49363 (N_49363,N_49148,N_49236);
and U49364 (N_49364,N_49082,N_49054);
or U49365 (N_49365,N_49223,N_49125);
nor U49366 (N_49366,N_49007,N_49085);
and U49367 (N_49367,N_49059,N_49150);
and U49368 (N_49368,N_49041,N_49038);
or U49369 (N_49369,N_49221,N_49179);
and U49370 (N_49370,N_49130,N_49168);
xor U49371 (N_49371,N_49004,N_49204);
nor U49372 (N_49372,N_49187,N_49006);
nor U49373 (N_49373,N_49135,N_49090);
nor U49374 (N_49374,N_49141,N_49034);
and U49375 (N_49375,N_49020,N_49233);
and U49376 (N_49376,N_49070,N_49236);
xnor U49377 (N_49377,N_49225,N_49150);
nand U49378 (N_49378,N_49089,N_49022);
xor U49379 (N_49379,N_49030,N_49130);
and U49380 (N_49380,N_49011,N_49027);
and U49381 (N_49381,N_49196,N_49205);
nor U49382 (N_49382,N_49132,N_49240);
and U49383 (N_49383,N_49043,N_49056);
and U49384 (N_49384,N_49106,N_49148);
xor U49385 (N_49385,N_49188,N_49115);
nor U49386 (N_49386,N_49029,N_49148);
or U49387 (N_49387,N_49105,N_49111);
nand U49388 (N_49388,N_49131,N_49146);
nor U49389 (N_49389,N_49133,N_49128);
nor U49390 (N_49390,N_49241,N_49123);
and U49391 (N_49391,N_49055,N_49216);
xor U49392 (N_49392,N_49111,N_49148);
or U49393 (N_49393,N_49069,N_49168);
or U49394 (N_49394,N_49226,N_49219);
nand U49395 (N_49395,N_49181,N_49213);
xnor U49396 (N_49396,N_49214,N_49166);
and U49397 (N_49397,N_49148,N_49152);
xnor U49398 (N_49398,N_49112,N_49170);
nor U49399 (N_49399,N_49000,N_49201);
xnor U49400 (N_49400,N_49144,N_49129);
xor U49401 (N_49401,N_49164,N_49143);
nand U49402 (N_49402,N_49215,N_49141);
and U49403 (N_49403,N_49139,N_49130);
xor U49404 (N_49404,N_49082,N_49020);
or U49405 (N_49405,N_49073,N_49189);
and U49406 (N_49406,N_49210,N_49228);
and U49407 (N_49407,N_49146,N_49136);
or U49408 (N_49408,N_49022,N_49101);
xor U49409 (N_49409,N_49170,N_49185);
xor U49410 (N_49410,N_49215,N_49082);
nand U49411 (N_49411,N_49003,N_49163);
or U49412 (N_49412,N_49149,N_49141);
or U49413 (N_49413,N_49012,N_49000);
xor U49414 (N_49414,N_49236,N_49142);
xor U49415 (N_49415,N_49237,N_49229);
xnor U49416 (N_49416,N_49219,N_49182);
nor U49417 (N_49417,N_49023,N_49243);
nor U49418 (N_49418,N_49121,N_49229);
and U49419 (N_49419,N_49232,N_49111);
nand U49420 (N_49420,N_49029,N_49146);
nand U49421 (N_49421,N_49162,N_49186);
or U49422 (N_49422,N_49246,N_49209);
or U49423 (N_49423,N_49170,N_49190);
nand U49424 (N_49424,N_49006,N_49177);
xor U49425 (N_49425,N_49206,N_49012);
or U49426 (N_49426,N_49086,N_49073);
or U49427 (N_49427,N_49160,N_49132);
xor U49428 (N_49428,N_49091,N_49127);
or U49429 (N_49429,N_49153,N_49047);
nor U49430 (N_49430,N_49174,N_49006);
xor U49431 (N_49431,N_49000,N_49014);
nor U49432 (N_49432,N_49023,N_49053);
nor U49433 (N_49433,N_49014,N_49096);
xnor U49434 (N_49434,N_49072,N_49047);
and U49435 (N_49435,N_49053,N_49001);
xor U49436 (N_49436,N_49182,N_49026);
xnor U49437 (N_49437,N_49098,N_49229);
nor U49438 (N_49438,N_49162,N_49114);
xor U49439 (N_49439,N_49215,N_49145);
nand U49440 (N_49440,N_49199,N_49223);
nand U49441 (N_49441,N_49095,N_49178);
nor U49442 (N_49442,N_49116,N_49007);
nor U49443 (N_49443,N_49043,N_49186);
xor U49444 (N_49444,N_49072,N_49178);
nand U49445 (N_49445,N_49206,N_49038);
nor U49446 (N_49446,N_49151,N_49160);
nor U49447 (N_49447,N_49146,N_49112);
xnor U49448 (N_49448,N_49197,N_49057);
nand U49449 (N_49449,N_49225,N_49230);
nand U49450 (N_49450,N_49090,N_49153);
nor U49451 (N_49451,N_49066,N_49018);
nand U49452 (N_49452,N_49106,N_49053);
xnor U49453 (N_49453,N_49176,N_49232);
nor U49454 (N_49454,N_49063,N_49232);
nor U49455 (N_49455,N_49043,N_49144);
nor U49456 (N_49456,N_49062,N_49140);
nor U49457 (N_49457,N_49234,N_49135);
nand U49458 (N_49458,N_49137,N_49058);
xnor U49459 (N_49459,N_49028,N_49232);
and U49460 (N_49460,N_49102,N_49205);
nand U49461 (N_49461,N_49113,N_49067);
nand U49462 (N_49462,N_49174,N_49199);
xor U49463 (N_49463,N_49172,N_49026);
nand U49464 (N_49464,N_49072,N_49057);
nand U49465 (N_49465,N_49000,N_49082);
xnor U49466 (N_49466,N_49197,N_49148);
nand U49467 (N_49467,N_49204,N_49189);
or U49468 (N_49468,N_49023,N_49045);
and U49469 (N_49469,N_49103,N_49205);
nand U49470 (N_49470,N_49178,N_49171);
nand U49471 (N_49471,N_49184,N_49121);
or U49472 (N_49472,N_49126,N_49130);
and U49473 (N_49473,N_49009,N_49099);
or U49474 (N_49474,N_49049,N_49214);
or U49475 (N_49475,N_49057,N_49133);
xnor U49476 (N_49476,N_49029,N_49130);
nor U49477 (N_49477,N_49059,N_49136);
nor U49478 (N_49478,N_49139,N_49092);
xor U49479 (N_49479,N_49033,N_49194);
or U49480 (N_49480,N_49164,N_49238);
xnor U49481 (N_49481,N_49013,N_49046);
xor U49482 (N_49482,N_49050,N_49069);
or U49483 (N_49483,N_49217,N_49233);
nor U49484 (N_49484,N_49124,N_49194);
nand U49485 (N_49485,N_49205,N_49064);
or U49486 (N_49486,N_49245,N_49043);
and U49487 (N_49487,N_49119,N_49231);
nand U49488 (N_49488,N_49180,N_49215);
xnor U49489 (N_49489,N_49030,N_49191);
and U49490 (N_49490,N_49043,N_49247);
or U49491 (N_49491,N_49248,N_49019);
and U49492 (N_49492,N_49157,N_49148);
xnor U49493 (N_49493,N_49059,N_49139);
or U49494 (N_49494,N_49122,N_49044);
nor U49495 (N_49495,N_49107,N_49056);
or U49496 (N_49496,N_49249,N_49219);
and U49497 (N_49497,N_49031,N_49194);
xnor U49498 (N_49498,N_49132,N_49172);
xnor U49499 (N_49499,N_49109,N_49022);
and U49500 (N_49500,N_49378,N_49263);
xor U49501 (N_49501,N_49377,N_49396);
or U49502 (N_49502,N_49340,N_49330);
and U49503 (N_49503,N_49269,N_49370);
nor U49504 (N_49504,N_49350,N_49275);
nand U49505 (N_49505,N_49361,N_49357);
nor U49506 (N_49506,N_49260,N_49472);
or U49507 (N_49507,N_49408,N_49446);
or U49508 (N_49508,N_49352,N_49414);
or U49509 (N_49509,N_49441,N_49462);
xor U49510 (N_49510,N_49264,N_49299);
nor U49511 (N_49511,N_49401,N_49322);
and U49512 (N_49512,N_49316,N_49307);
xor U49513 (N_49513,N_49418,N_49379);
nor U49514 (N_49514,N_49320,N_49423);
xor U49515 (N_49515,N_49256,N_49298);
xnor U49516 (N_49516,N_49312,N_49442);
or U49517 (N_49517,N_49397,N_49459);
nand U49518 (N_49518,N_49465,N_49427);
and U49519 (N_49519,N_49284,N_49468);
or U49520 (N_49520,N_49476,N_49280);
xnor U49521 (N_49521,N_49403,N_49258);
nor U49522 (N_49522,N_49317,N_49411);
nor U49523 (N_49523,N_49436,N_49486);
or U49524 (N_49524,N_49341,N_49376);
nand U49525 (N_49525,N_49428,N_49444);
and U49526 (N_49526,N_49419,N_49495);
or U49527 (N_49527,N_49321,N_49450);
or U49528 (N_49528,N_49254,N_49416);
nand U49529 (N_49529,N_49466,N_49457);
or U49530 (N_49530,N_49348,N_49386);
or U49531 (N_49531,N_49473,N_49480);
nand U49532 (N_49532,N_49309,N_49359);
or U49533 (N_49533,N_49366,N_49343);
and U49534 (N_49534,N_49491,N_49399);
or U49535 (N_49535,N_49400,N_49432);
nand U49536 (N_49536,N_49347,N_49328);
nand U49537 (N_49537,N_49291,N_49259);
or U49538 (N_49538,N_49308,N_49496);
nor U49539 (N_49539,N_49431,N_49406);
or U49540 (N_49540,N_49461,N_49391);
xnor U49541 (N_49541,N_49478,N_49329);
and U49542 (N_49542,N_49368,N_49374);
and U49543 (N_49543,N_49294,N_49314);
nor U49544 (N_49544,N_49306,N_49365);
nor U49545 (N_49545,N_49315,N_49429);
nor U49546 (N_49546,N_49296,N_49288);
nand U49547 (N_49547,N_49326,N_49430);
xnor U49548 (N_49548,N_49282,N_49498);
xnor U49549 (N_49549,N_49455,N_49351);
or U49550 (N_49550,N_49251,N_49272);
nand U49551 (N_49551,N_49354,N_49273);
nor U49552 (N_49552,N_49477,N_49485);
and U49553 (N_49553,N_49290,N_49448);
nand U49554 (N_49554,N_49393,N_49475);
or U49555 (N_49555,N_49277,N_49464);
and U49556 (N_49556,N_49369,N_49460);
or U49557 (N_49557,N_49454,N_49360);
nand U49558 (N_49558,N_49382,N_49426);
nor U49559 (N_49559,N_49482,N_49481);
and U49560 (N_49560,N_49458,N_49452);
or U49561 (N_49561,N_49345,N_49489);
nor U49562 (N_49562,N_49278,N_49437);
and U49563 (N_49563,N_49453,N_49479);
and U49564 (N_49564,N_49404,N_49388);
or U49565 (N_49565,N_49470,N_49385);
nor U49566 (N_49566,N_49331,N_49367);
and U49567 (N_49567,N_49443,N_49415);
and U49568 (N_49568,N_49405,N_49250);
nand U49569 (N_49569,N_49286,N_49355);
nand U49570 (N_49570,N_49371,N_49261);
or U49571 (N_49571,N_49417,N_49262);
and U49572 (N_49572,N_49467,N_49305);
or U49573 (N_49573,N_49300,N_49313);
and U49574 (N_49574,N_49325,N_49494);
nand U49575 (N_49575,N_49353,N_49412);
nor U49576 (N_49576,N_49270,N_49389);
nand U49577 (N_49577,N_49449,N_49497);
xor U49578 (N_49578,N_49488,N_49380);
nand U49579 (N_49579,N_49302,N_49279);
xnor U49580 (N_49580,N_49289,N_49281);
or U49581 (N_49581,N_49338,N_49363);
nand U49582 (N_49582,N_49292,N_49375);
nor U49583 (N_49583,N_49358,N_49346);
and U49584 (N_49584,N_49422,N_49407);
or U49585 (N_49585,N_49283,N_49297);
nand U49586 (N_49586,N_49333,N_49394);
and U49587 (N_49587,N_49356,N_49342);
nand U49588 (N_49588,N_49493,N_49276);
nor U49589 (N_49589,N_49271,N_49257);
or U49590 (N_49590,N_49372,N_49373);
nor U49591 (N_49591,N_49484,N_49253);
or U49592 (N_49592,N_49487,N_49295);
nor U49593 (N_49593,N_49438,N_49324);
nor U49594 (N_49594,N_49255,N_49327);
and U49595 (N_49595,N_49349,N_49310);
nand U49596 (N_49596,N_49364,N_49252);
xnor U49597 (N_49597,N_49344,N_49274);
or U49598 (N_49598,N_49335,N_49469);
xor U49599 (N_49599,N_49336,N_49413);
xor U49600 (N_49600,N_49409,N_49337);
xnor U49601 (N_49601,N_49445,N_49395);
nor U49602 (N_49602,N_49339,N_49433);
nand U49603 (N_49603,N_49435,N_49266);
or U49604 (N_49604,N_49392,N_49483);
or U49605 (N_49605,N_49293,N_49285);
nor U49606 (N_49606,N_49383,N_49387);
or U49607 (N_49607,N_49323,N_49402);
xnor U49608 (N_49608,N_49447,N_49424);
nand U49609 (N_49609,N_49362,N_49474);
and U49610 (N_49610,N_49304,N_49492);
nand U49611 (N_49611,N_49471,N_49439);
nand U49612 (N_49612,N_49332,N_49268);
or U49613 (N_49613,N_49421,N_49301);
or U49614 (N_49614,N_49398,N_49456);
nor U49615 (N_49615,N_49265,N_49490);
nor U49616 (N_49616,N_49381,N_49499);
or U49617 (N_49617,N_49303,N_49434);
and U49618 (N_49618,N_49420,N_49425);
nor U49619 (N_49619,N_49390,N_49440);
xnor U49620 (N_49620,N_49311,N_49451);
or U49621 (N_49621,N_49410,N_49463);
nor U49622 (N_49622,N_49318,N_49319);
nor U49623 (N_49623,N_49267,N_49287);
and U49624 (N_49624,N_49334,N_49384);
nor U49625 (N_49625,N_49349,N_49469);
nor U49626 (N_49626,N_49381,N_49490);
and U49627 (N_49627,N_49470,N_49442);
nor U49628 (N_49628,N_49297,N_49306);
xnor U49629 (N_49629,N_49379,N_49387);
nand U49630 (N_49630,N_49269,N_49448);
xor U49631 (N_49631,N_49259,N_49270);
nand U49632 (N_49632,N_49356,N_49434);
nor U49633 (N_49633,N_49356,N_49497);
and U49634 (N_49634,N_49456,N_49452);
and U49635 (N_49635,N_49477,N_49437);
nor U49636 (N_49636,N_49390,N_49337);
nand U49637 (N_49637,N_49337,N_49386);
or U49638 (N_49638,N_49416,N_49268);
and U49639 (N_49639,N_49432,N_49273);
nor U49640 (N_49640,N_49292,N_49367);
nand U49641 (N_49641,N_49382,N_49260);
nor U49642 (N_49642,N_49352,N_49474);
nor U49643 (N_49643,N_49492,N_49488);
nor U49644 (N_49644,N_49280,N_49264);
nand U49645 (N_49645,N_49404,N_49443);
or U49646 (N_49646,N_49339,N_49470);
nand U49647 (N_49647,N_49443,N_49364);
xor U49648 (N_49648,N_49487,N_49328);
nor U49649 (N_49649,N_49467,N_49388);
and U49650 (N_49650,N_49288,N_49282);
nand U49651 (N_49651,N_49417,N_49473);
or U49652 (N_49652,N_49349,N_49340);
xnor U49653 (N_49653,N_49265,N_49411);
nor U49654 (N_49654,N_49470,N_49282);
or U49655 (N_49655,N_49372,N_49400);
and U49656 (N_49656,N_49260,N_49306);
nand U49657 (N_49657,N_49413,N_49325);
nand U49658 (N_49658,N_49416,N_49368);
xnor U49659 (N_49659,N_49312,N_49349);
or U49660 (N_49660,N_49427,N_49387);
and U49661 (N_49661,N_49492,N_49323);
xor U49662 (N_49662,N_49460,N_49361);
nand U49663 (N_49663,N_49332,N_49308);
and U49664 (N_49664,N_49370,N_49304);
or U49665 (N_49665,N_49312,N_49276);
nor U49666 (N_49666,N_49265,N_49466);
nor U49667 (N_49667,N_49490,N_49253);
nand U49668 (N_49668,N_49360,N_49410);
and U49669 (N_49669,N_49442,N_49281);
nand U49670 (N_49670,N_49263,N_49317);
nand U49671 (N_49671,N_49260,N_49288);
nand U49672 (N_49672,N_49416,N_49390);
xor U49673 (N_49673,N_49350,N_49401);
xnor U49674 (N_49674,N_49289,N_49412);
nor U49675 (N_49675,N_49338,N_49487);
nor U49676 (N_49676,N_49349,N_49319);
and U49677 (N_49677,N_49333,N_49460);
xnor U49678 (N_49678,N_49254,N_49324);
xor U49679 (N_49679,N_49410,N_49389);
xnor U49680 (N_49680,N_49345,N_49444);
nor U49681 (N_49681,N_49369,N_49456);
nand U49682 (N_49682,N_49415,N_49283);
and U49683 (N_49683,N_49324,N_49306);
nor U49684 (N_49684,N_49345,N_49427);
nand U49685 (N_49685,N_49358,N_49330);
nand U49686 (N_49686,N_49262,N_49253);
and U49687 (N_49687,N_49290,N_49393);
and U49688 (N_49688,N_49358,N_49457);
or U49689 (N_49689,N_49404,N_49393);
xnor U49690 (N_49690,N_49332,N_49258);
or U49691 (N_49691,N_49370,N_49445);
nand U49692 (N_49692,N_49405,N_49451);
xor U49693 (N_49693,N_49492,N_49271);
nor U49694 (N_49694,N_49391,N_49297);
and U49695 (N_49695,N_49281,N_49359);
nor U49696 (N_49696,N_49378,N_49335);
nand U49697 (N_49697,N_49414,N_49361);
and U49698 (N_49698,N_49410,N_49443);
xnor U49699 (N_49699,N_49470,N_49392);
and U49700 (N_49700,N_49378,N_49480);
and U49701 (N_49701,N_49487,N_49459);
or U49702 (N_49702,N_49438,N_49336);
nand U49703 (N_49703,N_49285,N_49365);
nand U49704 (N_49704,N_49466,N_49284);
or U49705 (N_49705,N_49368,N_49265);
xnor U49706 (N_49706,N_49304,N_49313);
or U49707 (N_49707,N_49475,N_49497);
nor U49708 (N_49708,N_49267,N_49339);
or U49709 (N_49709,N_49490,N_49369);
nor U49710 (N_49710,N_49407,N_49388);
or U49711 (N_49711,N_49339,N_49257);
nand U49712 (N_49712,N_49277,N_49480);
xnor U49713 (N_49713,N_49384,N_49380);
nor U49714 (N_49714,N_49431,N_49408);
nand U49715 (N_49715,N_49326,N_49347);
xnor U49716 (N_49716,N_49311,N_49321);
nor U49717 (N_49717,N_49441,N_49453);
or U49718 (N_49718,N_49275,N_49356);
nand U49719 (N_49719,N_49314,N_49324);
xor U49720 (N_49720,N_49326,N_49332);
nand U49721 (N_49721,N_49495,N_49251);
nor U49722 (N_49722,N_49409,N_49300);
nor U49723 (N_49723,N_49320,N_49435);
xnor U49724 (N_49724,N_49421,N_49362);
or U49725 (N_49725,N_49372,N_49269);
or U49726 (N_49726,N_49431,N_49482);
xnor U49727 (N_49727,N_49392,N_49347);
nor U49728 (N_49728,N_49367,N_49267);
and U49729 (N_49729,N_49299,N_49307);
or U49730 (N_49730,N_49304,N_49459);
xnor U49731 (N_49731,N_49347,N_49493);
nand U49732 (N_49732,N_49294,N_49413);
nor U49733 (N_49733,N_49443,N_49278);
or U49734 (N_49734,N_49455,N_49441);
and U49735 (N_49735,N_49398,N_49353);
and U49736 (N_49736,N_49396,N_49270);
or U49737 (N_49737,N_49262,N_49430);
nor U49738 (N_49738,N_49394,N_49437);
or U49739 (N_49739,N_49272,N_49293);
or U49740 (N_49740,N_49270,N_49421);
xnor U49741 (N_49741,N_49307,N_49446);
and U49742 (N_49742,N_49357,N_49405);
xnor U49743 (N_49743,N_49362,N_49300);
nand U49744 (N_49744,N_49325,N_49264);
or U49745 (N_49745,N_49432,N_49305);
xnor U49746 (N_49746,N_49357,N_49492);
and U49747 (N_49747,N_49296,N_49353);
or U49748 (N_49748,N_49382,N_49407);
or U49749 (N_49749,N_49424,N_49409);
and U49750 (N_49750,N_49512,N_49659);
and U49751 (N_49751,N_49669,N_49652);
or U49752 (N_49752,N_49601,N_49570);
nor U49753 (N_49753,N_49510,N_49670);
and U49754 (N_49754,N_49746,N_49720);
and U49755 (N_49755,N_49710,N_49711);
and U49756 (N_49756,N_49591,N_49557);
or U49757 (N_49757,N_49515,N_49509);
nand U49758 (N_49758,N_49636,N_49641);
nand U49759 (N_49759,N_49527,N_49598);
or U49760 (N_49760,N_49645,N_49545);
and U49761 (N_49761,N_49686,N_49747);
and U49762 (N_49762,N_49602,N_49731);
xnor U49763 (N_49763,N_49648,N_49595);
xor U49764 (N_49764,N_49658,N_49718);
xor U49765 (N_49765,N_49672,N_49736);
xnor U49766 (N_49766,N_49541,N_49654);
nand U49767 (N_49767,N_49728,N_49631);
or U49768 (N_49768,N_49657,N_49574);
or U49769 (N_49769,N_49691,N_49576);
or U49770 (N_49770,N_49647,N_49707);
nor U49771 (N_49771,N_49606,N_49610);
nor U49772 (N_49772,N_49563,N_49725);
xor U49773 (N_49773,N_49585,N_49639);
xor U49774 (N_49774,N_49529,N_49705);
xor U49775 (N_49775,N_49717,N_49740);
and U49776 (N_49776,N_49612,N_49546);
and U49777 (N_49777,N_49554,N_49703);
or U49778 (N_49778,N_49644,N_49583);
nand U49779 (N_49779,N_49503,N_49607);
xor U49780 (N_49780,N_49558,N_49562);
or U49781 (N_49781,N_49540,N_49532);
nor U49782 (N_49782,N_49656,N_49568);
nor U49783 (N_49783,N_49613,N_49698);
xnor U49784 (N_49784,N_49716,N_49519);
and U49785 (N_49785,N_49697,N_49655);
and U49786 (N_49786,N_49577,N_49667);
and U49787 (N_49787,N_49664,N_49559);
or U49788 (N_49788,N_49632,N_49522);
or U49789 (N_49789,N_49708,N_49688);
or U49790 (N_49790,N_49500,N_49676);
nand U49791 (N_49791,N_49537,N_49694);
xor U49792 (N_49792,N_49525,N_49712);
and U49793 (N_49793,N_49508,N_49506);
or U49794 (N_49794,N_49704,N_49526);
nor U49795 (N_49795,N_49550,N_49682);
and U49796 (N_49796,N_49651,N_49739);
or U49797 (N_49797,N_49623,N_49617);
nor U49798 (N_49798,N_49530,N_49596);
nand U49799 (N_49799,N_49637,N_49600);
and U49800 (N_49800,N_49567,N_49531);
xor U49801 (N_49801,N_49744,N_49671);
xnor U49802 (N_49802,N_49544,N_49661);
nand U49803 (N_49803,N_49502,N_49706);
nand U49804 (N_49804,N_49517,N_49653);
and U49805 (N_49805,N_49719,N_49592);
xor U49806 (N_49806,N_49588,N_49741);
nand U49807 (N_49807,N_49735,N_49582);
nand U49808 (N_49808,N_49679,N_49742);
and U49809 (N_49809,N_49650,N_49553);
or U49810 (N_49810,N_49561,N_49572);
nor U49811 (N_49811,N_49727,N_49749);
nor U49812 (N_49812,N_49660,N_49638);
nand U49813 (N_49813,N_49732,N_49713);
and U49814 (N_49814,N_49681,N_49628);
nor U49815 (N_49815,N_49662,N_49715);
nor U49816 (N_49816,N_49643,N_49709);
or U49817 (N_49817,N_49624,N_49714);
nand U49818 (N_49818,N_49677,N_49565);
or U49819 (N_49819,N_49513,N_49528);
or U49820 (N_49820,N_49555,N_49571);
or U49821 (N_49821,N_49689,N_49594);
and U49822 (N_49822,N_49722,N_49552);
nor U49823 (N_49823,N_49548,N_49678);
or U49824 (N_49824,N_49587,N_49635);
nand U49825 (N_49825,N_49578,N_49683);
nor U49826 (N_49826,N_49608,N_49733);
or U49827 (N_49827,N_49564,N_49673);
nor U49828 (N_49828,N_49573,N_49543);
nand U49829 (N_49829,N_49629,N_49580);
nor U49830 (N_49830,N_49615,N_49748);
xor U49831 (N_49831,N_49685,N_49590);
nand U49832 (N_49832,N_49566,N_49724);
nand U49833 (N_49833,N_49589,N_49730);
and U49834 (N_49834,N_49521,N_49622);
or U49835 (N_49835,N_49663,N_49702);
nand U49836 (N_49836,N_49699,N_49619);
nand U49837 (N_49837,N_49723,N_49524);
or U49838 (N_49838,N_49640,N_49701);
or U49839 (N_49839,N_49535,N_49616);
nor U49840 (N_49840,N_49533,N_49507);
and U49841 (N_49841,N_49625,N_49556);
nand U49842 (N_49842,N_49549,N_49633);
and U49843 (N_49843,N_49693,N_49581);
nor U49844 (N_49844,N_49579,N_49551);
or U49845 (N_49845,N_49700,N_49649);
or U49846 (N_49846,N_49626,N_49627);
or U49847 (N_49847,N_49696,N_49611);
and U49848 (N_49848,N_49609,N_49534);
nor U49849 (N_49849,N_49618,N_49603);
xor U49850 (N_49850,N_49504,N_49620);
xnor U49851 (N_49851,N_49584,N_49674);
or U49852 (N_49852,N_49547,N_49634);
xnor U49853 (N_49853,N_49734,N_49687);
xnor U49854 (N_49854,N_49726,N_49738);
and U49855 (N_49855,N_49520,N_49597);
nand U49856 (N_49856,N_49586,N_49604);
nand U49857 (N_49857,N_49692,N_49599);
or U49858 (N_49858,N_49536,N_49539);
nand U49859 (N_49859,N_49523,N_49514);
and U49860 (N_49860,N_49501,N_49695);
or U49861 (N_49861,N_49743,N_49518);
or U49862 (N_49862,N_49721,N_49505);
nor U49863 (N_49863,N_49569,N_49614);
or U49864 (N_49864,N_49511,N_49680);
xnor U49865 (N_49865,N_49630,N_49666);
xor U49866 (N_49866,N_49668,N_49665);
nor U49867 (N_49867,N_49737,N_49675);
and U49868 (N_49868,N_49745,N_49684);
nor U49869 (N_49869,N_49646,N_49729);
and U49870 (N_49870,N_49516,N_49621);
or U49871 (N_49871,N_49593,N_49560);
nand U49872 (N_49872,N_49605,N_49642);
or U49873 (N_49873,N_49690,N_49538);
nand U49874 (N_49874,N_49575,N_49542);
nor U49875 (N_49875,N_49658,N_49678);
and U49876 (N_49876,N_49684,N_49719);
nand U49877 (N_49877,N_49723,N_49745);
nor U49878 (N_49878,N_49748,N_49556);
nand U49879 (N_49879,N_49616,N_49747);
xor U49880 (N_49880,N_49731,N_49674);
or U49881 (N_49881,N_49662,N_49529);
or U49882 (N_49882,N_49720,N_49667);
and U49883 (N_49883,N_49529,N_49695);
nand U49884 (N_49884,N_49601,N_49569);
and U49885 (N_49885,N_49594,N_49691);
nor U49886 (N_49886,N_49678,N_49692);
nor U49887 (N_49887,N_49548,N_49527);
nand U49888 (N_49888,N_49692,N_49654);
nor U49889 (N_49889,N_49568,N_49659);
nor U49890 (N_49890,N_49504,N_49703);
xnor U49891 (N_49891,N_49511,N_49690);
nand U49892 (N_49892,N_49554,N_49608);
xor U49893 (N_49893,N_49632,N_49605);
nor U49894 (N_49894,N_49688,N_49723);
nor U49895 (N_49895,N_49654,N_49575);
or U49896 (N_49896,N_49599,N_49620);
and U49897 (N_49897,N_49712,N_49508);
nand U49898 (N_49898,N_49684,N_49501);
xnor U49899 (N_49899,N_49615,N_49681);
nor U49900 (N_49900,N_49721,N_49625);
xor U49901 (N_49901,N_49692,N_49669);
xnor U49902 (N_49902,N_49629,N_49534);
nand U49903 (N_49903,N_49615,N_49715);
nor U49904 (N_49904,N_49548,N_49583);
and U49905 (N_49905,N_49587,N_49688);
nand U49906 (N_49906,N_49673,N_49666);
nand U49907 (N_49907,N_49621,N_49614);
or U49908 (N_49908,N_49727,N_49719);
and U49909 (N_49909,N_49568,N_49576);
xnor U49910 (N_49910,N_49623,N_49612);
nand U49911 (N_49911,N_49525,N_49566);
and U49912 (N_49912,N_49634,N_49643);
nor U49913 (N_49913,N_49620,N_49605);
xnor U49914 (N_49914,N_49521,N_49534);
and U49915 (N_49915,N_49694,N_49629);
or U49916 (N_49916,N_49647,N_49569);
xnor U49917 (N_49917,N_49675,N_49681);
nand U49918 (N_49918,N_49661,N_49654);
or U49919 (N_49919,N_49556,N_49513);
xor U49920 (N_49920,N_49602,N_49589);
xnor U49921 (N_49921,N_49747,N_49738);
nand U49922 (N_49922,N_49653,N_49556);
nor U49923 (N_49923,N_49516,N_49550);
nor U49924 (N_49924,N_49610,N_49718);
nand U49925 (N_49925,N_49655,N_49708);
or U49926 (N_49926,N_49610,N_49503);
nand U49927 (N_49927,N_49659,N_49602);
xnor U49928 (N_49928,N_49749,N_49741);
nor U49929 (N_49929,N_49568,N_49537);
nand U49930 (N_49930,N_49687,N_49527);
and U49931 (N_49931,N_49707,N_49705);
and U49932 (N_49932,N_49697,N_49624);
and U49933 (N_49933,N_49581,N_49641);
and U49934 (N_49934,N_49611,N_49636);
nand U49935 (N_49935,N_49704,N_49528);
nand U49936 (N_49936,N_49679,N_49588);
nand U49937 (N_49937,N_49570,N_49563);
and U49938 (N_49938,N_49536,N_49740);
nor U49939 (N_49939,N_49684,N_49505);
nand U49940 (N_49940,N_49699,N_49678);
nor U49941 (N_49941,N_49644,N_49651);
nor U49942 (N_49942,N_49749,N_49640);
and U49943 (N_49943,N_49501,N_49686);
nand U49944 (N_49944,N_49622,N_49518);
or U49945 (N_49945,N_49556,N_49614);
nand U49946 (N_49946,N_49657,N_49699);
and U49947 (N_49947,N_49664,N_49563);
xor U49948 (N_49948,N_49701,N_49607);
nand U49949 (N_49949,N_49526,N_49739);
xnor U49950 (N_49950,N_49667,N_49608);
nand U49951 (N_49951,N_49568,N_49711);
and U49952 (N_49952,N_49636,N_49680);
or U49953 (N_49953,N_49643,N_49599);
nor U49954 (N_49954,N_49637,N_49685);
or U49955 (N_49955,N_49694,N_49701);
nor U49956 (N_49956,N_49502,N_49734);
nand U49957 (N_49957,N_49583,N_49691);
nor U49958 (N_49958,N_49731,N_49721);
xnor U49959 (N_49959,N_49606,N_49663);
nor U49960 (N_49960,N_49585,N_49511);
nor U49961 (N_49961,N_49509,N_49601);
and U49962 (N_49962,N_49515,N_49690);
or U49963 (N_49963,N_49608,N_49632);
and U49964 (N_49964,N_49710,N_49689);
and U49965 (N_49965,N_49517,N_49600);
xnor U49966 (N_49966,N_49608,N_49601);
nand U49967 (N_49967,N_49699,N_49709);
nand U49968 (N_49968,N_49544,N_49574);
nor U49969 (N_49969,N_49630,N_49635);
or U49970 (N_49970,N_49606,N_49672);
nor U49971 (N_49971,N_49586,N_49710);
xnor U49972 (N_49972,N_49569,N_49586);
and U49973 (N_49973,N_49685,N_49623);
or U49974 (N_49974,N_49687,N_49515);
or U49975 (N_49975,N_49717,N_49645);
nand U49976 (N_49976,N_49505,N_49529);
or U49977 (N_49977,N_49657,N_49555);
nand U49978 (N_49978,N_49537,N_49625);
nor U49979 (N_49979,N_49593,N_49673);
xor U49980 (N_49980,N_49583,N_49636);
nor U49981 (N_49981,N_49712,N_49749);
or U49982 (N_49982,N_49514,N_49742);
nor U49983 (N_49983,N_49529,N_49644);
nand U49984 (N_49984,N_49641,N_49626);
nand U49985 (N_49985,N_49609,N_49677);
or U49986 (N_49986,N_49500,N_49571);
and U49987 (N_49987,N_49671,N_49627);
nand U49988 (N_49988,N_49519,N_49692);
nand U49989 (N_49989,N_49746,N_49649);
and U49990 (N_49990,N_49634,N_49699);
xnor U49991 (N_49991,N_49580,N_49518);
or U49992 (N_49992,N_49580,N_49673);
nand U49993 (N_49993,N_49612,N_49539);
and U49994 (N_49994,N_49703,N_49574);
and U49995 (N_49995,N_49627,N_49719);
nor U49996 (N_49996,N_49541,N_49663);
and U49997 (N_49997,N_49595,N_49621);
nand U49998 (N_49998,N_49617,N_49575);
and U49999 (N_49999,N_49652,N_49520);
and UO_0 (O_0,N_49752,N_49789);
or UO_1 (O_1,N_49940,N_49819);
nor UO_2 (O_2,N_49787,N_49923);
or UO_3 (O_3,N_49790,N_49841);
xor UO_4 (O_4,N_49769,N_49894);
and UO_5 (O_5,N_49813,N_49956);
and UO_6 (O_6,N_49948,N_49854);
nand UO_7 (O_7,N_49811,N_49802);
nor UO_8 (O_8,N_49960,N_49973);
nand UO_9 (O_9,N_49912,N_49836);
nand UO_10 (O_10,N_49991,N_49805);
nor UO_11 (O_11,N_49823,N_49829);
nor UO_12 (O_12,N_49903,N_49900);
nor UO_13 (O_13,N_49902,N_49750);
or UO_14 (O_14,N_49799,N_49883);
nand UO_15 (O_15,N_49881,N_49916);
xor UO_16 (O_16,N_49972,N_49822);
or UO_17 (O_17,N_49957,N_49807);
and UO_18 (O_18,N_49982,N_49803);
nand UO_19 (O_19,N_49832,N_49780);
nand UO_20 (O_20,N_49966,N_49756);
xnor UO_21 (O_21,N_49838,N_49824);
nand UO_22 (O_22,N_49758,N_49941);
and UO_23 (O_23,N_49840,N_49892);
or UO_24 (O_24,N_49926,N_49869);
nand UO_25 (O_25,N_49946,N_49971);
xnor UO_26 (O_26,N_49965,N_49884);
xnor UO_27 (O_27,N_49800,N_49889);
xnor UO_28 (O_28,N_49797,N_49874);
nor UO_29 (O_29,N_49981,N_49952);
and UO_30 (O_30,N_49766,N_49761);
and UO_31 (O_31,N_49939,N_49927);
xnor UO_32 (O_32,N_49950,N_49815);
nand UO_33 (O_33,N_49974,N_49977);
or UO_34 (O_34,N_49928,N_49901);
or UO_35 (O_35,N_49924,N_49954);
and UO_36 (O_36,N_49915,N_49938);
nand UO_37 (O_37,N_49909,N_49969);
nand UO_38 (O_38,N_49845,N_49868);
or UO_39 (O_39,N_49936,N_49996);
xnor UO_40 (O_40,N_49760,N_49904);
nor UO_41 (O_41,N_49784,N_49762);
and UO_42 (O_42,N_49994,N_49751);
nor UO_43 (O_43,N_49988,N_49967);
nand UO_44 (O_44,N_49828,N_49793);
nor UO_45 (O_45,N_49817,N_49961);
xor UO_46 (O_46,N_49871,N_49765);
and UO_47 (O_47,N_49825,N_49764);
nor UO_48 (O_48,N_49935,N_49872);
and UO_49 (O_49,N_49975,N_49873);
or UO_50 (O_50,N_49856,N_49899);
or UO_51 (O_51,N_49922,N_49771);
xor UO_52 (O_52,N_49920,N_49867);
or UO_53 (O_53,N_49942,N_49925);
nor UO_54 (O_54,N_49993,N_49933);
and UO_55 (O_55,N_49808,N_49979);
nor UO_56 (O_56,N_49830,N_49890);
nand UO_57 (O_57,N_49783,N_49932);
xnor UO_58 (O_58,N_49949,N_49853);
nor UO_59 (O_59,N_49806,N_49877);
nand UO_60 (O_60,N_49882,N_49918);
and UO_61 (O_61,N_49880,N_49908);
nand UO_62 (O_62,N_49992,N_49951);
nor UO_63 (O_63,N_49958,N_49847);
xnor UO_64 (O_64,N_49898,N_49755);
nor UO_65 (O_65,N_49879,N_49887);
nor UO_66 (O_66,N_49837,N_49970);
nand UO_67 (O_67,N_49917,N_49792);
nor UO_68 (O_68,N_49919,N_49911);
or UO_69 (O_69,N_49849,N_49987);
or UO_70 (O_70,N_49934,N_49767);
nand UO_71 (O_71,N_49997,N_49763);
or UO_72 (O_72,N_49774,N_49820);
nor UO_73 (O_73,N_49953,N_49779);
nor UO_74 (O_74,N_49857,N_49864);
nor UO_75 (O_75,N_49947,N_49843);
nand UO_76 (O_76,N_49851,N_49754);
nor UO_77 (O_77,N_49778,N_49798);
xnor UO_78 (O_78,N_49852,N_49955);
or UO_79 (O_79,N_49907,N_49968);
nand UO_80 (O_80,N_49846,N_49962);
and UO_81 (O_81,N_49844,N_49931);
nor UO_82 (O_82,N_49895,N_49804);
or UO_83 (O_83,N_49809,N_49818);
and UO_84 (O_84,N_49768,N_49786);
nand UO_85 (O_85,N_49810,N_49773);
nand UO_86 (O_86,N_49886,N_49980);
xnor UO_87 (O_87,N_49921,N_49855);
xor UO_88 (O_88,N_49861,N_49801);
and UO_89 (O_89,N_49929,N_49776);
and UO_90 (O_90,N_49772,N_49891);
nand UO_91 (O_91,N_49983,N_49860);
and UO_92 (O_92,N_49943,N_49876);
xnor UO_93 (O_93,N_49775,N_49976);
nand UO_94 (O_94,N_49888,N_49833);
or UO_95 (O_95,N_49753,N_49827);
nand UO_96 (O_96,N_49781,N_49905);
and UO_97 (O_97,N_49910,N_49757);
nand UO_98 (O_98,N_49893,N_49885);
and UO_99 (O_99,N_49782,N_49896);
and UO_100 (O_100,N_49821,N_49759);
nand UO_101 (O_101,N_49945,N_49897);
nand UO_102 (O_102,N_49995,N_49998);
and UO_103 (O_103,N_49986,N_49870);
or UO_104 (O_104,N_49839,N_49858);
nand UO_105 (O_105,N_49865,N_49866);
nor UO_106 (O_106,N_49862,N_49959);
nand UO_107 (O_107,N_49777,N_49944);
and UO_108 (O_108,N_49791,N_49978);
nor UO_109 (O_109,N_49999,N_49770);
nand UO_110 (O_110,N_49814,N_49906);
or UO_111 (O_111,N_49863,N_49984);
or UO_112 (O_112,N_49816,N_49850);
nand UO_113 (O_113,N_49859,N_49963);
or UO_114 (O_114,N_49875,N_49835);
xor UO_115 (O_115,N_49826,N_49990);
or UO_116 (O_116,N_49831,N_49842);
xnor UO_117 (O_117,N_49930,N_49937);
or UO_118 (O_118,N_49812,N_49795);
nand UO_119 (O_119,N_49913,N_49878);
or UO_120 (O_120,N_49989,N_49964);
or UO_121 (O_121,N_49788,N_49848);
xnor UO_122 (O_122,N_49796,N_49785);
or UO_123 (O_123,N_49914,N_49985);
xor UO_124 (O_124,N_49794,N_49834);
nor UO_125 (O_125,N_49947,N_49973);
nor UO_126 (O_126,N_49789,N_49969);
and UO_127 (O_127,N_49996,N_49853);
nor UO_128 (O_128,N_49972,N_49788);
and UO_129 (O_129,N_49800,N_49988);
or UO_130 (O_130,N_49861,N_49977);
or UO_131 (O_131,N_49905,N_49857);
nand UO_132 (O_132,N_49775,N_49888);
and UO_133 (O_133,N_49842,N_49893);
nor UO_134 (O_134,N_49773,N_49916);
nand UO_135 (O_135,N_49798,N_49866);
and UO_136 (O_136,N_49869,N_49829);
xnor UO_137 (O_137,N_49887,N_49813);
and UO_138 (O_138,N_49763,N_49897);
nor UO_139 (O_139,N_49991,N_49940);
and UO_140 (O_140,N_49839,N_49872);
nand UO_141 (O_141,N_49990,N_49831);
nand UO_142 (O_142,N_49822,N_49863);
and UO_143 (O_143,N_49950,N_49868);
and UO_144 (O_144,N_49883,N_49841);
nand UO_145 (O_145,N_49885,N_49949);
and UO_146 (O_146,N_49810,N_49850);
or UO_147 (O_147,N_49991,N_49771);
or UO_148 (O_148,N_49898,N_49768);
nor UO_149 (O_149,N_49810,N_49781);
nor UO_150 (O_150,N_49752,N_49986);
or UO_151 (O_151,N_49926,N_49992);
and UO_152 (O_152,N_49975,N_49904);
nor UO_153 (O_153,N_49899,N_49832);
xor UO_154 (O_154,N_49927,N_49921);
nand UO_155 (O_155,N_49763,N_49868);
nand UO_156 (O_156,N_49948,N_49974);
and UO_157 (O_157,N_49869,N_49958);
nand UO_158 (O_158,N_49794,N_49870);
nor UO_159 (O_159,N_49926,N_49840);
nor UO_160 (O_160,N_49955,N_49831);
or UO_161 (O_161,N_49826,N_49977);
or UO_162 (O_162,N_49807,N_49786);
nand UO_163 (O_163,N_49913,N_49811);
or UO_164 (O_164,N_49871,N_49976);
nor UO_165 (O_165,N_49797,N_49784);
xnor UO_166 (O_166,N_49772,N_49877);
xor UO_167 (O_167,N_49922,N_49853);
nor UO_168 (O_168,N_49788,N_49892);
or UO_169 (O_169,N_49792,N_49784);
or UO_170 (O_170,N_49956,N_49918);
xor UO_171 (O_171,N_49941,N_49936);
nand UO_172 (O_172,N_49921,N_49933);
nand UO_173 (O_173,N_49907,N_49862);
and UO_174 (O_174,N_49936,N_49947);
xnor UO_175 (O_175,N_49807,N_49776);
xor UO_176 (O_176,N_49938,N_49992);
nand UO_177 (O_177,N_49792,N_49956);
xnor UO_178 (O_178,N_49985,N_49953);
xor UO_179 (O_179,N_49951,N_49918);
or UO_180 (O_180,N_49976,N_49776);
xor UO_181 (O_181,N_49970,N_49922);
nor UO_182 (O_182,N_49827,N_49760);
and UO_183 (O_183,N_49757,N_49775);
xnor UO_184 (O_184,N_49766,N_49901);
nand UO_185 (O_185,N_49772,N_49956);
nand UO_186 (O_186,N_49922,N_49787);
nand UO_187 (O_187,N_49844,N_49800);
xnor UO_188 (O_188,N_49998,N_49938);
xnor UO_189 (O_189,N_49752,N_49878);
and UO_190 (O_190,N_49763,N_49860);
nand UO_191 (O_191,N_49854,N_49995);
or UO_192 (O_192,N_49773,N_49844);
or UO_193 (O_193,N_49990,N_49787);
nand UO_194 (O_194,N_49879,N_49906);
nand UO_195 (O_195,N_49884,N_49785);
or UO_196 (O_196,N_49819,N_49955);
nand UO_197 (O_197,N_49886,N_49819);
nand UO_198 (O_198,N_49994,N_49874);
xnor UO_199 (O_199,N_49933,N_49820);
and UO_200 (O_200,N_49896,N_49825);
xor UO_201 (O_201,N_49968,N_49986);
xnor UO_202 (O_202,N_49949,N_49805);
xnor UO_203 (O_203,N_49809,N_49856);
xor UO_204 (O_204,N_49998,N_49965);
or UO_205 (O_205,N_49986,N_49874);
or UO_206 (O_206,N_49836,N_49782);
and UO_207 (O_207,N_49826,N_49994);
xor UO_208 (O_208,N_49956,N_49830);
nand UO_209 (O_209,N_49797,N_49860);
xnor UO_210 (O_210,N_49806,N_49949);
and UO_211 (O_211,N_49923,N_49946);
nor UO_212 (O_212,N_49789,N_49914);
nand UO_213 (O_213,N_49772,N_49788);
xnor UO_214 (O_214,N_49815,N_49762);
nand UO_215 (O_215,N_49804,N_49827);
nor UO_216 (O_216,N_49799,N_49792);
xnor UO_217 (O_217,N_49955,N_49902);
nor UO_218 (O_218,N_49902,N_49808);
and UO_219 (O_219,N_49868,N_49758);
nor UO_220 (O_220,N_49781,N_49862);
or UO_221 (O_221,N_49810,N_49807);
nor UO_222 (O_222,N_49862,N_49916);
or UO_223 (O_223,N_49781,N_49966);
nor UO_224 (O_224,N_49790,N_49978);
or UO_225 (O_225,N_49814,N_49862);
nand UO_226 (O_226,N_49792,N_49822);
nor UO_227 (O_227,N_49786,N_49908);
or UO_228 (O_228,N_49808,N_49939);
nand UO_229 (O_229,N_49954,N_49856);
nor UO_230 (O_230,N_49966,N_49903);
nand UO_231 (O_231,N_49791,N_49830);
nor UO_232 (O_232,N_49825,N_49993);
and UO_233 (O_233,N_49809,N_49936);
nand UO_234 (O_234,N_49810,N_49906);
xnor UO_235 (O_235,N_49909,N_49937);
xor UO_236 (O_236,N_49879,N_49876);
and UO_237 (O_237,N_49909,N_49809);
and UO_238 (O_238,N_49890,N_49918);
and UO_239 (O_239,N_49989,N_49969);
nor UO_240 (O_240,N_49877,N_49892);
nor UO_241 (O_241,N_49972,N_49821);
and UO_242 (O_242,N_49822,N_49825);
nor UO_243 (O_243,N_49843,N_49902);
xnor UO_244 (O_244,N_49820,N_49981);
xor UO_245 (O_245,N_49846,N_49935);
and UO_246 (O_246,N_49925,N_49816);
nand UO_247 (O_247,N_49820,N_49984);
xnor UO_248 (O_248,N_49922,N_49858);
xor UO_249 (O_249,N_49982,N_49836);
nor UO_250 (O_250,N_49792,N_49805);
or UO_251 (O_251,N_49869,N_49761);
or UO_252 (O_252,N_49787,N_49993);
xor UO_253 (O_253,N_49791,N_49897);
or UO_254 (O_254,N_49823,N_49857);
nand UO_255 (O_255,N_49767,N_49883);
and UO_256 (O_256,N_49823,N_49938);
and UO_257 (O_257,N_49848,N_49865);
and UO_258 (O_258,N_49920,N_49768);
and UO_259 (O_259,N_49864,N_49787);
nand UO_260 (O_260,N_49797,N_49782);
nor UO_261 (O_261,N_49776,N_49882);
nor UO_262 (O_262,N_49923,N_49789);
and UO_263 (O_263,N_49947,N_49872);
and UO_264 (O_264,N_49840,N_49800);
xnor UO_265 (O_265,N_49992,N_49865);
xnor UO_266 (O_266,N_49755,N_49815);
nand UO_267 (O_267,N_49916,N_49844);
and UO_268 (O_268,N_49813,N_49979);
nor UO_269 (O_269,N_49947,N_49959);
or UO_270 (O_270,N_49775,N_49793);
or UO_271 (O_271,N_49940,N_49831);
or UO_272 (O_272,N_49830,N_49932);
and UO_273 (O_273,N_49771,N_49957);
or UO_274 (O_274,N_49842,N_49815);
nand UO_275 (O_275,N_49905,N_49814);
nor UO_276 (O_276,N_49873,N_49887);
or UO_277 (O_277,N_49814,N_49858);
xor UO_278 (O_278,N_49888,N_49875);
and UO_279 (O_279,N_49958,N_49929);
and UO_280 (O_280,N_49788,N_49939);
xnor UO_281 (O_281,N_49972,N_49855);
nor UO_282 (O_282,N_49921,N_49760);
nor UO_283 (O_283,N_49824,N_49841);
nor UO_284 (O_284,N_49938,N_49939);
nand UO_285 (O_285,N_49858,N_49892);
xor UO_286 (O_286,N_49791,N_49823);
nand UO_287 (O_287,N_49860,N_49901);
nor UO_288 (O_288,N_49848,N_49771);
or UO_289 (O_289,N_49767,N_49901);
nor UO_290 (O_290,N_49928,N_49985);
nand UO_291 (O_291,N_49899,N_49850);
nor UO_292 (O_292,N_49913,N_49843);
and UO_293 (O_293,N_49869,N_49965);
xor UO_294 (O_294,N_49843,N_49849);
xor UO_295 (O_295,N_49945,N_49805);
xnor UO_296 (O_296,N_49954,N_49846);
nor UO_297 (O_297,N_49904,N_49884);
nor UO_298 (O_298,N_49791,N_49892);
or UO_299 (O_299,N_49921,N_49883);
xnor UO_300 (O_300,N_49973,N_49752);
nor UO_301 (O_301,N_49937,N_49772);
nand UO_302 (O_302,N_49877,N_49968);
and UO_303 (O_303,N_49936,N_49852);
nor UO_304 (O_304,N_49760,N_49967);
xnor UO_305 (O_305,N_49984,N_49845);
nor UO_306 (O_306,N_49844,N_49954);
and UO_307 (O_307,N_49868,N_49880);
nor UO_308 (O_308,N_49787,N_49969);
nor UO_309 (O_309,N_49855,N_49893);
or UO_310 (O_310,N_49862,N_49825);
nor UO_311 (O_311,N_49925,N_49886);
and UO_312 (O_312,N_49860,N_49770);
nor UO_313 (O_313,N_49765,N_49976);
xor UO_314 (O_314,N_49794,N_49999);
and UO_315 (O_315,N_49859,N_49836);
nand UO_316 (O_316,N_49980,N_49976);
nor UO_317 (O_317,N_49815,N_49753);
and UO_318 (O_318,N_49973,N_49842);
nor UO_319 (O_319,N_49876,N_49763);
nand UO_320 (O_320,N_49904,N_49979);
and UO_321 (O_321,N_49947,N_49859);
and UO_322 (O_322,N_49824,N_49787);
xor UO_323 (O_323,N_49985,N_49825);
nor UO_324 (O_324,N_49957,N_49936);
and UO_325 (O_325,N_49849,N_49900);
xnor UO_326 (O_326,N_49828,N_49849);
xor UO_327 (O_327,N_49785,N_49819);
nand UO_328 (O_328,N_49941,N_49803);
or UO_329 (O_329,N_49870,N_49964);
or UO_330 (O_330,N_49884,N_49821);
or UO_331 (O_331,N_49940,N_49926);
nor UO_332 (O_332,N_49894,N_49810);
or UO_333 (O_333,N_49988,N_49759);
nor UO_334 (O_334,N_49891,N_49931);
xnor UO_335 (O_335,N_49857,N_49942);
xnor UO_336 (O_336,N_49788,N_49812);
nor UO_337 (O_337,N_49950,N_49982);
and UO_338 (O_338,N_49912,N_49919);
nor UO_339 (O_339,N_49964,N_49955);
or UO_340 (O_340,N_49973,N_49995);
nor UO_341 (O_341,N_49756,N_49947);
xnor UO_342 (O_342,N_49870,N_49868);
nand UO_343 (O_343,N_49983,N_49859);
or UO_344 (O_344,N_49969,N_49941);
and UO_345 (O_345,N_49811,N_49862);
xnor UO_346 (O_346,N_49792,N_49760);
or UO_347 (O_347,N_49859,N_49924);
xor UO_348 (O_348,N_49847,N_49981);
and UO_349 (O_349,N_49998,N_49755);
xor UO_350 (O_350,N_49818,N_49823);
xor UO_351 (O_351,N_49854,N_49981);
nor UO_352 (O_352,N_49928,N_49887);
and UO_353 (O_353,N_49937,N_49788);
xnor UO_354 (O_354,N_49899,N_49961);
nor UO_355 (O_355,N_49993,N_49828);
or UO_356 (O_356,N_49959,N_49816);
nor UO_357 (O_357,N_49807,N_49859);
nand UO_358 (O_358,N_49826,N_49974);
nand UO_359 (O_359,N_49790,N_49993);
and UO_360 (O_360,N_49770,N_49871);
and UO_361 (O_361,N_49907,N_49999);
nor UO_362 (O_362,N_49851,N_49855);
nor UO_363 (O_363,N_49926,N_49881);
and UO_364 (O_364,N_49880,N_49752);
nand UO_365 (O_365,N_49752,N_49857);
nand UO_366 (O_366,N_49870,N_49750);
nor UO_367 (O_367,N_49830,N_49785);
nor UO_368 (O_368,N_49851,N_49959);
nand UO_369 (O_369,N_49839,N_49848);
and UO_370 (O_370,N_49828,N_49870);
nor UO_371 (O_371,N_49787,N_49895);
xor UO_372 (O_372,N_49860,N_49784);
or UO_373 (O_373,N_49876,N_49812);
and UO_374 (O_374,N_49793,N_49779);
or UO_375 (O_375,N_49843,N_49762);
nor UO_376 (O_376,N_49822,N_49836);
and UO_377 (O_377,N_49930,N_49841);
nand UO_378 (O_378,N_49929,N_49963);
nand UO_379 (O_379,N_49826,N_49971);
nor UO_380 (O_380,N_49975,N_49760);
nand UO_381 (O_381,N_49854,N_49775);
and UO_382 (O_382,N_49833,N_49831);
xor UO_383 (O_383,N_49822,N_49880);
xor UO_384 (O_384,N_49759,N_49969);
and UO_385 (O_385,N_49773,N_49976);
nor UO_386 (O_386,N_49921,N_49953);
nand UO_387 (O_387,N_49985,N_49870);
nor UO_388 (O_388,N_49858,N_49983);
xnor UO_389 (O_389,N_49800,N_49986);
nand UO_390 (O_390,N_49777,N_49799);
and UO_391 (O_391,N_49827,N_49809);
xnor UO_392 (O_392,N_49818,N_49893);
or UO_393 (O_393,N_49980,N_49772);
nor UO_394 (O_394,N_49825,N_49805);
xnor UO_395 (O_395,N_49797,N_49781);
nand UO_396 (O_396,N_49949,N_49765);
xor UO_397 (O_397,N_49879,N_49932);
nand UO_398 (O_398,N_49778,N_49879);
xnor UO_399 (O_399,N_49797,N_49792);
xor UO_400 (O_400,N_49765,N_49807);
and UO_401 (O_401,N_49755,N_49840);
and UO_402 (O_402,N_49895,N_49835);
or UO_403 (O_403,N_49769,N_49933);
nor UO_404 (O_404,N_49818,N_49820);
nor UO_405 (O_405,N_49933,N_49997);
nor UO_406 (O_406,N_49940,N_49754);
xnor UO_407 (O_407,N_49881,N_49826);
xor UO_408 (O_408,N_49899,N_49922);
or UO_409 (O_409,N_49928,N_49925);
or UO_410 (O_410,N_49883,N_49914);
or UO_411 (O_411,N_49799,N_49915);
nor UO_412 (O_412,N_49888,N_49900);
or UO_413 (O_413,N_49921,N_49852);
or UO_414 (O_414,N_49781,N_49990);
nor UO_415 (O_415,N_49990,N_49983);
or UO_416 (O_416,N_49863,N_49820);
xor UO_417 (O_417,N_49915,N_49969);
xnor UO_418 (O_418,N_49967,N_49901);
nand UO_419 (O_419,N_49978,N_49904);
nor UO_420 (O_420,N_49765,N_49831);
and UO_421 (O_421,N_49841,N_49863);
and UO_422 (O_422,N_49852,N_49762);
nand UO_423 (O_423,N_49990,N_49961);
xor UO_424 (O_424,N_49990,N_49922);
nand UO_425 (O_425,N_49996,N_49926);
and UO_426 (O_426,N_49789,N_49998);
or UO_427 (O_427,N_49942,N_49802);
nand UO_428 (O_428,N_49767,N_49787);
nor UO_429 (O_429,N_49996,N_49890);
xor UO_430 (O_430,N_49880,N_49826);
nand UO_431 (O_431,N_49951,N_49835);
or UO_432 (O_432,N_49887,N_49910);
or UO_433 (O_433,N_49860,N_49918);
nand UO_434 (O_434,N_49823,N_49943);
and UO_435 (O_435,N_49751,N_49944);
xor UO_436 (O_436,N_49866,N_49999);
and UO_437 (O_437,N_49917,N_49758);
nor UO_438 (O_438,N_49849,N_49989);
or UO_439 (O_439,N_49830,N_49797);
nor UO_440 (O_440,N_49982,N_49789);
nor UO_441 (O_441,N_49833,N_49824);
nand UO_442 (O_442,N_49937,N_49942);
or UO_443 (O_443,N_49760,N_49891);
or UO_444 (O_444,N_49890,N_49813);
nand UO_445 (O_445,N_49952,N_49811);
xnor UO_446 (O_446,N_49998,N_49852);
and UO_447 (O_447,N_49786,N_49800);
nand UO_448 (O_448,N_49939,N_49891);
nor UO_449 (O_449,N_49776,N_49846);
nand UO_450 (O_450,N_49783,N_49863);
nor UO_451 (O_451,N_49950,N_49988);
and UO_452 (O_452,N_49940,N_49828);
and UO_453 (O_453,N_49815,N_49867);
xor UO_454 (O_454,N_49892,N_49940);
nand UO_455 (O_455,N_49820,N_49993);
nand UO_456 (O_456,N_49962,N_49783);
xnor UO_457 (O_457,N_49777,N_49997);
xor UO_458 (O_458,N_49773,N_49786);
nor UO_459 (O_459,N_49925,N_49835);
and UO_460 (O_460,N_49815,N_49883);
nand UO_461 (O_461,N_49940,N_49968);
nor UO_462 (O_462,N_49805,N_49767);
nand UO_463 (O_463,N_49960,N_49763);
nor UO_464 (O_464,N_49755,N_49951);
and UO_465 (O_465,N_49790,N_49965);
and UO_466 (O_466,N_49750,N_49855);
and UO_467 (O_467,N_49854,N_49927);
xor UO_468 (O_468,N_49794,N_49914);
and UO_469 (O_469,N_49956,N_49897);
or UO_470 (O_470,N_49833,N_49756);
or UO_471 (O_471,N_49763,N_49783);
xnor UO_472 (O_472,N_49962,N_49768);
and UO_473 (O_473,N_49844,N_49979);
nor UO_474 (O_474,N_49850,N_49844);
xor UO_475 (O_475,N_49760,N_49813);
or UO_476 (O_476,N_49858,N_49764);
xnor UO_477 (O_477,N_49766,N_49854);
or UO_478 (O_478,N_49869,N_49794);
and UO_479 (O_479,N_49933,N_49824);
nand UO_480 (O_480,N_49851,N_49876);
nand UO_481 (O_481,N_49843,N_49929);
nand UO_482 (O_482,N_49899,N_49847);
and UO_483 (O_483,N_49926,N_49993);
nor UO_484 (O_484,N_49828,N_49999);
xor UO_485 (O_485,N_49977,N_49840);
or UO_486 (O_486,N_49855,N_49946);
or UO_487 (O_487,N_49900,N_49980);
nor UO_488 (O_488,N_49894,N_49787);
xnor UO_489 (O_489,N_49758,N_49831);
nor UO_490 (O_490,N_49814,N_49925);
nor UO_491 (O_491,N_49968,N_49917);
or UO_492 (O_492,N_49897,N_49835);
nand UO_493 (O_493,N_49773,N_49769);
and UO_494 (O_494,N_49851,N_49784);
or UO_495 (O_495,N_49888,N_49799);
xnor UO_496 (O_496,N_49824,N_49893);
or UO_497 (O_497,N_49751,N_49926);
nor UO_498 (O_498,N_49865,N_49855);
or UO_499 (O_499,N_49760,N_49899);
nor UO_500 (O_500,N_49805,N_49765);
and UO_501 (O_501,N_49851,N_49770);
and UO_502 (O_502,N_49771,N_49994);
and UO_503 (O_503,N_49810,N_49794);
and UO_504 (O_504,N_49800,N_49985);
nand UO_505 (O_505,N_49956,N_49965);
xor UO_506 (O_506,N_49807,N_49803);
and UO_507 (O_507,N_49996,N_49882);
and UO_508 (O_508,N_49927,N_49863);
nand UO_509 (O_509,N_49915,N_49772);
or UO_510 (O_510,N_49939,N_49772);
nand UO_511 (O_511,N_49972,N_49852);
or UO_512 (O_512,N_49977,N_49893);
xor UO_513 (O_513,N_49962,N_49872);
nor UO_514 (O_514,N_49933,N_49849);
nand UO_515 (O_515,N_49872,N_49964);
nand UO_516 (O_516,N_49891,N_49761);
xnor UO_517 (O_517,N_49847,N_49890);
nand UO_518 (O_518,N_49956,N_49952);
nand UO_519 (O_519,N_49867,N_49964);
nand UO_520 (O_520,N_49804,N_49866);
nand UO_521 (O_521,N_49980,N_49791);
xor UO_522 (O_522,N_49982,N_49988);
nor UO_523 (O_523,N_49849,N_49816);
nor UO_524 (O_524,N_49998,N_49834);
and UO_525 (O_525,N_49903,N_49975);
xnor UO_526 (O_526,N_49997,N_49882);
nand UO_527 (O_527,N_49907,N_49960);
nor UO_528 (O_528,N_49753,N_49774);
or UO_529 (O_529,N_49912,N_49808);
nor UO_530 (O_530,N_49997,N_49833);
or UO_531 (O_531,N_49945,N_49914);
and UO_532 (O_532,N_49885,N_49986);
nor UO_533 (O_533,N_49842,N_49993);
xor UO_534 (O_534,N_49989,N_49832);
and UO_535 (O_535,N_49971,N_49885);
or UO_536 (O_536,N_49785,N_49966);
and UO_537 (O_537,N_49981,N_49940);
nor UO_538 (O_538,N_49941,N_49821);
xnor UO_539 (O_539,N_49797,N_49916);
or UO_540 (O_540,N_49891,N_49794);
nor UO_541 (O_541,N_49780,N_49916);
xnor UO_542 (O_542,N_49846,N_49952);
xnor UO_543 (O_543,N_49840,N_49887);
and UO_544 (O_544,N_49896,N_49817);
and UO_545 (O_545,N_49959,N_49871);
nor UO_546 (O_546,N_49777,N_49994);
xnor UO_547 (O_547,N_49918,N_49957);
nor UO_548 (O_548,N_49885,N_49770);
xnor UO_549 (O_549,N_49779,N_49835);
nand UO_550 (O_550,N_49795,N_49833);
or UO_551 (O_551,N_49920,N_49762);
nor UO_552 (O_552,N_49918,N_49841);
nand UO_553 (O_553,N_49806,N_49923);
nand UO_554 (O_554,N_49916,N_49838);
nand UO_555 (O_555,N_49800,N_49966);
nor UO_556 (O_556,N_49816,N_49765);
xor UO_557 (O_557,N_49875,N_49783);
nand UO_558 (O_558,N_49844,N_49867);
nor UO_559 (O_559,N_49792,N_49775);
xnor UO_560 (O_560,N_49912,N_49766);
or UO_561 (O_561,N_49871,N_49779);
and UO_562 (O_562,N_49834,N_49942);
or UO_563 (O_563,N_49919,N_49986);
nor UO_564 (O_564,N_49896,N_49958);
nand UO_565 (O_565,N_49937,N_49837);
or UO_566 (O_566,N_49825,N_49997);
and UO_567 (O_567,N_49776,N_49754);
or UO_568 (O_568,N_49775,N_49986);
and UO_569 (O_569,N_49897,N_49901);
nand UO_570 (O_570,N_49931,N_49760);
nor UO_571 (O_571,N_49763,N_49918);
xor UO_572 (O_572,N_49863,N_49852);
or UO_573 (O_573,N_49787,N_49913);
and UO_574 (O_574,N_49927,N_49963);
and UO_575 (O_575,N_49757,N_49873);
xnor UO_576 (O_576,N_49756,N_49840);
or UO_577 (O_577,N_49873,N_49936);
nand UO_578 (O_578,N_49792,N_49815);
nor UO_579 (O_579,N_49883,N_49998);
nor UO_580 (O_580,N_49854,N_49840);
nand UO_581 (O_581,N_49937,N_49985);
nand UO_582 (O_582,N_49885,N_49839);
nor UO_583 (O_583,N_49864,N_49756);
nand UO_584 (O_584,N_49979,N_49925);
nand UO_585 (O_585,N_49771,N_49797);
nor UO_586 (O_586,N_49940,N_49794);
and UO_587 (O_587,N_49862,N_49775);
nor UO_588 (O_588,N_49785,N_49835);
and UO_589 (O_589,N_49876,N_49819);
nor UO_590 (O_590,N_49826,N_49916);
and UO_591 (O_591,N_49869,N_49830);
xor UO_592 (O_592,N_49903,N_49909);
xnor UO_593 (O_593,N_49910,N_49940);
and UO_594 (O_594,N_49973,N_49869);
or UO_595 (O_595,N_49799,N_49856);
xnor UO_596 (O_596,N_49969,N_49872);
xor UO_597 (O_597,N_49775,N_49798);
nand UO_598 (O_598,N_49763,N_49778);
nand UO_599 (O_599,N_49918,N_49921);
or UO_600 (O_600,N_49917,N_49862);
nand UO_601 (O_601,N_49774,N_49945);
nor UO_602 (O_602,N_49773,N_49929);
nor UO_603 (O_603,N_49909,N_49858);
nor UO_604 (O_604,N_49852,N_49785);
nor UO_605 (O_605,N_49750,N_49769);
nor UO_606 (O_606,N_49761,N_49790);
and UO_607 (O_607,N_49757,N_49752);
and UO_608 (O_608,N_49752,N_49994);
and UO_609 (O_609,N_49957,N_49853);
xor UO_610 (O_610,N_49816,N_49899);
nor UO_611 (O_611,N_49800,N_49813);
or UO_612 (O_612,N_49921,N_49884);
or UO_613 (O_613,N_49977,N_49926);
nor UO_614 (O_614,N_49986,N_49790);
and UO_615 (O_615,N_49956,N_49798);
xor UO_616 (O_616,N_49943,N_49991);
nand UO_617 (O_617,N_49784,N_49786);
or UO_618 (O_618,N_49886,N_49875);
and UO_619 (O_619,N_49939,N_49865);
and UO_620 (O_620,N_49908,N_49981);
or UO_621 (O_621,N_49880,N_49893);
nand UO_622 (O_622,N_49905,N_49791);
and UO_623 (O_623,N_49807,N_49844);
or UO_624 (O_624,N_49901,N_49788);
or UO_625 (O_625,N_49850,N_49991);
xor UO_626 (O_626,N_49815,N_49870);
nor UO_627 (O_627,N_49885,N_49902);
xnor UO_628 (O_628,N_49951,N_49782);
and UO_629 (O_629,N_49842,N_49866);
nor UO_630 (O_630,N_49878,N_49945);
or UO_631 (O_631,N_49759,N_49842);
xor UO_632 (O_632,N_49993,N_49862);
xor UO_633 (O_633,N_49945,N_49824);
xor UO_634 (O_634,N_49887,N_49848);
nor UO_635 (O_635,N_49810,N_49840);
nor UO_636 (O_636,N_49942,N_49894);
nand UO_637 (O_637,N_49917,N_49796);
or UO_638 (O_638,N_49788,N_49883);
nor UO_639 (O_639,N_49877,N_49767);
nor UO_640 (O_640,N_49761,N_49960);
nand UO_641 (O_641,N_49780,N_49790);
nand UO_642 (O_642,N_49959,N_49771);
xor UO_643 (O_643,N_49829,N_49954);
nor UO_644 (O_644,N_49917,N_49993);
nor UO_645 (O_645,N_49951,N_49849);
xor UO_646 (O_646,N_49887,N_49945);
xnor UO_647 (O_647,N_49867,N_49898);
and UO_648 (O_648,N_49984,N_49843);
nand UO_649 (O_649,N_49996,N_49886);
xor UO_650 (O_650,N_49938,N_49842);
and UO_651 (O_651,N_49839,N_49788);
or UO_652 (O_652,N_49768,N_49760);
nor UO_653 (O_653,N_49868,N_49888);
nand UO_654 (O_654,N_49840,N_49846);
nor UO_655 (O_655,N_49848,N_49905);
or UO_656 (O_656,N_49986,N_49778);
nor UO_657 (O_657,N_49862,N_49882);
nor UO_658 (O_658,N_49966,N_49768);
nand UO_659 (O_659,N_49760,N_49856);
or UO_660 (O_660,N_49874,N_49759);
xnor UO_661 (O_661,N_49944,N_49871);
and UO_662 (O_662,N_49812,N_49983);
and UO_663 (O_663,N_49822,N_49831);
or UO_664 (O_664,N_49933,N_49904);
and UO_665 (O_665,N_49908,N_49797);
and UO_666 (O_666,N_49937,N_49851);
or UO_667 (O_667,N_49876,N_49779);
or UO_668 (O_668,N_49787,N_49919);
and UO_669 (O_669,N_49911,N_49860);
and UO_670 (O_670,N_49890,N_49801);
or UO_671 (O_671,N_49914,N_49983);
and UO_672 (O_672,N_49983,N_49806);
xor UO_673 (O_673,N_49785,N_49857);
or UO_674 (O_674,N_49981,N_49776);
nand UO_675 (O_675,N_49916,N_49891);
nand UO_676 (O_676,N_49956,N_49983);
or UO_677 (O_677,N_49959,N_49886);
nand UO_678 (O_678,N_49863,N_49794);
or UO_679 (O_679,N_49938,N_49901);
nor UO_680 (O_680,N_49934,N_49978);
nor UO_681 (O_681,N_49810,N_49784);
xor UO_682 (O_682,N_49890,N_49904);
xnor UO_683 (O_683,N_49956,N_49888);
xor UO_684 (O_684,N_49817,N_49800);
or UO_685 (O_685,N_49902,N_49827);
nor UO_686 (O_686,N_49847,N_49986);
nand UO_687 (O_687,N_49818,N_49875);
xor UO_688 (O_688,N_49892,N_49860);
and UO_689 (O_689,N_49853,N_49806);
xnor UO_690 (O_690,N_49960,N_49924);
and UO_691 (O_691,N_49793,N_49950);
nand UO_692 (O_692,N_49949,N_49903);
xor UO_693 (O_693,N_49836,N_49803);
xor UO_694 (O_694,N_49807,N_49797);
or UO_695 (O_695,N_49887,N_49769);
or UO_696 (O_696,N_49972,N_49790);
and UO_697 (O_697,N_49859,N_49921);
or UO_698 (O_698,N_49799,N_49919);
nor UO_699 (O_699,N_49949,N_49770);
nor UO_700 (O_700,N_49775,N_49995);
nor UO_701 (O_701,N_49873,N_49775);
xnor UO_702 (O_702,N_49785,N_49909);
and UO_703 (O_703,N_49963,N_49909);
and UO_704 (O_704,N_49981,N_49919);
xor UO_705 (O_705,N_49832,N_49818);
nand UO_706 (O_706,N_49955,N_49863);
nor UO_707 (O_707,N_49926,N_49800);
and UO_708 (O_708,N_49990,N_49938);
or UO_709 (O_709,N_49903,N_49870);
nand UO_710 (O_710,N_49934,N_49877);
xor UO_711 (O_711,N_49966,N_49957);
nor UO_712 (O_712,N_49965,N_49773);
or UO_713 (O_713,N_49983,N_49962);
and UO_714 (O_714,N_49989,N_49937);
and UO_715 (O_715,N_49856,N_49970);
and UO_716 (O_716,N_49811,N_49960);
nor UO_717 (O_717,N_49813,N_49971);
nand UO_718 (O_718,N_49963,N_49845);
or UO_719 (O_719,N_49848,N_49818);
xnor UO_720 (O_720,N_49918,N_49925);
nand UO_721 (O_721,N_49862,N_49766);
and UO_722 (O_722,N_49936,N_49978);
and UO_723 (O_723,N_49966,N_49886);
nor UO_724 (O_724,N_49838,N_49952);
xnor UO_725 (O_725,N_49986,N_49964);
nor UO_726 (O_726,N_49888,N_49860);
and UO_727 (O_727,N_49883,N_49978);
and UO_728 (O_728,N_49767,N_49844);
xnor UO_729 (O_729,N_49773,N_49991);
or UO_730 (O_730,N_49853,N_49890);
xor UO_731 (O_731,N_49774,N_49815);
and UO_732 (O_732,N_49769,N_49994);
xnor UO_733 (O_733,N_49942,N_49788);
xor UO_734 (O_734,N_49943,N_49848);
nor UO_735 (O_735,N_49812,N_49819);
nor UO_736 (O_736,N_49865,N_49938);
nor UO_737 (O_737,N_49791,N_49815);
nand UO_738 (O_738,N_49888,N_49789);
xor UO_739 (O_739,N_49781,N_49842);
nand UO_740 (O_740,N_49848,N_49938);
nand UO_741 (O_741,N_49933,N_49976);
or UO_742 (O_742,N_49778,N_49985);
and UO_743 (O_743,N_49942,N_49813);
or UO_744 (O_744,N_49861,N_49963);
nand UO_745 (O_745,N_49883,N_49819);
and UO_746 (O_746,N_49898,N_49887);
and UO_747 (O_747,N_49813,N_49957);
or UO_748 (O_748,N_49902,N_49797);
and UO_749 (O_749,N_49755,N_49792);
xnor UO_750 (O_750,N_49874,N_49843);
or UO_751 (O_751,N_49995,N_49978);
xor UO_752 (O_752,N_49876,N_49937);
or UO_753 (O_753,N_49823,N_49995);
nor UO_754 (O_754,N_49876,N_49786);
and UO_755 (O_755,N_49829,N_49926);
xor UO_756 (O_756,N_49967,N_49891);
or UO_757 (O_757,N_49847,N_49796);
xor UO_758 (O_758,N_49907,N_49911);
and UO_759 (O_759,N_49833,N_49925);
xor UO_760 (O_760,N_49999,N_49985);
nand UO_761 (O_761,N_49828,N_49883);
xnor UO_762 (O_762,N_49877,N_49793);
and UO_763 (O_763,N_49913,N_49914);
nor UO_764 (O_764,N_49846,N_49927);
and UO_765 (O_765,N_49938,N_49916);
xnor UO_766 (O_766,N_49977,N_49957);
and UO_767 (O_767,N_49836,N_49975);
and UO_768 (O_768,N_49879,N_49850);
nor UO_769 (O_769,N_49849,N_49838);
or UO_770 (O_770,N_49952,N_49807);
nor UO_771 (O_771,N_49988,N_49787);
nand UO_772 (O_772,N_49953,N_49765);
or UO_773 (O_773,N_49941,N_49811);
or UO_774 (O_774,N_49787,N_49852);
or UO_775 (O_775,N_49889,N_49854);
or UO_776 (O_776,N_49839,N_49922);
and UO_777 (O_777,N_49896,N_49867);
nand UO_778 (O_778,N_49823,N_49903);
or UO_779 (O_779,N_49754,N_49858);
or UO_780 (O_780,N_49927,N_49781);
nor UO_781 (O_781,N_49912,N_49778);
and UO_782 (O_782,N_49796,N_49945);
nand UO_783 (O_783,N_49881,N_49984);
and UO_784 (O_784,N_49951,N_49751);
nand UO_785 (O_785,N_49916,N_49989);
nand UO_786 (O_786,N_49767,N_49902);
xor UO_787 (O_787,N_49762,N_49856);
and UO_788 (O_788,N_49860,N_49787);
nand UO_789 (O_789,N_49897,N_49995);
nor UO_790 (O_790,N_49778,N_49916);
and UO_791 (O_791,N_49937,N_49967);
or UO_792 (O_792,N_49899,N_49855);
xnor UO_793 (O_793,N_49758,N_49870);
nor UO_794 (O_794,N_49945,N_49757);
nor UO_795 (O_795,N_49871,N_49918);
or UO_796 (O_796,N_49980,N_49919);
and UO_797 (O_797,N_49827,N_49929);
and UO_798 (O_798,N_49820,N_49911);
and UO_799 (O_799,N_49955,N_49768);
xnor UO_800 (O_800,N_49946,N_49786);
xnor UO_801 (O_801,N_49843,N_49821);
xor UO_802 (O_802,N_49861,N_49969);
and UO_803 (O_803,N_49885,N_49879);
and UO_804 (O_804,N_49817,N_49887);
xor UO_805 (O_805,N_49771,N_49900);
xor UO_806 (O_806,N_49956,N_49872);
and UO_807 (O_807,N_49765,N_49971);
and UO_808 (O_808,N_49850,N_49831);
and UO_809 (O_809,N_49988,N_49996);
or UO_810 (O_810,N_49947,N_49862);
xnor UO_811 (O_811,N_49771,N_49843);
nor UO_812 (O_812,N_49906,N_49872);
xnor UO_813 (O_813,N_49930,N_49795);
or UO_814 (O_814,N_49953,N_49846);
and UO_815 (O_815,N_49973,N_49941);
xor UO_816 (O_816,N_49844,N_49962);
nand UO_817 (O_817,N_49756,N_49801);
or UO_818 (O_818,N_49949,N_49775);
and UO_819 (O_819,N_49998,N_49795);
xor UO_820 (O_820,N_49883,N_49977);
or UO_821 (O_821,N_49928,N_49947);
or UO_822 (O_822,N_49992,N_49874);
xor UO_823 (O_823,N_49765,N_49849);
and UO_824 (O_824,N_49791,N_49887);
or UO_825 (O_825,N_49907,N_49949);
nand UO_826 (O_826,N_49915,N_49810);
nand UO_827 (O_827,N_49861,N_49829);
xnor UO_828 (O_828,N_49817,N_49882);
xnor UO_829 (O_829,N_49808,N_49862);
nor UO_830 (O_830,N_49978,N_49799);
nor UO_831 (O_831,N_49838,N_49778);
xor UO_832 (O_832,N_49889,N_49841);
and UO_833 (O_833,N_49757,N_49843);
nand UO_834 (O_834,N_49925,N_49879);
or UO_835 (O_835,N_49964,N_49916);
and UO_836 (O_836,N_49827,N_49820);
xor UO_837 (O_837,N_49967,N_49991);
nand UO_838 (O_838,N_49783,N_49886);
nand UO_839 (O_839,N_49988,N_49793);
or UO_840 (O_840,N_49897,N_49855);
nor UO_841 (O_841,N_49985,N_49904);
and UO_842 (O_842,N_49795,N_49898);
xor UO_843 (O_843,N_49905,N_49784);
nor UO_844 (O_844,N_49933,N_49788);
or UO_845 (O_845,N_49803,N_49762);
or UO_846 (O_846,N_49855,N_49881);
nor UO_847 (O_847,N_49972,N_49764);
and UO_848 (O_848,N_49789,N_49979);
nor UO_849 (O_849,N_49781,N_49783);
nor UO_850 (O_850,N_49965,N_49963);
or UO_851 (O_851,N_49771,N_49937);
nand UO_852 (O_852,N_49831,N_49755);
xnor UO_853 (O_853,N_49769,N_49957);
and UO_854 (O_854,N_49850,N_49790);
nor UO_855 (O_855,N_49972,N_49933);
or UO_856 (O_856,N_49938,N_49872);
nand UO_857 (O_857,N_49911,N_49905);
nand UO_858 (O_858,N_49761,N_49995);
xnor UO_859 (O_859,N_49949,N_49807);
nor UO_860 (O_860,N_49798,N_49804);
nor UO_861 (O_861,N_49788,N_49894);
nor UO_862 (O_862,N_49848,N_49919);
nor UO_863 (O_863,N_49840,N_49989);
nand UO_864 (O_864,N_49835,N_49820);
and UO_865 (O_865,N_49754,N_49846);
xnor UO_866 (O_866,N_49901,N_49822);
nand UO_867 (O_867,N_49978,N_49800);
and UO_868 (O_868,N_49998,N_49949);
xnor UO_869 (O_869,N_49919,N_49805);
or UO_870 (O_870,N_49877,N_49971);
nor UO_871 (O_871,N_49866,N_49787);
nor UO_872 (O_872,N_49849,N_49937);
nor UO_873 (O_873,N_49895,N_49969);
xor UO_874 (O_874,N_49767,N_49828);
xor UO_875 (O_875,N_49766,N_49967);
nor UO_876 (O_876,N_49789,N_49753);
nor UO_877 (O_877,N_49976,N_49994);
nor UO_878 (O_878,N_49918,N_49833);
nand UO_879 (O_879,N_49988,N_49955);
nor UO_880 (O_880,N_49924,N_49802);
xor UO_881 (O_881,N_49978,N_49871);
xor UO_882 (O_882,N_49809,N_49796);
nand UO_883 (O_883,N_49965,N_49947);
nor UO_884 (O_884,N_49977,N_49835);
and UO_885 (O_885,N_49893,N_49937);
xor UO_886 (O_886,N_49902,N_49874);
and UO_887 (O_887,N_49991,N_49880);
and UO_888 (O_888,N_49924,N_49897);
or UO_889 (O_889,N_49946,N_49763);
and UO_890 (O_890,N_49911,N_49876);
nor UO_891 (O_891,N_49877,N_49764);
and UO_892 (O_892,N_49893,N_49838);
nand UO_893 (O_893,N_49841,N_49853);
xor UO_894 (O_894,N_49840,N_49772);
nand UO_895 (O_895,N_49867,N_49771);
or UO_896 (O_896,N_49950,N_49763);
nor UO_897 (O_897,N_49870,N_49831);
and UO_898 (O_898,N_49765,N_49867);
nor UO_899 (O_899,N_49787,N_49843);
and UO_900 (O_900,N_49887,N_49807);
nor UO_901 (O_901,N_49830,N_49980);
nand UO_902 (O_902,N_49987,N_49854);
nor UO_903 (O_903,N_49849,N_49883);
and UO_904 (O_904,N_49952,N_49914);
and UO_905 (O_905,N_49879,N_49867);
or UO_906 (O_906,N_49906,N_49921);
nand UO_907 (O_907,N_49892,N_49828);
and UO_908 (O_908,N_49899,N_49924);
xnor UO_909 (O_909,N_49898,N_49814);
xor UO_910 (O_910,N_49751,N_49847);
or UO_911 (O_911,N_49899,N_49786);
or UO_912 (O_912,N_49834,N_49948);
nor UO_913 (O_913,N_49876,N_49988);
nor UO_914 (O_914,N_49978,N_49966);
xnor UO_915 (O_915,N_49911,N_49915);
nand UO_916 (O_916,N_49875,N_49957);
nor UO_917 (O_917,N_49911,N_49759);
nor UO_918 (O_918,N_49860,N_49853);
xnor UO_919 (O_919,N_49783,N_49920);
xor UO_920 (O_920,N_49947,N_49915);
nor UO_921 (O_921,N_49753,N_49811);
xor UO_922 (O_922,N_49971,N_49831);
and UO_923 (O_923,N_49769,N_49868);
or UO_924 (O_924,N_49933,N_49859);
xor UO_925 (O_925,N_49939,N_49787);
nor UO_926 (O_926,N_49959,N_49931);
nor UO_927 (O_927,N_49962,N_49793);
xnor UO_928 (O_928,N_49884,N_49810);
and UO_929 (O_929,N_49965,N_49901);
and UO_930 (O_930,N_49991,N_49977);
or UO_931 (O_931,N_49750,N_49882);
nor UO_932 (O_932,N_49803,N_49783);
xor UO_933 (O_933,N_49905,N_49920);
nor UO_934 (O_934,N_49837,N_49825);
nand UO_935 (O_935,N_49912,N_49956);
nor UO_936 (O_936,N_49825,N_49854);
xnor UO_937 (O_937,N_49768,N_49914);
and UO_938 (O_938,N_49818,N_49837);
and UO_939 (O_939,N_49832,N_49755);
and UO_940 (O_940,N_49835,N_49789);
and UO_941 (O_941,N_49855,N_49776);
xnor UO_942 (O_942,N_49860,N_49980);
nor UO_943 (O_943,N_49767,N_49978);
nor UO_944 (O_944,N_49820,N_49840);
or UO_945 (O_945,N_49750,N_49993);
and UO_946 (O_946,N_49973,N_49924);
and UO_947 (O_947,N_49904,N_49837);
xnor UO_948 (O_948,N_49814,N_49995);
or UO_949 (O_949,N_49955,N_49778);
nand UO_950 (O_950,N_49986,N_49920);
xor UO_951 (O_951,N_49948,N_49931);
and UO_952 (O_952,N_49788,N_49790);
nor UO_953 (O_953,N_49853,N_49815);
xnor UO_954 (O_954,N_49782,N_49788);
nand UO_955 (O_955,N_49811,N_49884);
xnor UO_956 (O_956,N_49969,N_49996);
nor UO_957 (O_957,N_49872,N_49831);
nor UO_958 (O_958,N_49824,N_49954);
nor UO_959 (O_959,N_49936,N_49841);
or UO_960 (O_960,N_49798,N_49933);
nand UO_961 (O_961,N_49909,N_49857);
xor UO_962 (O_962,N_49840,N_49944);
nand UO_963 (O_963,N_49759,N_49791);
nor UO_964 (O_964,N_49998,N_49777);
nand UO_965 (O_965,N_49904,N_49920);
and UO_966 (O_966,N_49758,N_49767);
xnor UO_967 (O_967,N_49922,N_49934);
xor UO_968 (O_968,N_49764,N_49969);
nand UO_969 (O_969,N_49839,N_49942);
or UO_970 (O_970,N_49897,N_49934);
or UO_971 (O_971,N_49870,N_49920);
nor UO_972 (O_972,N_49782,N_49804);
nand UO_973 (O_973,N_49837,N_49950);
nand UO_974 (O_974,N_49848,N_49752);
nand UO_975 (O_975,N_49906,N_49937);
nand UO_976 (O_976,N_49991,N_49961);
xnor UO_977 (O_977,N_49753,N_49981);
nand UO_978 (O_978,N_49824,N_49956);
nand UO_979 (O_979,N_49993,N_49773);
nor UO_980 (O_980,N_49755,N_49971);
nor UO_981 (O_981,N_49910,N_49784);
and UO_982 (O_982,N_49983,N_49756);
nand UO_983 (O_983,N_49787,N_49769);
or UO_984 (O_984,N_49905,N_49774);
xnor UO_985 (O_985,N_49836,N_49931);
or UO_986 (O_986,N_49933,N_49758);
xnor UO_987 (O_987,N_49973,N_49824);
or UO_988 (O_988,N_49849,N_49995);
and UO_989 (O_989,N_49831,N_49871);
and UO_990 (O_990,N_49798,N_49877);
and UO_991 (O_991,N_49999,N_49811);
nand UO_992 (O_992,N_49771,N_49872);
or UO_993 (O_993,N_49881,N_49752);
or UO_994 (O_994,N_49852,N_49953);
nand UO_995 (O_995,N_49795,N_49787);
xor UO_996 (O_996,N_49861,N_49956);
nand UO_997 (O_997,N_49813,N_49829);
and UO_998 (O_998,N_49908,N_49762);
and UO_999 (O_999,N_49872,N_49867);
nand UO_1000 (O_1000,N_49944,N_49752);
or UO_1001 (O_1001,N_49990,N_49847);
nand UO_1002 (O_1002,N_49828,N_49925);
or UO_1003 (O_1003,N_49901,N_49991);
or UO_1004 (O_1004,N_49901,N_49852);
nor UO_1005 (O_1005,N_49790,N_49974);
nor UO_1006 (O_1006,N_49928,N_49821);
nand UO_1007 (O_1007,N_49927,N_49916);
nand UO_1008 (O_1008,N_49926,N_49782);
nor UO_1009 (O_1009,N_49814,N_49891);
nand UO_1010 (O_1010,N_49965,N_49823);
nand UO_1011 (O_1011,N_49794,N_49983);
and UO_1012 (O_1012,N_49888,N_49962);
or UO_1013 (O_1013,N_49813,N_49875);
or UO_1014 (O_1014,N_49934,N_49962);
nor UO_1015 (O_1015,N_49773,N_49758);
nor UO_1016 (O_1016,N_49762,N_49751);
nand UO_1017 (O_1017,N_49876,N_49950);
and UO_1018 (O_1018,N_49937,N_49810);
and UO_1019 (O_1019,N_49949,N_49810);
or UO_1020 (O_1020,N_49992,N_49885);
nand UO_1021 (O_1021,N_49905,N_49961);
nand UO_1022 (O_1022,N_49950,N_49791);
xnor UO_1023 (O_1023,N_49890,N_49908);
and UO_1024 (O_1024,N_49955,N_49961);
and UO_1025 (O_1025,N_49829,N_49945);
nand UO_1026 (O_1026,N_49773,N_49906);
or UO_1027 (O_1027,N_49894,N_49757);
or UO_1028 (O_1028,N_49819,N_49781);
nor UO_1029 (O_1029,N_49832,N_49921);
and UO_1030 (O_1030,N_49922,N_49884);
nand UO_1031 (O_1031,N_49844,N_49802);
and UO_1032 (O_1032,N_49769,N_49801);
or UO_1033 (O_1033,N_49913,N_49922);
or UO_1034 (O_1034,N_49782,N_49880);
and UO_1035 (O_1035,N_49971,N_49883);
nor UO_1036 (O_1036,N_49768,N_49830);
nor UO_1037 (O_1037,N_49864,N_49816);
or UO_1038 (O_1038,N_49986,N_49917);
or UO_1039 (O_1039,N_49914,N_49863);
or UO_1040 (O_1040,N_49960,N_49860);
xnor UO_1041 (O_1041,N_49900,N_49763);
or UO_1042 (O_1042,N_49753,N_49884);
nand UO_1043 (O_1043,N_49765,N_49803);
nor UO_1044 (O_1044,N_49948,N_49941);
nor UO_1045 (O_1045,N_49840,N_49947);
xor UO_1046 (O_1046,N_49778,N_49782);
xnor UO_1047 (O_1047,N_49992,N_49919);
and UO_1048 (O_1048,N_49838,N_49930);
xnor UO_1049 (O_1049,N_49948,N_49762);
or UO_1050 (O_1050,N_49834,N_49980);
or UO_1051 (O_1051,N_49751,N_49991);
xor UO_1052 (O_1052,N_49856,N_49930);
nor UO_1053 (O_1053,N_49776,N_49990);
and UO_1054 (O_1054,N_49964,N_49960);
nand UO_1055 (O_1055,N_49973,N_49862);
and UO_1056 (O_1056,N_49816,N_49879);
or UO_1057 (O_1057,N_49786,N_49777);
xnor UO_1058 (O_1058,N_49957,N_49847);
nand UO_1059 (O_1059,N_49895,N_49947);
nor UO_1060 (O_1060,N_49888,N_49975);
or UO_1061 (O_1061,N_49862,N_49879);
nor UO_1062 (O_1062,N_49815,N_49932);
or UO_1063 (O_1063,N_49777,N_49932);
xnor UO_1064 (O_1064,N_49891,N_49836);
nand UO_1065 (O_1065,N_49898,N_49926);
or UO_1066 (O_1066,N_49860,N_49972);
xor UO_1067 (O_1067,N_49882,N_49839);
xnor UO_1068 (O_1068,N_49881,N_49755);
xor UO_1069 (O_1069,N_49908,N_49923);
and UO_1070 (O_1070,N_49932,N_49992);
and UO_1071 (O_1071,N_49796,N_49979);
xnor UO_1072 (O_1072,N_49833,N_49876);
and UO_1073 (O_1073,N_49787,N_49944);
or UO_1074 (O_1074,N_49839,N_49875);
xnor UO_1075 (O_1075,N_49778,N_49921);
xnor UO_1076 (O_1076,N_49803,N_49894);
nand UO_1077 (O_1077,N_49900,N_49780);
nor UO_1078 (O_1078,N_49861,N_49874);
and UO_1079 (O_1079,N_49776,N_49779);
or UO_1080 (O_1080,N_49954,N_49818);
nor UO_1081 (O_1081,N_49903,N_49886);
xor UO_1082 (O_1082,N_49793,N_49776);
xor UO_1083 (O_1083,N_49768,N_49767);
nor UO_1084 (O_1084,N_49851,N_49979);
nor UO_1085 (O_1085,N_49904,N_49929);
nand UO_1086 (O_1086,N_49912,N_49853);
nand UO_1087 (O_1087,N_49918,N_49842);
nor UO_1088 (O_1088,N_49863,N_49915);
xnor UO_1089 (O_1089,N_49839,N_49816);
or UO_1090 (O_1090,N_49906,N_49909);
nand UO_1091 (O_1091,N_49872,N_49932);
or UO_1092 (O_1092,N_49982,N_49865);
xor UO_1093 (O_1093,N_49961,N_49819);
nor UO_1094 (O_1094,N_49836,N_49999);
nand UO_1095 (O_1095,N_49990,N_49806);
xnor UO_1096 (O_1096,N_49973,N_49944);
xnor UO_1097 (O_1097,N_49864,N_49793);
and UO_1098 (O_1098,N_49852,N_49910);
nor UO_1099 (O_1099,N_49904,N_49944);
and UO_1100 (O_1100,N_49828,N_49760);
xnor UO_1101 (O_1101,N_49917,N_49766);
and UO_1102 (O_1102,N_49892,N_49753);
nand UO_1103 (O_1103,N_49842,N_49997);
and UO_1104 (O_1104,N_49999,N_49801);
or UO_1105 (O_1105,N_49804,N_49963);
nand UO_1106 (O_1106,N_49857,N_49976);
or UO_1107 (O_1107,N_49800,N_49766);
xnor UO_1108 (O_1108,N_49810,N_49853);
and UO_1109 (O_1109,N_49818,N_49963);
nand UO_1110 (O_1110,N_49864,N_49763);
or UO_1111 (O_1111,N_49932,N_49751);
or UO_1112 (O_1112,N_49780,N_49914);
nand UO_1113 (O_1113,N_49864,N_49853);
nor UO_1114 (O_1114,N_49945,N_49846);
nand UO_1115 (O_1115,N_49818,N_49937);
or UO_1116 (O_1116,N_49760,N_49836);
nand UO_1117 (O_1117,N_49800,N_49932);
or UO_1118 (O_1118,N_49765,N_49965);
nor UO_1119 (O_1119,N_49972,N_49906);
or UO_1120 (O_1120,N_49774,N_49789);
nor UO_1121 (O_1121,N_49848,N_49757);
or UO_1122 (O_1122,N_49920,N_49785);
xnor UO_1123 (O_1123,N_49979,N_49906);
and UO_1124 (O_1124,N_49765,N_49838);
nand UO_1125 (O_1125,N_49923,N_49918);
or UO_1126 (O_1126,N_49769,N_49959);
nand UO_1127 (O_1127,N_49981,N_49885);
xnor UO_1128 (O_1128,N_49824,N_49862);
or UO_1129 (O_1129,N_49920,N_49944);
and UO_1130 (O_1130,N_49787,N_49994);
xor UO_1131 (O_1131,N_49863,N_49860);
nor UO_1132 (O_1132,N_49828,N_49777);
or UO_1133 (O_1133,N_49872,N_49978);
nor UO_1134 (O_1134,N_49984,N_49850);
nor UO_1135 (O_1135,N_49754,N_49812);
or UO_1136 (O_1136,N_49974,N_49794);
nand UO_1137 (O_1137,N_49972,N_49779);
or UO_1138 (O_1138,N_49957,N_49864);
nor UO_1139 (O_1139,N_49761,N_49845);
xnor UO_1140 (O_1140,N_49883,N_49783);
and UO_1141 (O_1141,N_49927,N_49992);
nor UO_1142 (O_1142,N_49854,N_49793);
or UO_1143 (O_1143,N_49807,N_49815);
nand UO_1144 (O_1144,N_49987,N_49970);
and UO_1145 (O_1145,N_49990,N_49815);
xnor UO_1146 (O_1146,N_49812,N_49776);
nor UO_1147 (O_1147,N_49967,N_49873);
and UO_1148 (O_1148,N_49754,N_49887);
nand UO_1149 (O_1149,N_49857,N_49935);
xor UO_1150 (O_1150,N_49963,N_49920);
or UO_1151 (O_1151,N_49949,N_49978);
or UO_1152 (O_1152,N_49822,N_49864);
or UO_1153 (O_1153,N_49897,N_49967);
xnor UO_1154 (O_1154,N_49971,N_49951);
nand UO_1155 (O_1155,N_49994,N_49942);
xor UO_1156 (O_1156,N_49921,N_49868);
xnor UO_1157 (O_1157,N_49870,N_49953);
or UO_1158 (O_1158,N_49941,N_49825);
xor UO_1159 (O_1159,N_49917,N_49985);
nand UO_1160 (O_1160,N_49871,N_49952);
nor UO_1161 (O_1161,N_49777,N_49896);
nand UO_1162 (O_1162,N_49824,N_49813);
nand UO_1163 (O_1163,N_49915,N_49833);
and UO_1164 (O_1164,N_49877,N_49914);
nor UO_1165 (O_1165,N_49971,N_49875);
or UO_1166 (O_1166,N_49757,N_49763);
nand UO_1167 (O_1167,N_49930,N_49816);
xor UO_1168 (O_1168,N_49838,N_49968);
or UO_1169 (O_1169,N_49827,N_49771);
nor UO_1170 (O_1170,N_49884,N_49863);
xnor UO_1171 (O_1171,N_49958,N_49955);
xnor UO_1172 (O_1172,N_49923,N_49896);
xor UO_1173 (O_1173,N_49770,N_49868);
or UO_1174 (O_1174,N_49840,N_49850);
nand UO_1175 (O_1175,N_49819,N_49921);
or UO_1176 (O_1176,N_49796,N_49893);
or UO_1177 (O_1177,N_49789,N_49948);
xnor UO_1178 (O_1178,N_49835,N_49908);
nand UO_1179 (O_1179,N_49802,N_49933);
nor UO_1180 (O_1180,N_49999,N_49850);
xor UO_1181 (O_1181,N_49938,N_49907);
and UO_1182 (O_1182,N_49981,N_49893);
xor UO_1183 (O_1183,N_49835,N_49842);
xor UO_1184 (O_1184,N_49773,N_49796);
nand UO_1185 (O_1185,N_49978,N_49922);
or UO_1186 (O_1186,N_49758,N_49806);
nor UO_1187 (O_1187,N_49759,N_49868);
or UO_1188 (O_1188,N_49786,N_49970);
nand UO_1189 (O_1189,N_49895,N_49873);
and UO_1190 (O_1190,N_49881,N_49996);
and UO_1191 (O_1191,N_49752,N_49938);
nor UO_1192 (O_1192,N_49789,N_49776);
nor UO_1193 (O_1193,N_49838,N_49761);
and UO_1194 (O_1194,N_49774,N_49790);
or UO_1195 (O_1195,N_49913,N_49751);
nor UO_1196 (O_1196,N_49966,N_49778);
and UO_1197 (O_1197,N_49794,N_49821);
xor UO_1198 (O_1198,N_49904,N_49952);
xor UO_1199 (O_1199,N_49824,N_49836);
nand UO_1200 (O_1200,N_49870,N_49801);
and UO_1201 (O_1201,N_49752,N_49772);
or UO_1202 (O_1202,N_49879,N_49824);
nand UO_1203 (O_1203,N_49795,N_49907);
or UO_1204 (O_1204,N_49775,N_49893);
nand UO_1205 (O_1205,N_49801,N_49794);
xnor UO_1206 (O_1206,N_49855,N_49970);
and UO_1207 (O_1207,N_49979,N_49888);
and UO_1208 (O_1208,N_49938,N_49820);
and UO_1209 (O_1209,N_49843,N_49865);
and UO_1210 (O_1210,N_49818,N_49855);
and UO_1211 (O_1211,N_49951,N_49826);
xnor UO_1212 (O_1212,N_49950,N_49820);
nand UO_1213 (O_1213,N_49812,N_49962);
nand UO_1214 (O_1214,N_49984,N_49839);
and UO_1215 (O_1215,N_49790,N_49966);
nand UO_1216 (O_1216,N_49883,N_49867);
nor UO_1217 (O_1217,N_49755,N_49936);
nor UO_1218 (O_1218,N_49899,N_49883);
and UO_1219 (O_1219,N_49937,N_49792);
nor UO_1220 (O_1220,N_49900,N_49865);
and UO_1221 (O_1221,N_49998,N_49962);
and UO_1222 (O_1222,N_49799,N_49948);
xnor UO_1223 (O_1223,N_49837,N_49856);
nand UO_1224 (O_1224,N_49788,N_49834);
xnor UO_1225 (O_1225,N_49778,N_49971);
xor UO_1226 (O_1226,N_49929,N_49866);
or UO_1227 (O_1227,N_49848,N_49760);
and UO_1228 (O_1228,N_49942,N_49961);
or UO_1229 (O_1229,N_49830,N_49943);
and UO_1230 (O_1230,N_49977,N_49885);
or UO_1231 (O_1231,N_49754,N_49780);
xnor UO_1232 (O_1232,N_49930,N_49968);
nor UO_1233 (O_1233,N_49953,N_49837);
or UO_1234 (O_1234,N_49937,N_49959);
or UO_1235 (O_1235,N_49800,N_49980);
nand UO_1236 (O_1236,N_49833,N_49789);
or UO_1237 (O_1237,N_49981,N_49828);
nand UO_1238 (O_1238,N_49828,N_49759);
or UO_1239 (O_1239,N_49924,N_49951);
nand UO_1240 (O_1240,N_49954,N_49870);
or UO_1241 (O_1241,N_49762,N_49930);
and UO_1242 (O_1242,N_49931,N_49903);
nand UO_1243 (O_1243,N_49788,N_49830);
nor UO_1244 (O_1244,N_49832,N_49951);
and UO_1245 (O_1245,N_49752,N_49779);
xor UO_1246 (O_1246,N_49969,N_49970);
nor UO_1247 (O_1247,N_49755,N_49968);
and UO_1248 (O_1248,N_49814,N_49810);
nand UO_1249 (O_1249,N_49928,N_49795);
xor UO_1250 (O_1250,N_49849,N_49763);
and UO_1251 (O_1251,N_49960,N_49853);
nand UO_1252 (O_1252,N_49890,N_49779);
or UO_1253 (O_1253,N_49887,N_49951);
xor UO_1254 (O_1254,N_49993,N_49867);
nor UO_1255 (O_1255,N_49751,N_49852);
nand UO_1256 (O_1256,N_49830,N_49968);
or UO_1257 (O_1257,N_49974,N_49836);
xor UO_1258 (O_1258,N_49850,N_49961);
nor UO_1259 (O_1259,N_49784,N_49788);
xnor UO_1260 (O_1260,N_49869,N_49938);
and UO_1261 (O_1261,N_49785,N_49910);
xnor UO_1262 (O_1262,N_49876,N_49977);
and UO_1263 (O_1263,N_49799,N_49996);
nor UO_1264 (O_1264,N_49910,N_49991);
xnor UO_1265 (O_1265,N_49753,N_49859);
or UO_1266 (O_1266,N_49956,N_49942);
and UO_1267 (O_1267,N_49779,N_49921);
and UO_1268 (O_1268,N_49793,N_49827);
nand UO_1269 (O_1269,N_49811,N_49924);
nand UO_1270 (O_1270,N_49875,N_49800);
or UO_1271 (O_1271,N_49975,N_49892);
nor UO_1272 (O_1272,N_49843,N_49967);
and UO_1273 (O_1273,N_49887,N_49950);
nor UO_1274 (O_1274,N_49891,N_49886);
nand UO_1275 (O_1275,N_49971,N_49790);
nand UO_1276 (O_1276,N_49954,N_49960);
xor UO_1277 (O_1277,N_49892,N_49811);
nor UO_1278 (O_1278,N_49979,N_49810);
and UO_1279 (O_1279,N_49954,N_49833);
xnor UO_1280 (O_1280,N_49786,N_49918);
xor UO_1281 (O_1281,N_49825,N_49974);
or UO_1282 (O_1282,N_49884,N_49964);
nor UO_1283 (O_1283,N_49875,N_49959);
and UO_1284 (O_1284,N_49817,N_49936);
xor UO_1285 (O_1285,N_49919,N_49757);
and UO_1286 (O_1286,N_49957,N_49775);
or UO_1287 (O_1287,N_49913,N_49977);
nor UO_1288 (O_1288,N_49928,N_49883);
or UO_1289 (O_1289,N_49944,N_49939);
xnor UO_1290 (O_1290,N_49752,N_49766);
nand UO_1291 (O_1291,N_49906,N_49963);
and UO_1292 (O_1292,N_49998,N_49980);
or UO_1293 (O_1293,N_49860,N_49913);
nor UO_1294 (O_1294,N_49858,N_49900);
nor UO_1295 (O_1295,N_49790,N_49815);
or UO_1296 (O_1296,N_49821,N_49893);
or UO_1297 (O_1297,N_49994,N_49888);
or UO_1298 (O_1298,N_49903,N_49844);
and UO_1299 (O_1299,N_49912,N_49873);
or UO_1300 (O_1300,N_49770,N_49761);
nand UO_1301 (O_1301,N_49884,N_49820);
and UO_1302 (O_1302,N_49931,N_49798);
and UO_1303 (O_1303,N_49930,N_49903);
nor UO_1304 (O_1304,N_49941,N_49924);
nor UO_1305 (O_1305,N_49859,N_49996);
nand UO_1306 (O_1306,N_49827,N_49910);
and UO_1307 (O_1307,N_49758,N_49785);
nand UO_1308 (O_1308,N_49860,N_49969);
nor UO_1309 (O_1309,N_49782,N_49860);
xor UO_1310 (O_1310,N_49883,N_49947);
nand UO_1311 (O_1311,N_49866,N_49897);
nand UO_1312 (O_1312,N_49876,N_49781);
or UO_1313 (O_1313,N_49890,N_49823);
nor UO_1314 (O_1314,N_49761,N_49972);
nand UO_1315 (O_1315,N_49802,N_49856);
nand UO_1316 (O_1316,N_49952,N_49910);
xnor UO_1317 (O_1317,N_49790,N_49795);
nand UO_1318 (O_1318,N_49982,N_49815);
and UO_1319 (O_1319,N_49851,N_49900);
nor UO_1320 (O_1320,N_49852,N_49872);
or UO_1321 (O_1321,N_49903,N_49960);
nor UO_1322 (O_1322,N_49924,N_49876);
or UO_1323 (O_1323,N_49775,N_49895);
nand UO_1324 (O_1324,N_49817,N_49959);
nor UO_1325 (O_1325,N_49793,N_49981);
nor UO_1326 (O_1326,N_49780,N_49989);
nand UO_1327 (O_1327,N_49958,N_49814);
xor UO_1328 (O_1328,N_49912,N_49971);
or UO_1329 (O_1329,N_49836,N_49902);
xor UO_1330 (O_1330,N_49782,N_49950);
or UO_1331 (O_1331,N_49898,N_49955);
or UO_1332 (O_1332,N_49894,N_49978);
nor UO_1333 (O_1333,N_49909,N_49842);
nor UO_1334 (O_1334,N_49828,N_49820);
or UO_1335 (O_1335,N_49844,N_49856);
and UO_1336 (O_1336,N_49835,N_49921);
xnor UO_1337 (O_1337,N_49902,N_49762);
or UO_1338 (O_1338,N_49801,N_49776);
or UO_1339 (O_1339,N_49810,N_49834);
nand UO_1340 (O_1340,N_49894,N_49977);
and UO_1341 (O_1341,N_49904,N_49900);
or UO_1342 (O_1342,N_49768,N_49983);
nor UO_1343 (O_1343,N_49820,N_49853);
nand UO_1344 (O_1344,N_49885,N_49946);
nand UO_1345 (O_1345,N_49858,N_49844);
nor UO_1346 (O_1346,N_49819,N_49750);
nor UO_1347 (O_1347,N_49902,N_49872);
nand UO_1348 (O_1348,N_49971,N_49879);
nor UO_1349 (O_1349,N_49778,N_49776);
xor UO_1350 (O_1350,N_49989,N_49854);
or UO_1351 (O_1351,N_49787,N_49794);
xor UO_1352 (O_1352,N_49861,N_49763);
nor UO_1353 (O_1353,N_49925,N_49923);
or UO_1354 (O_1354,N_49766,N_49818);
xnor UO_1355 (O_1355,N_49752,N_49995);
nand UO_1356 (O_1356,N_49990,N_49981);
nand UO_1357 (O_1357,N_49921,N_49804);
nand UO_1358 (O_1358,N_49769,N_49873);
nor UO_1359 (O_1359,N_49866,N_49946);
xor UO_1360 (O_1360,N_49985,N_49970);
or UO_1361 (O_1361,N_49870,N_49938);
and UO_1362 (O_1362,N_49903,N_49836);
nor UO_1363 (O_1363,N_49929,N_49803);
nand UO_1364 (O_1364,N_49844,N_49921);
xnor UO_1365 (O_1365,N_49855,N_49817);
xor UO_1366 (O_1366,N_49806,N_49911);
nor UO_1367 (O_1367,N_49994,N_49878);
nor UO_1368 (O_1368,N_49873,N_49776);
nand UO_1369 (O_1369,N_49930,N_49825);
and UO_1370 (O_1370,N_49940,N_49816);
nor UO_1371 (O_1371,N_49948,N_49901);
nand UO_1372 (O_1372,N_49778,N_49825);
or UO_1373 (O_1373,N_49949,N_49838);
and UO_1374 (O_1374,N_49807,N_49762);
nand UO_1375 (O_1375,N_49899,N_49768);
or UO_1376 (O_1376,N_49912,N_49972);
nor UO_1377 (O_1377,N_49918,N_49856);
or UO_1378 (O_1378,N_49987,N_49892);
xnor UO_1379 (O_1379,N_49875,N_49969);
nand UO_1380 (O_1380,N_49755,N_49753);
nor UO_1381 (O_1381,N_49852,N_49947);
xnor UO_1382 (O_1382,N_49878,N_49938);
nand UO_1383 (O_1383,N_49864,N_49991);
or UO_1384 (O_1384,N_49924,N_49763);
and UO_1385 (O_1385,N_49808,N_49897);
nand UO_1386 (O_1386,N_49826,N_49975);
or UO_1387 (O_1387,N_49792,N_49883);
nor UO_1388 (O_1388,N_49770,N_49865);
xnor UO_1389 (O_1389,N_49898,N_49888);
xor UO_1390 (O_1390,N_49752,N_49805);
and UO_1391 (O_1391,N_49944,N_49938);
or UO_1392 (O_1392,N_49770,N_49916);
xor UO_1393 (O_1393,N_49790,N_49879);
or UO_1394 (O_1394,N_49972,N_49832);
nor UO_1395 (O_1395,N_49961,N_49827);
or UO_1396 (O_1396,N_49986,N_49801);
xor UO_1397 (O_1397,N_49810,N_49859);
or UO_1398 (O_1398,N_49810,N_49811);
nand UO_1399 (O_1399,N_49828,N_49787);
nand UO_1400 (O_1400,N_49980,N_49951);
nand UO_1401 (O_1401,N_49805,N_49987);
or UO_1402 (O_1402,N_49772,N_49953);
and UO_1403 (O_1403,N_49854,N_49769);
xnor UO_1404 (O_1404,N_49969,N_49878);
and UO_1405 (O_1405,N_49990,N_49818);
nor UO_1406 (O_1406,N_49982,N_49762);
and UO_1407 (O_1407,N_49987,N_49998);
xnor UO_1408 (O_1408,N_49918,N_49863);
and UO_1409 (O_1409,N_49856,N_49972);
nand UO_1410 (O_1410,N_49963,N_49942);
or UO_1411 (O_1411,N_49909,N_49931);
or UO_1412 (O_1412,N_49835,N_49801);
nand UO_1413 (O_1413,N_49977,N_49934);
nand UO_1414 (O_1414,N_49961,N_49877);
or UO_1415 (O_1415,N_49953,N_49788);
nor UO_1416 (O_1416,N_49898,N_49766);
and UO_1417 (O_1417,N_49850,N_49880);
and UO_1418 (O_1418,N_49926,N_49874);
nand UO_1419 (O_1419,N_49866,N_49944);
and UO_1420 (O_1420,N_49817,N_49856);
nand UO_1421 (O_1421,N_49799,N_49869);
and UO_1422 (O_1422,N_49918,N_49910);
nor UO_1423 (O_1423,N_49976,N_49850);
or UO_1424 (O_1424,N_49838,N_49936);
nor UO_1425 (O_1425,N_49892,N_49954);
nand UO_1426 (O_1426,N_49938,N_49921);
nand UO_1427 (O_1427,N_49834,N_49899);
or UO_1428 (O_1428,N_49787,N_49982);
or UO_1429 (O_1429,N_49879,N_49889);
xor UO_1430 (O_1430,N_49978,N_49847);
nor UO_1431 (O_1431,N_49995,N_49845);
or UO_1432 (O_1432,N_49972,N_49813);
and UO_1433 (O_1433,N_49858,N_49990);
or UO_1434 (O_1434,N_49812,N_49814);
xnor UO_1435 (O_1435,N_49861,N_49970);
nand UO_1436 (O_1436,N_49905,N_49821);
and UO_1437 (O_1437,N_49982,N_49915);
or UO_1438 (O_1438,N_49998,N_49975);
xnor UO_1439 (O_1439,N_49902,N_49832);
nor UO_1440 (O_1440,N_49946,N_49882);
xor UO_1441 (O_1441,N_49848,N_49858);
nand UO_1442 (O_1442,N_49917,N_49962);
nand UO_1443 (O_1443,N_49961,N_49786);
nand UO_1444 (O_1444,N_49823,N_49854);
and UO_1445 (O_1445,N_49778,N_49812);
or UO_1446 (O_1446,N_49993,N_49771);
nor UO_1447 (O_1447,N_49771,N_49979);
nor UO_1448 (O_1448,N_49884,N_49981);
or UO_1449 (O_1449,N_49926,N_49896);
nor UO_1450 (O_1450,N_49762,N_49978);
and UO_1451 (O_1451,N_49945,N_49847);
xor UO_1452 (O_1452,N_49844,N_49809);
or UO_1453 (O_1453,N_49828,N_49985);
nor UO_1454 (O_1454,N_49911,N_49762);
nand UO_1455 (O_1455,N_49920,N_49924);
and UO_1456 (O_1456,N_49848,N_49968);
and UO_1457 (O_1457,N_49854,N_49962);
and UO_1458 (O_1458,N_49777,N_49809);
and UO_1459 (O_1459,N_49776,N_49959);
nand UO_1460 (O_1460,N_49834,N_49910);
nand UO_1461 (O_1461,N_49883,N_49853);
nor UO_1462 (O_1462,N_49977,N_49853);
nor UO_1463 (O_1463,N_49821,N_49953);
or UO_1464 (O_1464,N_49956,N_49845);
nor UO_1465 (O_1465,N_49970,N_49993);
nor UO_1466 (O_1466,N_49928,N_49877);
xor UO_1467 (O_1467,N_49753,N_49960);
nand UO_1468 (O_1468,N_49750,N_49796);
nor UO_1469 (O_1469,N_49881,N_49882);
or UO_1470 (O_1470,N_49982,N_49956);
or UO_1471 (O_1471,N_49887,N_49812);
nand UO_1472 (O_1472,N_49950,N_49949);
nand UO_1473 (O_1473,N_49799,N_49793);
or UO_1474 (O_1474,N_49959,N_49998);
and UO_1475 (O_1475,N_49931,N_49837);
and UO_1476 (O_1476,N_49834,N_49799);
or UO_1477 (O_1477,N_49836,N_49986);
and UO_1478 (O_1478,N_49760,N_49928);
nor UO_1479 (O_1479,N_49828,N_49865);
xnor UO_1480 (O_1480,N_49760,N_49853);
or UO_1481 (O_1481,N_49911,N_49929);
xnor UO_1482 (O_1482,N_49830,N_49898);
or UO_1483 (O_1483,N_49943,N_49918);
nand UO_1484 (O_1484,N_49772,N_49844);
nor UO_1485 (O_1485,N_49870,N_49800);
nor UO_1486 (O_1486,N_49815,N_49875);
xor UO_1487 (O_1487,N_49913,N_49930);
nor UO_1488 (O_1488,N_49829,N_49935);
nor UO_1489 (O_1489,N_49779,N_49790);
xor UO_1490 (O_1490,N_49811,N_49788);
nor UO_1491 (O_1491,N_49995,N_49827);
xnor UO_1492 (O_1492,N_49756,N_49813);
nand UO_1493 (O_1493,N_49814,N_49763);
nor UO_1494 (O_1494,N_49929,N_49989);
and UO_1495 (O_1495,N_49991,N_49913);
or UO_1496 (O_1496,N_49960,N_49794);
nor UO_1497 (O_1497,N_49851,N_49853);
nor UO_1498 (O_1498,N_49999,N_49812);
xnor UO_1499 (O_1499,N_49792,N_49888);
or UO_1500 (O_1500,N_49808,N_49849);
xnor UO_1501 (O_1501,N_49892,N_49902);
nand UO_1502 (O_1502,N_49783,N_49991);
or UO_1503 (O_1503,N_49817,N_49973);
xnor UO_1504 (O_1504,N_49960,N_49809);
and UO_1505 (O_1505,N_49949,N_49938);
nand UO_1506 (O_1506,N_49860,N_49865);
xnor UO_1507 (O_1507,N_49856,N_49931);
nor UO_1508 (O_1508,N_49896,N_49871);
nand UO_1509 (O_1509,N_49909,N_49959);
nor UO_1510 (O_1510,N_49979,N_49843);
or UO_1511 (O_1511,N_49894,N_49881);
or UO_1512 (O_1512,N_49840,N_49920);
nand UO_1513 (O_1513,N_49764,N_49792);
and UO_1514 (O_1514,N_49801,N_49972);
or UO_1515 (O_1515,N_49773,N_49846);
nor UO_1516 (O_1516,N_49833,N_49964);
or UO_1517 (O_1517,N_49921,N_49822);
nor UO_1518 (O_1518,N_49883,N_49898);
and UO_1519 (O_1519,N_49784,N_49751);
xor UO_1520 (O_1520,N_49983,N_49834);
nor UO_1521 (O_1521,N_49993,N_49912);
nand UO_1522 (O_1522,N_49915,N_49858);
nand UO_1523 (O_1523,N_49895,N_49942);
and UO_1524 (O_1524,N_49899,N_49898);
nand UO_1525 (O_1525,N_49965,N_49819);
nor UO_1526 (O_1526,N_49769,N_49896);
xnor UO_1527 (O_1527,N_49895,N_49822);
xor UO_1528 (O_1528,N_49805,N_49937);
nor UO_1529 (O_1529,N_49824,N_49932);
nor UO_1530 (O_1530,N_49846,N_49979);
xor UO_1531 (O_1531,N_49964,N_49956);
nor UO_1532 (O_1532,N_49927,N_49896);
xnor UO_1533 (O_1533,N_49826,N_49849);
or UO_1534 (O_1534,N_49769,N_49843);
or UO_1535 (O_1535,N_49887,N_49952);
and UO_1536 (O_1536,N_49998,N_49799);
xnor UO_1537 (O_1537,N_49855,N_49939);
and UO_1538 (O_1538,N_49775,N_49761);
or UO_1539 (O_1539,N_49783,N_49871);
or UO_1540 (O_1540,N_49771,N_49814);
and UO_1541 (O_1541,N_49777,N_49872);
nand UO_1542 (O_1542,N_49868,N_49895);
or UO_1543 (O_1543,N_49824,N_49876);
xnor UO_1544 (O_1544,N_49978,N_49826);
or UO_1545 (O_1545,N_49986,N_49987);
or UO_1546 (O_1546,N_49954,N_49840);
nor UO_1547 (O_1547,N_49859,N_49904);
and UO_1548 (O_1548,N_49850,N_49960);
nand UO_1549 (O_1549,N_49882,N_49751);
nand UO_1550 (O_1550,N_49889,N_49774);
xnor UO_1551 (O_1551,N_49871,N_49807);
nand UO_1552 (O_1552,N_49769,N_49764);
nand UO_1553 (O_1553,N_49899,N_49919);
xor UO_1554 (O_1554,N_49812,N_49875);
and UO_1555 (O_1555,N_49787,N_49925);
and UO_1556 (O_1556,N_49766,N_49980);
nand UO_1557 (O_1557,N_49820,N_49971);
nand UO_1558 (O_1558,N_49871,N_49909);
xnor UO_1559 (O_1559,N_49999,N_49853);
xnor UO_1560 (O_1560,N_49936,N_49825);
nor UO_1561 (O_1561,N_49899,N_49779);
or UO_1562 (O_1562,N_49802,N_49786);
and UO_1563 (O_1563,N_49913,N_49903);
xor UO_1564 (O_1564,N_49779,N_49990);
xnor UO_1565 (O_1565,N_49906,N_49796);
xor UO_1566 (O_1566,N_49842,N_49826);
nand UO_1567 (O_1567,N_49918,N_49855);
and UO_1568 (O_1568,N_49946,N_49752);
nand UO_1569 (O_1569,N_49985,N_49926);
nand UO_1570 (O_1570,N_49832,N_49799);
nor UO_1571 (O_1571,N_49775,N_49931);
nand UO_1572 (O_1572,N_49912,N_49804);
and UO_1573 (O_1573,N_49960,N_49874);
and UO_1574 (O_1574,N_49858,N_49950);
xor UO_1575 (O_1575,N_49759,N_49883);
nor UO_1576 (O_1576,N_49750,N_49895);
xor UO_1577 (O_1577,N_49965,N_49864);
xor UO_1578 (O_1578,N_49756,N_49879);
nand UO_1579 (O_1579,N_49966,N_49822);
nand UO_1580 (O_1580,N_49840,N_49997);
and UO_1581 (O_1581,N_49953,N_49776);
nand UO_1582 (O_1582,N_49937,N_49987);
nand UO_1583 (O_1583,N_49941,N_49894);
and UO_1584 (O_1584,N_49812,N_49995);
or UO_1585 (O_1585,N_49960,N_49933);
xor UO_1586 (O_1586,N_49819,N_49962);
nor UO_1587 (O_1587,N_49971,N_49958);
nand UO_1588 (O_1588,N_49950,N_49816);
xnor UO_1589 (O_1589,N_49933,N_49799);
and UO_1590 (O_1590,N_49846,N_49957);
or UO_1591 (O_1591,N_49942,N_49863);
or UO_1592 (O_1592,N_49909,N_49884);
xnor UO_1593 (O_1593,N_49952,N_49777);
nand UO_1594 (O_1594,N_49848,N_49809);
nor UO_1595 (O_1595,N_49924,N_49847);
and UO_1596 (O_1596,N_49783,N_49814);
xnor UO_1597 (O_1597,N_49974,N_49920);
nand UO_1598 (O_1598,N_49923,N_49899);
nand UO_1599 (O_1599,N_49972,N_49989);
or UO_1600 (O_1600,N_49891,N_49789);
or UO_1601 (O_1601,N_49905,N_49981);
nor UO_1602 (O_1602,N_49966,N_49983);
xor UO_1603 (O_1603,N_49798,N_49795);
and UO_1604 (O_1604,N_49820,N_49762);
nand UO_1605 (O_1605,N_49847,N_49939);
or UO_1606 (O_1606,N_49954,N_49987);
or UO_1607 (O_1607,N_49766,N_49943);
xnor UO_1608 (O_1608,N_49790,N_49753);
or UO_1609 (O_1609,N_49994,N_49970);
or UO_1610 (O_1610,N_49761,N_49882);
or UO_1611 (O_1611,N_49799,N_49814);
nor UO_1612 (O_1612,N_49919,N_49892);
and UO_1613 (O_1613,N_49779,N_49995);
nor UO_1614 (O_1614,N_49854,N_49942);
nand UO_1615 (O_1615,N_49758,N_49990);
nand UO_1616 (O_1616,N_49945,N_49893);
xor UO_1617 (O_1617,N_49867,N_49987);
xnor UO_1618 (O_1618,N_49903,N_49932);
xnor UO_1619 (O_1619,N_49883,N_49777);
nand UO_1620 (O_1620,N_49951,N_49881);
nand UO_1621 (O_1621,N_49831,N_49845);
nor UO_1622 (O_1622,N_49956,N_49986);
or UO_1623 (O_1623,N_49824,N_49961);
or UO_1624 (O_1624,N_49902,N_49792);
or UO_1625 (O_1625,N_49953,N_49929);
or UO_1626 (O_1626,N_49932,N_49791);
and UO_1627 (O_1627,N_49961,N_49771);
or UO_1628 (O_1628,N_49885,N_49900);
or UO_1629 (O_1629,N_49955,N_49923);
or UO_1630 (O_1630,N_49958,N_49864);
xor UO_1631 (O_1631,N_49778,N_49997);
nor UO_1632 (O_1632,N_49872,N_49968);
and UO_1633 (O_1633,N_49902,N_49802);
nand UO_1634 (O_1634,N_49916,N_49956);
xor UO_1635 (O_1635,N_49955,N_49937);
nand UO_1636 (O_1636,N_49976,N_49999);
nand UO_1637 (O_1637,N_49843,N_49998);
nor UO_1638 (O_1638,N_49971,N_49864);
or UO_1639 (O_1639,N_49887,N_49931);
nand UO_1640 (O_1640,N_49821,N_49833);
nor UO_1641 (O_1641,N_49795,N_49778);
nor UO_1642 (O_1642,N_49812,N_49808);
and UO_1643 (O_1643,N_49808,N_49915);
nor UO_1644 (O_1644,N_49864,N_49879);
or UO_1645 (O_1645,N_49982,N_49798);
or UO_1646 (O_1646,N_49753,N_49793);
nor UO_1647 (O_1647,N_49919,N_49985);
nand UO_1648 (O_1648,N_49995,N_49776);
nand UO_1649 (O_1649,N_49840,N_49888);
nor UO_1650 (O_1650,N_49822,N_49907);
or UO_1651 (O_1651,N_49808,N_49961);
or UO_1652 (O_1652,N_49790,N_49982);
and UO_1653 (O_1653,N_49896,N_49820);
nor UO_1654 (O_1654,N_49893,N_49998);
and UO_1655 (O_1655,N_49945,N_49992);
nor UO_1656 (O_1656,N_49781,N_49770);
nand UO_1657 (O_1657,N_49968,N_49920);
nor UO_1658 (O_1658,N_49991,N_49927);
nor UO_1659 (O_1659,N_49968,N_49795);
or UO_1660 (O_1660,N_49806,N_49819);
xnor UO_1661 (O_1661,N_49787,N_49832);
or UO_1662 (O_1662,N_49928,N_49827);
xor UO_1663 (O_1663,N_49837,N_49778);
or UO_1664 (O_1664,N_49770,N_49958);
xnor UO_1665 (O_1665,N_49870,N_49899);
xnor UO_1666 (O_1666,N_49752,N_49786);
or UO_1667 (O_1667,N_49827,N_49879);
xor UO_1668 (O_1668,N_49936,N_49907);
xnor UO_1669 (O_1669,N_49901,N_49827);
xnor UO_1670 (O_1670,N_49902,N_49926);
nand UO_1671 (O_1671,N_49909,N_49872);
nand UO_1672 (O_1672,N_49856,N_49923);
xnor UO_1673 (O_1673,N_49897,N_49912);
nor UO_1674 (O_1674,N_49940,N_49904);
nor UO_1675 (O_1675,N_49907,N_49842);
xor UO_1676 (O_1676,N_49872,N_49994);
and UO_1677 (O_1677,N_49964,N_49980);
nand UO_1678 (O_1678,N_49976,N_49862);
or UO_1679 (O_1679,N_49983,N_49922);
nor UO_1680 (O_1680,N_49778,N_49761);
or UO_1681 (O_1681,N_49857,N_49937);
and UO_1682 (O_1682,N_49840,N_49928);
nand UO_1683 (O_1683,N_49830,N_49903);
or UO_1684 (O_1684,N_49828,N_49864);
nand UO_1685 (O_1685,N_49962,N_49836);
nand UO_1686 (O_1686,N_49871,N_49825);
and UO_1687 (O_1687,N_49876,N_49770);
xor UO_1688 (O_1688,N_49766,N_49958);
xor UO_1689 (O_1689,N_49766,N_49848);
xor UO_1690 (O_1690,N_49841,N_49880);
or UO_1691 (O_1691,N_49936,N_49990);
nand UO_1692 (O_1692,N_49843,N_49868);
or UO_1693 (O_1693,N_49835,N_49903);
nand UO_1694 (O_1694,N_49913,N_49776);
nor UO_1695 (O_1695,N_49759,N_49851);
and UO_1696 (O_1696,N_49976,N_49884);
nand UO_1697 (O_1697,N_49776,N_49769);
nor UO_1698 (O_1698,N_49815,N_49979);
xnor UO_1699 (O_1699,N_49754,N_49959);
nor UO_1700 (O_1700,N_49809,N_49767);
xor UO_1701 (O_1701,N_49844,N_49972);
or UO_1702 (O_1702,N_49768,N_49978);
nand UO_1703 (O_1703,N_49832,N_49938);
nand UO_1704 (O_1704,N_49922,N_49805);
nand UO_1705 (O_1705,N_49837,N_49983);
or UO_1706 (O_1706,N_49980,N_49876);
nor UO_1707 (O_1707,N_49994,N_49963);
xnor UO_1708 (O_1708,N_49972,N_49833);
or UO_1709 (O_1709,N_49863,N_49845);
nand UO_1710 (O_1710,N_49831,N_49794);
or UO_1711 (O_1711,N_49841,N_49870);
and UO_1712 (O_1712,N_49848,N_49774);
nand UO_1713 (O_1713,N_49981,N_49918);
nor UO_1714 (O_1714,N_49790,N_49916);
nor UO_1715 (O_1715,N_49871,N_49975);
xor UO_1716 (O_1716,N_49944,N_49996);
or UO_1717 (O_1717,N_49889,N_49791);
nand UO_1718 (O_1718,N_49948,N_49800);
nor UO_1719 (O_1719,N_49864,N_49917);
or UO_1720 (O_1720,N_49889,N_49995);
and UO_1721 (O_1721,N_49798,N_49940);
nor UO_1722 (O_1722,N_49892,N_49912);
xnor UO_1723 (O_1723,N_49756,N_49852);
nor UO_1724 (O_1724,N_49751,N_49763);
nor UO_1725 (O_1725,N_49804,N_49820);
and UO_1726 (O_1726,N_49841,N_49861);
or UO_1727 (O_1727,N_49842,N_49860);
xnor UO_1728 (O_1728,N_49824,N_49846);
or UO_1729 (O_1729,N_49900,N_49787);
nand UO_1730 (O_1730,N_49791,N_49819);
nand UO_1731 (O_1731,N_49906,N_49805);
xor UO_1732 (O_1732,N_49866,N_49810);
and UO_1733 (O_1733,N_49983,N_49975);
nor UO_1734 (O_1734,N_49850,N_49806);
nor UO_1735 (O_1735,N_49923,N_49830);
or UO_1736 (O_1736,N_49991,N_49971);
nand UO_1737 (O_1737,N_49961,N_49759);
or UO_1738 (O_1738,N_49796,N_49877);
and UO_1739 (O_1739,N_49847,N_49830);
nand UO_1740 (O_1740,N_49932,N_49980);
nor UO_1741 (O_1741,N_49915,N_49807);
and UO_1742 (O_1742,N_49903,N_49772);
or UO_1743 (O_1743,N_49858,N_49989);
nor UO_1744 (O_1744,N_49808,N_49817);
and UO_1745 (O_1745,N_49801,N_49887);
or UO_1746 (O_1746,N_49752,N_49783);
nor UO_1747 (O_1747,N_49948,N_49928);
or UO_1748 (O_1748,N_49811,N_49982);
nand UO_1749 (O_1749,N_49788,N_49948);
nor UO_1750 (O_1750,N_49864,N_49814);
and UO_1751 (O_1751,N_49867,N_49823);
nand UO_1752 (O_1752,N_49832,N_49805);
and UO_1753 (O_1753,N_49871,N_49987);
nor UO_1754 (O_1754,N_49790,N_49760);
nor UO_1755 (O_1755,N_49784,N_49820);
nand UO_1756 (O_1756,N_49919,N_49781);
nand UO_1757 (O_1757,N_49802,N_49849);
and UO_1758 (O_1758,N_49883,N_49761);
nor UO_1759 (O_1759,N_49765,N_49879);
or UO_1760 (O_1760,N_49882,N_49810);
nand UO_1761 (O_1761,N_49875,N_49877);
or UO_1762 (O_1762,N_49943,N_49811);
nor UO_1763 (O_1763,N_49779,N_49865);
xnor UO_1764 (O_1764,N_49829,N_49988);
nand UO_1765 (O_1765,N_49970,N_49983);
nand UO_1766 (O_1766,N_49768,N_49980);
nor UO_1767 (O_1767,N_49918,N_49886);
or UO_1768 (O_1768,N_49833,N_49856);
or UO_1769 (O_1769,N_49888,N_49788);
and UO_1770 (O_1770,N_49798,N_49857);
nor UO_1771 (O_1771,N_49847,N_49849);
nor UO_1772 (O_1772,N_49874,N_49828);
xor UO_1773 (O_1773,N_49924,N_49877);
or UO_1774 (O_1774,N_49948,N_49908);
or UO_1775 (O_1775,N_49863,N_49792);
xnor UO_1776 (O_1776,N_49948,N_49856);
and UO_1777 (O_1777,N_49989,N_49810);
nor UO_1778 (O_1778,N_49851,N_49837);
xnor UO_1779 (O_1779,N_49755,N_49843);
nand UO_1780 (O_1780,N_49806,N_49856);
and UO_1781 (O_1781,N_49839,N_49889);
or UO_1782 (O_1782,N_49825,N_49945);
xor UO_1783 (O_1783,N_49865,N_49797);
and UO_1784 (O_1784,N_49941,N_49997);
or UO_1785 (O_1785,N_49856,N_49975);
and UO_1786 (O_1786,N_49875,N_49755);
or UO_1787 (O_1787,N_49982,N_49885);
nand UO_1788 (O_1788,N_49915,N_49922);
and UO_1789 (O_1789,N_49837,N_49820);
nand UO_1790 (O_1790,N_49911,N_49775);
or UO_1791 (O_1791,N_49834,N_49870);
nor UO_1792 (O_1792,N_49888,N_49918);
or UO_1793 (O_1793,N_49882,N_49833);
and UO_1794 (O_1794,N_49905,N_49823);
or UO_1795 (O_1795,N_49936,N_49777);
xnor UO_1796 (O_1796,N_49799,N_49989);
xor UO_1797 (O_1797,N_49796,N_49839);
xor UO_1798 (O_1798,N_49779,N_49836);
xor UO_1799 (O_1799,N_49828,N_49796);
nor UO_1800 (O_1800,N_49906,N_49840);
nand UO_1801 (O_1801,N_49992,N_49811);
nand UO_1802 (O_1802,N_49897,N_49863);
or UO_1803 (O_1803,N_49766,N_49939);
nand UO_1804 (O_1804,N_49978,N_49751);
nor UO_1805 (O_1805,N_49819,N_49775);
nand UO_1806 (O_1806,N_49947,N_49781);
nand UO_1807 (O_1807,N_49900,N_49760);
nor UO_1808 (O_1808,N_49958,N_49833);
and UO_1809 (O_1809,N_49828,N_49922);
nor UO_1810 (O_1810,N_49922,N_49762);
nand UO_1811 (O_1811,N_49865,N_49778);
and UO_1812 (O_1812,N_49806,N_49810);
or UO_1813 (O_1813,N_49949,N_49928);
nand UO_1814 (O_1814,N_49796,N_49770);
xor UO_1815 (O_1815,N_49976,N_49913);
or UO_1816 (O_1816,N_49923,N_49884);
nand UO_1817 (O_1817,N_49933,N_49941);
xnor UO_1818 (O_1818,N_49843,N_49974);
or UO_1819 (O_1819,N_49926,N_49822);
xor UO_1820 (O_1820,N_49908,N_49993);
xor UO_1821 (O_1821,N_49990,N_49829);
or UO_1822 (O_1822,N_49973,N_49984);
and UO_1823 (O_1823,N_49841,N_49758);
or UO_1824 (O_1824,N_49803,N_49798);
or UO_1825 (O_1825,N_49758,N_49986);
xor UO_1826 (O_1826,N_49876,N_49931);
xnor UO_1827 (O_1827,N_49811,N_49987);
and UO_1828 (O_1828,N_49756,N_49834);
and UO_1829 (O_1829,N_49975,N_49855);
nor UO_1830 (O_1830,N_49995,N_49860);
xor UO_1831 (O_1831,N_49983,N_49969);
xor UO_1832 (O_1832,N_49909,N_49878);
nor UO_1833 (O_1833,N_49974,N_49927);
nor UO_1834 (O_1834,N_49756,N_49938);
xor UO_1835 (O_1835,N_49915,N_49795);
xor UO_1836 (O_1836,N_49871,N_49867);
or UO_1837 (O_1837,N_49770,N_49966);
xor UO_1838 (O_1838,N_49778,N_49783);
nor UO_1839 (O_1839,N_49923,N_49919);
xor UO_1840 (O_1840,N_49769,N_49829);
and UO_1841 (O_1841,N_49763,N_49886);
or UO_1842 (O_1842,N_49988,N_49910);
or UO_1843 (O_1843,N_49774,N_49910);
and UO_1844 (O_1844,N_49967,N_49889);
and UO_1845 (O_1845,N_49996,N_49863);
and UO_1846 (O_1846,N_49789,N_49751);
nor UO_1847 (O_1847,N_49761,N_49871);
nor UO_1848 (O_1848,N_49859,N_49832);
and UO_1849 (O_1849,N_49861,N_49859);
or UO_1850 (O_1850,N_49829,N_49774);
or UO_1851 (O_1851,N_49801,N_49895);
nor UO_1852 (O_1852,N_49777,N_49752);
nand UO_1853 (O_1853,N_49812,N_49908);
nor UO_1854 (O_1854,N_49984,N_49961);
or UO_1855 (O_1855,N_49809,N_49832);
and UO_1856 (O_1856,N_49857,N_49794);
and UO_1857 (O_1857,N_49963,N_49757);
nand UO_1858 (O_1858,N_49788,N_49837);
nand UO_1859 (O_1859,N_49750,N_49774);
xnor UO_1860 (O_1860,N_49887,N_49867);
xor UO_1861 (O_1861,N_49794,N_49997);
or UO_1862 (O_1862,N_49894,N_49772);
and UO_1863 (O_1863,N_49967,N_49769);
xor UO_1864 (O_1864,N_49936,N_49929);
and UO_1865 (O_1865,N_49866,N_49909);
nand UO_1866 (O_1866,N_49987,N_49950);
nor UO_1867 (O_1867,N_49814,N_49950);
or UO_1868 (O_1868,N_49785,N_49908);
and UO_1869 (O_1869,N_49758,N_49855);
nand UO_1870 (O_1870,N_49950,N_49786);
xor UO_1871 (O_1871,N_49990,N_49967);
nor UO_1872 (O_1872,N_49942,N_49883);
or UO_1873 (O_1873,N_49874,N_49917);
and UO_1874 (O_1874,N_49958,N_49891);
nor UO_1875 (O_1875,N_49988,N_49924);
nor UO_1876 (O_1876,N_49807,N_49938);
or UO_1877 (O_1877,N_49762,N_49789);
or UO_1878 (O_1878,N_49870,N_49808);
and UO_1879 (O_1879,N_49892,N_49866);
or UO_1880 (O_1880,N_49845,N_49918);
xor UO_1881 (O_1881,N_49930,N_49938);
and UO_1882 (O_1882,N_49819,N_49956);
nand UO_1883 (O_1883,N_49994,N_49948);
xnor UO_1884 (O_1884,N_49888,N_49988);
xor UO_1885 (O_1885,N_49914,N_49930);
nor UO_1886 (O_1886,N_49827,N_49911);
and UO_1887 (O_1887,N_49792,N_49930);
nor UO_1888 (O_1888,N_49922,N_49930);
or UO_1889 (O_1889,N_49980,N_49786);
and UO_1890 (O_1890,N_49962,N_49757);
and UO_1891 (O_1891,N_49989,N_49809);
or UO_1892 (O_1892,N_49973,N_49972);
and UO_1893 (O_1893,N_49882,N_49938);
and UO_1894 (O_1894,N_49990,N_49780);
nand UO_1895 (O_1895,N_49891,N_49871);
or UO_1896 (O_1896,N_49767,N_49775);
or UO_1897 (O_1897,N_49844,N_49837);
nor UO_1898 (O_1898,N_49936,N_49877);
nand UO_1899 (O_1899,N_49896,N_49783);
or UO_1900 (O_1900,N_49969,N_49990);
and UO_1901 (O_1901,N_49849,N_49952);
xnor UO_1902 (O_1902,N_49949,N_49828);
nand UO_1903 (O_1903,N_49822,N_49835);
and UO_1904 (O_1904,N_49891,N_49750);
or UO_1905 (O_1905,N_49915,N_49873);
nor UO_1906 (O_1906,N_49827,N_49917);
nand UO_1907 (O_1907,N_49892,N_49819);
and UO_1908 (O_1908,N_49836,N_49810);
nor UO_1909 (O_1909,N_49921,N_49991);
nor UO_1910 (O_1910,N_49949,N_49954);
nand UO_1911 (O_1911,N_49872,N_49789);
xnor UO_1912 (O_1912,N_49962,N_49815);
and UO_1913 (O_1913,N_49898,N_49936);
nand UO_1914 (O_1914,N_49803,N_49773);
and UO_1915 (O_1915,N_49876,N_49885);
or UO_1916 (O_1916,N_49820,N_49956);
nand UO_1917 (O_1917,N_49920,N_49990);
xor UO_1918 (O_1918,N_49900,N_49757);
or UO_1919 (O_1919,N_49941,N_49934);
and UO_1920 (O_1920,N_49793,N_49985);
and UO_1921 (O_1921,N_49810,N_49756);
and UO_1922 (O_1922,N_49944,N_49806);
nor UO_1923 (O_1923,N_49967,N_49877);
nand UO_1924 (O_1924,N_49940,N_49951);
and UO_1925 (O_1925,N_49834,N_49961);
and UO_1926 (O_1926,N_49906,N_49917);
nor UO_1927 (O_1927,N_49947,N_49785);
xor UO_1928 (O_1928,N_49958,N_49969);
nor UO_1929 (O_1929,N_49985,N_49886);
nor UO_1930 (O_1930,N_49793,N_49900);
and UO_1931 (O_1931,N_49899,N_49871);
and UO_1932 (O_1932,N_49912,N_49948);
or UO_1933 (O_1933,N_49935,N_49892);
nand UO_1934 (O_1934,N_49758,N_49922);
xnor UO_1935 (O_1935,N_49778,N_49860);
nand UO_1936 (O_1936,N_49753,N_49818);
and UO_1937 (O_1937,N_49972,N_49884);
or UO_1938 (O_1938,N_49793,N_49878);
nor UO_1939 (O_1939,N_49877,N_49814);
nand UO_1940 (O_1940,N_49964,N_49759);
nand UO_1941 (O_1941,N_49949,N_49896);
nand UO_1942 (O_1942,N_49750,N_49872);
nor UO_1943 (O_1943,N_49917,N_49979);
xor UO_1944 (O_1944,N_49759,N_49776);
xor UO_1945 (O_1945,N_49806,N_49901);
nor UO_1946 (O_1946,N_49908,N_49902);
or UO_1947 (O_1947,N_49750,N_49760);
nand UO_1948 (O_1948,N_49998,N_49859);
xnor UO_1949 (O_1949,N_49843,N_49815);
or UO_1950 (O_1950,N_49967,N_49917);
and UO_1951 (O_1951,N_49836,N_49938);
xnor UO_1952 (O_1952,N_49776,N_49975);
nor UO_1953 (O_1953,N_49751,N_49774);
xnor UO_1954 (O_1954,N_49773,N_49840);
xnor UO_1955 (O_1955,N_49956,N_49843);
and UO_1956 (O_1956,N_49953,N_49996);
nor UO_1957 (O_1957,N_49760,N_49977);
nand UO_1958 (O_1958,N_49751,N_49786);
nand UO_1959 (O_1959,N_49866,N_49945);
nand UO_1960 (O_1960,N_49983,N_49995);
xnor UO_1961 (O_1961,N_49762,N_49770);
nand UO_1962 (O_1962,N_49943,N_49979);
and UO_1963 (O_1963,N_49803,N_49787);
nand UO_1964 (O_1964,N_49980,N_49797);
and UO_1965 (O_1965,N_49863,N_49753);
nand UO_1966 (O_1966,N_49922,N_49932);
xor UO_1967 (O_1967,N_49819,N_49795);
xnor UO_1968 (O_1968,N_49765,N_49848);
nand UO_1969 (O_1969,N_49768,N_49788);
or UO_1970 (O_1970,N_49857,N_49769);
nand UO_1971 (O_1971,N_49894,N_49842);
and UO_1972 (O_1972,N_49841,N_49890);
nand UO_1973 (O_1973,N_49929,N_49835);
nand UO_1974 (O_1974,N_49876,N_49957);
xor UO_1975 (O_1975,N_49802,N_49775);
xnor UO_1976 (O_1976,N_49836,N_49873);
nor UO_1977 (O_1977,N_49751,N_49929);
or UO_1978 (O_1978,N_49943,N_49818);
or UO_1979 (O_1979,N_49896,N_49962);
nor UO_1980 (O_1980,N_49931,N_49932);
or UO_1981 (O_1981,N_49950,N_49940);
nand UO_1982 (O_1982,N_49871,N_49971);
nor UO_1983 (O_1983,N_49798,N_49962);
or UO_1984 (O_1984,N_49996,N_49903);
xor UO_1985 (O_1985,N_49888,N_49897);
and UO_1986 (O_1986,N_49866,N_49776);
or UO_1987 (O_1987,N_49759,N_49854);
nand UO_1988 (O_1988,N_49984,N_49859);
xor UO_1989 (O_1989,N_49911,N_49761);
and UO_1990 (O_1990,N_49875,N_49788);
and UO_1991 (O_1991,N_49961,N_49842);
and UO_1992 (O_1992,N_49756,N_49905);
nand UO_1993 (O_1993,N_49867,N_49997);
and UO_1994 (O_1994,N_49994,N_49779);
xor UO_1995 (O_1995,N_49804,N_49805);
and UO_1996 (O_1996,N_49978,N_49827);
nand UO_1997 (O_1997,N_49791,N_49786);
xor UO_1998 (O_1998,N_49945,N_49797);
nor UO_1999 (O_1999,N_49841,N_49872);
or UO_2000 (O_2000,N_49919,N_49825);
xnor UO_2001 (O_2001,N_49875,N_49908);
nor UO_2002 (O_2002,N_49890,N_49789);
or UO_2003 (O_2003,N_49820,N_49862);
and UO_2004 (O_2004,N_49975,N_49891);
and UO_2005 (O_2005,N_49838,N_49875);
or UO_2006 (O_2006,N_49761,N_49832);
nand UO_2007 (O_2007,N_49854,N_49772);
xnor UO_2008 (O_2008,N_49884,N_49873);
and UO_2009 (O_2009,N_49768,N_49919);
and UO_2010 (O_2010,N_49985,N_49911);
or UO_2011 (O_2011,N_49936,N_49827);
nand UO_2012 (O_2012,N_49818,N_49812);
xnor UO_2013 (O_2013,N_49896,N_49963);
and UO_2014 (O_2014,N_49972,N_49909);
and UO_2015 (O_2015,N_49851,N_49861);
and UO_2016 (O_2016,N_49852,N_49899);
and UO_2017 (O_2017,N_49867,N_49868);
nor UO_2018 (O_2018,N_49764,N_49852);
nand UO_2019 (O_2019,N_49982,N_49765);
xor UO_2020 (O_2020,N_49904,N_49780);
nand UO_2021 (O_2021,N_49774,N_49960);
or UO_2022 (O_2022,N_49892,N_49847);
nor UO_2023 (O_2023,N_49854,N_49996);
nor UO_2024 (O_2024,N_49946,N_49787);
and UO_2025 (O_2025,N_49857,N_49768);
nor UO_2026 (O_2026,N_49880,N_49846);
or UO_2027 (O_2027,N_49917,N_49923);
or UO_2028 (O_2028,N_49843,N_49816);
and UO_2029 (O_2029,N_49858,N_49943);
or UO_2030 (O_2030,N_49882,N_49780);
and UO_2031 (O_2031,N_49935,N_49773);
xnor UO_2032 (O_2032,N_49906,N_49926);
xnor UO_2033 (O_2033,N_49777,N_49995);
or UO_2034 (O_2034,N_49990,N_49941);
xor UO_2035 (O_2035,N_49872,N_49820);
and UO_2036 (O_2036,N_49785,N_49892);
nor UO_2037 (O_2037,N_49932,N_49816);
nor UO_2038 (O_2038,N_49984,N_49972);
xnor UO_2039 (O_2039,N_49902,N_49992);
and UO_2040 (O_2040,N_49973,N_49864);
nor UO_2041 (O_2041,N_49856,N_49834);
or UO_2042 (O_2042,N_49951,N_49917);
or UO_2043 (O_2043,N_49982,N_49821);
or UO_2044 (O_2044,N_49754,N_49801);
or UO_2045 (O_2045,N_49807,N_49983);
or UO_2046 (O_2046,N_49988,N_49822);
nand UO_2047 (O_2047,N_49908,N_49934);
or UO_2048 (O_2048,N_49781,N_49802);
or UO_2049 (O_2049,N_49788,N_49964);
nor UO_2050 (O_2050,N_49966,N_49808);
and UO_2051 (O_2051,N_49922,N_49880);
or UO_2052 (O_2052,N_49979,N_49957);
nor UO_2053 (O_2053,N_49971,N_49779);
xnor UO_2054 (O_2054,N_49881,N_49886);
and UO_2055 (O_2055,N_49846,N_49955);
or UO_2056 (O_2056,N_49894,N_49934);
and UO_2057 (O_2057,N_49952,N_49781);
xor UO_2058 (O_2058,N_49997,N_49800);
and UO_2059 (O_2059,N_49948,N_49962);
and UO_2060 (O_2060,N_49998,N_49750);
nand UO_2061 (O_2061,N_49869,N_49763);
xnor UO_2062 (O_2062,N_49981,N_49924);
and UO_2063 (O_2063,N_49803,N_49829);
xor UO_2064 (O_2064,N_49880,N_49970);
nand UO_2065 (O_2065,N_49807,N_49880);
or UO_2066 (O_2066,N_49928,N_49837);
xor UO_2067 (O_2067,N_49916,N_49894);
and UO_2068 (O_2068,N_49768,N_49885);
and UO_2069 (O_2069,N_49819,N_49888);
xnor UO_2070 (O_2070,N_49913,N_49936);
or UO_2071 (O_2071,N_49880,N_49881);
or UO_2072 (O_2072,N_49764,N_49963);
or UO_2073 (O_2073,N_49843,N_49800);
nor UO_2074 (O_2074,N_49768,N_49798);
and UO_2075 (O_2075,N_49917,N_49992);
xnor UO_2076 (O_2076,N_49895,N_49919);
and UO_2077 (O_2077,N_49875,N_49797);
xor UO_2078 (O_2078,N_49980,N_49762);
or UO_2079 (O_2079,N_49871,N_49937);
or UO_2080 (O_2080,N_49842,N_49960);
xor UO_2081 (O_2081,N_49880,N_49787);
nor UO_2082 (O_2082,N_49926,N_49964);
nor UO_2083 (O_2083,N_49943,N_49930);
and UO_2084 (O_2084,N_49762,N_49769);
and UO_2085 (O_2085,N_49981,N_49897);
or UO_2086 (O_2086,N_49993,N_49764);
and UO_2087 (O_2087,N_49982,N_49774);
or UO_2088 (O_2088,N_49890,N_49950);
nand UO_2089 (O_2089,N_49969,N_49904);
xnor UO_2090 (O_2090,N_49850,N_49764);
and UO_2091 (O_2091,N_49938,N_49905);
xnor UO_2092 (O_2092,N_49898,N_49824);
nor UO_2093 (O_2093,N_49830,N_49929);
nor UO_2094 (O_2094,N_49874,N_49894);
or UO_2095 (O_2095,N_49798,N_49800);
nand UO_2096 (O_2096,N_49947,N_49821);
nand UO_2097 (O_2097,N_49884,N_49768);
nand UO_2098 (O_2098,N_49996,N_49800);
xor UO_2099 (O_2099,N_49979,N_49900);
xor UO_2100 (O_2100,N_49922,N_49920);
and UO_2101 (O_2101,N_49761,N_49844);
nor UO_2102 (O_2102,N_49939,N_49771);
nor UO_2103 (O_2103,N_49885,N_49920);
nor UO_2104 (O_2104,N_49802,N_49797);
and UO_2105 (O_2105,N_49880,N_49992);
nor UO_2106 (O_2106,N_49923,N_49753);
and UO_2107 (O_2107,N_49865,N_49817);
and UO_2108 (O_2108,N_49828,N_49973);
or UO_2109 (O_2109,N_49930,N_49928);
nand UO_2110 (O_2110,N_49752,N_49792);
xor UO_2111 (O_2111,N_49840,N_49805);
xor UO_2112 (O_2112,N_49780,N_49842);
nand UO_2113 (O_2113,N_49975,N_49809);
nor UO_2114 (O_2114,N_49975,N_49950);
nand UO_2115 (O_2115,N_49910,N_49838);
and UO_2116 (O_2116,N_49750,N_49805);
and UO_2117 (O_2117,N_49815,N_49989);
nand UO_2118 (O_2118,N_49761,N_49914);
or UO_2119 (O_2119,N_49821,N_49977);
and UO_2120 (O_2120,N_49912,N_49968);
nor UO_2121 (O_2121,N_49956,N_49869);
nor UO_2122 (O_2122,N_49877,N_49986);
or UO_2123 (O_2123,N_49794,N_49927);
or UO_2124 (O_2124,N_49842,N_49888);
nor UO_2125 (O_2125,N_49884,N_49802);
nand UO_2126 (O_2126,N_49847,N_49868);
xor UO_2127 (O_2127,N_49952,N_49983);
nor UO_2128 (O_2128,N_49883,N_49873);
and UO_2129 (O_2129,N_49847,N_49921);
nor UO_2130 (O_2130,N_49790,N_49793);
and UO_2131 (O_2131,N_49915,N_49832);
and UO_2132 (O_2132,N_49831,N_49863);
or UO_2133 (O_2133,N_49794,N_49757);
xor UO_2134 (O_2134,N_49873,N_49842);
or UO_2135 (O_2135,N_49898,N_49868);
and UO_2136 (O_2136,N_49969,N_49849);
or UO_2137 (O_2137,N_49812,N_49900);
nand UO_2138 (O_2138,N_49789,N_49780);
xnor UO_2139 (O_2139,N_49990,N_49783);
xor UO_2140 (O_2140,N_49765,N_49922);
and UO_2141 (O_2141,N_49900,N_49970);
xor UO_2142 (O_2142,N_49958,N_49809);
nor UO_2143 (O_2143,N_49757,N_49830);
or UO_2144 (O_2144,N_49753,N_49861);
or UO_2145 (O_2145,N_49778,N_49849);
nand UO_2146 (O_2146,N_49825,N_49785);
nand UO_2147 (O_2147,N_49962,N_49930);
xor UO_2148 (O_2148,N_49752,N_49825);
nand UO_2149 (O_2149,N_49871,N_49991);
xor UO_2150 (O_2150,N_49750,N_49944);
xor UO_2151 (O_2151,N_49767,N_49958);
nand UO_2152 (O_2152,N_49847,N_49950);
nor UO_2153 (O_2153,N_49824,N_49935);
and UO_2154 (O_2154,N_49844,N_49835);
and UO_2155 (O_2155,N_49793,N_49831);
nand UO_2156 (O_2156,N_49842,N_49852);
or UO_2157 (O_2157,N_49844,N_49812);
nand UO_2158 (O_2158,N_49842,N_49765);
or UO_2159 (O_2159,N_49815,N_49999);
xnor UO_2160 (O_2160,N_49886,N_49834);
and UO_2161 (O_2161,N_49983,N_49957);
nand UO_2162 (O_2162,N_49841,N_49892);
nand UO_2163 (O_2163,N_49796,N_49811);
xor UO_2164 (O_2164,N_49798,N_49888);
nor UO_2165 (O_2165,N_49984,N_49956);
or UO_2166 (O_2166,N_49909,N_49998);
or UO_2167 (O_2167,N_49809,N_49871);
nor UO_2168 (O_2168,N_49934,N_49856);
xor UO_2169 (O_2169,N_49951,N_49757);
and UO_2170 (O_2170,N_49834,N_49781);
and UO_2171 (O_2171,N_49971,N_49963);
or UO_2172 (O_2172,N_49838,N_49897);
nor UO_2173 (O_2173,N_49875,N_49870);
nor UO_2174 (O_2174,N_49893,N_49765);
xnor UO_2175 (O_2175,N_49811,N_49951);
xnor UO_2176 (O_2176,N_49970,N_49932);
and UO_2177 (O_2177,N_49763,N_49917);
xor UO_2178 (O_2178,N_49769,N_49845);
or UO_2179 (O_2179,N_49853,N_49772);
nand UO_2180 (O_2180,N_49898,N_49920);
xnor UO_2181 (O_2181,N_49929,N_49867);
nand UO_2182 (O_2182,N_49846,N_49753);
xnor UO_2183 (O_2183,N_49875,N_49770);
xnor UO_2184 (O_2184,N_49972,N_49780);
xnor UO_2185 (O_2185,N_49753,N_49987);
and UO_2186 (O_2186,N_49859,N_49906);
nor UO_2187 (O_2187,N_49864,N_49797);
or UO_2188 (O_2188,N_49848,N_49822);
nor UO_2189 (O_2189,N_49951,N_49999);
nor UO_2190 (O_2190,N_49836,N_49963);
or UO_2191 (O_2191,N_49859,N_49939);
and UO_2192 (O_2192,N_49842,N_49981);
nand UO_2193 (O_2193,N_49998,N_49860);
or UO_2194 (O_2194,N_49908,N_49925);
nor UO_2195 (O_2195,N_49882,N_49798);
nand UO_2196 (O_2196,N_49999,N_49824);
and UO_2197 (O_2197,N_49978,N_49774);
nand UO_2198 (O_2198,N_49855,N_49961);
xor UO_2199 (O_2199,N_49807,N_49968);
or UO_2200 (O_2200,N_49882,N_49971);
or UO_2201 (O_2201,N_49773,N_49811);
xnor UO_2202 (O_2202,N_49939,N_49884);
xnor UO_2203 (O_2203,N_49963,N_49954);
nand UO_2204 (O_2204,N_49884,N_49849);
and UO_2205 (O_2205,N_49938,N_49860);
xnor UO_2206 (O_2206,N_49942,N_49845);
or UO_2207 (O_2207,N_49984,N_49791);
nor UO_2208 (O_2208,N_49869,N_49990);
or UO_2209 (O_2209,N_49920,N_49929);
or UO_2210 (O_2210,N_49831,N_49925);
and UO_2211 (O_2211,N_49840,N_49985);
or UO_2212 (O_2212,N_49838,N_49881);
xor UO_2213 (O_2213,N_49821,N_49934);
and UO_2214 (O_2214,N_49958,N_49885);
or UO_2215 (O_2215,N_49811,N_49955);
and UO_2216 (O_2216,N_49834,N_49941);
nor UO_2217 (O_2217,N_49830,N_49871);
nand UO_2218 (O_2218,N_49979,N_49750);
nor UO_2219 (O_2219,N_49789,N_49917);
nand UO_2220 (O_2220,N_49958,N_49874);
or UO_2221 (O_2221,N_49859,N_49848);
xor UO_2222 (O_2222,N_49971,N_49935);
and UO_2223 (O_2223,N_49934,N_49970);
nor UO_2224 (O_2224,N_49845,N_49833);
nor UO_2225 (O_2225,N_49919,N_49898);
and UO_2226 (O_2226,N_49753,N_49980);
or UO_2227 (O_2227,N_49922,N_49846);
nor UO_2228 (O_2228,N_49943,N_49758);
and UO_2229 (O_2229,N_49771,N_49807);
or UO_2230 (O_2230,N_49782,N_49833);
or UO_2231 (O_2231,N_49880,N_49869);
nand UO_2232 (O_2232,N_49977,N_49810);
nor UO_2233 (O_2233,N_49911,N_49887);
nor UO_2234 (O_2234,N_49820,N_49890);
or UO_2235 (O_2235,N_49896,N_49950);
and UO_2236 (O_2236,N_49772,N_49986);
nand UO_2237 (O_2237,N_49792,N_49893);
nand UO_2238 (O_2238,N_49998,N_49753);
or UO_2239 (O_2239,N_49817,N_49869);
nand UO_2240 (O_2240,N_49872,N_49899);
xnor UO_2241 (O_2241,N_49945,N_49761);
or UO_2242 (O_2242,N_49844,N_49872);
and UO_2243 (O_2243,N_49850,N_49845);
or UO_2244 (O_2244,N_49823,N_49881);
and UO_2245 (O_2245,N_49958,N_49771);
xor UO_2246 (O_2246,N_49929,N_49905);
and UO_2247 (O_2247,N_49854,N_49790);
xnor UO_2248 (O_2248,N_49979,N_49885);
nand UO_2249 (O_2249,N_49878,N_49997);
xnor UO_2250 (O_2250,N_49986,N_49969);
or UO_2251 (O_2251,N_49920,N_49941);
or UO_2252 (O_2252,N_49871,N_49920);
nor UO_2253 (O_2253,N_49824,N_49889);
and UO_2254 (O_2254,N_49755,N_49892);
nor UO_2255 (O_2255,N_49913,N_49886);
or UO_2256 (O_2256,N_49799,N_49945);
and UO_2257 (O_2257,N_49847,N_49836);
or UO_2258 (O_2258,N_49770,N_49982);
nand UO_2259 (O_2259,N_49815,N_49928);
nor UO_2260 (O_2260,N_49753,N_49937);
or UO_2261 (O_2261,N_49843,N_49964);
or UO_2262 (O_2262,N_49769,N_49804);
nand UO_2263 (O_2263,N_49800,N_49778);
nand UO_2264 (O_2264,N_49792,N_49979);
or UO_2265 (O_2265,N_49808,N_49852);
or UO_2266 (O_2266,N_49802,N_49939);
xor UO_2267 (O_2267,N_49847,N_49851);
nand UO_2268 (O_2268,N_49794,N_49779);
and UO_2269 (O_2269,N_49794,N_49768);
or UO_2270 (O_2270,N_49847,N_49980);
and UO_2271 (O_2271,N_49847,N_49959);
nor UO_2272 (O_2272,N_49765,N_49945);
nand UO_2273 (O_2273,N_49821,N_49902);
nand UO_2274 (O_2274,N_49754,N_49968);
nor UO_2275 (O_2275,N_49758,N_49750);
nor UO_2276 (O_2276,N_49999,N_49806);
and UO_2277 (O_2277,N_49912,N_49866);
or UO_2278 (O_2278,N_49766,N_49894);
xnor UO_2279 (O_2279,N_49847,N_49856);
xor UO_2280 (O_2280,N_49793,N_49973);
nor UO_2281 (O_2281,N_49851,N_49880);
and UO_2282 (O_2282,N_49768,N_49985);
nand UO_2283 (O_2283,N_49835,N_49765);
nor UO_2284 (O_2284,N_49943,N_49934);
or UO_2285 (O_2285,N_49940,N_49814);
and UO_2286 (O_2286,N_49876,N_49831);
or UO_2287 (O_2287,N_49807,N_49824);
xnor UO_2288 (O_2288,N_49793,N_49883);
xor UO_2289 (O_2289,N_49896,N_49995);
nand UO_2290 (O_2290,N_49819,N_49773);
nand UO_2291 (O_2291,N_49757,N_49899);
nor UO_2292 (O_2292,N_49984,N_49989);
and UO_2293 (O_2293,N_49839,N_49843);
and UO_2294 (O_2294,N_49979,N_49831);
or UO_2295 (O_2295,N_49824,N_49760);
nand UO_2296 (O_2296,N_49896,N_49796);
nor UO_2297 (O_2297,N_49759,N_49827);
xor UO_2298 (O_2298,N_49763,N_49812);
nor UO_2299 (O_2299,N_49985,N_49808);
nand UO_2300 (O_2300,N_49956,N_49804);
xor UO_2301 (O_2301,N_49875,N_49796);
and UO_2302 (O_2302,N_49868,N_49873);
or UO_2303 (O_2303,N_49914,N_49982);
nor UO_2304 (O_2304,N_49926,N_49781);
nand UO_2305 (O_2305,N_49852,N_49871);
and UO_2306 (O_2306,N_49878,N_49991);
nand UO_2307 (O_2307,N_49884,N_49945);
and UO_2308 (O_2308,N_49924,N_49994);
xnor UO_2309 (O_2309,N_49995,N_49869);
and UO_2310 (O_2310,N_49769,N_49941);
nor UO_2311 (O_2311,N_49992,N_49907);
and UO_2312 (O_2312,N_49751,N_49955);
or UO_2313 (O_2313,N_49933,N_49944);
nand UO_2314 (O_2314,N_49835,N_49860);
xnor UO_2315 (O_2315,N_49752,N_49755);
and UO_2316 (O_2316,N_49998,N_49787);
nor UO_2317 (O_2317,N_49901,N_49765);
and UO_2318 (O_2318,N_49945,N_49987);
and UO_2319 (O_2319,N_49819,N_49832);
nor UO_2320 (O_2320,N_49791,N_49810);
nor UO_2321 (O_2321,N_49894,N_49812);
xnor UO_2322 (O_2322,N_49831,N_49859);
nor UO_2323 (O_2323,N_49811,N_49934);
xnor UO_2324 (O_2324,N_49840,N_49915);
xor UO_2325 (O_2325,N_49804,N_49762);
nor UO_2326 (O_2326,N_49807,N_49868);
or UO_2327 (O_2327,N_49930,N_49983);
and UO_2328 (O_2328,N_49957,N_49943);
and UO_2329 (O_2329,N_49981,N_49986);
nor UO_2330 (O_2330,N_49813,N_49904);
nand UO_2331 (O_2331,N_49775,N_49851);
nor UO_2332 (O_2332,N_49863,N_49947);
nor UO_2333 (O_2333,N_49925,N_49810);
xnor UO_2334 (O_2334,N_49994,N_49754);
xnor UO_2335 (O_2335,N_49982,N_49832);
nor UO_2336 (O_2336,N_49913,N_49901);
nor UO_2337 (O_2337,N_49845,N_49855);
nand UO_2338 (O_2338,N_49752,N_49804);
xnor UO_2339 (O_2339,N_49770,N_49785);
and UO_2340 (O_2340,N_49912,N_49973);
xor UO_2341 (O_2341,N_49920,N_49980);
nand UO_2342 (O_2342,N_49818,N_49841);
nor UO_2343 (O_2343,N_49791,N_49761);
or UO_2344 (O_2344,N_49775,N_49751);
and UO_2345 (O_2345,N_49931,N_49851);
or UO_2346 (O_2346,N_49994,N_49930);
nand UO_2347 (O_2347,N_49788,N_49882);
nor UO_2348 (O_2348,N_49992,N_49912);
or UO_2349 (O_2349,N_49790,N_49786);
and UO_2350 (O_2350,N_49846,N_49785);
or UO_2351 (O_2351,N_49867,N_49827);
nor UO_2352 (O_2352,N_49772,N_49887);
and UO_2353 (O_2353,N_49911,N_49819);
nand UO_2354 (O_2354,N_49781,N_49824);
nor UO_2355 (O_2355,N_49834,N_49765);
xnor UO_2356 (O_2356,N_49876,N_49896);
xnor UO_2357 (O_2357,N_49892,N_49933);
nor UO_2358 (O_2358,N_49755,N_49759);
xor UO_2359 (O_2359,N_49999,N_49943);
nor UO_2360 (O_2360,N_49985,N_49821);
or UO_2361 (O_2361,N_49797,N_49766);
xnor UO_2362 (O_2362,N_49756,N_49876);
nand UO_2363 (O_2363,N_49833,N_49984);
nor UO_2364 (O_2364,N_49857,N_49872);
or UO_2365 (O_2365,N_49855,N_49969);
nand UO_2366 (O_2366,N_49767,N_49973);
nand UO_2367 (O_2367,N_49791,N_49866);
and UO_2368 (O_2368,N_49922,N_49900);
or UO_2369 (O_2369,N_49830,N_49862);
or UO_2370 (O_2370,N_49771,N_49871);
and UO_2371 (O_2371,N_49809,N_49778);
xor UO_2372 (O_2372,N_49839,N_49850);
and UO_2373 (O_2373,N_49959,N_49980);
nor UO_2374 (O_2374,N_49765,N_49841);
or UO_2375 (O_2375,N_49961,N_49962);
and UO_2376 (O_2376,N_49959,N_49996);
or UO_2377 (O_2377,N_49912,N_49977);
xor UO_2378 (O_2378,N_49878,N_49920);
nor UO_2379 (O_2379,N_49817,N_49839);
nor UO_2380 (O_2380,N_49859,N_49902);
xnor UO_2381 (O_2381,N_49953,N_49892);
xnor UO_2382 (O_2382,N_49858,N_49949);
nand UO_2383 (O_2383,N_49869,N_49865);
xnor UO_2384 (O_2384,N_49976,N_49809);
xor UO_2385 (O_2385,N_49846,N_49923);
or UO_2386 (O_2386,N_49912,N_49931);
nor UO_2387 (O_2387,N_49860,N_49796);
xor UO_2388 (O_2388,N_49961,N_49870);
nand UO_2389 (O_2389,N_49898,N_49776);
xnor UO_2390 (O_2390,N_49824,N_49794);
nand UO_2391 (O_2391,N_49897,N_49837);
nor UO_2392 (O_2392,N_49897,N_49828);
nor UO_2393 (O_2393,N_49943,N_49769);
and UO_2394 (O_2394,N_49841,N_49875);
nand UO_2395 (O_2395,N_49830,N_49858);
xor UO_2396 (O_2396,N_49987,N_49952);
xor UO_2397 (O_2397,N_49787,N_49943);
nand UO_2398 (O_2398,N_49965,N_49840);
nor UO_2399 (O_2399,N_49993,N_49795);
nor UO_2400 (O_2400,N_49865,N_49918);
nand UO_2401 (O_2401,N_49958,N_49798);
nand UO_2402 (O_2402,N_49983,N_49765);
or UO_2403 (O_2403,N_49767,N_49957);
and UO_2404 (O_2404,N_49928,N_49805);
and UO_2405 (O_2405,N_49792,N_49758);
or UO_2406 (O_2406,N_49779,N_49998);
and UO_2407 (O_2407,N_49956,N_49944);
nand UO_2408 (O_2408,N_49913,N_49813);
nor UO_2409 (O_2409,N_49834,N_49868);
or UO_2410 (O_2410,N_49898,N_49903);
and UO_2411 (O_2411,N_49845,N_49819);
nor UO_2412 (O_2412,N_49786,N_49870);
or UO_2413 (O_2413,N_49792,N_49769);
or UO_2414 (O_2414,N_49760,N_49980);
and UO_2415 (O_2415,N_49871,N_49803);
nand UO_2416 (O_2416,N_49875,N_49778);
nand UO_2417 (O_2417,N_49887,N_49824);
nand UO_2418 (O_2418,N_49755,N_49779);
or UO_2419 (O_2419,N_49865,N_49958);
and UO_2420 (O_2420,N_49953,N_49769);
nor UO_2421 (O_2421,N_49839,N_49857);
xor UO_2422 (O_2422,N_49758,N_49926);
and UO_2423 (O_2423,N_49782,N_49812);
or UO_2424 (O_2424,N_49843,N_49826);
nand UO_2425 (O_2425,N_49950,N_49829);
and UO_2426 (O_2426,N_49815,N_49942);
or UO_2427 (O_2427,N_49849,N_49901);
or UO_2428 (O_2428,N_49947,N_49817);
xnor UO_2429 (O_2429,N_49789,N_49965);
nor UO_2430 (O_2430,N_49800,N_49783);
or UO_2431 (O_2431,N_49774,N_49972);
or UO_2432 (O_2432,N_49863,N_49812);
nand UO_2433 (O_2433,N_49833,N_49874);
xnor UO_2434 (O_2434,N_49895,N_49870);
or UO_2435 (O_2435,N_49975,N_49790);
xor UO_2436 (O_2436,N_49949,N_49762);
xnor UO_2437 (O_2437,N_49858,N_49874);
nand UO_2438 (O_2438,N_49827,N_49934);
or UO_2439 (O_2439,N_49983,N_49813);
xnor UO_2440 (O_2440,N_49912,N_49937);
and UO_2441 (O_2441,N_49827,N_49865);
xor UO_2442 (O_2442,N_49996,N_49754);
or UO_2443 (O_2443,N_49797,N_49806);
and UO_2444 (O_2444,N_49921,N_49831);
and UO_2445 (O_2445,N_49805,N_49790);
nand UO_2446 (O_2446,N_49933,N_49965);
and UO_2447 (O_2447,N_49846,N_49797);
nand UO_2448 (O_2448,N_49784,N_49752);
and UO_2449 (O_2449,N_49936,N_49921);
xnor UO_2450 (O_2450,N_49935,N_49889);
nor UO_2451 (O_2451,N_49853,N_49946);
nand UO_2452 (O_2452,N_49844,N_49942);
nand UO_2453 (O_2453,N_49859,N_49874);
or UO_2454 (O_2454,N_49785,N_49813);
and UO_2455 (O_2455,N_49848,N_49871);
or UO_2456 (O_2456,N_49765,N_49972);
xor UO_2457 (O_2457,N_49881,N_49759);
xnor UO_2458 (O_2458,N_49901,N_49900);
nand UO_2459 (O_2459,N_49756,N_49891);
nor UO_2460 (O_2460,N_49983,N_49792);
or UO_2461 (O_2461,N_49891,N_49936);
xnor UO_2462 (O_2462,N_49790,N_49802);
and UO_2463 (O_2463,N_49990,N_49832);
nor UO_2464 (O_2464,N_49859,N_49972);
xnor UO_2465 (O_2465,N_49895,N_49968);
nand UO_2466 (O_2466,N_49937,N_49752);
nand UO_2467 (O_2467,N_49779,N_49958);
xor UO_2468 (O_2468,N_49874,N_49895);
and UO_2469 (O_2469,N_49929,N_49971);
and UO_2470 (O_2470,N_49806,N_49786);
and UO_2471 (O_2471,N_49881,N_49841);
xor UO_2472 (O_2472,N_49967,N_49961);
nor UO_2473 (O_2473,N_49968,N_49988);
xor UO_2474 (O_2474,N_49822,N_49869);
nor UO_2475 (O_2475,N_49998,N_49870);
xnor UO_2476 (O_2476,N_49825,N_49922);
xor UO_2477 (O_2477,N_49780,N_49865);
and UO_2478 (O_2478,N_49803,N_49793);
nand UO_2479 (O_2479,N_49794,N_49883);
or UO_2480 (O_2480,N_49921,N_49796);
or UO_2481 (O_2481,N_49796,N_49923);
xor UO_2482 (O_2482,N_49864,N_49782);
or UO_2483 (O_2483,N_49805,N_49847);
nand UO_2484 (O_2484,N_49940,N_49990);
or UO_2485 (O_2485,N_49794,N_49861);
or UO_2486 (O_2486,N_49765,N_49851);
nor UO_2487 (O_2487,N_49876,N_49987);
xor UO_2488 (O_2488,N_49953,N_49775);
or UO_2489 (O_2489,N_49854,N_49983);
and UO_2490 (O_2490,N_49780,N_49874);
nor UO_2491 (O_2491,N_49805,N_49993);
xor UO_2492 (O_2492,N_49965,N_49763);
or UO_2493 (O_2493,N_49803,N_49940);
xor UO_2494 (O_2494,N_49974,N_49995);
and UO_2495 (O_2495,N_49999,N_49924);
and UO_2496 (O_2496,N_49872,N_49946);
xnor UO_2497 (O_2497,N_49923,N_49881);
and UO_2498 (O_2498,N_49809,N_49843);
or UO_2499 (O_2499,N_49994,N_49757);
nand UO_2500 (O_2500,N_49882,N_49915);
nor UO_2501 (O_2501,N_49952,N_49966);
nor UO_2502 (O_2502,N_49762,N_49846);
nor UO_2503 (O_2503,N_49801,N_49841);
nor UO_2504 (O_2504,N_49940,N_49945);
xor UO_2505 (O_2505,N_49980,N_49936);
xor UO_2506 (O_2506,N_49789,N_49946);
and UO_2507 (O_2507,N_49824,N_49871);
nor UO_2508 (O_2508,N_49991,N_49857);
and UO_2509 (O_2509,N_49789,N_49812);
nor UO_2510 (O_2510,N_49806,N_49994);
and UO_2511 (O_2511,N_49806,N_49865);
nand UO_2512 (O_2512,N_49942,N_49989);
or UO_2513 (O_2513,N_49813,N_49834);
or UO_2514 (O_2514,N_49939,N_49863);
xor UO_2515 (O_2515,N_49910,N_49935);
xor UO_2516 (O_2516,N_49939,N_49910);
nand UO_2517 (O_2517,N_49905,N_49776);
nand UO_2518 (O_2518,N_49879,N_49994);
nand UO_2519 (O_2519,N_49983,N_49881);
nand UO_2520 (O_2520,N_49933,N_49828);
or UO_2521 (O_2521,N_49812,N_49948);
and UO_2522 (O_2522,N_49954,N_49970);
nor UO_2523 (O_2523,N_49835,N_49934);
nor UO_2524 (O_2524,N_49789,N_49791);
and UO_2525 (O_2525,N_49770,N_49909);
nand UO_2526 (O_2526,N_49881,N_49928);
and UO_2527 (O_2527,N_49856,N_49783);
and UO_2528 (O_2528,N_49999,N_49757);
and UO_2529 (O_2529,N_49775,N_49871);
nor UO_2530 (O_2530,N_49937,N_49932);
or UO_2531 (O_2531,N_49931,N_49840);
or UO_2532 (O_2532,N_49970,N_49791);
and UO_2533 (O_2533,N_49980,N_49912);
xor UO_2534 (O_2534,N_49900,N_49861);
and UO_2535 (O_2535,N_49931,N_49783);
nand UO_2536 (O_2536,N_49813,N_49941);
and UO_2537 (O_2537,N_49971,N_49866);
nand UO_2538 (O_2538,N_49860,N_49966);
nand UO_2539 (O_2539,N_49756,N_49826);
and UO_2540 (O_2540,N_49840,N_49753);
nand UO_2541 (O_2541,N_49800,N_49893);
nor UO_2542 (O_2542,N_49878,N_49772);
or UO_2543 (O_2543,N_49810,N_49910);
nand UO_2544 (O_2544,N_49972,N_49757);
nor UO_2545 (O_2545,N_49899,N_49857);
or UO_2546 (O_2546,N_49837,N_49821);
nand UO_2547 (O_2547,N_49965,N_49782);
or UO_2548 (O_2548,N_49991,N_49868);
or UO_2549 (O_2549,N_49824,N_49870);
and UO_2550 (O_2550,N_49794,N_49998);
xnor UO_2551 (O_2551,N_49907,N_49892);
nor UO_2552 (O_2552,N_49814,N_49848);
or UO_2553 (O_2553,N_49962,N_49924);
and UO_2554 (O_2554,N_49826,N_49760);
or UO_2555 (O_2555,N_49803,N_49834);
xnor UO_2556 (O_2556,N_49750,N_49813);
xnor UO_2557 (O_2557,N_49972,N_49986);
or UO_2558 (O_2558,N_49985,N_49839);
nand UO_2559 (O_2559,N_49981,N_49846);
or UO_2560 (O_2560,N_49882,N_49935);
xnor UO_2561 (O_2561,N_49896,N_49984);
xnor UO_2562 (O_2562,N_49974,N_49889);
nand UO_2563 (O_2563,N_49948,N_49841);
xor UO_2564 (O_2564,N_49856,N_49946);
and UO_2565 (O_2565,N_49862,N_49848);
and UO_2566 (O_2566,N_49779,N_49868);
nor UO_2567 (O_2567,N_49805,N_49794);
nor UO_2568 (O_2568,N_49829,N_49879);
or UO_2569 (O_2569,N_49970,N_49816);
nor UO_2570 (O_2570,N_49998,N_49903);
and UO_2571 (O_2571,N_49964,N_49903);
nand UO_2572 (O_2572,N_49814,N_49769);
or UO_2573 (O_2573,N_49956,N_49870);
and UO_2574 (O_2574,N_49944,N_49758);
nor UO_2575 (O_2575,N_49954,N_49852);
nor UO_2576 (O_2576,N_49999,N_49991);
and UO_2577 (O_2577,N_49929,N_49856);
or UO_2578 (O_2578,N_49858,N_49904);
nor UO_2579 (O_2579,N_49991,N_49969);
nand UO_2580 (O_2580,N_49798,N_49988);
or UO_2581 (O_2581,N_49967,N_49887);
xor UO_2582 (O_2582,N_49988,N_49756);
or UO_2583 (O_2583,N_49792,N_49791);
nand UO_2584 (O_2584,N_49914,N_49788);
nor UO_2585 (O_2585,N_49930,N_49948);
and UO_2586 (O_2586,N_49952,N_49989);
and UO_2587 (O_2587,N_49967,N_49796);
nor UO_2588 (O_2588,N_49790,N_49897);
and UO_2589 (O_2589,N_49915,N_49923);
xor UO_2590 (O_2590,N_49997,N_49850);
and UO_2591 (O_2591,N_49883,N_49856);
nand UO_2592 (O_2592,N_49761,N_49807);
and UO_2593 (O_2593,N_49857,N_49984);
nor UO_2594 (O_2594,N_49975,N_49880);
xnor UO_2595 (O_2595,N_49853,N_49926);
nand UO_2596 (O_2596,N_49919,N_49887);
nand UO_2597 (O_2597,N_49926,N_49930);
nand UO_2598 (O_2598,N_49866,N_49838);
xnor UO_2599 (O_2599,N_49856,N_49859);
nand UO_2600 (O_2600,N_49751,N_49872);
or UO_2601 (O_2601,N_49862,N_49895);
and UO_2602 (O_2602,N_49947,N_49935);
xor UO_2603 (O_2603,N_49922,N_49952);
and UO_2604 (O_2604,N_49764,N_49833);
nand UO_2605 (O_2605,N_49852,N_49898);
nand UO_2606 (O_2606,N_49886,N_49940);
xor UO_2607 (O_2607,N_49864,N_49890);
nand UO_2608 (O_2608,N_49837,N_49754);
nand UO_2609 (O_2609,N_49949,N_49774);
xor UO_2610 (O_2610,N_49789,N_49861);
nand UO_2611 (O_2611,N_49834,N_49931);
xor UO_2612 (O_2612,N_49987,N_49782);
or UO_2613 (O_2613,N_49906,N_49971);
or UO_2614 (O_2614,N_49877,N_49881);
or UO_2615 (O_2615,N_49830,N_49846);
nor UO_2616 (O_2616,N_49784,N_49785);
and UO_2617 (O_2617,N_49772,N_49837);
xor UO_2618 (O_2618,N_49924,N_49934);
and UO_2619 (O_2619,N_49919,N_49793);
nor UO_2620 (O_2620,N_49880,N_49990);
or UO_2621 (O_2621,N_49849,N_49938);
xnor UO_2622 (O_2622,N_49950,N_49842);
nor UO_2623 (O_2623,N_49770,N_49995);
nand UO_2624 (O_2624,N_49959,N_49933);
nand UO_2625 (O_2625,N_49914,N_49935);
nand UO_2626 (O_2626,N_49887,N_49980);
nor UO_2627 (O_2627,N_49936,N_49897);
and UO_2628 (O_2628,N_49861,N_49850);
nor UO_2629 (O_2629,N_49985,N_49944);
nor UO_2630 (O_2630,N_49894,N_49960);
nand UO_2631 (O_2631,N_49920,N_49981);
nand UO_2632 (O_2632,N_49858,N_49805);
or UO_2633 (O_2633,N_49755,N_49932);
nand UO_2634 (O_2634,N_49833,N_49875);
and UO_2635 (O_2635,N_49868,N_49825);
nand UO_2636 (O_2636,N_49759,N_49892);
xor UO_2637 (O_2637,N_49995,N_49817);
nor UO_2638 (O_2638,N_49920,N_49761);
xnor UO_2639 (O_2639,N_49882,N_49843);
nor UO_2640 (O_2640,N_49817,N_49971);
and UO_2641 (O_2641,N_49854,N_49778);
nor UO_2642 (O_2642,N_49850,N_49938);
xnor UO_2643 (O_2643,N_49853,N_49763);
or UO_2644 (O_2644,N_49761,N_49904);
nor UO_2645 (O_2645,N_49809,N_49845);
and UO_2646 (O_2646,N_49817,N_49909);
or UO_2647 (O_2647,N_49808,N_49842);
nor UO_2648 (O_2648,N_49909,N_49913);
nand UO_2649 (O_2649,N_49860,N_49822);
nor UO_2650 (O_2650,N_49779,N_49922);
xor UO_2651 (O_2651,N_49750,N_49896);
nor UO_2652 (O_2652,N_49934,N_49984);
nand UO_2653 (O_2653,N_49790,N_49785);
and UO_2654 (O_2654,N_49919,N_49935);
nand UO_2655 (O_2655,N_49799,N_49825);
nor UO_2656 (O_2656,N_49915,N_49972);
and UO_2657 (O_2657,N_49890,N_49939);
nand UO_2658 (O_2658,N_49775,N_49993);
or UO_2659 (O_2659,N_49879,N_49874);
nand UO_2660 (O_2660,N_49814,N_49861);
nand UO_2661 (O_2661,N_49793,N_49954);
xor UO_2662 (O_2662,N_49941,N_49868);
or UO_2663 (O_2663,N_49979,N_49756);
xor UO_2664 (O_2664,N_49754,N_49865);
nor UO_2665 (O_2665,N_49979,N_49922);
or UO_2666 (O_2666,N_49815,N_49836);
or UO_2667 (O_2667,N_49763,N_49833);
and UO_2668 (O_2668,N_49876,N_49752);
or UO_2669 (O_2669,N_49954,N_49994);
nor UO_2670 (O_2670,N_49916,N_49930);
xor UO_2671 (O_2671,N_49961,N_49956);
and UO_2672 (O_2672,N_49929,N_49820);
or UO_2673 (O_2673,N_49846,N_49875);
nor UO_2674 (O_2674,N_49872,N_49942);
or UO_2675 (O_2675,N_49797,N_49761);
nor UO_2676 (O_2676,N_49920,N_49999);
xnor UO_2677 (O_2677,N_49764,N_49950);
or UO_2678 (O_2678,N_49933,N_49808);
nor UO_2679 (O_2679,N_49950,N_49959);
and UO_2680 (O_2680,N_49868,N_49793);
and UO_2681 (O_2681,N_49891,N_49977);
nor UO_2682 (O_2682,N_49928,N_49844);
and UO_2683 (O_2683,N_49995,N_49982);
nand UO_2684 (O_2684,N_49976,N_49937);
and UO_2685 (O_2685,N_49842,N_49861);
nor UO_2686 (O_2686,N_49804,N_49953);
nand UO_2687 (O_2687,N_49977,N_49805);
nor UO_2688 (O_2688,N_49988,N_49809);
or UO_2689 (O_2689,N_49775,N_49758);
and UO_2690 (O_2690,N_49835,N_49959);
xor UO_2691 (O_2691,N_49912,N_49945);
nor UO_2692 (O_2692,N_49860,N_49929);
and UO_2693 (O_2693,N_49779,N_49821);
nand UO_2694 (O_2694,N_49848,N_49885);
nor UO_2695 (O_2695,N_49903,N_49767);
or UO_2696 (O_2696,N_49935,N_49803);
and UO_2697 (O_2697,N_49756,N_49968);
nand UO_2698 (O_2698,N_49838,N_49879);
or UO_2699 (O_2699,N_49901,N_49979);
nand UO_2700 (O_2700,N_49851,N_49830);
and UO_2701 (O_2701,N_49980,N_49943);
xnor UO_2702 (O_2702,N_49820,N_49841);
nor UO_2703 (O_2703,N_49764,N_49945);
xnor UO_2704 (O_2704,N_49893,N_49916);
nor UO_2705 (O_2705,N_49864,N_49826);
nor UO_2706 (O_2706,N_49751,N_49945);
xor UO_2707 (O_2707,N_49786,N_49767);
and UO_2708 (O_2708,N_49993,N_49927);
or UO_2709 (O_2709,N_49963,N_49956);
nand UO_2710 (O_2710,N_49955,N_49903);
nand UO_2711 (O_2711,N_49818,N_49774);
nand UO_2712 (O_2712,N_49957,N_49984);
or UO_2713 (O_2713,N_49973,N_49894);
nand UO_2714 (O_2714,N_49849,N_49755);
nand UO_2715 (O_2715,N_49839,N_49879);
nand UO_2716 (O_2716,N_49970,N_49838);
and UO_2717 (O_2717,N_49774,N_49762);
and UO_2718 (O_2718,N_49860,N_49981);
xnor UO_2719 (O_2719,N_49850,N_49990);
xor UO_2720 (O_2720,N_49918,N_49808);
xnor UO_2721 (O_2721,N_49914,N_49937);
xor UO_2722 (O_2722,N_49762,N_49950);
or UO_2723 (O_2723,N_49778,N_49756);
xor UO_2724 (O_2724,N_49942,N_49781);
nand UO_2725 (O_2725,N_49983,N_49789);
xor UO_2726 (O_2726,N_49989,N_49897);
or UO_2727 (O_2727,N_49912,N_49909);
and UO_2728 (O_2728,N_49845,N_49992);
and UO_2729 (O_2729,N_49796,N_49814);
nand UO_2730 (O_2730,N_49756,N_49946);
nor UO_2731 (O_2731,N_49820,N_49899);
nand UO_2732 (O_2732,N_49828,N_49979);
nor UO_2733 (O_2733,N_49979,N_49793);
nor UO_2734 (O_2734,N_49821,N_49957);
nor UO_2735 (O_2735,N_49763,N_49786);
or UO_2736 (O_2736,N_49856,N_49919);
or UO_2737 (O_2737,N_49982,N_49891);
xnor UO_2738 (O_2738,N_49942,N_49778);
xnor UO_2739 (O_2739,N_49876,N_49765);
nor UO_2740 (O_2740,N_49771,N_49783);
xor UO_2741 (O_2741,N_49892,N_49885);
nand UO_2742 (O_2742,N_49931,N_49785);
xnor UO_2743 (O_2743,N_49815,N_49833);
xnor UO_2744 (O_2744,N_49937,N_49829);
and UO_2745 (O_2745,N_49965,N_49859);
nor UO_2746 (O_2746,N_49792,N_49783);
or UO_2747 (O_2747,N_49984,N_49967);
nand UO_2748 (O_2748,N_49983,N_49802);
xnor UO_2749 (O_2749,N_49967,N_49856);
nand UO_2750 (O_2750,N_49940,N_49883);
xor UO_2751 (O_2751,N_49824,N_49977);
nand UO_2752 (O_2752,N_49849,N_49837);
and UO_2753 (O_2753,N_49794,N_49802);
and UO_2754 (O_2754,N_49901,N_49995);
and UO_2755 (O_2755,N_49954,N_49784);
nand UO_2756 (O_2756,N_49919,N_49865);
or UO_2757 (O_2757,N_49767,N_49986);
and UO_2758 (O_2758,N_49992,N_49949);
or UO_2759 (O_2759,N_49893,N_49854);
and UO_2760 (O_2760,N_49888,N_49766);
and UO_2761 (O_2761,N_49896,N_49808);
nand UO_2762 (O_2762,N_49760,N_49895);
and UO_2763 (O_2763,N_49771,N_49876);
xor UO_2764 (O_2764,N_49982,N_49984);
nor UO_2765 (O_2765,N_49902,N_49869);
or UO_2766 (O_2766,N_49889,N_49964);
nor UO_2767 (O_2767,N_49876,N_49767);
nand UO_2768 (O_2768,N_49917,N_49810);
nor UO_2769 (O_2769,N_49796,N_49936);
nand UO_2770 (O_2770,N_49986,N_49777);
nor UO_2771 (O_2771,N_49938,N_49801);
xnor UO_2772 (O_2772,N_49998,N_49988);
xnor UO_2773 (O_2773,N_49781,N_49761);
or UO_2774 (O_2774,N_49817,N_49978);
nor UO_2775 (O_2775,N_49812,N_49793);
or UO_2776 (O_2776,N_49854,N_49856);
or UO_2777 (O_2777,N_49767,N_49854);
nor UO_2778 (O_2778,N_49932,N_49814);
nand UO_2779 (O_2779,N_49782,N_49770);
and UO_2780 (O_2780,N_49793,N_49995);
xor UO_2781 (O_2781,N_49809,N_49762);
xor UO_2782 (O_2782,N_49937,N_49919);
nand UO_2783 (O_2783,N_49806,N_49802);
and UO_2784 (O_2784,N_49960,N_49904);
nand UO_2785 (O_2785,N_49791,N_49936);
nand UO_2786 (O_2786,N_49878,N_49904);
and UO_2787 (O_2787,N_49790,N_49923);
xnor UO_2788 (O_2788,N_49756,N_49804);
nand UO_2789 (O_2789,N_49918,N_49776);
and UO_2790 (O_2790,N_49847,N_49962);
nand UO_2791 (O_2791,N_49912,N_49942);
and UO_2792 (O_2792,N_49809,N_49957);
nor UO_2793 (O_2793,N_49973,N_49831);
xor UO_2794 (O_2794,N_49848,N_49817);
and UO_2795 (O_2795,N_49940,N_49759);
nor UO_2796 (O_2796,N_49801,N_49897);
and UO_2797 (O_2797,N_49894,N_49773);
nand UO_2798 (O_2798,N_49804,N_49893);
nand UO_2799 (O_2799,N_49802,N_49750);
nor UO_2800 (O_2800,N_49807,N_49939);
or UO_2801 (O_2801,N_49808,N_49923);
and UO_2802 (O_2802,N_49805,N_49889);
or UO_2803 (O_2803,N_49831,N_49788);
xor UO_2804 (O_2804,N_49878,N_49757);
nand UO_2805 (O_2805,N_49853,N_49764);
nor UO_2806 (O_2806,N_49927,N_49981);
or UO_2807 (O_2807,N_49930,N_49978);
or UO_2808 (O_2808,N_49805,N_49828);
nand UO_2809 (O_2809,N_49863,N_49764);
nor UO_2810 (O_2810,N_49840,N_49760);
xnor UO_2811 (O_2811,N_49851,N_49941);
xnor UO_2812 (O_2812,N_49963,N_49868);
or UO_2813 (O_2813,N_49967,N_49846);
nand UO_2814 (O_2814,N_49918,N_49971);
and UO_2815 (O_2815,N_49862,N_49872);
nand UO_2816 (O_2816,N_49750,N_49885);
or UO_2817 (O_2817,N_49996,N_49841);
nor UO_2818 (O_2818,N_49983,N_49879);
and UO_2819 (O_2819,N_49991,N_49830);
xor UO_2820 (O_2820,N_49930,N_49781);
nand UO_2821 (O_2821,N_49756,N_49895);
and UO_2822 (O_2822,N_49805,N_49844);
nor UO_2823 (O_2823,N_49831,N_49953);
or UO_2824 (O_2824,N_49809,N_49999);
xor UO_2825 (O_2825,N_49949,N_49956);
xor UO_2826 (O_2826,N_49859,N_49868);
and UO_2827 (O_2827,N_49943,N_49895);
nand UO_2828 (O_2828,N_49880,N_49873);
xnor UO_2829 (O_2829,N_49942,N_49835);
nand UO_2830 (O_2830,N_49913,N_49795);
xor UO_2831 (O_2831,N_49920,N_49964);
or UO_2832 (O_2832,N_49864,N_49947);
or UO_2833 (O_2833,N_49928,N_49783);
nor UO_2834 (O_2834,N_49775,N_49982);
nor UO_2835 (O_2835,N_49834,N_49985);
nand UO_2836 (O_2836,N_49799,N_49900);
or UO_2837 (O_2837,N_49894,N_49922);
and UO_2838 (O_2838,N_49958,N_49852);
or UO_2839 (O_2839,N_49906,N_49867);
and UO_2840 (O_2840,N_49866,N_49860);
nand UO_2841 (O_2841,N_49908,N_49851);
xnor UO_2842 (O_2842,N_49960,N_49790);
nand UO_2843 (O_2843,N_49893,N_49820);
xnor UO_2844 (O_2844,N_49819,N_49920);
or UO_2845 (O_2845,N_49975,N_49906);
nand UO_2846 (O_2846,N_49773,N_49855);
nor UO_2847 (O_2847,N_49871,N_49808);
nor UO_2848 (O_2848,N_49900,N_49776);
and UO_2849 (O_2849,N_49900,N_49921);
or UO_2850 (O_2850,N_49966,N_49927);
and UO_2851 (O_2851,N_49969,N_49887);
and UO_2852 (O_2852,N_49802,N_49986);
nand UO_2853 (O_2853,N_49820,N_49934);
nor UO_2854 (O_2854,N_49965,N_49768);
or UO_2855 (O_2855,N_49991,N_49800);
or UO_2856 (O_2856,N_49802,N_49880);
xnor UO_2857 (O_2857,N_49889,N_49859);
nand UO_2858 (O_2858,N_49862,N_49785);
and UO_2859 (O_2859,N_49864,N_49799);
or UO_2860 (O_2860,N_49769,N_49788);
nor UO_2861 (O_2861,N_49805,N_49774);
and UO_2862 (O_2862,N_49897,N_49761);
nor UO_2863 (O_2863,N_49870,N_49799);
nand UO_2864 (O_2864,N_49783,N_49753);
or UO_2865 (O_2865,N_49952,N_49954);
and UO_2866 (O_2866,N_49860,N_49903);
or UO_2867 (O_2867,N_49827,N_49796);
nor UO_2868 (O_2868,N_49996,N_49910);
or UO_2869 (O_2869,N_49885,N_49822);
and UO_2870 (O_2870,N_49875,N_49787);
and UO_2871 (O_2871,N_49895,N_49950);
nor UO_2872 (O_2872,N_49946,N_49902);
and UO_2873 (O_2873,N_49993,N_49941);
or UO_2874 (O_2874,N_49853,N_49797);
and UO_2875 (O_2875,N_49827,N_49894);
or UO_2876 (O_2876,N_49884,N_49789);
nor UO_2877 (O_2877,N_49806,N_49958);
nor UO_2878 (O_2878,N_49883,N_49907);
nand UO_2879 (O_2879,N_49773,N_49862);
and UO_2880 (O_2880,N_49857,N_49986);
or UO_2881 (O_2881,N_49935,N_49860);
nand UO_2882 (O_2882,N_49780,N_49796);
nand UO_2883 (O_2883,N_49863,N_49941);
xnor UO_2884 (O_2884,N_49971,N_49821);
xnor UO_2885 (O_2885,N_49984,N_49911);
or UO_2886 (O_2886,N_49929,N_49825);
or UO_2887 (O_2887,N_49833,N_49805);
nor UO_2888 (O_2888,N_49956,N_49930);
xnor UO_2889 (O_2889,N_49957,N_49752);
xnor UO_2890 (O_2890,N_49760,N_49966);
nand UO_2891 (O_2891,N_49785,N_49776);
or UO_2892 (O_2892,N_49952,N_49900);
xnor UO_2893 (O_2893,N_49788,N_49970);
xor UO_2894 (O_2894,N_49978,N_49794);
and UO_2895 (O_2895,N_49824,N_49751);
xor UO_2896 (O_2896,N_49862,N_49859);
xor UO_2897 (O_2897,N_49841,N_49767);
nand UO_2898 (O_2898,N_49858,N_49838);
and UO_2899 (O_2899,N_49789,N_49883);
nor UO_2900 (O_2900,N_49893,N_49907);
xor UO_2901 (O_2901,N_49879,N_49978);
and UO_2902 (O_2902,N_49817,N_49891);
nor UO_2903 (O_2903,N_49856,N_49987);
xnor UO_2904 (O_2904,N_49808,N_49886);
and UO_2905 (O_2905,N_49946,N_49750);
or UO_2906 (O_2906,N_49961,N_49981);
xor UO_2907 (O_2907,N_49817,N_49819);
nand UO_2908 (O_2908,N_49890,N_49769);
and UO_2909 (O_2909,N_49988,N_49801);
nor UO_2910 (O_2910,N_49819,N_49790);
nor UO_2911 (O_2911,N_49903,N_49782);
nor UO_2912 (O_2912,N_49768,N_49854);
xnor UO_2913 (O_2913,N_49756,N_49978);
and UO_2914 (O_2914,N_49912,N_49955);
xor UO_2915 (O_2915,N_49903,N_49856);
or UO_2916 (O_2916,N_49843,N_49923);
nand UO_2917 (O_2917,N_49981,N_49937);
and UO_2918 (O_2918,N_49985,N_49758);
or UO_2919 (O_2919,N_49907,N_49924);
and UO_2920 (O_2920,N_49855,N_49926);
nor UO_2921 (O_2921,N_49756,N_49757);
xnor UO_2922 (O_2922,N_49849,N_49866);
and UO_2923 (O_2923,N_49992,N_49934);
or UO_2924 (O_2924,N_49884,N_49885);
nand UO_2925 (O_2925,N_49872,N_49759);
xnor UO_2926 (O_2926,N_49883,N_49835);
xor UO_2927 (O_2927,N_49902,N_49789);
xnor UO_2928 (O_2928,N_49909,N_49982);
nor UO_2929 (O_2929,N_49935,N_49826);
xor UO_2930 (O_2930,N_49996,N_49921);
nand UO_2931 (O_2931,N_49971,N_49756);
xnor UO_2932 (O_2932,N_49974,N_49985);
and UO_2933 (O_2933,N_49905,N_49794);
nor UO_2934 (O_2934,N_49939,N_49793);
and UO_2935 (O_2935,N_49826,N_49898);
xor UO_2936 (O_2936,N_49863,N_49809);
xor UO_2937 (O_2937,N_49927,N_49815);
nor UO_2938 (O_2938,N_49963,N_49878);
nand UO_2939 (O_2939,N_49836,N_49898);
and UO_2940 (O_2940,N_49826,N_49949);
and UO_2941 (O_2941,N_49780,N_49885);
and UO_2942 (O_2942,N_49873,N_49865);
and UO_2943 (O_2943,N_49906,N_49757);
nor UO_2944 (O_2944,N_49875,N_49999);
nor UO_2945 (O_2945,N_49869,N_49821);
or UO_2946 (O_2946,N_49870,N_49892);
nand UO_2947 (O_2947,N_49867,N_49830);
nand UO_2948 (O_2948,N_49897,N_49809);
and UO_2949 (O_2949,N_49966,N_49829);
xnor UO_2950 (O_2950,N_49905,N_49958);
or UO_2951 (O_2951,N_49898,N_49750);
or UO_2952 (O_2952,N_49898,N_49833);
nor UO_2953 (O_2953,N_49780,N_49896);
xor UO_2954 (O_2954,N_49755,N_49805);
xor UO_2955 (O_2955,N_49965,N_49757);
and UO_2956 (O_2956,N_49898,N_49999);
nor UO_2957 (O_2957,N_49868,N_49977);
xnor UO_2958 (O_2958,N_49833,N_49993);
or UO_2959 (O_2959,N_49939,N_49761);
and UO_2960 (O_2960,N_49819,N_49924);
and UO_2961 (O_2961,N_49813,N_49789);
or UO_2962 (O_2962,N_49781,N_49893);
and UO_2963 (O_2963,N_49967,N_49763);
xnor UO_2964 (O_2964,N_49976,N_49961);
and UO_2965 (O_2965,N_49807,N_49987);
or UO_2966 (O_2966,N_49888,N_49980);
and UO_2967 (O_2967,N_49870,N_49885);
and UO_2968 (O_2968,N_49926,N_49978);
xnor UO_2969 (O_2969,N_49989,N_49785);
or UO_2970 (O_2970,N_49839,N_49905);
nand UO_2971 (O_2971,N_49779,N_49992);
xor UO_2972 (O_2972,N_49816,N_49878);
or UO_2973 (O_2973,N_49926,N_49839);
xnor UO_2974 (O_2974,N_49988,N_49790);
and UO_2975 (O_2975,N_49770,N_49881);
or UO_2976 (O_2976,N_49777,N_49762);
or UO_2977 (O_2977,N_49965,N_49780);
xor UO_2978 (O_2978,N_49993,N_49940);
or UO_2979 (O_2979,N_49945,N_49827);
or UO_2980 (O_2980,N_49751,N_49904);
nand UO_2981 (O_2981,N_49899,N_49794);
xnor UO_2982 (O_2982,N_49811,N_49912);
nor UO_2983 (O_2983,N_49810,N_49856);
nor UO_2984 (O_2984,N_49772,N_49822);
or UO_2985 (O_2985,N_49891,N_49863);
nand UO_2986 (O_2986,N_49866,N_49931);
nand UO_2987 (O_2987,N_49790,N_49797);
xnor UO_2988 (O_2988,N_49777,N_49850);
nor UO_2989 (O_2989,N_49779,N_49853);
nor UO_2990 (O_2990,N_49952,N_49820);
and UO_2991 (O_2991,N_49885,N_49965);
and UO_2992 (O_2992,N_49845,N_49852);
nor UO_2993 (O_2993,N_49859,N_49813);
xor UO_2994 (O_2994,N_49999,N_49964);
and UO_2995 (O_2995,N_49750,N_49869);
xor UO_2996 (O_2996,N_49985,N_49903);
xor UO_2997 (O_2997,N_49822,N_49924);
or UO_2998 (O_2998,N_49952,N_49930);
xnor UO_2999 (O_2999,N_49788,N_49868);
and UO_3000 (O_3000,N_49995,N_49936);
or UO_3001 (O_3001,N_49850,N_49759);
nand UO_3002 (O_3002,N_49810,N_49804);
nand UO_3003 (O_3003,N_49947,N_49875);
xor UO_3004 (O_3004,N_49936,N_49869);
xor UO_3005 (O_3005,N_49833,N_49775);
or UO_3006 (O_3006,N_49779,N_49856);
nor UO_3007 (O_3007,N_49787,N_49818);
or UO_3008 (O_3008,N_49840,N_49759);
nand UO_3009 (O_3009,N_49889,N_49794);
and UO_3010 (O_3010,N_49976,N_49890);
nand UO_3011 (O_3011,N_49824,N_49991);
or UO_3012 (O_3012,N_49838,N_49856);
nand UO_3013 (O_3013,N_49962,N_49766);
nand UO_3014 (O_3014,N_49923,N_49926);
nor UO_3015 (O_3015,N_49873,N_49762);
nand UO_3016 (O_3016,N_49919,N_49771);
and UO_3017 (O_3017,N_49908,N_49842);
and UO_3018 (O_3018,N_49880,N_49848);
or UO_3019 (O_3019,N_49751,N_49856);
and UO_3020 (O_3020,N_49753,N_49751);
or UO_3021 (O_3021,N_49949,N_49979);
and UO_3022 (O_3022,N_49885,N_49799);
and UO_3023 (O_3023,N_49965,N_49913);
or UO_3024 (O_3024,N_49782,N_49976);
xnor UO_3025 (O_3025,N_49911,N_49922);
or UO_3026 (O_3026,N_49980,N_49945);
and UO_3027 (O_3027,N_49954,N_49843);
or UO_3028 (O_3028,N_49818,N_49816);
nor UO_3029 (O_3029,N_49833,N_49966);
nand UO_3030 (O_3030,N_49872,N_49943);
and UO_3031 (O_3031,N_49784,N_49835);
and UO_3032 (O_3032,N_49912,N_49933);
xor UO_3033 (O_3033,N_49953,N_49891);
xnor UO_3034 (O_3034,N_49896,N_49763);
nor UO_3035 (O_3035,N_49753,N_49791);
xor UO_3036 (O_3036,N_49927,N_49999);
and UO_3037 (O_3037,N_49751,N_49887);
nand UO_3038 (O_3038,N_49918,N_49938);
and UO_3039 (O_3039,N_49980,N_49859);
xnor UO_3040 (O_3040,N_49905,N_49925);
and UO_3041 (O_3041,N_49803,N_49992);
or UO_3042 (O_3042,N_49900,N_49961);
and UO_3043 (O_3043,N_49921,N_49912);
xor UO_3044 (O_3044,N_49797,N_49934);
and UO_3045 (O_3045,N_49798,N_49967);
or UO_3046 (O_3046,N_49769,N_49821);
xor UO_3047 (O_3047,N_49872,N_49963);
and UO_3048 (O_3048,N_49771,N_49941);
and UO_3049 (O_3049,N_49956,N_49905);
xnor UO_3050 (O_3050,N_49839,N_49820);
nor UO_3051 (O_3051,N_49861,N_49766);
xor UO_3052 (O_3052,N_49984,N_49766);
xnor UO_3053 (O_3053,N_49844,N_49943);
xnor UO_3054 (O_3054,N_49952,N_49853);
or UO_3055 (O_3055,N_49760,N_49961);
nor UO_3056 (O_3056,N_49827,N_49823);
xor UO_3057 (O_3057,N_49833,N_49988);
xnor UO_3058 (O_3058,N_49754,N_49960);
nor UO_3059 (O_3059,N_49939,N_49930);
or UO_3060 (O_3060,N_49764,N_49755);
and UO_3061 (O_3061,N_49896,N_49789);
nor UO_3062 (O_3062,N_49936,N_49774);
nor UO_3063 (O_3063,N_49974,N_49820);
nor UO_3064 (O_3064,N_49810,N_49900);
or UO_3065 (O_3065,N_49934,N_49832);
nor UO_3066 (O_3066,N_49955,N_49895);
and UO_3067 (O_3067,N_49909,N_49897);
nand UO_3068 (O_3068,N_49797,N_49750);
nand UO_3069 (O_3069,N_49921,N_49897);
or UO_3070 (O_3070,N_49957,N_49866);
xnor UO_3071 (O_3071,N_49814,N_49908);
xnor UO_3072 (O_3072,N_49919,N_49788);
nand UO_3073 (O_3073,N_49831,N_49862);
xnor UO_3074 (O_3074,N_49809,N_49984);
and UO_3075 (O_3075,N_49917,N_49950);
or UO_3076 (O_3076,N_49829,N_49943);
xnor UO_3077 (O_3077,N_49757,N_49881);
or UO_3078 (O_3078,N_49954,N_49797);
nand UO_3079 (O_3079,N_49928,N_49966);
and UO_3080 (O_3080,N_49922,N_49999);
nand UO_3081 (O_3081,N_49956,N_49987);
xnor UO_3082 (O_3082,N_49964,N_49813);
nand UO_3083 (O_3083,N_49860,N_49812);
or UO_3084 (O_3084,N_49872,N_49945);
nand UO_3085 (O_3085,N_49926,N_49877);
xor UO_3086 (O_3086,N_49990,N_49751);
nor UO_3087 (O_3087,N_49887,N_49845);
and UO_3088 (O_3088,N_49941,N_49983);
and UO_3089 (O_3089,N_49999,N_49817);
xnor UO_3090 (O_3090,N_49829,N_49883);
or UO_3091 (O_3091,N_49752,N_49813);
nand UO_3092 (O_3092,N_49848,N_49879);
nand UO_3093 (O_3093,N_49792,N_49955);
or UO_3094 (O_3094,N_49825,N_49820);
nand UO_3095 (O_3095,N_49889,N_49767);
nor UO_3096 (O_3096,N_49765,N_49990);
or UO_3097 (O_3097,N_49990,N_49801);
nand UO_3098 (O_3098,N_49797,N_49778);
and UO_3099 (O_3099,N_49881,N_49780);
or UO_3100 (O_3100,N_49981,N_49845);
xor UO_3101 (O_3101,N_49980,N_49884);
or UO_3102 (O_3102,N_49775,N_49755);
nor UO_3103 (O_3103,N_49972,N_49818);
nand UO_3104 (O_3104,N_49933,N_49940);
xor UO_3105 (O_3105,N_49985,N_49951);
nand UO_3106 (O_3106,N_49846,N_49771);
nand UO_3107 (O_3107,N_49999,N_49849);
and UO_3108 (O_3108,N_49951,N_49937);
and UO_3109 (O_3109,N_49948,N_49964);
nand UO_3110 (O_3110,N_49773,N_49971);
and UO_3111 (O_3111,N_49985,N_49770);
nand UO_3112 (O_3112,N_49977,N_49973);
nand UO_3113 (O_3113,N_49759,N_49899);
nor UO_3114 (O_3114,N_49865,N_49926);
nand UO_3115 (O_3115,N_49825,N_49859);
xor UO_3116 (O_3116,N_49807,N_49806);
nor UO_3117 (O_3117,N_49929,N_49941);
or UO_3118 (O_3118,N_49914,N_49817);
nor UO_3119 (O_3119,N_49803,N_49960);
xor UO_3120 (O_3120,N_49965,N_49788);
nor UO_3121 (O_3121,N_49868,N_49761);
nor UO_3122 (O_3122,N_49790,N_49895);
or UO_3123 (O_3123,N_49759,N_49944);
xor UO_3124 (O_3124,N_49908,N_49959);
and UO_3125 (O_3125,N_49960,N_49899);
nand UO_3126 (O_3126,N_49915,N_49910);
and UO_3127 (O_3127,N_49752,N_49840);
nor UO_3128 (O_3128,N_49754,N_49836);
xor UO_3129 (O_3129,N_49764,N_49836);
or UO_3130 (O_3130,N_49827,N_49931);
or UO_3131 (O_3131,N_49760,N_49844);
nor UO_3132 (O_3132,N_49836,N_49775);
or UO_3133 (O_3133,N_49799,N_49821);
nor UO_3134 (O_3134,N_49962,N_49904);
nor UO_3135 (O_3135,N_49995,N_49997);
nor UO_3136 (O_3136,N_49954,N_49871);
and UO_3137 (O_3137,N_49911,N_49813);
nand UO_3138 (O_3138,N_49819,N_49982);
nor UO_3139 (O_3139,N_49773,N_49750);
and UO_3140 (O_3140,N_49995,N_49824);
or UO_3141 (O_3141,N_49795,N_49952);
nor UO_3142 (O_3142,N_49967,N_49794);
nand UO_3143 (O_3143,N_49849,N_49821);
nor UO_3144 (O_3144,N_49757,N_49777);
or UO_3145 (O_3145,N_49849,N_49772);
and UO_3146 (O_3146,N_49835,N_49876);
nand UO_3147 (O_3147,N_49933,N_49805);
xor UO_3148 (O_3148,N_49902,N_49915);
and UO_3149 (O_3149,N_49913,N_49894);
nand UO_3150 (O_3150,N_49761,N_49943);
nor UO_3151 (O_3151,N_49995,N_49847);
nand UO_3152 (O_3152,N_49804,N_49883);
or UO_3153 (O_3153,N_49846,N_49929);
or UO_3154 (O_3154,N_49858,N_49834);
and UO_3155 (O_3155,N_49759,N_49879);
xnor UO_3156 (O_3156,N_49919,N_49801);
and UO_3157 (O_3157,N_49763,N_49858);
xor UO_3158 (O_3158,N_49993,N_49818);
xnor UO_3159 (O_3159,N_49810,N_49797);
and UO_3160 (O_3160,N_49985,N_49881);
and UO_3161 (O_3161,N_49819,N_49882);
and UO_3162 (O_3162,N_49818,N_49861);
nand UO_3163 (O_3163,N_49921,N_49955);
nor UO_3164 (O_3164,N_49993,N_49753);
nand UO_3165 (O_3165,N_49862,N_49832);
nor UO_3166 (O_3166,N_49852,N_49795);
and UO_3167 (O_3167,N_49833,N_49812);
nor UO_3168 (O_3168,N_49823,N_49788);
or UO_3169 (O_3169,N_49889,N_49989);
xnor UO_3170 (O_3170,N_49890,N_49914);
xor UO_3171 (O_3171,N_49898,N_49817);
nor UO_3172 (O_3172,N_49773,N_49956);
nand UO_3173 (O_3173,N_49766,N_49937);
or UO_3174 (O_3174,N_49794,N_49894);
or UO_3175 (O_3175,N_49772,N_49950);
and UO_3176 (O_3176,N_49954,N_49881);
xor UO_3177 (O_3177,N_49993,N_49910);
nor UO_3178 (O_3178,N_49836,N_49900);
and UO_3179 (O_3179,N_49788,N_49979);
or UO_3180 (O_3180,N_49756,N_49755);
nor UO_3181 (O_3181,N_49967,N_49775);
xor UO_3182 (O_3182,N_49843,N_49838);
nor UO_3183 (O_3183,N_49895,N_49887);
nand UO_3184 (O_3184,N_49998,N_49971);
and UO_3185 (O_3185,N_49861,N_49770);
and UO_3186 (O_3186,N_49896,N_49934);
xnor UO_3187 (O_3187,N_49816,N_49952);
nand UO_3188 (O_3188,N_49878,N_49755);
nor UO_3189 (O_3189,N_49786,N_49756);
nor UO_3190 (O_3190,N_49856,N_49824);
nand UO_3191 (O_3191,N_49816,N_49770);
nor UO_3192 (O_3192,N_49833,N_49868);
nand UO_3193 (O_3193,N_49803,N_49867);
xnor UO_3194 (O_3194,N_49918,N_49827);
or UO_3195 (O_3195,N_49815,N_49897);
xor UO_3196 (O_3196,N_49923,N_49961);
or UO_3197 (O_3197,N_49989,N_49885);
and UO_3198 (O_3198,N_49961,N_49959);
xnor UO_3199 (O_3199,N_49883,N_49852);
nand UO_3200 (O_3200,N_49997,N_49795);
or UO_3201 (O_3201,N_49775,N_49827);
nor UO_3202 (O_3202,N_49773,N_49832);
xnor UO_3203 (O_3203,N_49873,N_49935);
nor UO_3204 (O_3204,N_49851,N_49789);
and UO_3205 (O_3205,N_49752,N_49809);
or UO_3206 (O_3206,N_49973,N_49845);
nor UO_3207 (O_3207,N_49774,N_49929);
nor UO_3208 (O_3208,N_49784,N_49875);
and UO_3209 (O_3209,N_49914,N_49950);
or UO_3210 (O_3210,N_49901,N_49814);
nand UO_3211 (O_3211,N_49883,N_49969);
nand UO_3212 (O_3212,N_49787,N_49906);
xor UO_3213 (O_3213,N_49967,N_49878);
nand UO_3214 (O_3214,N_49997,N_49804);
or UO_3215 (O_3215,N_49879,N_49886);
xnor UO_3216 (O_3216,N_49775,N_49864);
and UO_3217 (O_3217,N_49790,N_49953);
or UO_3218 (O_3218,N_49995,N_49996);
nand UO_3219 (O_3219,N_49990,N_49788);
xnor UO_3220 (O_3220,N_49906,N_49848);
and UO_3221 (O_3221,N_49810,N_49782);
or UO_3222 (O_3222,N_49812,N_49790);
nand UO_3223 (O_3223,N_49756,N_49912);
xor UO_3224 (O_3224,N_49770,N_49802);
nor UO_3225 (O_3225,N_49952,N_49892);
xnor UO_3226 (O_3226,N_49799,N_49850);
or UO_3227 (O_3227,N_49868,N_49943);
and UO_3228 (O_3228,N_49911,N_49872);
and UO_3229 (O_3229,N_49803,N_49989);
and UO_3230 (O_3230,N_49843,N_49926);
xor UO_3231 (O_3231,N_49968,N_49964);
xnor UO_3232 (O_3232,N_49884,N_49767);
nand UO_3233 (O_3233,N_49999,N_49751);
and UO_3234 (O_3234,N_49810,N_49787);
and UO_3235 (O_3235,N_49944,N_49852);
nand UO_3236 (O_3236,N_49874,N_49916);
nand UO_3237 (O_3237,N_49769,N_49915);
or UO_3238 (O_3238,N_49853,N_49895);
or UO_3239 (O_3239,N_49859,N_49880);
and UO_3240 (O_3240,N_49823,N_49964);
xnor UO_3241 (O_3241,N_49765,N_49943);
and UO_3242 (O_3242,N_49884,N_49808);
nor UO_3243 (O_3243,N_49916,N_49828);
xnor UO_3244 (O_3244,N_49762,N_49848);
and UO_3245 (O_3245,N_49987,N_49779);
and UO_3246 (O_3246,N_49818,N_49874);
nand UO_3247 (O_3247,N_49753,N_49807);
nor UO_3248 (O_3248,N_49821,N_49930);
nor UO_3249 (O_3249,N_49991,N_49793);
nor UO_3250 (O_3250,N_49796,N_49788);
and UO_3251 (O_3251,N_49845,N_49955);
xor UO_3252 (O_3252,N_49882,N_49948);
xor UO_3253 (O_3253,N_49940,N_49895);
and UO_3254 (O_3254,N_49783,N_49897);
or UO_3255 (O_3255,N_49972,N_49990);
nor UO_3256 (O_3256,N_49888,N_49783);
or UO_3257 (O_3257,N_49942,N_49967);
xor UO_3258 (O_3258,N_49964,N_49919);
nand UO_3259 (O_3259,N_49759,N_49806);
xnor UO_3260 (O_3260,N_49755,N_49823);
xnor UO_3261 (O_3261,N_49971,N_49878);
or UO_3262 (O_3262,N_49956,N_49840);
xnor UO_3263 (O_3263,N_49838,N_49828);
and UO_3264 (O_3264,N_49833,N_49781);
and UO_3265 (O_3265,N_49862,N_49779);
xnor UO_3266 (O_3266,N_49846,N_49971);
nand UO_3267 (O_3267,N_49891,N_49937);
and UO_3268 (O_3268,N_49793,N_49761);
and UO_3269 (O_3269,N_49859,N_49929);
xor UO_3270 (O_3270,N_49941,N_49906);
nand UO_3271 (O_3271,N_49973,N_49990);
nand UO_3272 (O_3272,N_49988,N_49825);
and UO_3273 (O_3273,N_49800,N_49822);
nor UO_3274 (O_3274,N_49903,N_49997);
nand UO_3275 (O_3275,N_49841,N_49756);
and UO_3276 (O_3276,N_49891,N_49847);
or UO_3277 (O_3277,N_49898,N_49791);
or UO_3278 (O_3278,N_49801,N_49959);
and UO_3279 (O_3279,N_49906,N_49771);
and UO_3280 (O_3280,N_49766,N_49886);
or UO_3281 (O_3281,N_49896,N_49766);
nor UO_3282 (O_3282,N_49777,N_49942);
nor UO_3283 (O_3283,N_49984,N_49917);
and UO_3284 (O_3284,N_49981,N_49941);
and UO_3285 (O_3285,N_49781,N_49803);
nand UO_3286 (O_3286,N_49803,N_49842);
xor UO_3287 (O_3287,N_49824,N_49786);
xor UO_3288 (O_3288,N_49868,N_49969);
or UO_3289 (O_3289,N_49761,N_49760);
nand UO_3290 (O_3290,N_49929,N_49838);
nor UO_3291 (O_3291,N_49985,N_49822);
nand UO_3292 (O_3292,N_49892,N_49778);
or UO_3293 (O_3293,N_49995,N_49864);
and UO_3294 (O_3294,N_49844,N_49788);
xor UO_3295 (O_3295,N_49928,N_49942);
xor UO_3296 (O_3296,N_49848,N_49895);
nor UO_3297 (O_3297,N_49856,N_49980);
nor UO_3298 (O_3298,N_49866,N_49809);
xnor UO_3299 (O_3299,N_49951,N_49802);
and UO_3300 (O_3300,N_49760,N_49879);
nand UO_3301 (O_3301,N_49810,N_49933);
nor UO_3302 (O_3302,N_49961,N_49965);
and UO_3303 (O_3303,N_49853,N_49903);
and UO_3304 (O_3304,N_49866,N_49958);
and UO_3305 (O_3305,N_49930,N_49818);
nand UO_3306 (O_3306,N_49914,N_49875);
nor UO_3307 (O_3307,N_49792,N_49795);
xor UO_3308 (O_3308,N_49762,N_49850);
or UO_3309 (O_3309,N_49922,N_49973);
and UO_3310 (O_3310,N_49930,N_49958);
and UO_3311 (O_3311,N_49886,N_49860);
nor UO_3312 (O_3312,N_49779,N_49800);
and UO_3313 (O_3313,N_49754,N_49874);
and UO_3314 (O_3314,N_49916,N_49784);
xor UO_3315 (O_3315,N_49772,N_49890);
nand UO_3316 (O_3316,N_49858,N_49934);
xnor UO_3317 (O_3317,N_49793,N_49860);
and UO_3318 (O_3318,N_49779,N_49807);
nand UO_3319 (O_3319,N_49930,N_49855);
and UO_3320 (O_3320,N_49764,N_49937);
and UO_3321 (O_3321,N_49812,N_49772);
and UO_3322 (O_3322,N_49781,N_49852);
nor UO_3323 (O_3323,N_49907,N_49922);
xnor UO_3324 (O_3324,N_49900,N_49902);
and UO_3325 (O_3325,N_49971,N_49816);
xor UO_3326 (O_3326,N_49966,N_49986);
nand UO_3327 (O_3327,N_49928,N_49954);
or UO_3328 (O_3328,N_49789,N_49868);
nand UO_3329 (O_3329,N_49867,N_49768);
nand UO_3330 (O_3330,N_49893,N_49786);
and UO_3331 (O_3331,N_49951,N_49776);
and UO_3332 (O_3332,N_49913,N_49759);
and UO_3333 (O_3333,N_49904,N_49857);
or UO_3334 (O_3334,N_49804,N_49821);
nand UO_3335 (O_3335,N_49954,N_49896);
xnor UO_3336 (O_3336,N_49871,N_49985);
xor UO_3337 (O_3337,N_49820,N_49769);
nor UO_3338 (O_3338,N_49814,N_49979);
or UO_3339 (O_3339,N_49949,N_49803);
nand UO_3340 (O_3340,N_49817,N_49827);
and UO_3341 (O_3341,N_49956,N_49750);
nor UO_3342 (O_3342,N_49906,N_49924);
or UO_3343 (O_3343,N_49905,N_49770);
or UO_3344 (O_3344,N_49916,N_49764);
or UO_3345 (O_3345,N_49859,N_49801);
and UO_3346 (O_3346,N_49922,N_49918);
or UO_3347 (O_3347,N_49782,N_49768);
nor UO_3348 (O_3348,N_49759,N_49999);
xnor UO_3349 (O_3349,N_49930,N_49770);
xor UO_3350 (O_3350,N_49870,N_49894);
and UO_3351 (O_3351,N_49879,N_49830);
or UO_3352 (O_3352,N_49919,N_49995);
and UO_3353 (O_3353,N_49849,N_49911);
nor UO_3354 (O_3354,N_49969,N_49841);
nor UO_3355 (O_3355,N_49906,N_49986);
nand UO_3356 (O_3356,N_49965,N_49858);
or UO_3357 (O_3357,N_49779,N_49944);
nand UO_3358 (O_3358,N_49917,N_49856);
nand UO_3359 (O_3359,N_49780,N_49814);
or UO_3360 (O_3360,N_49776,N_49845);
or UO_3361 (O_3361,N_49814,N_49775);
xor UO_3362 (O_3362,N_49923,N_49821);
nand UO_3363 (O_3363,N_49753,N_49852);
and UO_3364 (O_3364,N_49755,N_49979);
nand UO_3365 (O_3365,N_49795,N_49969);
or UO_3366 (O_3366,N_49913,N_49858);
and UO_3367 (O_3367,N_49829,N_49827);
or UO_3368 (O_3368,N_49973,N_49998);
or UO_3369 (O_3369,N_49822,N_49813);
nor UO_3370 (O_3370,N_49771,N_49793);
and UO_3371 (O_3371,N_49861,N_49911);
nor UO_3372 (O_3372,N_49851,N_49866);
nor UO_3373 (O_3373,N_49989,N_49956);
and UO_3374 (O_3374,N_49806,N_49801);
and UO_3375 (O_3375,N_49988,N_49764);
or UO_3376 (O_3376,N_49752,N_49847);
or UO_3377 (O_3377,N_49864,N_49922);
nand UO_3378 (O_3378,N_49778,N_49930);
xnor UO_3379 (O_3379,N_49754,N_49905);
nand UO_3380 (O_3380,N_49809,N_49783);
xor UO_3381 (O_3381,N_49851,N_49854);
nor UO_3382 (O_3382,N_49829,N_49759);
and UO_3383 (O_3383,N_49998,N_49944);
nand UO_3384 (O_3384,N_49883,N_49929);
or UO_3385 (O_3385,N_49849,N_49946);
nand UO_3386 (O_3386,N_49902,N_49826);
nor UO_3387 (O_3387,N_49776,N_49843);
or UO_3388 (O_3388,N_49988,N_49945);
xnor UO_3389 (O_3389,N_49990,N_49998);
and UO_3390 (O_3390,N_49986,N_49953);
nor UO_3391 (O_3391,N_49919,N_49871);
nor UO_3392 (O_3392,N_49987,N_49996);
xnor UO_3393 (O_3393,N_49768,N_49855);
nand UO_3394 (O_3394,N_49940,N_49963);
or UO_3395 (O_3395,N_49938,N_49863);
or UO_3396 (O_3396,N_49829,N_49944);
and UO_3397 (O_3397,N_49831,N_49967);
and UO_3398 (O_3398,N_49810,N_49981);
and UO_3399 (O_3399,N_49825,N_49787);
xnor UO_3400 (O_3400,N_49873,N_49861);
or UO_3401 (O_3401,N_49767,N_49969);
or UO_3402 (O_3402,N_49978,N_49788);
nor UO_3403 (O_3403,N_49902,N_49845);
xnor UO_3404 (O_3404,N_49987,N_49960);
nor UO_3405 (O_3405,N_49786,N_49823);
nand UO_3406 (O_3406,N_49776,N_49863);
or UO_3407 (O_3407,N_49932,N_49845);
and UO_3408 (O_3408,N_49784,N_49928);
or UO_3409 (O_3409,N_49983,N_49840);
and UO_3410 (O_3410,N_49935,N_49881);
nor UO_3411 (O_3411,N_49813,N_49832);
and UO_3412 (O_3412,N_49823,N_49931);
nor UO_3413 (O_3413,N_49988,N_49853);
nand UO_3414 (O_3414,N_49837,N_49934);
and UO_3415 (O_3415,N_49790,N_49801);
or UO_3416 (O_3416,N_49870,N_49837);
and UO_3417 (O_3417,N_49891,N_49981);
or UO_3418 (O_3418,N_49862,N_49944);
nor UO_3419 (O_3419,N_49970,N_49944);
nor UO_3420 (O_3420,N_49912,N_49962);
xor UO_3421 (O_3421,N_49884,N_49836);
or UO_3422 (O_3422,N_49785,N_49943);
or UO_3423 (O_3423,N_49754,N_49800);
nor UO_3424 (O_3424,N_49842,N_49974);
nand UO_3425 (O_3425,N_49952,N_49799);
xor UO_3426 (O_3426,N_49842,N_49807);
nor UO_3427 (O_3427,N_49822,N_49986);
nand UO_3428 (O_3428,N_49919,N_49803);
or UO_3429 (O_3429,N_49912,N_49869);
xnor UO_3430 (O_3430,N_49822,N_49963);
xnor UO_3431 (O_3431,N_49840,N_49829);
nor UO_3432 (O_3432,N_49776,N_49774);
nor UO_3433 (O_3433,N_49785,N_49903);
nor UO_3434 (O_3434,N_49905,N_49953);
and UO_3435 (O_3435,N_49993,N_49856);
or UO_3436 (O_3436,N_49874,N_49787);
and UO_3437 (O_3437,N_49945,N_49815);
xor UO_3438 (O_3438,N_49848,N_49988);
nor UO_3439 (O_3439,N_49943,N_49866);
or UO_3440 (O_3440,N_49925,N_49873);
nor UO_3441 (O_3441,N_49896,N_49889);
nand UO_3442 (O_3442,N_49910,N_49801);
nand UO_3443 (O_3443,N_49943,N_49860);
and UO_3444 (O_3444,N_49886,N_49840);
and UO_3445 (O_3445,N_49871,N_49897);
xor UO_3446 (O_3446,N_49975,N_49771);
nand UO_3447 (O_3447,N_49946,N_49806);
nand UO_3448 (O_3448,N_49796,N_49835);
and UO_3449 (O_3449,N_49857,N_49912);
nor UO_3450 (O_3450,N_49800,N_49819);
xnor UO_3451 (O_3451,N_49888,N_49986);
nor UO_3452 (O_3452,N_49948,N_49988);
nand UO_3453 (O_3453,N_49995,N_49926);
and UO_3454 (O_3454,N_49930,N_49807);
or UO_3455 (O_3455,N_49921,N_49917);
nand UO_3456 (O_3456,N_49964,N_49995);
xor UO_3457 (O_3457,N_49759,N_49936);
nand UO_3458 (O_3458,N_49826,N_49789);
xor UO_3459 (O_3459,N_49964,N_49777);
nand UO_3460 (O_3460,N_49917,N_49769);
and UO_3461 (O_3461,N_49850,N_49829);
nor UO_3462 (O_3462,N_49815,N_49793);
nor UO_3463 (O_3463,N_49917,N_49998);
or UO_3464 (O_3464,N_49929,N_49833);
nor UO_3465 (O_3465,N_49920,N_49844);
nor UO_3466 (O_3466,N_49872,N_49827);
nand UO_3467 (O_3467,N_49981,N_49774);
and UO_3468 (O_3468,N_49766,N_49750);
and UO_3469 (O_3469,N_49917,N_49836);
nand UO_3470 (O_3470,N_49997,N_49908);
nor UO_3471 (O_3471,N_49982,N_49957);
nand UO_3472 (O_3472,N_49876,N_49773);
or UO_3473 (O_3473,N_49953,N_49963);
nor UO_3474 (O_3474,N_49990,N_49978);
nand UO_3475 (O_3475,N_49909,N_49870);
xnor UO_3476 (O_3476,N_49787,N_49911);
and UO_3477 (O_3477,N_49839,N_49937);
and UO_3478 (O_3478,N_49782,N_49835);
and UO_3479 (O_3479,N_49838,N_49790);
nor UO_3480 (O_3480,N_49797,N_49791);
nor UO_3481 (O_3481,N_49773,N_49967);
nand UO_3482 (O_3482,N_49826,N_49758);
xor UO_3483 (O_3483,N_49787,N_49949);
xor UO_3484 (O_3484,N_49870,N_49926);
nor UO_3485 (O_3485,N_49767,N_49914);
nand UO_3486 (O_3486,N_49827,N_49992);
nor UO_3487 (O_3487,N_49872,N_49990);
and UO_3488 (O_3488,N_49884,N_49853);
and UO_3489 (O_3489,N_49992,N_49790);
nand UO_3490 (O_3490,N_49824,N_49913);
xnor UO_3491 (O_3491,N_49811,N_49873);
nor UO_3492 (O_3492,N_49889,N_49915);
xor UO_3493 (O_3493,N_49815,N_49844);
nor UO_3494 (O_3494,N_49834,N_49959);
xor UO_3495 (O_3495,N_49983,N_49973);
nand UO_3496 (O_3496,N_49928,N_49879);
nand UO_3497 (O_3497,N_49834,N_49962);
or UO_3498 (O_3498,N_49924,N_49892);
nand UO_3499 (O_3499,N_49808,N_49791);
or UO_3500 (O_3500,N_49834,N_49971);
or UO_3501 (O_3501,N_49891,N_49999);
xor UO_3502 (O_3502,N_49919,N_49961);
or UO_3503 (O_3503,N_49980,N_49957);
and UO_3504 (O_3504,N_49780,N_49951);
or UO_3505 (O_3505,N_49796,N_49759);
xnor UO_3506 (O_3506,N_49904,N_49788);
and UO_3507 (O_3507,N_49923,N_49953);
xnor UO_3508 (O_3508,N_49939,N_49998);
nand UO_3509 (O_3509,N_49993,N_49819);
nand UO_3510 (O_3510,N_49892,N_49965);
nand UO_3511 (O_3511,N_49920,N_49896);
or UO_3512 (O_3512,N_49981,N_49922);
nand UO_3513 (O_3513,N_49817,N_49931);
xor UO_3514 (O_3514,N_49808,N_49920);
nor UO_3515 (O_3515,N_49859,N_49764);
and UO_3516 (O_3516,N_49942,N_49793);
and UO_3517 (O_3517,N_49917,N_49851);
nand UO_3518 (O_3518,N_49893,N_49967);
or UO_3519 (O_3519,N_49928,N_49750);
xor UO_3520 (O_3520,N_49807,N_49804);
and UO_3521 (O_3521,N_49920,N_49810);
nand UO_3522 (O_3522,N_49956,N_49900);
and UO_3523 (O_3523,N_49835,N_49843);
nand UO_3524 (O_3524,N_49987,N_49928);
xor UO_3525 (O_3525,N_49775,N_49846);
and UO_3526 (O_3526,N_49930,N_49845);
xnor UO_3527 (O_3527,N_49837,N_49941);
nand UO_3528 (O_3528,N_49812,N_49967);
nor UO_3529 (O_3529,N_49909,N_49910);
nand UO_3530 (O_3530,N_49846,N_49786);
or UO_3531 (O_3531,N_49854,N_49755);
and UO_3532 (O_3532,N_49760,N_49910);
xnor UO_3533 (O_3533,N_49886,N_49836);
and UO_3534 (O_3534,N_49934,N_49909);
nor UO_3535 (O_3535,N_49831,N_49857);
or UO_3536 (O_3536,N_49941,N_49989);
xnor UO_3537 (O_3537,N_49958,N_49895);
nor UO_3538 (O_3538,N_49992,N_49787);
nor UO_3539 (O_3539,N_49875,N_49794);
nand UO_3540 (O_3540,N_49943,N_49955);
xnor UO_3541 (O_3541,N_49812,N_49769);
nand UO_3542 (O_3542,N_49957,N_49992);
and UO_3543 (O_3543,N_49774,N_49885);
and UO_3544 (O_3544,N_49781,N_49962);
xnor UO_3545 (O_3545,N_49928,N_49979);
xnor UO_3546 (O_3546,N_49809,N_49937);
and UO_3547 (O_3547,N_49853,N_49759);
or UO_3548 (O_3548,N_49782,N_49891);
xnor UO_3549 (O_3549,N_49893,N_49957);
or UO_3550 (O_3550,N_49881,N_49900);
and UO_3551 (O_3551,N_49782,N_49943);
and UO_3552 (O_3552,N_49815,N_49971);
xnor UO_3553 (O_3553,N_49808,N_49774);
and UO_3554 (O_3554,N_49879,N_49852);
nand UO_3555 (O_3555,N_49831,N_49984);
nand UO_3556 (O_3556,N_49966,N_49902);
and UO_3557 (O_3557,N_49812,N_49993);
or UO_3558 (O_3558,N_49922,N_49877);
or UO_3559 (O_3559,N_49885,N_49805);
nor UO_3560 (O_3560,N_49794,N_49837);
nor UO_3561 (O_3561,N_49987,N_49969);
nor UO_3562 (O_3562,N_49884,N_49938);
nor UO_3563 (O_3563,N_49968,N_49977);
xor UO_3564 (O_3564,N_49819,N_49848);
nor UO_3565 (O_3565,N_49920,N_49826);
nand UO_3566 (O_3566,N_49930,N_49851);
and UO_3567 (O_3567,N_49910,N_49816);
nand UO_3568 (O_3568,N_49898,N_49986);
nand UO_3569 (O_3569,N_49992,N_49821);
nand UO_3570 (O_3570,N_49752,N_49818);
or UO_3571 (O_3571,N_49911,N_49854);
or UO_3572 (O_3572,N_49863,N_49802);
and UO_3573 (O_3573,N_49798,N_49910);
nand UO_3574 (O_3574,N_49910,N_49877);
nand UO_3575 (O_3575,N_49813,N_49961);
and UO_3576 (O_3576,N_49914,N_49850);
and UO_3577 (O_3577,N_49880,N_49797);
nand UO_3578 (O_3578,N_49874,N_49953);
xor UO_3579 (O_3579,N_49873,N_49897);
nand UO_3580 (O_3580,N_49784,N_49768);
nand UO_3581 (O_3581,N_49897,N_49947);
or UO_3582 (O_3582,N_49755,N_49851);
nand UO_3583 (O_3583,N_49783,N_49976);
or UO_3584 (O_3584,N_49913,N_49839);
and UO_3585 (O_3585,N_49883,N_49765);
nand UO_3586 (O_3586,N_49841,N_49944);
or UO_3587 (O_3587,N_49818,N_49862);
or UO_3588 (O_3588,N_49787,N_49871);
nor UO_3589 (O_3589,N_49991,N_49837);
nor UO_3590 (O_3590,N_49859,N_49898);
nor UO_3591 (O_3591,N_49957,N_49753);
nor UO_3592 (O_3592,N_49975,N_49949);
or UO_3593 (O_3593,N_49826,N_49957);
and UO_3594 (O_3594,N_49872,N_49836);
or UO_3595 (O_3595,N_49891,N_49929);
nor UO_3596 (O_3596,N_49969,N_49790);
or UO_3597 (O_3597,N_49892,N_49783);
nor UO_3598 (O_3598,N_49899,N_49752);
and UO_3599 (O_3599,N_49813,N_49874);
and UO_3600 (O_3600,N_49849,N_49985);
nand UO_3601 (O_3601,N_49754,N_49806);
and UO_3602 (O_3602,N_49776,N_49925);
nor UO_3603 (O_3603,N_49833,N_49780);
xor UO_3604 (O_3604,N_49877,N_49920);
xnor UO_3605 (O_3605,N_49807,N_49962);
xor UO_3606 (O_3606,N_49930,N_49853);
xnor UO_3607 (O_3607,N_49874,N_49758);
nor UO_3608 (O_3608,N_49995,N_49940);
xor UO_3609 (O_3609,N_49882,N_49891);
nor UO_3610 (O_3610,N_49929,N_49965);
xnor UO_3611 (O_3611,N_49991,N_49811);
or UO_3612 (O_3612,N_49884,N_49993);
nand UO_3613 (O_3613,N_49962,N_49931);
xor UO_3614 (O_3614,N_49914,N_49815);
nand UO_3615 (O_3615,N_49979,N_49854);
or UO_3616 (O_3616,N_49879,N_49927);
nor UO_3617 (O_3617,N_49759,N_49750);
nor UO_3618 (O_3618,N_49975,N_49761);
and UO_3619 (O_3619,N_49751,N_49900);
xor UO_3620 (O_3620,N_49821,N_49854);
or UO_3621 (O_3621,N_49882,N_49885);
nand UO_3622 (O_3622,N_49891,N_49818);
nor UO_3623 (O_3623,N_49750,N_49788);
nor UO_3624 (O_3624,N_49928,N_49982);
and UO_3625 (O_3625,N_49837,N_49954);
nand UO_3626 (O_3626,N_49962,N_49883);
nand UO_3627 (O_3627,N_49966,N_49820);
or UO_3628 (O_3628,N_49900,N_49845);
xor UO_3629 (O_3629,N_49956,N_49899);
nor UO_3630 (O_3630,N_49900,N_49869);
nand UO_3631 (O_3631,N_49845,N_49765);
nand UO_3632 (O_3632,N_49917,N_49905);
xnor UO_3633 (O_3633,N_49966,N_49933);
and UO_3634 (O_3634,N_49944,N_49816);
xnor UO_3635 (O_3635,N_49976,N_49812);
or UO_3636 (O_3636,N_49883,N_49983);
nand UO_3637 (O_3637,N_49778,N_49819);
and UO_3638 (O_3638,N_49828,N_49980);
nor UO_3639 (O_3639,N_49826,N_49855);
and UO_3640 (O_3640,N_49994,N_49914);
or UO_3641 (O_3641,N_49753,N_49777);
xnor UO_3642 (O_3642,N_49848,N_49861);
nor UO_3643 (O_3643,N_49794,N_49956);
and UO_3644 (O_3644,N_49750,N_49970);
nand UO_3645 (O_3645,N_49832,N_49946);
and UO_3646 (O_3646,N_49899,N_49776);
or UO_3647 (O_3647,N_49960,N_49769);
nor UO_3648 (O_3648,N_49757,N_49810);
or UO_3649 (O_3649,N_49961,N_49979);
nor UO_3650 (O_3650,N_49889,N_49835);
or UO_3651 (O_3651,N_49927,N_49962);
and UO_3652 (O_3652,N_49846,N_49802);
nor UO_3653 (O_3653,N_49818,N_49849);
nand UO_3654 (O_3654,N_49997,N_49930);
nand UO_3655 (O_3655,N_49774,N_49864);
or UO_3656 (O_3656,N_49756,N_49991);
or UO_3657 (O_3657,N_49863,N_49937);
xor UO_3658 (O_3658,N_49933,N_49929);
or UO_3659 (O_3659,N_49902,N_49754);
and UO_3660 (O_3660,N_49842,N_49940);
xor UO_3661 (O_3661,N_49771,N_49761);
nor UO_3662 (O_3662,N_49874,N_49905);
nor UO_3663 (O_3663,N_49778,N_49919);
or UO_3664 (O_3664,N_49851,N_49846);
xor UO_3665 (O_3665,N_49881,N_49891);
nand UO_3666 (O_3666,N_49977,N_49859);
nor UO_3667 (O_3667,N_49940,N_49934);
nor UO_3668 (O_3668,N_49954,N_49828);
xor UO_3669 (O_3669,N_49996,N_49981);
nor UO_3670 (O_3670,N_49937,N_49910);
xnor UO_3671 (O_3671,N_49757,N_49984);
and UO_3672 (O_3672,N_49763,N_49856);
nand UO_3673 (O_3673,N_49858,N_49846);
nand UO_3674 (O_3674,N_49814,N_49770);
and UO_3675 (O_3675,N_49873,N_49806);
and UO_3676 (O_3676,N_49966,N_49765);
nor UO_3677 (O_3677,N_49905,N_49969);
nand UO_3678 (O_3678,N_49971,N_49999);
or UO_3679 (O_3679,N_49868,N_49890);
or UO_3680 (O_3680,N_49757,N_49917);
or UO_3681 (O_3681,N_49889,N_49837);
or UO_3682 (O_3682,N_49801,N_49816);
nand UO_3683 (O_3683,N_49798,N_49987);
xnor UO_3684 (O_3684,N_49903,N_49991);
xnor UO_3685 (O_3685,N_49835,N_49794);
and UO_3686 (O_3686,N_49925,N_49772);
or UO_3687 (O_3687,N_49935,N_49756);
or UO_3688 (O_3688,N_49976,N_49869);
and UO_3689 (O_3689,N_49980,N_49925);
and UO_3690 (O_3690,N_49828,N_49969);
nand UO_3691 (O_3691,N_49775,N_49977);
or UO_3692 (O_3692,N_49836,N_49805);
nand UO_3693 (O_3693,N_49927,N_49956);
or UO_3694 (O_3694,N_49971,N_49787);
or UO_3695 (O_3695,N_49964,N_49918);
nor UO_3696 (O_3696,N_49944,N_49861);
or UO_3697 (O_3697,N_49938,N_49911);
xor UO_3698 (O_3698,N_49808,N_49839);
or UO_3699 (O_3699,N_49989,N_49881);
or UO_3700 (O_3700,N_49762,N_49958);
nor UO_3701 (O_3701,N_49892,N_49986);
and UO_3702 (O_3702,N_49782,N_49874);
and UO_3703 (O_3703,N_49860,N_49870);
nand UO_3704 (O_3704,N_49923,N_49827);
or UO_3705 (O_3705,N_49822,N_49903);
xnor UO_3706 (O_3706,N_49898,N_49796);
xnor UO_3707 (O_3707,N_49756,N_49812);
nor UO_3708 (O_3708,N_49864,N_49975);
nor UO_3709 (O_3709,N_49929,N_49987);
nor UO_3710 (O_3710,N_49768,N_49922);
nand UO_3711 (O_3711,N_49865,N_49832);
nor UO_3712 (O_3712,N_49912,N_49991);
nand UO_3713 (O_3713,N_49929,N_49792);
xnor UO_3714 (O_3714,N_49946,N_49804);
nor UO_3715 (O_3715,N_49769,N_49895);
xnor UO_3716 (O_3716,N_49847,N_49785);
and UO_3717 (O_3717,N_49987,N_49792);
or UO_3718 (O_3718,N_49956,N_49936);
or UO_3719 (O_3719,N_49836,N_49770);
xnor UO_3720 (O_3720,N_49898,N_49809);
xor UO_3721 (O_3721,N_49815,N_49985);
or UO_3722 (O_3722,N_49933,N_49957);
or UO_3723 (O_3723,N_49997,N_49830);
and UO_3724 (O_3724,N_49990,N_49974);
xor UO_3725 (O_3725,N_49820,N_49856);
nor UO_3726 (O_3726,N_49860,N_49912);
or UO_3727 (O_3727,N_49844,N_49853);
and UO_3728 (O_3728,N_49962,N_49964);
xor UO_3729 (O_3729,N_49814,N_49850);
or UO_3730 (O_3730,N_49890,N_49955);
nand UO_3731 (O_3731,N_49783,N_49984);
nor UO_3732 (O_3732,N_49998,N_49901);
nor UO_3733 (O_3733,N_49787,N_49947);
or UO_3734 (O_3734,N_49782,N_49845);
and UO_3735 (O_3735,N_49866,N_49942);
nor UO_3736 (O_3736,N_49787,N_49938);
nand UO_3737 (O_3737,N_49964,N_49996);
nor UO_3738 (O_3738,N_49785,N_49839);
nor UO_3739 (O_3739,N_49928,N_49846);
and UO_3740 (O_3740,N_49877,N_49995);
or UO_3741 (O_3741,N_49914,N_49965);
and UO_3742 (O_3742,N_49959,N_49859);
nand UO_3743 (O_3743,N_49834,N_49925);
xnor UO_3744 (O_3744,N_49752,N_49794);
nor UO_3745 (O_3745,N_49824,N_49810);
nor UO_3746 (O_3746,N_49777,N_49781);
or UO_3747 (O_3747,N_49890,N_49921);
xnor UO_3748 (O_3748,N_49790,N_49983);
nor UO_3749 (O_3749,N_49853,N_49788);
nand UO_3750 (O_3750,N_49783,N_49802);
or UO_3751 (O_3751,N_49922,N_49885);
nor UO_3752 (O_3752,N_49752,N_49864);
xor UO_3753 (O_3753,N_49960,N_49862);
or UO_3754 (O_3754,N_49913,N_49856);
nand UO_3755 (O_3755,N_49941,N_49959);
xnor UO_3756 (O_3756,N_49849,N_49758);
nand UO_3757 (O_3757,N_49969,N_49997);
nor UO_3758 (O_3758,N_49980,N_49950);
nand UO_3759 (O_3759,N_49816,N_49855);
nand UO_3760 (O_3760,N_49858,N_49996);
nor UO_3761 (O_3761,N_49990,N_49942);
or UO_3762 (O_3762,N_49809,N_49786);
nor UO_3763 (O_3763,N_49820,N_49812);
or UO_3764 (O_3764,N_49985,N_49788);
xnor UO_3765 (O_3765,N_49962,N_49786);
and UO_3766 (O_3766,N_49803,N_49975);
or UO_3767 (O_3767,N_49835,N_49922);
nand UO_3768 (O_3768,N_49892,N_49879);
nand UO_3769 (O_3769,N_49894,N_49796);
xnor UO_3770 (O_3770,N_49959,N_49758);
nor UO_3771 (O_3771,N_49893,N_49975);
nor UO_3772 (O_3772,N_49840,N_49868);
and UO_3773 (O_3773,N_49794,N_49777);
nor UO_3774 (O_3774,N_49884,N_49977);
or UO_3775 (O_3775,N_49771,N_49789);
and UO_3776 (O_3776,N_49994,N_49847);
nand UO_3777 (O_3777,N_49856,N_49785);
xor UO_3778 (O_3778,N_49862,N_49962);
or UO_3779 (O_3779,N_49990,N_49842);
nand UO_3780 (O_3780,N_49978,N_49951);
xnor UO_3781 (O_3781,N_49860,N_49917);
and UO_3782 (O_3782,N_49908,N_49883);
nor UO_3783 (O_3783,N_49753,N_49946);
xor UO_3784 (O_3784,N_49913,N_49941);
nor UO_3785 (O_3785,N_49797,N_49825);
or UO_3786 (O_3786,N_49925,N_49927);
and UO_3787 (O_3787,N_49816,N_49951);
or UO_3788 (O_3788,N_49866,N_49877);
or UO_3789 (O_3789,N_49992,N_49826);
nand UO_3790 (O_3790,N_49967,N_49945);
nand UO_3791 (O_3791,N_49944,N_49897);
and UO_3792 (O_3792,N_49856,N_49953);
nor UO_3793 (O_3793,N_49777,N_49970);
nand UO_3794 (O_3794,N_49780,N_49876);
nor UO_3795 (O_3795,N_49948,N_49849);
or UO_3796 (O_3796,N_49843,N_49888);
xor UO_3797 (O_3797,N_49785,N_49783);
nor UO_3798 (O_3798,N_49979,N_49908);
nand UO_3799 (O_3799,N_49883,N_49866);
xor UO_3800 (O_3800,N_49855,N_49801);
or UO_3801 (O_3801,N_49994,N_49867);
xnor UO_3802 (O_3802,N_49804,N_49923);
xor UO_3803 (O_3803,N_49820,N_49987);
and UO_3804 (O_3804,N_49880,N_49877);
and UO_3805 (O_3805,N_49815,N_49934);
or UO_3806 (O_3806,N_49855,N_49858);
xor UO_3807 (O_3807,N_49943,N_49770);
nand UO_3808 (O_3808,N_49853,N_49775);
nand UO_3809 (O_3809,N_49992,N_49997);
and UO_3810 (O_3810,N_49820,N_49886);
nor UO_3811 (O_3811,N_49972,N_49773);
nor UO_3812 (O_3812,N_49823,N_49752);
nor UO_3813 (O_3813,N_49870,N_49817);
xnor UO_3814 (O_3814,N_49967,N_49880);
nor UO_3815 (O_3815,N_49928,N_49756);
xor UO_3816 (O_3816,N_49877,N_49830);
or UO_3817 (O_3817,N_49802,N_49787);
or UO_3818 (O_3818,N_49753,N_49841);
xor UO_3819 (O_3819,N_49758,N_49981);
and UO_3820 (O_3820,N_49843,N_49770);
or UO_3821 (O_3821,N_49918,N_49872);
nor UO_3822 (O_3822,N_49838,N_49757);
nor UO_3823 (O_3823,N_49865,N_49932);
or UO_3824 (O_3824,N_49816,N_49893);
nor UO_3825 (O_3825,N_49798,N_49925);
nor UO_3826 (O_3826,N_49757,N_49977);
and UO_3827 (O_3827,N_49892,N_49909);
xor UO_3828 (O_3828,N_49896,N_49902);
or UO_3829 (O_3829,N_49909,N_49826);
and UO_3830 (O_3830,N_49759,N_49897);
nand UO_3831 (O_3831,N_49824,N_49877);
nor UO_3832 (O_3832,N_49879,N_49831);
nor UO_3833 (O_3833,N_49896,N_49969);
nand UO_3834 (O_3834,N_49840,N_49890);
nor UO_3835 (O_3835,N_49997,N_49843);
nor UO_3836 (O_3836,N_49792,N_49862);
and UO_3837 (O_3837,N_49903,N_49889);
and UO_3838 (O_3838,N_49753,N_49763);
nor UO_3839 (O_3839,N_49790,N_49874);
and UO_3840 (O_3840,N_49814,N_49986);
nor UO_3841 (O_3841,N_49789,N_49828);
xor UO_3842 (O_3842,N_49964,N_49811);
and UO_3843 (O_3843,N_49829,N_49794);
nand UO_3844 (O_3844,N_49962,N_49958);
and UO_3845 (O_3845,N_49990,N_49786);
nand UO_3846 (O_3846,N_49904,N_49767);
nand UO_3847 (O_3847,N_49750,N_49782);
and UO_3848 (O_3848,N_49789,N_49770);
nor UO_3849 (O_3849,N_49924,N_49780);
or UO_3850 (O_3850,N_49974,N_49936);
nor UO_3851 (O_3851,N_49908,N_49921);
nand UO_3852 (O_3852,N_49859,N_49967);
or UO_3853 (O_3853,N_49831,N_49808);
nand UO_3854 (O_3854,N_49771,N_49831);
xnor UO_3855 (O_3855,N_49983,N_49876);
xnor UO_3856 (O_3856,N_49820,N_49833);
xnor UO_3857 (O_3857,N_49854,N_49867);
and UO_3858 (O_3858,N_49979,N_49937);
xnor UO_3859 (O_3859,N_49834,N_49930);
and UO_3860 (O_3860,N_49793,N_49862);
nand UO_3861 (O_3861,N_49975,N_49942);
and UO_3862 (O_3862,N_49874,N_49955);
nand UO_3863 (O_3863,N_49869,N_49968);
xnor UO_3864 (O_3864,N_49863,N_49906);
nor UO_3865 (O_3865,N_49858,N_49876);
nand UO_3866 (O_3866,N_49835,N_49828);
nand UO_3867 (O_3867,N_49765,N_49788);
xnor UO_3868 (O_3868,N_49967,N_49968);
xnor UO_3869 (O_3869,N_49951,N_49923);
nand UO_3870 (O_3870,N_49816,N_49761);
xnor UO_3871 (O_3871,N_49987,N_49812);
nand UO_3872 (O_3872,N_49769,N_49751);
and UO_3873 (O_3873,N_49828,N_49923);
nand UO_3874 (O_3874,N_49807,N_49862);
or UO_3875 (O_3875,N_49899,N_49995);
and UO_3876 (O_3876,N_49987,N_49930);
and UO_3877 (O_3877,N_49822,N_49994);
or UO_3878 (O_3878,N_49962,N_49775);
xnor UO_3879 (O_3879,N_49957,N_49922);
and UO_3880 (O_3880,N_49789,N_49975);
nor UO_3881 (O_3881,N_49981,N_49910);
nand UO_3882 (O_3882,N_49934,N_49987);
and UO_3883 (O_3883,N_49896,N_49781);
or UO_3884 (O_3884,N_49902,N_49981);
nor UO_3885 (O_3885,N_49792,N_49855);
nand UO_3886 (O_3886,N_49938,N_49902);
or UO_3887 (O_3887,N_49914,N_49762);
or UO_3888 (O_3888,N_49893,N_49941);
or UO_3889 (O_3889,N_49881,N_49800);
nor UO_3890 (O_3890,N_49763,N_49819);
and UO_3891 (O_3891,N_49987,N_49823);
or UO_3892 (O_3892,N_49856,N_49818);
and UO_3893 (O_3893,N_49809,N_49801);
xnor UO_3894 (O_3894,N_49777,N_49906);
or UO_3895 (O_3895,N_49985,N_49952);
xor UO_3896 (O_3896,N_49934,N_49913);
xnor UO_3897 (O_3897,N_49925,N_49914);
xnor UO_3898 (O_3898,N_49951,N_49897);
nor UO_3899 (O_3899,N_49950,N_49884);
or UO_3900 (O_3900,N_49984,N_49980);
or UO_3901 (O_3901,N_49957,N_49878);
or UO_3902 (O_3902,N_49788,N_49994);
nand UO_3903 (O_3903,N_49791,N_49760);
nand UO_3904 (O_3904,N_49820,N_49979);
or UO_3905 (O_3905,N_49943,N_49790);
and UO_3906 (O_3906,N_49850,N_49818);
and UO_3907 (O_3907,N_49972,N_49777);
and UO_3908 (O_3908,N_49772,N_49977);
or UO_3909 (O_3909,N_49895,N_49781);
nor UO_3910 (O_3910,N_49991,N_49932);
nand UO_3911 (O_3911,N_49769,N_49879);
xnor UO_3912 (O_3912,N_49889,N_49830);
nor UO_3913 (O_3913,N_49798,N_49826);
or UO_3914 (O_3914,N_49913,N_49862);
xnor UO_3915 (O_3915,N_49819,N_49801);
xnor UO_3916 (O_3916,N_49794,N_49911);
nor UO_3917 (O_3917,N_49882,N_49773);
nor UO_3918 (O_3918,N_49806,N_49937);
and UO_3919 (O_3919,N_49861,N_49865);
and UO_3920 (O_3920,N_49985,N_49806);
and UO_3921 (O_3921,N_49754,N_49899);
nand UO_3922 (O_3922,N_49762,N_49988);
nand UO_3923 (O_3923,N_49879,N_49751);
nor UO_3924 (O_3924,N_49798,N_49954);
nor UO_3925 (O_3925,N_49905,N_49867);
nor UO_3926 (O_3926,N_49770,N_49788);
nand UO_3927 (O_3927,N_49876,N_49869);
nor UO_3928 (O_3928,N_49849,N_49857);
xor UO_3929 (O_3929,N_49840,N_49832);
or UO_3930 (O_3930,N_49770,N_49983);
or UO_3931 (O_3931,N_49899,N_49986);
nand UO_3932 (O_3932,N_49901,N_49819);
and UO_3933 (O_3933,N_49883,N_49785);
xnor UO_3934 (O_3934,N_49812,N_49858);
xnor UO_3935 (O_3935,N_49774,N_49869);
xnor UO_3936 (O_3936,N_49868,N_49882);
or UO_3937 (O_3937,N_49936,N_49931);
or UO_3938 (O_3938,N_49968,N_49874);
xor UO_3939 (O_3939,N_49947,N_49926);
nand UO_3940 (O_3940,N_49825,N_49849);
xor UO_3941 (O_3941,N_49991,N_49828);
nor UO_3942 (O_3942,N_49988,N_49819);
nor UO_3943 (O_3943,N_49892,N_49830);
nand UO_3944 (O_3944,N_49788,N_49761);
or UO_3945 (O_3945,N_49781,N_49858);
and UO_3946 (O_3946,N_49775,N_49970);
nand UO_3947 (O_3947,N_49907,N_49970);
and UO_3948 (O_3948,N_49807,N_49827);
nor UO_3949 (O_3949,N_49855,N_49863);
xnor UO_3950 (O_3950,N_49841,N_49807);
nor UO_3951 (O_3951,N_49790,N_49926);
xor UO_3952 (O_3952,N_49884,N_49932);
nor UO_3953 (O_3953,N_49930,N_49886);
xnor UO_3954 (O_3954,N_49882,N_49880);
and UO_3955 (O_3955,N_49862,N_49822);
nor UO_3956 (O_3956,N_49796,N_49934);
and UO_3957 (O_3957,N_49759,N_49971);
nand UO_3958 (O_3958,N_49870,N_49942);
nand UO_3959 (O_3959,N_49896,N_49942);
or UO_3960 (O_3960,N_49818,N_49858);
and UO_3961 (O_3961,N_49945,N_49783);
and UO_3962 (O_3962,N_49841,N_49799);
or UO_3963 (O_3963,N_49803,N_49901);
nand UO_3964 (O_3964,N_49912,N_49984);
nor UO_3965 (O_3965,N_49985,N_49774);
nand UO_3966 (O_3966,N_49821,N_49999);
and UO_3967 (O_3967,N_49988,N_49874);
or UO_3968 (O_3968,N_49811,N_49900);
and UO_3969 (O_3969,N_49949,N_49980);
and UO_3970 (O_3970,N_49956,N_49815);
or UO_3971 (O_3971,N_49832,N_49863);
or UO_3972 (O_3972,N_49913,N_49870);
or UO_3973 (O_3973,N_49969,N_49782);
or UO_3974 (O_3974,N_49792,N_49922);
xnor UO_3975 (O_3975,N_49812,N_49807);
nor UO_3976 (O_3976,N_49912,N_49916);
xor UO_3977 (O_3977,N_49809,N_49855);
or UO_3978 (O_3978,N_49821,N_49937);
nor UO_3979 (O_3979,N_49882,N_49806);
nor UO_3980 (O_3980,N_49869,N_49917);
or UO_3981 (O_3981,N_49762,N_49868);
nor UO_3982 (O_3982,N_49858,N_49859);
or UO_3983 (O_3983,N_49799,N_49859);
and UO_3984 (O_3984,N_49855,N_49812);
nand UO_3985 (O_3985,N_49967,N_49927);
or UO_3986 (O_3986,N_49767,N_49997);
nand UO_3987 (O_3987,N_49872,N_49940);
nand UO_3988 (O_3988,N_49879,N_49781);
nor UO_3989 (O_3989,N_49984,N_49847);
or UO_3990 (O_3990,N_49755,N_49905);
nor UO_3991 (O_3991,N_49799,N_49892);
xnor UO_3992 (O_3992,N_49768,N_49881);
xnor UO_3993 (O_3993,N_49917,N_49762);
nor UO_3994 (O_3994,N_49786,N_49929);
or UO_3995 (O_3995,N_49905,N_49990);
or UO_3996 (O_3996,N_49772,N_49863);
nor UO_3997 (O_3997,N_49877,N_49810);
xnor UO_3998 (O_3998,N_49999,N_49975);
or UO_3999 (O_3999,N_49845,N_49759);
or UO_4000 (O_4000,N_49768,N_49916);
and UO_4001 (O_4001,N_49885,N_49814);
xnor UO_4002 (O_4002,N_49934,N_49914);
and UO_4003 (O_4003,N_49941,N_49855);
nor UO_4004 (O_4004,N_49818,N_49773);
nor UO_4005 (O_4005,N_49769,N_49920);
xnor UO_4006 (O_4006,N_49785,N_49809);
nand UO_4007 (O_4007,N_49770,N_49771);
xor UO_4008 (O_4008,N_49881,N_49921);
and UO_4009 (O_4009,N_49982,N_49758);
xnor UO_4010 (O_4010,N_49839,N_49894);
xor UO_4011 (O_4011,N_49916,N_49860);
xor UO_4012 (O_4012,N_49983,N_49870);
nor UO_4013 (O_4013,N_49905,N_49866);
or UO_4014 (O_4014,N_49792,N_49803);
nand UO_4015 (O_4015,N_49964,N_49752);
or UO_4016 (O_4016,N_49780,N_49760);
nand UO_4017 (O_4017,N_49862,N_49927);
xnor UO_4018 (O_4018,N_49905,N_49800);
and UO_4019 (O_4019,N_49943,N_49842);
and UO_4020 (O_4020,N_49844,N_49981);
nand UO_4021 (O_4021,N_49981,N_49967);
nor UO_4022 (O_4022,N_49775,N_49872);
or UO_4023 (O_4023,N_49830,N_49780);
nor UO_4024 (O_4024,N_49765,N_49804);
nor UO_4025 (O_4025,N_49967,N_49830);
xnor UO_4026 (O_4026,N_49924,N_49931);
nor UO_4027 (O_4027,N_49948,N_49863);
and UO_4028 (O_4028,N_49846,N_49993);
and UO_4029 (O_4029,N_49772,N_49911);
nor UO_4030 (O_4030,N_49999,N_49859);
nor UO_4031 (O_4031,N_49943,N_49826);
or UO_4032 (O_4032,N_49820,N_49830);
nand UO_4033 (O_4033,N_49977,N_49938);
nand UO_4034 (O_4034,N_49975,N_49963);
xnor UO_4035 (O_4035,N_49916,N_49819);
or UO_4036 (O_4036,N_49931,N_49986);
nor UO_4037 (O_4037,N_49797,N_49960);
xor UO_4038 (O_4038,N_49806,N_49965);
nand UO_4039 (O_4039,N_49783,N_49797);
or UO_4040 (O_4040,N_49845,N_49998);
nand UO_4041 (O_4041,N_49904,N_49931);
or UO_4042 (O_4042,N_49993,N_49770);
xnor UO_4043 (O_4043,N_49843,N_49953);
or UO_4044 (O_4044,N_49912,N_49891);
xor UO_4045 (O_4045,N_49884,N_49960);
nand UO_4046 (O_4046,N_49891,N_49954);
or UO_4047 (O_4047,N_49968,N_49882);
nand UO_4048 (O_4048,N_49936,N_49856);
and UO_4049 (O_4049,N_49795,N_49909);
nand UO_4050 (O_4050,N_49809,N_49766);
nand UO_4051 (O_4051,N_49751,N_49953);
nand UO_4052 (O_4052,N_49805,N_49865);
xor UO_4053 (O_4053,N_49930,N_49919);
xnor UO_4054 (O_4054,N_49779,N_49798);
and UO_4055 (O_4055,N_49889,N_49973);
and UO_4056 (O_4056,N_49793,N_49800);
xnor UO_4057 (O_4057,N_49887,N_49883);
or UO_4058 (O_4058,N_49930,N_49812);
or UO_4059 (O_4059,N_49979,N_49849);
nand UO_4060 (O_4060,N_49833,N_49855);
nor UO_4061 (O_4061,N_49985,N_49797);
nand UO_4062 (O_4062,N_49827,N_49761);
nand UO_4063 (O_4063,N_49996,N_49889);
nor UO_4064 (O_4064,N_49937,N_49915);
and UO_4065 (O_4065,N_49931,N_49991);
nand UO_4066 (O_4066,N_49860,N_49895);
nand UO_4067 (O_4067,N_49993,N_49810);
and UO_4068 (O_4068,N_49830,N_49813);
nand UO_4069 (O_4069,N_49880,N_49790);
nor UO_4070 (O_4070,N_49873,N_49803);
or UO_4071 (O_4071,N_49946,N_49779);
nand UO_4072 (O_4072,N_49871,N_49845);
xnor UO_4073 (O_4073,N_49771,N_49786);
or UO_4074 (O_4074,N_49886,N_49780);
and UO_4075 (O_4075,N_49969,N_49951);
or UO_4076 (O_4076,N_49962,N_49754);
or UO_4077 (O_4077,N_49952,N_49947);
xnor UO_4078 (O_4078,N_49824,N_49865);
or UO_4079 (O_4079,N_49851,N_49849);
or UO_4080 (O_4080,N_49952,N_49945);
xnor UO_4081 (O_4081,N_49831,N_49775);
nand UO_4082 (O_4082,N_49840,N_49909);
and UO_4083 (O_4083,N_49939,N_49997);
nand UO_4084 (O_4084,N_49888,N_49905);
xnor UO_4085 (O_4085,N_49869,N_49955);
or UO_4086 (O_4086,N_49830,N_49984);
or UO_4087 (O_4087,N_49813,N_49901);
nor UO_4088 (O_4088,N_49814,N_49781);
nor UO_4089 (O_4089,N_49798,N_49784);
and UO_4090 (O_4090,N_49999,N_49791);
nand UO_4091 (O_4091,N_49852,N_49801);
nand UO_4092 (O_4092,N_49906,N_49786);
nor UO_4093 (O_4093,N_49844,N_49993);
or UO_4094 (O_4094,N_49772,N_49943);
nor UO_4095 (O_4095,N_49758,N_49916);
xnor UO_4096 (O_4096,N_49913,N_49777);
and UO_4097 (O_4097,N_49916,N_49998);
or UO_4098 (O_4098,N_49959,N_49923);
xnor UO_4099 (O_4099,N_49978,N_49985);
or UO_4100 (O_4100,N_49939,N_49957);
and UO_4101 (O_4101,N_49808,N_49926);
or UO_4102 (O_4102,N_49952,N_49967);
nand UO_4103 (O_4103,N_49894,N_49780);
xor UO_4104 (O_4104,N_49779,N_49848);
and UO_4105 (O_4105,N_49971,N_49763);
nand UO_4106 (O_4106,N_49904,N_49897);
nand UO_4107 (O_4107,N_49992,N_49858);
nor UO_4108 (O_4108,N_49840,N_49808);
nand UO_4109 (O_4109,N_49769,N_49837);
xnor UO_4110 (O_4110,N_49786,N_49983);
nand UO_4111 (O_4111,N_49775,N_49941);
xor UO_4112 (O_4112,N_49777,N_49815);
nor UO_4113 (O_4113,N_49860,N_49950);
and UO_4114 (O_4114,N_49979,N_49769);
nand UO_4115 (O_4115,N_49827,N_49984);
xor UO_4116 (O_4116,N_49840,N_49814);
nand UO_4117 (O_4117,N_49807,N_49935);
and UO_4118 (O_4118,N_49997,N_49762);
or UO_4119 (O_4119,N_49926,N_49942);
and UO_4120 (O_4120,N_49778,N_49847);
or UO_4121 (O_4121,N_49896,N_49953);
xnor UO_4122 (O_4122,N_49999,N_49893);
nand UO_4123 (O_4123,N_49885,N_49934);
or UO_4124 (O_4124,N_49858,N_49986);
or UO_4125 (O_4125,N_49881,N_49967);
or UO_4126 (O_4126,N_49917,N_49955);
or UO_4127 (O_4127,N_49970,N_49889);
xnor UO_4128 (O_4128,N_49769,N_49934);
or UO_4129 (O_4129,N_49975,N_49793);
nand UO_4130 (O_4130,N_49752,N_49862);
nand UO_4131 (O_4131,N_49778,N_49948);
and UO_4132 (O_4132,N_49901,N_49771);
nor UO_4133 (O_4133,N_49867,N_49940);
and UO_4134 (O_4134,N_49826,N_49976);
xnor UO_4135 (O_4135,N_49830,N_49826);
xor UO_4136 (O_4136,N_49969,N_49847);
xor UO_4137 (O_4137,N_49857,N_49809);
and UO_4138 (O_4138,N_49807,N_49967);
and UO_4139 (O_4139,N_49947,N_49833);
nor UO_4140 (O_4140,N_49830,N_49845);
nand UO_4141 (O_4141,N_49814,N_49968);
and UO_4142 (O_4142,N_49920,N_49869);
nor UO_4143 (O_4143,N_49958,N_49815);
or UO_4144 (O_4144,N_49753,N_49797);
nand UO_4145 (O_4145,N_49816,N_49802);
nor UO_4146 (O_4146,N_49851,N_49947);
nor UO_4147 (O_4147,N_49841,N_49956);
nand UO_4148 (O_4148,N_49809,N_49932);
nor UO_4149 (O_4149,N_49895,N_49817);
nand UO_4150 (O_4150,N_49911,N_49999);
nand UO_4151 (O_4151,N_49955,N_49995);
xnor UO_4152 (O_4152,N_49867,N_49792);
or UO_4153 (O_4153,N_49809,N_49862);
nor UO_4154 (O_4154,N_49918,N_49926);
and UO_4155 (O_4155,N_49925,N_49894);
or UO_4156 (O_4156,N_49918,N_49820);
nor UO_4157 (O_4157,N_49919,N_49833);
or UO_4158 (O_4158,N_49904,N_49935);
nor UO_4159 (O_4159,N_49852,N_49752);
or UO_4160 (O_4160,N_49784,N_49811);
and UO_4161 (O_4161,N_49889,N_49985);
xor UO_4162 (O_4162,N_49842,N_49791);
xnor UO_4163 (O_4163,N_49880,N_49825);
or UO_4164 (O_4164,N_49752,N_49802);
xnor UO_4165 (O_4165,N_49910,N_49936);
nand UO_4166 (O_4166,N_49818,N_49884);
nand UO_4167 (O_4167,N_49938,N_49924);
and UO_4168 (O_4168,N_49751,N_49918);
nand UO_4169 (O_4169,N_49836,N_49908);
and UO_4170 (O_4170,N_49966,N_49881);
xnor UO_4171 (O_4171,N_49768,N_49930);
nor UO_4172 (O_4172,N_49797,N_49919);
nand UO_4173 (O_4173,N_49844,N_49769);
nor UO_4174 (O_4174,N_49773,N_49801);
and UO_4175 (O_4175,N_49901,N_49796);
or UO_4176 (O_4176,N_49965,N_49845);
nand UO_4177 (O_4177,N_49864,N_49771);
nand UO_4178 (O_4178,N_49867,N_49925);
nor UO_4179 (O_4179,N_49828,N_49975);
nand UO_4180 (O_4180,N_49752,N_49962);
or UO_4181 (O_4181,N_49769,N_49904);
nor UO_4182 (O_4182,N_49987,N_49931);
xor UO_4183 (O_4183,N_49997,N_49811);
xnor UO_4184 (O_4184,N_49861,N_49796);
nor UO_4185 (O_4185,N_49904,N_49785);
nand UO_4186 (O_4186,N_49944,N_49992);
nand UO_4187 (O_4187,N_49974,N_49922);
nand UO_4188 (O_4188,N_49786,N_49842);
or UO_4189 (O_4189,N_49966,N_49769);
and UO_4190 (O_4190,N_49765,N_49964);
and UO_4191 (O_4191,N_49763,N_49988);
nand UO_4192 (O_4192,N_49792,N_49787);
xnor UO_4193 (O_4193,N_49845,N_49917);
xor UO_4194 (O_4194,N_49956,N_49862);
nand UO_4195 (O_4195,N_49793,N_49976);
and UO_4196 (O_4196,N_49780,N_49797);
xor UO_4197 (O_4197,N_49897,N_49784);
xor UO_4198 (O_4198,N_49959,N_49857);
or UO_4199 (O_4199,N_49801,N_49911);
nand UO_4200 (O_4200,N_49918,N_49778);
nor UO_4201 (O_4201,N_49808,N_49965);
and UO_4202 (O_4202,N_49867,N_49972);
xnor UO_4203 (O_4203,N_49892,N_49983);
and UO_4204 (O_4204,N_49876,N_49908);
and UO_4205 (O_4205,N_49851,N_49960);
nor UO_4206 (O_4206,N_49840,N_49771);
nand UO_4207 (O_4207,N_49980,N_49982);
nor UO_4208 (O_4208,N_49851,N_49802);
nand UO_4209 (O_4209,N_49945,N_49998);
nor UO_4210 (O_4210,N_49990,N_49935);
xor UO_4211 (O_4211,N_49794,N_49885);
nor UO_4212 (O_4212,N_49804,N_49836);
xnor UO_4213 (O_4213,N_49790,N_49936);
nor UO_4214 (O_4214,N_49903,N_49849);
nand UO_4215 (O_4215,N_49851,N_49826);
or UO_4216 (O_4216,N_49966,N_49893);
nand UO_4217 (O_4217,N_49903,N_49791);
and UO_4218 (O_4218,N_49912,N_49772);
nand UO_4219 (O_4219,N_49948,N_49782);
or UO_4220 (O_4220,N_49831,N_49858);
nor UO_4221 (O_4221,N_49998,N_49981);
xor UO_4222 (O_4222,N_49768,N_49944);
nand UO_4223 (O_4223,N_49850,N_49766);
nor UO_4224 (O_4224,N_49935,N_49851);
xor UO_4225 (O_4225,N_49858,N_49817);
nor UO_4226 (O_4226,N_49789,N_49804);
nand UO_4227 (O_4227,N_49766,N_49954);
xnor UO_4228 (O_4228,N_49789,N_49855);
or UO_4229 (O_4229,N_49851,N_49793);
nand UO_4230 (O_4230,N_49921,N_49882);
nor UO_4231 (O_4231,N_49894,N_49933);
and UO_4232 (O_4232,N_49900,N_49848);
and UO_4233 (O_4233,N_49873,N_49770);
xnor UO_4234 (O_4234,N_49842,N_49904);
or UO_4235 (O_4235,N_49968,N_49888);
or UO_4236 (O_4236,N_49848,N_49922);
xnor UO_4237 (O_4237,N_49866,N_49911);
or UO_4238 (O_4238,N_49943,N_49983);
nor UO_4239 (O_4239,N_49949,N_49973);
nand UO_4240 (O_4240,N_49898,N_49913);
xor UO_4241 (O_4241,N_49761,N_49944);
nor UO_4242 (O_4242,N_49837,N_49995);
nor UO_4243 (O_4243,N_49967,N_49935);
or UO_4244 (O_4244,N_49951,N_49767);
xor UO_4245 (O_4245,N_49805,N_49803);
or UO_4246 (O_4246,N_49830,N_49750);
and UO_4247 (O_4247,N_49760,N_49994);
or UO_4248 (O_4248,N_49906,N_49874);
and UO_4249 (O_4249,N_49783,N_49981);
nand UO_4250 (O_4250,N_49940,N_49810);
nor UO_4251 (O_4251,N_49842,N_49969);
and UO_4252 (O_4252,N_49927,N_49807);
nand UO_4253 (O_4253,N_49833,N_49825);
nor UO_4254 (O_4254,N_49833,N_49917);
or UO_4255 (O_4255,N_49998,N_49774);
and UO_4256 (O_4256,N_49877,N_49819);
xor UO_4257 (O_4257,N_49789,N_49761);
xnor UO_4258 (O_4258,N_49960,N_49905);
or UO_4259 (O_4259,N_49889,N_49801);
xnor UO_4260 (O_4260,N_49811,N_49760);
or UO_4261 (O_4261,N_49871,N_49782);
nor UO_4262 (O_4262,N_49784,N_49893);
and UO_4263 (O_4263,N_49817,N_49990);
or UO_4264 (O_4264,N_49948,N_49913);
xnor UO_4265 (O_4265,N_49976,N_49750);
nand UO_4266 (O_4266,N_49979,N_49870);
nand UO_4267 (O_4267,N_49867,N_49888);
and UO_4268 (O_4268,N_49912,N_49750);
nand UO_4269 (O_4269,N_49842,N_49810);
xor UO_4270 (O_4270,N_49932,N_49813);
nand UO_4271 (O_4271,N_49763,N_49954);
xor UO_4272 (O_4272,N_49963,N_49983);
nand UO_4273 (O_4273,N_49840,N_49922);
nor UO_4274 (O_4274,N_49932,N_49939);
nor UO_4275 (O_4275,N_49896,N_49837);
or UO_4276 (O_4276,N_49932,N_49774);
or UO_4277 (O_4277,N_49779,N_49866);
nor UO_4278 (O_4278,N_49981,N_49865);
or UO_4279 (O_4279,N_49789,N_49836);
nand UO_4280 (O_4280,N_49933,N_49905);
or UO_4281 (O_4281,N_49956,N_49852);
xnor UO_4282 (O_4282,N_49752,N_49987);
nand UO_4283 (O_4283,N_49842,N_49764);
xor UO_4284 (O_4284,N_49994,N_49825);
or UO_4285 (O_4285,N_49772,N_49843);
nand UO_4286 (O_4286,N_49879,N_49880);
and UO_4287 (O_4287,N_49911,N_49992);
and UO_4288 (O_4288,N_49895,N_49759);
xnor UO_4289 (O_4289,N_49985,N_49843);
nor UO_4290 (O_4290,N_49823,N_49923);
nor UO_4291 (O_4291,N_49816,N_49796);
and UO_4292 (O_4292,N_49902,N_49876);
nor UO_4293 (O_4293,N_49888,N_49809);
nor UO_4294 (O_4294,N_49791,N_49756);
or UO_4295 (O_4295,N_49985,N_49837);
or UO_4296 (O_4296,N_49783,N_49969);
xor UO_4297 (O_4297,N_49893,N_49936);
xor UO_4298 (O_4298,N_49866,N_49914);
nand UO_4299 (O_4299,N_49780,N_49771);
or UO_4300 (O_4300,N_49904,N_49957);
and UO_4301 (O_4301,N_49815,N_49752);
xor UO_4302 (O_4302,N_49898,N_49802);
nor UO_4303 (O_4303,N_49813,N_49993);
or UO_4304 (O_4304,N_49957,N_49886);
or UO_4305 (O_4305,N_49802,N_49839);
or UO_4306 (O_4306,N_49801,N_49947);
nor UO_4307 (O_4307,N_49839,N_49813);
nor UO_4308 (O_4308,N_49837,N_49900);
nor UO_4309 (O_4309,N_49839,N_49959);
nand UO_4310 (O_4310,N_49762,N_49915);
nor UO_4311 (O_4311,N_49987,N_49982);
nor UO_4312 (O_4312,N_49836,N_49893);
or UO_4313 (O_4313,N_49905,N_49818);
and UO_4314 (O_4314,N_49903,N_49984);
or UO_4315 (O_4315,N_49951,N_49779);
xor UO_4316 (O_4316,N_49776,N_49750);
or UO_4317 (O_4317,N_49962,N_49764);
and UO_4318 (O_4318,N_49893,N_49856);
xor UO_4319 (O_4319,N_49996,N_49787);
and UO_4320 (O_4320,N_49885,N_49771);
nand UO_4321 (O_4321,N_49864,N_49998);
and UO_4322 (O_4322,N_49976,N_49904);
xnor UO_4323 (O_4323,N_49954,N_49786);
or UO_4324 (O_4324,N_49872,N_49773);
or UO_4325 (O_4325,N_49838,N_49950);
nand UO_4326 (O_4326,N_49829,N_49791);
xnor UO_4327 (O_4327,N_49812,N_49767);
nor UO_4328 (O_4328,N_49834,N_49754);
nor UO_4329 (O_4329,N_49768,N_49917);
nor UO_4330 (O_4330,N_49796,N_49873);
nand UO_4331 (O_4331,N_49899,N_49854);
nand UO_4332 (O_4332,N_49983,N_49961);
or UO_4333 (O_4333,N_49881,N_49956);
nor UO_4334 (O_4334,N_49800,N_49795);
and UO_4335 (O_4335,N_49906,N_49829);
nor UO_4336 (O_4336,N_49783,N_49999);
xnor UO_4337 (O_4337,N_49921,N_49785);
xnor UO_4338 (O_4338,N_49897,N_49930);
and UO_4339 (O_4339,N_49766,N_49842);
nor UO_4340 (O_4340,N_49855,N_49997);
nor UO_4341 (O_4341,N_49792,N_49832);
and UO_4342 (O_4342,N_49854,N_49844);
or UO_4343 (O_4343,N_49901,N_49797);
or UO_4344 (O_4344,N_49768,N_49815);
and UO_4345 (O_4345,N_49905,N_49826);
xor UO_4346 (O_4346,N_49932,N_49927);
xnor UO_4347 (O_4347,N_49866,N_49888);
nand UO_4348 (O_4348,N_49918,N_49825);
nor UO_4349 (O_4349,N_49786,N_49850);
xor UO_4350 (O_4350,N_49880,N_49966);
and UO_4351 (O_4351,N_49870,N_49914);
or UO_4352 (O_4352,N_49919,N_49798);
xnor UO_4353 (O_4353,N_49860,N_49832);
nor UO_4354 (O_4354,N_49871,N_49835);
nor UO_4355 (O_4355,N_49852,N_49991);
xor UO_4356 (O_4356,N_49765,N_49955);
xor UO_4357 (O_4357,N_49820,N_49946);
or UO_4358 (O_4358,N_49841,N_49899);
nor UO_4359 (O_4359,N_49792,N_49943);
nor UO_4360 (O_4360,N_49807,N_49808);
xor UO_4361 (O_4361,N_49758,N_49998);
xnor UO_4362 (O_4362,N_49968,N_49863);
nand UO_4363 (O_4363,N_49988,N_49898);
nand UO_4364 (O_4364,N_49844,N_49777);
nor UO_4365 (O_4365,N_49903,N_49862);
nor UO_4366 (O_4366,N_49816,N_49852);
nor UO_4367 (O_4367,N_49903,N_49989);
nor UO_4368 (O_4368,N_49946,N_49934);
xnor UO_4369 (O_4369,N_49929,N_49795);
nor UO_4370 (O_4370,N_49901,N_49961);
or UO_4371 (O_4371,N_49802,N_49798);
nand UO_4372 (O_4372,N_49926,N_49928);
and UO_4373 (O_4373,N_49845,N_49977);
or UO_4374 (O_4374,N_49845,N_49926);
or UO_4375 (O_4375,N_49903,N_49901);
nor UO_4376 (O_4376,N_49890,N_49846);
nor UO_4377 (O_4377,N_49863,N_49870);
xnor UO_4378 (O_4378,N_49991,N_49826);
xnor UO_4379 (O_4379,N_49814,N_49829);
nor UO_4380 (O_4380,N_49850,N_49774);
and UO_4381 (O_4381,N_49756,N_49817);
nor UO_4382 (O_4382,N_49945,N_49890);
xor UO_4383 (O_4383,N_49795,N_49808);
xnor UO_4384 (O_4384,N_49965,N_49993);
nand UO_4385 (O_4385,N_49996,N_49888);
or UO_4386 (O_4386,N_49979,N_49776);
xor UO_4387 (O_4387,N_49815,N_49992);
and UO_4388 (O_4388,N_49926,N_49754);
and UO_4389 (O_4389,N_49901,N_49908);
xnor UO_4390 (O_4390,N_49887,N_49956);
and UO_4391 (O_4391,N_49984,N_49806);
xor UO_4392 (O_4392,N_49885,N_49751);
nand UO_4393 (O_4393,N_49918,N_49766);
or UO_4394 (O_4394,N_49894,N_49931);
nand UO_4395 (O_4395,N_49929,N_49770);
nor UO_4396 (O_4396,N_49937,N_49904);
or UO_4397 (O_4397,N_49792,N_49944);
and UO_4398 (O_4398,N_49951,N_49910);
and UO_4399 (O_4399,N_49907,N_49998);
nand UO_4400 (O_4400,N_49847,N_49761);
xnor UO_4401 (O_4401,N_49850,N_49819);
and UO_4402 (O_4402,N_49968,N_49753);
xor UO_4403 (O_4403,N_49752,N_49936);
nand UO_4404 (O_4404,N_49817,N_49787);
or UO_4405 (O_4405,N_49750,N_49860);
and UO_4406 (O_4406,N_49813,N_49795);
and UO_4407 (O_4407,N_49866,N_49922);
xnor UO_4408 (O_4408,N_49917,N_49837);
xor UO_4409 (O_4409,N_49802,N_49757);
or UO_4410 (O_4410,N_49759,N_49966);
xor UO_4411 (O_4411,N_49824,N_49909);
and UO_4412 (O_4412,N_49927,N_49984);
nand UO_4413 (O_4413,N_49815,N_49817);
xnor UO_4414 (O_4414,N_49822,N_49753);
nor UO_4415 (O_4415,N_49887,N_49902);
xnor UO_4416 (O_4416,N_49800,N_49826);
and UO_4417 (O_4417,N_49815,N_49764);
nor UO_4418 (O_4418,N_49860,N_49955);
and UO_4419 (O_4419,N_49973,N_49813);
xor UO_4420 (O_4420,N_49810,N_49753);
xnor UO_4421 (O_4421,N_49783,N_49933);
nand UO_4422 (O_4422,N_49859,N_49886);
or UO_4423 (O_4423,N_49794,N_49994);
and UO_4424 (O_4424,N_49877,N_49773);
nor UO_4425 (O_4425,N_49774,N_49947);
and UO_4426 (O_4426,N_49905,N_49772);
xor UO_4427 (O_4427,N_49849,N_49993);
or UO_4428 (O_4428,N_49877,N_49843);
and UO_4429 (O_4429,N_49808,N_49758);
or UO_4430 (O_4430,N_49887,N_49888);
xnor UO_4431 (O_4431,N_49911,N_49960);
xnor UO_4432 (O_4432,N_49998,N_49914);
and UO_4433 (O_4433,N_49768,N_49907);
xnor UO_4434 (O_4434,N_49986,N_49850);
nand UO_4435 (O_4435,N_49790,N_49840);
nand UO_4436 (O_4436,N_49847,N_49848);
or UO_4437 (O_4437,N_49768,N_49909);
xor UO_4438 (O_4438,N_49866,N_49940);
or UO_4439 (O_4439,N_49807,N_49923);
nand UO_4440 (O_4440,N_49908,N_49976);
and UO_4441 (O_4441,N_49853,N_49837);
and UO_4442 (O_4442,N_49857,N_49850);
and UO_4443 (O_4443,N_49996,N_49930);
and UO_4444 (O_4444,N_49908,N_49858);
or UO_4445 (O_4445,N_49783,N_49935);
xnor UO_4446 (O_4446,N_49783,N_49947);
nor UO_4447 (O_4447,N_49861,N_49756);
or UO_4448 (O_4448,N_49878,N_49845);
nor UO_4449 (O_4449,N_49912,N_49785);
nor UO_4450 (O_4450,N_49787,N_49934);
nor UO_4451 (O_4451,N_49883,N_49886);
nor UO_4452 (O_4452,N_49856,N_49784);
nand UO_4453 (O_4453,N_49852,N_49811);
and UO_4454 (O_4454,N_49919,N_49829);
xnor UO_4455 (O_4455,N_49849,N_49801);
nor UO_4456 (O_4456,N_49888,N_49758);
nand UO_4457 (O_4457,N_49971,N_49785);
nand UO_4458 (O_4458,N_49963,N_49807);
or UO_4459 (O_4459,N_49988,N_49789);
and UO_4460 (O_4460,N_49893,N_49753);
xnor UO_4461 (O_4461,N_49801,N_49750);
and UO_4462 (O_4462,N_49953,N_49783);
and UO_4463 (O_4463,N_49988,N_49942);
nor UO_4464 (O_4464,N_49800,N_49949);
xor UO_4465 (O_4465,N_49907,N_49872);
or UO_4466 (O_4466,N_49794,N_49867);
nor UO_4467 (O_4467,N_49920,N_49866);
xnor UO_4468 (O_4468,N_49854,N_49970);
xnor UO_4469 (O_4469,N_49807,N_49788);
nor UO_4470 (O_4470,N_49818,N_49885);
nor UO_4471 (O_4471,N_49758,N_49819);
nand UO_4472 (O_4472,N_49765,N_49932);
or UO_4473 (O_4473,N_49928,N_49960);
nand UO_4474 (O_4474,N_49970,N_49787);
nand UO_4475 (O_4475,N_49996,N_49931);
nand UO_4476 (O_4476,N_49969,N_49810);
nor UO_4477 (O_4477,N_49877,N_49876);
xor UO_4478 (O_4478,N_49968,N_49942);
or UO_4479 (O_4479,N_49845,N_49851);
nand UO_4480 (O_4480,N_49941,N_49777);
xor UO_4481 (O_4481,N_49903,N_49815);
nor UO_4482 (O_4482,N_49941,N_49914);
xnor UO_4483 (O_4483,N_49829,N_49911);
nand UO_4484 (O_4484,N_49838,N_49818);
xnor UO_4485 (O_4485,N_49925,N_49917);
xor UO_4486 (O_4486,N_49958,N_49928);
xnor UO_4487 (O_4487,N_49838,N_49865);
nor UO_4488 (O_4488,N_49965,N_49932);
or UO_4489 (O_4489,N_49830,N_49981);
and UO_4490 (O_4490,N_49994,N_49782);
nand UO_4491 (O_4491,N_49817,N_49832);
and UO_4492 (O_4492,N_49939,N_49913);
or UO_4493 (O_4493,N_49899,N_49877);
nor UO_4494 (O_4494,N_49843,N_49920);
or UO_4495 (O_4495,N_49795,N_49878);
and UO_4496 (O_4496,N_49852,N_49858);
or UO_4497 (O_4497,N_49873,N_49929);
or UO_4498 (O_4498,N_49846,N_49938);
nand UO_4499 (O_4499,N_49826,N_49844);
nor UO_4500 (O_4500,N_49887,N_49870);
or UO_4501 (O_4501,N_49914,N_49825);
xor UO_4502 (O_4502,N_49936,N_49799);
nand UO_4503 (O_4503,N_49879,N_49999);
and UO_4504 (O_4504,N_49982,N_49877);
and UO_4505 (O_4505,N_49798,N_49900);
or UO_4506 (O_4506,N_49951,N_49762);
xor UO_4507 (O_4507,N_49881,N_49756);
nor UO_4508 (O_4508,N_49809,N_49928);
or UO_4509 (O_4509,N_49791,N_49809);
and UO_4510 (O_4510,N_49868,N_49862);
nand UO_4511 (O_4511,N_49793,N_49923);
nand UO_4512 (O_4512,N_49863,N_49828);
or UO_4513 (O_4513,N_49772,N_49791);
nor UO_4514 (O_4514,N_49760,N_49925);
nand UO_4515 (O_4515,N_49997,N_49758);
and UO_4516 (O_4516,N_49930,N_49871);
nor UO_4517 (O_4517,N_49868,N_49937);
nand UO_4518 (O_4518,N_49957,N_49916);
nor UO_4519 (O_4519,N_49790,N_49915);
nand UO_4520 (O_4520,N_49991,N_49829);
nor UO_4521 (O_4521,N_49813,N_49807);
or UO_4522 (O_4522,N_49846,N_49970);
or UO_4523 (O_4523,N_49873,N_49876);
or UO_4524 (O_4524,N_49895,N_49910);
xor UO_4525 (O_4525,N_49843,N_49930);
or UO_4526 (O_4526,N_49854,N_49765);
nand UO_4527 (O_4527,N_49788,N_49825);
and UO_4528 (O_4528,N_49758,N_49848);
nor UO_4529 (O_4529,N_49785,N_49891);
and UO_4530 (O_4530,N_49870,N_49936);
xnor UO_4531 (O_4531,N_49939,N_49754);
or UO_4532 (O_4532,N_49807,N_49882);
xnor UO_4533 (O_4533,N_49898,N_49770);
and UO_4534 (O_4534,N_49855,N_49780);
xnor UO_4535 (O_4535,N_49954,N_49827);
nand UO_4536 (O_4536,N_49900,N_49895);
xnor UO_4537 (O_4537,N_49795,N_49804);
nand UO_4538 (O_4538,N_49886,N_49752);
xnor UO_4539 (O_4539,N_49845,N_49920);
and UO_4540 (O_4540,N_49806,N_49823);
and UO_4541 (O_4541,N_49803,N_49797);
nor UO_4542 (O_4542,N_49959,N_49971);
xnor UO_4543 (O_4543,N_49779,N_49788);
or UO_4544 (O_4544,N_49901,N_49946);
nand UO_4545 (O_4545,N_49868,N_49936);
xnor UO_4546 (O_4546,N_49958,N_49805);
or UO_4547 (O_4547,N_49765,N_49778);
xnor UO_4548 (O_4548,N_49865,N_49807);
xnor UO_4549 (O_4549,N_49881,N_49802);
or UO_4550 (O_4550,N_49821,N_49881);
nor UO_4551 (O_4551,N_49932,N_49823);
and UO_4552 (O_4552,N_49768,N_49820);
nand UO_4553 (O_4553,N_49873,N_49818);
or UO_4554 (O_4554,N_49973,N_49765);
xnor UO_4555 (O_4555,N_49972,N_49976);
and UO_4556 (O_4556,N_49752,N_49761);
nand UO_4557 (O_4557,N_49845,N_49903);
nor UO_4558 (O_4558,N_49974,N_49814);
nand UO_4559 (O_4559,N_49901,N_49886);
xor UO_4560 (O_4560,N_49802,N_49755);
nand UO_4561 (O_4561,N_49794,N_49874);
and UO_4562 (O_4562,N_49931,N_49898);
or UO_4563 (O_4563,N_49982,N_49848);
and UO_4564 (O_4564,N_49906,N_49845);
nand UO_4565 (O_4565,N_49971,N_49772);
or UO_4566 (O_4566,N_49803,N_49963);
xnor UO_4567 (O_4567,N_49930,N_49885);
or UO_4568 (O_4568,N_49935,N_49791);
nor UO_4569 (O_4569,N_49819,N_49994);
nor UO_4570 (O_4570,N_49755,N_49855);
and UO_4571 (O_4571,N_49902,N_49804);
nand UO_4572 (O_4572,N_49901,N_49862);
nor UO_4573 (O_4573,N_49904,N_49778);
xor UO_4574 (O_4574,N_49759,N_49834);
and UO_4575 (O_4575,N_49937,N_49877);
xor UO_4576 (O_4576,N_49965,N_49753);
nand UO_4577 (O_4577,N_49966,N_49752);
nor UO_4578 (O_4578,N_49869,N_49934);
or UO_4579 (O_4579,N_49940,N_49973);
nand UO_4580 (O_4580,N_49945,N_49786);
xnor UO_4581 (O_4581,N_49902,N_49927);
nand UO_4582 (O_4582,N_49887,N_49889);
xor UO_4583 (O_4583,N_49944,N_49934);
nand UO_4584 (O_4584,N_49791,N_49847);
and UO_4585 (O_4585,N_49888,N_49972);
nor UO_4586 (O_4586,N_49774,N_49768);
and UO_4587 (O_4587,N_49988,N_49946);
nor UO_4588 (O_4588,N_49781,N_49756);
or UO_4589 (O_4589,N_49934,N_49829);
and UO_4590 (O_4590,N_49945,N_49785);
xor UO_4591 (O_4591,N_49764,N_49923);
or UO_4592 (O_4592,N_49855,N_49861);
or UO_4593 (O_4593,N_49786,N_49774);
nor UO_4594 (O_4594,N_49956,N_49951);
nand UO_4595 (O_4595,N_49818,N_49845);
xnor UO_4596 (O_4596,N_49864,N_49899);
or UO_4597 (O_4597,N_49767,N_49890);
xor UO_4598 (O_4598,N_49867,N_49922);
nor UO_4599 (O_4599,N_49757,N_49769);
nor UO_4600 (O_4600,N_49837,N_49812);
xor UO_4601 (O_4601,N_49946,N_49776);
nand UO_4602 (O_4602,N_49830,N_49770);
or UO_4603 (O_4603,N_49985,N_49909);
xor UO_4604 (O_4604,N_49958,N_49804);
nand UO_4605 (O_4605,N_49955,N_49931);
nand UO_4606 (O_4606,N_49793,N_49937);
nand UO_4607 (O_4607,N_49927,N_49982);
nand UO_4608 (O_4608,N_49849,N_49931);
or UO_4609 (O_4609,N_49920,N_49880);
and UO_4610 (O_4610,N_49961,N_49756);
nor UO_4611 (O_4611,N_49993,N_49794);
nand UO_4612 (O_4612,N_49771,N_49768);
nor UO_4613 (O_4613,N_49884,N_49967);
xnor UO_4614 (O_4614,N_49990,N_49899);
and UO_4615 (O_4615,N_49889,N_49992);
xnor UO_4616 (O_4616,N_49944,N_49849);
and UO_4617 (O_4617,N_49810,N_49889);
xor UO_4618 (O_4618,N_49905,N_49999);
xor UO_4619 (O_4619,N_49853,N_49962);
nor UO_4620 (O_4620,N_49811,N_49977);
nor UO_4621 (O_4621,N_49927,N_49867);
nand UO_4622 (O_4622,N_49787,N_49833);
or UO_4623 (O_4623,N_49929,N_49881);
nand UO_4624 (O_4624,N_49782,N_49898);
and UO_4625 (O_4625,N_49948,N_49925);
xor UO_4626 (O_4626,N_49950,N_49784);
nor UO_4627 (O_4627,N_49955,N_49812);
and UO_4628 (O_4628,N_49820,N_49787);
nor UO_4629 (O_4629,N_49759,N_49860);
nand UO_4630 (O_4630,N_49859,N_49910);
and UO_4631 (O_4631,N_49932,N_49938);
nand UO_4632 (O_4632,N_49830,N_49801);
xnor UO_4633 (O_4633,N_49888,N_49989);
nor UO_4634 (O_4634,N_49857,N_49801);
or UO_4635 (O_4635,N_49978,N_49974);
nor UO_4636 (O_4636,N_49939,N_49912);
or UO_4637 (O_4637,N_49862,N_49835);
xor UO_4638 (O_4638,N_49800,N_49916);
nor UO_4639 (O_4639,N_49750,N_49837);
xnor UO_4640 (O_4640,N_49797,N_49774);
and UO_4641 (O_4641,N_49888,N_49878);
xnor UO_4642 (O_4642,N_49951,N_49914);
and UO_4643 (O_4643,N_49918,N_49799);
or UO_4644 (O_4644,N_49760,N_49907);
nand UO_4645 (O_4645,N_49918,N_49857);
xnor UO_4646 (O_4646,N_49895,N_49813);
nor UO_4647 (O_4647,N_49804,N_49813);
xnor UO_4648 (O_4648,N_49777,N_49999);
or UO_4649 (O_4649,N_49895,N_49867);
or UO_4650 (O_4650,N_49958,N_49817);
nor UO_4651 (O_4651,N_49914,N_49811);
and UO_4652 (O_4652,N_49915,N_49854);
nor UO_4653 (O_4653,N_49851,N_49958);
nor UO_4654 (O_4654,N_49965,N_49899);
or UO_4655 (O_4655,N_49995,N_49965);
and UO_4656 (O_4656,N_49909,N_49873);
xnor UO_4657 (O_4657,N_49827,N_49941);
and UO_4658 (O_4658,N_49839,N_49962);
nand UO_4659 (O_4659,N_49881,N_49865);
xor UO_4660 (O_4660,N_49809,N_49967);
xor UO_4661 (O_4661,N_49823,N_49856);
nand UO_4662 (O_4662,N_49900,N_49809);
nor UO_4663 (O_4663,N_49918,N_49769);
nand UO_4664 (O_4664,N_49810,N_49985);
or UO_4665 (O_4665,N_49816,N_49921);
nand UO_4666 (O_4666,N_49858,N_49840);
xor UO_4667 (O_4667,N_49764,N_49961);
xnor UO_4668 (O_4668,N_49793,N_49974);
or UO_4669 (O_4669,N_49996,N_49873);
and UO_4670 (O_4670,N_49978,N_49988);
xor UO_4671 (O_4671,N_49755,N_49989);
and UO_4672 (O_4672,N_49832,N_49752);
xor UO_4673 (O_4673,N_49931,N_49757);
nand UO_4674 (O_4674,N_49930,N_49760);
nor UO_4675 (O_4675,N_49750,N_49757);
nand UO_4676 (O_4676,N_49793,N_49778);
and UO_4677 (O_4677,N_49836,N_49885);
nor UO_4678 (O_4678,N_49906,N_49900);
or UO_4679 (O_4679,N_49874,N_49891);
nor UO_4680 (O_4680,N_49823,N_49896);
and UO_4681 (O_4681,N_49887,N_49758);
nand UO_4682 (O_4682,N_49765,N_49928);
nor UO_4683 (O_4683,N_49932,N_49907);
xnor UO_4684 (O_4684,N_49962,N_49974);
or UO_4685 (O_4685,N_49830,N_49805);
or UO_4686 (O_4686,N_49784,N_49781);
xor UO_4687 (O_4687,N_49970,N_49851);
or UO_4688 (O_4688,N_49909,N_49898);
or UO_4689 (O_4689,N_49926,N_49787);
xor UO_4690 (O_4690,N_49814,N_49778);
xor UO_4691 (O_4691,N_49949,N_49827);
nand UO_4692 (O_4692,N_49842,N_49976);
or UO_4693 (O_4693,N_49956,N_49993);
or UO_4694 (O_4694,N_49995,N_49855);
or UO_4695 (O_4695,N_49858,N_49907);
or UO_4696 (O_4696,N_49853,N_49839);
or UO_4697 (O_4697,N_49954,N_49814);
and UO_4698 (O_4698,N_49872,N_49842);
or UO_4699 (O_4699,N_49940,N_49989);
nand UO_4700 (O_4700,N_49796,N_49806);
nor UO_4701 (O_4701,N_49773,N_49776);
nor UO_4702 (O_4702,N_49903,N_49807);
or UO_4703 (O_4703,N_49795,N_49888);
nor UO_4704 (O_4704,N_49891,N_49801);
and UO_4705 (O_4705,N_49850,N_49891);
nor UO_4706 (O_4706,N_49878,N_49877);
or UO_4707 (O_4707,N_49871,N_49992);
nor UO_4708 (O_4708,N_49943,N_49861);
and UO_4709 (O_4709,N_49998,N_49833);
nor UO_4710 (O_4710,N_49936,N_49845);
and UO_4711 (O_4711,N_49977,N_49819);
and UO_4712 (O_4712,N_49983,N_49931);
and UO_4713 (O_4713,N_49802,N_49772);
xor UO_4714 (O_4714,N_49807,N_49965);
or UO_4715 (O_4715,N_49868,N_49823);
or UO_4716 (O_4716,N_49958,N_49944);
and UO_4717 (O_4717,N_49766,N_49816);
or UO_4718 (O_4718,N_49907,N_49868);
and UO_4719 (O_4719,N_49927,N_49842);
and UO_4720 (O_4720,N_49887,N_49779);
nand UO_4721 (O_4721,N_49849,N_49998);
xnor UO_4722 (O_4722,N_49886,N_49993);
nor UO_4723 (O_4723,N_49981,N_49771);
nor UO_4724 (O_4724,N_49771,N_49775);
xnor UO_4725 (O_4725,N_49941,N_49853);
or UO_4726 (O_4726,N_49897,N_49806);
xnor UO_4727 (O_4727,N_49848,N_49959);
or UO_4728 (O_4728,N_49888,N_49773);
and UO_4729 (O_4729,N_49889,N_49900);
or UO_4730 (O_4730,N_49831,N_49802);
xnor UO_4731 (O_4731,N_49860,N_49894);
and UO_4732 (O_4732,N_49841,N_49980);
or UO_4733 (O_4733,N_49964,N_49890);
or UO_4734 (O_4734,N_49976,N_49897);
nand UO_4735 (O_4735,N_49758,N_49964);
xnor UO_4736 (O_4736,N_49808,N_49834);
and UO_4737 (O_4737,N_49847,N_49821);
or UO_4738 (O_4738,N_49802,N_49789);
and UO_4739 (O_4739,N_49807,N_49770);
or UO_4740 (O_4740,N_49940,N_49752);
nand UO_4741 (O_4741,N_49859,N_49958);
nor UO_4742 (O_4742,N_49921,N_49842);
nand UO_4743 (O_4743,N_49951,N_49946);
or UO_4744 (O_4744,N_49958,N_49844);
and UO_4745 (O_4745,N_49867,N_49878);
nor UO_4746 (O_4746,N_49818,N_49962);
nor UO_4747 (O_4747,N_49892,N_49963);
or UO_4748 (O_4748,N_49806,N_49753);
or UO_4749 (O_4749,N_49934,N_49810);
nand UO_4750 (O_4750,N_49913,N_49762);
nand UO_4751 (O_4751,N_49994,N_49803);
nand UO_4752 (O_4752,N_49807,N_49918);
xnor UO_4753 (O_4753,N_49926,N_49836);
and UO_4754 (O_4754,N_49754,N_49823);
xnor UO_4755 (O_4755,N_49813,N_49871);
or UO_4756 (O_4756,N_49873,N_49805);
nand UO_4757 (O_4757,N_49849,N_49893);
or UO_4758 (O_4758,N_49997,N_49894);
nor UO_4759 (O_4759,N_49779,N_49785);
nand UO_4760 (O_4760,N_49938,N_49843);
and UO_4761 (O_4761,N_49856,N_49984);
nand UO_4762 (O_4762,N_49809,N_49933);
or UO_4763 (O_4763,N_49990,N_49923);
xor UO_4764 (O_4764,N_49864,N_49807);
or UO_4765 (O_4765,N_49837,N_49869);
nand UO_4766 (O_4766,N_49820,N_49992);
nor UO_4767 (O_4767,N_49910,N_49989);
xnor UO_4768 (O_4768,N_49949,N_49847);
nor UO_4769 (O_4769,N_49948,N_49758);
nand UO_4770 (O_4770,N_49785,N_49815);
or UO_4771 (O_4771,N_49866,N_49816);
nor UO_4772 (O_4772,N_49943,N_49931);
xnor UO_4773 (O_4773,N_49944,N_49807);
nand UO_4774 (O_4774,N_49999,N_49955);
or UO_4775 (O_4775,N_49783,N_49965);
xnor UO_4776 (O_4776,N_49824,N_49859);
and UO_4777 (O_4777,N_49910,N_49897);
xnor UO_4778 (O_4778,N_49988,N_49973);
and UO_4779 (O_4779,N_49965,N_49809);
nand UO_4780 (O_4780,N_49943,N_49752);
and UO_4781 (O_4781,N_49875,N_49807);
nand UO_4782 (O_4782,N_49756,N_49867);
and UO_4783 (O_4783,N_49755,N_49829);
or UO_4784 (O_4784,N_49817,N_49908);
and UO_4785 (O_4785,N_49950,N_49850);
or UO_4786 (O_4786,N_49967,N_49801);
and UO_4787 (O_4787,N_49757,N_49807);
and UO_4788 (O_4788,N_49986,N_49846);
and UO_4789 (O_4789,N_49941,N_49865);
nand UO_4790 (O_4790,N_49758,N_49993);
and UO_4791 (O_4791,N_49878,N_49906);
and UO_4792 (O_4792,N_49773,N_49763);
or UO_4793 (O_4793,N_49772,N_49778);
or UO_4794 (O_4794,N_49879,N_49813);
or UO_4795 (O_4795,N_49763,N_49877);
nor UO_4796 (O_4796,N_49828,N_49816);
nor UO_4797 (O_4797,N_49953,N_49756);
and UO_4798 (O_4798,N_49923,N_49954);
xor UO_4799 (O_4799,N_49759,N_49822);
nand UO_4800 (O_4800,N_49915,N_49874);
nand UO_4801 (O_4801,N_49765,N_49963);
xnor UO_4802 (O_4802,N_49774,N_49836);
nand UO_4803 (O_4803,N_49931,N_49793);
and UO_4804 (O_4804,N_49870,N_49759);
or UO_4805 (O_4805,N_49858,N_49770);
and UO_4806 (O_4806,N_49923,N_49805);
nand UO_4807 (O_4807,N_49784,N_49965);
nand UO_4808 (O_4808,N_49898,N_49821);
and UO_4809 (O_4809,N_49751,N_49889);
or UO_4810 (O_4810,N_49963,N_49919);
and UO_4811 (O_4811,N_49859,N_49750);
xor UO_4812 (O_4812,N_49756,N_49920);
or UO_4813 (O_4813,N_49890,N_49946);
xor UO_4814 (O_4814,N_49917,N_49919);
nor UO_4815 (O_4815,N_49934,N_49764);
and UO_4816 (O_4816,N_49800,N_49900);
xnor UO_4817 (O_4817,N_49898,N_49862);
xor UO_4818 (O_4818,N_49844,N_49755);
xor UO_4819 (O_4819,N_49872,N_49960);
and UO_4820 (O_4820,N_49893,N_49940);
xnor UO_4821 (O_4821,N_49779,N_49880);
nor UO_4822 (O_4822,N_49997,N_49919);
nand UO_4823 (O_4823,N_49783,N_49974);
nand UO_4824 (O_4824,N_49896,N_49800);
and UO_4825 (O_4825,N_49812,N_49871);
nor UO_4826 (O_4826,N_49917,N_49991);
xor UO_4827 (O_4827,N_49907,N_49866);
or UO_4828 (O_4828,N_49783,N_49948);
xnor UO_4829 (O_4829,N_49948,N_49803);
xor UO_4830 (O_4830,N_49893,N_49859);
nor UO_4831 (O_4831,N_49869,N_49940);
and UO_4832 (O_4832,N_49803,N_49983);
xnor UO_4833 (O_4833,N_49870,N_49966);
and UO_4834 (O_4834,N_49762,N_49817);
or UO_4835 (O_4835,N_49880,N_49836);
and UO_4836 (O_4836,N_49957,N_49762);
nor UO_4837 (O_4837,N_49795,N_49757);
or UO_4838 (O_4838,N_49790,N_49939);
nor UO_4839 (O_4839,N_49780,N_49763);
nand UO_4840 (O_4840,N_49931,N_49964);
xnor UO_4841 (O_4841,N_49861,N_49806);
or UO_4842 (O_4842,N_49966,N_49913);
or UO_4843 (O_4843,N_49831,N_49893);
or UO_4844 (O_4844,N_49818,N_49785);
nor UO_4845 (O_4845,N_49905,N_49855);
and UO_4846 (O_4846,N_49883,N_49957);
xor UO_4847 (O_4847,N_49801,N_49989);
nand UO_4848 (O_4848,N_49784,N_49876);
nor UO_4849 (O_4849,N_49947,N_49802);
and UO_4850 (O_4850,N_49847,N_49925);
nand UO_4851 (O_4851,N_49933,N_49855);
and UO_4852 (O_4852,N_49930,N_49826);
nor UO_4853 (O_4853,N_49947,N_49967);
nand UO_4854 (O_4854,N_49948,N_49914);
and UO_4855 (O_4855,N_49912,N_49796);
and UO_4856 (O_4856,N_49772,N_49951);
xor UO_4857 (O_4857,N_49795,N_49871);
nor UO_4858 (O_4858,N_49995,N_49927);
and UO_4859 (O_4859,N_49781,N_49993);
nand UO_4860 (O_4860,N_49850,N_49928);
nand UO_4861 (O_4861,N_49955,N_49897);
or UO_4862 (O_4862,N_49873,N_49795);
nor UO_4863 (O_4863,N_49848,N_49830);
or UO_4864 (O_4864,N_49895,N_49909);
or UO_4865 (O_4865,N_49996,N_49870);
nor UO_4866 (O_4866,N_49928,N_49886);
xor UO_4867 (O_4867,N_49792,N_49911);
and UO_4868 (O_4868,N_49782,N_49929);
or UO_4869 (O_4869,N_49979,N_49965);
nand UO_4870 (O_4870,N_49780,N_49853);
and UO_4871 (O_4871,N_49782,N_49877);
xnor UO_4872 (O_4872,N_49894,N_49797);
nor UO_4873 (O_4873,N_49885,N_49810);
nor UO_4874 (O_4874,N_49921,N_49850);
nor UO_4875 (O_4875,N_49793,N_49977);
nor UO_4876 (O_4876,N_49842,N_49763);
xor UO_4877 (O_4877,N_49992,N_49977);
nor UO_4878 (O_4878,N_49756,N_49795);
nand UO_4879 (O_4879,N_49789,N_49766);
xor UO_4880 (O_4880,N_49933,N_49937);
xnor UO_4881 (O_4881,N_49893,N_49968);
and UO_4882 (O_4882,N_49937,N_49918);
or UO_4883 (O_4883,N_49875,N_49759);
nor UO_4884 (O_4884,N_49914,N_49967);
nand UO_4885 (O_4885,N_49924,N_49754);
nor UO_4886 (O_4886,N_49999,N_49873);
or UO_4887 (O_4887,N_49973,N_49796);
and UO_4888 (O_4888,N_49788,N_49900);
or UO_4889 (O_4889,N_49878,N_49975);
nor UO_4890 (O_4890,N_49784,N_49923);
or UO_4891 (O_4891,N_49817,N_49803);
nand UO_4892 (O_4892,N_49791,N_49940);
and UO_4893 (O_4893,N_49935,N_49830);
or UO_4894 (O_4894,N_49961,N_49882);
nand UO_4895 (O_4895,N_49837,N_49877);
xor UO_4896 (O_4896,N_49849,N_49872);
xnor UO_4897 (O_4897,N_49946,N_49863);
nor UO_4898 (O_4898,N_49951,N_49913);
nor UO_4899 (O_4899,N_49906,N_49779);
or UO_4900 (O_4900,N_49812,N_49982);
nand UO_4901 (O_4901,N_49876,N_49855);
or UO_4902 (O_4902,N_49843,N_49949);
nand UO_4903 (O_4903,N_49876,N_49889);
nor UO_4904 (O_4904,N_49893,N_49917);
and UO_4905 (O_4905,N_49853,N_49819);
or UO_4906 (O_4906,N_49906,N_49780);
or UO_4907 (O_4907,N_49786,N_49911);
and UO_4908 (O_4908,N_49793,N_49921);
xnor UO_4909 (O_4909,N_49787,N_49804);
xnor UO_4910 (O_4910,N_49777,N_49792);
nand UO_4911 (O_4911,N_49929,N_49781);
nand UO_4912 (O_4912,N_49998,N_49827);
nor UO_4913 (O_4913,N_49994,N_49952);
nand UO_4914 (O_4914,N_49921,N_49787);
or UO_4915 (O_4915,N_49813,N_49799);
or UO_4916 (O_4916,N_49933,N_49917);
nor UO_4917 (O_4917,N_49923,N_49950);
nand UO_4918 (O_4918,N_49971,N_49967);
and UO_4919 (O_4919,N_49905,N_49897);
and UO_4920 (O_4920,N_49994,N_49849);
nand UO_4921 (O_4921,N_49945,N_49763);
nor UO_4922 (O_4922,N_49959,N_49843);
and UO_4923 (O_4923,N_49832,N_49878);
nand UO_4924 (O_4924,N_49984,N_49798);
and UO_4925 (O_4925,N_49913,N_49967);
and UO_4926 (O_4926,N_49878,N_49853);
nor UO_4927 (O_4927,N_49831,N_49792);
nand UO_4928 (O_4928,N_49826,N_49783);
nor UO_4929 (O_4929,N_49776,N_49967);
nor UO_4930 (O_4930,N_49893,N_49988);
nor UO_4931 (O_4931,N_49867,N_49957);
nor UO_4932 (O_4932,N_49839,N_49794);
or UO_4933 (O_4933,N_49805,N_49956);
xor UO_4934 (O_4934,N_49869,N_49975);
nand UO_4935 (O_4935,N_49878,N_49810);
or UO_4936 (O_4936,N_49785,N_49983);
nor UO_4937 (O_4937,N_49790,N_49873);
or UO_4938 (O_4938,N_49994,N_49885);
xnor UO_4939 (O_4939,N_49787,N_49762);
xor UO_4940 (O_4940,N_49954,N_49811);
or UO_4941 (O_4941,N_49990,N_49956);
and UO_4942 (O_4942,N_49823,N_49800);
nor UO_4943 (O_4943,N_49961,N_49781);
nand UO_4944 (O_4944,N_49894,N_49999);
and UO_4945 (O_4945,N_49797,N_49800);
xnor UO_4946 (O_4946,N_49941,N_49778);
nor UO_4947 (O_4947,N_49984,N_49858);
or UO_4948 (O_4948,N_49916,N_49799);
xor UO_4949 (O_4949,N_49756,N_49770);
xor UO_4950 (O_4950,N_49761,N_49956);
nand UO_4951 (O_4951,N_49801,N_49762);
xnor UO_4952 (O_4952,N_49945,N_49845);
or UO_4953 (O_4953,N_49778,N_49925);
or UO_4954 (O_4954,N_49807,N_49869);
and UO_4955 (O_4955,N_49895,N_49859);
xnor UO_4956 (O_4956,N_49977,N_49998);
nand UO_4957 (O_4957,N_49987,N_49915);
nor UO_4958 (O_4958,N_49861,N_49761);
nor UO_4959 (O_4959,N_49976,N_49875);
xor UO_4960 (O_4960,N_49883,N_49817);
or UO_4961 (O_4961,N_49882,N_49765);
xnor UO_4962 (O_4962,N_49910,N_49923);
nor UO_4963 (O_4963,N_49777,N_49775);
nor UO_4964 (O_4964,N_49943,N_49877);
xnor UO_4965 (O_4965,N_49895,N_49807);
nor UO_4966 (O_4966,N_49924,N_49762);
xnor UO_4967 (O_4967,N_49861,N_49871);
nor UO_4968 (O_4968,N_49923,N_49938);
nand UO_4969 (O_4969,N_49933,N_49832);
nor UO_4970 (O_4970,N_49991,N_49801);
xnor UO_4971 (O_4971,N_49904,N_49810);
and UO_4972 (O_4972,N_49995,N_49853);
and UO_4973 (O_4973,N_49819,N_49807);
nand UO_4974 (O_4974,N_49828,N_49814);
or UO_4975 (O_4975,N_49844,N_49995);
nor UO_4976 (O_4976,N_49911,N_49927);
xor UO_4977 (O_4977,N_49920,N_49818);
nor UO_4978 (O_4978,N_49778,N_49872);
xor UO_4979 (O_4979,N_49874,N_49779);
or UO_4980 (O_4980,N_49838,N_49942);
nand UO_4981 (O_4981,N_49816,N_49898);
nand UO_4982 (O_4982,N_49980,N_49844);
or UO_4983 (O_4983,N_49941,N_49871);
nor UO_4984 (O_4984,N_49878,N_49978);
xor UO_4985 (O_4985,N_49847,N_49759);
nor UO_4986 (O_4986,N_49915,N_49866);
xnor UO_4987 (O_4987,N_49922,N_49893);
nor UO_4988 (O_4988,N_49936,N_49896);
and UO_4989 (O_4989,N_49934,N_49875);
nor UO_4990 (O_4990,N_49931,N_49794);
xnor UO_4991 (O_4991,N_49827,N_49912);
nor UO_4992 (O_4992,N_49900,N_49821);
or UO_4993 (O_4993,N_49958,N_49927);
nor UO_4994 (O_4994,N_49943,N_49759);
nand UO_4995 (O_4995,N_49846,N_49852);
xor UO_4996 (O_4996,N_49887,N_49790);
or UO_4997 (O_4997,N_49871,N_49984);
xnor UO_4998 (O_4998,N_49777,N_49852);
or UO_4999 (O_4999,N_49798,N_49758);
endmodule