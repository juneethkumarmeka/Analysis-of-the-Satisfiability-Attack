module basic_2500_25000_3000_5_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_607,In_1790);
nand U1 (N_1,In_806,In_1020);
nand U2 (N_2,In_220,In_1886);
xnor U3 (N_3,In_92,In_911);
and U4 (N_4,In_644,In_395);
nand U5 (N_5,In_1255,In_889);
nand U6 (N_6,In_1594,In_590);
and U7 (N_7,In_693,In_1172);
or U8 (N_8,In_1111,In_13);
nand U9 (N_9,In_198,In_379);
nor U10 (N_10,In_1998,In_652);
nand U11 (N_11,In_1977,In_1689);
or U12 (N_12,In_1694,In_879);
and U13 (N_13,In_1713,In_1603);
and U14 (N_14,In_859,In_1029);
or U15 (N_15,In_2335,In_144);
nor U16 (N_16,In_2403,In_2427);
or U17 (N_17,In_1753,In_417);
xnor U18 (N_18,In_1884,In_172);
xnor U19 (N_19,In_1326,In_545);
xnor U20 (N_20,In_2434,In_1641);
and U21 (N_21,In_1631,In_360);
and U22 (N_22,In_355,In_1161);
and U23 (N_23,In_118,In_2375);
and U24 (N_24,In_840,In_2090);
nor U25 (N_25,In_527,In_1692);
nand U26 (N_26,In_2162,In_737);
xnor U27 (N_27,In_622,In_839);
and U28 (N_28,In_59,In_194);
and U29 (N_29,In_812,In_1240);
nor U30 (N_30,In_1916,In_305);
nor U31 (N_31,In_2017,In_209);
xnor U32 (N_32,In_913,In_1218);
or U33 (N_33,In_1460,In_2024);
xnor U34 (N_34,In_82,In_1080);
nand U35 (N_35,In_1992,In_893);
nand U36 (N_36,In_797,In_106);
xor U37 (N_37,In_1438,In_6);
or U38 (N_38,In_1766,In_2059);
and U39 (N_39,In_555,In_1173);
xnor U40 (N_40,In_566,In_1510);
xor U41 (N_41,In_272,In_1138);
nor U42 (N_42,In_2450,In_727);
xnor U43 (N_43,In_1671,In_1423);
nor U44 (N_44,In_427,In_2301);
nand U45 (N_45,In_618,In_2094);
xor U46 (N_46,In_1588,In_139);
xnor U47 (N_47,In_562,In_474);
xor U48 (N_48,In_1368,In_1182);
and U49 (N_49,In_1573,In_621);
nand U50 (N_50,In_179,In_1527);
xor U51 (N_51,In_2231,In_1842);
and U52 (N_52,In_1462,In_1150);
or U53 (N_53,In_270,In_1476);
xor U54 (N_54,In_2440,In_1523);
nor U55 (N_55,In_1037,In_2068);
xnor U56 (N_56,In_479,In_2437);
nand U57 (N_57,In_2001,In_196);
or U58 (N_58,In_809,In_1880);
nor U59 (N_59,In_292,In_1890);
nand U60 (N_60,In_1968,In_698);
nor U61 (N_61,In_1467,In_192);
and U62 (N_62,In_2370,In_1762);
xnor U63 (N_63,In_1204,In_1958);
nand U64 (N_64,In_1908,In_2239);
and U65 (N_65,In_959,In_1373);
and U66 (N_66,In_154,In_1954);
nor U67 (N_67,In_313,In_21);
or U68 (N_68,In_1948,In_1714);
nand U69 (N_69,In_1291,In_2291);
xnor U70 (N_70,In_447,In_814);
nor U71 (N_71,In_359,In_1817);
nor U72 (N_72,In_707,In_1961);
nand U73 (N_73,In_764,In_1361);
and U74 (N_74,In_132,In_1508);
xor U75 (N_75,In_356,In_964);
nor U76 (N_76,In_1096,In_2117);
nor U77 (N_77,In_925,In_1823);
nand U78 (N_78,In_1385,In_1808);
nor U79 (N_79,In_1678,In_51);
nand U80 (N_80,In_1261,In_1016);
nand U81 (N_81,In_1760,In_967);
or U82 (N_82,In_1354,In_1412);
or U83 (N_83,In_300,In_941);
xnor U84 (N_84,In_1820,In_960);
nor U85 (N_85,In_1146,In_2438);
and U86 (N_86,In_1101,In_1801);
nand U87 (N_87,In_1128,In_1792);
xnor U88 (N_88,In_1976,In_467);
and U89 (N_89,In_1812,In_1562);
xor U90 (N_90,In_931,In_884);
xnor U91 (N_91,In_2246,In_1468);
and U92 (N_92,In_1337,In_2148);
nor U93 (N_93,In_469,In_1089);
or U94 (N_94,In_1061,In_483);
xor U95 (N_95,In_2142,In_748);
or U96 (N_96,In_1439,In_643);
xor U97 (N_97,In_1814,In_749);
and U98 (N_98,In_337,In_244);
and U99 (N_99,In_181,In_2075);
and U100 (N_100,In_1800,In_902);
xor U101 (N_101,In_1860,In_1311);
nand U102 (N_102,In_2421,In_150);
nand U103 (N_103,In_1127,In_1033);
or U104 (N_104,In_1498,In_369);
and U105 (N_105,In_2460,In_391);
nand U106 (N_106,In_890,In_1009);
and U107 (N_107,In_1421,In_325);
xnor U108 (N_108,In_1899,In_2404);
nor U109 (N_109,In_1684,In_821);
nor U110 (N_110,In_920,In_824);
or U111 (N_111,In_938,In_668);
nand U112 (N_112,In_431,In_2402);
nand U113 (N_113,In_1153,In_275);
xnor U114 (N_114,In_2235,In_1879);
xnor U115 (N_115,In_1515,In_2369);
nand U116 (N_116,In_1489,In_145);
nand U117 (N_117,In_1869,In_2425);
or U118 (N_118,In_531,In_974);
xor U119 (N_119,In_1268,In_1363);
nor U120 (N_120,In_1565,In_1491);
xnor U121 (N_121,In_1953,In_1608);
nand U122 (N_122,In_1630,In_1873);
nor U123 (N_123,In_1551,In_2385);
or U124 (N_124,In_2398,In_9);
xor U125 (N_125,In_567,In_745);
or U126 (N_126,In_757,In_301);
nand U127 (N_127,In_1446,In_1648);
or U128 (N_128,In_2222,In_532);
xnor U129 (N_129,In_684,In_1081);
nor U130 (N_130,In_278,In_2112);
nand U131 (N_131,In_58,In_250);
xor U132 (N_132,In_947,In_1169);
and U133 (N_133,In_682,In_2061);
xnor U134 (N_134,In_1633,In_1442);
xor U135 (N_135,In_1226,In_171);
nor U136 (N_136,In_1050,In_2417);
xor U137 (N_137,In_719,In_2035);
nand U138 (N_138,In_1465,In_239);
nand U139 (N_139,In_1095,In_731);
xnor U140 (N_140,In_2359,In_819);
xor U141 (N_141,In_38,In_783);
nor U142 (N_142,In_1358,In_559);
and U143 (N_143,In_1167,In_1160);
nor U144 (N_144,In_1207,In_1286);
nor U145 (N_145,In_1166,In_1698);
or U146 (N_146,In_1712,In_1872);
and U147 (N_147,In_213,In_2211);
nand U148 (N_148,In_2317,In_1148);
xor U149 (N_149,In_1735,In_1816);
nor U150 (N_150,In_1829,In_217);
or U151 (N_151,In_579,In_1939);
nor U152 (N_152,In_1509,In_86);
nor U153 (N_153,In_1942,In_414);
and U154 (N_154,In_1856,In_695);
xnor U155 (N_155,In_1092,In_357);
xnor U156 (N_156,In_1934,In_1659);
and U157 (N_157,In_1483,In_97);
nand U158 (N_158,In_1564,In_2092);
nand U159 (N_159,In_1568,In_1099);
or U160 (N_160,In_16,In_2120);
nand U161 (N_161,In_124,In_2210);
or U162 (N_162,In_113,In_1691);
or U163 (N_163,In_976,In_1929);
or U164 (N_164,In_2049,In_415);
xor U165 (N_165,In_2103,In_2178);
and U166 (N_166,In_1068,In_587);
nand U167 (N_167,In_956,In_766);
nand U168 (N_168,In_1120,In_2319);
and U169 (N_169,In_2000,In_625);
or U170 (N_170,In_2444,In_1521);
or U171 (N_171,In_324,In_768);
nand U172 (N_172,In_219,In_221);
and U173 (N_173,In_787,In_1482);
nor U174 (N_174,In_413,In_1711);
nand U175 (N_175,In_1485,In_1918);
or U176 (N_176,In_1821,In_2029);
xnor U177 (N_177,In_2048,In_2219);
xnor U178 (N_178,In_1021,In_2127);
nand U179 (N_179,In_680,In_2253);
xor U180 (N_180,In_1676,In_384);
xnor U181 (N_181,In_2153,In_810);
or U182 (N_182,In_1355,In_230);
xor U183 (N_183,In_1357,In_461);
nor U184 (N_184,In_1706,In_1771);
nand U185 (N_185,In_1078,In_1528);
and U186 (N_186,In_1619,In_1827);
or U187 (N_187,In_2361,In_282);
nor U188 (N_188,In_1310,In_1846);
nor U189 (N_189,In_2135,In_342);
xor U190 (N_190,In_1212,In_1917);
nor U191 (N_191,In_23,In_1674);
nor U192 (N_192,In_267,In_1947);
nor U193 (N_193,In_481,In_310);
or U194 (N_194,In_1071,In_560);
nor U195 (N_195,In_442,In_463);
and U196 (N_196,In_1470,In_283);
nor U197 (N_197,In_492,In_1469);
xnor U198 (N_198,In_2078,In_362);
nand U199 (N_199,In_1333,In_591);
nor U200 (N_200,In_1404,In_1459);
nand U201 (N_201,In_1072,In_1795);
and U202 (N_202,In_1539,In_677);
and U203 (N_203,In_233,In_99);
or U204 (N_204,In_1,In_2464);
or U205 (N_205,In_999,In_2028);
or U206 (N_206,In_1230,In_2077);
and U207 (N_207,In_2489,In_1253);
and U208 (N_208,In_571,In_4);
xor U209 (N_209,In_1054,In_1013);
nand U210 (N_210,In_226,In_436);
or U211 (N_211,In_1654,In_898);
nor U212 (N_212,In_844,In_1126);
nor U213 (N_213,In_1436,In_27);
and U214 (N_214,In_1930,In_249);
or U215 (N_215,In_1875,In_770);
or U216 (N_216,In_491,In_550);
xnor U217 (N_217,In_1964,In_936);
or U218 (N_218,In_174,In_2108);
nand U219 (N_219,In_1598,In_830);
nor U220 (N_220,In_261,In_1466);
and U221 (N_221,In_248,In_374);
xnor U222 (N_222,In_2129,In_437);
and U223 (N_223,In_1955,In_1755);
and U224 (N_224,In_1191,In_441);
nor U225 (N_225,In_1116,In_2229);
nor U226 (N_226,In_1220,In_1962);
nor U227 (N_227,In_2083,In_1904);
xor U228 (N_228,In_2188,In_2125);
or U229 (N_229,In_700,In_2259);
nand U230 (N_230,In_210,In_2151);
or U231 (N_231,In_180,In_576);
nor U232 (N_232,In_2258,In_860);
xnor U233 (N_233,In_1275,In_2388);
or U234 (N_234,In_537,In_2172);
nand U235 (N_235,In_2157,In_403);
nor U236 (N_236,In_1414,In_1301);
nor U237 (N_237,In_2080,In_1171);
or U238 (N_238,In_1536,In_2101);
and U239 (N_239,In_274,In_970);
nor U240 (N_240,In_2067,In_2303);
and U241 (N_241,In_661,In_1702);
nand U242 (N_242,In_166,In_1577);
or U243 (N_243,In_2429,In_109);
xor U244 (N_244,In_524,In_2063);
xnor U245 (N_245,In_1915,In_990);
nor U246 (N_246,In_50,In_1243);
nor U247 (N_247,In_871,In_1086);
and U248 (N_248,In_2087,In_1943);
nor U249 (N_249,In_817,In_402);
xnor U250 (N_250,In_1656,In_409);
xnor U251 (N_251,In_1923,In_259);
or U252 (N_252,In_1767,In_1234);
xor U253 (N_253,In_1062,In_1777);
xor U254 (N_254,In_1746,In_377);
or U255 (N_255,In_515,In_2128);
nand U256 (N_256,In_1710,In_1300);
nand U257 (N_257,In_2423,In_47);
nand U258 (N_258,In_1122,In_1993);
nand U259 (N_259,In_2300,In_934);
nor U260 (N_260,In_1197,In_921);
and U261 (N_261,In_43,In_1448);
nor U262 (N_262,In_123,In_2312);
nand U263 (N_263,In_1229,In_472);
and U264 (N_264,In_188,In_2478);
nor U265 (N_265,In_1883,In_1709);
nor U266 (N_266,In_1369,In_72);
nor U267 (N_267,In_853,In_279);
xnor U268 (N_268,In_1660,In_1592);
or U269 (N_269,In_1107,In_205);
nand U270 (N_270,In_1293,In_338);
and U271 (N_271,In_90,In_746);
xnor U272 (N_272,In_2256,In_1380);
nor U273 (N_273,In_1644,In_1501);
xnor U274 (N_274,In_392,In_598);
nand U275 (N_275,In_1718,In_1039);
nand U276 (N_276,In_525,In_2395);
xnor U277 (N_277,In_1497,In_743);
or U278 (N_278,In_1957,In_229);
nor U279 (N_279,In_335,In_443);
or U280 (N_280,In_1587,In_800);
nand U281 (N_281,In_1926,In_1051);
xnor U282 (N_282,In_1558,In_163);
or U283 (N_283,In_1210,In_1666);
nand U284 (N_284,In_19,In_71);
or U285 (N_285,In_1773,In_2472);
nor U286 (N_286,In_734,In_231);
nor U287 (N_287,In_613,In_364);
nor U288 (N_288,In_517,In_588);
or U289 (N_289,In_1832,In_1517);
nand U290 (N_290,In_471,In_1600);
nand U291 (N_291,In_1499,In_2147);
nand U292 (N_292,In_720,In_759);
nor U293 (N_293,In_2409,In_7);
xor U294 (N_294,In_674,In_1925);
and U295 (N_295,In_554,In_1217);
or U296 (N_296,In_1905,In_408);
or U297 (N_297,In_1305,In_77);
nor U298 (N_298,In_361,In_1208);
and U299 (N_299,In_1428,In_1833);
xor U300 (N_300,In_2072,In_2175);
nand U301 (N_301,In_168,In_1283);
and U302 (N_302,In_1487,In_862);
nor U303 (N_303,In_782,In_1403);
nand U304 (N_304,In_155,In_33);
or U305 (N_305,In_2036,In_2060);
or U306 (N_306,In_75,In_1578);
nor U307 (N_307,In_1584,In_833);
nand U308 (N_308,In_1841,In_1813);
xor U309 (N_309,In_2405,In_1077);
or U310 (N_310,In_1559,In_779);
nand U311 (N_311,In_733,In_284);
or U312 (N_312,In_2309,In_1541);
nand U313 (N_313,In_95,In_1650);
nor U314 (N_314,In_851,In_401);
nand U315 (N_315,In_1108,In_924);
nand U316 (N_316,In_1911,In_946);
nor U317 (N_317,In_983,In_183);
nand U318 (N_318,In_1110,In_2380);
xnor U319 (N_319,In_1896,In_801);
and U320 (N_320,In_1566,In_2307);
nand U321 (N_321,In_2284,In_994);
nand U322 (N_322,In_119,In_697);
xor U323 (N_323,In_1885,In_396);
or U324 (N_324,In_1567,In_1410);
and U325 (N_325,In_1511,In_32);
nor U326 (N_326,In_475,In_1049);
nand U327 (N_327,In_2226,In_1473);
nor U328 (N_328,In_892,In_1347);
or U329 (N_329,In_912,In_1325);
nor U330 (N_330,In_1242,In_573);
and U331 (N_331,In_147,In_2428);
nand U332 (N_332,In_1002,In_1944);
nand U333 (N_333,In_1149,In_1717);
nor U334 (N_334,In_2463,In_660);
and U335 (N_335,In_1209,In_2378);
and U336 (N_336,In_2170,In_1235);
and U337 (N_337,In_2293,In_2058);
and U338 (N_338,In_2089,In_1471);
xnor U339 (N_339,In_2116,In_1434);
nand U340 (N_340,In_771,In_1996);
xnor U341 (N_341,In_2313,In_751);
and U342 (N_342,In_1190,In_1854);
xor U343 (N_343,In_1290,In_2396);
nor U344 (N_344,In_1011,In_1625);
or U345 (N_345,In_286,In_786);
xnor U346 (N_346,In_796,In_1699);
and U347 (N_347,In_971,In_1774);
nor U348 (N_348,In_1927,In_1500);
or U349 (N_349,In_1323,In_2111);
nor U350 (N_350,In_997,In_923);
xor U351 (N_351,In_2011,In_662);
or U352 (N_352,In_1091,In_1835);
or U353 (N_353,In_406,In_1478);
xor U354 (N_354,In_304,In_2371);
and U355 (N_355,In_2419,In_69);
nor U356 (N_356,In_1249,In_2267);
nand U357 (N_357,In_55,In_949);
xor U358 (N_358,In_1019,In_204);
and U359 (N_359,In_1087,In_572);
nor U360 (N_360,In_404,In_1067);
nor U361 (N_361,In_1505,In_842);
nor U362 (N_362,In_1184,In_1602);
or U363 (N_363,In_741,In_2454);
nand U364 (N_364,In_2243,In_874);
nand U365 (N_365,In_1682,In_1623);
xnor U366 (N_366,In_103,In_1321);
and U367 (N_367,In_2104,In_722);
xnor U368 (N_368,In_858,In_1102);
nand U369 (N_369,In_61,In_1317);
nand U370 (N_370,In_1028,In_1507);
nand U371 (N_371,In_708,In_2353);
nand U372 (N_372,In_780,In_1740);
or U373 (N_373,In_1681,In_2456);
nand U374 (N_374,In_170,In_3);
xnor U375 (N_375,In_227,In_1940);
nand U376 (N_376,In_235,In_1533);
xor U377 (N_377,In_1607,In_1806);
xnor U378 (N_378,In_2121,In_1481);
nand U379 (N_379,In_616,In_1308);
or U380 (N_380,In_49,In_1141);
xor U381 (N_381,In_1583,In_1553);
nor U382 (N_382,In_314,In_1134);
xnor U383 (N_383,In_1315,In_2411);
xor U384 (N_384,In_493,In_679);
nor U385 (N_385,In_433,In_683);
and U386 (N_386,In_1552,In_1259);
xor U387 (N_387,In_280,In_189);
nor U388 (N_388,In_1341,In_928);
nand U389 (N_389,In_2206,In_1895);
and U390 (N_390,In_888,In_2110);
and U391 (N_391,In_1661,In_2399);
xnor U392 (N_392,In_1012,In_52);
nor U393 (N_393,In_1647,In_2469);
nand U394 (N_394,In_2299,In_1165);
or U395 (N_395,In_987,In_548);
or U396 (N_396,In_813,In_1636);
nand U397 (N_397,In_1722,In_1272);
and U398 (N_398,In_1180,In_240);
nand U399 (N_399,In_1254,In_629);
or U400 (N_400,In_916,In_444);
nor U401 (N_401,In_758,In_1335);
xor U402 (N_402,In_1512,In_482);
xor U403 (N_403,In_659,In_666);
or U404 (N_404,In_2288,In_2123);
xnor U405 (N_405,In_2362,In_1398);
nand U406 (N_406,In_829,In_85);
nor U407 (N_407,In_637,In_1857);
or U408 (N_408,In_825,In_1237);
xor U409 (N_409,In_2114,In_2187);
nor U410 (N_410,In_1973,In_608);
nor U411 (N_411,In_1529,In_2273);
nor U412 (N_412,In_728,In_141);
nand U413 (N_413,In_1267,In_1725);
xor U414 (N_414,In_2167,In_1838);
nor U415 (N_415,In_701,In_464);
and U416 (N_416,In_378,In_1601);
nand U417 (N_417,In_232,In_1745);
nor U418 (N_418,In_1822,In_945);
xor U419 (N_419,In_1383,In_2248);
xor U420 (N_420,In_1309,In_381);
nand U421 (N_421,In_116,In_2071);
and U422 (N_422,In_1131,In_1922);
and U423 (N_423,In_316,In_2037);
xnor U424 (N_424,In_615,In_2333);
or U425 (N_425,In_2155,In_803);
or U426 (N_426,In_339,In_2455);
and U427 (N_427,In_1324,In_162);
and U428 (N_428,In_1549,In_117);
or U429 (N_429,In_1495,In_1667);
and U430 (N_430,In_958,In_866);
and U431 (N_431,In_295,In_1595);
xor U432 (N_432,In_789,In_729);
and U433 (N_433,In_1910,In_838);
nor U434 (N_434,In_744,In_1280);
nand U435 (N_435,In_2384,In_1130);
xnor U436 (N_436,In_1085,In_1359);
and U437 (N_437,In_1177,In_1336);
nand U438 (N_438,In_142,In_647);
nor U439 (N_439,In_136,In_1298);
and U440 (N_440,In_405,In_1544);
or U441 (N_441,In_557,In_28);
nand U442 (N_442,In_2325,In_306);
or U443 (N_443,In_1036,In_687);
nand U444 (N_444,In_1959,In_1990);
and U445 (N_445,In_2480,In_1859);
and U446 (N_446,In_1024,In_1479);
and U447 (N_447,In_320,In_2485);
and U448 (N_448,In_1979,In_1213);
and U449 (N_449,In_614,In_508);
nor U450 (N_450,In_539,In_25);
and U451 (N_451,In_1391,In_1981);
and U452 (N_452,In_952,In_2373);
nand U453 (N_453,In_1787,In_247);
and U454 (N_454,In_2287,In_2466);
or U455 (N_455,In_1646,In_792);
nand U456 (N_456,In_2199,In_484);
nor U457 (N_457,In_955,In_1431);
nor U458 (N_458,In_2310,In_1727);
nor U459 (N_459,In_238,In_108);
nor U460 (N_460,In_1198,In_1450);
and U461 (N_461,In_594,In_2021);
nor U462 (N_462,In_658,In_1451);
and U463 (N_463,In_46,In_293);
or U464 (N_464,In_1728,In_1464);
nor U465 (N_465,In_2131,In_702);
xor U466 (N_466,In_2368,In_1375);
nor U467 (N_467,In_585,In_756);
or U468 (N_468,In_2013,In_2230);
nor U469 (N_469,In_2462,In_2073);
and U470 (N_470,In_981,In_856);
xnor U471 (N_471,In_380,In_826);
and U472 (N_472,In_1965,In_2415);
nand U473 (N_473,In_1258,In_937);
nor U474 (N_474,In_1804,In_1840);
or U475 (N_475,In_1420,In_2130);
or U476 (N_476,In_143,In_1117);
or U477 (N_477,In_635,In_1989);
or U478 (N_478,In_129,In_961);
nand U479 (N_479,In_1794,In_1613);
xnor U480 (N_480,In_399,In_1339);
and U481 (N_481,In_1991,In_2268);
or U482 (N_482,In_445,In_513);
or U483 (N_483,In_299,In_2420);
nor U484 (N_484,In_977,In_1704);
nand U485 (N_485,In_775,In_78);
nor U486 (N_486,In_2053,In_966);
nand U487 (N_487,In_2099,In_1986);
nand U488 (N_488,In_1247,In_896);
and U489 (N_489,In_1316,In_907);
or U490 (N_490,In_257,In_939);
or U491 (N_491,In_182,In_1027);
and U492 (N_492,In_915,In_1901);
nand U493 (N_493,In_1271,In_735);
nand U494 (N_494,In_847,In_452);
nor U495 (N_495,In_2347,In_1152);
nand U496 (N_496,In_1007,In_91);
xnor U497 (N_497,In_2134,In_1532);
or U498 (N_498,In_289,In_2326);
nand U499 (N_499,In_953,In_2198);
and U500 (N_500,In_1980,In_899);
nand U501 (N_501,In_1651,In_1673);
or U502 (N_502,In_2144,In_1045);
nand U503 (N_503,In_37,In_1069);
nand U504 (N_504,In_135,In_715);
and U505 (N_505,In_430,In_1778);
nand U506 (N_506,In_1294,In_1256);
xnor U507 (N_507,In_623,In_1852);
nor U508 (N_508,In_327,In_506);
and U509 (N_509,In_965,In_691);
and U510 (N_510,In_843,In_1265);
xor U511 (N_511,In_1724,In_1189);
and U512 (N_512,In_1589,In_241);
and U513 (N_513,In_1845,In_2336);
and U514 (N_514,In_2193,In_1987);
xnor U515 (N_515,In_1836,In_717);
xor U516 (N_516,In_2047,In_2493);
xnor U517 (N_517,In_2088,In_2424);
or U518 (N_518,In_1893,In_1297);
and U519 (N_519,In_1006,In_1737);
nand U520 (N_520,In_505,In_863);
xnor U521 (N_521,In_1731,In_252);
xnor U522 (N_522,In_1877,In_2497);
nor U523 (N_523,In_185,In_564);
and U524 (N_524,In_940,In_2171);
or U525 (N_525,In_2100,In_45);
or U526 (N_526,In_954,In_64);
xnor U527 (N_527,In_2311,In_1252);
nor U528 (N_528,In_1983,In_1455);
or U529 (N_529,In_487,In_1867);
nand U530 (N_530,In_638,In_2194);
and U531 (N_531,In_112,In_602);
and U532 (N_532,In_2449,In_1227);
and U533 (N_533,In_1312,In_1221);
and U534 (N_534,In_1570,In_561);
nand U535 (N_535,In_1395,In_1585);
nor U536 (N_536,In_2394,In_2446);
nand U537 (N_537,In_1605,In_1104);
or U538 (N_538,In_1394,In_1032);
and U539 (N_539,In_1035,In_269);
nand U540 (N_540,In_930,In_114);
xnor U541 (N_541,In_536,In_1811);
and U542 (N_542,In_1534,In_122);
nor U543 (N_543,In_2279,In_2146);
xor U544 (N_544,In_2156,In_1454);
nand U545 (N_545,In_2338,In_2316);
nand U546 (N_546,In_26,In_520);
and U547 (N_547,In_1898,In_1396);
nor U548 (N_548,In_1136,In_351);
xnor U549 (N_549,In_1748,In_1304);
nand U550 (N_550,In_460,In_1984);
nand U551 (N_551,In_1582,In_656);
and U552 (N_552,In_1475,In_2260);
nand U553 (N_553,In_788,In_2124);
nand U554 (N_554,In_1417,In_126);
and U555 (N_555,In_1550,In_1397);
xor U556 (N_556,In_975,In_973);
and U557 (N_557,In_434,In_1658);
nor U558 (N_558,In_2458,In_1075);
xnor U559 (N_559,In_593,In_2366);
nor U560 (N_560,In_2250,In_1429);
xnor U561 (N_561,In_1634,In_1196);
nand U562 (N_562,In_2138,In_1518);
or U563 (N_563,In_2225,In_2341);
xor U564 (N_564,In_330,In_2498);
nand U565 (N_565,In_1502,In_79);
nor U566 (N_566,In_558,In_2018);
and U567 (N_567,In_872,In_1803);
nand U568 (N_568,In_822,In_1569);
or U569 (N_569,In_1931,In_1245);
or U570 (N_570,In_836,In_2033);
or U571 (N_571,In_1723,In_2056);
or U572 (N_572,In_1427,In_137);
nand U573 (N_573,In_578,In_2038);
xor U574 (N_574,In_918,In_102);
nand U575 (N_575,In_2050,In_2332);
or U576 (N_576,In_197,In_1044);
nor U577 (N_577,In_332,In_1616);
nand U578 (N_578,In_2292,In_2096);
or U579 (N_579,In_2228,In_1393);
nand U580 (N_580,In_1798,In_2006);
or U581 (N_581,In_942,In_849);
and U582 (N_582,In_762,In_688);
xnor U583 (N_583,In_1690,In_774);
or U584 (N_584,In_1211,In_1266);
and U585 (N_585,In_2245,In_1837);
or U586 (N_586,In_699,In_2270);
or U587 (N_587,In_1657,In_2295);
or U588 (N_588,In_2345,In_979);
nand U589 (N_589,In_2025,In_76);
or U590 (N_590,In_2247,In_2145);
and U591 (N_591,In_1381,In_905);
or U592 (N_592,In_15,In_1195);
or U593 (N_593,In_2467,In_795);
nand U594 (N_594,In_1088,In_2254);
or U595 (N_595,In_1574,In_127);
nand U596 (N_596,In_1408,In_820);
or U597 (N_597,In_721,In_1070);
or U598 (N_598,In_2190,In_904);
nand U599 (N_599,In_583,In_2183);
xnor U600 (N_600,In_1768,In_563);
or U601 (N_601,In_1338,In_619);
nand U602 (N_602,In_1178,In_2282);
and U603 (N_603,In_152,In_2214);
or U604 (N_604,In_1815,In_2278);
and U605 (N_605,In_501,In_927);
or U606 (N_606,In_258,In_1705);
or U607 (N_607,In_597,In_1364);
or U608 (N_608,In_1611,In_30);
nand U609 (N_609,In_919,In_529);
and U610 (N_610,In_456,In_827);
or U611 (N_611,In_24,In_218);
nand U612 (N_612,In_1121,In_1000);
xnor U613 (N_613,In_429,In_148);
nor U614 (N_614,In_1862,In_1118);
and U615 (N_615,In_291,In_2031);
or U616 (N_616,In_665,In_1853);
and U617 (N_617,In_1264,In_521);
xnor U618 (N_618,In_419,In_1741);
nand U619 (N_619,In_989,In_2386);
xnor U620 (N_620,In_1073,In_1525);
nand U621 (N_621,In_2499,In_0);
nor U622 (N_622,In_1972,In_1621);
xor U623 (N_623,In_211,In_2026);
nand U624 (N_624,In_2164,In_1225);
nand U625 (N_625,In_577,In_1618);
or U626 (N_626,In_1456,In_885);
and U627 (N_627,In_31,In_2457);
nor U628 (N_628,In_2391,In_2122);
or U629 (N_629,In_2351,In_393);
xor U630 (N_630,In_1769,In_2354);
or U631 (N_631,In_382,In_1575);
and U632 (N_632,In_186,In_767);
nor U633 (N_633,In_83,In_2158);
xor U634 (N_634,In_1340,In_1861);
nand U635 (N_635,In_1026,In_53);
or U636 (N_636,In_111,In_1995);
xor U637 (N_637,In_1248,In_2132);
nand U638 (N_638,In_1484,In_251);
or U639 (N_639,In_880,In_1453);
xor U640 (N_640,In_1941,In_569);
nand U641 (N_641,In_2126,In_1215);
nand U642 (N_642,In_773,In_673);
or U643 (N_643,In_1825,In_823);
and U644 (N_644,In_245,In_1683);
nor U645 (N_645,In_2358,In_1010);
nor U646 (N_646,In_1332,In_1186);
xnor U647 (N_647,In_465,In_2179);
and U648 (N_648,In_1192,In_2376);
nor U649 (N_649,In_781,In_2477);
and U650 (N_650,In_1418,In_951);
or U651 (N_651,In_1432,In_646);
or U652 (N_652,In_1906,In_1384);
nor U653 (N_653,In_1677,In_2027);
or U654 (N_654,In_2065,In_2002);
nor U655 (N_655,In_1982,In_1887);
or U656 (N_656,In_2052,In_2074);
xnor U657 (N_657,In_121,In_2109);
nand U658 (N_658,In_2383,In_1720);
nand U659 (N_659,In_664,In_2197);
or U660 (N_660,In_1571,In_207);
and U661 (N_661,In_804,In_1876);
nand U662 (N_662,In_1374,In_1530);
nor U663 (N_663,In_540,In_1156);
nor U664 (N_664,In_523,In_1376);
and U665 (N_665,In_344,In_739);
nor U666 (N_666,In_1206,In_1238);
and U667 (N_667,In_802,In_1668);
nand U668 (N_668,In_2323,In_657);
nand U669 (N_669,In_1330,In_627);
and U670 (N_670,In_519,In_1693);
nand U671 (N_671,In_1366,In_1974);
xor U672 (N_672,In_948,In_2189);
and U673 (N_673,In_589,In_1334);
nor U674 (N_674,In_932,In_478);
or U675 (N_675,In_1685,In_1458);
and U676 (N_676,In_1174,In_1865);
xnor U677 (N_677,In_1306,In_2285);
nand U678 (N_678,In_2283,In_1796);
and U679 (N_679,In_1343,In_1739);
and U680 (N_680,In_497,In_454);
or U681 (N_681,In_1703,In_2019);
xnor U682 (N_682,In_534,In_586);
nand U683 (N_683,In_1406,In_1715);
nor U684 (N_684,In_400,In_1262);
or U685 (N_685,In_841,In_2168);
nand U686 (N_686,In_1302,In_808);
and U687 (N_687,In_365,In_234);
xor U688 (N_688,In_1726,In_1747);
xnor U689 (N_689,In_689,In_2076);
or U690 (N_690,In_256,In_1834);
nand U691 (N_691,In_2496,In_1907);
xor U692 (N_692,In_1679,In_1350);
xnor U693 (N_693,In_831,In_710);
nand U694 (N_694,In_2360,In_755);
or U695 (N_695,In_832,In_1932);
nand U696 (N_696,In_1185,In_1277);
and U697 (N_697,In_1203,In_290);
nand U698 (N_698,In_988,In_2329);
or U699 (N_699,In_1219,In_1610);
and U700 (N_700,In_2304,In_169);
nand U701 (N_701,In_2085,In_2091);
and U702 (N_702,In_1236,In_1194);
xnor U703 (N_703,In_761,In_1307);
xor U704 (N_704,In_2272,In_510);
or U705 (N_705,In_547,In_633);
xnor U706 (N_706,In_617,In_321);
nand U707 (N_707,In_1850,In_1617);
nand U708 (N_708,In_886,In_1839);
nand U709 (N_709,In_476,In_326);
xnor U710 (N_710,In_1945,In_1535);
xnor U711 (N_711,In_1094,In_1556);
or U712 (N_712,In_703,In_425);
xor U713 (N_713,In_1729,In_1017);
and U714 (N_714,In_850,In_184);
nor U715 (N_715,In_2113,In_363);
or U716 (N_716,In_2034,In_329);
and U717 (N_717,In_2445,In_1750);
xor U718 (N_718,In_2340,In_1409);
nor U719 (N_719,In_2265,In_1785);
nand U720 (N_720,In_315,In_2393);
and U721 (N_721,In_2356,In_1349);
nand U722 (N_722,In_488,In_1642);
xor U723 (N_723,In_1098,In_2173);
or U724 (N_724,In_2079,In_2334);
and U725 (N_725,In_906,In_551);
and U726 (N_726,In_2069,In_496);
xnor U727 (N_727,In_570,In_2451);
or U728 (N_728,In_1132,In_1526);
xor U729 (N_729,In_2381,In_394);
xor U730 (N_730,In_969,In_65);
or U731 (N_731,In_2165,In_323);
xnor U732 (N_732,In_1545,In_312);
nand U733 (N_733,In_2294,In_1274);
nor U734 (N_734,In_848,In_1554);
and U735 (N_735,In_1319,In_1791);
xnor U736 (N_736,In_66,In_1193);
and U737 (N_737,In_1057,In_153);
and U738 (N_738,In_1670,In_1513);
nand U739 (N_739,In_1251,In_1415);
nor U740 (N_740,In_167,In_1824);
or U741 (N_741,In_2045,In_1537);
nand U742 (N_742,In_2015,In_271);
nand U743 (N_743,In_1066,In_260);
nand U744 (N_744,In_544,In_882);
xnor U745 (N_745,In_1956,In_1719);
nor U746 (N_746,In_855,In_645);
or U747 (N_747,In_798,In_765);
nor U748 (N_748,In_2004,In_2266);
xnor U749 (N_749,In_2492,In_190);
xor U750 (N_750,In_448,In_2297);
nor U751 (N_751,In_1022,In_507);
or U752 (N_752,In_176,In_1288);
or U753 (N_753,In_2486,In_747);
nor U754 (N_754,In_2461,In_1147);
and U755 (N_755,In_2084,In_908);
nor U756 (N_756,In_985,In_878);
nor U757 (N_757,In_1721,In_1579);
nand U758 (N_758,In_2296,In_502);
nand U759 (N_759,In_74,In_754);
and U760 (N_760,In_1688,In_120);
and U761 (N_761,In_173,In_2406);
xor U762 (N_762,In_328,In_317);
or U763 (N_763,In_996,In_1960);
nand U764 (N_764,In_39,In_2224);
and U765 (N_765,In_671,In_753);
xor U766 (N_766,In_1700,In_1214);
and U767 (N_767,In_2344,In_68);
nor U768 (N_768,In_477,In_1273);
nor U769 (N_769,In_1752,In_2220);
nor U770 (N_770,In_2352,In_2339);
nand U771 (N_771,In_35,In_1179);
and U772 (N_772,In_1858,In_1232);
xor U773 (N_773,In_2476,In_193);
nand U774 (N_774,In_273,In_2475);
xor U775 (N_775,In_322,In_388);
nor U776 (N_776,In_917,In_1056);
xnor U777 (N_777,In_1488,In_2184);
nor U778 (N_778,In_1496,In_962);
nand U779 (N_779,In_175,In_432);
nand U780 (N_780,In_978,In_1040);
or U781 (N_781,In_1680,In_2160);
xor U782 (N_782,In_2481,In_1951);
nand U783 (N_783,In_980,In_157);
xnor U784 (N_784,In_837,In_2479);
or U785 (N_785,In_255,In_2217);
and U786 (N_786,In_277,In_1367);
xnor U787 (N_787,In_8,In_1318);
nand U788 (N_788,In_1200,In_2261);
xnor U789 (N_789,In_2223,In_1443);
or U790 (N_790,In_963,In_1697);
and U791 (N_791,In_1843,In_1758);
nor U792 (N_792,In_867,In_1912);
or U793 (N_793,In_2263,In_1538);
or U794 (N_794,In_341,In_1866);
and U795 (N_795,In_582,In_1604);
nor U796 (N_796,In_2314,In_2412);
and U797 (N_797,In_2422,In_2276);
nor U798 (N_798,In_1924,In_1233);
nor U799 (N_799,In_992,In_1257);
or U800 (N_800,In_1937,In_1114);
xnor U801 (N_801,In_740,In_2152);
nor U802 (N_802,In_1145,In_2234);
and U803 (N_803,In_2390,In_266);
xnor U804 (N_804,In_1733,In_1743);
or U805 (N_805,In_712,In_1855);
or U806 (N_806,In_1868,In_713);
and U807 (N_807,In_1606,In_385);
and U808 (N_808,In_1162,In_1014);
xnor U809 (N_809,In_1378,In_2255);
xnor U810 (N_810,In_1201,In_1894);
and U811 (N_811,In_2014,In_2364);
or U812 (N_812,In_346,In_2020);
or U813 (N_813,In_370,In_1506);
or U814 (N_814,In_449,In_96);
and U815 (N_815,In_22,In_1100);
and U816 (N_816,In_2097,In_1155);
and U817 (N_817,In_435,In_1105);
nand U818 (N_818,In_1356,In_1643);
nand U819 (N_819,In_1749,In_1615);
and U820 (N_820,In_692,In_1493);
nor U821 (N_821,In_349,In_2046);
or U822 (N_822,In_1738,In_2169);
nor U823 (N_823,In_1047,In_1377);
nor U824 (N_824,In_1919,In_1669);
xor U825 (N_825,In_298,In_2308);
and U826 (N_826,In_1555,In_1490);
and U827 (N_827,In_1175,In_1038);
or U828 (N_828,In_2470,In_1730);
or U829 (N_829,In_48,In_653);
nand U830 (N_830,In_1831,In_2349);
nand U831 (N_831,In_495,In_1756);
nor U832 (N_832,In_489,In_2262);
nor U833 (N_833,In_922,In_606);
xor U834 (N_834,In_1362,In_1935);
and U835 (N_835,In_1520,In_2041);
xnor U836 (N_836,In_2275,In_1222);
xor U837 (N_837,In_2,In_1181);
nor U838 (N_838,In_1327,In_2441);
and U839 (N_839,In_1563,In_2216);
and U840 (N_840,In_1246,In_1614);
nor U841 (N_841,In_910,In_528);
and U842 (N_842,In_1881,In_1370);
xor U843 (N_843,In_208,In_678);
nor U844 (N_844,In_914,In_228);
nand U845 (N_845,In_543,In_2379);
xnor U846 (N_846,In_730,In_368);
nor U847 (N_847,In_732,In_1001);
nor U848 (N_848,In_900,In_2443);
nand U849 (N_849,In_1576,In_2185);
nand U850 (N_850,In_1844,In_34);
nor U851 (N_851,In_2414,In_20);
nand U852 (N_852,In_1761,In_2442);
or U853 (N_853,In_1902,In_1270);
nor U854 (N_854,In_294,In_1282);
and U855 (N_855,In_1205,In_968);
xnor U856 (N_856,In_1540,In_1387);
nor U857 (N_857,In_457,In_309);
or U858 (N_858,In_2473,In_1742);
xor U859 (N_859,In_846,In_2119);
and U860 (N_860,In_651,In_2328);
or U861 (N_861,In_1652,In_1591);
nand U862 (N_862,In_626,In_36);
and U863 (N_863,In_2453,In_2357);
nor U864 (N_864,In_929,In_1663);
nor U865 (N_865,In_2269,In_158);
and U866 (N_866,In_1142,In_340);
nand U867 (N_867,In_1672,In_14);
nand U868 (N_868,In_2102,In_1133);
and U869 (N_869,In_1407,In_2212);
nor U870 (N_870,In_752,In_490);
nand U871 (N_871,In_995,In_2070);
and U872 (N_872,In_1348,In_1920);
nand U873 (N_873,In_511,In_580);
and U874 (N_874,In_2432,In_1437);
nor U875 (N_875,In_1379,In_1422);
nand U876 (N_876,In_2487,In_2161);
or U877 (N_877,In_828,In_1653);
nor U878 (N_878,In_1952,In_1093);
or U879 (N_879,In_742,In_1351);
or U880 (N_880,In_640,In_438);
nand U881 (N_881,In_56,In_556);
and U882 (N_882,In_2318,In_1765);
nor U883 (N_883,In_685,In_2010);
and U884 (N_884,In_620,In_986);
nor U885 (N_885,In_140,In_2040);
xnor U886 (N_886,In_654,In_1163);
and U887 (N_887,In_2342,In_10);
nand U888 (N_888,In_418,In_2374);
and U889 (N_889,In_2081,In_87);
xor U890 (N_890,In_1696,In_1871);
xor U891 (N_891,In_2348,In_516);
and U892 (N_892,In_818,In_1776);
xnor U893 (N_893,In_1732,In_353);
nor U894 (N_894,In_535,In_2154);
xor U895 (N_895,In_215,In_1135);
and U896 (N_896,In_1628,In_1851);
xnor U897 (N_897,In_2435,In_624);
and U898 (N_898,In_264,In_2274);
xor U899 (N_899,In_17,In_1441);
nor U900 (N_900,In_81,In_2377);
and U901 (N_901,In_187,In_1140);
nor U902 (N_902,In_2277,In_2459);
nand U903 (N_903,In_287,In_428);
nor U904 (N_904,In_2066,In_2436);
nor U905 (N_905,In_1260,In_1516);
nor U906 (N_906,In_1284,In_485);
nand U907 (N_907,In_852,In_2430);
and U908 (N_908,In_1645,In_470);
or U909 (N_909,In_1797,In_612);
xnor U910 (N_910,In_2186,In_736);
xnor U911 (N_911,In_857,In_1278);
nor U912 (N_912,In_2166,In_63);
nor U913 (N_913,In_2474,In_1328);
nand U914 (N_914,In_546,In_861);
or U915 (N_915,In_1015,In_1313);
nand U916 (N_916,In_115,In_214);
and U917 (N_917,In_1314,In_1971);
nand U918 (N_918,In_372,In_2468);
and U919 (N_919,In_2387,In_634);
and U920 (N_920,In_1322,In_420);
and U921 (N_921,In_2343,In_1477);
xor U922 (N_922,In_599,In_319);
and U923 (N_923,In_199,In_2054);
nor U924 (N_924,In_2163,In_991);
and U925 (N_925,In_648,In_574);
nor U926 (N_926,In_2400,In_1269);
nand U927 (N_927,In_2242,In_1878);
and U928 (N_928,In_165,In_223);
nor U929 (N_929,In_1074,In_354);
nand U930 (N_930,In_2215,In_2490);
nor U931 (N_931,In_1053,In_881);
and U932 (N_932,In_1624,In_1764);
nor U933 (N_933,In_603,In_1686);
and U934 (N_934,In_29,In_1938);
nand U935 (N_935,In_1119,In_373);
xnor U936 (N_936,In_1346,In_609);
and U937 (N_937,In_641,In_161);
xor U938 (N_938,In_1780,In_1581);
xor U939 (N_939,In_1597,In_2093);
and U940 (N_940,In_2482,In_450);
nand U941 (N_941,In_302,In_73);
nand U942 (N_942,In_1928,In_2057);
xor U943 (N_943,In_1287,In_1064);
and U944 (N_944,In_984,In_2431);
or U945 (N_945,In_60,In_1848);
and U946 (N_946,In_1372,In_2252);
or U947 (N_947,In_2401,In_1041);
nand U948 (N_948,In_1168,In_2195);
or U949 (N_949,In_565,In_2177);
nand U950 (N_950,In_128,In_1426);
nor U951 (N_951,In_2062,In_1400);
and U952 (N_952,In_191,In_1199);
nand U953 (N_953,In_738,In_793);
xor U954 (N_954,In_446,In_2327);
nand U955 (N_955,In_714,In_711);
or U956 (N_956,In_2012,In_486);
xnor U957 (N_957,In_1903,In_2238);
nor U958 (N_958,In_1444,In_1411);
and U959 (N_959,In_2320,In_42);
nor U960 (N_960,In_352,In_1137);
and U961 (N_961,In_397,In_1151);
nor U962 (N_962,In_98,In_610);
nand U963 (N_963,In_2139,In_1967);
and U964 (N_964,In_1048,In_1388);
nand U965 (N_965,In_1392,In_2271);
and U966 (N_966,In_1303,In_1586);
nor U967 (N_967,In_2465,In_1994);
nand U968 (N_968,In_2003,In_750);
nand U969 (N_969,In_1139,In_366);
or U970 (N_970,In_455,In_2098);
nor U971 (N_971,In_134,In_1744);
and U972 (N_972,In_84,In_1365);
xor U973 (N_973,In_894,In_2321);
and U974 (N_974,In_1492,In_1457);
and U975 (N_975,In_935,In_281);
xnor U976 (N_976,In_1106,In_1472);
or U977 (N_977,In_2483,In_243);
nand U978 (N_978,In_347,In_67);
nand U979 (N_979,In_784,In_1548);
nand U980 (N_980,In_345,In_667);
and U981 (N_981,In_553,In_1781);
and U982 (N_982,In_2022,In_2204);
nand U983 (N_983,In_1751,In_216);
and U984 (N_984,In_1224,In_285);
nor U985 (N_985,In_2418,In_1599);
xnor U986 (N_986,In_650,In_2032);
and U987 (N_987,In_2221,In_303);
nor U988 (N_988,In_778,In_222);
xnor U989 (N_989,In_2350,In_835);
nand U990 (N_990,In_110,In_864);
nand U991 (N_991,In_675,In_1183);
and U992 (N_992,In_1695,In_1082);
or U993 (N_993,In_1590,In_131);
nor U994 (N_994,In_706,In_2150);
xor U995 (N_995,In_254,In_877);
nand U996 (N_996,In_1244,In_887);
and U997 (N_997,In_2305,In_130);
or U998 (N_998,In_1123,In_1043);
xnor U999 (N_999,In_2180,In_44);
nor U1000 (N_1000,In_1830,In_628);
and U1001 (N_1001,In_1999,In_1143);
and U1002 (N_1002,In_1416,In_632);
xor U1003 (N_1003,In_718,In_639);
and U1004 (N_1004,In_1063,In_468);
and U1005 (N_1005,In_1440,In_2023);
nor U1006 (N_1006,In_2181,In_1557);
and U1007 (N_1007,In_891,In_2392);
or U1008 (N_1008,In_1596,In_1775);
xnor U1009 (N_1009,In_1401,In_2452);
nor U1010 (N_1010,In_57,In_2264);
nand U1011 (N_1011,In_1424,In_195);
nand U1012 (N_1012,In_1084,In_1810);
or U1013 (N_1013,In_1786,In_2007);
xnor U1014 (N_1014,In_224,In_1546);
or U1015 (N_1015,In_769,In_1042);
nand U1016 (N_1016,In_777,In_1933);
nor U1017 (N_1017,In_331,In_2363);
and U1018 (N_1018,In_263,In_242);
xor U1019 (N_1019,In_512,In_799);
or U1020 (N_1020,In_1847,In_1344);
nand U1021 (N_1021,In_1030,In_202);
or U1022 (N_1022,In_1480,In_1640);
nor U1023 (N_1023,In_873,In_2484);
xor U1024 (N_1024,In_2205,In_1449);
and U1025 (N_1025,In_1687,In_541);
or U1026 (N_1026,In_2337,In_383);
xnor U1027 (N_1027,In_1701,In_605);
or U1028 (N_1028,In_549,In_1626);
nand U1029 (N_1029,In_1463,In_1083);
nor U1030 (N_1030,In_54,In_149);
or U1031 (N_1031,In_390,In_268);
nand U1032 (N_1032,In_630,In_1874);
nor U1033 (N_1033,In_201,In_1863);
nand U1034 (N_1034,In_2397,In_1946);
xor U1035 (N_1035,In_1320,In_1950);
nor U1036 (N_1036,In_499,In_1818);
xnor U1037 (N_1037,In_2064,In_297);
nand U1038 (N_1038,In_94,In_318);
xor U1039 (N_1039,In_854,In_1125);
and U1040 (N_1040,In_870,In_1514);
nand U1041 (N_1041,In_2016,In_1170);
nand U1042 (N_1042,In_514,In_2213);
xnor U1043 (N_1043,In_655,In_2286);
xnor U1044 (N_1044,In_2426,In_2005);
or U1045 (N_1045,In_1662,In_160);
nor U1046 (N_1046,In_426,In_1103);
or U1047 (N_1047,In_2218,In_1004);
nand U1048 (N_1048,In_811,In_89);
nand U1049 (N_1049,In_1144,In_705);
and U1050 (N_1050,In_458,In_1560);
nor U1051 (N_1051,In_1664,In_480);
xor U1052 (N_1052,In_1281,In_1390);
nor U1053 (N_1053,In_203,In_2095);
or U1054 (N_1054,In_1782,In_1921);
nand U1055 (N_1055,In_2009,In_1736);
xnor U1056 (N_1056,In_62,In_410);
nor U1057 (N_1057,In_2106,In_1295);
and U1058 (N_1058,In_1461,In_1352);
xor U1059 (N_1059,In_526,In_2237);
or U1060 (N_1060,In_411,In_1060);
nand U1061 (N_1061,In_2324,In_663);
xor U1062 (N_1062,In_1988,In_709);
xor U1063 (N_1063,In_1891,In_2176);
and U1064 (N_1064,In_440,In_1216);
or U1065 (N_1065,In_412,In_875);
or U1066 (N_1066,In_1793,In_957);
xor U1067 (N_1067,In_1159,In_398);
and U1068 (N_1068,In_575,In_600);
and U1069 (N_1069,In_262,In_1113);
xnor U1070 (N_1070,In_1524,In_389);
and U1071 (N_1071,In_146,In_581);
and U1072 (N_1072,In_451,In_1329);
nor U1073 (N_1073,In_1296,In_2236);
nor U1074 (N_1074,In_865,In_225);
and U1075 (N_1075,In_1870,In_1864);
and U1076 (N_1076,In_498,In_101);
or U1077 (N_1077,In_901,In_1949);
and U1078 (N_1078,In_1353,In_1772);
nor U1079 (N_1079,In_386,In_1799);
and U1080 (N_1080,In_807,In_2043);
nor U1081 (N_1081,In_2448,In_2192);
nand U1082 (N_1082,In_1109,In_1285);
or U1083 (N_1083,In_2416,In_1202);
nand U1084 (N_1084,In_595,In_1985);
nor U1085 (N_1085,In_794,In_2207);
xor U1086 (N_1086,In_1637,In_1788);
xnor U1087 (N_1087,In_177,In_1580);
xnor U1088 (N_1088,In_522,In_1649);
and U1089 (N_1089,In_1547,In_1900);
nor U1090 (N_1090,In_104,In_107);
or U1091 (N_1091,In_676,In_1176);
nor U1092 (N_1092,In_1241,In_156);
or U1093 (N_1093,In_5,In_1503);
and U1094 (N_1094,In_1978,In_237);
nor U1095 (N_1095,In_2257,In_311);
and U1096 (N_1096,In_1079,In_1627);
nand U1097 (N_1097,In_1963,In_530);
nand U1098 (N_1098,In_1008,In_933);
nor U1099 (N_1099,In_1779,In_1819);
xor U1100 (N_1100,In_2306,In_236);
or U1101 (N_1101,In_1292,In_672);
nand U1102 (N_1102,In_138,In_1445);
and U1103 (N_1103,In_845,In_1447);
and U1104 (N_1104,In_2232,In_1675);
xnor U1105 (N_1105,In_1572,In_2137);
xnor U1106 (N_1106,In_2182,In_1371);
nor U1107 (N_1107,In_1639,In_1975);
xnor U1108 (N_1108,In_2410,In_2302);
nand U1109 (N_1109,In_1188,In_376);
and U1110 (N_1110,In_12,In_2298);
and U1111 (N_1111,In_1065,In_2209);
nor U1112 (N_1112,In_1629,In_1809);
or U1113 (N_1113,In_1936,In_1784);
xnor U1114 (N_1114,In_694,In_1228);
nand U1115 (N_1115,In_2471,In_704);
and U1116 (N_1116,In_288,In_246);
or U1117 (N_1117,In_133,In_1909);
nand U1118 (N_1118,In_1826,In_125);
or U1119 (N_1119,In_2174,In_869);
xor U1120 (N_1120,In_2055,In_763);
or U1121 (N_1121,In_690,In_868);
nor U1122 (N_1122,In_1789,In_1486);
nand U1123 (N_1123,In_18,In_422);
nand U1124 (N_1124,In_88,In_2115);
xor U1125 (N_1125,In_1331,In_816);
nor U1126 (N_1126,In_1289,In_1609);
or U1127 (N_1127,In_998,In_1154);
or U1128 (N_1128,In_1805,In_1425);
nor U1129 (N_1129,In_2281,In_358);
nor U1130 (N_1130,In_307,In_2495);
or U1131 (N_1131,In_1046,In_253);
or U1132 (N_1132,In_815,In_611);
and U1133 (N_1133,In_1622,In_533);
xor U1134 (N_1134,In_1382,In_276);
nand U1135 (N_1135,In_1757,In_2346);
nor U1136 (N_1136,In_2488,In_1345);
and U1137 (N_1137,In_1018,In_336);
xnor U1138 (N_1138,In_686,In_1519);
xor U1139 (N_1139,In_1435,In_1966);
xnor U1140 (N_1140,In_2249,In_333);
nand U1141 (N_1141,In_1707,In_669);
or U1142 (N_1142,In_1997,In_1655);
nor U1143 (N_1143,In_1969,In_1115);
nand U1144 (N_1144,In_897,In_584);
or U1145 (N_1145,In_462,In_1076);
and U1146 (N_1146,In_2389,In_926);
and U1147 (N_1147,In_1754,In_387);
or U1148 (N_1148,In_883,In_1389);
nand U1149 (N_1149,In_2240,In_1402);
nand U1150 (N_1150,In_1708,In_1807);
xor U1151 (N_1151,In_944,In_1504);
nor U1152 (N_1152,In_2447,In_371);
nor U1153 (N_1153,In_1914,In_334);
and U1154 (N_1154,In_453,In_1828);
or U1155 (N_1155,In_1665,In_164);
nor U1156 (N_1156,In_2140,In_2191);
and U1157 (N_1157,In_2136,In_1231);
and U1158 (N_1158,In_1494,In_1561);
or U1159 (N_1159,In_416,In_1522);
xor U1160 (N_1160,In_423,In_1005);
or U1161 (N_1161,In_1276,In_407);
or U1162 (N_1162,In_642,In_1299);
and U1163 (N_1163,In_2330,In_1452);
nor U1164 (N_1164,In_459,In_1360);
and U1165 (N_1165,In_1055,In_367);
xor U1166 (N_1166,In_670,In_1034);
and U1167 (N_1167,In_776,In_1058);
or U1168 (N_1168,In_348,In_2494);
and U1169 (N_1169,In_1112,In_1531);
nor U1170 (N_1170,In_681,In_1090);
or U1171 (N_1171,In_696,In_716);
nand U1172 (N_1172,In_2322,In_943);
nor U1173 (N_1173,In_1882,In_2196);
nand U1174 (N_1174,In_1542,In_631);
nand U1175 (N_1175,In_494,In_2491);
and U1176 (N_1176,In_2133,In_1158);
nand U1177 (N_1177,In_1632,In_2042);
nand U1178 (N_1178,In_466,In_1783);
nor U1179 (N_1179,In_1250,In_2227);
nor U1180 (N_1180,In_1263,In_1635);
and U1181 (N_1181,In_1003,In_950);
nand U1182 (N_1182,In_601,In_80);
or U1183 (N_1183,In_2355,In_159);
nand U1184 (N_1184,In_649,In_2233);
or U1185 (N_1185,In_2086,In_439);
nor U1186 (N_1186,In_473,In_903);
and U1187 (N_1187,In_791,In_93);
nor U1188 (N_1188,In_509,In_2372);
nor U1189 (N_1189,In_2200,In_178);
nor U1190 (N_1190,In_2107,In_1770);
and U1191 (N_1191,In_725,In_596);
or U1192 (N_1192,In_876,In_1342);
and U1193 (N_1193,In_538,In_552);
and U1194 (N_1194,In_2433,In_2030);
nand U1195 (N_1195,In_1405,In_2082);
nand U1196 (N_1196,In_2201,In_2105);
or U1197 (N_1197,In_1430,In_1433);
xor U1198 (N_1198,In_2141,In_1279);
and U1199 (N_1199,In_1802,In_1025);
xnor U1200 (N_1200,In_1059,In_212);
nand U1201 (N_1201,In_1889,In_2331);
or U1202 (N_1202,In_2244,In_1638);
nand U1203 (N_1203,In_424,In_1620);
and U1204 (N_1204,In_723,In_993);
nor U1205 (N_1205,In_1023,In_568);
nand U1206 (N_1206,In_1474,In_1399);
and U1207 (N_1207,In_1031,In_2408);
or U1208 (N_1208,In_1763,In_504);
xor U1209 (N_1209,In_2407,In_2289);
and U1210 (N_1210,In_834,In_542);
nand U1211 (N_1211,In_2413,In_2143);
xnor U1212 (N_1212,In_343,In_805);
xnor U1213 (N_1213,In_421,In_70);
nor U1214 (N_1214,In_1593,In_206);
or U1215 (N_1215,In_2290,In_296);
xnor U1216 (N_1216,In_2008,In_772);
and U1217 (N_1217,In_2202,In_760);
or U1218 (N_1218,In_785,In_1734);
and U1219 (N_1219,In_1097,In_1223);
and U1220 (N_1220,In_375,In_726);
or U1221 (N_1221,In_1913,In_972);
nand U1222 (N_1222,In_1129,In_1759);
or U1223 (N_1223,In_2251,In_1052);
nand U1224 (N_1224,In_100,In_1970);
nand U1225 (N_1225,In_1157,In_2208);
xnor U1226 (N_1226,In_895,In_1164);
xor U1227 (N_1227,In_724,In_2044);
nor U1228 (N_1228,In_2039,In_2365);
and U1229 (N_1229,In_1413,In_1543);
xor U1230 (N_1230,In_1386,In_1124);
nor U1231 (N_1231,In_1716,In_518);
or U1232 (N_1232,In_1892,In_11);
nand U1233 (N_1233,In_636,In_2241);
and U1234 (N_1234,In_2149,In_2051);
nor U1235 (N_1235,In_2280,In_2439);
and U1236 (N_1236,In_1419,In_151);
nand U1237 (N_1237,In_982,In_604);
xnor U1238 (N_1238,In_909,In_41);
nor U1239 (N_1239,In_1187,In_2203);
xor U1240 (N_1240,In_105,In_1897);
nor U1241 (N_1241,In_500,In_2159);
nand U1242 (N_1242,In_200,In_592);
nand U1243 (N_1243,In_350,In_1849);
and U1244 (N_1244,In_1612,In_1888);
nand U1245 (N_1245,In_790,In_1239);
or U1246 (N_1246,In_40,In_265);
and U1247 (N_1247,In_2382,In_308);
xor U1248 (N_1248,In_503,In_2367);
or U1249 (N_1249,In_2118,In_2315);
or U1250 (N_1250,In_1261,In_2121);
nand U1251 (N_1251,In_2151,In_1031);
nand U1252 (N_1252,In_1274,In_1491);
and U1253 (N_1253,In_2264,In_2066);
and U1254 (N_1254,In_527,In_2109);
nor U1255 (N_1255,In_422,In_414);
or U1256 (N_1256,In_620,In_458);
xnor U1257 (N_1257,In_145,In_105);
xnor U1258 (N_1258,In_2354,In_1918);
nor U1259 (N_1259,In_964,In_1542);
or U1260 (N_1260,In_328,In_341);
xor U1261 (N_1261,In_157,In_1631);
nand U1262 (N_1262,In_1394,In_1972);
nor U1263 (N_1263,In_436,In_1265);
xor U1264 (N_1264,In_1872,In_1569);
and U1265 (N_1265,In_1584,In_2216);
xnor U1266 (N_1266,In_1454,In_1382);
xnor U1267 (N_1267,In_906,In_2056);
or U1268 (N_1268,In_1075,In_1585);
xor U1269 (N_1269,In_2217,In_586);
xor U1270 (N_1270,In_2083,In_1978);
or U1271 (N_1271,In_956,In_2389);
and U1272 (N_1272,In_322,In_384);
and U1273 (N_1273,In_1093,In_470);
nor U1274 (N_1274,In_158,In_2069);
nor U1275 (N_1275,In_1604,In_445);
and U1276 (N_1276,In_298,In_898);
nand U1277 (N_1277,In_1431,In_2404);
nor U1278 (N_1278,In_1159,In_687);
or U1279 (N_1279,In_1888,In_361);
and U1280 (N_1280,In_521,In_1687);
and U1281 (N_1281,In_1546,In_747);
and U1282 (N_1282,In_1140,In_207);
xor U1283 (N_1283,In_895,In_2057);
and U1284 (N_1284,In_391,In_1952);
and U1285 (N_1285,In_1811,In_218);
or U1286 (N_1286,In_2044,In_609);
and U1287 (N_1287,In_2481,In_1685);
nand U1288 (N_1288,In_1646,In_1351);
and U1289 (N_1289,In_973,In_2093);
and U1290 (N_1290,In_329,In_2405);
xor U1291 (N_1291,In_1135,In_951);
nor U1292 (N_1292,In_307,In_1432);
xor U1293 (N_1293,In_1738,In_650);
nor U1294 (N_1294,In_575,In_2495);
nand U1295 (N_1295,In_1903,In_369);
xnor U1296 (N_1296,In_1349,In_156);
or U1297 (N_1297,In_847,In_2250);
nand U1298 (N_1298,In_1704,In_473);
or U1299 (N_1299,In_1168,In_1638);
nor U1300 (N_1300,In_10,In_1421);
nor U1301 (N_1301,In_314,In_1486);
nand U1302 (N_1302,In_1416,In_2376);
nand U1303 (N_1303,In_527,In_1730);
and U1304 (N_1304,In_1933,In_196);
nand U1305 (N_1305,In_1583,In_1835);
nand U1306 (N_1306,In_2054,In_1121);
nand U1307 (N_1307,In_1567,In_2309);
and U1308 (N_1308,In_2074,In_902);
and U1309 (N_1309,In_300,In_1368);
and U1310 (N_1310,In_2176,In_1985);
nand U1311 (N_1311,In_340,In_1561);
nand U1312 (N_1312,In_1315,In_2174);
nand U1313 (N_1313,In_1735,In_450);
or U1314 (N_1314,In_1869,In_790);
or U1315 (N_1315,In_1606,In_449);
or U1316 (N_1316,In_195,In_1561);
xnor U1317 (N_1317,In_467,In_58);
or U1318 (N_1318,In_2395,In_383);
and U1319 (N_1319,In_2020,In_1593);
nand U1320 (N_1320,In_899,In_365);
and U1321 (N_1321,In_1887,In_1963);
nor U1322 (N_1322,In_1107,In_751);
or U1323 (N_1323,In_597,In_1261);
nand U1324 (N_1324,In_1451,In_1916);
nor U1325 (N_1325,In_54,In_826);
xor U1326 (N_1326,In_1211,In_2191);
xnor U1327 (N_1327,In_1095,In_1676);
or U1328 (N_1328,In_2294,In_103);
or U1329 (N_1329,In_610,In_422);
xnor U1330 (N_1330,In_1868,In_2125);
nand U1331 (N_1331,In_219,In_1698);
or U1332 (N_1332,In_734,In_2181);
xor U1333 (N_1333,In_263,In_323);
xor U1334 (N_1334,In_1879,In_1551);
nand U1335 (N_1335,In_963,In_1025);
and U1336 (N_1336,In_1077,In_652);
nor U1337 (N_1337,In_1951,In_2269);
nor U1338 (N_1338,In_968,In_1065);
xor U1339 (N_1339,In_746,In_181);
nand U1340 (N_1340,In_1473,In_866);
or U1341 (N_1341,In_1071,In_349);
nor U1342 (N_1342,In_970,In_154);
nand U1343 (N_1343,In_1017,In_522);
and U1344 (N_1344,In_1748,In_1160);
nor U1345 (N_1345,In_1161,In_640);
and U1346 (N_1346,In_1868,In_1937);
nand U1347 (N_1347,In_1329,In_591);
or U1348 (N_1348,In_40,In_2252);
or U1349 (N_1349,In_2235,In_2414);
or U1350 (N_1350,In_997,In_317);
or U1351 (N_1351,In_1389,In_808);
or U1352 (N_1352,In_923,In_102);
nor U1353 (N_1353,In_2163,In_2278);
xor U1354 (N_1354,In_2259,In_678);
or U1355 (N_1355,In_643,In_1845);
nor U1356 (N_1356,In_213,In_1067);
nand U1357 (N_1357,In_1497,In_590);
or U1358 (N_1358,In_2415,In_1535);
and U1359 (N_1359,In_750,In_760);
nand U1360 (N_1360,In_1269,In_2484);
and U1361 (N_1361,In_897,In_774);
and U1362 (N_1362,In_1135,In_636);
nor U1363 (N_1363,In_1105,In_1160);
and U1364 (N_1364,In_1850,In_602);
nand U1365 (N_1365,In_1590,In_1627);
xor U1366 (N_1366,In_1773,In_1176);
or U1367 (N_1367,In_1814,In_31);
xor U1368 (N_1368,In_1394,In_1082);
and U1369 (N_1369,In_1729,In_1625);
xor U1370 (N_1370,In_663,In_640);
nand U1371 (N_1371,In_2420,In_1589);
xnor U1372 (N_1372,In_91,In_1338);
and U1373 (N_1373,In_212,In_847);
nor U1374 (N_1374,In_2335,In_1749);
xor U1375 (N_1375,In_1519,In_734);
nor U1376 (N_1376,In_876,In_464);
or U1377 (N_1377,In_139,In_60);
and U1378 (N_1378,In_2366,In_749);
and U1379 (N_1379,In_649,In_464);
xnor U1380 (N_1380,In_2085,In_1);
nor U1381 (N_1381,In_1149,In_120);
or U1382 (N_1382,In_509,In_1643);
and U1383 (N_1383,In_707,In_1514);
nand U1384 (N_1384,In_187,In_1826);
nand U1385 (N_1385,In_343,In_420);
and U1386 (N_1386,In_1044,In_425);
nor U1387 (N_1387,In_1761,In_43);
and U1388 (N_1388,In_23,In_465);
xnor U1389 (N_1389,In_1717,In_1311);
or U1390 (N_1390,In_948,In_1240);
or U1391 (N_1391,In_788,In_692);
nor U1392 (N_1392,In_2485,In_587);
and U1393 (N_1393,In_2417,In_183);
and U1394 (N_1394,In_914,In_737);
and U1395 (N_1395,In_1122,In_923);
xor U1396 (N_1396,In_2218,In_228);
nor U1397 (N_1397,In_1364,In_1027);
and U1398 (N_1398,In_1929,In_1005);
nor U1399 (N_1399,In_1933,In_507);
and U1400 (N_1400,In_2108,In_1153);
xnor U1401 (N_1401,In_1746,In_71);
nand U1402 (N_1402,In_1536,In_1477);
and U1403 (N_1403,In_2314,In_212);
and U1404 (N_1404,In_142,In_1952);
nand U1405 (N_1405,In_1323,In_1507);
and U1406 (N_1406,In_2444,In_194);
nand U1407 (N_1407,In_1733,In_327);
or U1408 (N_1408,In_2276,In_2403);
or U1409 (N_1409,In_2107,In_2054);
xor U1410 (N_1410,In_577,In_578);
or U1411 (N_1411,In_1961,In_1059);
nand U1412 (N_1412,In_2302,In_814);
nor U1413 (N_1413,In_157,In_733);
xor U1414 (N_1414,In_2433,In_849);
or U1415 (N_1415,In_1858,In_1245);
nand U1416 (N_1416,In_1953,In_11);
nor U1417 (N_1417,In_508,In_1028);
nand U1418 (N_1418,In_1239,In_2070);
nor U1419 (N_1419,In_203,In_1699);
nand U1420 (N_1420,In_355,In_2438);
or U1421 (N_1421,In_789,In_730);
nor U1422 (N_1422,In_1997,In_1634);
or U1423 (N_1423,In_305,In_2158);
or U1424 (N_1424,In_463,In_905);
nand U1425 (N_1425,In_509,In_1771);
or U1426 (N_1426,In_2133,In_677);
nor U1427 (N_1427,In_2309,In_13);
nor U1428 (N_1428,In_905,In_1409);
nor U1429 (N_1429,In_890,In_2133);
xnor U1430 (N_1430,In_2341,In_1263);
and U1431 (N_1431,In_1881,In_280);
or U1432 (N_1432,In_798,In_463);
and U1433 (N_1433,In_2320,In_250);
nor U1434 (N_1434,In_444,In_1385);
nor U1435 (N_1435,In_935,In_1443);
and U1436 (N_1436,In_260,In_613);
xnor U1437 (N_1437,In_2252,In_1272);
xor U1438 (N_1438,In_1729,In_831);
and U1439 (N_1439,In_1509,In_2424);
and U1440 (N_1440,In_543,In_2153);
nand U1441 (N_1441,In_2,In_2149);
and U1442 (N_1442,In_205,In_1318);
nor U1443 (N_1443,In_1299,In_728);
and U1444 (N_1444,In_520,In_1762);
or U1445 (N_1445,In_1491,In_2190);
and U1446 (N_1446,In_1108,In_1002);
or U1447 (N_1447,In_756,In_1284);
and U1448 (N_1448,In_156,In_317);
or U1449 (N_1449,In_1321,In_2493);
nand U1450 (N_1450,In_1239,In_669);
nand U1451 (N_1451,In_2032,In_613);
nand U1452 (N_1452,In_1890,In_1264);
nor U1453 (N_1453,In_1344,In_298);
and U1454 (N_1454,In_2182,In_183);
nand U1455 (N_1455,In_1194,In_88);
nor U1456 (N_1456,In_183,In_891);
nor U1457 (N_1457,In_2024,In_918);
xor U1458 (N_1458,In_572,In_353);
or U1459 (N_1459,In_1476,In_664);
nor U1460 (N_1460,In_697,In_892);
nor U1461 (N_1461,In_180,In_764);
nand U1462 (N_1462,In_187,In_1650);
xnor U1463 (N_1463,In_1608,In_912);
nor U1464 (N_1464,In_1640,In_1982);
and U1465 (N_1465,In_612,In_588);
xor U1466 (N_1466,In_2492,In_1815);
nor U1467 (N_1467,In_964,In_1106);
and U1468 (N_1468,In_1063,In_41);
or U1469 (N_1469,In_2123,In_1795);
xor U1470 (N_1470,In_669,In_714);
nor U1471 (N_1471,In_613,In_2467);
nand U1472 (N_1472,In_509,In_331);
xnor U1473 (N_1473,In_2010,In_2038);
nor U1474 (N_1474,In_2394,In_1714);
nand U1475 (N_1475,In_1945,In_2245);
nor U1476 (N_1476,In_104,In_2233);
and U1477 (N_1477,In_1728,In_1199);
or U1478 (N_1478,In_757,In_1488);
or U1479 (N_1479,In_1469,In_1268);
and U1480 (N_1480,In_1516,In_2386);
and U1481 (N_1481,In_1947,In_431);
or U1482 (N_1482,In_2471,In_1538);
or U1483 (N_1483,In_1452,In_235);
and U1484 (N_1484,In_147,In_1388);
or U1485 (N_1485,In_304,In_590);
nor U1486 (N_1486,In_2245,In_1126);
and U1487 (N_1487,In_266,In_56);
xnor U1488 (N_1488,In_2218,In_738);
xor U1489 (N_1489,In_2165,In_1061);
nand U1490 (N_1490,In_1832,In_2317);
or U1491 (N_1491,In_1302,In_449);
xor U1492 (N_1492,In_1307,In_577);
and U1493 (N_1493,In_812,In_1484);
nand U1494 (N_1494,In_2403,In_1323);
or U1495 (N_1495,In_2309,In_1945);
and U1496 (N_1496,In_1820,In_1584);
nor U1497 (N_1497,In_2124,In_2430);
nand U1498 (N_1498,In_507,In_474);
nand U1499 (N_1499,In_1761,In_197);
nand U1500 (N_1500,In_1572,In_2219);
and U1501 (N_1501,In_2264,In_1690);
or U1502 (N_1502,In_2363,In_930);
nand U1503 (N_1503,In_1799,In_411);
or U1504 (N_1504,In_1764,In_395);
and U1505 (N_1505,In_2010,In_600);
xor U1506 (N_1506,In_1323,In_399);
xnor U1507 (N_1507,In_1992,In_1309);
nand U1508 (N_1508,In_1877,In_718);
and U1509 (N_1509,In_698,In_658);
and U1510 (N_1510,In_1891,In_724);
nor U1511 (N_1511,In_144,In_357);
xnor U1512 (N_1512,In_940,In_1530);
nor U1513 (N_1513,In_211,In_1593);
xnor U1514 (N_1514,In_1862,In_286);
nand U1515 (N_1515,In_2017,In_892);
nand U1516 (N_1516,In_2261,In_532);
and U1517 (N_1517,In_971,In_1055);
xor U1518 (N_1518,In_621,In_2233);
and U1519 (N_1519,In_2109,In_259);
and U1520 (N_1520,In_1902,In_894);
xor U1521 (N_1521,In_2043,In_1879);
nand U1522 (N_1522,In_456,In_435);
xnor U1523 (N_1523,In_359,In_2030);
and U1524 (N_1524,In_292,In_2081);
nor U1525 (N_1525,In_728,In_1087);
nor U1526 (N_1526,In_1834,In_731);
xnor U1527 (N_1527,In_1527,In_967);
nand U1528 (N_1528,In_1888,In_1902);
xnor U1529 (N_1529,In_842,In_841);
nand U1530 (N_1530,In_411,In_762);
or U1531 (N_1531,In_1165,In_2268);
nand U1532 (N_1532,In_663,In_2094);
or U1533 (N_1533,In_1362,In_244);
nand U1534 (N_1534,In_1252,In_233);
or U1535 (N_1535,In_2454,In_2163);
nor U1536 (N_1536,In_1186,In_435);
nand U1537 (N_1537,In_1948,In_797);
or U1538 (N_1538,In_1641,In_1726);
or U1539 (N_1539,In_1145,In_2459);
and U1540 (N_1540,In_991,In_1835);
nor U1541 (N_1541,In_2460,In_720);
nand U1542 (N_1542,In_2239,In_1860);
or U1543 (N_1543,In_1615,In_2497);
and U1544 (N_1544,In_1346,In_1709);
nor U1545 (N_1545,In_373,In_1839);
or U1546 (N_1546,In_292,In_1407);
xnor U1547 (N_1547,In_1693,In_996);
and U1548 (N_1548,In_2183,In_1683);
nor U1549 (N_1549,In_424,In_682);
nor U1550 (N_1550,In_1218,In_311);
nand U1551 (N_1551,In_665,In_1277);
or U1552 (N_1552,In_1654,In_467);
nor U1553 (N_1553,In_2190,In_691);
nor U1554 (N_1554,In_1947,In_1217);
xnor U1555 (N_1555,In_2356,In_2234);
nor U1556 (N_1556,In_2000,In_918);
and U1557 (N_1557,In_248,In_379);
and U1558 (N_1558,In_1782,In_148);
nand U1559 (N_1559,In_502,In_2120);
and U1560 (N_1560,In_2100,In_44);
and U1561 (N_1561,In_1294,In_1718);
or U1562 (N_1562,In_1626,In_880);
xnor U1563 (N_1563,In_1821,In_744);
nand U1564 (N_1564,In_2421,In_2373);
nor U1565 (N_1565,In_1522,In_815);
nand U1566 (N_1566,In_917,In_2263);
or U1567 (N_1567,In_2314,In_1371);
nor U1568 (N_1568,In_1329,In_10);
nor U1569 (N_1569,In_1026,In_893);
or U1570 (N_1570,In_608,In_1739);
and U1571 (N_1571,In_2293,In_1280);
nand U1572 (N_1572,In_2006,In_593);
nand U1573 (N_1573,In_459,In_1567);
xor U1574 (N_1574,In_1625,In_934);
nand U1575 (N_1575,In_2148,In_2431);
and U1576 (N_1576,In_1048,In_1536);
nand U1577 (N_1577,In_2433,In_2424);
or U1578 (N_1578,In_2300,In_778);
and U1579 (N_1579,In_1947,In_603);
nor U1580 (N_1580,In_583,In_1004);
nor U1581 (N_1581,In_785,In_827);
nor U1582 (N_1582,In_1981,In_2161);
and U1583 (N_1583,In_1919,In_1123);
and U1584 (N_1584,In_1781,In_2106);
nand U1585 (N_1585,In_1569,In_467);
xor U1586 (N_1586,In_2053,In_1393);
nor U1587 (N_1587,In_1713,In_2235);
and U1588 (N_1588,In_1975,In_1469);
and U1589 (N_1589,In_1563,In_430);
nor U1590 (N_1590,In_59,In_1420);
or U1591 (N_1591,In_463,In_2243);
or U1592 (N_1592,In_2401,In_886);
xor U1593 (N_1593,In_152,In_336);
nor U1594 (N_1594,In_365,In_887);
and U1595 (N_1595,In_469,In_639);
nor U1596 (N_1596,In_1132,In_1925);
nand U1597 (N_1597,In_748,In_1297);
and U1598 (N_1598,In_953,In_1523);
and U1599 (N_1599,In_942,In_756);
nand U1600 (N_1600,In_715,In_1585);
nor U1601 (N_1601,In_763,In_1);
xnor U1602 (N_1602,In_637,In_1847);
and U1603 (N_1603,In_791,In_502);
or U1604 (N_1604,In_1611,In_1093);
and U1605 (N_1605,In_1837,In_1482);
or U1606 (N_1606,In_2311,In_697);
or U1607 (N_1607,In_987,In_1009);
nand U1608 (N_1608,In_1142,In_2308);
nor U1609 (N_1609,In_1663,In_355);
nand U1610 (N_1610,In_2072,In_1248);
or U1611 (N_1611,In_2457,In_84);
or U1612 (N_1612,In_995,In_2080);
and U1613 (N_1613,In_838,In_1057);
and U1614 (N_1614,In_174,In_2072);
nor U1615 (N_1615,In_1378,In_95);
or U1616 (N_1616,In_1333,In_2283);
nand U1617 (N_1617,In_1554,In_1787);
and U1618 (N_1618,In_1451,In_1791);
nor U1619 (N_1619,In_2020,In_705);
and U1620 (N_1620,In_1365,In_679);
and U1621 (N_1621,In_950,In_389);
nor U1622 (N_1622,In_354,In_1785);
xor U1623 (N_1623,In_152,In_1517);
nand U1624 (N_1624,In_1743,In_1634);
and U1625 (N_1625,In_1944,In_2148);
or U1626 (N_1626,In_2043,In_1795);
or U1627 (N_1627,In_91,In_836);
or U1628 (N_1628,In_1644,In_158);
or U1629 (N_1629,In_1128,In_1604);
nor U1630 (N_1630,In_1019,In_2242);
and U1631 (N_1631,In_351,In_1105);
or U1632 (N_1632,In_1981,In_326);
nand U1633 (N_1633,In_1542,In_1846);
or U1634 (N_1634,In_1634,In_531);
nor U1635 (N_1635,In_526,In_1896);
nand U1636 (N_1636,In_100,In_1396);
or U1637 (N_1637,In_822,In_1682);
or U1638 (N_1638,In_1685,In_1199);
nor U1639 (N_1639,In_1825,In_1795);
and U1640 (N_1640,In_743,In_419);
xor U1641 (N_1641,In_942,In_1269);
xor U1642 (N_1642,In_1649,In_645);
nand U1643 (N_1643,In_2296,In_2092);
nor U1644 (N_1644,In_835,In_2054);
xor U1645 (N_1645,In_861,In_434);
or U1646 (N_1646,In_796,In_1311);
and U1647 (N_1647,In_1952,In_406);
and U1648 (N_1648,In_880,In_2174);
and U1649 (N_1649,In_696,In_822);
xnor U1650 (N_1650,In_1559,In_1447);
nor U1651 (N_1651,In_2337,In_1706);
and U1652 (N_1652,In_399,In_618);
xnor U1653 (N_1653,In_1096,In_278);
and U1654 (N_1654,In_2154,In_1100);
xnor U1655 (N_1655,In_1036,In_596);
or U1656 (N_1656,In_2368,In_998);
or U1657 (N_1657,In_869,In_1965);
xnor U1658 (N_1658,In_389,In_816);
nor U1659 (N_1659,In_2326,In_514);
and U1660 (N_1660,In_1012,In_1142);
nand U1661 (N_1661,In_2044,In_1731);
nand U1662 (N_1662,In_2365,In_512);
nand U1663 (N_1663,In_1523,In_1310);
xor U1664 (N_1664,In_2033,In_2104);
nor U1665 (N_1665,In_677,In_1668);
nor U1666 (N_1666,In_1045,In_1906);
nand U1667 (N_1667,In_666,In_1781);
or U1668 (N_1668,In_1549,In_1688);
nor U1669 (N_1669,In_1671,In_718);
xnor U1670 (N_1670,In_562,In_117);
nand U1671 (N_1671,In_1332,In_2199);
and U1672 (N_1672,In_886,In_1460);
nor U1673 (N_1673,In_2298,In_405);
nor U1674 (N_1674,In_1723,In_702);
nand U1675 (N_1675,In_2298,In_2234);
nand U1676 (N_1676,In_2115,In_2394);
nand U1677 (N_1677,In_432,In_1564);
and U1678 (N_1678,In_1296,In_191);
nand U1679 (N_1679,In_742,In_1186);
xor U1680 (N_1680,In_1804,In_2262);
and U1681 (N_1681,In_722,In_2437);
xnor U1682 (N_1682,In_2129,In_2263);
nor U1683 (N_1683,In_1354,In_1524);
nand U1684 (N_1684,In_2243,In_439);
xnor U1685 (N_1685,In_853,In_2254);
or U1686 (N_1686,In_337,In_608);
xnor U1687 (N_1687,In_1062,In_335);
nor U1688 (N_1688,In_1885,In_1521);
and U1689 (N_1689,In_236,In_343);
xor U1690 (N_1690,In_672,In_1654);
nand U1691 (N_1691,In_1026,In_1185);
nor U1692 (N_1692,In_2201,In_1277);
nor U1693 (N_1693,In_1296,In_1456);
and U1694 (N_1694,In_1957,In_2040);
or U1695 (N_1695,In_1739,In_371);
xor U1696 (N_1696,In_1602,In_1127);
nand U1697 (N_1697,In_852,In_1532);
and U1698 (N_1698,In_1172,In_71);
or U1699 (N_1699,In_395,In_278);
xnor U1700 (N_1700,In_58,In_1768);
nor U1701 (N_1701,In_2405,In_129);
and U1702 (N_1702,In_2014,In_2021);
xnor U1703 (N_1703,In_1060,In_1112);
or U1704 (N_1704,In_942,In_2080);
and U1705 (N_1705,In_1517,In_2496);
nand U1706 (N_1706,In_2311,In_1634);
nand U1707 (N_1707,In_1993,In_288);
nand U1708 (N_1708,In_285,In_770);
xnor U1709 (N_1709,In_597,In_380);
xnor U1710 (N_1710,In_1877,In_1051);
xor U1711 (N_1711,In_636,In_2361);
nor U1712 (N_1712,In_2312,In_1636);
xnor U1713 (N_1713,In_707,In_992);
and U1714 (N_1714,In_1108,In_78);
or U1715 (N_1715,In_2331,In_715);
nand U1716 (N_1716,In_1165,In_2312);
nand U1717 (N_1717,In_2468,In_2430);
xnor U1718 (N_1718,In_233,In_739);
and U1719 (N_1719,In_921,In_171);
xor U1720 (N_1720,In_1637,In_2303);
or U1721 (N_1721,In_2119,In_943);
or U1722 (N_1722,In_1371,In_2452);
or U1723 (N_1723,In_1681,In_2399);
nand U1724 (N_1724,In_85,In_166);
and U1725 (N_1725,In_381,In_2083);
nand U1726 (N_1726,In_2434,In_68);
nand U1727 (N_1727,In_401,In_1019);
or U1728 (N_1728,In_278,In_693);
nand U1729 (N_1729,In_345,In_813);
nand U1730 (N_1730,In_503,In_637);
nor U1731 (N_1731,In_640,In_466);
or U1732 (N_1732,In_791,In_780);
and U1733 (N_1733,In_535,In_2226);
nor U1734 (N_1734,In_1339,In_1219);
and U1735 (N_1735,In_862,In_767);
or U1736 (N_1736,In_381,In_294);
nand U1737 (N_1737,In_2150,In_1781);
nor U1738 (N_1738,In_2162,In_316);
and U1739 (N_1739,In_2498,In_108);
xor U1740 (N_1740,In_1668,In_2468);
or U1741 (N_1741,In_774,In_1226);
xor U1742 (N_1742,In_1994,In_1694);
nor U1743 (N_1743,In_1096,In_2443);
nor U1744 (N_1744,In_283,In_1242);
or U1745 (N_1745,In_550,In_2442);
xor U1746 (N_1746,In_534,In_623);
xnor U1747 (N_1747,In_372,In_493);
and U1748 (N_1748,In_997,In_916);
nor U1749 (N_1749,In_1553,In_1311);
or U1750 (N_1750,In_5,In_2352);
and U1751 (N_1751,In_732,In_1607);
nor U1752 (N_1752,In_1965,In_730);
xor U1753 (N_1753,In_58,In_1337);
nand U1754 (N_1754,In_1099,In_1347);
and U1755 (N_1755,In_1315,In_1641);
nor U1756 (N_1756,In_2375,In_681);
nor U1757 (N_1757,In_1776,In_1301);
and U1758 (N_1758,In_82,In_1669);
or U1759 (N_1759,In_2422,In_913);
xor U1760 (N_1760,In_884,In_1910);
or U1761 (N_1761,In_306,In_2382);
and U1762 (N_1762,In_189,In_100);
nand U1763 (N_1763,In_643,In_1327);
nor U1764 (N_1764,In_613,In_1586);
nor U1765 (N_1765,In_2212,In_309);
xnor U1766 (N_1766,In_288,In_2319);
and U1767 (N_1767,In_867,In_1704);
xor U1768 (N_1768,In_1675,In_889);
nand U1769 (N_1769,In_1131,In_1609);
and U1770 (N_1770,In_638,In_58);
nor U1771 (N_1771,In_889,In_888);
and U1772 (N_1772,In_2117,In_350);
nor U1773 (N_1773,In_267,In_1409);
and U1774 (N_1774,In_2165,In_169);
nand U1775 (N_1775,In_561,In_640);
nand U1776 (N_1776,In_2390,In_1696);
xnor U1777 (N_1777,In_1013,In_844);
or U1778 (N_1778,In_1540,In_2173);
nand U1779 (N_1779,In_757,In_1125);
and U1780 (N_1780,In_228,In_2320);
nor U1781 (N_1781,In_1553,In_1127);
or U1782 (N_1782,In_1019,In_2371);
nand U1783 (N_1783,In_1866,In_1799);
xor U1784 (N_1784,In_263,In_1959);
nand U1785 (N_1785,In_789,In_195);
nor U1786 (N_1786,In_347,In_1521);
nand U1787 (N_1787,In_850,In_1199);
or U1788 (N_1788,In_438,In_665);
nor U1789 (N_1789,In_2187,In_669);
nand U1790 (N_1790,In_562,In_862);
nand U1791 (N_1791,In_1399,In_1200);
nor U1792 (N_1792,In_852,In_1230);
nand U1793 (N_1793,In_1534,In_2493);
or U1794 (N_1794,In_1086,In_601);
xnor U1795 (N_1795,In_405,In_1897);
and U1796 (N_1796,In_1470,In_530);
nand U1797 (N_1797,In_1457,In_1322);
and U1798 (N_1798,In_428,In_1202);
or U1799 (N_1799,In_1915,In_1187);
xor U1800 (N_1800,In_2167,In_2217);
xor U1801 (N_1801,In_1043,In_1206);
nand U1802 (N_1802,In_254,In_2158);
nand U1803 (N_1803,In_1554,In_2077);
nor U1804 (N_1804,In_227,In_2395);
and U1805 (N_1805,In_1767,In_1847);
nand U1806 (N_1806,In_1620,In_1316);
nand U1807 (N_1807,In_1403,In_2255);
nand U1808 (N_1808,In_900,In_225);
xor U1809 (N_1809,In_2351,In_48);
or U1810 (N_1810,In_2411,In_2053);
nor U1811 (N_1811,In_1137,In_498);
xor U1812 (N_1812,In_1091,In_1004);
nor U1813 (N_1813,In_1785,In_1231);
and U1814 (N_1814,In_1182,In_176);
and U1815 (N_1815,In_75,In_1598);
nor U1816 (N_1816,In_1297,In_1933);
nor U1817 (N_1817,In_1872,In_1847);
xnor U1818 (N_1818,In_927,In_87);
or U1819 (N_1819,In_1355,In_1972);
or U1820 (N_1820,In_2469,In_660);
and U1821 (N_1821,In_1123,In_945);
nor U1822 (N_1822,In_37,In_433);
nand U1823 (N_1823,In_1944,In_800);
and U1824 (N_1824,In_102,In_2393);
nand U1825 (N_1825,In_373,In_1164);
or U1826 (N_1826,In_1398,In_522);
nor U1827 (N_1827,In_1940,In_972);
xnor U1828 (N_1828,In_2449,In_1299);
xor U1829 (N_1829,In_1010,In_1547);
or U1830 (N_1830,In_100,In_2336);
nand U1831 (N_1831,In_1640,In_12);
and U1832 (N_1832,In_2259,In_1434);
and U1833 (N_1833,In_2017,In_52);
and U1834 (N_1834,In_2312,In_2214);
nand U1835 (N_1835,In_1601,In_42);
nor U1836 (N_1836,In_2041,In_640);
or U1837 (N_1837,In_2121,In_1172);
nor U1838 (N_1838,In_2093,In_1280);
or U1839 (N_1839,In_270,In_817);
and U1840 (N_1840,In_598,In_1171);
or U1841 (N_1841,In_151,In_447);
or U1842 (N_1842,In_879,In_501);
and U1843 (N_1843,In_327,In_1097);
or U1844 (N_1844,In_2141,In_1085);
or U1845 (N_1845,In_2242,In_401);
or U1846 (N_1846,In_1398,In_2385);
or U1847 (N_1847,In_113,In_2100);
nand U1848 (N_1848,In_2126,In_63);
or U1849 (N_1849,In_1383,In_1725);
nand U1850 (N_1850,In_1315,In_168);
nand U1851 (N_1851,In_409,In_1315);
and U1852 (N_1852,In_2063,In_1448);
and U1853 (N_1853,In_434,In_1125);
nand U1854 (N_1854,In_1547,In_638);
nand U1855 (N_1855,In_282,In_704);
or U1856 (N_1856,In_1530,In_1572);
and U1857 (N_1857,In_2223,In_2487);
nor U1858 (N_1858,In_170,In_552);
xnor U1859 (N_1859,In_1895,In_902);
nand U1860 (N_1860,In_1858,In_2369);
nor U1861 (N_1861,In_1195,In_67);
nor U1862 (N_1862,In_53,In_2315);
xor U1863 (N_1863,In_2427,In_1286);
nor U1864 (N_1864,In_589,In_1302);
xnor U1865 (N_1865,In_1988,In_1991);
and U1866 (N_1866,In_1762,In_811);
nor U1867 (N_1867,In_1543,In_192);
nor U1868 (N_1868,In_1458,In_1955);
or U1869 (N_1869,In_1614,In_660);
nor U1870 (N_1870,In_529,In_1170);
nor U1871 (N_1871,In_1247,In_2293);
or U1872 (N_1872,In_942,In_702);
nor U1873 (N_1873,In_2450,In_540);
nor U1874 (N_1874,In_2439,In_1626);
and U1875 (N_1875,In_393,In_439);
nor U1876 (N_1876,In_243,In_1318);
nand U1877 (N_1877,In_150,In_1443);
nand U1878 (N_1878,In_911,In_2048);
nor U1879 (N_1879,In_564,In_1754);
nand U1880 (N_1880,In_956,In_1981);
or U1881 (N_1881,In_1092,In_1611);
nand U1882 (N_1882,In_1971,In_196);
nor U1883 (N_1883,In_1386,In_1946);
xnor U1884 (N_1884,In_795,In_138);
or U1885 (N_1885,In_1879,In_1719);
xor U1886 (N_1886,In_836,In_2051);
nand U1887 (N_1887,In_1875,In_1155);
nor U1888 (N_1888,In_2478,In_1907);
and U1889 (N_1889,In_1524,In_497);
xor U1890 (N_1890,In_470,In_858);
nor U1891 (N_1891,In_2230,In_1708);
xnor U1892 (N_1892,In_1986,In_608);
and U1893 (N_1893,In_695,In_1237);
xor U1894 (N_1894,In_122,In_1043);
or U1895 (N_1895,In_2171,In_2021);
nand U1896 (N_1896,In_263,In_1640);
or U1897 (N_1897,In_212,In_1219);
nor U1898 (N_1898,In_1058,In_1100);
nand U1899 (N_1899,In_1234,In_1105);
nand U1900 (N_1900,In_2349,In_17);
nor U1901 (N_1901,In_174,In_107);
or U1902 (N_1902,In_1387,In_2408);
xnor U1903 (N_1903,In_37,In_1823);
and U1904 (N_1904,In_2469,In_2066);
xor U1905 (N_1905,In_1277,In_137);
xnor U1906 (N_1906,In_2354,In_1978);
nand U1907 (N_1907,In_2326,In_2109);
and U1908 (N_1908,In_2300,In_1409);
xnor U1909 (N_1909,In_1640,In_2305);
and U1910 (N_1910,In_433,In_1263);
nand U1911 (N_1911,In_1822,In_1776);
and U1912 (N_1912,In_1575,In_2119);
nor U1913 (N_1913,In_1709,In_497);
or U1914 (N_1914,In_1565,In_105);
nor U1915 (N_1915,In_2416,In_1370);
nand U1916 (N_1916,In_2398,In_622);
and U1917 (N_1917,In_1388,In_1998);
and U1918 (N_1918,In_1607,In_1667);
or U1919 (N_1919,In_60,In_804);
nor U1920 (N_1920,In_1965,In_868);
or U1921 (N_1921,In_2327,In_1116);
nor U1922 (N_1922,In_1977,In_2273);
xor U1923 (N_1923,In_2052,In_2124);
or U1924 (N_1924,In_520,In_994);
and U1925 (N_1925,In_1736,In_2400);
nand U1926 (N_1926,In_500,In_1342);
xor U1927 (N_1927,In_35,In_282);
xor U1928 (N_1928,In_2258,In_984);
nand U1929 (N_1929,In_390,In_2307);
or U1930 (N_1930,In_799,In_147);
and U1931 (N_1931,In_1306,In_722);
and U1932 (N_1932,In_924,In_1167);
nor U1933 (N_1933,In_628,In_1087);
xor U1934 (N_1934,In_1170,In_496);
nand U1935 (N_1935,In_1782,In_1662);
nand U1936 (N_1936,In_1743,In_2438);
xnor U1937 (N_1937,In_2258,In_529);
nand U1938 (N_1938,In_224,In_2117);
or U1939 (N_1939,In_1639,In_2441);
nor U1940 (N_1940,In_2062,In_493);
xor U1941 (N_1941,In_2145,In_629);
or U1942 (N_1942,In_1261,In_2048);
nand U1943 (N_1943,In_448,In_219);
xnor U1944 (N_1944,In_872,In_2030);
nand U1945 (N_1945,In_615,In_1708);
nand U1946 (N_1946,In_302,In_1268);
nor U1947 (N_1947,In_2496,In_1316);
nor U1948 (N_1948,In_1332,In_759);
or U1949 (N_1949,In_1948,In_2189);
or U1950 (N_1950,In_632,In_1383);
and U1951 (N_1951,In_1043,In_1956);
nor U1952 (N_1952,In_1338,In_614);
nand U1953 (N_1953,In_307,In_1614);
xnor U1954 (N_1954,In_1161,In_711);
and U1955 (N_1955,In_121,In_538);
nand U1956 (N_1956,In_1642,In_1763);
and U1957 (N_1957,In_596,In_72);
nand U1958 (N_1958,In_1640,In_794);
and U1959 (N_1959,In_752,In_3);
or U1960 (N_1960,In_459,In_36);
and U1961 (N_1961,In_590,In_231);
or U1962 (N_1962,In_184,In_533);
and U1963 (N_1963,In_1718,In_2162);
nand U1964 (N_1964,In_1014,In_525);
or U1965 (N_1965,In_1398,In_1109);
and U1966 (N_1966,In_2197,In_858);
and U1967 (N_1967,In_854,In_123);
or U1968 (N_1968,In_1984,In_191);
nor U1969 (N_1969,In_236,In_1019);
xor U1970 (N_1970,In_6,In_1597);
and U1971 (N_1971,In_1405,In_753);
nand U1972 (N_1972,In_652,In_1790);
nor U1973 (N_1973,In_1949,In_2278);
or U1974 (N_1974,In_1430,In_1255);
xor U1975 (N_1975,In_1707,In_1829);
xnor U1976 (N_1976,In_1371,In_488);
nand U1977 (N_1977,In_1636,In_2220);
xor U1978 (N_1978,In_515,In_1269);
nor U1979 (N_1979,In_701,In_657);
xnor U1980 (N_1980,In_46,In_555);
nand U1981 (N_1981,In_2259,In_1498);
or U1982 (N_1982,In_2083,In_995);
xnor U1983 (N_1983,In_1609,In_73);
nand U1984 (N_1984,In_2191,In_1735);
xor U1985 (N_1985,In_2337,In_1070);
nand U1986 (N_1986,In_1374,In_1007);
or U1987 (N_1987,In_1876,In_1326);
nand U1988 (N_1988,In_1320,In_1376);
xor U1989 (N_1989,In_271,In_1397);
xor U1990 (N_1990,In_1401,In_1598);
or U1991 (N_1991,In_359,In_745);
or U1992 (N_1992,In_1020,In_1437);
or U1993 (N_1993,In_134,In_1349);
or U1994 (N_1994,In_1864,In_1279);
xnor U1995 (N_1995,In_614,In_1300);
and U1996 (N_1996,In_289,In_1912);
xor U1997 (N_1997,In_1216,In_1297);
xor U1998 (N_1998,In_768,In_2203);
nor U1999 (N_1999,In_43,In_1693);
xnor U2000 (N_2000,In_1219,In_1451);
or U2001 (N_2001,In_2445,In_1379);
and U2002 (N_2002,In_1,In_368);
nand U2003 (N_2003,In_2466,In_2451);
xor U2004 (N_2004,In_1350,In_232);
nand U2005 (N_2005,In_235,In_1459);
and U2006 (N_2006,In_1265,In_2393);
nor U2007 (N_2007,In_2228,In_581);
or U2008 (N_2008,In_44,In_1466);
nand U2009 (N_2009,In_2074,In_1986);
or U2010 (N_2010,In_760,In_1125);
and U2011 (N_2011,In_1314,In_1087);
or U2012 (N_2012,In_844,In_296);
or U2013 (N_2013,In_1664,In_1883);
or U2014 (N_2014,In_2282,In_710);
nand U2015 (N_2015,In_1198,In_257);
nand U2016 (N_2016,In_379,In_1586);
xnor U2017 (N_2017,In_188,In_317);
nor U2018 (N_2018,In_750,In_1227);
nand U2019 (N_2019,In_918,In_370);
nor U2020 (N_2020,In_1628,In_1691);
or U2021 (N_2021,In_1659,In_727);
nor U2022 (N_2022,In_1653,In_1832);
nor U2023 (N_2023,In_1774,In_2166);
nor U2024 (N_2024,In_1812,In_1953);
nor U2025 (N_2025,In_2058,In_1143);
xor U2026 (N_2026,In_1466,In_1282);
nand U2027 (N_2027,In_852,In_284);
nor U2028 (N_2028,In_2153,In_195);
and U2029 (N_2029,In_1797,In_351);
and U2030 (N_2030,In_223,In_1017);
nand U2031 (N_2031,In_129,In_2374);
nand U2032 (N_2032,In_2061,In_2309);
or U2033 (N_2033,In_1931,In_456);
and U2034 (N_2034,In_431,In_1425);
nand U2035 (N_2035,In_501,In_487);
nand U2036 (N_2036,In_211,In_584);
nor U2037 (N_2037,In_298,In_1987);
or U2038 (N_2038,In_1121,In_260);
or U2039 (N_2039,In_1702,In_2464);
xor U2040 (N_2040,In_2041,In_852);
nand U2041 (N_2041,In_1794,In_649);
or U2042 (N_2042,In_2296,In_1131);
xor U2043 (N_2043,In_265,In_2095);
nand U2044 (N_2044,In_200,In_2327);
nor U2045 (N_2045,In_171,In_783);
nor U2046 (N_2046,In_371,In_484);
or U2047 (N_2047,In_242,In_2158);
or U2048 (N_2048,In_1489,In_710);
nor U2049 (N_2049,In_1857,In_243);
and U2050 (N_2050,In_11,In_402);
and U2051 (N_2051,In_1135,In_210);
nand U2052 (N_2052,In_231,In_297);
and U2053 (N_2053,In_2339,In_266);
xor U2054 (N_2054,In_1000,In_934);
or U2055 (N_2055,In_1508,In_450);
or U2056 (N_2056,In_2264,In_2410);
xor U2057 (N_2057,In_1590,In_2438);
or U2058 (N_2058,In_1731,In_821);
nand U2059 (N_2059,In_1245,In_1406);
and U2060 (N_2060,In_685,In_1235);
xor U2061 (N_2061,In_730,In_2005);
and U2062 (N_2062,In_344,In_1095);
nand U2063 (N_2063,In_948,In_224);
and U2064 (N_2064,In_1046,In_108);
or U2065 (N_2065,In_249,In_721);
or U2066 (N_2066,In_381,In_431);
and U2067 (N_2067,In_1256,In_1161);
or U2068 (N_2068,In_633,In_889);
nand U2069 (N_2069,In_1612,In_417);
and U2070 (N_2070,In_1128,In_330);
and U2071 (N_2071,In_2091,In_2361);
xnor U2072 (N_2072,In_286,In_1607);
nand U2073 (N_2073,In_1523,In_1371);
and U2074 (N_2074,In_409,In_659);
or U2075 (N_2075,In_1151,In_2044);
or U2076 (N_2076,In_1745,In_195);
xor U2077 (N_2077,In_688,In_1347);
nor U2078 (N_2078,In_221,In_2245);
or U2079 (N_2079,In_41,In_417);
xnor U2080 (N_2080,In_908,In_1172);
nor U2081 (N_2081,In_1787,In_278);
nor U2082 (N_2082,In_1658,In_1702);
nand U2083 (N_2083,In_1662,In_1154);
nor U2084 (N_2084,In_548,In_1333);
or U2085 (N_2085,In_45,In_1936);
xnor U2086 (N_2086,In_2017,In_1045);
and U2087 (N_2087,In_575,In_46);
nor U2088 (N_2088,In_1447,In_2316);
or U2089 (N_2089,In_1533,In_437);
or U2090 (N_2090,In_620,In_89);
and U2091 (N_2091,In_2471,In_294);
or U2092 (N_2092,In_1907,In_221);
and U2093 (N_2093,In_337,In_1450);
or U2094 (N_2094,In_2383,In_1181);
and U2095 (N_2095,In_2238,In_1397);
and U2096 (N_2096,In_995,In_304);
nor U2097 (N_2097,In_1020,In_331);
or U2098 (N_2098,In_649,In_2151);
nand U2099 (N_2099,In_2097,In_12);
nand U2100 (N_2100,In_801,In_2184);
nor U2101 (N_2101,In_133,In_2331);
nor U2102 (N_2102,In_1359,In_516);
nor U2103 (N_2103,In_1140,In_890);
and U2104 (N_2104,In_1112,In_942);
or U2105 (N_2105,In_2223,In_753);
nand U2106 (N_2106,In_2155,In_264);
xnor U2107 (N_2107,In_345,In_859);
or U2108 (N_2108,In_1849,In_1630);
nand U2109 (N_2109,In_2268,In_401);
nand U2110 (N_2110,In_488,In_81);
or U2111 (N_2111,In_2235,In_218);
or U2112 (N_2112,In_50,In_155);
xor U2113 (N_2113,In_555,In_1679);
or U2114 (N_2114,In_1121,In_2418);
nor U2115 (N_2115,In_2206,In_2453);
nor U2116 (N_2116,In_1527,In_1019);
or U2117 (N_2117,In_19,In_1842);
and U2118 (N_2118,In_1026,In_643);
or U2119 (N_2119,In_670,In_1991);
and U2120 (N_2120,In_1383,In_98);
nor U2121 (N_2121,In_429,In_2120);
nand U2122 (N_2122,In_1706,In_2380);
nor U2123 (N_2123,In_888,In_1070);
or U2124 (N_2124,In_680,In_1878);
or U2125 (N_2125,In_411,In_32);
nor U2126 (N_2126,In_1617,In_2143);
nor U2127 (N_2127,In_909,In_508);
or U2128 (N_2128,In_1027,In_2165);
xnor U2129 (N_2129,In_1385,In_282);
and U2130 (N_2130,In_1133,In_121);
and U2131 (N_2131,In_960,In_1027);
xnor U2132 (N_2132,In_1876,In_2450);
nand U2133 (N_2133,In_1667,In_1232);
nor U2134 (N_2134,In_821,In_2419);
or U2135 (N_2135,In_750,In_1835);
nor U2136 (N_2136,In_1992,In_1438);
nor U2137 (N_2137,In_1205,In_2226);
or U2138 (N_2138,In_2106,In_2079);
xnor U2139 (N_2139,In_912,In_970);
and U2140 (N_2140,In_2085,In_1921);
or U2141 (N_2141,In_1981,In_869);
or U2142 (N_2142,In_357,In_1672);
nor U2143 (N_2143,In_388,In_647);
nand U2144 (N_2144,In_298,In_1990);
xnor U2145 (N_2145,In_2429,In_1948);
xor U2146 (N_2146,In_1483,In_1852);
and U2147 (N_2147,In_487,In_373);
or U2148 (N_2148,In_1386,In_2152);
or U2149 (N_2149,In_2366,In_1368);
nor U2150 (N_2150,In_1596,In_2146);
or U2151 (N_2151,In_1682,In_2394);
xnor U2152 (N_2152,In_899,In_2372);
nand U2153 (N_2153,In_2438,In_460);
and U2154 (N_2154,In_244,In_2235);
nor U2155 (N_2155,In_1569,In_207);
and U2156 (N_2156,In_2034,In_230);
xnor U2157 (N_2157,In_1569,In_889);
and U2158 (N_2158,In_954,In_572);
xor U2159 (N_2159,In_2284,In_420);
nor U2160 (N_2160,In_1539,In_176);
and U2161 (N_2161,In_146,In_401);
and U2162 (N_2162,In_582,In_1722);
nor U2163 (N_2163,In_1920,In_557);
nor U2164 (N_2164,In_1627,In_2261);
xor U2165 (N_2165,In_1346,In_1509);
and U2166 (N_2166,In_1689,In_1117);
and U2167 (N_2167,In_315,In_995);
or U2168 (N_2168,In_193,In_961);
and U2169 (N_2169,In_2384,In_1180);
or U2170 (N_2170,In_1884,In_414);
nor U2171 (N_2171,In_80,In_1412);
xnor U2172 (N_2172,In_1041,In_1321);
nor U2173 (N_2173,In_1519,In_714);
xor U2174 (N_2174,In_2476,In_1995);
nor U2175 (N_2175,In_1460,In_674);
xor U2176 (N_2176,In_206,In_684);
nor U2177 (N_2177,In_1578,In_1823);
nand U2178 (N_2178,In_1057,In_1910);
and U2179 (N_2179,In_645,In_450);
nand U2180 (N_2180,In_1367,In_313);
nand U2181 (N_2181,In_20,In_1339);
nor U2182 (N_2182,In_213,In_2053);
xor U2183 (N_2183,In_1309,In_2409);
xor U2184 (N_2184,In_1761,In_2296);
or U2185 (N_2185,In_365,In_2499);
nand U2186 (N_2186,In_752,In_2117);
nand U2187 (N_2187,In_289,In_753);
nor U2188 (N_2188,In_310,In_81);
and U2189 (N_2189,In_1097,In_228);
nor U2190 (N_2190,In_766,In_2424);
and U2191 (N_2191,In_1563,In_2199);
nand U2192 (N_2192,In_2451,In_1704);
and U2193 (N_2193,In_992,In_180);
xnor U2194 (N_2194,In_995,In_1199);
and U2195 (N_2195,In_1171,In_2308);
nor U2196 (N_2196,In_511,In_2457);
nor U2197 (N_2197,In_2086,In_1366);
nand U2198 (N_2198,In_2208,In_1781);
or U2199 (N_2199,In_1386,In_936);
xor U2200 (N_2200,In_1229,In_2453);
nor U2201 (N_2201,In_109,In_1632);
xor U2202 (N_2202,In_74,In_2216);
nor U2203 (N_2203,In_382,In_476);
xnor U2204 (N_2204,In_1435,In_1192);
xor U2205 (N_2205,In_737,In_1327);
nor U2206 (N_2206,In_733,In_1631);
or U2207 (N_2207,In_2063,In_447);
and U2208 (N_2208,In_399,In_299);
and U2209 (N_2209,In_1691,In_2004);
nor U2210 (N_2210,In_2210,In_1608);
xor U2211 (N_2211,In_94,In_1177);
or U2212 (N_2212,In_198,In_2260);
and U2213 (N_2213,In_2495,In_2376);
and U2214 (N_2214,In_621,In_785);
nor U2215 (N_2215,In_16,In_1916);
nor U2216 (N_2216,In_1827,In_591);
nor U2217 (N_2217,In_1193,In_2374);
nor U2218 (N_2218,In_2354,In_1851);
nand U2219 (N_2219,In_779,In_1785);
xor U2220 (N_2220,In_2294,In_1592);
nand U2221 (N_2221,In_2383,In_266);
and U2222 (N_2222,In_1014,In_2298);
nor U2223 (N_2223,In_2004,In_1409);
and U2224 (N_2224,In_742,In_1100);
nor U2225 (N_2225,In_2237,In_2482);
or U2226 (N_2226,In_2462,In_1860);
or U2227 (N_2227,In_1302,In_364);
nor U2228 (N_2228,In_1519,In_2424);
xnor U2229 (N_2229,In_2239,In_1437);
or U2230 (N_2230,In_2310,In_1686);
nor U2231 (N_2231,In_2022,In_2445);
nor U2232 (N_2232,In_270,In_969);
nor U2233 (N_2233,In_127,In_1052);
or U2234 (N_2234,In_145,In_2040);
nor U2235 (N_2235,In_43,In_1794);
nor U2236 (N_2236,In_1446,In_1339);
and U2237 (N_2237,In_985,In_326);
xnor U2238 (N_2238,In_398,In_956);
xor U2239 (N_2239,In_2038,In_2103);
and U2240 (N_2240,In_1075,In_2350);
and U2241 (N_2241,In_888,In_2468);
or U2242 (N_2242,In_2463,In_679);
and U2243 (N_2243,In_634,In_905);
nand U2244 (N_2244,In_2285,In_369);
nand U2245 (N_2245,In_407,In_2021);
xor U2246 (N_2246,In_243,In_19);
nor U2247 (N_2247,In_1335,In_215);
or U2248 (N_2248,In_2119,In_610);
nand U2249 (N_2249,In_1246,In_131);
or U2250 (N_2250,In_2486,In_665);
and U2251 (N_2251,In_446,In_1343);
nand U2252 (N_2252,In_1775,In_2168);
xor U2253 (N_2253,In_2484,In_646);
or U2254 (N_2254,In_1240,In_154);
or U2255 (N_2255,In_1894,In_666);
nand U2256 (N_2256,In_2068,In_1647);
nand U2257 (N_2257,In_244,In_817);
xor U2258 (N_2258,In_2030,In_1904);
nor U2259 (N_2259,In_1528,In_1883);
nor U2260 (N_2260,In_2173,In_180);
xor U2261 (N_2261,In_1724,In_685);
or U2262 (N_2262,In_2093,In_2386);
and U2263 (N_2263,In_1111,In_2023);
and U2264 (N_2264,In_175,In_1776);
nand U2265 (N_2265,In_21,In_698);
xnor U2266 (N_2266,In_1259,In_872);
and U2267 (N_2267,In_1856,In_758);
nand U2268 (N_2268,In_2050,In_1181);
and U2269 (N_2269,In_1388,In_1392);
xor U2270 (N_2270,In_1863,In_2266);
or U2271 (N_2271,In_2131,In_35);
nor U2272 (N_2272,In_2127,In_3);
nor U2273 (N_2273,In_172,In_2246);
nand U2274 (N_2274,In_314,In_2449);
and U2275 (N_2275,In_1954,In_222);
and U2276 (N_2276,In_907,In_746);
xnor U2277 (N_2277,In_773,In_104);
xor U2278 (N_2278,In_1574,In_2257);
and U2279 (N_2279,In_406,In_1672);
and U2280 (N_2280,In_1412,In_1273);
nand U2281 (N_2281,In_1102,In_470);
nand U2282 (N_2282,In_2,In_54);
and U2283 (N_2283,In_302,In_1552);
or U2284 (N_2284,In_2124,In_2321);
nand U2285 (N_2285,In_922,In_1929);
nand U2286 (N_2286,In_95,In_2251);
nand U2287 (N_2287,In_720,In_543);
and U2288 (N_2288,In_1281,In_20);
nor U2289 (N_2289,In_2354,In_932);
nand U2290 (N_2290,In_551,In_2053);
nand U2291 (N_2291,In_2137,In_1876);
nand U2292 (N_2292,In_2300,In_365);
or U2293 (N_2293,In_559,In_879);
nor U2294 (N_2294,In_835,In_1560);
and U2295 (N_2295,In_881,In_1175);
or U2296 (N_2296,In_1018,In_1230);
nand U2297 (N_2297,In_1839,In_923);
nor U2298 (N_2298,In_1530,In_2253);
or U2299 (N_2299,In_1287,In_1688);
and U2300 (N_2300,In_996,In_173);
xor U2301 (N_2301,In_1538,In_2451);
nor U2302 (N_2302,In_364,In_2182);
and U2303 (N_2303,In_1476,In_1078);
nor U2304 (N_2304,In_338,In_2271);
xor U2305 (N_2305,In_121,In_1033);
nand U2306 (N_2306,In_2212,In_431);
and U2307 (N_2307,In_1650,In_612);
nand U2308 (N_2308,In_2338,In_1798);
nand U2309 (N_2309,In_361,In_1409);
and U2310 (N_2310,In_1747,In_1733);
xnor U2311 (N_2311,In_1179,In_638);
and U2312 (N_2312,In_2448,In_1884);
and U2313 (N_2313,In_95,In_324);
xor U2314 (N_2314,In_54,In_1021);
and U2315 (N_2315,In_767,In_1058);
nand U2316 (N_2316,In_162,In_363);
and U2317 (N_2317,In_1265,In_2055);
or U2318 (N_2318,In_186,In_2044);
or U2319 (N_2319,In_1519,In_725);
nand U2320 (N_2320,In_2479,In_1323);
nand U2321 (N_2321,In_860,In_438);
or U2322 (N_2322,In_2420,In_1454);
and U2323 (N_2323,In_1730,In_525);
and U2324 (N_2324,In_994,In_1320);
nor U2325 (N_2325,In_877,In_639);
nor U2326 (N_2326,In_969,In_1914);
nand U2327 (N_2327,In_1345,In_1755);
and U2328 (N_2328,In_2320,In_918);
nand U2329 (N_2329,In_959,In_1068);
or U2330 (N_2330,In_1589,In_726);
nor U2331 (N_2331,In_1748,In_1507);
and U2332 (N_2332,In_1711,In_1935);
nor U2333 (N_2333,In_379,In_2403);
xor U2334 (N_2334,In_1786,In_2014);
and U2335 (N_2335,In_1971,In_1658);
and U2336 (N_2336,In_1643,In_519);
and U2337 (N_2337,In_156,In_1705);
and U2338 (N_2338,In_1222,In_1473);
xor U2339 (N_2339,In_350,In_1743);
xor U2340 (N_2340,In_1735,In_2127);
nand U2341 (N_2341,In_1334,In_1225);
and U2342 (N_2342,In_2055,In_929);
or U2343 (N_2343,In_773,In_987);
and U2344 (N_2344,In_570,In_1016);
or U2345 (N_2345,In_1493,In_1359);
or U2346 (N_2346,In_1214,In_985);
and U2347 (N_2347,In_1195,In_626);
xor U2348 (N_2348,In_83,In_2060);
or U2349 (N_2349,In_683,In_1838);
and U2350 (N_2350,In_389,In_1071);
xor U2351 (N_2351,In_1450,In_299);
nand U2352 (N_2352,In_580,In_2271);
and U2353 (N_2353,In_455,In_2402);
and U2354 (N_2354,In_1302,In_1138);
or U2355 (N_2355,In_2400,In_2005);
nand U2356 (N_2356,In_1992,In_276);
or U2357 (N_2357,In_785,In_2315);
nand U2358 (N_2358,In_822,In_737);
nor U2359 (N_2359,In_622,In_581);
nand U2360 (N_2360,In_442,In_2252);
nand U2361 (N_2361,In_725,In_1882);
nand U2362 (N_2362,In_991,In_1576);
xnor U2363 (N_2363,In_2263,In_1947);
nor U2364 (N_2364,In_945,In_832);
nor U2365 (N_2365,In_2257,In_1513);
nand U2366 (N_2366,In_1890,In_1748);
nand U2367 (N_2367,In_1141,In_195);
and U2368 (N_2368,In_439,In_1087);
or U2369 (N_2369,In_1792,In_2416);
nand U2370 (N_2370,In_1871,In_1943);
nor U2371 (N_2371,In_372,In_1195);
nand U2372 (N_2372,In_975,In_1692);
nor U2373 (N_2373,In_1619,In_2164);
or U2374 (N_2374,In_459,In_2174);
or U2375 (N_2375,In_1586,In_819);
nor U2376 (N_2376,In_638,In_215);
or U2377 (N_2377,In_1580,In_304);
and U2378 (N_2378,In_74,In_1388);
nand U2379 (N_2379,In_231,In_1503);
nor U2380 (N_2380,In_1819,In_2420);
and U2381 (N_2381,In_2321,In_134);
and U2382 (N_2382,In_286,In_2489);
or U2383 (N_2383,In_2364,In_1702);
xor U2384 (N_2384,In_580,In_1498);
and U2385 (N_2385,In_2303,In_470);
nand U2386 (N_2386,In_174,In_2391);
nand U2387 (N_2387,In_405,In_1739);
and U2388 (N_2388,In_2108,In_640);
xor U2389 (N_2389,In_2289,In_204);
and U2390 (N_2390,In_1715,In_1400);
nor U2391 (N_2391,In_18,In_2048);
nor U2392 (N_2392,In_2028,In_2447);
xor U2393 (N_2393,In_96,In_2042);
nand U2394 (N_2394,In_1879,In_1699);
and U2395 (N_2395,In_1610,In_2045);
or U2396 (N_2396,In_466,In_2102);
nand U2397 (N_2397,In_2209,In_2220);
nor U2398 (N_2398,In_2250,In_2038);
and U2399 (N_2399,In_2296,In_2139);
nand U2400 (N_2400,In_1002,In_531);
or U2401 (N_2401,In_657,In_2492);
or U2402 (N_2402,In_1653,In_1714);
xor U2403 (N_2403,In_1348,In_1848);
and U2404 (N_2404,In_1016,In_178);
and U2405 (N_2405,In_1378,In_2059);
or U2406 (N_2406,In_1675,In_1027);
nor U2407 (N_2407,In_1236,In_182);
and U2408 (N_2408,In_2480,In_772);
nor U2409 (N_2409,In_2172,In_94);
or U2410 (N_2410,In_29,In_1486);
nor U2411 (N_2411,In_105,In_2395);
and U2412 (N_2412,In_1503,In_865);
nor U2413 (N_2413,In_392,In_928);
nand U2414 (N_2414,In_1124,In_2327);
and U2415 (N_2415,In_1440,In_1631);
xor U2416 (N_2416,In_1901,In_1750);
and U2417 (N_2417,In_1583,In_168);
nor U2418 (N_2418,In_2164,In_44);
or U2419 (N_2419,In_1764,In_364);
or U2420 (N_2420,In_1416,In_1891);
xnor U2421 (N_2421,In_1528,In_1334);
nand U2422 (N_2422,In_2442,In_1726);
nor U2423 (N_2423,In_2412,In_1996);
xor U2424 (N_2424,In_2234,In_2285);
and U2425 (N_2425,In_2164,In_351);
and U2426 (N_2426,In_1375,In_1317);
and U2427 (N_2427,In_1798,In_2011);
and U2428 (N_2428,In_2202,In_2209);
xnor U2429 (N_2429,In_1418,In_2328);
and U2430 (N_2430,In_597,In_281);
and U2431 (N_2431,In_96,In_817);
nor U2432 (N_2432,In_816,In_1597);
nand U2433 (N_2433,In_2032,In_211);
and U2434 (N_2434,In_713,In_1885);
and U2435 (N_2435,In_153,In_1497);
xnor U2436 (N_2436,In_2201,In_1252);
xor U2437 (N_2437,In_1942,In_670);
and U2438 (N_2438,In_1729,In_193);
nor U2439 (N_2439,In_2494,In_1028);
and U2440 (N_2440,In_320,In_977);
xor U2441 (N_2441,In_218,In_1850);
xnor U2442 (N_2442,In_2241,In_490);
and U2443 (N_2443,In_2334,In_996);
or U2444 (N_2444,In_1545,In_1045);
nand U2445 (N_2445,In_2186,In_1331);
nand U2446 (N_2446,In_688,In_821);
or U2447 (N_2447,In_650,In_193);
xnor U2448 (N_2448,In_273,In_84);
xor U2449 (N_2449,In_1350,In_1013);
and U2450 (N_2450,In_2357,In_597);
xor U2451 (N_2451,In_94,In_1095);
or U2452 (N_2452,In_592,In_1504);
or U2453 (N_2453,In_648,In_338);
and U2454 (N_2454,In_1596,In_2484);
nor U2455 (N_2455,In_435,In_2434);
or U2456 (N_2456,In_2015,In_1753);
xor U2457 (N_2457,In_1248,In_2313);
xnor U2458 (N_2458,In_1968,In_1682);
or U2459 (N_2459,In_1182,In_2297);
and U2460 (N_2460,In_2366,In_1570);
and U2461 (N_2461,In_502,In_1971);
or U2462 (N_2462,In_2050,In_1165);
or U2463 (N_2463,In_993,In_404);
and U2464 (N_2464,In_669,In_1383);
and U2465 (N_2465,In_1268,In_924);
or U2466 (N_2466,In_1921,In_422);
or U2467 (N_2467,In_1874,In_86);
and U2468 (N_2468,In_121,In_1427);
and U2469 (N_2469,In_1629,In_2168);
xor U2470 (N_2470,In_1500,In_62);
xnor U2471 (N_2471,In_688,In_1449);
xnor U2472 (N_2472,In_611,In_1919);
xor U2473 (N_2473,In_145,In_309);
xor U2474 (N_2474,In_504,In_1259);
and U2475 (N_2475,In_1249,In_57);
nor U2476 (N_2476,In_69,In_1689);
or U2477 (N_2477,In_1855,In_624);
and U2478 (N_2478,In_2219,In_1072);
or U2479 (N_2479,In_2142,In_1478);
and U2480 (N_2480,In_1126,In_640);
nand U2481 (N_2481,In_2258,In_188);
nand U2482 (N_2482,In_1543,In_1322);
and U2483 (N_2483,In_2480,In_961);
and U2484 (N_2484,In_762,In_1995);
and U2485 (N_2485,In_26,In_1765);
nor U2486 (N_2486,In_1480,In_1376);
or U2487 (N_2487,In_1202,In_1587);
or U2488 (N_2488,In_2047,In_1155);
xnor U2489 (N_2489,In_529,In_944);
nor U2490 (N_2490,In_331,In_1825);
nor U2491 (N_2491,In_2369,In_658);
or U2492 (N_2492,In_984,In_922);
or U2493 (N_2493,In_2451,In_1607);
xnor U2494 (N_2494,In_2184,In_619);
nor U2495 (N_2495,In_1072,In_542);
nor U2496 (N_2496,In_1404,In_1679);
or U2497 (N_2497,In_2050,In_541);
xor U2498 (N_2498,In_1609,In_2105);
nand U2499 (N_2499,In_1291,In_2184);
or U2500 (N_2500,In_910,In_2409);
xor U2501 (N_2501,In_146,In_174);
xor U2502 (N_2502,In_2020,In_1115);
or U2503 (N_2503,In_1355,In_660);
nor U2504 (N_2504,In_679,In_532);
nor U2505 (N_2505,In_1520,In_247);
nor U2506 (N_2506,In_878,In_1125);
and U2507 (N_2507,In_607,In_308);
xor U2508 (N_2508,In_347,In_1110);
xor U2509 (N_2509,In_1803,In_1728);
and U2510 (N_2510,In_42,In_2215);
nor U2511 (N_2511,In_1953,In_593);
or U2512 (N_2512,In_721,In_2306);
and U2513 (N_2513,In_2008,In_1739);
nor U2514 (N_2514,In_1199,In_777);
nand U2515 (N_2515,In_1171,In_997);
or U2516 (N_2516,In_627,In_270);
or U2517 (N_2517,In_642,In_745);
and U2518 (N_2518,In_1439,In_1343);
nor U2519 (N_2519,In_428,In_1227);
nand U2520 (N_2520,In_612,In_229);
nor U2521 (N_2521,In_2460,In_1661);
nand U2522 (N_2522,In_111,In_1039);
or U2523 (N_2523,In_1631,In_1708);
and U2524 (N_2524,In_2170,In_268);
and U2525 (N_2525,In_2152,In_776);
xnor U2526 (N_2526,In_448,In_672);
and U2527 (N_2527,In_2438,In_1942);
or U2528 (N_2528,In_950,In_135);
xor U2529 (N_2529,In_199,In_125);
nand U2530 (N_2530,In_511,In_2315);
or U2531 (N_2531,In_731,In_302);
nand U2532 (N_2532,In_153,In_577);
xor U2533 (N_2533,In_1668,In_1754);
nand U2534 (N_2534,In_2440,In_2365);
nand U2535 (N_2535,In_81,In_505);
nor U2536 (N_2536,In_7,In_1201);
nor U2537 (N_2537,In_645,In_1451);
or U2538 (N_2538,In_727,In_1798);
xor U2539 (N_2539,In_105,In_1657);
nand U2540 (N_2540,In_214,In_395);
and U2541 (N_2541,In_536,In_762);
xor U2542 (N_2542,In_2037,In_317);
nand U2543 (N_2543,In_2177,In_2124);
and U2544 (N_2544,In_1334,In_2118);
and U2545 (N_2545,In_1553,In_2314);
nand U2546 (N_2546,In_196,In_684);
nor U2547 (N_2547,In_1931,In_1696);
nor U2548 (N_2548,In_912,In_1718);
nor U2549 (N_2549,In_235,In_1967);
or U2550 (N_2550,In_915,In_611);
nor U2551 (N_2551,In_2149,In_873);
nor U2552 (N_2552,In_288,In_1799);
or U2553 (N_2553,In_334,In_1311);
or U2554 (N_2554,In_1843,In_645);
or U2555 (N_2555,In_1676,In_78);
and U2556 (N_2556,In_249,In_1347);
nor U2557 (N_2557,In_1810,In_30);
nand U2558 (N_2558,In_654,In_1072);
and U2559 (N_2559,In_2245,In_2107);
and U2560 (N_2560,In_307,In_691);
and U2561 (N_2561,In_558,In_988);
nand U2562 (N_2562,In_1019,In_1896);
nand U2563 (N_2563,In_1697,In_1077);
nor U2564 (N_2564,In_117,In_734);
and U2565 (N_2565,In_1510,In_1717);
xor U2566 (N_2566,In_1094,In_2460);
nor U2567 (N_2567,In_2081,In_2489);
nor U2568 (N_2568,In_356,In_877);
nand U2569 (N_2569,In_1354,In_2018);
xor U2570 (N_2570,In_2292,In_355);
and U2571 (N_2571,In_2389,In_24);
xnor U2572 (N_2572,In_1343,In_796);
nand U2573 (N_2573,In_484,In_1471);
xnor U2574 (N_2574,In_2293,In_1026);
or U2575 (N_2575,In_2458,In_2133);
nor U2576 (N_2576,In_1740,In_1223);
and U2577 (N_2577,In_2323,In_663);
nor U2578 (N_2578,In_379,In_2445);
nand U2579 (N_2579,In_2176,In_1583);
or U2580 (N_2580,In_1029,In_2131);
nor U2581 (N_2581,In_2480,In_685);
and U2582 (N_2582,In_588,In_2384);
nor U2583 (N_2583,In_1732,In_2070);
nand U2584 (N_2584,In_2013,In_106);
nand U2585 (N_2585,In_2118,In_406);
nand U2586 (N_2586,In_2253,In_881);
xor U2587 (N_2587,In_179,In_2226);
nor U2588 (N_2588,In_1494,In_1584);
and U2589 (N_2589,In_1151,In_1562);
xnor U2590 (N_2590,In_1676,In_1541);
and U2591 (N_2591,In_421,In_883);
nand U2592 (N_2592,In_1644,In_713);
or U2593 (N_2593,In_992,In_1260);
nor U2594 (N_2594,In_2009,In_1510);
nor U2595 (N_2595,In_974,In_1429);
or U2596 (N_2596,In_529,In_1609);
nand U2597 (N_2597,In_1306,In_2413);
nor U2598 (N_2598,In_1554,In_101);
and U2599 (N_2599,In_2247,In_83);
xnor U2600 (N_2600,In_1666,In_2489);
or U2601 (N_2601,In_1024,In_398);
xor U2602 (N_2602,In_2198,In_725);
and U2603 (N_2603,In_949,In_168);
nand U2604 (N_2604,In_470,In_1611);
and U2605 (N_2605,In_1577,In_1913);
nand U2606 (N_2606,In_507,In_2398);
xnor U2607 (N_2607,In_1390,In_2330);
nor U2608 (N_2608,In_1411,In_1761);
nand U2609 (N_2609,In_1569,In_1223);
and U2610 (N_2610,In_1661,In_1472);
nor U2611 (N_2611,In_691,In_2214);
xnor U2612 (N_2612,In_451,In_527);
xor U2613 (N_2613,In_151,In_807);
nor U2614 (N_2614,In_1596,In_333);
nor U2615 (N_2615,In_1949,In_933);
or U2616 (N_2616,In_134,In_241);
xnor U2617 (N_2617,In_2156,In_97);
nor U2618 (N_2618,In_1675,In_2237);
nand U2619 (N_2619,In_718,In_1648);
xor U2620 (N_2620,In_1316,In_1112);
xor U2621 (N_2621,In_2,In_927);
or U2622 (N_2622,In_1666,In_1980);
and U2623 (N_2623,In_89,In_868);
nor U2624 (N_2624,In_1123,In_1719);
nor U2625 (N_2625,In_999,In_2136);
and U2626 (N_2626,In_203,In_2365);
or U2627 (N_2627,In_1015,In_917);
or U2628 (N_2628,In_250,In_2267);
or U2629 (N_2629,In_897,In_1897);
nand U2630 (N_2630,In_1012,In_1451);
nand U2631 (N_2631,In_2256,In_886);
nand U2632 (N_2632,In_698,In_366);
or U2633 (N_2633,In_1193,In_1500);
and U2634 (N_2634,In_884,In_1965);
nor U2635 (N_2635,In_467,In_2159);
or U2636 (N_2636,In_941,In_1409);
nor U2637 (N_2637,In_1921,In_745);
nand U2638 (N_2638,In_49,In_1318);
xor U2639 (N_2639,In_2288,In_1332);
nor U2640 (N_2640,In_1591,In_1961);
nand U2641 (N_2641,In_1557,In_1716);
xnor U2642 (N_2642,In_664,In_1394);
nand U2643 (N_2643,In_961,In_647);
and U2644 (N_2644,In_873,In_646);
and U2645 (N_2645,In_1696,In_502);
xnor U2646 (N_2646,In_66,In_899);
xor U2647 (N_2647,In_753,In_1422);
nor U2648 (N_2648,In_1530,In_1527);
nor U2649 (N_2649,In_162,In_2227);
xor U2650 (N_2650,In_407,In_2086);
nand U2651 (N_2651,In_1823,In_2466);
nor U2652 (N_2652,In_11,In_1003);
nand U2653 (N_2653,In_1772,In_451);
xor U2654 (N_2654,In_288,In_1290);
nand U2655 (N_2655,In_2040,In_1443);
nor U2656 (N_2656,In_1851,In_621);
nand U2657 (N_2657,In_2391,In_823);
nor U2658 (N_2658,In_2236,In_2197);
nand U2659 (N_2659,In_126,In_627);
and U2660 (N_2660,In_1837,In_442);
nand U2661 (N_2661,In_1137,In_2175);
xnor U2662 (N_2662,In_931,In_854);
nand U2663 (N_2663,In_779,In_18);
nor U2664 (N_2664,In_1809,In_444);
or U2665 (N_2665,In_1020,In_2379);
or U2666 (N_2666,In_2127,In_793);
nor U2667 (N_2667,In_247,In_2065);
and U2668 (N_2668,In_542,In_772);
xor U2669 (N_2669,In_157,In_1309);
nor U2670 (N_2670,In_1879,In_1792);
nand U2671 (N_2671,In_2227,In_1158);
xnor U2672 (N_2672,In_13,In_2041);
nor U2673 (N_2673,In_1395,In_523);
nor U2674 (N_2674,In_1738,In_1778);
nor U2675 (N_2675,In_684,In_988);
xor U2676 (N_2676,In_2075,In_74);
nand U2677 (N_2677,In_1747,In_231);
nand U2678 (N_2678,In_1040,In_2286);
xnor U2679 (N_2679,In_1713,In_2076);
xor U2680 (N_2680,In_998,In_58);
and U2681 (N_2681,In_177,In_1324);
or U2682 (N_2682,In_2305,In_2321);
and U2683 (N_2683,In_493,In_1049);
xor U2684 (N_2684,In_1157,In_1832);
nor U2685 (N_2685,In_1911,In_1519);
and U2686 (N_2686,In_1762,In_1416);
and U2687 (N_2687,In_2480,In_1503);
and U2688 (N_2688,In_2094,In_1321);
or U2689 (N_2689,In_608,In_1830);
nor U2690 (N_2690,In_1851,In_148);
nand U2691 (N_2691,In_132,In_2112);
nand U2692 (N_2692,In_1483,In_1857);
nand U2693 (N_2693,In_587,In_1957);
nand U2694 (N_2694,In_120,In_1480);
nor U2695 (N_2695,In_305,In_1463);
nand U2696 (N_2696,In_2109,In_85);
or U2697 (N_2697,In_714,In_1050);
or U2698 (N_2698,In_1280,In_704);
nand U2699 (N_2699,In_2212,In_2416);
xnor U2700 (N_2700,In_2188,In_471);
and U2701 (N_2701,In_2400,In_1807);
nand U2702 (N_2702,In_1727,In_2365);
xnor U2703 (N_2703,In_1669,In_1872);
or U2704 (N_2704,In_1388,In_1412);
and U2705 (N_2705,In_1268,In_1495);
xor U2706 (N_2706,In_2460,In_1632);
nand U2707 (N_2707,In_2061,In_1891);
xor U2708 (N_2708,In_2382,In_718);
and U2709 (N_2709,In_196,In_444);
or U2710 (N_2710,In_2418,In_1573);
xnor U2711 (N_2711,In_1421,In_1885);
and U2712 (N_2712,In_397,In_400);
nand U2713 (N_2713,In_575,In_105);
nor U2714 (N_2714,In_484,In_2037);
or U2715 (N_2715,In_1344,In_1317);
xnor U2716 (N_2716,In_2398,In_108);
and U2717 (N_2717,In_204,In_1912);
nor U2718 (N_2718,In_490,In_416);
and U2719 (N_2719,In_2074,In_2034);
nor U2720 (N_2720,In_2354,In_2156);
and U2721 (N_2721,In_2389,In_321);
xor U2722 (N_2722,In_1905,In_1582);
and U2723 (N_2723,In_2423,In_1029);
or U2724 (N_2724,In_687,In_2431);
and U2725 (N_2725,In_598,In_1787);
nand U2726 (N_2726,In_1654,In_79);
and U2727 (N_2727,In_1612,In_640);
xnor U2728 (N_2728,In_187,In_64);
nor U2729 (N_2729,In_1070,In_860);
nand U2730 (N_2730,In_525,In_2277);
or U2731 (N_2731,In_1221,In_1151);
and U2732 (N_2732,In_1656,In_2230);
or U2733 (N_2733,In_943,In_1405);
and U2734 (N_2734,In_88,In_1663);
and U2735 (N_2735,In_2013,In_1309);
nand U2736 (N_2736,In_2487,In_2116);
or U2737 (N_2737,In_632,In_683);
and U2738 (N_2738,In_2112,In_1757);
nand U2739 (N_2739,In_1208,In_2270);
or U2740 (N_2740,In_2210,In_244);
and U2741 (N_2741,In_1216,In_1452);
and U2742 (N_2742,In_747,In_2337);
nand U2743 (N_2743,In_1990,In_2414);
and U2744 (N_2744,In_759,In_2292);
nand U2745 (N_2745,In_1733,In_1049);
xnor U2746 (N_2746,In_641,In_1624);
nor U2747 (N_2747,In_1247,In_1515);
nor U2748 (N_2748,In_1768,In_813);
nor U2749 (N_2749,In_2236,In_511);
xor U2750 (N_2750,In_536,In_1037);
xor U2751 (N_2751,In_1783,In_806);
nand U2752 (N_2752,In_1620,In_699);
nand U2753 (N_2753,In_908,In_1255);
nand U2754 (N_2754,In_1972,In_827);
nand U2755 (N_2755,In_2124,In_155);
xor U2756 (N_2756,In_1457,In_2300);
nor U2757 (N_2757,In_875,In_1949);
nand U2758 (N_2758,In_811,In_1097);
or U2759 (N_2759,In_601,In_2184);
nor U2760 (N_2760,In_842,In_107);
nand U2761 (N_2761,In_1958,In_144);
nor U2762 (N_2762,In_1321,In_1628);
nor U2763 (N_2763,In_1239,In_466);
nor U2764 (N_2764,In_1632,In_1122);
nand U2765 (N_2765,In_176,In_670);
or U2766 (N_2766,In_2313,In_1477);
nand U2767 (N_2767,In_1363,In_1228);
nand U2768 (N_2768,In_603,In_1365);
and U2769 (N_2769,In_2463,In_863);
or U2770 (N_2770,In_1604,In_48);
nor U2771 (N_2771,In_1223,In_2078);
nand U2772 (N_2772,In_438,In_1918);
xnor U2773 (N_2773,In_2377,In_2403);
and U2774 (N_2774,In_1023,In_654);
and U2775 (N_2775,In_1400,In_1800);
nor U2776 (N_2776,In_1448,In_308);
and U2777 (N_2777,In_2479,In_2002);
nor U2778 (N_2778,In_1056,In_323);
or U2779 (N_2779,In_2332,In_252);
and U2780 (N_2780,In_658,In_2448);
nor U2781 (N_2781,In_2137,In_1096);
xnor U2782 (N_2782,In_2449,In_1198);
nand U2783 (N_2783,In_765,In_2008);
or U2784 (N_2784,In_1264,In_1777);
or U2785 (N_2785,In_1861,In_90);
xnor U2786 (N_2786,In_591,In_447);
nor U2787 (N_2787,In_1542,In_2246);
xor U2788 (N_2788,In_873,In_949);
or U2789 (N_2789,In_1,In_595);
xor U2790 (N_2790,In_672,In_247);
xnor U2791 (N_2791,In_2126,In_813);
nor U2792 (N_2792,In_2313,In_1451);
or U2793 (N_2793,In_498,In_2284);
and U2794 (N_2794,In_191,In_2251);
or U2795 (N_2795,In_1035,In_1796);
nor U2796 (N_2796,In_1259,In_628);
nor U2797 (N_2797,In_1254,In_794);
nand U2798 (N_2798,In_226,In_711);
nor U2799 (N_2799,In_1732,In_1745);
xor U2800 (N_2800,In_1913,In_1876);
and U2801 (N_2801,In_1515,In_422);
xnor U2802 (N_2802,In_299,In_20);
nand U2803 (N_2803,In_373,In_1306);
nor U2804 (N_2804,In_209,In_138);
nor U2805 (N_2805,In_1419,In_1063);
nand U2806 (N_2806,In_750,In_2323);
xnor U2807 (N_2807,In_1092,In_847);
and U2808 (N_2808,In_1756,In_6);
or U2809 (N_2809,In_736,In_1972);
nor U2810 (N_2810,In_1667,In_1240);
and U2811 (N_2811,In_1630,In_2224);
nor U2812 (N_2812,In_2018,In_1698);
xnor U2813 (N_2813,In_1267,In_1112);
nand U2814 (N_2814,In_1402,In_484);
nor U2815 (N_2815,In_2037,In_1339);
nor U2816 (N_2816,In_1855,In_2285);
or U2817 (N_2817,In_1246,In_2205);
xor U2818 (N_2818,In_907,In_1795);
nand U2819 (N_2819,In_150,In_603);
xor U2820 (N_2820,In_911,In_1934);
nor U2821 (N_2821,In_324,In_2271);
or U2822 (N_2822,In_158,In_569);
or U2823 (N_2823,In_110,In_550);
nand U2824 (N_2824,In_1127,In_1597);
xnor U2825 (N_2825,In_1533,In_962);
and U2826 (N_2826,In_2127,In_183);
xor U2827 (N_2827,In_523,In_1408);
nand U2828 (N_2828,In_308,In_2447);
nand U2829 (N_2829,In_802,In_330);
xnor U2830 (N_2830,In_287,In_2146);
xor U2831 (N_2831,In_1765,In_744);
nand U2832 (N_2832,In_78,In_1737);
nand U2833 (N_2833,In_1566,In_712);
nor U2834 (N_2834,In_2358,In_353);
or U2835 (N_2835,In_2438,In_2228);
nand U2836 (N_2836,In_2426,In_169);
nand U2837 (N_2837,In_1522,In_302);
or U2838 (N_2838,In_2287,In_1715);
or U2839 (N_2839,In_1089,In_2087);
xnor U2840 (N_2840,In_1453,In_2375);
nor U2841 (N_2841,In_2002,In_1208);
and U2842 (N_2842,In_1701,In_1651);
nor U2843 (N_2843,In_645,In_1104);
and U2844 (N_2844,In_857,In_2489);
nand U2845 (N_2845,In_1013,In_1830);
and U2846 (N_2846,In_2316,In_539);
nand U2847 (N_2847,In_51,In_282);
nand U2848 (N_2848,In_1305,In_134);
xnor U2849 (N_2849,In_1374,In_2138);
and U2850 (N_2850,In_2225,In_1288);
and U2851 (N_2851,In_1580,In_297);
nand U2852 (N_2852,In_1424,In_863);
nor U2853 (N_2853,In_1187,In_1083);
or U2854 (N_2854,In_1204,In_1569);
nor U2855 (N_2855,In_2295,In_750);
xor U2856 (N_2856,In_1884,In_626);
and U2857 (N_2857,In_1806,In_2408);
and U2858 (N_2858,In_1312,In_868);
and U2859 (N_2859,In_2336,In_1916);
nand U2860 (N_2860,In_1292,In_661);
nor U2861 (N_2861,In_492,In_632);
or U2862 (N_2862,In_94,In_2343);
nand U2863 (N_2863,In_1758,In_2107);
xor U2864 (N_2864,In_1297,In_2482);
or U2865 (N_2865,In_971,In_240);
and U2866 (N_2866,In_1196,In_973);
nor U2867 (N_2867,In_1233,In_2069);
xor U2868 (N_2868,In_2169,In_976);
or U2869 (N_2869,In_2023,In_1554);
nand U2870 (N_2870,In_850,In_895);
or U2871 (N_2871,In_617,In_21);
or U2872 (N_2872,In_681,In_1934);
xnor U2873 (N_2873,In_312,In_1827);
and U2874 (N_2874,In_1183,In_2232);
nand U2875 (N_2875,In_643,In_336);
nand U2876 (N_2876,In_2485,In_1425);
and U2877 (N_2877,In_2285,In_552);
nor U2878 (N_2878,In_1490,In_1960);
xor U2879 (N_2879,In_494,In_2359);
nor U2880 (N_2880,In_2065,In_388);
or U2881 (N_2881,In_129,In_77);
nor U2882 (N_2882,In_305,In_1277);
or U2883 (N_2883,In_1513,In_157);
nand U2884 (N_2884,In_1524,In_1371);
and U2885 (N_2885,In_1341,In_921);
xnor U2886 (N_2886,In_1441,In_2201);
nor U2887 (N_2887,In_450,In_1513);
nor U2888 (N_2888,In_701,In_1831);
and U2889 (N_2889,In_442,In_1849);
or U2890 (N_2890,In_872,In_2486);
nor U2891 (N_2891,In_940,In_454);
nand U2892 (N_2892,In_2027,In_1873);
nand U2893 (N_2893,In_786,In_840);
or U2894 (N_2894,In_1463,In_1258);
nand U2895 (N_2895,In_200,In_1282);
xnor U2896 (N_2896,In_819,In_2249);
nor U2897 (N_2897,In_1781,In_1398);
or U2898 (N_2898,In_1581,In_1482);
nand U2899 (N_2899,In_1154,In_1416);
nor U2900 (N_2900,In_1313,In_720);
nor U2901 (N_2901,In_1449,In_902);
nor U2902 (N_2902,In_1063,In_1617);
nand U2903 (N_2903,In_233,In_564);
or U2904 (N_2904,In_1751,In_488);
or U2905 (N_2905,In_440,In_1352);
nor U2906 (N_2906,In_2178,In_926);
or U2907 (N_2907,In_1829,In_1069);
and U2908 (N_2908,In_352,In_1121);
and U2909 (N_2909,In_2232,In_1819);
xor U2910 (N_2910,In_584,In_183);
nor U2911 (N_2911,In_972,In_1404);
nand U2912 (N_2912,In_1033,In_682);
or U2913 (N_2913,In_2406,In_1081);
or U2914 (N_2914,In_1077,In_554);
nor U2915 (N_2915,In_181,In_1810);
xnor U2916 (N_2916,In_27,In_197);
and U2917 (N_2917,In_1660,In_636);
or U2918 (N_2918,In_160,In_1918);
and U2919 (N_2919,In_1988,In_418);
and U2920 (N_2920,In_1609,In_298);
nor U2921 (N_2921,In_1050,In_848);
nor U2922 (N_2922,In_1481,In_239);
nand U2923 (N_2923,In_1283,In_254);
nor U2924 (N_2924,In_1784,In_1782);
nor U2925 (N_2925,In_127,In_1002);
nand U2926 (N_2926,In_102,In_22);
xnor U2927 (N_2927,In_1667,In_767);
xnor U2928 (N_2928,In_103,In_1925);
nand U2929 (N_2929,In_784,In_190);
or U2930 (N_2930,In_1364,In_524);
nor U2931 (N_2931,In_2017,In_990);
and U2932 (N_2932,In_1883,In_1667);
or U2933 (N_2933,In_1795,In_1869);
or U2934 (N_2934,In_1737,In_320);
nand U2935 (N_2935,In_828,In_2268);
nand U2936 (N_2936,In_2434,In_2379);
nor U2937 (N_2937,In_1383,In_1525);
nor U2938 (N_2938,In_300,In_2144);
xnor U2939 (N_2939,In_974,In_1971);
xor U2940 (N_2940,In_1657,In_328);
or U2941 (N_2941,In_2060,In_1409);
or U2942 (N_2942,In_660,In_39);
nand U2943 (N_2943,In_343,In_1649);
nor U2944 (N_2944,In_1784,In_1861);
nand U2945 (N_2945,In_2339,In_337);
or U2946 (N_2946,In_707,In_157);
nor U2947 (N_2947,In_707,In_84);
nand U2948 (N_2948,In_713,In_884);
xor U2949 (N_2949,In_357,In_488);
nand U2950 (N_2950,In_1416,In_2393);
nor U2951 (N_2951,In_1428,In_458);
nand U2952 (N_2952,In_1576,In_1358);
xor U2953 (N_2953,In_1724,In_2333);
or U2954 (N_2954,In_919,In_1062);
or U2955 (N_2955,In_1403,In_1491);
nor U2956 (N_2956,In_2196,In_672);
nor U2957 (N_2957,In_1244,In_605);
or U2958 (N_2958,In_2376,In_1938);
or U2959 (N_2959,In_2361,In_1322);
or U2960 (N_2960,In_459,In_2235);
nand U2961 (N_2961,In_1653,In_2469);
xor U2962 (N_2962,In_2111,In_1844);
xnor U2963 (N_2963,In_1590,In_1278);
or U2964 (N_2964,In_223,In_1986);
xnor U2965 (N_2965,In_2190,In_352);
nor U2966 (N_2966,In_863,In_1453);
nor U2967 (N_2967,In_1647,In_519);
and U2968 (N_2968,In_1638,In_1059);
nand U2969 (N_2969,In_360,In_2056);
or U2970 (N_2970,In_1533,In_2078);
and U2971 (N_2971,In_632,In_1238);
or U2972 (N_2972,In_343,In_847);
nor U2973 (N_2973,In_2201,In_439);
xnor U2974 (N_2974,In_2175,In_852);
xnor U2975 (N_2975,In_1391,In_1518);
nor U2976 (N_2976,In_889,In_477);
xnor U2977 (N_2977,In_1298,In_1641);
xor U2978 (N_2978,In_968,In_276);
and U2979 (N_2979,In_1341,In_1809);
nand U2980 (N_2980,In_434,In_708);
or U2981 (N_2981,In_1885,In_723);
nor U2982 (N_2982,In_1337,In_1012);
xnor U2983 (N_2983,In_957,In_2329);
nor U2984 (N_2984,In_1397,In_864);
and U2985 (N_2985,In_871,In_914);
or U2986 (N_2986,In_8,In_2253);
or U2987 (N_2987,In_501,In_1809);
xnor U2988 (N_2988,In_1102,In_388);
or U2989 (N_2989,In_2105,In_1720);
and U2990 (N_2990,In_1408,In_1373);
xnor U2991 (N_2991,In_941,In_1416);
nand U2992 (N_2992,In_316,In_1129);
and U2993 (N_2993,In_1144,In_93);
nor U2994 (N_2994,In_1874,In_913);
and U2995 (N_2995,In_433,In_2397);
nand U2996 (N_2996,In_664,In_1530);
nand U2997 (N_2997,In_2389,In_2314);
and U2998 (N_2998,In_2027,In_858);
xnor U2999 (N_2999,In_1503,In_1706);
xor U3000 (N_3000,In_1404,In_1984);
xor U3001 (N_3001,In_1456,In_378);
or U3002 (N_3002,In_2203,In_1183);
and U3003 (N_3003,In_1678,In_1342);
and U3004 (N_3004,In_312,In_1434);
and U3005 (N_3005,In_877,In_438);
and U3006 (N_3006,In_1135,In_312);
nor U3007 (N_3007,In_2385,In_224);
xnor U3008 (N_3008,In_213,In_1547);
xor U3009 (N_3009,In_511,In_822);
nor U3010 (N_3010,In_1981,In_1440);
xor U3011 (N_3011,In_2151,In_283);
nand U3012 (N_3012,In_1216,In_2171);
nand U3013 (N_3013,In_659,In_72);
xor U3014 (N_3014,In_2246,In_2187);
nand U3015 (N_3015,In_2009,In_1288);
nor U3016 (N_3016,In_2113,In_2140);
and U3017 (N_3017,In_1254,In_672);
nand U3018 (N_3018,In_1839,In_2186);
and U3019 (N_3019,In_621,In_1545);
nor U3020 (N_3020,In_322,In_1565);
xnor U3021 (N_3021,In_894,In_452);
nor U3022 (N_3022,In_682,In_1491);
and U3023 (N_3023,In_1602,In_795);
or U3024 (N_3024,In_2496,In_2452);
and U3025 (N_3025,In_2064,In_817);
and U3026 (N_3026,In_1813,In_2052);
or U3027 (N_3027,In_1632,In_458);
nand U3028 (N_3028,In_2291,In_737);
nand U3029 (N_3029,In_2331,In_2134);
nand U3030 (N_3030,In_1402,In_1825);
xor U3031 (N_3031,In_811,In_2025);
or U3032 (N_3032,In_865,In_2469);
nand U3033 (N_3033,In_896,In_1968);
nand U3034 (N_3034,In_2438,In_1783);
and U3035 (N_3035,In_1763,In_228);
nor U3036 (N_3036,In_2360,In_257);
or U3037 (N_3037,In_1049,In_1730);
and U3038 (N_3038,In_155,In_382);
nand U3039 (N_3039,In_166,In_438);
and U3040 (N_3040,In_2381,In_31);
or U3041 (N_3041,In_1296,In_1687);
or U3042 (N_3042,In_489,In_60);
nand U3043 (N_3043,In_890,In_27);
nand U3044 (N_3044,In_372,In_886);
or U3045 (N_3045,In_554,In_1100);
nand U3046 (N_3046,In_301,In_1264);
and U3047 (N_3047,In_402,In_35);
xnor U3048 (N_3048,In_507,In_2198);
or U3049 (N_3049,In_1587,In_409);
nor U3050 (N_3050,In_700,In_1548);
nand U3051 (N_3051,In_788,In_81);
and U3052 (N_3052,In_1553,In_1202);
xor U3053 (N_3053,In_673,In_1959);
xnor U3054 (N_3054,In_1844,In_1454);
xor U3055 (N_3055,In_1972,In_955);
and U3056 (N_3056,In_550,In_181);
xnor U3057 (N_3057,In_2373,In_1844);
nand U3058 (N_3058,In_739,In_521);
or U3059 (N_3059,In_287,In_1871);
nand U3060 (N_3060,In_34,In_158);
or U3061 (N_3061,In_2456,In_27);
nor U3062 (N_3062,In_987,In_1532);
nor U3063 (N_3063,In_1016,In_254);
nand U3064 (N_3064,In_1347,In_573);
xnor U3065 (N_3065,In_2011,In_2314);
nand U3066 (N_3066,In_357,In_2148);
or U3067 (N_3067,In_592,In_2311);
or U3068 (N_3068,In_1654,In_1293);
nor U3069 (N_3069,In_1796,In_2322);
or U3070 (N_3070,In_1365,In_2380);
xnor U3071 (N_3071,In_521,In_1025);
or U3072 (N_3072,In_244,In_2171);
nand U3073 (N_3073,In_2459,In_475);
and U3074 (N_3074,In_1353,In_1433);
and U3075 (N_3075,In_309,In_327);
or U3076 (N_3076,In_247,In_158);
and U3077 (N_3077,In_240,In_1357);
xnor U3078 (N_3078,In_240,In_2022);
or U3079 (N_3079,In_88,In_1798);
nor U3080 (N_3080,In_2167,In_2168);
or U3081 (N_3081,In_923,In_74);
nor U3082 (N_3082,In_1320,In_1481);
and U3083 (N_3083,In_72,In_1714);
and U3084 (N_3084,In_459,In_1820);
xnor U3085 (N_3085,In_694,In_21);
nor U3086 (N_3086,In_655,In_2253);
nor U3087 (N_3087,In_87,In_765);
and U3088 (N_3088,In_14,In_2327);
xor U3089 (N_3089,In_2454,In_758);
and U3090 (N_3090,In_2114,In_1311);
xnor U3091 (N_3091,In_244,In_1759);
nand U3092 (N_3092,In_2180,In_486);
nand U3093 (N_3093,In_875,In_1600);
nor U3094 (N_3094,In_2471,In_1979);
xor U3095 (N_3095,In_2222,In_1584);
and U3096 (N_3096,In_2256,In_459);
xnor U3097 (N_3097,In_1890,In_1110);
xor U3098 (N_3098,In_869,In_2456);
xnor U3099 (N_3099,In_764,In_1262);
xnor U3100 (N_3100,In_117,In_725);
or U3101 (N_3101,In_719,In_304);
nor U3102 (N_3102,In_1342,In_1176);
xor U3103 (N_3103,In_1940,In_1899);
xnor U3104 (N_3104,In_1230,In_1282);
and U3105 (N_3105,In_55,In_664);
or U3106 (N_3106,In_190,In_389);
and U3107 (N_3107,In_2029,In_543);
nand U3108 (N_3108,In_792,In_2360);
and U3109 (N_3109,In_1181,In_2267);
nor U3110 (N_3110,In_1506,In_458);
and U3111 (N_3111,In_1323,In_932);
nand U3112 (N_3112,In_729,In_1795);
nand U3113 (N_3113,In_148,In_1476);
nor U3114 (N_3114,In_1314,In_55);
and U3115 (N_3115,In_739,In_20);
nand U3116 (N_3116,In_1122,In_2126);
nor U3117 (N_3117,In_793,In_396);
and U3118 (N_3118,In_1900,In_1240);
xor U3119 (N_3119,In_103,In_1705);
xnor U3120 (N_3120,In_1654,In_2284);
xor U3121 (N_3121,In_130,In_327);
nor U3122 (N_3122,In_42,In_1047);
nand U3123 (N_3123,In_1837,In_2346);
xnor U3124 (N_3124,In_858,In_323);
xor U3125 (N_3125,In_618,In_501);
and U3126 (N_3126,In_1318,In_526);
or U3127 (N_3127,In_227,In_1806);
and U3128 (N_3128,In_2112,In_2323);
nor U3129 (N_3129,In_1582,In_138);
or U3130 (N_3130,In_2076,In_760);
nand U3131 (N_3131,In_1162,In_257);
nand U3132 (N_3132,In_5,In_225);
xnor U3133 (N_3133,In_1553,In_1444);
or U3134 (N_3134,In_1696,In_1164);
and U3135 (N_3135,In_2414,In_163);
nand U3136 (N_3136,In_2389,In_1450);
and U3137 (N_3137,In_1500,In_671);
xnor U3138 (N_3138,In_1421,In_1707);
or U3139 (N_3139,In_40,In_1704);
xor U3140 (N_3140,In_2280,In_1610);
xnor U3141 (N_3141,In_2126,In_250);
xor U3142 (N_3142,In_1197,In_996);
xnor U3143 (N_3143,In_1785,In_1705);
and U3144 (N_3144,In_1019,In_1865);
nand U3145 (N_3145,In_1559,In_2381);
or U3146 (N_3146,In_7,In_1746);
or U3147 (N_3147,In_790,In_843);
nand U3148 (N_3148,In_2210,In_1279);
nor U3149 (N_3149,In_206,In_1255);
nand U3150 (N_3150,In_1725,In_1179);
nor U3151 (N_3151,In_2130,In_167);
or U3152 (N_3152,In_688,In_282);
nor U3153 (N_3153,In_1234,In_1590);
xnor U3154 (N_3154,In_206,In_441);
nor U3155 (N_3155,In_2431,In_1348);
xnor U3156 (N_3156,In_1186,In_1909);
or U3157 (N_3157,In_1172,In_13);
xor U3158 (N_3158,In_227,In_602);
and U3159 (N_3159,In_1752,In_1872);
xnor U3160 (N_3160,In_649,In_896);
or U3161 (N_3161,In_553,In_1648);
or U3162 (N_3162,In_1223,In_594);
nor U3163 (N_3163,In_524,In_432);
and U3164 (N_3164,In_37,In_90);
xnor U3165 (N_3165,In_234,In_1169);
nor U3166 (N_3166,In_111,In_527);
or U3167 (N_3167,In_1725,In_1477);
xnor U3168 (N_3168,In_1917,In_452);
or U3169 (N_3169,In_175,In_1982);
nand U3170 (N_3170,In_2155,In_594);
nand U3171 (N_3171,In_667,In_290);
nand U3172 (N_3172,In_1903,In_329);
nor U3173 (N_3173,In_1166,In_905);
nand U3174 (N_3174,In_1836,In_2201);
xor U3175 (N_3175,In_1680,In_2022);
nand U3176 (N_3176,In_803,In_1618);
xor U3177 (N_3177,In_1443,In_394);
nand U3178 (N_3178,In_1795,In_2460);
xor U3179 (N_3179,In_2267,In_794);
nor U3180 (N_3180,In_436,In_2490);
or U3181 (N_3181,In_1427,In_1582);
xor U3182 (N_3182,In_2120,In_2440);
xnor U3183 (N_3183,In_2199,In_491);
and U3184 (N_3184,In_1645,In_1495);
nor U3185 (N_3185,In_2450,In_1235);
nor U3186 (N_3186,In_1407,In_841);
nand U3187 (N_3187,In_2044,In_1140);
nand U3188 (N_3188,In_1713,In_1223);
or U3189 (N_3189,In_947,In_757);
nor U3190 (N_3190,In_1326,In_414);
or U3191 (N_3191,In_136,In_1345);
and U3192 (N_3192,In_1562,In_51);
or U3193 (N_3193,In_1240,In_757);
nand U3194 (N_3194,In_1778,In_533);
xor U3195 (N_3195,In_2185,In_2014);
nor U3196 (N_3196,In_1706,In_1258);
and U3197 (N_3197,In_2210,In_1412);
or U3198 (N_3198,In_1222,In_1801);
and U3199 (N_3199,In_132,In_2159);
and U3200 (N_3200,In_1272,In_1811);
nor U3201 (N_3201,In_1441,In_1054);
or U3202 (N_3202,In_279,In_2068);
nand U3203 (N_3203,In_765,In_1898);
nand U3204 (N_3204,In_292,In_374);
nor U3205 (N_3205,In_1796,In_947);
or U3206 (N_3206,In_932,In_1506);
xor U3207 (N_3207,In_369,In_2060);
or U3208 (N_3208,In_999,In_569);
and U3209 (N_3209,In_1903,In_544);
nand U3210 (N_3210,In_1393,In_1257);
nor U3211 (N_3211,In_51,In_1579);
xnor U3212 (N_3212,In_432,In_1362);
and U3213 (N_3213,In_2445,In_975);
or U3214 (N_3214,In_1857,In_99);
and U3215 (N_3215,In_1299,In_1748);
or U3216 (N_3216,In_1890,In_2116);
or U3217 (N_3217,In_1114,In_1421);
nand U3218 (N_3218,In_68,In_2046);
xor U3219 (N_3219,In_2280,In_2241);
nor U3220 (N_3220,In_938,In_1815);
nand U3221 (N_3221,In_2272,In_566);
xor U3222 (N_3222,In_1701,In_2031);
nor U3223 (N_3223,In_898,In_1049);
or U3224 (N_3224,In_1145,In_839);
and U3225 (N_3225,In_1028,In_786);
nand U3226 (N_3226,In_1224,In_2385);
nor U3227 (N_3227,In_1597,In_2226);
and U3228 (N_3228,In_602,In_1984);
and U3229 (N_3229,In_529,In_2253);
or U3230 (N_3230,In_2450,In_1805);
and U3231 (N_3231,In_1108,In_1281);
and U3232 (N_3232,In_1790,In_705);
xor U3233 (N_3233,In_1964,In_1225);
and U3234 (N_3234,In_1859,In_965);
or U3235 (N_3235,In_26,In_1777);
and U3236 (N_3236,In_180,In_1413);
nand U3237 (N_3237,In_1345,In_2479);
nor U3238 (N_3238,In_2485,In_1679);
or U3239 (N_3239,In_1690,In_2217);
and U3240 (N_3240,In_1165,In_1526);
xor U3241 (N_3241,In_4,In_1632);
nand U3242 (N_3242,In_2465,In_1186);
and U3243 (N_3243,In_1955,In_303);
nor U3244 (N_3244,In_425,In_1491);
nor U3245 (N_3245,In_758,In_1681);
xnor U3246 (N_3246,In_1544,In_382);
nand U3247 (N_3247,In_867,In_413);
nor U3248 (N_3248,In_54,In_716);
nor U3249 (N_3249,In_761,In_401);
and U3250 (N_3250,In_2309,In_350);
nor U3251 (N_3251,In_1882,In_2251);
nand U3252 (N_3252,In_1877,In_51);
and U3253 (N_3253,In_1329,In_1456);
xor U3254 (N_3254,In_667,In_2180);
xnor U3255 (N_3255,In_1445,In_1803);
xor U3256 (N_3256,In_2118,In_1811);
xor U3257 (N_3257,In_1668,In_1860);
nor U3258 (N_3258,In_1020,In_572);
nand U3259 (N_3259,In_2383,In_1499);
nor U3260 (N_3260,In_1782,In_1483);
nor U3261 (N_3261,In_1948,In_252);
nor U3262 (N_3262,In_2318,In_284);
xnor U3263 (N_3263,In_173,In_957);
nor U3264 (N_3264,In_1576,In_72);
nor U3265 (N_3265,In_595,In_749);
nor U3266 (N_3266,In_1972,In_329);
nand U3267 (N_3267,In_2075,In_1496);
and U3268 (N_3268,In_1455,In_1178);
and U3269 (N_3269,In_1044,In_102);
nand U3270 (N_3270,In_310,In_704);
xnor U3271 (N_3271,In_1206,In_606);
nor U3272 (N_3272,In_1442,In_1798);
nor U3273 (N_3273,In_2253,In_1165);
nand U3274 (N_3274,In_1089,In_1421);
nor U3275 (N_3275,In_1204,In_429);
and U3276 (N_3276,In_2416,In_2053);
or U3277 (N_3277,In_1965,In_1715);
xor U3278 (N_3278,In_89,In_69);
nor U3279 (N_3279,In_1243,In_156);
or U3280 (N_3280,In_243,In_2203);
and U3281 (N_3281,In_42,In_774);
xnor U3282 (N_3282,In_1197,In_407);
nand U3283 (N_3283,In_1294,In_2328);
nand U3284 (N_3284,In_839,In_1574);
xor U3285 (N_3285,In_1379,In_766);
or U3286 (N_3286,In_2276,In_2318);
xnor U3287 (N_3287,In_73,In_1892);
nor U3288 (N_3288,In_1594,In_2156);
or U3289 (N_3289,In_2152,In_557);
nand U3290 (N_3290,In_2389,In_2249);
nor U3291 (N_3291,In_1386,In_646);
nand U3292 (N_3292,In_1570,In_694);
nor U3293 (N_3293,In_2288,In_387);
nor U3294 (N_3294,In_2436,In_2075);
and U3295 (N_3295,In_151,In_213);
nor U3296 (N_3296,In_899,In_979);
xnor U3297 (N_3297,In_65,In_597);
and U3298 (N_3298,In_1987,In_1134);
nor U3299 (N_3299,In_986,In_65);
and U3300 (N_3300,In_590,In_364);
nor U3301 (N_3301,In_1633,In_89);
nor U3302 (N_3302,In_183,In_537);
nor U3303 (N_3303,In_747,In_159);
nand U3304 (N_3304,In_1475,In_896);
and U3305 (N_3305,In_2238,In_335);
and U3306 (N_3306,In_1985,In_465);
or U3307 (N_3307,In_1173,In_226);
nand U3308 (N_3308,In_639,In_42);
nor U3309 (N_3309,In_1321,In_1315);
xnor U3310 (N_3310,In_36,In_571);
xnor U3311 (N_3311,In_2487,In_177);
xnor U3312 (N_3312,In_1651,In_98);
nand U3313 (N_3313,In_1080,In_1651);
nor U3314 (N_3314,In_1863,In_174);
nor U3315 (N_3315,In_699,In_1346);
or U3316 (N_3316,In_2449,In_354);
or U3317 (N_3317,In_750,In_1364);
or U3318 (N_3318,In_1201,In_1964);
or U3319 (N_3319,In_1207,In_1487);
or U3320 (N_3320,In_69,In_23);
nand U3321 (N_3321,In_2019,In_2426);
or U3322 (N_3322,In_1942,In_826);
and U3323 (N_3323,In_1067,In_83);
nand U3324 (N_3324,In_459,In_2406);
nor U3325 (N_3325,In_904,In_501);
or U3326 (N_3326,In_1093,In_1143);
or U3327 (N_3327,In_27,In_1303);
and U3328 (N_3328,In_1955,In_1521);
nor U3329 (N_3329,In_2341,In_1357);
and U3330 (N_3330,In_1396,In_1843);
and U3331 (N_3331,In_1127,In_1952);
and U3332 (N_3332,In_1473,In_2022);
xor U3333 (N_3333,In_2397,In_1462);
xor U3334 (N_3334,In_2157,In_2060);
nand U3335 (N_3335,In_2420,In_2445);
and U3336 (N_3336,In_45,In_240);
nand U3337 (N_3337,In_2378,In_531);
or U3338 (N_3338,In_556,In_1103);
nor U3339 (N_3339,In_922,In_977);
nor U3340 (N_3340,In_1048,In_644);
or U3341 (N_3341,In_1519,In_1401);
xor U3342 (N_3342,In_263,In_366);
nand U3343 (N_3343,In_1713,In_628);
nand U3344 (N_3344,In_2128,In_107);
xor U3345 (N_3345,In_895,In_1821);
and U3346 (N_3346,In_626,In_1938);
and U3347 (N_3347,In_1341,In_1626);
or U3348 (N_3348,In_1832,In_1211);
nor U3349 (N_3349,In_2281,In_442);
and U3350 (N_3350,In_975,In_569);
and U3351 (N_3351,In_1415,In_1118);
xor U3352 (N_3352,In_1590,In_683);
xor U3353 (N_3353,In_2290,In_847);
nor U3354 (N_3354,In_1312,In_1136);
and U3355 (N_3355,In_1402,In_1613);
or U3356 (N_3356,In_300,In_279);
and U3357 (N_3357,In_1430,In_374);
nand U3358 (N_3358,In_688,In_1189);
and U3359 (N_3359,In_139,In_1116);
and U3360 (N_3360,In_830,In_1425);
nand U3361 (N_3361,In_1539,In_486);
nand U3362 (N_3362,In_2108,In_160);
nand U3363 (N_3363,In_867,In_321);
nand U3364 (N_3364,In_984,In_1227);
nand U3365 (N_3365,In_2396,In_909);
xnor U3366 (N_3366,In_1569,In_641);
or U3367 (N_3367,In_2494,In_1182);
xnor U3368 (N_3368,In_1680,In_2330);
nand U3369 (N_3369,In_1985,In_1341);
nand U3370 (N_3370,In_1095,In_2401);
nand U3371 (N_3371,In_1211,In_115);
nor U3372 (N_3372,In_1852,In_167);
nor U3373 (N_3373,In_911,In_985);
or U3374 (N_3374,In_205,In_575);
nor U3375 (N_3375,In_1833,In_428);
xor U3376 (N_3376,In_1746,In_541);
nand U3377 (N_3377,In_2283,In_1965);
and U3378 (N_3378,In_2014,In_412);
xnor U3379 (N_3379,In_2254,In_2000);
and U3380 (N_3380,In_1759,In_929);
nand U3381 (N_3381,In_1770,In_1508);
nor U3382 (N_3382,In_162,In_1966);
xnor U3383 (N_3383,In_282,In_1149);
and U3384 (N_3384,In_61,In_515);
nand U3385 (N_3385,In_1770,In_2063);
xor U3386 (N_3386,In_100,In_1574);
or U3387 (N_3387,In_1693,In_851);
xnor U3388 (N_3388,In_2028,In_2204);
nor U3389 (N_3389,In_46,In_159);
xnor U3390 (N_3390,In_2058,In_2182);
or U3391 (N_3391,In_2361,In_1415);
nand U3392 (N_3392,In_416,In_1378);
xnor U3393 (N_3393,In_2258,In_503);
or U3394 (N_3394,In_638,In_930);
nand U3395 (N_3395,In_764,In_1149);
nand U3396 (N_3396,In_349,In_1506);
nor U3397 (N_3397,In_1227,In_1859);
and U3398 (N_3398,In_2092,In_1761);
or U3399 (N_3399,In_310,In_1337);
or U3400 (N_3400,In_68,In_500);
and U3401 (N_3401,In_2115,In_255);
xnor U3402 (N_3402,In_619,In_1430);
xor U3403 (N_3403,In_674,In_177);
nand U3404 (N_3404,In_1663,In_1273);
or U3405 (N_3405,In_2242,In_1360);
xor U3406 (N_3406,In_174,In_1011);
nor U3407 (N_3407,In_191,In_2420);
and U3408 (N_3408,In_935,In_1441);
or U3409 (N_3409,In_1399,In_1557);
nand U3410 (N_3410,In_821,In_1824);
and U3411 (N_3411,In_800,In_1141);
or U3412 (N_3412,In_1361,In_1647);
nor U3413 (N_3413,In_508,In_2330);
nand U3414 (N_3414,In_560,In_1052);
nor U3415 (N_3415,In_2340,In_313);
xor U3416 (N_3416,In_2223,In_315);
or U3417 (N_3417,In_1544,In_1024);
nand U3418 (N_3418,In_1777,In_1680);
and U3419 (N_3419,In_1586,In_697);
or U3420 (N_3420,In_1757,In_102);
nand U3421 (N_3421,In_2494,In_1559);
nand U3422 (N_3422,In_670,In_1952);
xnor U3423 (N_3423,In_949,In_2379);
and U3424 (N_3424,In_2199,In_111);
nor U3425 (N_3425,In_1657,In_502);
xor U3426 (N_3426,In_2165,In_1351);
or U3427 (N_3427,In_1738,In_1444);
and U3428 (N_3428,In_442,In_316);
nor U3429 (N_3429,In_89,In_180);
nor U3430 (N_3430,In_1485,In_1680);
nor U3431 (N_3431,In_455,In_1626);
xor U3432 (N_3432,In_1068,In_384);
xnor U3433 (N_3433,In_497,In_1708);
nor U3434 (N_3434,In_598,In_736);
nand U3435 (N_3435,In_1738,In_2419);
nand U3436 (N_3436,In_162,In_444);
xnor U3437 (N_3437,In_733,In_2300);
nand U3438 (N_3438,In_710,In_960);
or U3439 (N_3439,In_955,In_1824);
or U3440 (N_3440,In_1999,In_1607);
or U3441 (N_3441,In_1873,In_1633);
nor U3442 (N_3442,In_963,In_2352);
or U3443 (N_3443,In_2152,In_1992);
xnor U3444 (N_3444,In_1368,In_2364);
xor U3445 (N_3445,In_2167,In_1007);
xor U3446 (N_3446,In_182,In_2184);
or U3447 (N_3447,In_774,In_1424);
xor U3448 (N_3448,In_2185,In_535);
or U3449 (N_3449,In_2317,In_1543);
and U3450 (N_3450,In_484,In_2357);
xor U3451 (N_3451,In_78,In_905);
xnor U3452 (N_3452,In_1649,In_1738);
and U3453 (N_3453,In_1506,In_1750);
and U3454 (N_3454,In_1558,In_304);
xnor U3455 (N_3455,In_301,In_27);
xor U3456 (N_3456,In_861,In_1728);
or U3457 (N_3457,In_1966,In_726);
and U3458 (N_3458,In_1866,In_1686);
or U3459 (N_3459,In_2173,In_2478);
and U3460 (N_3460,In_548,In_560);
xor U3461 (N_3461,In_533,In_228);
or U3462 (N_3462,In_789,In_451);
xor U3463 (N_3463,In_2079,In_1656);
xnor U3464 (N_3464,In_66,In_1481);
xnor U3465 (N_3465,In_2487,In_354);
and U3466 (N_3466,In_649,In_1422);
nor U3467 (N_3467,In_177,In_1347);
nor U3468 (N_3468,In_758,In_2130);
and U3469 (N_3469,In_1778,In_1442);
nor U3470 (N_3470,In_1,In_1341);
nand U3471 (N_3471,In_169,In_1978);
nand U3472 (N_3472,In_1760,In_169);
nor U3473 (N_3473,In_2203,In_719);
and U3474 (N_3474,In_1536,In_831);
and U3475 (N_3475,In_1303,In_155);
xnor U3476 (N_3476,In_652,In_2314);
and U3477 (N_3477,In_2086,In_1468);
or U3478 (N_3478,In_24,In_1358);
or U3479 (N_3479,In_671,In_709);
nor U3480 (N_3480,In_885,In_1796);
xor U3481 (N_3481,In_2096,In_31);
and U3482 (N_3482,In_1738,In_1579);
nor U3483 (N_3483,In_1737,In_462);
or U3484 (N_3484,In_876,In_120);
xnor U3485 (N_3485,In_842,In_937);
nand U3486 (N_3486,In_121,In_66);
or U3487 (N_3487,In_2302,In_666);
nand U3488 (N_3488,In_417,In_1547);
and U3489 (N_3489,In_1488,In_736);
nor U3490 (N_3490,In_2431,In_2211);
or U3491 (N_3491,In_833,In_2434);
xnor U3492 (N_3492,In_1641,In_874);
nand U3493 (N_3493,In_30,In_1540);
nor U3494 (N_3494,In_1948,In_1472);
or U3495 (N_3495,In_1844,In_1930);
nor U3496 (N_3496,In_1230,In_165);
and U3497 (N_3497,In_341,In_1884);
xor U3498 (N_3498,In_221,In_1045);
nor U3499 (N_3499,In_298,In_906);
nand U3500 (N_3500,In_1881,In_1613);
xnor U3501 (N_3501,In_705,In_643);
xor U3502 (N_3502,In_1436,In_404);
or U3503 (N_3503,In_566,In_2216);
nand U3504 (N_3504,In_904,In_81);
and U3505 (N_3505,In_3,In_354);
nor U3506 (N_3506,In_823,In_1441);
or U3507 (N_3507,In_764,In_436);
nand U3508 (N_3508,In_1779,In_281);
or U3509 (N_3509,In_2208,In_261);
xnor U3510 (N_3510,In_1373,In_847);
or U3511 (N_3511,In_1599,In_2456);
nand U3512 (N_3512,In_2450,In_1309);
nor U3513 (N_3513,In_303,In_2080);
or U3514 (N_3514,In_2250,In_2295);
and U3515 (N_3515,In_1830,In_70);
or U3516 (N_3516,In_664,In_1971);
xnor U3517 (N_3517,In_1312,In_867);
or U3518 (N_3518,In_885,In_713);
nor U3519 (N_3519,In_779,In_1411);
nand U3520 (N_3520,In_218,In_268);
xor U3521 (N_3521,In_1381,In_88);
nor U3522 (N_3522,In_699,In_605);
and U3523 (N_3523,In_2334,In_604);
and U3524 (N_3524,In_1792,In_142);
nand U3525 (N_3525,In_1805,In_1392);
or U3526 (N_3526,In_2390,In_1298);
xnor U3527 (N_3527,In_516,In_778);
or U3528 (N_3528,In_661,In_338);
nor U3529 (N_3529,In_189,In_528);
and U3530 (N_3530,In_587,In_358);
xnor U3531 (N_3531,In_1529,In_2366);
nand U3532 (N_3532,In_880,In_2408);
and U3533 (N_3533,In_961,In_1418);
or U3534 (N_3534,In_1822,In_826);
or U3535 (N_3535,In_1983,In_2134);
or U3536 (N_3536,In_972,In_1141);
nor U3537 (N_3537,In_1288,In_1258);
nand U3538 (N_3538,In_2347,In_399);
and U3539 (N_3539,In_1902,In_2456);
xor U3540 (N_3540,In_153,In_1179);
nand U3541 (N_3541,In_1718,In_481);
and U3542 (N_3542,In_802,In_2212);
or U3543 (N_3543,In_130,In_2005);
nor U3544 (N_3544,In_789,In_1078);
nor U3545 (N_3545,In_1150,In_799);
or U3546 (N_3546,In_1383,In_257);
nand U3547 (N_3547,In_1791,In_15);
nor U3548 (N_3548,In_51,In_1798);
xnor U3549 (N_3549,In_1798,In_115);
nor U3550 (N_3550,In_2106,In_1596);
and U3551 (N_3551,In_1415,In_615);
or U3552 (N_3552,In_517,In_134);
nor U3553 (N_3553,In_1480,In_1363);
nor U3554 (N_3554,In_972,In_372);
and U3555 (N_3555,In_1216,In_1725);
nand U3556 (N_3556,In_1811,In_1589);
nor U3557 (N_3557,In_1632,In_2438);
xnor U3558 (N_3558,In_1,In_1034);
xor U3559 (N_3559,In_630,In_2262);
and U3560 (N_3560,In_1846,In_2015);
nor U3561 (N_3561,In_2344,In_479);
nor U3562 (N_3562,In_1374,In_2266);
nor U3563 (N_3563,In_1520,In_239);
or U3564 (N_3564,In_876,In_758);
nand U3565 (N_3565,In_1786,In_1550);
xnor U3566 (N_3566,In_797,In_1822);
and U3567 (N_3567,In_377,In_2341);
and U3568 (N_3568,In_857,In_1752);
and U3569 (N_3569,In_623,In_1831);
or U3570 (N_3570,In_2053,In_1892);
xor U3571 (N_3571,In_46,In_7);
xnor U3572 (N_3572,In_763,In_1154);
nand U3573 (N_3573,In_1819,In_137);
xnor U3574 (N_3574,In_364,In_859);
nor U3575 (N_3575,In_153,In_48);
nor U3576 (N_3576,In_1751,In_632);
and U3577 (N_3577,In_1914,In_984);
and U3578 (N_3578,In_2485,In_476);
or U3579 (N_3579,In_529,In_615);
xnor U3580 (N_3580,In_1358,In_49);
nor U3581 (N_3581,In_286,In_912);
and U3582 (N_3582,In_1278,In_1516);
xnor U3583 (N_3583,In_854,In_1568);
and U3584 (N_3584,In_1239,In_1476);
or U3585 (N_3585,In_2440,In_1652);
nor U3586 (N_3586,In_433,In_1063);
and U3587 (N_3587,In_1819,In_1718);
nand U3588 (N_3588,In_1071,In_331);
or U3589 (N_3589,In_745,In_11);
or U3590 (N_3590,In_2189,In_1437);
nand U3591 (N_3591,In_1391,In_1266);
and U3592 (N_3592,In_1342,In_2428);
nor U3593 (N_3593,In_1228,In_1446);
xnor U3594 (N_3594,In_2333,In_2196);
nor U3595 (N_3595,In_218,In_878);
nand U3596 (N_3596,In_1153,In_500);
xor U3597 (N_3597,In_841,In_1456);
nor U3598 (N_3598,In_1369,In_2179);
xor U3599 (N_3599,In_16,In_1227);
nand U3600 (N_3600,In_1192,In_2178);
xor U3601 (N_3601,In_1734,In_1398);
nor U3602 (N_3602,In_640,In_76);
and U3603 (N_3603,In_386,In_2352);
nand U3604 (N_3604,In_2279,In_15);
or U3605 (N_3605,In_2452,In_594);
nand U3606 (N_3606,In_934,In_2334);
or U3607 (N_3607,In_798,In_557);
xor U3608 (N_3608,In_2385,In_470);
nor U3609 (N_3609,In_2431,In_1417);
xor U3610 (N_3610,In_1726,In_1459);
nand U3611 (N_3611,In_540,In_121);
and U3612 (N_3612,In_337,In_1093);
nand U3613 (N_3613,In_654,In_292);
xnor U3614 (N_3614,In_1876,In_352);
or U3615 (N_3615,In_2161,In_2155);
nor U3616 (N_3616,In_933,In_331);
or U3617 (N_3617,In_2072,In_2056);
nand U3618 (N_3618,In_2314,In_491);
and U3619 (N_3619,In_188,In_782);
nand U3620 (N_3620,In_2108,In_42);
or U3621 (N_3621,In_1470,In_1572);
nor U3622 (N_3622,In_1963,In_1997);
nor U3623 (N_3623,In_1224,In_2345);
xor U3624 (N_3624,In_1119,In_406);
or U3625 (N_3625,In_1852,In_694);
and U3626 (N_3626,In_529,In_1354);
nor U3627 (N_3627,In_1333,In_1851);
nand U3628 (N_3628,In_1797,In_145);
and U3629 (N_3629,In_1392,In_1122);
xor U3630 (N_3630,In_893,In_130);
xnor U3631 (N_3631,In_2152,In_268);
nor U3632 (N_3632,In_2185,In_1829);
nor U3633 (N_3633,In_955,In_428);
xor U3634 (N_3634,In_2138,In_1578);
nor U3635 (N_3635,In_976,In_638);
xnor U3636 (N_3636,In_2023,In_194);
nor U3637 (N_3637,In_1143,In_434);
nand U3638 (N_3638,In_791,In_905);
nand U3639 (N_3639,In_1350,In_1763);
xor U3640 (N_3640,In_2311,In_1275);
nor U3641 (N_3641,In_1241,In_680);
nand U3642 (N_3642,In_1610,In_309);
nor U3643 (N_3643,In_113,In_238);
or U3644 (N_3644,In_1025,In_1926);
and U3645 (N_3645,In_1260,In_2002);
nand U3646 (N_3646,In_748,In_1040);
xor U3647 (N_3647,In_872,In_1263);
or U3648 (N_3648,In_2078,In_136);
and U3649 (N_3649,In_270,In_317);
nand U3650 (N_3650,In_188,In_1185);
or U3651 (N_3651,In_2279,In_54);
and U3652 (N_3652,In_1037,In_1854);
or U3653 (N_3653,In_929,In_144);
and U3654 (N_3654,In_2107,In_1193);
nor U3655 (N_3655,In_1019,In_24);
xnor U3656 (N_3656,In_1866,In_61);
or U3657 (N_3657,In_873,In_670);
and U3658 (N_3658,In_706,In_2112);
and U3659 (N_3659,In_1555,In_719);
nand U3660 (N_3660,In_1184,In_875);
nand U3661 (N_3661,In_220,In_411);
or U3662 (N_3662,In_456,In_1786);
or U3663 (N_3663,In_2342,In_250);
nand U3664 (N_3664,In_91,In_535);
or U3665 (N_3665,In_295,In_2396);
xnor U3666 (N_3666,In_614,In_1535);
or U3667 (N_3667,In_1428,In_1511);
or U3668 (N_3668,In_2263,In_1337);
nand U3669 (N_3669,In_157,In_2054);
xnor U3670 (N_3670,In_886,In_676);
nor U3671 (N_3671,In_1736,In_1174);
or U3672 (N_3672,In_2082,In_1581);
nor U3673 (N_3673,In_1350,In_2291);
nand U3674 (N_3674,In_1897,In_2279);
and U3675 (N_3675,In_1657,In_31);
xnor U3676 (N_3676,In_198,In_2125);
nor U3677 (N_3677,In_648,In_831);
and U3678 (N_3678,In_465,In_1430);
xnor U3679 (N_3679,In_2018,In_1076);
nor U3680 (N_3680,In_1107,In_1101);
and U3681 (N_3681,In_841,In_332);
nand U3682 (N_3682,In_512,In_1624);
nor U3683 (N_3683,In_137,In_1240);
nor U3684 (N_3684,In_1367,In_2209);
or U3685 (N_3685,In_1403,In_2279);
xnor U3686 (N_3686,In_76,In_2348);
nor U3687 (N_3687,In_95,In_1851);
xor U3688 (N_3688,In_1919,In_1199);
or U3689 (N_3689,In_1582,In_581);
or U3690 (N_3690,In_678,In_232);
and U3691 (N_3691,In_561,In_2379);
and U3692 (N_3692,In_2483,In_58);
and U3693 (N_3693,In_381,In_2000);
xnor U3694 (N_3694,In_1831,In_401);
nor U3695 (N_3695,In_1371,In_2154);
nand U3696 (N_3696,In_22,In_1298);
or U3697 (N_3697,In_472,In_2416);
xor U3698 (N_3698,In_709,In_1919);
nand U3699 (N_3699,In_2495,In_2233);
and U3700 (N_3700,In_894,In_1072);
nand U3701 (N_3701,In_102,In_1876);
nor U3702 (N_3702,In_2035,In_521);
xnor U3703 (N_3703,In_2251,In_1116);
and U3704 (N_3704,In_1222,In_1941);
or U3705 (N_3705,In_1859,In_1344);
and U3706 (N_3706,In_1923,In_291);
nor U3707 (N_3707,In_173,In_1581);
and U3708 (N_3708,In_1903,In_1932);
xor U3709 (N_3709,In_1390,In_1076);
or U3710 (N_3710,In_951,In_400);
nand U3711 (N_3711,In_678,In_2099);
xnor U3712 (N_3712,In_78,In_1176);
nand U3713 (N_3713,In_2031,In_798);
or U3714 (N_3714,In_1536,In_1532);
and U3715 (N_3715,In_505,In_1802);
and U3716 (N_3716,In_1765,In_2141);
nor U3717 (N_3717,In_761,In_2338);
and U3718 (N_3718,In_1706,In_2379);
and U3719 (N_3719,In_558,In_2447);
xnor U3720 (N_3720,In_41,In_1109);
xor U3721 (N_3721,In_933,In_381);
nor U3722 (N_3722,In_1370,In_2032);
nand U3723 (N_3723,In_434,In_1547);
nor U3724 (N_3724,In_2473,In_2399);
and U3725 (N_3725,In_1763,In_821);
xor U3726 (N_3726,In_1868,In_2118);
nor U3727 (N_3727,In_2441,In_1811);
nor U3728 (N_3728,In_1702,In_337);
and U3729 (N_3729,In_483,In_284);
nor U3730 (N_3730,In_803,In_2320);
nor U3731 (N_3731,In_1857,In_1855);
xor U3732 (N_3732,In_550,In_2372);
nor U3733 (N_3733,In_113,In_1036);
xnor U3734 (N_3734,In_770,In_1012);
nor U3735 (N_3735,In_85,In_1179);
nor U3736 (N_3736,In_299,In_557);
nor U3737 (N_3737,In_253,In_404);
nand U3738 (N_3738,In_751,In_1139);
and U3739 (N_3739,In_714,In_2323);
nor U3740 (N_3740,In_1090,In_992);
or U3741 (N_3741,In_2488,In_1192);
nor U3742 (N_3742,In_1673,In_1648);
or U3743 (N_3743,In_1821,In_1331);
or U3744 (N_3744,In_913,In_1701);
nand U3745 (N_3745,In_404,In_2431);
xnor U3746 (N_3746,In_2090,In_2486);
xor U3747 (N_3747,In_1026,In_960);
or U3748 (N_3748,In_1901,In_1808);
nand U3749 (N_3749,In_1208,In_1346);
and U3750 (N_3750,In_568,In_1170);
and U3751 (N_3751,In_1743,In_982);
nor U3752 (N_3752,In_590,In_1607);
and U3753 (N_3753,In_1143,In_193);
nand U3754 (N_3754,In_1088,In_1848);
nor U3755 (N_3755,In_1467,In_737);
nor U3756 (N_3756,In_225,In_1731);
and U3757 (N_3757,In_667,In_320);
and U3758 (N_3758,In_2416,In_1462);
nand U3759 (N_3759,In_297,In_1655);
nor U3760 (N_3760,In_1439,In_209);
or U3761 (N_3761,In_1742,In_1491);
xnor U3762 (N_3762,In_1652,In_856);
or U3763 (N_3763,In_1246,In_2108);
xor U3764 (N_3764,In_1911,In_517);
nor U3765 (N_3765,In_2254,In_831);
and U3766 (N_3766,In_419,In_2014);
xor U3767 (N_3767,In_590,In_1561);
or U3768 (N_3768,In_1176,In_36);
xor U3769 (N_3769,In_1421,In_985);
nor U3770 (N_3770,In_1818,In_2157);
nand U3771 (N_3771,In_1820,In_2299);
nand U3772 (N_3772,In_66,In_2372);
nor U3773 (N_3773,In_1397,In_59);
xor U3774 (N_3774,In_1137,In_275);
nand U3775 (N_3775,In_1348,In_1954);
nand U3776 (N_3776,In_318,In_1511);
nand U3777 (N_3777,In_423,In_262);
nand U3778 (N_3778,In_269,In_1090);
or U3779 (N_3779,In_2439,In_519);
nor U3780 (N_3780,In_2451,In_480);
and U3781 (N_3781,In_818,In_1552);
xor U3782 (N_3782,In_1599,In_1539);
nand U3783 (N_3783,In_475,In_1221);
or U3784 (N_3784,In_1226,In_1756);
nand U3785 (N_3785,In_2304,In_2300);
or U3786 (N_3786,In_726,In_2476);
nand U3787 (N_3787,In_2210,In_1923);
or U3788 (N_3788,In_1411,In_93);
nor U3789 (N_3789,In_996,In_2330);
xor U3790 (N_3790,In_1352,In_1440);
and U3791 (N_3791,In_514,In_44);
and U3792 (N_3792,In_727,In_2257);
xnor U3793 (N_3793,In_1777,In_1204);
nor U3794 (N_3794,In_209,In_1389);
nand U3795 (N_3795,In_2355,In_1056);
and U3796 (N_3796,In_1136,In_2114);
nor U3797 (N_3797,In_156,In_1294);
and U3798 (N_3798,In_1220,In_1219);
nand U3799 (N_3799,In_1978,In_998);
or U3800 (N_3800,In_1066,In_642);
nor U3801 (N_3801,In_1786,In_1490);
nand U3802 (N_3802,In_2244,In_1573);
nor U3803 (N_3803,In_568,In_1050);
or U3804 (N_3804,In_1735,In_2490);
nand U3805 (N_3805,In_766,In_1381);
and U3806 (N_3806,In_1948,In_571);
nor U3807 (N_3807,In_2373,In_1593);
nor U3808 (N_3808,In_122,In_963);
and U3809 (N_3809,In_1886,In_1654);
xnor U3810 (N_3810,In_1372,In_1717);
nand U3811 (N_3811,In_351,In_2403);
nand U3812 (N_3812,In_2393,In_529);
xnor U3813 (N_3813,In_1104,In_2023);
and U3814 (N_3814,In_22,In_411);
nand U3815 (N_3815,In_760,In_1784);
nor U3816 (N_3816,In_237,In_1417);
nor U3817 (N_3817,In_167,In_427);
nor U3818 (N_3818,In_1789,In_798);
nor U3819 (N_3819,In_479,In_947);
nor U3820 (N_3820,In_61,In_2371);
and U3821 (N_3821,In_1683,In_682);
nand U3822 (N_3822,In_1020,In_2205);
or U3823 (N_3823,In_410,In_189);
nand U3824 (N_3824,In_2425,In_164);
xnor U3825 (N_3825,In_818,In_205);
xnor U3826 (N_3826,In_2425,In_1302);
and U3827 (N_3827,In_1902,In_365);
nand U3828 (N_3828,In_446,In_247);
nand U3829 (N_3829,In_2125,In_1166);
xnor U3830 (N_3830,In_1001,In_1687);
nand U3831 (N_3831,In_2338,In_234);
nor U3832 (N_3832,In_1317,In_2267);
nand U3833 (N_3833,In_2490,In_164);
nor U3834 (N_3834,In_1935,In_1630);
or U3835 (N_3835,In_327,In_1997);
and U3836 (N_3836,In_2339,In_17);
nor U3837 (N_3837,In_1130,In_1445);
xor U3838 (N_3838,In_643,In_409);
or U3839 (N_3839,In_1877,In_507);
or U3840 (N_3840,In_1428,In_767);
xor U3841 (N_3841,In_1898,In_1804);
nor U3842 (N_3842,In_436,In_1402);
nand U3843 (N_3843,In_844,In_2191);
and U3844 (N_3844,In_994,In_919);
and U3845 (N_3845,In_1594,In_2418);
and U3846 (N_3846,In_2167,In_1999);
nand U3847 (N_3847,In_1694,In_2140);
nor U3848 (N_3848,In_1789,In_2356);
and U3849 (N_3849,In_469,In_939);
or U3850 (N_3850,In_922,In_2298);
or U3851 (N_3851,In_2337,In_1691);
nor U3852 (N_3852,In_2032,In_245);
and U3853 (N_3853,In_1838,In_2075);
xnor U3854 (N_3854,In_2162,In_1522);
nand U3855 (N_3855,In_1108,In_168);
nand U3856 (N_3856,In_1001,In_437);
or U3857 (N_3857,In_234,In_977);
or U3858 (N_3858,In_221,In_820);
or U3859 (N_3859,In_241,In_29);
xnor U3860 (N_3860,In_1938,In_420);
xor U3861 (N_3861,In_1670,In_247);
and U3862 (N_3862,In_2230,In_2027);
xnor U3863 (N_3863,In_1646,In_189);
and U3864 (N_3864,In_328,In_1060);
and U3865 (N_3865,In_1193,In_1369);
nand U3866 (N_3866,In_589,In_1933);
nor U3867 (N_3867,In_65,In_553);
nor U3868 (N_3868,In_782,In_819);
nor U3869 (N_3869,In_1502,In_1071);
nor U3870 (N_3870,In_923,In_199);
xor U3871 (N_3871,In_2230,In_1647);
nor U3872 (N_3872,In_416,In_520);
nor U3873 (N_3873,In_16,In_1998);
nor U3874 (N_3874,In_1889,In_1203);
nor U3875 (N_3875,In_2192,In_1357);
nand U3876 (N_3876,In_1970,In_1407);
nor U3877 (N_3877,In_1881,In_81);
nand U3878 (N_3878,In_1181,In_1414);
or U3879 (N_3879,In_313,In_1132);
nor U3880 (N_3880,In_1318,In_1596);
nand U3881 (N_3881,In_1515,In_2156);
or U3882 (N_3882,In_1814,In_1049);
and U3883 (N_3883,In_670,In_1832);
nand U3884 (N_3884,In_171,In_1056);
nor U3885 (N_3885,In_2356,In_1230);
nand U3886 (N_3886,In_444,In_202);
xor U3887 (N_3887,In_621,In_1255);
nor U3888 (N_3888,In_314,In_2413);
nand U3889 (N_3889,In_2324,In_243);
nand U3890 (N_3890,In_1781,In_1927);
and U3891 (N_3891,In_2167,In_345);
and U3892 (N_3892,In_1656,In_1272);
and U3893 (N_3893,In_2220,In_2029);
xnor U3894 (N_3894,In_1588,In_1899);
or U3895 (N_3895,In_1254,In_1740);
or U3896 (N_3896,In_1025,In_88);
xor U3897 (N_3897,In_2459,In_1290);
and U3898 (N_3898,In_2282,In_2168);
or U3899 (N_3899,In_676,In_1672);
nand U3900 (N_3900,In_2244,In_2158);
and U3901 (N_3901,In_2289,In_1520);
nand U3902 (N_3902,In_1198,In_884);
nand U3903 (N_3903,In_665,In_1759);
or U3904 (N_3904,In_1035,In_482);
or U3905 (N_3905,In_1795,In_2302);
or U3906 (N_3906,In_2136,In_790);
nand U3907 (N_3907,In_35,In_1897);
nor U3908 (N_3908,In_1977,In_2189);
xor U3909 (N_3909,In_1559,In_2281);
and U3910 (N_3910,In_2260,In_487);
xor U3911 (N_3911,In_0,In_2399);
or U3912 (N_3912,In_949,In_1820);
or U3913 (N_3913,In_533,In_915);
nor U3914 (N_3914,In_306,In_421);
xnor U3915 (N_3915,In_39,In_980);
and U3916 (N_3916,In_527,In_833);
nand U3917 (N_3917,In_530,In_1103);
nand U3918 (N_3918,In_2472,In_1554);
or U3919 (N_3919,In_1813,In_1839);
nand U3920 (N_3920,In_707,In_827);
nand U3921 (N_3921,In_612,In_1775);
nand U3922 (N_3922,In_1108,In_887);
nand U3923 (N_3923,In_1959,In_545);
xor U3924 (N_3924,In_2461,In_824);
nor U3925 (N_3925,In_1132,In_1418);
xnor U3926 (N_3926,In_1683,In_1473);
or U3927 (N_3927,In_756,In_1814);
and U3928 (N_3928,In_1401,In_1104);
and U3929 (N_3929,In_2320,In_457);
xnor U3930 (N_3930,In_931,In_1516);
nor U3931 (N_3931,In_19,In_2463);
or U3932 (N_3932,In_2443,In_663);
nor U3933 (N_3933,In_1758,In_1344);
nor U3934 (N_3934,In_2043,In_1487);
nor U3935 (N_3935,In_933,In_788);
xor U3936 (N_3936,In_909,In_1442);
nand U3937 (N_3937,In_1451,In_381);
xor U3938 (N_3938,In_1571,In_2366);
and U3939 (N_3939,In_151,In_1768);
nand U3940 (N_3940,In_710,In_2455);
xnor U3941 (N_3941,In_27,In_2137);
xnor U3942 (N_3942,In_2177,In_1240);
or U3943 (N_3943,In_1392,In_1087);
xnor U3944 (N_3944,In_302,In_650);
nor U3945 (N_3945,In_2352,In_267);
xor U3946 (N_3946,In_1487,In_1050);
or U3947 (N_3947,In_2155,In_9);
and U3948 (N_3948,In_2171,In_1623);
xor U3949 (N_3949,In_648,In_1749);
and U3950 (N_3950,In_1823,In_325);
and U3951 (N_3951,In_2275,In_824);
or U3952 (N_3952,In_2145,In_489);
and U3953 (N_3953,In_1061,In_1242);
nor U3954 (N_3954,In_272,In_746);
and U3955 (N_3955,In_1639,In_2199);
and U3956 (N_3956,In_1409,In_525);
nand U3957 (N_3957,In_1325,In_2487);
nand U3958 (N_3958,In_2373,In_1475);
or U3959 (N_3959,In_1231,In_1250);
and U3960 (N_3960,In_221,In_1400);
nand U3961 (N_3961,In_1545,In_1759);
xor U3962 (N_3962,In_1615,In_1342);
and U3963 (N_3963,In_712,In_2411);
or U3964 (N_3964,In_2057,In_934);
or U3965 (N_3965,In_901,In_51);
nand U3966 (N_3966,In_497,In_1113);
or U3967 (N_3967,In_1676,In_2446);
xor U3968 (N_3968,In_1451,In_1774);
nand U3969 (N_3969,In_99,In_877);
and U3970 (N_3970,In_365,In_544);
or U3971 (N_3971,In_2224,In_275);
or U3972 (N_3972,In_1959,In_337);
xor U3973 (N_3973,In_2106,In_1520);
nand U3974 (N_3974,In_738,In_511);
nand U3975 (N_3975,In_984,In_2404);
nand U3976 (N_3976,In_2319,In_1443);
nand U3977 (N_3977,In_611,In_393);
nor U3978 (N_3978,In_2085,In_2437);
nand U3979 (N_3979,In_1735,In_1617);
and U3980 (N_3980,In_1300,In_1396);
and U3981 (N_3981,In_340,In_72);
nor U3982 (N_3982,In_1156,In_909);
nor U3983 (N_3983,In_468,In_366);
or U3984 (N_3984,In_503,In_183);
and U3985 (N_3985,In_174,In_1521);
and U3986 (N_3986,In_1781,In_1913);
and U3987 (N_3987,In_199,In_1161);
xnor U3988 (N_3988,In_1597,In_1993);
and U3989 (N_3989,In_1461,In_2015);
or U3990 (N_3990,In_1044,In_193);
nand U3991 (N_3991,In_2067,In_42);
xor U3992 (N_3992,In_2472,In_210);
xnor U3993 (N_3993,In_599,In_1283);
xor U3994 (N_3994,In_1633,In_65);
nand U3995 (N_3995,In_553,In_2204);
and U3996 (N_3996,In_572,In_183);
or U3997 (N_3997,In_2070,In_2327);
xnor U3998 (N_3998,In_256,In_313);
nor U3999 (N_3999,In_677,In_1219);
nand U4000 (N_4000,In_1078,In_629);
xnor U4001 (N_4001,In_1362,In_478);
xor U4002 (N_4002,In_122,In_1948);
xor U4003 (N_4003,In_2326,In_462);
xor U4004 (N_4004,In_378,In_634);
and U4005 (N_4005,In_1145,In_362);
and U4006 (N_4006,In_1133,In_354);
and U4007 (N_4007,In_2170,In_434);
or U4008 (N_4008,In_1028,In_90);
nand U4009 (N_4009,In_552,In_2187);
nand U4010 (N_4010,In_2439,In_2334);
xor U4011 (N_4011,In_413,In_663);
or U4012 (N_4012,In_1175,In_1354);
nor U4013 (N_4013,In_1432,In_654);
xnor U4014 (N_4014,In_1222,In_2124);
nor U4015 (N_4015,In_171,In_454);
or U4016 (N_4016,In_1329,In_264);
or U4017 (N_4017,In_947,In_94);
nor U4018 (N_4018,In_1588,In_2133);
xnor U4019 (N_4019,In_422,In_1010);
xor U4020 (N_4020,In_1105,In_278);
and U4021 (N_4021,In_320,In_2068);
and U4022 (N_4022,In_472,In_1289);
nor U4023 (N_4023,In_1860,In_2163);
nor U4024 (N_4024,In_2136,In_105);
xnor U4025 (N_4025,In_213,In_920);
or U4026 (N_4026,In_1011,In_1672);
xor U4027 (N_4027,In_909,In_2251);
xnor U4028 (N_4028,In_2427,In_1990);
or U4029 (N_4029,In_1283,In_1930);
nor U4030 (N_4030,In_1665,In_1530);
or U4031 (N_4031,In_206,In_178);
nand U4032 (N_4032,In_409,In_827);
and U4033 (N_4033,In_2381,In_1497);
nor U4034 (N_4034,In_313,In_69);
nand U4035 (N_4035,In_1838,In_1711);
nand U4036 (N_4036,In_2499,In_2283);
nor U4037 (N_4037,In_506,In_576);
nor U4038 (N_4038,In_498,In_224);
and U4039 (N_4039,In_158,In_343);
nor U4040 (N_4040,In_2427,In_1763);
nand U4041 (N_4041,In_764,In_2303);
and U4042 (N_4042,In_412,In_1908);
nand U4043 (N_4043,In_1848,In_1272);
nor U4044 (N_4044,In_313,In_561);
or U4045 (N_4045,In_1227,In_229);
xnor U4046 (N_4046,In_2190,In_847);
nand U4047 (N_4047,In_1821,In_2394);
xor U4048 (N_4048,In_254,In_1240);
nor U4049 (N_4049,In_1772,In_948);
or U4050 (N_4050,In_1536,In_1744);
or U4051 (N_4051,In_1131,In_2186);
xor U4052 (N_4052,In_1733,In_2076);
xor U4053 (N_4053,In_400,In_1145);
or U4054 (N_4054,In_2081,In_1461);
or U4055 (N_4055,In_969,In_2304);
nand U4056 (N_4056,In_1149,In_329);
xnor U4057 (N_4057,In_1855,In_1695);
nand U4058 (N_4058,In_908,In_1094);
and U4059 (N_4059,In_1159,In_364);
nand U4060 (N_4060,In_719,In_1232);
nor U4061 (N_4061,In_1568,In_1235);
nand U4062 (N_4062,In_413,In_130);
nand U4063 (N_4063,In_86,In_2425);
xor U4064 (N_4064,In_2275,In_548);
or U4065 (N_4065,In_1762,In_2235);
or U4066 (N_4066,In_1285,In_570);
nor U4067 (N_4067,In_2202,In_1922);
nand U4068 (N_4068,In_1825,In_2113);
or U4069 (N_4069,In_950,In_859);
or U4070 (N_4070,In_1471,In_1864);
or U4071 (N_4071,In_1581,In_1857);
nor U4072 (N_4072,In_2121,In_1590);
nand U4073 (N_4073,In_1342,In_1046);
nor U4074 (N_4074,In_653,In_1881);
and U4075 (N_4075,In_137,In_1670);
or U4076 (N_4076,In_351,In_299);
nor U4077 (N_4077,In_1837,In_975);
xnor U4078 (N_4078,In_2212,In_573);
or U4079 (N_4079,In_2466,In_1593);
and U4080 (N_4080,In_2025,In_2458);
and U4081 (N_4081,In_37,In_1295);
nand U4082 (N_4082,In_1337,In_2003);
nor U4083 (N_4083,In_2200,In_1371);
and U4084 (N_4084,In_1249,In_802);
or U4085 (N_4085,In_324,In_1683);
nor U4086 (N_4086,In_2213,In_2335);
nand U4087 (N_4087,In_1074,In_1398);
nand U4088 (N_4088,In_953,In_2037);
or U4089 (N_4089,In_845,In_849);
and U4090 (N_4090,In_296,In_83);
nor U4091 (N_4091,In_1496,In_2152);
xnor U4092 (N_4092,In_374,In_385);
nand U4093 (N_4093,In_2133,In_710);
nand U4094 (N_4094,In_1808,In_948);
or U4095 (N_4095,In_2161,In_36);
xnor U4096 (N_4096,In_355,In_246);
xor U4097 (N_4097,In_1709,In_2143);
nor U4098 (N_4098,In_2154,In_1714);
nor U4099 (N_4099,In_980,In_2310);
and U4100 (N_4100,In_1467,In_2283);
xor U4101 (N_4101,In_605,In_2449);
xor U4102 (N_4102,In_2021,In_1411);
or U4103 (N_4103,In_1041,In_2157);
nor U4104 (N_4104,In_1808,In_2041);
and U4105 (N_4105,In_2196,In_912);
xnor U4106 (N_4106,In_816,In_1025);
or U4107 (N_4107,In_409,In_2181);
nor U4108 (N_4108,In_2042,In_1367);
xnor U4109 (N_4109,In_293,In_1296);
or U4110 (N_4110,In_2196,In_2453);
xor U4111 (N_4111,In_2186,In_741);
and U4112 (N_4112,In_1161,In_1284);
or U4113 (N_4113,In_286,In_744);
xor U4114 (N_4114,In_2068,In_885);
or U4115 (N_4115,In_1946,In_1328);
xor U4116 (N_4116,In_1491,In_2204);
nor U4117 (N_4117,In_359,In_1114);
nand U4118 (N_4118,In_2428,In_1186);
nand U4119 (N_4119,In_1218,In_922);
nand U4120 (N_4120,In_526,In_1602);
nand U4121 (N_4121,In_137,In_902);
nor U4122 (N_4122,In_2461,In_1885);
nand U4123 (N_4123,In_945,In_1311);
nor U4124 (N_4124,In_1039,In_670);
or U4125 (N_4125,In_727,In_974);
nor U4126 (N_4126,In_1601,In_259);
or U4127 (N_4127,In_2164,In_126);
or U4128 (N_4128,In_2034,In_1423);
nand U4129 (N_4129,In_693,In_1338);
xor U4130 (N_4130,In_2380,In_1710);
xor U4131 (N_4131,In_2241,In_2438);
nor U4132 (N_4132,In_752,In_1576);
and U4133 (N_4133,In_823,In_1818);
nand U4134 (N_4134,In_777,In_135);
nand U4135 (N_4135,In_442,In_1778);
and U4136 (N_4136,In_2488,In_533);
or U4137 (N_4137,In_594,In_1495);
or U4138 (N_4138,In_654,In_16);
nor U4139 (N_4139,In_1184,In_762);
xnor U4140 (N_4140,In_750,In_733);
or U4141 (N_4141,In_1759,In_2080);
nand U4142 (N_4142,In_900,In_1655);
nand U4143 (N_4143,In_293,In_2403);
xnor U4144 (N_4144,In_1543,In_1918);
xor U4145 (N_4145,In_1252,In_861);
nor U4146 (N_4146,In_1416,In_1296);
and U4147 (N_4147,In_603,In_1584);
and U4148 (N_4148,In_1149,In_340);
xnor U4149 (N_4149,In_936,In_491);
nor U4150 (N_4150,In_1404,In_296);
or U4151 (N_4151,In_1227,In_1174);
or U4152 (N_4152,In_2104,In_2210);
nand U4153 (N_4153,In_413,In_1544);
nand U4154 (N_4154,In_2416,In_655);
xor U4155 (N_4155,In_860,In_1154);
nor U4156 (N_4156,In_1488,In_2171);
nand U4157 (N_4157,In_1182,In_2026);
xor U4158 (N_4158,In_2496,In_2360);
or U4159 (N_4159,In_1854,In_2304);
xnor U4160 (N_4160,In_1713,In_2124);
nand U4161 (N_4161,In_315,In_701);
and U4162 (N_4162,In_1554,In_719);
nor U4163 (N_4163,In_403,In_1316);
nand U4164 (N_4164,In_268,In_1220);
and U4165 (N_4165,In_1125,In_1083);
xnor U4166 (N_4166,In_2247,In_2120);
xor U4167 (N_4167,In_659,In_1088);
xor U4168 (N_4168,In_1414,In_2069);
or U4169 (N_4169,In_1986,In_160);
nand U4170 (N_4170,In_2262,In_2186);
xnor U4171 (N_4171,In_1397,In_885);
or U4172 (N_4172,In_2150,In_991);
xnor U4173 (N_4173,In_940,In_2017);
nor U4174 (N_4174,In_354,In_631);
or U4175 (N_4175,In_1820,In_2010);
or U4176 (N_4176,In_51,In_2400);
xnor U4177 (N_4177,In_1715,In_479);
nand U4178 (N_4178,In_2384,In_2131);
or U4179 (N_4179,In_300,In_1416);
xor U4180 (N_4180,In_1268,In_1011);
nor U4181 (N_4181,In_1230,In_1475);
or U4182 (N_4182,In_428,In_307);
and U4183 (N_4183,In_1869,In_2496);
xnor U4184 (N_4184,In_938,In_677);
nand U4185 (N_4185,In_79,In_1515);
or U4186 (N_4186,In_599,In_745);
xnor U4187 (N_4187,In_1681,In_1468);
xnor U4188 (N_4188,In_672,In_2213);
nand U4189 (N_4189,In_234,In_691);
nand U4190 (N_4190,In_2434,In_1242);
nand U4191 (N_4191,In_2060,In_1750);
nor U4192 (N_4192,In_2266,In_1141);
nor U4193 (N_4193,In_1134,In_380);
xor U4194 (N_4194,In_5,In_1425);
or U4195 (N_4195,In_1454,In_1762);
or U4196 (N_4196,In_1932,In_2102);
and U4197 (N_4197,In_1667,In_1746);
or U4198 (N_4198,In_1273,In_1880);
nand U4199 (N_4199,In_1492,In_466);
or U4200 (N_4200,In_1261,In_83);
nor U4201 (N_4201,In_1501,In_2472);
and U4202 (N_4202,In_921,In_2439);
nor U4203 (N_4203,In_552,In_1112);
and U4204 (N_4204,In_190,In_484);
nand U4205 (N_4205,In_796,In_53);
nor U4206 (N_4206,In_1873,In_2482);
nor U4207 (N_4207,In_2482,In_2287);
and U4208 (N_4208,In_1501,In_1831);
or U4209 (N_4209,In_1010,In_1072);
and U4210 (N_4210,In_1179,In_1097);
or U4211 (N_4211,In_1827,In_838);
xnor U4212 (N_4212,In_260,In_2362);
and U4213 (N_4213,In_2087,In_1385);
nand U4214 (N_4214,In_1124,In_1184);
xor U4215 (N_4215,In_870,In_472);
nand U4216 (N_4216,In_1720,In_1133);
and U4217 (N_4217,In_1269,In_1252);
nor U4218 (N_4218,In_1863,In_153);
xnor U4219 (N_4219,In_774,In_927);
or U4220 (N_4220,In_2077,In_1673);
nand U4221 (N_4221,In_1758,In_2466);
and U4222 (N_4222,In_515,In_1653);
or U4223 (N_4223,In_1614,In_1801);
and U4224 (N_4224,In_2469,In_1915);
nor U4225 (N_4225,In_595,In_170);
or U4226 (N_4226,In_1973,In_994);
nand U4227 (N_4227,In_1923,In_2026);
or U4228 (N_4228,In_1468,In_707);
xnor U4229 (N_4229,In_1889,In_614);
and U4230 (N_4230,In_1819,In_2242);
nand U4231 (N_4231,In_123,In_27);
and U4232 (N_4232,In_599,In_2298);
xor U4233 (N_4233,In_503,In_1679);
xnor U4234 (N_4234,In_474,In_559);
nand U4235 (N_4235,In_1006,In_276);
and U4236 (N_4236,In_1957,In_2494);
or U4237 (N_4237,In_2397,In_1780);
or U4238 (N_4238,In_1393,In_2308);
or U4239 (N_4239,In_762,In_2162);
and U4240 (N_4240,In_2420,In_861);
and U4241 (N_4241,In_1447,In_2116);
or U4242 (N_4242,In_663,In_1338);
or U4243 (N_4243,In_1024,In_2088);
nor U4244 (N_4244,In_6,In_1503);
or U4245 (N_4245,In_726,In_737);
or U4246 (N_4246,In_114,In_800);
nor U4247 (N_4247,In_2249,In_2107);
xnor U4248 (N_4248,In_22,In_1730);
or U4249 (N_4249,In_2098,In_1304);
or U4250 (N_4250,In_766,In_1467);
or U4251 (N_4251,In_256,In_379);
and U4252 (N_4252,In_784,In_1185);
and U4253 (N_4253,In_113,In_1482);
nand U4254 (N_4254,In_626,In_2348);
or U4255 (N_4255,In_1044,In_1348);
and U4256 (N_4256,In_1140,In_1319);
nand U4257 (N_4257,In_1887,In_1504);
nand U4258 (N_4258,In_1643,In_494);
nor U4259 (N_4259,In_86,In_1898);
nand U4260 (N_4260,In_1098,In_1916);
nand U4261 (N_4261,In_699,In_505);
and U4262 (N_4262,In_2090,In_1653);
or U4263 (N_4263,In_1754,In_1717);
nor U4264 (N_4264,In_2062,In_518);
or U4265 (N_4265,In_2342,In_335);
or U4266 (N_4266,In_2156,In_361);
or U4267 (N_4267,In_1073,In_1418);
and U4268 (N_4268,In_1516,In_110);
or U4269 (N_4269,In_1760,In_143);
nor U4270 (N_4270,In_1449,In_1088);
or U4271 (N_4271,In_1102,In_2180);
xor U4272 (N_4272,In_750,In_1350);
nand U4273 (N_4273,In_196,In_941);
or U4274 (N_4274,In_2071,In_1705);
nor U4275 (N_4275,In_2147,In_712);
nand U4276 (N_4276,In_1936,In_1764);
nor U4277 (N_4277,In_1302,In_928);
nand U4278 (N_4278,In_1410,In_1554);
and U4279 (N_4279,In_1077,In_787);
or U4280 (N_4280,In_421,In_37);
or U4281 (N_4281,In_2068,In_1502);
xnor U4282 (N_4282,In_1355,In_1769);
nor U4283 (N_4283,In_137,In_508);
and U4284 (N_4284,In_1927,In_1135);
xnor U4285 (N_4285,In_804,In_304);
or U4286 (N_4286,In_1468,In_604);
nor U4287 (N_4287,In_1095,In_2053);
nand U4288 (N_4288,In_2385,In_1828);
nand U4289 (N_4289,In_1783,In_1337);
nor U4290 (N_4290,In_2251,In_1910);
xnor U4291 (N_4291,In_1737,In_406);
nand U4292 (N_4292,In_704,In_1645);
nand U4293 (N_4293,In_873,In_1055);
nand U4294 (N_4294,In_1655,In_1142);
or U4295 (N_4295,In_1436,In_698);
and U4296 (N_4296,In_1967,In_576);
or U4297 (N_4297,In_1281,In_1996);
nand U4298 (N_4298,In_2154,In_2355);
nand U4299 (N_4299,In_157,In_858);
xor U4300 (N_4300,In_432,In_1466);
nor U4301 (N_4301,In_94,In_297);
nor U4302 (N_4302,In_907,In_1263);
xnor U4303 (N_4303,In_1935,In_1109);
nand U4304 (N_4304,In_1476,In_21);
nor U4305 (N_4305,In_433,In_1497);
or U4306 (N_4306,In_2176,In_468);
and U4307 (N_4307,In_1192,In_1924);
xnor U4308 (N_4308,In_1514,In_2116);
and U4309 (N_4309,In_1814,In_1486);
nor U4310 (N_4310,In_88,In_750);
xor U4311 (N_4311,In_1438,In_1101);
nor U4312 (N_4312,In_1130,In_1734);
or U4313 (N_4313,In_2283,In_1629);
nor U4314 (N_4314,In_501,In_1483);
xor U4315 (N_4315,In_1538,In_1645);
and U4316 (N_4316,In_763,In_2388);
nand U4317 (N_4317,In_824,In_1421);
and U4318 (N_4318,In_1044,In_1717);
nand U4319 (N_4319,In_1474,In_727);
and U4320 (N_4320,In_901,In_1802);
xnor U4321 (N_4321,In_2168,In_1494);
nor U4322 (N_4322,In_2335,In_1626);
or U4323 (N_4323,In_938,In_1996);
and U4324 (N_4324,In_712,In_765);
xor U4325 (N_4325,In_346,In_2158);
xnor U4326 (N_4326,In_149,In_650);
and U4327 (N_4327,In_971,In_823);
or U4328 (N_4328,In_541,In_1465);
nor U4329 (N_4329,In_1041,In_1103);
nor U4330 (N_4330,In_44,In_1259);
xnor U4331 (N_4331,In_1266,In_1414);
or U4332 (N_4332,In_1893,In_2394);
and U4333 (N_4333,In_2212,In_560);
or U4334 (N_4334,In_2181,In_433);
or U4335 (N_4335,In_2479,In_1286);
and U4336 (N_4336,In_1010,In_2056);
or U4337 (N_4337,In_2262,In_2209);
nand U4338 (N_4338,In_1644,In_496);
nor U4339 (N_4339,In_555,In_730);
or U4340 (N_4340,In_1154,In_1340);
and U4341 (N_4341,In_2170,In_2296);
and U4342 (N_4342,In_803,In_1385);
nor U4343 (N_4343,In_1751,In_1743);
nand U4344 (N_4344,In_299,In_1398);
nor U4345 (N_4345,In_865,In_1294);
nor U4346 (N_4346,In_294,In_1566);
nand U4347 (N_4347,In_485,In_1186);
nand U4348 (N_4348,In_1861,In_890);
nor U4349 (N_4349,In_1272,In_1319);
or U4350 (N_4350,In_1033,In_2147);
or U4351 (N_4351,In_2199,In_1600);
or U4352 (N_4352,In_2323,In_83);
and U4353 (N_4353,In_990,In_32);
nor U4354 (N_4354,In_1060,In_1750);
and U4355 (N_4355,In_1400,In_1946);
nor U4356 (N_4356,In_2069,In_2151);
nand U4357 (N_4357,In_1582,In_1225);
nand U4358 (N_4358,In_452,In_552);
xnor U4359 (N_4359,In_890,In_2160);
nand U4360 (N_4360,In_2464,In_1229);
xnor U4361 (N_4361,In_768,In_914);
xnor U4362 (N_4362,In_1367,In_710);
nor U4363 (N_4363,In_1270,In_1712);
nor U4364 (N_4364,In_219,In_2090);
and U4365 (N_4365,In_2295,In_670);
and U4366 (N_4366,In_1828,In_2432);
nor U4367 (N_4367,In_1935,In_1075);
or U4368 (N_4368,In_1941,In_576);
nand U4369 (N_4369,In_842,In_601);
nor U4370 (N_4370,In_1603,In_2306);
xor U4371 (N_4371,In_2362,In_2076);
nand U4372 (N_4372,In_779,In_2094);
xnor U4373 (N_4373,In_1170,In_717);
nor U4374 (N_4374,In_203,In_1821);
nor U4375 (N_4375,In_2346,In_1416);
nand U4376 (N_4376,In_898,In_1101);
and U4377 (N_4377,In_487,In_2474);
nand U4378 (N_4378,In_1955,In_518);
or U4379 (N_4379,In_27,In_262);
xor U4380 (N_4380,In_486,In_2224);
or U4381 (N_4381,In_2086,In_1771);
xor U4382 (N_4382,In_2002,In_1624);
nand U4383 (N_4383,In_2026,In_2040);
or U4384 (N_4384,In_1344,In_2052);
xnor U4385 (N_4385,In_1941,In_1848);
nand U4386 (N_4386,In_81,In_1255);
xor U4387 (N_4387,In_1760,In_735);
nand U4388 (N_4388,In_1421,In_1149);
xnor U4389 (N_4389,In_850,In_2358);
nand U4390 (N_4390,In_2113,In_200);
xnor U4391 (N_4391,In_1229,In_330);
or U4392 (N_4392,In_630,In_1372);
xnor U4393 (N_4393,In_2131,In_288);
xor U4394 (N_4394,In_2207,In_1828);
or U4395 (N_4395,In_1755,In_1321);
nand U4396 (N_4396,In_1015,In_1585);
nand U4397 (N_4397,In_991,In_2084);
nor U4398 (N_4398,In_1540,In_427);
or U4399 (N_4399,In_1613,In_1690);
nand U4400 (N_4400,In_2275,In_1030);
nand U4401 (N_4401,In_2466,In_63);
and U4402 (N_4402,In_2040,In_2100);
nor U4403 (N_4403,In_1061,In_366);
nand U4404 (N_4404,In_13,In_263);
nand U4405 (N_4405,In_1292,In_218);
and U4406 (N_4406,In_1980,In_744);
and U4407 (N_4407,In_821,In_1388);
and U4408 (N_4408,In_799,In_894);
nor U4409 (N_4409,In_629,In_2494);
or U4410 (N_4410,In_1634,In_1051);
and U4411 (N_4411,In_237,In_259);
xnor U4412 (N_4412,In_471,In_672);
or U4413 (N_4413,In_1206,In_429);
nand U4414 (N_4414,In_434,In_2402);
nor U4415 (N_4415,In_1262,In_204);
and U4416 (N_4416,In_1148,In_1080);
or U4417 (N_4417,In_2012,In_2395);
nand U4418 (N_4418,In_1096,In_2453);
nand U4419 (N_4419,In_1797,In_16);
or U4420 (N_4420,In_1976,In_1446);
nand U4421 (N_4421,In_898,In_2293);
or U4422 (N_4422,In_697,In_1561);
nor U4423 (N_4423,In_147,In_1704);
nor U4424 (N_4424,In_1313,In_1523);
nand U4425 (N_4425,In_1695,In_2027);
xor U4426 (N_4426,In_927,In_1919);
nor U4427 (N_4427,In_1765,In_174);
or U4428 (N_4428,In_1410,In_1422);
nand U4429 (N_4429,In_750,In_2169);
xor U4430 (N_4430,In_1321,In_2314);
nor U4431 (N_4431,In_538,In_567);
or U4432 (N_4432,In_2087,In_2071);
nand U4433 (N_4433,In_807,In_109);
nor U4434 (N_4434,In_2150,In_1086);
nand U4435 (N_4435,In_1760,In_1865);
nor U4436 (N_4436,In_346,In_2113);
xnor U4437 (N_4437,In_957,In_991);
or U4438 (N_4438,In_520,In_559);
nand U4439 (N_4439,In_1062,In_35);
xor U4440 (N_4440,In_246,In_649);
xnor U4441 (N_4441,In_1986,In_484);
xor U4442 (N_4442,In_2049,In_1321);
or U4443 (N_4443,In_2016,In_577);
and U4444 (N_4444,In_379,In_2093);
xnor U4445 (N_4445,In_24,In_70);
xor U4446 (N_4446,In_1989,In_2279);
or U4447 (N_4447,In_626,In_1961);
xnor U4448 (N_4448,In_2426,In_2171);
xnor U4449 (N_4449,In_589,In_808);
or U4450 (N_4450,In_1592,In_1492);
nor U4451 (N_4451,In_1883,In_819);
xnor U4452 (N_4452,In_841,In_72);
and U4453 (N_4453,In_1431,In_1407);
and U4454 (N_4454,In_340,In_2335);
xor U4455 (N_4455,In_24,In_564);
nand U4456 (N_4456,In_2407,In_2449);
xor U4457 (N_4457,In_975,In_1859);
and U4458 (N_4458,In_2496,In_318);
xnor U4459 (N_4459,In_744,In_21);
and U4460 (N_4460,In_1660,In_369);
nor U4461 (N_4461,In_2246,In_2307);
and U4462 (N_4462,In_184,In_739);
xnor U4463 (N_4463,In_938,In_664);
and U4464 (N_4464,In_1526,In_944);
nor U4465 (N_4465,In_191,In_1698);
nor U4466 (N_4466,In_991,In_90);
or U4467 (N_4467,In_1900,In_2436);
and U4468 (N_4468,In_2164,In_1278);
and U4469 (N_4469,In_1197,In_441);
nand U4470 (N_4470,In_2130,In_1782);
and U4471 (N_4471,In_140,In_2065);
nand U4472 (N_4472,In_2110,In_1914);
xnor U4473 (N_4473,In_142,In_1760);
nor U4474 (N_4474,In_1619,In_1630);
nand U4475 (N_4475,In_2460,In_1645);
xor U4476 (N_4476,In_17,In_1691);
or U4477 (N_4477,In_886,In_464);
xnor U4478 (N_4478,In_1679,In_772);
and U4479 (N_4479,In_1325,In_1941);
nor U4480 (N_4480,In_2205,In_1620);
or U4481 (N_4481,In_2095,In_783);
nor U4482 (N_4482,In_1027,In_2190);
nor U4483 (N_4483,In_1530,In_379);
nand U4484 (N_4484,In_367,In_286);
nand U4485 (N_4485,In_972,In_569);
nand U4486 (N_4486,In_2486,In_1819);
nor U4487 (N_4487,In_1315,In_2294);
or U4488 (N_4488,In_336,In_2465);
nor U4489 (N_4489,In_596,In_1622);
xor U4490 (N_4490,In_1972,In_2416);
nor U4491 (N_4491,In_856,In_1970);
xnor U4492 (N_4492,In_100,In_1347);
or U4493 (N_4493,In_618,In_2261);
nand U4494 (N_4494,In_957,In_867);
and U4495 (N_4495,In_25,In_27);
and U4496 (N_4496,In_1253,In_260);
and U4497 (N_4497,In_357,In_312);
nand U4498 (N_4498,In_1117,In_2045);
or U4499 (N_4499,In_12,In_229);
nand U4500 (N_4500,In_23,In_1282);
nand U4501 (N_4501,In_1426,In_1355);
nor U4502 (N_4502,In_219,In_141);
xor U4503 (N_4503,In_1196,In_2404);
and U4504 (N_4504,In_2006,In_1812);
xnor U4505 (N_4505,In_93,In_1348);
nand U4506 (N_4506,In_1710,In_196);
or U4507 (N_4507,In_601,In_1277);
nand U4508 (N_4508,In_2372,In_702);
or U4509 (N_4509,In_1385,In_465);
and U4510 (N_4510,In_1564,In_794);
or U4511 (N_4511,In_937,In_1944);
and U4512 (N_4512,In_1598,In_2473);
xnor U4513 (N_4513,In_2109,In_1226);
nor U4514 (N_4514,In_1038,In_1412);
nor U4515 (N_4515,In_1876,In_1202);
nand U4516 (N_4516,In_1568,In_2427);
and U4517 (N_4517,In_2108,In_1579);
or U4518 (N_4518,In_1133,In_1356);
xor U4519 (N_4519,In_1733,In_963);
or U4520 (N_4520,In_966,In_1344);
nand U4521 (N_4521,In_2154,In_1231);
nand U4522 (N_4522,In_66,In_1556);
nor U4523 (N_4523,In_76,In_2182);
and U4524 (N_4524,In_1665,In_2409);
or U4525 (N_4525,In_1844,In_1200);
nor U4526 (N_4526,In_2242,In_2020);
and U4527 (N_4527,In_724,In_487);
nor U4528 (N_4528,In_703,In_966);
nand U4529 (N_4529,In_1129,In_1589);
or U4530 (N_4530,In_595,In_2023);
or U4531 (N_4531,In_734,In_970);
nand U4532 (N_4532,In_827,In_912);
or U4533 (N_4533,In_1481,In_693);
nand U4534 (N_4534,In_258,In_1208);
and U4535 (N_4535,In_2000,In_2489);
nor U4536 (N_4536,In_365,In_975);
and U4537 (N_4537,In_2272,In_1921);
xor U4538 (N_4538,In_1479,In_333);
xnor U4539 (N_4539,In_1402,In_270);
nor U4540 (N_4540,In_1269,In_230);
nor U4541 (N_4541,In_2310,In_1857);
and U4542 (N_4542,In_1008,In_58);
nor U4543 (N_4543,In_2115,In_1652);
nand U4544 (N_4544,In_1610,In_30);
xor U4545 (N_4545,In_1523,In_1583);
xnor U4546 (N_4546,In_1371,In_665);
and U4547 (N_4547,In_790,In_777);
nand U4548 (N_4548,In_904,In_1169);
and U4549 (N_4549,In_1591,In_1783);
or U4550 (N_4550,In_1012,In_2472);
xor U4551 (N_4551,In_1455,In_1585);
nor U4552 (N_4552,In_2233,In_2159);
nand U4553 (N_4553,In_1562,In_1773);
nor U4554 (N_4554,In_1602,In_916);
xor U4555 (N_4555,In_701,In_1288);
nor U4556 (N_4556,In_540,In_942);
nand U4557 (N_4557,In_522,In_151);
and U4558 (N_4558,In_2110,In_1566);
xnor U4559 (N_4559,In_1738,In_2018);
nand U4560 (N_4560,In_2483,In_66);
nor U4561 (N_4561,In_2354,In_2230);
nor U4562 (N_4562,In_863,In_557);
nand U4563 (N_4563,In_368,In_1239);
nand U4564 (N_4564,In_2142,In_1171);
xnor U4565 (N_4565,In_742,In_547);
nor U4566 (N_4566,In_660,In_910);
and U4567 (N_4567,In_110,In_1316);
or U4568 (N_4568,In_1806,In_1416);
or U4569 (N_4569,In_2110,In_1399);
or U4570 (N_4570,In_1720,In_2467);
and U4571 (N_4571,In_1945,In_103);
nor U4572 (N_4572,In_1296,In_1233);
xnor U4573 (N_4573,In_2001,In_1365);
xnor U4574 (N_4574,In_1280,In_834);
xor U4575 (N_4575,In_1048,In_2457);
xor U4576 (N_4576,In_864,In_216);
nor U4577 (N_4577,In_429,In_1180);
nand U4578 (N_4578,In_1376,In_2244);
xnor U4579 (N_4579,In_1540,In_760);
or U4580 (N_4580,In_2320,In_2326);
xnor U4581 (N_4581,In_114,In_443);
and U4582 (N_4582,In_705,In_1983);
xnor U4583 (N_4583,In_1621,In_1575);
and U4584 (N_4584,In_2387,In_1854);
nand U4585 (N_4585,In_1137,In_505);
and U4586 (N_4586,In_818,In_2292);
nor U4587 (N_4587,In_2200,In_2013);
and U4588 (N_4588,In_766,In_1373);
or U4589 (N_4589,In_1311,In_1823);
and U4590 (N_4590,In_1385,In_1937);
xnor U4591 (N_4591,In_850,In_1065);
or U4592 (N_4592,In_2271,In_1030);
or U4593 (N_4593,In_601,In_125);
xor U4594 (N_4594,In_1352,In_1962);
xnor U4595 (N_4595,In_1690,In_1989);
or U4596 (N_4596,In_2240,In_922);
nand U4597 (N_4597,In_1819,In_741);
xnor U4598 (N_4598,In_1178,In_1243);
nand U4599 (N_4599,In_1434,In_1828);
and U4600 (N_4600,In_1512,In_1547);
nor U4601 (N_4601,In_1898,In_1256);
and U4602 (N_4602,In_2086,In_2090);
or U4603 (N_4603,In_1815,In_1324);
nand U4604 (N_4604,In_2226,In_1678);
and U4605 (N_4605,In_2018,In_2323);
or U4606 (N_4606,In_1347,In_1662);
nand U4607 (N_4607,In_2031,In_591);
nand U4608 (N_4608,In_428,In_1500);
nor U4609 (N_4609,In_1462,In_1099);
and U4610 (N_4610,In_1878,In_1389);
nor U4611 (N_4611,In_726,In_2216);
xor U4612 (N_4612,In_134,In_1591);
xor U4613 (N_4613,In_2373,In_1411);
nand U4614 (N_4614,In_326,In_2203);
or U4615 (N_4615,In_1658,In_1083);
and U4616 (N_4616,In_1185,In_1142);
and U4617 (N_4617,In_757,In_1566);
nand U4618 (N_4618,In_1467,In_333);
nor U4619 (N_4619,In_2225,In_1238);
xor U4620 (N_4620,In_1256,In_2129);
nor U4621 (N_4621,In_367,In_1565);
nand U4622 (N_4622,In_1107,In_1938);
nand U4623 (N_4623,In_1728,In_2414);
and U4624 (N_4624,In_1500,In_2060);
and U4625 (N_4625,In_333,In_1452);
nor U4626 (N_4626,In_784,In_1868);
xor U4627 (N_4627,In_1129,In_1113);
nor U4628 (N_4628,In_1884,In_695);
or U4629 (N_4629,In_2261,In_1339);
and U4630 (N_4630,In_855,In_37);
nand U4631 (N_4631,In_59,In_1636);
or U4632 (N_4632,In_1232,In_417);
xnor U4633 (N_4633,In_2280,In_962);
nor U4634 (N_4634,In_63,In_174);
and U4635 (N_4635,In_2064,In_1801);
or U4636 (N_4636,In_853,In_557);
xnor U4637 (N_4637,In_2452,In_1654);
or U4638 (N_4638,In_571,In_559);
nor U4639 (N_4639,In_201,In_697);
xnor U4640 (N_4640,In_63,In_2434);
nor U4641 (N_4641,In_1835,In_424);
nand U4642 (N_4642,In_2285,In_135);
xnor U4643 (N_4643,In_530,In_17);
xor U4644 (N_4644,In_805,In_2160);
and U4645 (N_4645,In_1148,In_2203);
xnor U4646 (N_4646,In_277,In_2472);
or U4647 (N_4647,In_1317,In_1691);
or U4648 (N_4648,In_933,In_1591);
and U4649 (N_4649,In_199,In_928);
nor U4650 (N_4650,In_230,In_879);
or U4651 (N_4651,In_407,In_703);
nand U4652 (N_4652,In_1779,In_1201);
or U4653 (N_4653,In_716,In_1175);
or U4654 (N_4654,In_450,In_1403);
and U4655 (N_4655,In_759,In_901);
nor U4656 (N_4656,In_2040,In_2476);
xnor U4657 (N_4657,In_1918,In_427);
and U4658 (N_4658,In_124,In_1589);
nor U4659 (N_4659,In_1116,In_488);
nand U4660 (N_4660,In_918,In_516);
nor U4661 (N_4661,In_2134,In_1620);
nor U4662 (N_4662,In_2499,In_136);
or U4663 (N_4663,In_1567,In_2043);
xor U4664 (N_4664,In_1637,In_808);
xnor U4665 (N_4665,In_397,In_1637);
or U4666 (N_4666,In_2218,In_1133);
nor U4667 (N_4667,In_317,In_1137);
or U4668 (N_4668,In_686,In_620);
nand U4669 (N_4669,In_1040,In_1104);
or U4670 (N_4670,In_2326,In_1506);
nor U4671 (N_4671,In_761,In_1317);
nor U4672 (N_4672,In_1333,In_2121);
nor U4673 (N_4673,In_54,In_1327);
xnor U4674 (N_4674,In_1682,In_1353);
nand U4675 (N_4675,In_1239,In_646);
xor U4676 (N_4676,In_2326,In_1900);
nor U4677 (N_4677,In_745,In_1209);
nor U4678 (N_4678,In_2067,In_204);
xnor U4679 (N_4679,In_754,In_2142);
nand U4680 (N_4680,In_127,In_2122);
nor U4681 (N_4681,In_307,In_2297);
xor U4682 (N_4682,In_2143,In_549);
xor U4683 (N_4683,In_1245,In_1658);
nor U4684 (N_4684,In_1599,In_2140);
and U4685 (N_4685,In_1240,In_1056);
nor U4686 (N_4686,In_1371,In_1775);
nand U4687 (N_4687,In_2293,In_316);
and U4688 (N_4688,In_438,In_672);
and U4689 (N_4689,In_2478,In_2266);
nor U4690 (N_4690,In_298,In_1042);
nand U4691 (N_4691,In_2215,In_2289);
or U4692 (N_4692,In_1274,In_2306);
or U4693 (N_4693,In_1718,In_1843);
nand U4694 (N_4694,In_74,In_2473);
nand U4695 (N_4695,In_186,In_1622);
nand U4696 (N_4696,In_559,In_625);
nor U4697 (N_4697,In_940,In_1396);
xnor U4698 (N_4698,In_491,In_385);
xnor U4699 (N_4699,In_1770,In_1865);
and U4700 (N_4700,In_1583,In_493);
nor U4701 (N_4701,In_1687,In_1584);
nor U4702 (N_4702,In_366,In_1738);
nand U4703 (N_4703,In_2458,In_275);
nor U4704 (N_4704,In_2245,In_881);
and U4705 (N_4705,In_2384,In_482);
nand U4706 (N_4706,In_1706,In_1264);
and U4707 (N_4707,In_1016,In_139);
xnor U4708 (N_4708,In_1286,In_689);
and U4709 (N_4709,In_635,In_1272);
nand U4710 (N_4710,In_1290,In_2252);
nor U4711 (N_4711,In_534,In_2009);
nand U4712 (N_4712,In_1633,In_162);
xor U4713 (N_4713,In_425,In_1781);
nor U4714 (N_4714,In_1876,In_2464);
or U4715 (N_4715,In_979,In_1892);
nor U4716 (N_4716,In_224,In_704);
nand U4717 (N_4717,In_588,In_2359);
xor U4718 (N_4718,In_757,In_2460);
and U4719 (N_4719,In_2002,In_2242);
xor U4720 (N_4720,In_340,In_373);
xnor U4721 (N_4721,In_1792,In_2355);
xor U4722 (N_4722,In_163,In_1445);
xnor U4723 (N_4723,In_1605,In_10);
or U4724 (N_4724,In_1249,In_1634);
and U4725 (N_4725,In_20,In_1023);
nand U4726 (N_4726,In_2435,In_2388);
nand U4727 (N_4727,In_1527,In_213);
or U4728 (N_4728,In_924,In_674);
nand U4729 (N_4729,In_529,In_642);
and U4730 (N_4730,In_464,In_2209);
xor U4731 (N_4731,In_2457,In_55);
or U4732 (N_4732,In_2269,In_1438);
and U4733 (N_4733,In_2250,In_1171);
or U4734 (N_4734,In_908,In_146);
or U4735 (N_4735,In_43,In_1655);
and U4736 (N_4736,In_726,In_2256);
and U4737 (N_4737,In_1610,In_1826);
or U4738 (N_4738,In_1317,In_38);
and U4739 (N_4739,In_1545,In_343);
nor U4740 (N_4740,In_1370,In_2265);
and U4741 (N_4741,In_1075,In_2060);
xnor U4742 (N_4742,In_1921,In_1289);
nor U4743 (N_4743,In_118,In_168);
xnor U4744 (N_4744,In_895,In_948);
xnor U4745 (N_4745,In_412,In_1133);
or U4746 (N_4746,In_1432,In_1463);
nand U4747 (N_4747,In_2287,In_1916);
nand U4748 (N_4748,In_1684,In_844);
or U4749 (N_4749,In_2103,In_2426);
nand U4750 (N_4750,In_1418,In_1029);
nor U4751 (N_4751,In_2138,In_347);
xor U4752 (N_4752,In_179,In_981);
and U4753 (N_4753,In_1782,In_707);
nor U4754 (N_4754,In_1934,In_2059);
nor U4755 (N_4755,In_2409,In_1869);
or U4756 (N_4756,In_1287,In_2358);
and U4757 (N_4757,In_2418,In_1651);
or U4758 (N_4758,In_1038,In_1899);
nor U4759 (N_4759,In_1117,In_164);
nor U4760 (N_4760,In_785,In_1280);
or U4761 (N_4761,In_338,In_515);
or U4762 (N_4762,In_1150,In_1277);
nand U4763 (N_4763,In_1904,In_769);
and U4764 (N_4764,In_1561,In_2244);
nor U4765 (N_4765,In_1150,In_1330);
xnor U4766 (N_4766,In_107,In_817);
nand U4767 (N_4767,In_38,In_863);
nor U4768 (N_4768,In_1159,In_966);
nand U4769 (N_4769,In_1403,In_579);
nand U4770 (N_4770,In_1338,In_328);
nor U4771 (N_4771,In_999,In_406);
or U4772 (N_4772,In_121,In_1878);
xor U4773 (N_4773,In_304,In_2258);
and U4774 (N_4774,In_751,In_1692);
or U4775 (N_4775,In_1627,In_1512);
and U4776 (N_4776,In_1488,In_681);
xnor U4777 (N_4777,In_1892,In_1084);
xnor U4778 (N_4778,In_906,In_937);
or U4779 (N_4779,In_1987,In_2323);
nand U4780 (N_4780,In_1603,In_2001);
or U4781 (N_4781,In_1416,In_1187);
nor U4782 (N_4782,In_195,In_2129);
or U4783 (N_4783,In_811,In_1759);
nor U4784 (N_4784,In_952,In_2185);
nand U4785 (N_4785,In_722,In_785);
nor U4786 (N_4786,In_1912,In_2269);
nor U4787 (N_4787,In_673,In_2210);
nor U4788 (N_4788,In_318,In_1116);
and U4789 (N_4789,In_2177,In_1798);
nor U4790 (N_4790,In_574,In_1852);
and U4791 (N_4791,In_1871,In_2458);
nand U4792 (N_4792,In_578,In_1583);
nor U4793 (N_4793,In_955,In_610);
and U4794 (N_4794,In_934,In_219);
or U4795 (N_4795,In_1694,In_2242);
xnor U4796 (N_4796,In_359,In_207);
nor U4797 (N_4797,In_2104,In_54);
xor U4798 (N_4798,In_2423,In_662);
and U4799 (N_4799,In_1890,In_671);
xnor U4800 (N_4800,In_194,In_450);
or U4801 (N_4801,In_886,In_330);
nor U4802 (N_4802,In_2045,In_335);
and U4803 (N_4803,In_555,In_2247);
and U4804 (N_4804,In_2158,In_2269);
and U4805 (N_4805,In_2132,In_143);
xnor U4806 (N_4806,In_2388,In_102);
and U4807 (N_4807,In_1360,In_1855);
nor U4808 (N_4808,In_2044,In_579);
nand U4809 (N_4809,In_879,In_1833);
nand U4810 (N_4810,In_2456,In_926);
and U4811 (N_4811,In_580,In_1651);
xnor U4812 (N_4812,In_1001,In_993);
xnor U4813 (N_4813,In_1892,In_2090);
nor U4814 (N_4814,In_723,In_1769);
and U4815 (N_4815,In_556,In_743);
and U4816 (N_4816,In_590,In_1712);
nor U4817 (N_4817,In_825,In_1665);
nor U4818 (N_4818,In_784,In_1951);
nand U4819 (N_4819,In_1998,In_1754);
nor U4820 (N_4820,In_1211,In_635);
xnor U4821 (N_4821,In_1468,In_2208);
xor U4822 (N_4822,In_1807,In_391);
nand U4823 (N_4823,In_2451,In_1915);
nor U4824 (N_4824,In_1780,In_17);
nand U4825 (N_4825,In_1296,In_276);
nand U4826 (N_4826,In_1312,In_1676);
or U4827 (N_4827,In_536,In_837);
and U4828 (N_4828,In_1243,In_501);
and U4829 (N_4829,In_478,In_1035);
xor U4830 (N_4830,In_1185,In_559);
nand U4831 (N_4831,In_2251,In_623);
nor U4832 (N_4832,In_1242,In_228);
xnor U4833 (N_4833,In_997,In_1186);
or U4834 (N_4834,In_1769,In_1359);
or U4835 (N_4835,In_349,In_987);
nor U4836 (N_4836,In_1052,In_826);
nor U4837 (N_4837,In_1568,In_2009);
nand U4838 (N_4838,In_1165,In_880);
nor U4839 (N_4839,In_2327,In_454);
and U4840 (N_4840,In_1194,In_1430);
or U4841 (N_4841,In_1778,In_1940);
or U4842 (N_4842,In_1939,In_1768);
or U4843 (N_4843,In_533,In_1365);
xnor U4844 (N_4844,In_381,In_1752);
or U4845 (N_4845,In_1314,In_1178);
and U4846 (N_4846,In_1816,In_2393);
or U4847 (N_4847,In_1439,In_916);
or U4848 (N_4848,In_1201,In_724);
nor U4849 (N_4849,In_616,In_173);
nand U4850 (N_4850,In_1074,In_2026);
nor U4851 (N_4851,In_1864,In_959);
nor U4852 (N_4852,In_149,In_738);
or U4853 (N_4853,In_1323,In_2248);
and U4854 (N_4854,In_319,In_2108);
nor U4855 (N_4855,In_726,In_2406);
nor U4856 (N_4856,In_975,In_2093);
xor U4857 (N_4857,In_754,In_118);
and U4858 (N_4858,In_231,In_522);
or U4859 (N_4859,In_2386,In_1995);
nor U4860 (N_4860,In_1739,In_2195);
or U4861 (N_4861,In_129,In_182);
nor U4862 (N_4862,In_2064,In_26);
nand U4863 (N_4863,In_526,In_1007);
and U4864 (N_4864,In_2259,In_2294);
xor U4865 (N_4865,In_956,In_307);
nand U4866 (N_4866,In_97,In_1302);
nand U4867 (N_4867,In_1745,In_1479);
nand U4868 (N_4868,In_706,In_2426);
and U4869 (N_4869,In_2054,In_1027);
nor U4870 (N_4870,In_1433,In_628);
nand U4871 (N_4871,In_1312,In_1524);
and U4872 (N_4872,In_934,In_2062);
or U4873 (N_4873,In_2099,In_1582);
nor U4874 (N_4874,In_166,In_304);
xnor U4875 (N_4875,In_443,In_384);
xor U4876 (N_4876,In_1734,In_1074);
or U4877 (N_4877,In_66,In_2133);
or U4878 (N_4878,In_2159,In_1689);
nand U4879 (N_4879,In_1272,In_1915);
or U4880 (N_4880,In_2456,In_296);
and U4881 (N_4881,In_633,In_264);
nand U4882 (N_4882,In_2218,In_1555);
nand U4883 (N_4883,In_2326,In_2381);
or U4884 (N_4884,In_888,In_507);
or U4885 (N_4885,In_1973,In_1689);
nand U4886 (N_4886,In_1896,In_838);
or U4887 (N_4887,In_1919,In_876);
nand U4888 (N_4888,In_1410,In_1649);
nor U4889 (N_4889,In_1085,In_1530);
nor U4890 (N_4890,In_1468,In_191);
or U4891 (N_4891,In_531,In_277);
or U4892 (N_4892,In_707,In_1256);
nor U4893 (N_4893,In_1011,In_1657);
and U4894 (N_4894,In_270,In_673);
nor U4895 (N_4895,In_2211,In_2157);
or U4896 (N_4896,In_1718,In_1832);
or U4897 (N_4897,In_2106,In_1040);
or U4898 (N_4898,In_997,In_761);
or U4899 (N_4899,In_1270,In_330);
and U4900 (N_4900,In_220,In_2153);
xnor U4901 (N_4901,In_591,In_1010);
nand U4902 (N_4902,In_243,In_360);
nand U4903 (N_4903,In_899,In_1547);
xnor U4904 (N_4904,In_1574,In_2012);
nor U4905 (N_4905,In_1319,In_284);
nor U4906 (N_4906,In_1096,In_57);
or U4907 (N_4907,In_402,In_941);
nor U4908 (N_4908,In_525,In_1233);
nand U4909 (N_4909,In_683,In_721);
nand U4910 (N_4910,In_1295,In_914);
nor U4911 (N_4911,In_1569,In_1466);
nor U4912 (N_4912,In_2201,In_2266);
or U4913 (N_4913,In_1558,In_2460);
and U4914 (N_4914,In_1995,In_1067);
and U4915 (N_4915,In_1958,In_1436);
or U4916 (N_4916,In_2126,In_2170);
xor U4917 (N_4917,In_403,In_1100);
nand U4918 (N_4918,In_1772,In_1456);
or U4919 (N_4919,In_142,In_569);
xnor U4920 (N_4920,In_1286,In_1619);
or U4921 (N_4921,In_1598,In_2375);
or U4922 (N_4922,In_189,In_22);
nor U4923 (N_4923,In_598,In_1899);
xor U4924 (N_4924,In_1983,In_441);
xnor U4925 (N_4925,In_2384,In_363);
nor U4926 (N_4926,In_621,In_2004);
or U4927 (N_4927,In_1070,In_1254);
or U4928 (N_4928,In_437,In_926);
or U4929 (N_4929,In_376,In_113);
or U4930 (N_4930,In_812,In_2071);
and U4931 (N_4931,In_1079,In_2398);
xnor U4932 (N_4932,In_1998,In_1300);
xnor U4933 (N_4933,In_1488,In_1431);
nor U4934 (N_4934,In_2341,In_1382);
and U4935 (N_4935,In_630,In_2365);
or U4936 (N_4936,In_1998,In_1753);
xnor U4937 (N_4937,In_1756,In_1745);
and U4938 (N_4938,In_1935,In_2206);
nor U4939 (N_4939,In_1558,In_893);
or U4940 (N_4940,In_2074,In_1211);
or U4941 (N_4941,In_1791,In_1245);
and U4942 (N_4942,In_2070,In_1174);
or U4943 (N_4943,In_130,In_2450);
nand U4944 (N_4944,In_208,In_949);
nand U4945 (N_4945,In_1078,In_1864);
nand U4946 (N_4946,In_81,In_709);
and U4947 (N_4947,In_547,In_820);
and U4948 (N_4948,In_1902,In_2034);
and U4949 (N_4949,In_1317,In_516);
nor U4950 (N_4950,In_1470,In_750);
and U4951 (N_4951,In_1096,In_451);
xnor U4952 (N_4952,In_2427,In_1710);
nor U4953 (N_4953,In_1010,In_1143);
or U4954 (N_4954,In_1454,In_1375);
and U4955 (N_4955,In_1599,In_2314);
and U4956 (N_4956,In_1235,In_1992);
or U4957 (N_4957,In_1498,In_1916);
and U4958 (N_4958,In_2105,In_1006);
nand U4959 (N_4959,In_789,In_901);
nand U4960 (N_4960,In_1902,In_351);
nor U4961 (N_4961,In_1867,In_596);
or U4962 (N_4962,In_2235,In_1450);
and U4963 (N_4963,In_704,In_1826);
nor U4964 (N_4964,In_2275,In_2425);
and U4965 (N_4965,In_492,In_243);
nand U4966 (N_4966,In_2268,In_2493);
or U4967 (N_4967,In_2493,In_484);
nand U4968 (N_4968,In_1127,In_2083);
xnor U4969 (N_4969,In_935,In_254);
nor U4970 (N_4970,In_1746,In_681);
and U4971 (N_4971,In_1510,In_1995);
nand U4972 (N_4972,In_1579,In_751);
or U4973 (N_4973,In_1606,In_2340);
nand U4974 (N_4974,In_1343,In_1092);
and U4975 (N_4975,In_622,In_1963);
or U4976 (N_4976,In_2100,In_2216);
and U4977 (N_4977,In_457,In_2472);
xor U4978 (N_4978,In_1153,In_1951);
xnor U4979 (N_4979,In_255,In_1320);
nor U4980 (N_4980,In_1721,In_547);
or U4981 (N_4981,In_1846,In_2322);
or U4982 (N_4982,In_2163,In_2127);
xnor U4983 (N_4983,In_819,In_2253);
nand U4984 (N_4984,In_2463,In_1325);
nand U4985 (N_4985,In_1230,In_2118);
nand U4986 (N_4986,In_1311,In_1339);
or U4987 (N_4987,In_142,In_2372);
xnor U4988 (N_4988,In_2168,In_1854);
or U4989 (N_4989,In_1221,In_608);
and U4990 (N_4990,In_2411,In_2259);
or U4991 (N_4991,In_2194,In_749);
xnor U4992 (N_4992,In_826,In_189);
xnor U4993 (N_4993,In_1094,In_2142);
xor U4994 (N_4994,In_296,In_393);
or U4995 (N_4995,In_1866,In_2141);
and U4996 (N_4996,In_1782,In_2375);
xor U4997 (N_4997,In_875,In_1209);
xor U4998 (N_4998,In_11,In_775);
nor U4999 (N_4999,In_1777,In_673);
and U5000 (N_5000,N_4821,N_4747);
and U5001 (N_5001,N_600,N_1512);
or U5002 (N_5002,N_3307,N_978);
and U5003 (N_5003,N_1879,N_2414);
nand U5004 (N_5004,N_2653,N_3164);
nor U5005 (N_5005,N_4256,N_3831);
xor U5006 (N_5006,N_316,N_1833);
and U5007 (N_5007,N_630,N_3341);
nand U5008 (N_5008,N_4074,N_3953);
xnor U5009 (N_5009,N_749,N_1725);
xor U5010 (N_5010,N_3515,N_3658);
xnor U5011 (N_5011,N_2637,N_3118);
xor U5012 (N_5012,N_510,N_2994);
nand U5013 (N_5013,N_4158,N_1251);
nor U5014 (N_5014,N_2323,N_3866);
nand U5015 (N_5015,N_2718,N_1488);
xor U5016 (N_5016,N_4282,N_3322);
xor U5017 (N_5017,N_4626,N_57);
xor U5018 (N_5018,N_1942,N_3744);
nand U5019 (N_5019,N_1401,N_1418);
xnor U5020 (N_5020,N_4101,N_1231);
nand U5021 (N_5021,N_4011,N_705);
nor U5022 (N_5022,N_1151,N_335);
and U5023 (N_5023,N_2121,N_1069);
nand U5024 (N_5024,N_2353,N_2838);
nor U5025 (N_5025,N_4830,N_2768);
nand U5026 (N_5026,N_2343,N_4612);
nand U5027 (N_5027,N_2177,N_4871);
and U5028 (N_5028,N_3146,N_2828);
xnor U5029 (N_5029,N_2633,N_3149);
or U5030 (N_5030,N_912,N_1756);
nand U5031 (N_5031,N_1557,N_4810);
or U5032 (N_5032,N_3226,N_2801);
and U5033 (N_5033,N_1701,N_2008);
nor U5034 (N_5034,N_1502,N_4763);
nand U5035 (N_5035,N_2825,N_4765);
and U5036 (N_5036,N_3043,N_2341);
nand U5037 (N_5037,N_1332,N_713);
and U5038 (N_5038,N_1883,N_3134);
nor U5039 (N_5039,N_1227,N_1195);
and U5040 (N_5040,N_893,N_2473);
nor U5041 (N_5041,N_2829,N_97);
nand U5042 (N_5042,N_408,N_1885);
and U5043 (N_5043,N_3429,N_449);
nor U5044 (N_5044,N_200,N_568);
nor U5045 (N_5045,N_1853,N_3668);
or U5046 (N_5046,N_3313,N_107);
or U5047 (N_5047,N_3385,N_2329);
nand U5048 (N_5048,N_3034,N_423);
nor U5049 (N_5049,N_1472,N_2203);
xor U5050 (N_5050,N_3378,N_686);
xnor U5051 (N_5051,N_721,N_3985);
nand U5052 (N_5052,N_730,N_1580);
nor U5053 (N_5053,N_4990,N_3690);
or U5054 (N_5054,N_2227,N_254);
nand U5055 (N_5055,N_2101,N_711);
nand U5056 (N_5056,N_2474,N_4286);
nand U5057 (N_5057,N_4588,N_532);
and U5058 (N_5058,N_3003,N_3440);
xor U5059 (N_5059,N_3267,N_2907);
and U5060 (N_5060,N_2578,N_4002);
nand U5061 (N_5061,N_1789,N_2159);
and U5062 (N_5062,N_1666,N_4346);
or U5063 (N_5063,N_3035,N_1090);
and U5064 (N_5064,N_3206,N_4882);
nand U5065 (N_5065,N_2822,N_4958);
nand U5066 (N_5066,N_221,N_1587);
or U5067 (N_5067,N_2767,N_253);
or U5068 (N_5068,N_4215,N_2927);
and U5069 (N_5069,N_4940,N_3589);
nand U5070 (N_5070,N_645,N_351);
or U5071 (N_5071,N_4505,N_1830);
nor U5072 (N_5072,N_3350,N_661);
and U5073 (N_5073,N_3527,N_4644);
and U5074 (N_5074,N_3664,N_2076);
nand U5075 (N_5075,N_3305,N_3203);
nand U5076 (N_5076,N_4000,N_4760);
or U5077 (N_5077,N_2193,N_2562);
nand U5078 (N_5078,N_3768,N_601);
and U5079 (N_5079,N_1282,N_352);
nor U5080 (N_5080,N_387,N_3033);
or U5081 (N_5081,N_3657,N_3020);
nor U5082 (N_5082,N_2461,N_2097);
or U5083 (N_5083,N_548,N_4337);
and U5084 (N_5084,N_4849,N_1687);
nor U5085 (N_5085,N_65,N_4850);
and U5086 (N_5086,N_4417,N_672);
and U5087 (N_5087,N_608,N_1003);
nand U5088 (N_5088,N_806,N_823);
and U5089 (N_5089,N_3218,N_1422);
or U5090 (N_5090,N_3826,N_3158);
or U5091 (N_5091,N_265,N_4455);
nor U5092 (N_5092,N_4986,N_2873);
xnor U5093 (N_5093,N_2805,N_847);
nor U5094 (N_5094,N_4997,N_100);
xnor U5095 (N_5095,N_1364,N_4598);
and U5096 (N_5096,N_945,N_1530);
and U5097 (N_5097,N_3469,N_3063);
or U5098 (N_5098,N_4557,N_3078);
nand U5099 (N_5099,N_2627,N_1333);
or U5100 (N_5100,N_614,N_4895);
nand U5101 (N_5101,N_1609,N_3488);
or U5102 (N_5102,N_965,N_300);
or U5103 (N_5103,N_3924,N_4085);
or U5104 (N_5104,N_1057,N_3095);
nand U5105 (N_5105,N_2889,N_783);
and U5106 (N_5106,N_676,N_1178);
nand U5107 (N_5107,N_4229,N_3029);
nand U5108 (N_5108,N_1309,N_3789);
nor U5109 (N_5109,N_1420,N_500);
or U5110 (N_5110,N_1058,N_333);
xor U5111 (N_5111,N_790,N_2979);
xor U5112 (N_5112,N_2634,N_593);
and U5113 (N_5113,N_4679,N_1901);
nor U5114 (N_5114,N_952,N_4052);
nor U5115 (N_5115,N_577,N_1529);
or U5116 (N_5116,N_3448,N_1767);
or U5117 (N_5117,N_2275,N_491);
nand U5118 (N_5118,N_1636,N_4316);
or U5119 (N_5119,N_4336,N_620);
nand U5120 (N_5120,N_3685,N_1871);
or U5121 (N_5121,N_3144,N_3865);
nor U5122 (N_5122,N_3824,N_812);
and U5123 (N_5123,N_3625,N_3727);
xor U5124 (N_5124,N_4154,N_3002);
or U5125 (N_5125,N_505,N_3596);
nor U5126 (N_5126,N_2770,N_2220);
xnor U5127 (N_5127,N_281,N_1486);
nor U5128 (N_5128,N_2250,N_3537);
and U5129 (N_5129,N_3976,N_2245);
nor U5130 (N_5130,N_455,N_3004);
nor U5131 (N_5131,N_4613,N_739);
xnor U5132 (N_5132,N_2790,N_3266);
and U5133 (N_5133,N_305,N_4808);
and U5134 (N_5134,N_1367,N_2237);
xnor U5135 (N_5135,N_3125,N_218);
nor U5136 (N_5136,N_2964,N_2151);
nor U5137 (N_5137,N_4759,N_2643);
or U5138 (N_5138,N_2224,N_206);
and U5139 (N_5139,N_3573,N_4955);
and U5140 (N_5140,N_3918,N_1366);
xor U5141 (N_5141,N_3514,N_4624);
or U5142 (N_5142,N_3877,N_76);
or U5143 (N_5143,N_2863,N_4746);
nor U5144 (N_5144,N_1941,N_4929);
or U5145 (N_5145,N_781,N_5);
nor U5146 (N_5146,N_2748,N_2882);
or U5147 (N_5147,N_4996,N_181);
nand U5148 (N_5148,N_4192,N_1660);
and U5149 (N_5149,N_1320,N_2978);
xor U5150 (N_5150,N_1298,N_4711);
nand U5151 (N_5151,N_2750,N_557);
nand U5152 (N_5152,N_2688,N_3993);
xnor U5153 (N_5153,N_4903,N_2929);
and U5154 (N_5154,N_4174,N_1297);
or U5155 (N_5155,N_3421,N_2600);
and U5156 (N_5156,N_4607,N_309);
or U5157 (N_5157,N_3697,N_1435);
or U5158 (N_5158,N_4220,N_4800);
and U5159 (N_5159,N_89,N_1899);
xnor U5160 (N_5160,N_3108,N_59);
or U5161 (N_5161,N_4243,N_2904);
and U5162 (N_5162,N_2609,N_584);
nor U5163 (N_5163,N_3576,N_1188);
nor U5164 (N_5164,N_1338,N_1200);
nand U5165 (N_5165,N_2527,N_1651);
xor U5166 (N_5166,N_4031,N_451);
or U5167 (N_5167,N_764,N_2939);
nor U5168 (N_5168,N_255,N_1464);
nor U5169 (N_5169,N_3317,N_2854);
and U5170 (N_5170,N_4548,N_2467);
nor U5171 (N_5171,N_613,N_1475);
and U5172 (N_5172,N_483,N_3279);
xor U5173 (N_5173,N_1140,N_3446);
nand U5174 (N_5174,N_2523,N_656);
and U5175 (N_5175,N_4070,N_3060);
nand U5176 (N_5176,N_2859,N_2060);
nor U5177 (N_5177,N_3153,N_4604);
nand U5178 (N_5178,N_1874,N_4231);
or U5179 (N_5179,N_1841,N_343);
nand U5180 (N_5180,N_202,N_4854);
or U5181 (N_5181,N_3500,N_974);
xor U5182 (N_5182,N_27,N_4457);
xnor U5183 (N_5183,N_177,N_2);
and U5184 (N_5184,N_3368,N_4259);
and U5185 (N_5185,N_129,N_2355);
nor U5186 (N_5186,N_3339,N_2928);
nand U5187 (N_5187,N_1004,N_2447);
nand U5188 (N_5188,N_829,N_3445);
or U5189 (N_5189,N_2759,N_3601);
and U5190 (N_5190,N_2356,N_897);
and U5191 (N_5191,N_3564,N_391);
and U5192 (N_5192,N_4798,N_1768);
nor U5193 (N_5193,N_3869,N_2672);
or U5194 (N_5194,N_196,N_2552);
xor U5195 (N_5195,N_118,N_4780);
or U5196 (N_5196,N_4827,N_1116);
xnor U5197 (N_5197,N_3067,N_3502);
nand U5198 (N_5198,N_4384,N_2154);
and U5199 (N_5199,N_3324,N_1561);
nor U5200 (N_5200,N_3217,N_4556);
nand U5201 (N_5201,N_2391,N_1267);
and U5202 (N_5202,N_2708,N_1412);
xor U5203 (N_5203,N_3431,N_1066);
nand U5204 (N_5204,N_4773,N_719);
nor U5205 (N_5205,N_1832,N_2229);
nor U5206 (N_5206,N_2499,N_2235);
or U5207 (N_5207,N_150,N_3923);
xnor U5208 (N_5208,N_2170,N_4493);
nand U5209 (N_5209,N_1911,N_1797);
or U5210 (N_5210,N_4039,N_4839);
nand U5211 (N_5211,N_2367,N_2487);
nand U5212 (N_5212,N_4441,N_354);
or U5213 (N_5213,N_4866,N_1331);
nand U5214 (N_5214,N_1536,N_3273);
and U5215 (N_5215,N_1695,N_26);
nor U5216 (N_5216,N_2596,N_3762);
and U5217 (N_5217,N_296,N_4942);
xnor U5218 (N_5218,N_3830,N_3748);
nor U5219 (N_5219,N_1918,N_3375);
xor U5220 (N_5220,N_3129,N_2424);
nor U5221 (N_5221,N_3315,N_3997);
nor U5222 (N_5222,N_2302,N_1230);
and U5223 (N_5223,N_3000,N_3509);
and U5224 (N_5224,N_3813,N_2493);
nand U5225 (N_5225,N_4855,N_3906);
and U5226 (N_5226,N_2923,N_2427);
nor U5227 (N_5227,N_4660,N_1358);
or U5228 (N_5228,N_4889,N_2754);
or U5229 (N_5229,N_1658,N_3632);
nand U5230 (N_5230,N_3948,N_720);
nor U5231 (N_5231,N_4435,N_4312);
xnor U5232 (N_5232,N_2817,N_1744);
or U5233 (N_5233,N_1510,N_112);
and U5234 (N_5234,N_3525,N_4667);
and U5235 (N_5235,N_2268,N_8);
nor U5236 (N_5236,N_1008,N_498);
or U5237 (N_5237,N_2209,N_3362);
or U5238 (N_5238,N_4590,N_4285);
nand U5239 (N_5239,N_4552,N_507);
or U5240 (N_5240,N_2563,N_1137);
nand U5241 (N_5241,N_3926,N_2619);
or U5242 (N_5242,N_2912,N_1970);
or U5243 (N_5243,N_4573,N_1122);
nand U5244 (N_5244,N_4017,N_2622);
xnor U5245 (N_5245,N_4999,N_2146);
nor U5246 (N_5246,N_1946,N_2894);
and U5247 (N_5247,N_1934,N_1414);
nor U5248 (N_5248,N_589,N_4066);
nor U5249 (N_5249,N_12,N_1754);
or U5250 (N_5250,N_2061,N_1958);
and U5251 (N_5251,N_4720,N_3947);
nand U5252 (N_5252,N_4092,N_1608);
and U5253 (N_5253,N_1342,N_4529);
nand U5254 (N_5254,N_1873,N_4943);
nand U5255 (N_5255,N_1152,N_4257);
or U5256 (N_5256,N_1318,N_2326);
nand U5257 (N_5257,N_2078,N_2835);
nand U5258 (N_5258,N_375,N_2645);
or U5259 (N_5259,N_4994,N_3710);
nand U5260 (N_5260,N_844,N_1405);
or U5261 (N_5261,N_1181,N_1481);
or U5262 (N_5262,N_1631,N_402);
nor U5263 (N_5263,N_2707,N_3101);
nor U5264 (N_5264,N_2175,N_3970);
nand U5265 (N_5265,N_446,N_4722);
or U5266 (N_5266,N_4513,N_4246);
nand U5267 (N_5267,N_4891,N_3680);
and U5268 (N_5268,N_4753,N_3667);
nor U5269 (N_5269,N_2599,N_122);
xnor U5270 (N_5270,N_3794,N_867);
xor U5271 (N_5271,N_513,N_2819);
xnor U5272 (N_5272,N_184,N_2298);
nand U5273 (N_5273,N_3716,N_2335);
and U5274 (N_5274,N_1498,N_180);
or U5275 (N_5275,N_2568,N_923);
xor U5276 (N_5276,N_3374,N_3890);
xor U5277 (N_5277,N_521,N_4715);
and U5278 (N_5278,N_2837,N_143);
nand U5279 (N_5279,N_1712,N_430);
and U5280 (N_5280,N_678,N_68);
or U5281 (N_5281,N_2216,N_3428);
nand U5282 (N_5282,N_2350,N_2071);
and U5283 (N_5283,N_1107,N_1953);
xor U5284 (N_5284,N_4050,N_4376);
and U5285 (N_5285,N_2525,N_4291);
or U5286 (N_5286,N_658,N_3696);
and U5287 (N_5287,N_2033,N_2372);
and U5288 (N_5288,N_511,N_3371);
xor U5289 (N_5289,N_349,N_821);
xnor U5290 (N_5290,N_2520,N_2236);
xor U5291 (N_5291,N_1362,N_2199);
or U5292 (N_5292,N_3262,N_470);
nand U5293 (N_5293,N_4770,N_1549);
and U5294 (N_5294,N_3246,N_1275);
nand U5295 (N_5295,N_2558,N_1849);
nor U5296 (N_5296,N_928,N_90);
nor U5297 (N_5297,N_924,N_2287);
nor U5298 (N_5298,N_4248,N_1949);
or U5299 (N_5299,N_3471,N_3087);
and U5300 (N_5300,N_2363,N_4620);
or U5301 (N_5301,N_295,N_1905);
xor U5302 (N_5302,N_3767,N_1588);
xnor U5303 (N_5303,N_3086,N_1858);
nor U5304 (N_5304,N_2976,N_2710);
nand U5305 (N_5305,N_2984,N_4139);
nor U5306 (N_5306,N_2899,N_1735);
nand U5307 (N_5307,N_4743,N_3402);
nand U5308 (N_5308,N_1465,N_1395);
nor U5309 (N_5309,N_3764,N_1955);
nor U5310 (N_5310,N_793,N_2215);
nor U5311 (N_5311,N_4856,N_3641);
nor U5312 (N_5312,N_182,N_489);
or U5313 (N_5313,N_2387,N_1308);
nor U5314 (N_5314,N_4811,N_640);
xor U5315 (N_5315,N_4437,N_3136);
xor U5316 (N_5316,N_3450,N_2821);
nor U5317 (N_5317,N_3560,N_3230);
nand U5318 (N_5318,N_3623,N_1023);
or U5319 (N_5319,N_1150,N_92);
nand U5320 (N_5320,N_685,N_2187);
or U5321 (N_5321,N_1820,N_2704);
nor U5322 (N_5322,N_4899,N_1457);
and U5323 (N_5323,N_1581,N_963);
nor U5324 (N_5324,N_30,N_75);
nor U5325 (N_5325,N_1697,N_3009);
xnor U5326 (N_5326,N_2077,N_4102);
xnor U5327 (N_5327,N_4253,N_1114);
or U5328 (N_5328,N_1972,N_3836);
xnor U5329 (N_5329,N_2294,N_938);
xor U5330 (N_5330,N_4462,N_137);
xor U5331 (N_5331,N_2756,N_187);
xor U5332 (N_5332,N_3308,N_860);
nor U5333 (N_5333,N_684,N_516);
or U5334 (N_5334,N_2226,N_1431);
and U5335 (N_5335,N_492,N_1460);
nor U5336 (N_5336,N_120,N_2885);
or U5337 (N_5337,N_2351,N_2306);
nand U5338 (N_5338,N_881,N_1593);
nor U5339 (N_5339,N_2789,N_4272);
nor U5340 (N_5340,N_1146,N_2941);
xnor U5341 (N_5341,N_818,N_4095);
nor U5342 (N_5342,N_2065,N_3635);
xor U5343 (N_5343,N_2985,N_4813);
nor U5344 (N_5344,N_1506,N_2451);
nor U5345 (N_5345,N_3379,N_2997);
xnor U5346 (N_5346,N_4984,N_1156);
nor U5347 (N_5347,N_535,N_969);
nand U5348 (N_5348,N_2860,N_4670);
and U5349 (N_5349,N_2655,N_2004);
nor U5350 (N_5350,N_2377,N_759);
xor U5351 (N_5351,N_662,N_4518);
nand U5352 (N_5352,N_1037,N_826);
nor U5353 (N_5353,N_1430,N_2105);
xnor U5354 (N_5354,N_742,N_4864);
xor U5355 (N_5355,N_401,N_590);
and U5356 (N_5356,N_2331,N_1816);
nor U5357 (N_5357,N_443,N_3850);
nor U5358 (N_5358,N_1139,N_3994);
and U5359 (N_5359,N_361,N_2875);
nor U5360 (N_5360,N_4047,N_2549);
or U5361 (N_5361,N_3757,N_2066);
and U5362 (N_5362,N_2174,N_3507);
and U5363 (N_5363,N_4569,N_2153);
xnor U5364 (N_5364,N_4580,N_3345);
nor U5365 (N_5365,N_1924,N_506);
xor U5366 (N_5366,N_144,N_1049);
nor U5367 (N_5367,N_4407,N_3666);
xor U5368 (N_5368,N_2724,N_2257);
nor U5369 (N_5369,N_1862,N_527);
nor U5370 (N_5370,N_729,N_341);
and U5371 (N_5371,N_2253,N_55);
xnor U5372 (N_5372,N_1274,N_251);
and U5373 (N_5373,N_1912,N_4225);
nand U5374 (N_5374,N_356,N_2299);
nor U5375 (N_5375,N_4290,N_1542);
xnor U5376 (N_5376,N_2908,N_3352);
nand U5377 (N_5377,N_79,N_3232);
or U5378 (N_5378,N_2920,N_1594);
or U5379 (N_5379,N_1825,N_2644);
nor U5380 (N_5380,N_38,N_4171);
nand U5381 (N_5381,N_3529,N_4848);
nor U5382 (N_5382,N_3570,N_4965);
nand U5383 (N_5383,N_3921,N_3018);
and U5384 (N_5384,N_39,N_3594);
and U5385 (N_5385,N_2273,N_1761);
nand U5386 (N_5386,N_1855,N_4609);
or U5387 (N_5387,N_4795,N_3832);
nand U5388 (N_5388,N_2662,N_1326);
xor U5389 (N_5389,N_701,N_4834);
nor U5390 (N_5390,N_176,N_3460);
and U5391 (N_5391,N_3925,N_32);
and U5392 (N_5392,N_4551,N_424);
or U5393 (N_5393,N_4003,N_799);
nor U5394 (N_5394,N_3883,N_3543);
nor U5395 (N_5395,N_989,N_3911);
nand U5396 (N_5396,N_249,N_1638);
and U5397 (N_5397,N_4547,N_2715);
and U5398 (N_5398,N_4324,N_988);
or U5399 (N_5399,N_3211,N_871);
nand U5400 (N_5400,N_1672,N_3945);
xnor U5401 (N_5401,N_3404,N_1680);
nand U5402 (N_5402,N_1904,N_4915);
or U5403 (N_5403,N_816,N_4657);
nand U5404 (N_5404,N_4845,N_2039);
nand U5405 (N_5405,N_3039,N_4414);
nand U5406 (N_5406,N_2531,N_2385);
or U5407 (N_5407,N_4621,N_1348);
nand U5408 (N_5408,N_3302,N_914);
nor U5409 (N_5409,N_2263,N_2936);
or U5410 (N_5410,N_1208,N_3376);
nand U5411 (N_5411,N_4390,N_1528);
nor U5412 (N_5412,N_2364,N_746);
xor U5413 (N_5413,N_4566,N_1264);
nand U5414 (N_5414,N_297,N_328);
xnor U5415 (N_5415,N_1847,N_4639);
and U5416 (N_5416,N_4939,N_536);
xnor U5417 (N_5417,N_999,N_3319);
or U5418 (N_5418,N_668,N_1798);
nor U5419 (N_5419,N_1526,N_1284);
and U5420 (N_5420,N_1368,N_743);
or U5421 (N_5421,N_4387,N_565);
xnor U5422 (N_5422,N_304,N_3733);
nor U5423 (N_5423,N_2416,N_9);
nand U5424 (N_5424,N_4106,N_28);
and U5425 (N_5425,N_1184,N_1673);
or U5426 (N_5426,N_2902,N_2853);
nand U5427 (N_5427,N_1961,N_3897);
xnor U5428 (N_5428,N_805,N_4824);
or U5429 (N_5429,N_2689,N_162);
xnor U5430 (N_5430,N_287,N_3090);
and U5431 (N_5431,N_4732,N_1930);
xnor U5432 (N_5432,N_3597,N_707);
nand U5433 (N_5433,N_4966,N_3739);
and U5434 (N_5434,N_4415,N_145);
nor U5435 (N_5435,N_514,N_3606);
xor U5436 (N_5436,N_44,N_4704);
and U5437 (N_5437,N_562,N_1777);
or U5438 (N_5438,N_437,N_1810);
and U5439 (N_5439,N_2987,N_271);
and U5440 (N_5440,N_798,N_4197);
xor U5441 (N_5441,N_902,N_2966);
and U5442 (N_5442,N_215,N_1917);
and U5443 (N_5443,N_3637,N_3476);
nor U5444 (N_5444,N_1271,N_1385);
xnor U5445 (N_5445,N_298,N_1094);
xor U5446 (N_5446,N_1117,N_155);
or U5447 (N_5447,N_1689,N_4534);
nand U5448 (N_5448,N_1407,N_66);
nor U5449 (N_5449,N_3718,N_1852);
nor U5450 (N_5450,N_4306,N_4164);
and U5451 (N_5451,N_4427,N_1908);
nand U5452 (N_5452,N_2940,N_2011);
xor U5453 (N_5453,N_1714,N_689);
nor U5454 (N_5454,N_153,N_283);
nor U5455 (N_5455,N_4389,N_3477);
or U5456 (N_5456,N_2606,N_558);
or U5457 (N_5457,N_231,N_986);
nor U5458 (N_5458,N_2733,N_3453);
xor U5459 (N_5459,N_755,N_2109);
or U5460 (N_5460,N_1990,N_88);
nand U5461 (N_5461,N_54,N_931);
nor U5462 (N_5462,N_4788,N_3027);
nand U5463 (N_5463,N_2646,N_2477);
xnor U5464 (N_5464,N_898,N_433);
or U5465 (N_5465,N_4614,N_4701);
and U5466 (N_5466,N_2652,N_2613);
and U5467 (N_5467,N_4124,N_1109);
or U5468 (N_5468,N_1487,N_4623);
nor U5469 (N_5469,N_4433,N_2083);
nand U5470 (N_5470,N_2583,N_2573);
nor U5471 (N_5471,N_450,N_2827);
and U5472 (N_5472,N_2629,N_3892);
xnor U5473 (N_5473,N_2266,N_2423);
and U5474 (N_5474,N_655,N_2535);
and U5475 (N_5475,N_3709,N_3998);
xor U5476 (N_5476,N_2876,N_1586);
xnor U5477 (N_5477,N_1383,N_499);
nand U5478 (N_5478,N_2031,N_2388);
xnor U5479 (N_5479,N_1900,N_580);
nand U5480 (N_5480,N_585,N_2591);
nor U5481 (N_5481,N_4490,N_2228);
xor U5482 (N_5482,N_3530,N_1288);
and U5483 (N_5483,N_2571,N_3126);
nand U5484 (N_5484,N_1179,N_4244);
nor U5485 (N_5485,N_3834,N_4951);
nor U5486 (N_5486,N_4467,N_554);
xnor U5487 (N_5487,N_1202,N_3200);
nor U5488 (N_5488,N_4251,N_3728);
or U5489 (N_5489,N_2589,N_1730);
or U5490 (N_5490,N_4183,N_4029);
nor U5491 (N_5491,N_1163,N_1717);
and U5492 (N_5492,N_4077,N_3551);
nand U5493 (N_5493,N_10,N_1083);
and U5494 (N_5494,N_4906,N_3557);
nand U5495 (N_5495,N_1445,N_1525);
nor U5496 (N_5496,N_501,N_4198);
or U5497 (N_5497,N_3451,N_1618);
or U5498 (N_5498,N_4071,N_2974);
or U5499 (N_5499,N_4509,N_4969);
or U5500 (N_5500,N_3829,N_292);
xor U5501 (N_5501,N_487,N_3343);
and U5502 (N_5502,N_957,N_4252);
nand U5503 (N_5503,N_2594,N_3111);
or U5504 (N_5504,N_2909,N_432);
nand U5505 (N_5505,N_4697,N_4649);
nand U5506 (N_5506,N_1940,N_2556);
or U5507 (N_5507,N_3942,N_2204);
and U5508 (N_5508,N_4946,N_264);
and U5509 (N_5509,N_2405,N_158);
xnor U5510 (N_5510,N_2991,N_626);
xnor U5511 (N_5511,N_1423,N_4249);
nor U5512 (N_5512,N_808,N_4035);
nor U5513 (N_5513,N_802,N_2171);
nand U5514 (N_5514,N_900,N_3595);
nand U5515 (N_5515,N_2210,N_1884);
and U5516 (N_5516,N_1016,N_4874);
xor U5517 (N_5517,N_4671,N_708);
nand U5518 (N_5518,N_1299,N_486);
and U5519 (N_5519,N_4195,N_2284);
or U5520 (N_5520,N_3974,N_4494);
and U5521 (N_5521,N_728,N_4964);
nor U5522 (N_5522,N_4216,N_35);
or U5523 (N_5523,N_2258,N_4468);
xor U5524 (N_5524,N_3373,N_2037);
nor U5525 (N_5525,N_2489,N_2453);
xor U5526 (N_5526,N_1962,N_220);
or U5527 (N_5527,N_1982,N_4936);
and U5528 (N_5528,N_3270,N_56);
and U5529 (N_5529,N_4430,N_1644);
nor U5530 (N_5530,N_1760,N_116);
or U5531 (N_5531,N_1543,N_2013);
and U5532 (N_5532,N_4,N_936);
nand U5533 (N_5533,N_262,N_1876);
xnor U5534 (N_5534,N_4525,N_3380);
and U5535 (N_5535,N_2392,N_3912);
nor U5536 (N_5536,N_3386,N_3123);
and U5537 (N_5537,N_3568,N_1684);
or U5538 (N_5538,N_1729,N_2120);
nand U5539 (N_5539,N_1044,N_3628);
and U5540 (N_5540,N_1329,N_3265);
xor U5541 (N_5541,N_2484,N_3639);
or U5542 (N_5542,N_3258,N_2519);
nand U5543 (N_5543,N_2744,N_1653);
nor U5544 (N_5544,N_2900,N_273);
or U5545 (N_5545,N_2296,N_875);
and U5546 (N_5546,N_2683,N_628);
xor U5547 (N_5547,N_4661,N_2816);
nor U5548 (N_5548,N_4258,N_2534);
nand U5549 (N_5549,N_2475,N_175);
or U5550 (N_5550,N_3745,N_586);
nand U5551 (N_5551,N_515,N_1377);
nand U5552 (N_5552,N_2108,N_1111);
nand U5553 (N_5553,N_168,N_916);
or U5554 (N_5554,N_169,N_1694);
nand U5555 (N_5555,N_4113,N_1601);
nand U5556 (N_5556,N_3293,N_4783);
or U5557 (N_5557,N_3318,N_2721);
nor U5558 (N_5558,N_2581,N_1315);
nand U5559 (N_5559,N_642,N_2935);
nand U5560 (N_5560,N_1713,N_80);
nand U5561 (N_5561,N_4776,N_2205);
xor U5562 (N_5562,N_1102,N_1926);
or U5563 (N_5563,N_4893,N_926);
and U5564 (N_5564,N_2554,N_2132);
xor U5565 (N_5565,N_4072,N_2305);
nand U5566 (N_5566,N_346,N_2530);
and U5567 (N_5567,N_2545,N_3225);
and U5568 (N_5568,N_3403,N_3181);
and U5569 (N_5569,N_1563,N_1373);
nand U5570 (N_5570,N_2064,N_4125);
or U5571 (N_5571,N_4083,N_3975);
or U5572 (N_5572,N_4097,N_2942);
nand U5573 (N_5573,N_229,N_1939);
or U5574 (N_5574,N_243,N_3995);
nand U5575 (N_5575,N_2124,N_2810);
xnor U5576 (N_5576,N_4726,N_1389);
or U5577 (N_5577,N_966,N_1708);
and U5578 (N_5578,N_4592,N_1865);
or U5579 (N_5579,N_3938,N_3100);
and U5580 (N_5580,N_1468,N_4761);
and U5581 (N_5581,N_3775,N_2677);
or U5582 (N_5582,N_1513,N_1133);
and U5583 (N_5583,N_2457,N_3383);
or U5584 (N_5584,N_3022,N_3627);
nand U5585 (N_5585,N_4712,N_3548);
or U5586 (N_5586,N_2524,N_1492);
nand U5587 (N_5587,N_4618,N_4281);
and U5588 (N_5588,N_3424,N_2667);
xor U5589 (N_5589,N_602,N_481);
xor U5590 (N_5590,N_2533,N_3492);
nand U5591 (N_5591,N_1080,N_1799);
nand U5592 (N_5592,N_1787,N_3889);
and U5593 (N_5593,N_18,N_2604);
nand U5594 (N_5594,N_2503,N_1570);
nand U5595 (N_5595,N_1300,N_4033);
or U5596 (N_5596,N_1317,N_1145);
nand U5597 (N_5597,N_1296,N_964);
nand U5598 (N_5598,N_224,N_2823);
nand U5599 (N_5599,N_2802,N_3005);
nor U5600 (N_5600,N_1266,N_1629);
and U5601 (N_5601,N_1471,N_1025);
and U5602 (N_5602,N_1305,N_3746);
or U5603 (N_5603,N_597,N_3905);
nand U5604 (N_5604,N_1566,N_43);
and U5605 (N_5605,N_2129,N_2763);
xor U5606 (N_5606,N_4527,N_939);
nor U5607 (N_5607,N_1161,N_4819);
nor U5608 (N_5608,N_982,N_3705);
or U5609 (N_5609,N_873,N_1944);
nor U5610 (N_5610,N_4413,N_3210);
nor U5611 (N_5611,N_1535,N_4060);
or U5612 (N_5612,N_2274,N_576);
and U5613 (N_5613,N_3068,N_330);
nor U5614 (N_5614,N_4968,N_4146);
and U5615 (N_5615,N_252,N_303);
or U5616 (N_5616,N_4179,N_1157);
or U5617 (N_5617,N_3239,N_4163);
nand U5618 (N_5618,N_4374,N_452);
or U5619 (N_5619,N_2022,N_4320);
and U5620 (N_5620,N_4184,N_3184);
nor U5621 (N_5621,N_2560,N_3359);
xor U5622 (N_5622,N_4656,N_850);
and U5623 (N_5623,N_2851,N_1011);
xnor U5624 (N_5624,N_191,N_2468);
nor U5625 (N_5625,N_4967,N_4807);
nor U5626 (N_5626,N_1577,N_2088);
nand U5627 (N_5627,N_427,N_3964);
or U5628 (N_5628,N_234,N_4107);
and U5629 (N_5629,N_508,N_1870);
nand U5630 (N_5630,N_3853,N_2264);
nor U5631 (N_5631,N_4166,N_766);
and U5632 (N_5632,N_2251,N_4325);
and U5633 (N_5633,N_2207,N_3042);
xor U5634 (N_5634,N_1683,N_3268);
nor U5635 (N_5635,N_3967,N_2651);
and U5636 (N_5636,N_2764,N_396);
xor U5637 (N_5637,N_2543,N_366);
nand U5638 (N_5638,N_6,N_2189);
xnor U5639 (N_5639,N_3684,N_409);
and U5640 (N_5640,N_734,N_2675);
or U5641 (N_5641,N_3006,N_1916);
nor U5642 (N_5642,N_1194,N_3336);
nand U5643 (N_5643,N_2417,N_3245);
and U5644 (N_5644,N_136,N_2232);
nor U5645 (N_5645,N_1214,N_4181);
and U5646 (N_5646,N_3828,N_2926);
or U5647 (N_5647,N_2521,N_4189);
xnor U5648 (N_5648,N_3808,N_4010);
nor U5649 (N_5649,N_164,N_533);
nor U5650 (N_5650,N_2701,N_3556);
nand U5651 (N_5651,N_3001,N_3290);
and U5652 (N_5652,N_2532,N_104);
xnor U5653 (N_5653,N_1088,N_3074);
nand U5654 (N_5654,N_1670,N_435);
and U5655 (N_5655,N_1428,N_3452);
and U5656 (N_5656,N_1106,N_2219);
xor U5657 (N_5657,N_2818,N_3390);
nor U5658 (N_5658,N_2297,N_1796);
and U5659 (N_5659,N_605,N_1746);
xor U5660 (N_5660,N_4648,N_2930);
nand U5661 (N_5661,N_4226,N_270);
and U5662 (N_5662,N_3099,N_2133);
and U5663 (N_5663,N_1518,N_3903);
nor U5664 (N_5664,N_4591,N_2098);
or U5665 (N_5665,N_389,N_4067);
nor U5666 (N_5666,N_210,N_1914);
nor U5667 (N_5667,N_4313,N_3822);
xnor U5668 (N_5668,N_2538,N_4283);
nor U5669 (N_5669,N_4918,N_2443);
nand U5670 (N_5670,N_1301,N_4075);
nand U5671 (N_5671,N_4519,N_570);
xnor U5672 (N_5672,N_1923,N_2542);
nand U5673 (N_5673,N_199,N_4062);
nand U5674 (N_5674,N_3949,N_1656);
and U5675 (N_5675,N_1424,N_2390);
nor U5676 (N_5676,N_4960,N_559);
and U5677 (N_5677,N_1056,N_2505);
and U5678 (N_5678,N_2579,N_3687);
xnor U5679 (N_5679,N_4710,N_3493);
and U5680 (N_5680,N_845,N_998);
or U5681 (N_5681,N_4079,N_4109);
and U5682 (N_5682,N_3941,N_1606);
or U5683 (N_5683,N_1806,N_2114);
xnor U5684 (N_5684,N_318,N_1867);
nor U5685 (N_5685,N_3357,N_1845);
xnor U5686 (N_5686,N_2806,N_1285);
or U5687 (N_5687,N_4108,N_3172);
and U5688 (N_5688,N_4363,N_3989);
nand U5689 (N_5689,N_4935,N_4267);
xnor U5690 (N_5690,N_42,N_2905);
and U5691 (N_5691,N_2621,N_1257);
and U5692 (N_5692,N_3197,N_17);
nand U5693 (N_5693,N_4749,N_3772);
or U5694 (N_5694,N_3183,N_4175);
nor U5695 (N_5695,N_2256,N_3057);
and U5696 (N_5696,N_4400,N_2127);
xor U5697 (N_5697,N_3405,N_3962);
xor U5698 (N_5698,N_2735,N_637);
xor U5699 (N_5699,N_3769,N_3052);
nor U5700 (N_5700,N_3940,N_2044);
nor U5701 (N_5701,N_2408,N_2168);
xor U5702 (N_5702,N_4944,N_1120);
or U5703 (N_5703,N_2537,N_3377);
xor U5704 (N_5704,N_384,N_3089);
and U5705 (N_5705,N_3481,N_3770);
and U5706 (N_5706,N_956,N_372);
nand U5707 (N_5707,N_2485,N_418);
nand U5708 (N_5708,N_2670,N_3138);
or U5709 (N_5709,N_4814,N_2144);
and U5710 (N_5710,N_3706,N_4584);
or U5711 (N_5711,N_1352,N_2780);
xor U5712 (N_5712,N_3464,N_2142);
and U5713 (N_5713,N_71,N_3151);
xor U5714 (N_5714,N_3731,N_4919);
xnor U5715 (N_5715,N_1124,N_649);
nand U5716 (N_5716,N_2290,N_1749);
xor U5717 (N_5717,N_2771,N_1576);
nor U5718 (N_5718,N_2354,N_3721);
nand U5719 (N_5719,N_3037,N_4589);
and U5720 (N_5720,N_3264,N_1623);
nor U5721 (N_5721,N_4222,N_546);
and U5722 (N_5722,N_67,N_4703);
or U5723 (N_5723,N_3935,N_503);
nor U5724 (N_5724,N_2466,N_528);
nand U5725 (N_5725,N_417,N_1119);
xnor U5726 (N_5726,N_1255,N_2901);
nand U5727 (N_5727,N_1063,N_4831);
nor U5728 (N_5728,N_3192,N_2518);
or U5729 (N_5729,N_4064,N_3292);
xnor U5730 (N_5730,N_4168,N_103);
or U5731 (N_5731,N_289,N_4068);
or U5732 (N_5732,N_3602,N_4296);
or U5733 (N_5733,N_3854,N_1721);
or U5734 (N_5734,N_3864,N_4937);
nand U5735 (N_5735,N_748,N_4817);
nand U5736 (N_5736,N_4739,N_2781);
or U5737 (N_5737,N_4535,N_4924);
xnor U5738 (N_5738,N_185,N_2431);
xnor U5739 (N_5739,N_1980,N_3426);
nand U5740 (N_5740,N_2973,N_258);
nor U5741 (N_5741,N_2470,N_3702);
or U5742 (N_5742,N_2711,N_3839);
and U5743 (N_5743,N_3331,N_4276);
and U5744 (N_5744,N_2725,N_1743);
nor U5745 (N_5745,N_3486,N_4851);
or U5746 (N_5746,N_1533,N_2202);
xor U5747 (N_5747,N_753,N_468);
xor U5748 (N_5748,N_4913,N_4578);
nor U5749 (N_5749,N_1440,N_1007);
nor U5750 (N_5750,N_712,N_2002);
nand U5751 (N_5751,N_1928,N_667);
nand U5752 (N_5752,N_4112,N_946);
nand U5753 (N_5753,N_1527,N_440);
nand U5754 (N_5754,N_2799,N_1344);
or U5755 (N_5755,N_3954,N_4912);
nor U5756 (N_5756,N_2319,N_4897);
xor U5757 (N_5757,N_2638,N_2191);
or U5758 (N_5758,N_4448,N_3024);
or U5759 (N_5759,N_373,N_2369);
nor U5760 (N_5760,N_690,N_2380);
nor U5761 (N_5761,N_1322,N_2448);
or U5762 (N_5762,N_4887,N_2564);
nor U5763 (N_5763,N_414,N_2868);
and U5764 (N_5764,N_2867,N_1391);
nand U5765 (N_5765,N_4130,N_4221);
nor U5766 (N_5766,N_2865,N_1821);
nand U5767 (N_5767,N_2691,N_237);
xnor U5768 (N_5768,N_4988,N_3521);
and U5769 (N_5769,N_2115,N_4344);
nor U5770 (N_5770,N_2320,N_4330);
and U5771 (N_5771,N_852,N_2450);
or U5772 (N_5772,N_1863,N_3051);
and U5773 (N_5773,N_131,N_2288);
or U5774 (N_5774,N_1144,N_189);
nor U5775 (N_5775,N_1261,N_4521);
nor U5776 (N_5776,N_467,N_2397);
xor U5777 (N_5777,N_541,N_1493);
and U5778 (N_5778,N_4403,N_286);
xor U5779 (N_5779,N_4892,N_3584);
nor U5780 (N_5780,N_2110,N_242);
or U5781 (N_5781,N_1355,N_1782);
nand U5782 (N_5782,N_4745,N_3306);
nand U5783 (N_5783,N_955,N_1603);
nor U5784 (N_5784,N_3332,N_386);
nand U5785 (N_5785,N_1886,N_392);
nor U5786 (N_5786,N_2986,N_4907);
and U5787 (N_5787,N_3815,N_727);
and U5788 (N_5788,N_2988,N_2016);
xor U5789 (N_5789,N_474,N_4635);
or U5790 (N_5790,N_2893,N_2947);
nand U5791 (N_5791,N_4804,N_2544);
nand U5792 (N_5792,N_4089,N_3939);
nor U5793 (N_5793,N_2248,N_4698);
and U5794 (N_5794,N_4150,N_828);
or U5795 (N_5795,N_1134,N_4926);
xor U5796 (N_5796,N_2785,N_3812);
or U5797 (N_5797,N_2244,N_2042);
nor U5798 (N_5798,N_2325,N_3170);
or U5799 (N_5799,N_1341,N_3870);
or U5800 (N_5800,N_1010,N_1968);
xor U5801 (N_5801,N_523,N_3185);
nor U5802 (N_5802,N_744,N_4122);
xor U5803 (N_5803,N_2745,N_3630);
nand U5804 (N_5804,N_2309,N_3683);
or U5805 (N_5805,N_4013,N_1203);
or U5806 (N_5806,N_473,N_269);
or U5807 (N_5807,N_3809,N_3061);
nor U5808 (N_5808,N_617,N_4921);
xnor U5809 (N_5809,N_420,N_899);
nor U5810 (N_5810,N_3987,N_2051);
nand U5811 (N_5811,N_3400,N_3653);
or U5812 (N_5812,N_2800,N_485);
and U5813 (N_5813,N_3780,N_3801);
or U5814 (N_5814,N_3176,N_390);
and U5815 (N_5815,N_1218,N_360);
nor U5816 (N_5816,N_1100,N_621);
or U5817 (N_5817,N_4972,N_1545);
nand U5818 (N_5818,N_3247,N_1198);
xor U5819 (N_5819,N_4998,N_3803);
and U5820 (N_5820,N_1966,N_3790);
nor U5821 (N_5821,N_3283,N_587);
and U5822 (N_5822,N_4615,N_434);
or U5823 (N_5823,N_2483,N_663);
xor U5824 (N_5824,N_851,N_3563);
or U5825 (N_5825,N_4707,N_4875);
nand U5826 (N_5826,N_3013,N_3021);
or U5827 (N_5827,N_4847,N_1408);
and U5828 (N_5828,N_3566,N_3473);
nor U5829 (N_5829,N_4001,N_4345);
nand U5830 (N_5830,N_3725,N_4261);
nand U5831 (N_5831,N_1764,N_1851);
nand U5832 (N_5832,N_1602,N_1532);
xor U5833 (N_5833,N_1677,N_3820);
nor U5834 (N_5834,N_740,N_2255);
or U5835 (N_5835,N_37,N_4898);
nor U5836 (N_5836,N_788,N_1985);
or U5837 (N_5837,N_2093,N_3025);
nor U5838 (N_5838,N_2585,N_869);
or U5839 (N_5839,N_2073,N_906);
nand U5840 (N_5840,N_4452,N_3774);
xnor U5841 (N_5841,N_4806,N_1840);
nand U5842 (N_5842,N_1273,N_2000);
nand U5843 (N_5843,N_1135,N_718);
xor U5844 (N_5844,N_48,N_1148);
xor U5845 (N_5845,N_4602,N_4461);
xnor U5846 (N_5846,N_288,N_1068);
and U5847 (N_5847,N_1164,N_735);
and U5848 (N_5848,N_94,N_1197);
xnor U5849 (N_5849,N_1473,N_3092);
nand U5850 (N_5850,N_2318,N_2762);
nand U5851 (N_5851,N_3455,N_4134);
and U5852 (N_5852,N_1382,N_616);
nand U5853 (N_5853,N_3895,N_3048);
or U5854 (N_5854,N_299,N_997);
and U5855 (N_5855,N_3807,N_4708);
nor U5856 (N_5856,N_172,N_16);
xor U5857 (N_5857,N_4205,N_2308);
xor U5858 (N_5858,N_3694,N_878);
nor U5859 (N_5859,N_4310,N_4869);
xor U5860 (N_5860,N_2874,N_4420);
xnor U5861 (N_5861,N_385,N_2025);
nor U5862 (N_5862,N_4818,N_722);
nor U5863 (N_5863,N_1219,N_4916);
or U5864 (N_5864,N_4242,N_556);
nor U5865 (N_5865,N_4372,N_4786);
nor U5866 (N_5866,N_2739,N_20);
nor U5867 (N_5867,N_3642,N_466);
nor U5868 (N_5868,N_1559,N_688);
xor U5869 (N_5869,N_2280,N_2428);
and U5870 (N_5870,N_3439,N_3861);
and U5871 (N_5871,N_1771,N_190);
and U5872 (N_5872,N_3558,N_3960);
xnor U5873 (N_5873,N_2310,N_3130);
or U5874 (N_5874,N_4880,N_245);
or U5875 (N_5875,N_3722,N_33);
or U5876 (N_5876,N_2162,N_932);
xor U5877 (N_5877,N_1828,N_3294);
and U5878 (N_5878,N_1872,N_3648);
nor U5879 (N_5879,N_1829,N_1790);
and U5880 (N_5880,N_2963,N_1732);
or U5881 (N_5881,N_1013,N_4843);
and U5882 (N_5882,N_3213,N_1458);
nor U5883 (N_5883,N_623,N_886);
nand U5884 (N_5884,N_4365,N_3387);
nand U5885 (N_5885,N_3016,N_3805);
and U5886 (N_5886,N_2494,N_174);
and U5887 (N_5887,N_4133,N_4332);
nand U5888 (N_5888,N_4512,N_4114);
and U5889 (N_5889,N_4317,N_1974);
nor U5890 (N_5890,N_1668,N_2620);
and U5891 (N_5891,N_1544,N_4920);
nor U5892 (N_5892,N_323,N_1279);
xnor U5893 (N_5893,N_2186,N_4974);
nand U5894 (N_5894,N_469,N_1172);
xor U5895 (N_5895,N_3083,N_2131);
and U5896 (N_5896,N_3433,N_1598);
xnor U5897 (N_5897,N_159,N_1036);
nor U5898 (N_5898,N_3478,N_84);
nand U5899 (N_5899,N_2081,N_1042);
xor U5900 (N_5900,N_3715,N_4514);
or U5901 (N_5901,N_3075,N_441);
nor U5902 (N_5902,N_2316,N_1328);
nor U5903 (N_5903,N_4785,N_3346);
xor U5904 (N_5904,N_911,N_314);
nand U5905 (N_5905,N_933,N_1050);
or U5906 (N_5906,N_4503,N_542);
xor U5907 (N_5907,N_2289,N_1741);
or U5908 (N_5908,N_3561,N_1875);
nor U5909 (N_5909,N_3096,N_2459);
and U5910 (N_5910,N_2811,N_1446);
nor U5911 (N_5911,N_313,N_4212);
and U5912 (N_5912,N_1758,N_436);
nor U5913 (N_5913,N_4260,N_4245);
or U5914 (N_5914,N_4837,N_813);
nor U5915 (N_5915,N_4676,N_477);
or U5916 (N_5916,N_3631,N_7);
xnor U5917 (N_5917,N_4662,N_3157);
xor U5918 (N_5918,N_765,N_786);
xnor U5919 (N_5919,N_3105,N_2658);
or U5920 (N_5920,N_4129,N_78);
nor U5921 (N_5921,N_331,N_2660);
and U5922 (N_5922,N_45,N_671);
or U5923 (N_5923,N_3040,N_2307);
nand U5924 (N_5924,N_2176,N_4279);
or U5925 (N_5925,N_1323,N_646);
or U5926 (N_5926,N_4504,N_3417);
and U5927 (N_5927,N_1878,N_3115);
or U5928 (N_5928,N_2743,N_4809);
nand U5929 (N_5929,N_1937,N_1705);
or U5930 (N_5930,N_670,N_4397);
and U5931 (N_5931,N_4793,N_3978);
nand U5932 (N_5932,N_4978,N_4696);
nand U5933 (N_5933,N_285,N_60);
nor U5934 (N_5934,N_2587,N_913);
xnor U5935 (N_5935,N_2999,N_3104);
nand U5936 (N_5936,N_2507,N_2425);
nand U5937 (N_5937,N_497,N_4668);
nor U5938 (N_5938,N_3855,N_4219);
nor U5939 (N_5939,N_2616,N_1217);
or U5940 (N_5940,N_2046,N_3881);
nand U5941 (N_5941,N_863,N_4632);
and U5942 (N_5942,N_3884,N_4187);
or U5943 (N_5943,N_832,N_3432);
or U5944 (N_5944,N_3155,N_1349);
and U5945 (N_5945,N_991,N_3131);
or U5946 (N_5946,N_3064,N_2378);
or U5947 (N_5947,N_3041,N_4741);
nand U5948 (N_5948,N_4797,N_4438);
nor U5949 (N_5949,N_807,N_4466);
nor U5950 (N_5950,N_1584,N_4019);
xnor U5951 (N_5951,N_1243,N_1232);
and U5952 (N_5952,N_4729,N_1932);
and U5953 (N_5953,N_615,N_3145);
xor U5954 (N_5954,N_3888,N_2855);
nor U5955 (N_5955,N_3340,N_552);
xor U5956 (N_5956,N_2846,N_2026);
and U5957 (N_5957,N_3849,N_1571);
and U5958 (N_5958,N_1979,N_4160);
nor U5959 (N_5959,N_4439,N_1943);
nand U5960 (N_5960,N_3327,N_1084);
nand U5961 (N_5961,N_2808,N_4501);
nor U5962 (N_5962,N_3982,N_944);
and U5963 (N_5963,N_3920,N_4331);
xnor U5964 (N_5964,N_3285,N_971);
and U5965 (N_5965,N_4391,N_4091);
nand U5966 (N_5966,N_3845,N_2626);
nand U5967 (N_5967,N_217,N_3827);
xor U5968 (N_5968,N_2797,N_3878);
or U5969 (N_5969,N_4949,N_774);
and U5970 (N_5970,N_4032,N_1426);
xor U5971 (N_5971,N_4057,N_2370);
or U5972 (N_5972,N_4616,N_4568);
and U5973 (N_5973,N_1248,N_4540);
nor U5974 (N_5974,N_4901,N_2769);
xor U5975 (N_5975,N_1000,N_1268);
and U5976 (N_5976,N_980,N_3943);
nor U5977 (N_5977,N_4208,N_4735);
nand U5978 (N_5978,N_2444,N_3799);
or U5979 (N_5979,N_3103,N_1553);
or U5980 (N_5980,N_416,N_3044);
nand U5981 (N_5981,N_3147,N_4434);
nor U5982 (N_5982,N_603,N_2446);
nand U5983 (N_5983,N_529,N_1534);
nor U5984 (N_5984,N_3863,N_412);
or U5985 (N_5985,N_3531,N_238);
nor U5986 (N_5986,N_650,N_2595);
nor U5987 (N_5987,N_3382,N_3071);
xnor U5988 (N_5988,N_2281,N_4952);
or U5989 (N_5989,N_618,N_495);
nor U5990 (N_5990,N_1736,N_588);
xnor U5991 (N_5991,N_4595,N_208);
and U5992 (N_5992,N_1020,N_1850);
or U5993 (N_5993,N_3655,N_896);
or U5994 (N_5994,N_170,N_4480);
xnor U5995 (N_5995,N_1277,N_2482);
xnor U5996 (N_5996,N_1515,N_1201);
xnor U5997 (N_5997,N_429,N_2182);
and U5998 (N_5998,N_2134,N_1538);
nand U5999 (N_5999,N_3466,N_3786);
nor U6000 (N_6000,N_2731,N_3516);
xnor U6001 (N_6001,N_2282,N_1614);
nor U6002 (N_6002,N_2030,N_4883);
xor U6003 (N_6003,N_1834,N_152);
nand U6004 (N_6004,N_2035,N_3615);
nor U6005 (N_6005,N_1225,N_3669);
nand U6006 (N_6006,N_2211,N_4694);
nand U6007 (N_6007,N_3779,N_4379);
nand U6008 (N_6008,N_2895,N_2147);
nand U6009 (N_6009,N_4309,N_1919);
nand U6010 (N_6010,N_1483,N_479);
and U6011 (N_6011,N_673,N_2714);
and U6012 (N_6012,N_225,N_2382);
nor U6013 (N_6013,N_3711,N_4475);
nand U6014 (N_6014,N_4254,N_4586);
xor U6015 (N_6015,N_4182,N_2332);
xor U6016 (N_6016,N_4459,N_4059);
nor U6017 (N_6017,N_4489,N_3510);
or U6018 (N_6018,N_1997,N_1354);
nor U6019 (N_6019,N_25,N_1822);
nand U6020 (N_6020,N_1973,N_1171);
and U6021 (N_6021,N_1501,N_4853);
and U6022 (N_6022,N_2514,N_1808);
xor U6023 (N_6023,N_3030,N_4233);
xor U6024 (N_6024,N_894,N_2139);
xnor U6025 (N_6025,N_4911,N_3250);
nand U6026 (N_6026,N_19,N_3795);
or U6027 (N_6027,N_3234,N_1967);
nor U6028 (N_6028,N_648,N_1321);
and U6029 (N_6029,N_4597,N_2934);
and U6030 (N_6030,N_1903,N_891);
xnor U6031 (N_6031,N_194,N_567);
xnor U6032 (N_6032,N_1938,N_3065);
and U6033 (N_6033,N_1192,N_1604);
xnor U6034 (N_6034,N_3399,N_3260);
or U6035 (N_6035,N_2359,N_1592);
nand U6036 (N_6036,N_3575,N_3593);
nor U6037 (N_6037,N_1703,N_4128);
or U6038 (N_6038,N_4799,N_4037);
nand U6039 (N_6039,N_1902,N_4672);
nor U6040 (N_6040,N_50,N_2352);
nor U6041 (N_6041,N_995,N_1560);
or U6042 (N_6042,N_683,N_3301);
or U6043 (N_6043,N_3462,N_4255);
and U6044 (N_6044,N_1753,N_4265);
xor U6045 (N_6045,N_1964,N_1089);
or U6046 (N_6046,N_1607,N_4178);
or U6047 (N_6047,N_1253,N_611);
xor U6048 (N_6048,N_2249,N_2041);
and U6049 (N_6049,N_4411,N_1051);
nor U6050 (N_6050,N_3053,N_2590);
nor U6051 (N_6051,N_3366,N_4061);
or U6052 (N_6052,N_3406,N_2850);
nor U6053 (N_6053,N_1314,N_4633);
xor U6054 (N_6054,N_4931,N_151);
xnor U6055 (N_6055,N_226,N_1794);
nand U6056 (N_6056,N_415,N_1079);
and U6057 (N_6057,N_3724,N_3553);
nand U6058 (N_6058,N_2541,N_3216);
nor U6059 (N_6059,N_4792,N_3188);
or U6060 (N_6060,N_3309,N_140);
xnor U6061 (N_6061,N_4177,N_2160);
nor U6062 (N_6062,N_779,N_2238);
or U6063 (N_6063,N_2155,N_4815);
nand U6064 (N_6064,N_4750,N_4894);
nand U6065 (N_6065,N_4247,N_1627);
and U6066 (N_6066,N_3806,N_4823);
or U6067 (N_6067,N_2055,N_439);
or U6068 (N_6068,N_368,N_4323);
or U6069 (N_6069,N_1578,N_2338);
or U6070 (N_6070,N_3656,N_1960);
and U6071 (N_6071,N_4930,N_2557);
and U6072 (N_6072,N_3480,N_519);
or U6073 (N_6073,N_448,N_2887);
xor U6074 (N_6074,N_941,N_2028);
and U6075 (N_6075,N_1427,N_1149);
and U6076 (N_6076,N_1661,N_1463);
nand U6077 (N_6077,N_4541,N_2791);
xor U6078 (N_6078,N_1131,N_347);
xnor U6079 (N_6079,N_4980,N_1679);
xor U6080 (N_6080,N_3166,N_3852);
or U6081 (N_6081,N_827,N_1421);
or U6082 (N_6082,N_3528,N_3326);
or U6083 (N_6083,N_3116,N_4399);
or U6084 (N_6084,N_951,N_2983);
nand U6085 (N_6085,N_2009,N_2669);
or U6086 (N_6086,N_3054,N_1241);
nor U6087 (N_6087,N_1945,N_3407);
and U6088 (N_6088,N_815,N_201);
nor U6089 (N_6089,N_2285,N_2032);
or U6090 (N_6090,N_142,N_3017);
xor U6091 (N_6091,N_3599,N_2478);
and U6092 (N_6092,N_1868,N_1877);
nand U6093 (N_6093,N_3999,N_2410);
and U6094 (N_6094,N_4300,N_1126);
xor U6095 (N_6095,N_1409,N_1999);
nand U6096 (N_6096,N_4368,N_1196);
xnor U6097 (N_6097,N_4954,N_3689);
or U6098 (N_6098,N_1698,N_195);
and U6099 (N_6099,N_977,N_659);
or U6100 (N_6100,N_3334,N_1880);
xor U6101 (N_6101,N_641,N_109);
nand U6102 (N_6102,N_4030,N_2357);
or U6103 (N_6103,N_4141,N_4678);
xor U6104 (N_6104,N_2087,N_4473);
or U6105 (N_6105,N_3634,N_2059);
or U6106 (N_6106,N_2057,N_3233);
or U6107 (N_6107,N_2661,N_4167);
nand U6108 (N_6108,N_3148,N_1819);
nand U6109 (N_6109,N_2106,N_3354);
or U6110 (N_6110,N_3484,N_1129);
or U6111 (N_6111,N_1402,N_4395);
and U6112 (N_6112,N_1017,N_4043);
and U6113 (N_6113,N_2719,N_4169);
xor U6114 (N_6114,N_3278,N_2454);
xnor U6115 (N_6115,N_3496,N_3755);
xor U6116 (N_6116,N_2916,N_1387);
and U6117 (N_6117,N_1951,N_4896);
xnor U6118 (N_6118,N_3540,N_4733);
and U6119 (N_6119,N_1204,N_4135);
or U6120 (N_6120,N_2726,N_883);
and U6121 (N_6121,N_3875,N_1803);
nand U6122 (N_6122,N_2692,N_4117);
nand U6123 (N_6123,N_4273,N_3555);
nor U6124 (N_6124,N_1617,N_2074);
xor U6125 (N_6125,N_1099,N_3010);
xnor U6126 (N_6126,N_22,N_24);
and U6127 (N_6127,N_223,N_547);
nor U6128 (N_6128,N_2877,N_4446);
and U6129 (N_6129,N_2194,N_1726);
nor U6130 (N_6130,N_3621,N_4594);
nor U6131 (N_6131,N_2099,N_2360);
or U6132 (N_6132,N_992,N_3494);
and U6133 (N_6133,N_4844,N_2663);
nand U6134 (N_6134,N_3640,N_2898);
and U6135 (N_6135,N_3303,N_2697);
or U6136 (N_6136,N_835,N_2717);
or U6137 (N_6137,N_4046,N_3814);
xor U6138 (N_6138,N_3654,N_3497);
nand U6139 (N_6139,N_4873,N_3311);
nor U6140 (N_6140,N_302,N_171);
nand U6141 (N_6141,N_2365,N_2389);
nand U6142 (N_6142,N_4305,N_4409);
nor U6143 (N_6143,N_3825,N_1372);
and U6144 (N_6144,N_756,N_3073);
and U6145 (N_6145,N_2148,N_394);
nor U6146 (N_6146,N_4396,N_4375);
nor U6147 (N_6147,N_2180,N_571);
xor U6148 (N_6148,N_1476,N_3236);
xnor U6149 (N_6149,N_3580,N_2206);
or U6150 (N_6150,N_758,N_4239);
and U6151 (N_6151,N_14,N_4491);
and U6152 (N_6152,N_367,N_3436);
xnor U6153 (N_6153,N_4132,N_2852);
nand U6154 (N_6154,N_569,N_4719);
xnor U6155 (N_6155,N_3408,N_2014);
nor U6156 (N_6156,N_4718,N_1813);
nor U6157 (N_6157,N_771,N_1166);
or U6158 (N_6158,N_1078,N_905);
and U6159 (N_6159,N_3644,N_1450);
and U6160 (N_6160,N_1639,N_2593);
or U6161 (N_6161,N_378,N_3140);
and U6162 (N_6162,N_3393,N_2502);
and U6163 (N_6163,N_1818,N_4364);
and U6164 (N_6164,N_1324,N_4716);
and U6165 (N_6165,N_146,N_654);
and U6166 (N_6166,N_509,N_1226);
nand U6167 (N_6167,N_2779,N_4582);
or U6168 (N_6168,N_698,N_636);
nor U6169 (N_6169,N_3102,N_3841);
xnor U6170 (N_6170,N_2413,N_4398);
nor U6171 (N_6171,N_1686,N_4538);
or U6172 (N_6172,N_789,N_4058);
nor U6173 (N_6173,N_2755,N_544);
nor U6174 (N_6174,N_1640,N_1077);
or U6175 (N_6175,N_3165,N_2575);
or U6176 (N_6176,N_2079,N_2442);
nor U6177 (N_6177,N_1573,N_3818);
nand U6178 (N_6178,N_710,N_91);
and U6179 (N_6179,N_3659,N_2261);
nand U6180 (N_6180,N_2831,N_2774);
and U6181 (N_6181,N_3591,N_4460);
and U6182 (N_6182,N_1759,N_3713);
and U6183 (N_6183,N_4654,N_345);
and U6184 (N_6184,N_4572,N_3524);
or U6185 (N_6185,N_1415,N_4373);
nand U6186 (N_6186,N_4659,N_3858);
and U6187 (N_6187,N_3173,N_1734);
and U6188 (N_6188,N_4983,N_846);
nand U6189 (N_6189,N_1993,N_2401);
nand U6190 (N_6190,N_1456,N_1189);
and U6191 (N_6191,N_4051,N_4284);
and U6192 (N_6192,N_1992,N_2167);
nand U6193 (N_6193,N_1574,N_4280);
or U6194 (N_6194,N_1785,N_4600);
xor U6195 (N_6195,N_4110,N_4675);
and U6196 (N_6196,N_4764,N_1462);
or U6197 (N_6197,N_522,N_4382);
xor U6198 (N_6198,N_4235,N_1921);
or U6199 (N_6199,N_2611,N_2982);
xnor U6200 (N_6200,N_2295,N_1276);
nor U6201 (N_6201,N_3280,N_4832);
or U6202 (N_6202,N_4725,N_2486);
nor U6203 (N_6203,N_1029,N_3485);
nand U6204 (N_6204,N_733,N_2508);
xor U6205 (N_6205,N_1127,N_2551);
and U6206 (N_6206,N_1086,N_4605);
and U6207 (N_6207,N_3552,N_3784);
or U6208 (N_6208,N_822,N_524);
xor U6209 (N_6209,N_796,N_3121);
or U6210 (N_6210,N_2376,N_2891);
xor U6211 (N_6211,N_4655,N_1971);
xnor U6212 (N_6212,N_1554,N_340);
or U6213 (N_6213,N_2671,N_2624);
nor U6214 (N_6214,N_4495,N_518);
xnor U6215 (N_6215,N_3120,N_3094);
nor U6216 (N_6216,N_3212,N_324);
and U6217 (N_6217,N_3660,N_1551);
and U6218 (N_6218,N_3676,N_2751);
nand U6219 (N_6219,N_4794,N_2856);
and U6220 (N_6220,N_3518,N_227);
and U6221 (N_6221,N_1384,N_3785);
and U6222 (N_6222,N_817,N_2687);
and U6223 (N_6223,N_4677,N_1959);
nand U6224 (N_6224,N_1562,N_4370);
nor U6225 (N_6225,N_4202,N_4981);
xor U6226 (N_6226,N_3743,N_1334);
and U6227 (N_6227,N_996,N_3291);
nor U6228 (N_6228,N_1240,N_4706);
nor U6229 (N_6229,N_3972,N_4485);
nor U6230 (N_6230,N_2509,N_4523);
nor U6231 (N_6231,N_1747,N_3459);
xnor U6232 (N_6232,N_4536,N_1541);
nor U6233 (N_6233,N_291,N_3154);
nor U6234 (N_6234,N_3609,N_2218);
nor U6235 (N_6235,N_2565,N_1718);
nor U6236 (N_6236,N_1466,N_4428);
nand U6237 (N_6237,N_1369,N_4018);
nand U6238 (N_6238,N_4690,N_51);
or U6239 (N_6239,N_4186,N_4422);
or U6240 (N_6240,N_574,N_4762);
xor U6241 (N_6241,N_3117,N_338);
nor U6242 (N_6242,N_751,N_3562);
nand U6243 (N_6243,N_4991,N_98);
or U6244 (N_6244,N_950,N_3224);
nor U6245 (N_6245,N_4016,N_2381);
or U6246 (N_6246,N_4268,N_3295);
nor U6247 (N_6247,N_1444,N_3396);
xnor U6248 (N_6248,N_892,N_163);
or U6249 (N_6249,N_3365,N_4078);
xnor U6250 (N_6250,N_573,N_2504);
or U6251 (N_6251,N_3996,N_757);
or U6252 (N_6252,N_1836,N_3254);
nor U6253 (N_6253,N_3800,N_4223);
xor U6254 (N_6254,N_1147,N_3603);
nand U6255 (N_6255,N_3626,N_651);
nand U6256 (N_6256,N_1881,N_165);
and U6257 (N_6257,N_1521,N_2971);
nand U6258 (N_6258,N_3098,N_1065);
xor U6259 (N_6259,N_293,N_2516);
or U6260 (N_6260,N_2166,N_1589);
and U6261 (N_6261,N_2213,N_2924);
xnor U6262 (N_6262,N_2946,N_2362);
nor U6263 (N_6263,N_2641,N_3209);
and U6264 (N_6264,N_3141,N_447);
and U6265 (N_6265,N_2913,N_261);
or U6266 (N_6266,N_4118,N_4987);
nor U6267 (N_6267,N_2036,N_463);
and U6268 (N_6268,N_3862,N_3712);
nor U6269 (N_6269,N_1448,N_1012);
nor U6270 (N_6270,N_4241,N_1750);
xor U6271 (N_6271,N_4405,N_1263);
and U6272 (N_6272,N_36,N_1018);
xor U6273 (N_6273,N_4962,N_138);
and U6274 (N_6274,N_4599,N_2892);
and U6275 (N_6275,N_1508,N_2430);
nor U6276 (N_6276,N_193,N_407);
nand U6277 (N_6277,N_1495,N_4877);
xor U6278 (N_6278,N_239,N_1652);
nor U6279 (N_6279,N_1610,N_4822);
nand U6280 (N_6280,N_3662,N_1626);
and U6281 (N_6281,N_4036,N_4329);
or U6282 (N_6282,N_1641,N_606);
xor U6283 (N_6283,N_1752,N_2117);
or U6284 (N_6284,N_4663,N_4629);
or U6285 (N_6285,N_2631,N_4045);
nor U6286 (N_6286,N_4610,N_1805);
xnor U6287 (N_6287,N_1357,N_2018);
and U6288 (N_6288,N_2312,N_1438);
xor U6289 (N_6289,N_993,N_2648);
nor U6290 (N_6290,N_1339,N_4574);
nor U6291 (N_6291,N_1633,N_3347);
or U6292 (N_6292,N_910,N_2003);
or U6293 (N_6293,N_2217,N_4367);
or U6294 (N_6294,N_3220,N_537);
or U6295 (N_6295,N_2112,N_970);
nor U6296 (N_6296,N_4549,N_4567);
nand U6297 (N_6297,N_4888,N_3598);
nand U6298 (N_6298,N_3614,N_903);
and U6299 (N_6299,N_3479,N_1991);
nand U6300 (N_6300,N_1470,N_675);
nand U6301 (N_6301,N_4695,N_2024);
or U6302 (N_6302,N_2313,N_2490);
nor U6303 (N_6303,N_4938,N_961);
or U6304 (N_6304,N_4349,N_2917);
nor U6305 (N_6305,N_2234,N_1613);
and U6306 (N_6306,N_4423,N_2328);
nor U6307 (N_6307,N_723,N_3605);
nand U6308 (N_6308,N_2498,N_1469);
nor U6309 (N_6309,N_1925,N_462);
and U6310 (N_6310,N_1702,N_2842);
or U6311 (N_6311,N_2632,N_3189);
nor U6312 (N_6312,N_3522,N_1256);
or U6313 (N_6313,N_3032,N_1210);
and U6314 (N_6314,N_624,N_1027);
or U6315 (N_6315,N_4299,N_1392);
nor U6316 (N_6316,N_3257,N_4724);
nand U6317 (N_6317,N_2472,N_2185);
nand U6318 (N_6318,N_3356,N_3588);
nor U6319 (N_6319,N_1039,N_2426);
or U6320 (N_6320,N_2178,N_2539);
xnor U6321 (N_6321,N_4196,N_4471);
or U6322 (N_6322,N_1801,N_3501);
or U6323 (N_6323,N_695,N_4959);
or U6324 (N_6324,N_866,N_4026);
nand U6325 (N_6325,N_907,N_1507);
nor U6326 (N_6326,N_3913,N_1325);
nor U6327 (N_6327,N_4717,N_2659);
nor U6328 (N_6328,N_141,N_4914);
xnor U6329 (N_6329,N_525,N_1215);
xnor U6330 (N_6330,N_257,N_979);
xor U6331 (N_6331,N_2330,N_3330);
nor U6332 (N_6332,N_2023,N_773);
nor U6333 (N_6333,N_3804,N_1784);
nor U6334 (N_6334,N_3958,N_2069);
and U6335 (N_6335,N_973,N_3182);
and U6336 (N_6336,N_3296,N_2736);
nand U6337 (N_6337,N_4341,N_1005);
nand U6338 (N_6338,N_3113,N_1711);
xor U6339 (N_6339,N_279,N_3663);
nand U6340 (N_6340,N_1844,N_2062);
nor U6341 (N_6341,N_2996,N_4751);
xnor U6342 (N_6342,N_3719,N_4357);
or U6343 (N_6343,N_1975,N_2456);
xnor U6344 (N_6344,N_480,N_4315);
and U6345 (N_6345,N_4044,N_4714);
or U6346 (N_6346,N_2695,N_890);
or U6347 (N_6347,N_2393,N_836);
nor U6348 (N_6348,N_2951,N_4862);
xnor U6349 (N_6349,N_3708,N_3571);
xor U6350 (N_6350,N_4378,N_3569);
nand U6351 (N_6351,N_108,N_459);
nor U6352 (N_6352,N_2292,N_3495);
and U6353 (N_6353,N_126,N_3868);
nor U6354 (N_6354,N_3886,N_3328);
and U6355 (N_6355,N_2787,N_3782);
nor U6356 (N_6356,N_3076,N_4507);
nor U6357 (N_6357,N_3314,N_3752);
nand U6358 (N_6358,N_769,N_3581);
or U6359 (N_6359,N_3456,N_3856);
xnor U6360 (N_6360,N_4476,N_4385);
xnor U6361 (N_6361,N_1522,N_1138);
nor U6362 (N_6362,N_3896,N_3773);
and U6363 (N_6363,N_3435,N_563);
or U6364 (N_6364,N_203,N_2639);
or U6365 (N_6365,N_1236,N_1692);
nand U6366 (N_6366,N_3414,N_3929);
nor U6367 (N_6367,N_4784,N_149);
xnor U6368 (N_6368,N_3014,N_3990);
nor U6369 (N_6369,N_496,N_256);
nand U6370 (N_6370,N_2547,N_369);
nor U6371 (N_6371,N_1031,N_3874);
or U6372 (N_6372,N_1663,N_4440);
and U6373 (N_6373,N_2021,N_3277);
nand U6374 (N_6374,N_2561,N_3235);
xor U6375 (N_6375,N_186,N_179);
xnor U6376 (N_6376,N_4563,N_365);
and U6377 (N_6377,N_953,N_2607);
nand U6378 (N_6378,N_1306,N_3848);
nor U6379 (N_6379,N_2501,N_1087);
or U6380 (N_6380,N_2713,N_428);
xnor U6381 (N_6381,N_2123,N_3397);
xnor U6382 (N_6382,N_4705,N_767);
xor U6383 (N_6383,N_1619,N_53);
nand U6384 (N_6384,N_3391,N_4934);
nor U6385 (N_6385,N_4436,N_1467);
and U6386 (N_6386,N_3610,N_2126);
xnor U6387 (N_6387,N_4199,N_2143);
xor U6388 (N_6388,N_1624,N_4294);
and U6389 (N_6389,N_687,N_4840);
nor U6390 (N_6390,N_2140,N_4992);
nand U6391 (N_6391,N_4142,N_3645);
or U6392 (N_6392,N_2183,N_1654);
or U6393 (N_6393,N_581,N_1497);
and U6394 (N_6394,N_4472,N_566);
nor U6395 (N_6395,N_1316,N_2029);
or U6396 (N_6396,N_1699,N_1371);
nand U6397 (N_6397,N_2967,N_3607);
xnor U6398 (N_6398,N_1484,N_909);
xnor U6399 (N_6399,N_1605,N_4425);
and U6400 (N_6400,N_4781,N_3447);
and U6401 (N_6401,N_4333,N_4176);
xnor U6402 (N_6402,N_1909,N_1731);
and U6403 (N_6403,N_460,N_4564);
or U6404 (N_6404,N_1433,N_442);
nand U6405 (N_6405,N_2840,N_622);
nor U6406 (N_6406,N_3928,N_1404);
nor U6407 (N_6407,N_3271,N_1252);
nor U6408 (N_6408,N_1082,N_3885);
xor U6409 (N_6409,N_1045,N_2100);
nor U6410 (N_6410,N_4731,N_2200);
and U6411 (N_6411,N_4520,N_3344);
and U6412 (N_6412,N_1978,N_4115);
nor U6413 (N_6413,N_1814,N_2375);
and U6414 (N_6414,N_653,N_1597);
nand U6415 (N_6415,N_1118,N_1546);
nand U6416 (N_6416,N_2150,N_1477);
xor U6417 (N_6417,N_858,N_3251);
and U6418 (N_6418,N_1915,N_3988);
xnor U6419 (N_6419,N_4401,N_3122);
or U6420 (N_6420,N_4470,N_2157);
nand U6421 (N_6421,N_3867,N_2636);
nor U6422 (N_6422,N_4213,N_2409);
and U6423 (N_6423,N_2513,N_3263);
xnor U6424 (N_6424,N_4348,N_3193);
and U6425 (N_6425,N_2625,N_3523);
and U6426 (N_6426,N_1857,N_233);
and U6427 (N_6427,N_2793,N_2919);
xnor U6428 (N_6428,N_4104,N_4234);
and U6429 (N_6429,N_1896,N_4362);
nor U6430 (N_6430,N_1350,N_2839);
and U6431 (N_6431,N_4236,N_2559);
or U6432 (N_6432,N_2314,N_4127);
nor U6433 (N_6433,N_458,N_4689);
and U6434 (N_6434,N_3367,N_930);
xnor U6435 (N_6435,N_4577,N_706);
nand U6436 (N_6436,N_4302,N_1206);
nand U6437 (N_6437,N_2809,N_3190);
xnor U6438 (N_6438,N_2301,N_1920);
nand U6439 (N_6439,N_0,N_575);
nor U6440 (N_6440,N_652,N_3717);
and U6441 (N_6441,N_2572,N_2221);
nand U6442 (N_6442,N_2773,N_1933);
xor U6443 (N_6443,N_3287,N_929);
or U6444 (N_6444,N_4693,N_2247);
or U6445 (N_6445,N_3992,N_1983);
nand U6446 (N_6446,N_2705,N_2267);
nand U6447 (N_6447,N_3846,N_2642);
or U6448 (N_6448,N_4319,N_3542);
and U6449 (N_6449,N_2043,N_3196);
nor U6450 (N_6450,N_1041,N_1807);
nor U6451 (N_6451,N_2794,N_3066);
nand U6452 (N_6452,N_282,N_631);
nor U6453 (N_6453,N_1009,N_596);
nor U6454 (N_6454,N_3107,N_2886);
xor U6455 (N_6455,N_2830,N_4230);
nand U6456 (N_6456,N_4024,N_4905);
nand U6457 (N_6457,N_1646,N_599);
or U6458 (N_6458,N_2434,N_380);
or U6459 (N_6459,N_604,N_3221);
or U6460 (N_6460,N_1649,N_213);
nand U6461 (N_6461,N_3316,N_482);
or U6462 (N_6462,N_3612,N_4554);
and U6463 (N_6463,N_1390,N_3353);
xor U6464 (N_6464,N_2804,N_2104);
nand U6465 (N_6465,N_4338,N_2776);
nand U6466 (N_6466,N_4497,N_1449);
nor U6467 (N_6467,N_2492,N_259);
or U6468 (N_6468,N_4100,N_3766);
and U6469 (N_6469,N_4638,N_2775);
or U6470 (N_6470,N_904,N_406);
or U6471 (N_6471,N_1105,N_46);
xor U6472 (N_6472,N_2614,N_1489);
nand U6473 (N_6473,N_2598,N_2820);
xnor U6474 (N_6474,N_803,N_4355);
and U6475 (N_6475,N_4857,N_4442);
nand U6476 (N_6476,N_2152,N_4579);
and U6477 (N_6477,N_2758,N_1453);
xor U6478 (N_6478,N_472,N_1380);
and U6479 (N_6479,N_1667,N_4350);
and U6480 (N_6480,N_4054,N_3286);
nand U6481 (N_6481,N_2784,N_4867);
nor U6482 (N_6482,N_3046,N_2959);
and U6483 (N_6483,N_2336,N_1410);
or U6484 (N_6484,N_2278,N_797);
or U6485 (N_6485,N_976,N_494);
or U6486 (N_6486,N_3080,N_3127);
or U6487 (N_6487,N_147,N_2612);
nand U6488 (N_6488,N_2411,N_4528);
or U6489 (N_6489,N_2664,N_4418);
or U6490 (N_6490,N_1676,N_3771);
or U6491 (N_6491,N_3237,N_2481);
xnor U6492 (N_6492,N_276,N_3730);
nor U6493 (N_6493,N_4779,N_4238);
nand U6494 (N_6494,N_204,N_3821);
nand U6495 (N_6495,N_3608,N_4841);
nor U6496 (N_6496,N_3699,N_3734);
and U6497 (N_6497,N_3859,N_1893);
xnor U6498 (N_6498,N_411,N_4771);
or U6499 (N_6499,N_3487,N_274);
and U6500 (N_6500,N_3698,N_2223);
and U6501 (N_6501,N_4526,N_272);
or U6502 (N_6502,N_4692,N_3671);
and U6503 (N_6503,N_2807,N_627);
or U6504 (N_6504,N_2897,N_4828);
and U6505 (N_6505,N_4151,N_3276);
xor U6506 (N_6506,N_1719,N_1728);
nand U6507 (N_6507,N_2786,N_1612);
nand U6508 (N_6508,N_4664,N_1259);
xor U6509 (N_6509,N_3384,N_3394);
nor U6510 (N_6510,N_1894,N_4744);
nand U6511 (N_6511,N_134,N_4860);
nor U6512 (N_6512,N_1304,N_1378);
nand U6513 (N_6513,N_2053,N_2878);
or U6514 (N_6514,N_3934,N_2528);
nand U6515 (N_6515,N_2566,N_4478);
xor U6516 (N_6516,N_4449,N_2866);
and U6517 (N_6517,N_3649,N_3427);
xnor U6518 (N_6518,N_1110,N_1292);
xor U6519 (N_6519,N_1419,N_382);
and U6520 (N_6520,N_4314,N_1447);
nand U6521 (N_6521,N_2195,N_3418);
or U6522 (N_6522,N_3650,N_431);
nor U6523 (N_6523,N_4207,N_1442);
xor U6524 (N_6524,N_250,N_4769);
xnor U6525 (N_6525,N_334,N_317);
or U6526 (N_6526,N_2582,N_2734);
or U6527 (N_6527,N_2732,N_1076);
or U6528 (N_6528,N_1989,N_1910);
or U6529 (N_6529,N_1186,N_4264);
and U6530 (N_6530,N_2512,N_702);
nand U6531 (N_6531,N_1229,N_520);
nand U6532 (N_6532,N_1053,N_4451);
nor U6533 (N_6533,N_3179,N_2615);
nor U6534 (N_6534,N_1678,N_277);
nand U6535 (N_6535,N_2862,N_1363);
nand U6536 (N_6536,N_942,N_2628);
and U6537 (N_6537,N_1788,N_990);
and U6538 (N_6538,N_3797,N_1176);
and U6539 (N_6539,N_1310,N_4298);
xnor U6540 (N_6540,N_2291,N_128);
xnor U6541 (N_6541,N_4713,N_2699);
nand U6542 (N_6542,N_3651,N_3879);
xor U6543 (N_6543,N_3168,N_2243);
nor U6544 (N_6544,N_3914,N_3872);
or U6545 (N_6545,N_4432,N_4340);
and U6546 (N_6546,N_3927,N_2608);
and U6547 (N_6547,N_2952,N_4288);
nor U6548 (N_6548,N_4516,N_1707);
nor U6549 (N_6549,N_1591,N_703);
and U6550 (N_6550,N_1046,N_2550);
and U6551 (N_6551,N_4287,N_2436);
nand U6552 (N_6552,N_3282,N_879);
or U6553 (N_6553,N_3536,N_4361);
and U6554 (N_6554,N_1965,N_1376);
nand U6555 (N_6555,N_647,N_1258);
or U6556 (N_6556,N_2778,N_3751);
or U6557 (N_6557,N_290,N_3323);
or U6558 (N_6558,N_3409,N_634);
nand U6559 (N_6559,N_4685,N_2765);
or U6560 (N_6560,N_1565,N_4730);
nor U6561 (N_6561,N_679,N_1681);
and U6562 (N_6562,N_1669,N_1891);
nor U6563 (N_6563,N_1246,N_1159);
and U6564 (N_6564,N_2164,N_3844);
or U6565 (N_6565,N_86,N_124);
nor U6566 (N_6566,N_4443,N_3909);
and U6567 (N_6567,N_629,N_791);
nor U6568 (N_6568,N_2230,N_1295);
nor U6569 (N_6569,N_3756,N_2276);
nand U6570 (N_6570,N_657,N_2990);
nor U6571 (N_6571,N_4861,N_2358);
xor U6572 (N_6572,N_3298,N_1155);
or U6573 (N_6573,N_1882,N_4852);
nor U6574 (N_6574,N_310,N_1859);
or U6575 (N_6575,N_582,N_934);
xnor U6576 (N_6576,N_4571,N_1947);
nand U6577 (N_6577,N_1351,N_2303);
nand U6578 (N_6578,N_660,N_3019);
nor U6579 (N_6579,N_3412,N_1696);
or U6580 (N_6580,N_1199,N_1216);
xnor U6581 (N_6581,N_1763,N_4295);
nor U6582 (N_6582,N_4289,N_2989);
nand U6583 (N_6583,N_555,N_2569);
xnor U6584 (N_6584,N_4206,N_2346);
and U6585 (N_6585,N_4224,N_4087);
or U6586 (N_6586,N_526,N_4069);
xor U6587 (N_6587,N_1751,N_1499);
and U6588 (N_6588,N_1564,N_868);
and U6589 (N_6589,N_3070,N_4335);
xor U6590 (N_6590,N_543,N_454);
nand U6591 (N_6591,N_1173,N_1906);
and U6592 (N_6592,N_1375,N_1417);
and U6593 (N_6593,N_4301,N_861);
or U6594 (N_6594,N_2921,N_2749);
nand U6595 (N_6595,N_1092,N_2965);
nor U6596 (N_6596,N_1160,N_3559);
nand U6597 (N_6597,N_1478,N_3139);
xor U6598 (N_6598,N_1095,N_3675);
nor U6599 (N_6599,N_1403,N_4218);
nand U6600 (N_6600,N_3275,N_1393);
and U6601 (N_6601,N_888,N_404);
nand U6602 (N_6602,N_105,N_1211);
nand U6603 (N_6603,N_374,N_1047);
xor U6604 (N_6604,N_2082,N_819);
nand U6605 (N_6605,N_2922,N_2286);
or U6606 (N_6606,N_1439,N_3093);
nor U6607 (N_6607,N_1628,N_915);
and U6608 (N_6608,N_3638,N_2190);
and U6609 (N_6609,N_3119,N_422);
nor U6610 (N_6610,N_2654,N_457);
or U6611 (N_6611,N_2597,N_3777);
nand U6612 (N_6612,N_1722,N_1451);
and U6613 (N_6613,N_2406,N_85);
nand U6614 (N_6614,N_3381,N_3944);
nand U6615 (N_6615,N_1142,N_3468);
and U6616 (N_6616,N_2738,N_4870);
nand U6617 (N_6617,N_3238,N_4469);
nor U6618 (N_6618,N_3369,N_1479);
xor U6619 (N_6619,N_561,N_326);
nand U6620 (N_6620,N_2975,N_4098);
xor U6621 (N_6621,N_1645,N_1706);
nor U6622 (N_6622,N_1568,N_1399);
nand U6623 (N_6623,N_3582,N_4159);
nor U6624 (N_6624,N_3059,N_1727);
xor U6625 (N_6625,N_4351,N_2196);
nand U6626 (N_6626,N_1616,N_1434);
xnor U6627 (N_6627,N_4868,N_2440);
or U6628 (N_6628,N_4829,N_2948);
nand U6629 (N_6629,N_2052,N_4270);
nand U6630 (N_6630,N_2995,N_1748);
nor U6631 (N_6631,N_166,N_2694);
nor U6632 (N_6632,N_3504,N_4041);
and U6633 (N_6633,N_3438,N_937);
or U6634 (N_6634,N_1436,N_2340);
xor U6635 (N_6635,N_2702,N_2834);
or U6636 (N_6636,N_4756,N_1128);
or U6637 (N_6637,N_476,N_4532);
nor U6638 (N_6638,N_1519,N_1927);
nor U6639 (N_6639,N_2283,N_4950);
xor U6640 (N_6640,N_3031,N_61);
and U6641 (N_6641,N_714,N_3714);
nor U6642 (N_6642,N_972,N_1406);
nor U6643 (N_6643,N_2746,N_2311);
nand U6644 (N_6644,N_1030,N_3177);
or U6645 (N_6645,N_3796,N_4450);
and U6646 (N_6646,N_1455,N_3351);
xnor U6647 (N_6647,N_2063,N_1347);
nor U6648 (N_6648,N_2954,N_488);
xor U6649 (N_6649,N_3252,N_1720);
or U6650 (N_6650,N_3355,N_3415);
nand U6651 (N_6651,N_1485,N_397);
and U6652 (N_6652,N_1033,N_3798);
or U6653 (N_6653,N_2696,N_947);
nand U6654 (N_6654,N_2617,N_1585);
and U6655 (N_6655,N_2968,N_133);
xor U6656 (N_6656,N_1075,N_329);
or U6657 (N_6657,N_1733,N_2548);
or U6658 (N_6658,N_1400,N_785);
nor U6659 (N_6659,N_4111,N_4742);
nand U6660 (N_6660,N_4228,N_3490);
xnor U6661 (N_6661,N_1929,N_820);
or U6662 (N_6662,N_4049,N_3692);
xnor U6663 (N_6663,N_1052,N_4347);
and U6664 (N_6664,N_1558,N_664);
nand U6665 (N_6665,N_106,N_4211);
nor U6666 (N_6666,N_922,N_3578);
nor U6667 (N_6667,N_2137,N_2981);
xnor U6668 (N_6668,N_564,N_4499);
nor U6669 (N_6669,N_862,N_1913);
nand U6670 (N_6670,N_1353,N_3162);
xor U6671 (N_6671,N_4474,N_3901);
and U6672 (N_6672,N_1249,N_3916);
nor U6673 (N_6673,N_278,N_207);
nand U6674 (N_6674,N_853,N_2950);
nor U6675 (N_6675,N_1599,N_3517);
or U6676 (N_6676,N_1866,N_3842);
and U6677 (N_6677,N_1024,N_260);
and U6678 (N_6678,N_3036,N_4558);
or U6679 (N_6679,N_960,N_1019);
or U6680 (N_6680,N_3701,N_3726);
xor U6681 (N_6681,N_1062,N_4023);
or U6682 (N_6682,N_1103,N_4642);
nor U6683 (N_6683,N_3227,N_21);
nand U6684 (N_6684,N_3572,N_3321);
nor U6685 (N_6685,N_677,N_4805);
nand U6686 (N_6686,N_4136,N_3028);
nand U6687 (N_6687,N_3961,N_3180);
nor U6688 (N_6688,N_583,N_4752);
and U6689 (N_6689,N_198,N_4073);
nor U6690 (N_6690,N_2510,N_3792);
and U6691 (N_6691,N_1432,N_2239);
and U6692 (N_6692,N_388,N_834);
or U6693 (N_6693,N_2324,N_1397);
or U6694 (N_6694,N_512,N_2700);
nand U6695 (N_6695,N_4123,N_681);
nand U6696 (N_6696,N_2910,N_3360);
nand U6697 (N_6697,N_2394,N_3735);
nand U6698 (N_6698,N_4575,N_2208);
and U6699 (N_6699,N_2246,N_47);
nand U6700 (N_6700,N_919,N_383);
nand U6701 (N_6701,N_3682,N_4486);
nor U6702 (N_6702,N_2693,N_3201);
or U6703 (N_6703,N_1474,N_3214);
and U6704 (N_6704,N_4038,N_2333);
xor U6705 (N_6705,N_2955,N_4539);
xnor U6706 (N_6706,N_2458,N_3413);
xnor U6707 (N_6707,N_1381,N_1520);
nand U6708 (N_6708,N_1800,N_1831);
nand U6709 (N_6709,N_2511,N_2322);
and U6710 (N_6710,N_1611,N_1289);
xor U6711 (N_6711,N_2012,N_3973);
and U6712 (N_6712,N_2441,N_4581);
and U6713 (N_6713,N_1572,N_1642);
nand U6714 (N_6714,N_2803,N_1791);
or U6715 (N_6715,N_4277,N_1340);
nand U6716 (N_6716,N_538,N_2896);
nand U6717 (N_6717,N_4933,N_1398);
nor U6718 (N_6718,N_810,N_3150);
nor U6719 (N_6719,N_4042,N_4099);
nor U6720 (N_6720,N_2118,N_665);
and U6721 (N_6721,N_2496,N_1242);
or U6722 (N_6722,N_2602,N_2480);
xnor U6723 (N_6723,N_1311,N_776);
or U6724 (N_6724,N_1021,N_1988);
nand U6725 (N_6725,N_4565,N_3050);
xnor U6726 (N_6726,N_4416,N_967);
and U6727 (N_6727,N_1783,N_1765);
nand U6728 (N_6728,N_1265,N_4699);
xnor U6729 (N_6729,N_3673,N_410);
or U6730 (N_6730,N_235,N_4327);
and U6731 (N_6731,N_4028,N_1664);
nand U6732 (N_6732,N_4910,N_692);
xor U6733 (N_6733,N_3965,N_3951);
nand U6734 (N_6734,N_266,N_2847);
nor U6735 (N_6735,N_2681,N_4201);
and U6736 (N_6736,N_209,N_4767);
or U6737 (N_6737,N_2684,N_3085);
nand U6738 (N_6738,N_2737,N_3565);
and U6739 (N_6739,N_1793,N_4957);
and U6740 (N_6740,N_4293,N_4625);
or U6741 (N_6741,N_1675,N_1222);
nor U6742 (N_6742,N_2601,N_4702);
nor U6743 (N_6743,N_2998,N_3187);
and U6744 (N_6744,N_3681,N_2279);
nand U6745 (N_6745,N_445,N_4269);
or U6746 (N_6746,N_4056,N_4737);
or U6747 (N_6747,N_2315,N_4787);
nor U6748 (N_6748,N_2826,N_1073);
xnor U6749 (N_6749,N_716,N_3590);
or U6750 (N_6750,N_3338,N_1665);
or U6751 (N_6751,N_3622,N_1234);
and U6752 (N_6752,N_4297,N_3624);
xor U6753 (N_6753,N_3458,N_3161);
and U6754 (N_6754,N_1892,N_4647);
or U6755 (N_6755,N_3506,N_2858);
and U6756 (N_6756,N_1700,N_1742);
or U6757 (N_6757,N_358,N_1709);
xnor U6758 (N_6758,N_2798,N_2864);
nand U6759 (N_6759,N_4885,N_717);
nor U6760 (N_6760,N_553,N_357);
or U6761 (N_6761,N_173,N_4953);
or U6762 (N_6762,N_342,N_1907);
xor U6763 (N_6763,N_607,N_1590);
nand U6764 (N_6764,N_1238,N_1130);
and U6765 (N_6765,N_704,N_2782);
or U6766 (N_6766,N_3765,N_1235);
nor U6767 (N_6767,N_3983,N_465);
nand U6768 (N_6768,N_531,N_4454);
nand U6769 (N_6769,N_2753,N_726);
and U6770 (N_6770,N_3679,N_4191);
nand U6771 (N_6771,N_921,N_2783);
nand U6772 (N_6772,N_2371,N_3072);
or U6773 (N_6773,N_3788,N_4458);
xor U6774 (N_6774,N_3986,N_4065);
and U6775 (N_6775,N_205,N_1098);
or U6776 (N_6776,N_3457,N_1500);
nand U6777 (N_6777,N_23,N_2546);
nor U6778 (N_6778,N_1637,N_762);
nand U6779 (N_6779,N_456,N_3289);
and U6780 (N_6780,N_1737,N_3299);
nor U6781 (N_6781,N_4772,N_2418);
and U6782 (N_6782,N_1302,N_1630);
or U6783 (N_6783,N_3454,N_13);
or U6784 (N_6784,N_4021,N_2075);
nor U6785 (N_6785,N_4641,N_2522);
nor U6786 (N_6786,N_1994,N_1595);
nand U6787 (N_6787,N_2577,N_1187);
nand U6788 (N_6788,N_3284,N_1583);
and U6789 (N_6789,N_4022,N_3723);
nor U6790 (N_6790,N_1509,N_2116);
xor U6791 (N_6791,N_3652,N_4007);
nor U6792 (N_6792,N_188,N_4237);
nand U6793 (N_6793,N_4961,N_4140);
nor U6794 (N_6794,N_4080,N_4686);
or U6795 (N_6795,N_4748,N_3787);
or U6796 (N_6796,N_3620,N_4637);
or U6797 (N_6797,N_4537,N_2188);
and U6798 (N_6798,N_4126,N_1346);
nor U6799 (N_6799,N_246,N_3907);
and U6800 (N_6800,N_3325,N_517);
xnor U6801 (N_6801,N_3971,N_1895);
nor U6802 (N_6802,N_117,N_4995);
nand U6803 (N_6803,N_2567,N_4369);
nand U6804 (N_6804,N_2679,N_1115);
or U6805 (N_6805,N_578,N_490);
and U6806 (N_6806,N_1922,N_2690);
nor U6807 (N_6807,N_4630,N_2015);
xor U6808 (N_6808,N_3223,N_882);
or U6809 (N_6809,N_752,N_3955);
nor U6810 (N_6810,N_2795,N_315);
nor U6811 (N_6811,N_4105,N_4859);
and U6812 (N_6812,N_3081,N_4606);
or U6813 (N_6813,N_551,N_4353);
xnor U6814 (N_6814,N_1067,N_4006);
nand U6815 (N_6815,N_4791,N_4484);
nor U6816 (N_6816,N_4250,N_3616);
or U6817 (N_6817,N_4040,N_62);
or U6818 (N_6818,N_493,N_4342);
and U6819 (N_6819,N_4170,N_3759);
nor U6820 (N_6820,N_2960,N_2067);
nor U6821 (N_6821,N_3461,N_1995);
xor U6822 (N_6822,N_4650,N_4682);
xnor U6823 (N_6823,N_3358,N_34);
nor U6824 (N_6824,N_1662,N_1169);
nor U6825 (N_6825,N_1336,N_4157);
nand U6826 (N_6826,N_984,N_2437);
and U6827 (N_6827,N_3693,N_2961);
nor U6828 (N_6828,N_2321,N_73);
xor U6829 (N_6829,N_949,N_232);
nor U6830 (N_6830,N_1170,N_1290);
and U6831 (N_6831,N_4464,N_320);
nand U6832 (N_6832,N_157,N_3112);
and U6833 (N_6833,N_119,N_4502);
nand U6834 (N_6834,N_1762,N_3248);
or U6835 (N_6835,N_2673,N_4524);
nor U6836 (N_6836,N_2495,N_2460);
nand U6837 (N_6837,N_2674,N_2455);
nand U6838 (N_6838,N_4203,N_2464);
and U6839 (N_6839,N_3069,N_3840);
and U6840 (N_6840,N_1280,N_1224);
or U6841 (N_6841,N_804,N_1770);
xor U6842 (N_6842,N_363,N_4093);
or U6843 (N_6843,N_3135,N_4927);
xor U6844 (N_6844,N_4782,N_4890);
nand U6845 (N_6845,N_4292,N_399);
nor U6846 (N_6846,N_1193,N_3337);
or U6847 (N_6847,N_4055,N_4680);
or U6848 (N_6848,N_3106,N_3441);
nor U6849 (N_6849,N_1827,N_4012);
and U6850 (N_6850,N_2588,N_2949);
nor U6851 (N_6851,N_833,N_2163);
and U6852 (N_6852,N_3062,N_3191);
xor U6853 (N_6853,N_4576,N_3586);
nor U6854 (N_6854,N_4148,N_540);
nand U6855 (N_6855,N_1854,N_4691);
xor U6856 (N_6856,N_777,N_2635);
nand U6857 (N_6857,N_4755,N_1824);
nor U6858 (N_6858,N_3567,N_1600);
or U6859 (N_6859,N_3957,N_1632);
or U6860 (N_6860,N_3672,N_4917);
nor U6861 (N_6861,N_775,N_2465);
and U6862 (N_6862,N_3617,N_160);
or U6863 (N_6863,N_311,N_4009);
xor U6864 (N_6864,N_3893,N_4200);
or U6865 (N_6865,N_855,N_1776);
and U6866 (N_6866,N_1278,N_4147);
nand U6867 (N_6867,N_4754,N_1898);
nand U6868 (N_6868,N_1071,N_4976);
xor U6869 (N_6869,N_2222,N_592);
nor U6870 (N_6870,N_1112,N_1006);
xor U6871 (N_6871,N_1165,N_3899);
nor U6872 (N_6872,N_4094,N_3171);
nand U6873 (N_6873,N_3661,N_1307);
nand U6874 (N_6874,N_4121,N_1579);
nand U6875 (N_6875,N_2630,N_1848);
and U6876 (N_6876,N_2649,N_1459);
nor U6877 (N_6877,N_2792,N_4209);
and U6878 (N_6878,N_859,N_985);
xnor U6879 (N_6879,N_3629,N_737);
nand U6880 (N_6880,N_4790,N_954);
and U6881 (N_6881,N_987,N_3851);
nand U6882 (N_6882,N_63,N_4496);
xnor U6883 (N_6883,N_4881,N_572);
and U6884 (N_6884,N_1097,N_49);
and U6885 (N_6885,N_1034,N_4956);
xnor U6886 (N_6886,N_4334,N_1778);
xnor U6887 (N_6887,N_3977,N_74);
xor U6888 (N_6888,N_839,N_4985);
nor U6889 (N_6889,N_4768,N_3372);
nor U6890 (N_6890,N_2925,N_267);
or U6891 (N_6891,N_2640,N_3174);
xnor U6892 (N_6892,N_228,N_99);
and U6893 (N_6893,N_3823,N_4904);
xnor U6894 (N_6894,N_87,N_4778);
nor U6895 (N_6895,N_1182,N_3538);
nand U6896 (N_6896,N_222,N_4561);
nor U6897 (N_6897,N_3793,N_2665);
xnor U6898 (N_6898,N_1779,N_2192);
nand U6899 (N_6899,N_2540,N_4973);
and U6900 (N_6900,N_598,N_4948);
nand U6901 (N_6901,N_4758,N_784);
nand U6902 (N_6902,N_2317,N_1374);
nand U6903 (N_6903,N_1093,N_4090);
and U6904 (N_6904,N_4081,N_3811);
nand U6905 (N_6905,N_3574,N_666);
or U6906 (N_6906,N_4631,N_1548);
nand U6907 (N_6907,N_1291,N_2084);
or U6908 (N_6908,N_3133,N_4371);
nor U6909 (N_6909,N_1740,N_4227);
xnor U6910 (N_6910,N_3288,N_1413);
nor U6911 (N_6911,N_3269,N_4596);
or U6912 (N_6912,N_3175,N_700);
and U6913 (N_6913,N_4922,N_111);
and U6914 (N_6914,N_3549,N_1123);
and U6915 (N_6915,N_2080,N_4008);
xor U6916 (N_6916,N_2165,N_3695);
nor U6917 (N_6917,N_1262,N_444);
nor U6918 (N_6918,N_3791,N_2843);
xnor U6919 (N_6919,N_3747,N_2049);
and U6920 (N_6920,N_2412,N_419);
or U6921 (N_6921,N_1950,N_1839);
and U6922 (N_6922,N_935,N_4149);
nor U6923 (N_6923,N_2119,N_2610);
nor U6924 (N_6924,N_1154,N_1622);
and U6925 (N_6925,N_3422,N_3707);
nand U6926 (N_6926,N_2111,N_4321);
nor U6927 (N_6927,N_1191,N_4445);
and U6928 (N_6928,N_2422,N_1757);
and U6929 (N_6929,N_2240,N_3084);
nor U6930 (N_6930,N_1889,N_4825);
nand U6931 (N_6931,N_534,N_1054);
or U6932 (N_6932,N_2957,N_2327);
nand U6933 (N_6933,N_1688,N_2915);
xor U6934 (N_6934,N_1167,N_4034);
nand U6935 (N_6935,N_3585,N_958);
or U6936 (N_6936,N_2141,N_3420);
xnor U6937 (N_6937,N_1984,N_3281);
nor U6938 (N_6938,N_2815,N_3968);
and U6939 (N_6939,N_2396,N_3008);
and U6940 (N_6940,N_4383,N_3776);
nor U6941 (N_6941,N_4392,N_2384);
xor U6942 (N_6942,N_2383,N_1575);
and U6943 (N_6943,N_2752,N_3917);
or U6944 (N_6944,N_699,N_1269);
and U6945 (N_6945,N_3613,N_247);
and U6946 (N_6946,N_4982,N_4928);
nand U6947 (N_6947,N_3491,N_4014);
nand U6948 (N_6948,N_2404,N_4408);
xnor U6949 (N_6949,N_1775,N_4271);
or U6950 (N_6950,N_3891,N_2870);
xor U6951 (N_6951,N_4757,N_3361);
xor U6952 (N_6952,N_4517,N_1843);
and U6953 (N_6953,N_4651,N_2980);
xnor U6954 (N_6954,N_2871,N_348);
nor U6955 (N_6955,N_4204,N_3643);
xnor U6956 (N_6956,N_4386,N_2678);
nor U6957 (N_6957,N_2476,N_3205);
nand U6958 (N_6958,N_284,N_3364);
xnor U6959 (N_6959,N_738,N_2515);
xnor U6960 (N_6960,N_3539,N_4232);
and U6961 (N_6961,N_3915,N_2172);
and U6962 (N_6962,N_3007,N_4683);
or U6963 (N_6963,N_4531,N_3342);
or U6964 (N_6964,N_2757,N_4587);
or U6965 (N_6965,N_3686,N_2914);
nor U6966 (N_6966,N_3691,N_2058);
xnor U6967 (N_6967,N_4424,N_1780);
and U6968 (N_6968,N_355,N_4533);
nand U6969 (N_6969,N_3272,N_29);
xor U6970 (N_6970,N_4908,N_1260);
or U6971 (N_6971,N_4456,N_644);
and U6972 (N_6972,N_2007,N_322);
xor U6973 (N_6973,N_77,N_3980);
xnor U6974 (N_6974,N_2584,N_2339);
and U6975 (N_6975,N_3398,N_248);
xnor U6976 (N_6976,N_2136,N_132);
nor U6977 (N_6977,N_2685,N_2918);
xnor U6978 (N_6978,N_1330,N_4172);
or U6979 (N_6979,N_3837,N_3919);
nor U6980 (N_6980,N_1826,N_1716);
nand U6981 (N_6981,N_4636,N_2334);
nor U6982 (N_6982,N_4736,N_1957);
or U6983 (N_6983,N_4820,N_3674);
xnor U6984 (N_6984,N_854,N_2085);
and U6985 (N_6985,N_2300,N_3910);
xnor U6986 (N_6986,N_332,N_4103);
nor U6987 (N_6987,N_4876,N_2666);
nor U6988 (N_6988,N_2225,N_959);
nand U6989 (N_6989,N_3700,N_4646);
and U6990 (N_6990,N_2956,N_413);
nor U6991 (N_6991,N_3256,N_4412);
and U6992 (N_6992,N_2970,N_1294);
and U6993 (N_6993,N_3198,N_4878);
and U6994 (N_6994,N_2832,N_3249);
and U6995 (N_6995,N_1846,N_3754);
nor U6996 (N_6996,N_2027,N_2345);
and U6997 (N_6997,N_1582,N_1055);
nor U6998 (N_6998,N_4274,N_1693);
and U6999 (N_6999,N_761,N_975);
xor U7000 (N_7000,N_1074,N_72);
nand U7001 (N_7001,N_1802,N_4838);
nand U7002 (N_7002,N_2169,N_4836);
xor U7003 (N_7003,N_732,N_4511);
and U7004 (N_7004,N_3860,N_2198);
nand U7005 (N_7005,N_674,N_814);
nand U7006 (N_7006,N_2398,N_3499);
nand U7007 (N_7007,N_4543,N_3843);
xnor U7008 (N_7008,N_2034,N_876);
and U7009 (N_7009,N_1312,N_2777);
and U7010 (N_7010,N_4608,N_1416);
nor U7011 (N_7011,N_3,N_438);
nand U7012 (N_7012,N_3047,N_4214);
nor U7013 (N_7013,N_560,N_4145);
or U7014 (N_7014,N_1064,N_4359);
nand U7015 (N_7015,N_3611,N_4796);
nor U7016 (N_7016,N_3633,N_2138);
nand U7017 (N_7017,N_1244,N_908);
nand U7018 (N_7018,N_4429,N_619);
nand U7019 (N_7019,N_1313,N_1739);
and U7020 (N_7020,N_3363,N_2361);
or U7021 (N_7021,N_130,N_3857);
nand U7022 (N_7022,N_1370,N_2135);
nor U7023 (N_7023,N_4015,N_1360);
and U7024 (N_7024,N_4738,N_3335);
nand U7025 (N_7025,N_2038,N_2814);
and U7026 (N_7026,N_2969,N_211);
and U7027 (N_7027,N_4669,N_377);
and U7028 (N_7028,N_4508,N_1738);
and U7029 (N_7029,N_3959,N_4617);
and U7030 (N_7030,N_4366,N_809);
and U7031 (N_7031,N_1773,N_1327);
xor U7032 (N_7032,N_1221,N_4977);
nand U7033 (N_7033,N_1104,N_2386);
nor U7034 (N_7034,N_895,N_2841);
nor U7035 (N_7035,N_3760,N_1437);
xnor U7036 (N_7036,N_2373,N_889);
and U7037 (N_7037,N_2730,N_2091);
and U7038 (N_7038,N_4188,N_1132);
nand U7039 (N_7039,N_4932,N_884);
xnor U7040 (N_7040,N_3833,N_2747);
or U7041 (N_7041,N_3738,N_3465);
or U7042 (N_7042,N_2020,N_2890);
xor U7043 (N_7043,N_4628,N_3761);
nor U7044 (N_7044,N_1657,N_2201);
or U7045 (N_7045,N_754,N_2720);
nor U7046 (N_7046,N_2740,N_2128);
nand U7047 (N_7047,N_3946,N_1615);
and U7048 (N_7048,N_2047,N_3936);
xor U7049 (N_7049,N_1537,N_3512);
and U7050 (N_7050,N_1856,N_1890);
nand U7051 (N_7051,N_178,N_2056);
and U7052 (N_7052,N_3167,N_1491);
nor U7053 (N_7053,N_2445,N_1625);
and U7054 (N_7054,N_3922,N_1809);
nor U7055 (N_7055,N_824,N_4923);
or U7056 (N_7056,N_2943,N_2488);
and U7057 (N_7057,N_4487,N_3470);
xor U7058 (N_7058,N_2156,N_3472);
or U7059 (N_7059,N_4481,N_610);
or U7060 (N_7060,N_167,N_3600);
or U7061 (N_7061,N_3244,N_4381);
xnor U7062 (N_7062,N_230,N_2953);
xnor U7063 (N_7063,N_872,N_3778);
nand U7064 (N_7064,N_3541,N_4453);
and U7065 (N_7065,N_2054,N_3038);
and U7066 (N_7066,N_4510,N_4900);
or U7067 (N_7067,N_58,N_2944);
nor U7068 (N_7068,N_635,N_4463);
nand U7069 (N_7069,N_1514,N_95);
or U7070 (N_7070,N_1190,N_4727);
or U7071 (N_7071,N_3242,N_4611);
and U7072 (N_7072,N_920,N_2727);
nor U7073 (N_7073,N_321,N_1952);
or U7074 (N_7074,N_3742,N_350);
nor U7075 (N_7075,N_1503,N_4560);
and U7076 (N_7076,N_64,N_1969);
xor U7077 (N_7077,N_1620,N_3816);
xnor U7078 (N_7078,N_2812,N_2813);
nor U7079 (N_7079,N_948,N_244);
nor U7080 (N_7080,N_4356,N_856);
or U7081 (N_7081,N_2262,N_3533);
and U7082 (N_7082,N_3545,N_1815);
and U7083 (N_7083,N_3729,N_3577);
or U7084 (N_7084,N_4652,N_3142);
nand U7085 (N_7085,N_2019,N_2680);
nand U7086 (N_7086,N_4846,N_694);
or U7087 (N_7087,N_69,N_4165);
nand U7088 (N_7088,N_4553,N_2420);
xnor U7089 (N_7089,N_3297,N_2254);
xnor U7090 (N_7090,N_4410,N_4947);
and U7091 (N_7091,N_2603,N_4721);
or U7092 (N_7092,N_3547,N_3444);
nor U7093 (N_7093,N_2676,N_2972);
and U7094 (N_7094,N_1096,N_3349);
nor U7095 (N_7095,N_3049,N_4674);
nand U7096 (N_7096,N_3508,N_1935);
and U7097 (N_7097,N_1567,N_4388);
or U7098 (N_7098,N_3348,N_3156);
nand U7099 (N_7099,N_1153,N_1755);
nand U7100 (N_7100,N_1704,N_4483);
or U7101 (N_7101,N_2001,N_1804);
nor U7102 (N_7102,N_3950,N_4086);
and U7103 (N_7103,N_1774,N_4970);
xor U7104 (N_7104,N_4210,N_3932);
nand U7105 (N_7105,N_1212,N_2766);
or U7106 (N_7106,N_1162,N_31);
nor U7107 (N_7107,N_3437,N_4137);
xor U7108 (N_7108,N_4653,N_594);
xnor U7109 (N_7109,N_156,N_2259);
nor U7110 (N_7110,N_4658,N_2722);
or U7111 (N_7111,N_2570,N_1948);
and U7112 (N_7112,N_1723,N_4506);
xnor U7113 (N_7113,N_4775,N_2337);
nand U7114 (N_7114,N_1038,N_1070);
or U7115 (N_7115,N_2017,N_3253);
or U7116 (N_7116,N_693,N_4979);
or U7117 (N_7117,N_364,N_633);
xor U7118 (N_7118,N_3215,N_1842);
or U7119 (N_7119,N_4360,N_2698);
xor U7120 (N_7120,N_3114,N_3554);
and U7121 (N_7121,N_3056,N_1480);
or U7122 (N_7122,N_4835,N_4025);
or U7123 (N_7123,N_4131,N_219);
xor U7124 (N_7124,N_2741,N_4096);
nor U7125 (N_7125,N_306,N_3688);
nor U7126 (N_7126,N_747,N_530);
or U7127 (N_7127,N_4723,N_3579);
nor U7128 (N_7128,N_426,N_2712);
xnor U7129 (N_7129,N_3132,N_3109);
nor U7130 (N_7130,N_121,N_4404);
nor U7131 (N_7131,N_3482,N_2050);
xnor U7132 (N_7132,N_4622,N_308);
xnor U7133 (N_7133,N_4156,N_3513);
nor U7134 (N_7134,N_918,N_750);
nand U7135 (N_7135,N_4119,N_1655);
nand U7136 (N_7136,N_1209,N_4262);
and U7137 (N_7137,N_4812,N_3310);
nor U7138 (N_7138,N_101,N_3758);
or U7139 (N_7139,N_632,N_1635);
or U7140 (N_7140,N_1356,N_2095);
and U7141 (N_7141,N_4886,N_2836);
nor U7142 (N_7142,N_1710,N_2576);
or U7143 (N_7143,N_4709,N_3511);
or U7144 (N_7144,N_403,N_2347);
and U7145 (N_7145,N_4546,N_1035);
nor U7146 (N_7146,N_3741,N_4545);
xnor U7147 (N_7147,N_1540,N_1247);
nor U7148 (N_7148,N_2435,N_3966);
nand U7149 (N_7149,N_691,N_3231);
or U7150 (N_7150,N_3876,N_4803);
nand U7151 (N_7151,N_1531,N_2574);
or U7152 (N_7152,N_4585,N_1143);
xor U7153 (N_7153,N_2366,N_1303);
or U7154 (N_7154,N_478,N_114);
xor U7155 (N_7155,N_1552,N_682);
or U7156 (N_7156,N_216,N_864);
nor U7157 (N_7157,N_3646,N_2703);
nor U7158 (N_7158,N_3665,N_579);
nor U7159 (N_7159,N_3740,N_3434);
xor U7160 (N_7160,N_3763,N_1028);
and U7161 (N_7161,N_3952,N_2107);
or U7162 (N_7162,N_1517,N_4684);
or U7163 (N_7163,N_2090,N_425);
or U7164 (N_7164,N_400,N_1015);
nand U7165 (N_7165,N_4993,N_1795);
xor U7166 (N_7166,N_2438,N_3519);
nor U7167 (N_7167,N_4542,N_2113);
nor U7168 (N_7168,N_2500,N_1002);
xor U7169 (N_7169,N_3410,N_2429);
or U7170 (N_7170,N_3535,N_2400);
and U7171 (N_7171,N_1121,N_840);
nor U7172 (N_7172,N_3882,N_1650);
nand U7173 (N_7173,N_2872,N_1425);
xor U7174 (N_7174,N_3956,N_2555);
xnor U7175 (N_7175,N_2796,N_4498);
and U7176 (N_7176,N_1032,N_848);
nor U7177 (N_7177,N_1125,N_1272);
or U7178 (N_7178,N_4076,N_504);
nor U7179 (N_7179,N_4522,N_4544);
xor U7180 (N_7180,N_1523,N_3159);
nor U7181 (N_7181,N_4082,N_1223);
nor U7182 (N_7182,N_3963,N_1569);
nand U7183 (N_7183,N_3152,N_127);
nor U7184 (N_7184,N_337,N_3647);
nand U7185 (N_7185,N_2788,N_376);
xnor U7186 (N_7186,N_2706,N_1547);
or U7187 (N_7187,N_3781,N_1956);
and U7188 (N_7188,N_887,N_2880);
xnor U7189 (N_7189,N_115,N_2145);
nand U7190 (N_7190,N_2344,N_1977);
and U7191 (N_7191,N_3243,N_2993);
and U7192 (N_7192,N_4634,N_3300);
and U7193 (N_7193,N_294,N_981);
nand U7194 (N_7194,N_1283,N_2271);
nand U7195 (N_7195,N_4740,N_1319);
and U7196 (N_7196,N_3208,N_638);
xor U7197 (N_7197,N_763,N_800);
nand U7198 (N_7198,N_1986,N_1936);
or U7199 (N_7199,N_2348,N_917);
and U7200 (N_7200,N_3219,N_1647);
nor U7201 (N_7201,N_3430,N_4816);
and U7202 (N_7202,N_841,N_4326);
nor U7203 (N_7203,N_1365,N_1724);
nor U7204 (N_7204,N_3583,N_940);
or U7205 (N_7205,N_3783,N_4989);
nor U7206 (N_7206,N_3873,N_240);
and U7207 (N_7207,N_3894,N_41);
nand U7208 (N_7208,N_4144,N_2958);
and U7209 (N_7209,N_4562,N_1496);
nor U7210 (N_7210,N_4088,N_3320);
nand U7211 (N_7211,N_139,N_843);
nand U7212 (N_7212,N_135,N_696);
xor U7213 (N_7213,N_782,N_795);
nor U7214 (N_7214,N_307,N_2977);
xnor U7215 (N_7215,N_4872,N_1239);
nor U7216 (N_7216,N_1040,N_241);
or U7217 (N_7217,N_1690,N_2491);
xor U7218 (N_7218,N_4005,N_370);
nor U7219 (N_7219,N_1648,N_1685);
or U7220 (N_7220,N_3838,N_2092);
nor U7221 (N_7221,N_3163,N_102);
nand U7222 (N_7222,N_2086,N_2407);
nand U7223 (N_7223,N_1621,N_3082);
or U7224 (N_7224,N_3186,N_4444);
xnor U7225 (N_7225,N_4482,N_2931);
or U7226 (N_7226,N_2937,N_2869);
nor U7227 (N_7227,N_4774,N_2506);
nand U7228 (N_7228,N_1228,N_2439);
or U7229 (N_7229,N_1766,N_2342);
xor U7230 (N_7230,N_2686,N_4728);
and U7231 (N_7231,N_2260,N_2845);
and U7232 (N_7232,N_4048,N_1386);
nand U7233 (N_7233,N_3930,N_4308);
or U7234 (N_7234,N_3991,N_697);
nor U7235 (N_7235,N_3636,N_1281);
nand U7236 (N_7236,N_1812,N_591);
xor U7237 (N_7237,N_1887,N_4339);
nand U7238 (N_7238,N_52,N_4500);
nand U7239 (N_7239,N_2605,N_4879);
and U7240 (N_7240,N_4555,N_3442);
and U7241 (N_7241,N_2040,N_3423);
nand U7242 (N_7242,N_4645,N_885);
or U7243 (N_7243,N_4963,N_874);
nand U7244 (N_7244,N_1811,N_3737);
nor U7245 (N_7245,N_1987,N_1287);
and U7246 (N_7246,N_2623,N_2349);
or U7247 (N_7247,N_371,N_2122);
nand U7248 (N_7248,N_1250,N_336);
nor U7249 (N_7249,N_4863,N_880);
nand U7250 (N_7250,N_870,N_1634);
and U7251 (N_7251,N_4488,N_2161);
or U7252 (N_7252,N_3091,N_1361);
and U7253 (N_7253,N_2668,N_680);
or U7254 (N_7254,N_2888,N_4673);
nor U7255 (N_7255,N_2772,N_1838);
nand U7256 (N_7256,N_1443,N_2181);
or U7257 (N_7257,N_1359,N_353);
xnor U7258 (N_7258,N_1177,N_3370);
and U7259 (N_7259,N_3544,N_1837);
or U7260 (N_7260,N_1524,N_2179);
xnor U7261 (N_7261,N_3937,N_1411);
nand U7262 (N_7262,N_4559,N_3534);
and U7263 (N_7263,N_4138,N_1931);
nor U7264 (N_7264,N_4173,N_842);
nand U7265 (N_7265,N_4153,N_1596);
and U7266 (N_7266,N_4570,N_1001);
and U7267 (N_7267,N_3984,N_4603);
nand U7268 (N_7268,N_379,N_3312);
and U7269 (N_7269,N_4394,N_3489);
xor U7270 (N_7270,N_11,N_471);
or U7271 (N_7271,N_4665,N_398);
nand U7272 (N_7272,N_709,N_1043);
and U7273 (N_7273,N_4975,N_197);
or U7274 (N_7274,N_3137,N_3160);
nor U7275 (N_7275,N_2479,N_359);
and U7276 (N_7276,N_780,N_15);
nand U7277 (N_7277,N_2265,N_1671);
and U7278 (N_7278,N_2884,N_3904);
nand U7279 (N_7279,N_2068,N_1550);
or U7280 (N_7280,N_639,N_1897);
and U7281 (N_7281,N_268,N_1674);
xor U7282 (N_7282,N_3704,N_4777);
and U7283 (N_7283,N_2072,N_3475);
and U7284 (N_7284,N_1293,N_3199);
nand U7285 (N_7285,N_3546,N_2452);
xor U7286 (N_7286,N_4909,N_2006);
nand U7287 (N_7287,N_3419,N_4700);
or U7288 (N_7288,N_4311,N_3749);
and U7289 (N_7289,N_4120,N_475);
nor U7290 (N_7290,N_1072,N_3255);
or U7291 (N_7291,N_1,N_943);
nor U7292 (N_7292,N_1396,N_4492);
nor U7293 (N_7293,N_1335,N_4217);
xor U7294 (N_7294,N_2277,N_994);
nand U7295 (N_7295,N_3026,N_4515);
xor U7296 (N_7296,N_3753,N_393);
xnor U7297 (N_7297,N_3012,N_1220);
xnor U7298 (N_7298,N_4687,N_1061);
or U7299 (N_7299,N_968,N_1556);
xor U7300 (N_7300,N_725,N_3677);
nor U7301 (N_7301,N_2304,N_3389);
nand U7302 (N_7302,N_1963,N_1996);
nand U7303 (N_7303,N_4020,N_96);
or U7304 (N_7304,N_3969,N_3933);
or U7305 (N_7305,N_1823,N_4240);
xnor U7306 (N_7306,N_4479,N_3483);
and U7307 (N_7307,N_3810,N_1286);
and U7308 (N_7308,N_4053,N_1183);
nor U7309 (N_7309,N_549,N_2729);
or U7310 (N_7310,N_4842,N_857);
and U7311 (N_7311,N_212,N_2433);
nand U7312 (N_7312,N_3678,N_838);
xnor U7313 (N_7313,N_3817,N_792);
nand U7314 (N_7314,N_4688,N_801);
or U7315 (N_7315,N_3079,N_4666);
nor U7316 (N_7316,N_3333,N_1981);
xnor U7317 (N_7317,N_2656,N_4945);
xor U7318 (N_7318,N_70,N_3178);
and U7319 (N_7319,N_4766,N_2432);
nand U7320 (N_7320,N_280,N_161);
and U7321 (N_7321,N_1379,N_2580);
or U7322 (N_7322,N_3222,N_3750);
or U7323 (N_7323,N_1022,N_625);
nand U7324 (N_7324,N_344,N_1388);
nand U7325 (N_7325,N_1136,N_2517);
nand U7326 (N_7326,N_4278,N_93);
and U7327 (N_7327,N_1014,N_3329);
xnor U7328 (N_7328,N_3505,N_2368);
nand U7329 (N_7329,N_1682,N_3463);
nand U7330 (N_7330,N_1185,N_1516);
xnor U7331 (N_7331,N_83,N_1745);
nor U7332 (N_7332,N_1175,N_831);
xor U7333 (N_7333,N_192,N_2911);
and U7334 (N_7334,N_3110,N_4352);
or U7335 (N_7335,N_849,N_1101);
nand U7336 (N_7336,N_609,N_502);
or U7337 (N_7337,N_2096,N_4941);
xnor U7338 (N_7338,N_4307,N_1715);
or U7339 (N_7339,N_1954,N_669);
xnor U7340 (N_7340,N_3443,N_405);
nor U7341 (N_7341,N_2760,N_3259);
or U7342 (N_7342,N_2184,N_2536);
nor U7343 (N_7343,N_3395,N_3077);
nor U7344 (N_7344,N_1085,N_453);
xor U7345 (N_7345,N_4601,N_3204);
nor U7346 (N_7346,N_4465,N_1869);
and U7347 (N_7347,N_3207,N_4116);
xnor U7348 (N_7348,N_4084,N_741);
and U7349 (N_7349,N_4377,N_3532);
xor U7350 (N_7350,N_4152,N_325);
and U7351 (N_7351,N_3703,N_2650);
nor U7352 (N_7352,N_3392,N_2833);
or U7353 (N_7353,N_1060,N_2402);
and U7354 (N_7354,N_3304,N_381);
xor U7355 (N_7355,N_110,N_4303);
nand U7356 (N_7356,N_2824,N_461);
nand U7357 (N_7357,N_3261,N_3195);
nor U7358 (N_7358,N_4789,N_2421);
nor U7359 (N_7359,N_1270,N_4858);
nand U7360 (N_7360,N_3425,N_4318);
or U7361 (N_7361,N_2529,N_327);
xnor U7362 (N_7362,N_421,N_301);
and U7363 (N_7363,N_2844,N_2233);
nor U7364 (N_7364,N_3887,N_2379);
and U7365 (N_7365,N_395,N_925);
nand U7366 (N_7366,N_2883,N_3880);
and U7367 (N_7367,N_4971,N_4826);
xor U7368 (N_7368,N_2395,N_2158);
nand U7369 (N_7369,N_3550,N_4193);
nor U7370 (N_7370,N_1059,N_2241);
and U7371 (N_7371,N_2469,N_4884);
and U7372 (N_7372,N_1659,N_1769);
or U7373 (N_7373,N_4640,N_2089);
nor U7374 (N_7374,N_4925,N_464);
nor U7375 (N_7375,N_1237,N_830);
nor U7376 (N_7376,N_2647,N_3736);
or U7377 (N_7377,N_724,N_3819);
and U7378 (N_7378,N_2197,N_183);
xor U7379 (N_7379,N_1860,N_1168);
or U7380 (N_7380,N_736,N_312);
nor U7381 (N_7381,N_4194,N_2048);
nand U7382 (N_7382,N_2723,N_1345);
nand U7383 (N_7383,N_2849,N_2103);
or U7384 (N_7384,N_2102,N_1337);
or U7385 (N_7385,N_2932,N_4275);
or U7386 (N_7386,N_3835,N_962);
and U7387 (N_7387,N_1254,N_2906);
or U7388 (N_7388,N_1792,N_4734);
xnor U7389 (N_7389,N_2045,N_2231);
and U7390 (N_7390,N_2861,N_1781);
xor U7391 (N_7391,N_2399,N_4143);
nor U7392 (N_7392,N_3732,N_3592);
nand U7393 (N_7393,N_2094,N_3401);
or U7394 (N_7394,N_3097,N_2553);
and U7395 (N_7395,N_3055,N_2716);
or U7396 (N_7396,N_770,N_545);
nand U7397 (N_7397,N_3503,N_595);
or U7398 (N_7398,N_4402,N_2269);
nor U7399 (N_7399,N_4328,N_319);
or U7400 (N_7400,N_4185,N_3143);
or U7401 (N_7401,N_4358,N_1494);
nor U7402 (N_7402,N_1511,N_1643);
nor U7403 (N_7403,N_4550,N_1174);
nand U7404 (N_7404,N_4419,N_4322);
or U7405 (N_7405,N_362,N_2618);
or U7406 (N_7406,N_3229,N_2005);
or U7407 (N_7407,N_1180,N_1429);
xnor U7408 (N_7408,N_1441,N_2848);
nor U7409 (N_7409,N_1861,N_2374);
or U7410 (N_7410,N_484,N_811);
or U7411 (N_7411,N_3720,N_1213);
nor U7412 (N_7412,N_1207,N_82);
or U7413 (N_7413,N_263,N_3124);
xor U7414 (N_7414,N_1026,N_3240);
nand U7415 (N_7415,N_1081,N_2742);
and U7416 (N_7416,N_3274,N_4627);
xnor U7417 (N_7417,N_3931,N_1998);
or U7418 (N_7418,N_1394,N_3388);
xnor U7419 (N_7419,N_3228,N_4190);
xnor U7420 (N_7420,N_760,N_3520);
xnor U7421 (N_7421,N_4263,N_4161);
or U7422 (N_7422,N_794,N_4027);
nand U7423 (N_7423,N_3587,N_236);
or U7424 (N_7424,N_4431,N_612);
and U7425 (N_7425,N_1452,N_4477);
xnor U7426 (N_7426,N_1786,N_3128);
and U7427 (N_7427,N_715,N_1555);
nor U7428 (N_7428,N_4530,N_3449);
nor U7429 (N_7429,N_4447,N_4266);
or U7430 (N_7430,N_643,N_3618);
and U7431 (N_7431,N_3871,N_2463);
and U7432 (N_7432,N_3045,N_4902);
or U7433 (N_7433,N_539,N_4380);
nand U7434 (N_7434,N_275,N_3604);
xnor U7435 (N_7435,N_1482,N_2419);
and U7436 (N_7436,N_123,N_837);
or U7437 (N_7437,N_1976,N_2070);
and U7438 (N_7438,N_3619,N_4180);
nor U7439 (N_7439,N_3498,N_1454);
xor U7440 (N_7440,N_148,N_772);
xnor U7441 (N_7441,N_901,N_1691);
xnor U7442 (N_7442,N_3908,N_3202);
and U7443 (N_7443,N_2471,N_4681);
and U7444 (N_7444,N_1233,N_4004);
or U7445 (N_7445,N_4343,N_4421);
or U7446 (N_7446,N_2857,N_2592);
and U7447 (N_7447,N_1113,N_745);
xor U7448 (N_7448,N_2449,N_3981);
and U7449 (N_7449,N_4619,N_4643);
nor U7450 (N_7450,N_3979,N_3802);
nor U7451 (N_7451,N_3900,N_2149);
nor U7452 (N_7452,N_3474,N_4802);
and U7453 (N_7453,N_125,N_4801);
and U7454 (N_7454,N_2252,N_2903);
and U7455 (N_7455,N_4583,N_2462);
xor U7456 (N_7456,N_1141,N_2938);
or U7457 (N_7457,N_2415,N_550);
nand U7458 (N_7458,N_2761,N_4354);
and U7459 (N_7459,N_3416,N_2010);
and U7460 (N_7460,N_1888,N_2497);
nand U7461 (N_7461,N_2272,N_2945);
xor U7462 (N_7462,N_1091,N_3467);
and U7463 (N_7463,N_4162,N_1245);
nor U7464 (N_7464,N_3194,N_2657);
nor U7465 (N_7465,N_4155,N_1048);
xnor U7466 (N_7466,N_2125,N_877);
or U7467 (N_7467,N_865,N_339);
nor U7468 (N_7468,N_2270,N_4865);
or U7469 (N_7469,N_4304,N_1205);
xor U7470 (N_7470,N_2881,N_1158);
nor U7471 (N_7471,N_787,N_778);
or U7472 (N_7472,N_1772,N_3241);
xnor U7473 (N_7473,N_3898,N_2879);
or U7474 (N_7474,N_2293,N_927);
and U7475 (N_7475,N_768,N_154);
nor U7476 (N_7476,N_2212,N_1343);
nor U7477 (N_7477,N_2173,N_2403);
and U7478 (N_7478,N_3011,N_4426);
nor U7479 (N_7479,N_3015,N_113);
nand U7480 (N_7480,N_3023,N_983);
xnor U7481 (N_7481,N_1835,N_2992);
nor U7482 (N_7482,N_40,N_1539);
and U7483 (N_7483,N_825,N_2586);
nand U7484 (N_7484,N_4593,N_3670);
or U7485 (N_7485,N_1461,N_1490);
xor U7486 (N_7486,N_3902,N_1108);
xor U7487 (N_7487,N_2526,N_81);
nand U7488 (N_7488,N_3058,N_2933);
and U7489 (N_7489,N_4063,N_2728);
nor U7490 (N_7490,N_3526,N_4393);
and U7491 (N_7491,N_1504,N_2962);
xnor U7492 (N_7492,N_3411,N_3847);
or U7493 (N_7493,N_2130,N_2709);
nor U7494 (N_7494,N_2242,N_1505);
nand U7495 (N_7495,N_4406,N_3169);
and U7496 (N_7496,N_2214,N_731);
nor U7497 (N_7497,N_214,N_3088);
and U7498 (N_7498,N_4833,N_1864);
or U7499 (N_7499,N_2682,N_1817);
and U7500 (N_7500,N_2328,N_3297);
nand U7501 (N_7501,N_4636,N_1578);
nand U7502 (N_7502,N_4860,N_3319);
and U7503 (N_7503,N_3880,N_1145);
nor U7504 (N_7504,N_579,N_62);
xnor U7505 (N_7505,N_4122,N_1345);
or U7506 (N_7506,N_1057,N_107);
xor U7507 (N_7507,N_4338,N_4849);
or U7508 (N_7508,N_837,N_1389);
or U7509 (N_7509,N_544,N_2218);
xor U7510 (N_7510,N_4256,N_2477);
xnor U7511 (N_7511,N_2488,N_2441);
nor U7512 (N_7512,N_1845,N_3);
or U7513 (N_7513,N_3582,N_48);
nor U7514 (N_7514,N_3061,N_1993);
and U7515 (N_7515,N_4107,N_4928);
or U7516 (N_7516,N_1589,N_2596);
and U7517 (N_7517,N_214,N_1490);
nand U7518 (N_7518,N_416,N_1361);
nor U7519 (N_7519,N_2413,N_2873);
nand U7520 (N_7520,N_4718,N_4856);
xor U7521 (N_7521,N_3977,N_876);
nand U7522 (N_7522,N_775,N_4006);
and U7523 (N_7523,N_1027,N_1240);
xnor U7524 (N_7524,N_3853,N_541);
nand U7525 (N_7525,N_857,N_2400);
nand U7526 (N_7526,N_2098,N_686);
nor U7527 (N_7527,N_4128,N_3495);
and U7528 (N_7528,N_746,N_2679);
or U7529 (N_7529,N_478,N_2721);
and U7530 (N_7530,N_1502,N_1025);
or U7531 (N_7531,N_1314,N_1709);
or U7532 (N_7532,N_4398,N_4806);
nor U7533 (N_7533,N_319,N_4451);
nand U7534 (N_7534,N_2894,N_797);
nand U7535 (N_7535,N_3334,N_2036);
xor U7536 (N_7536,N_4153,N_3096);
nand U7537 (N_7537,N_4518,N_2377);
nand U7538 (N_7538,N_164,N_2444);
nor U7539 (N_7539,N_961,N_1901);
and U7540 (N_7540,N_3666,N_1146);
xor U7541 (N_7541,N_2849,N_3774);
nor U7542 (N_7542,N_2575,N_1989);
xor U7543 (N_7543,N_1399,N_2343);
nand U7544 (N_7544,N_439,N_4898);
or U7545 (N_7545,N_620,N_1880);
or U7546 (N_7546,N_1175,N_2126);
nand U7547 (N_7547,N_2362,N_4758);
xor U7548 (N_7548,N_155,N_4678);
nor U7549 (N_7549,N_2047,N_2157);
and U7550 (N_7550,N_3575,N_1558);
xor U7551 (N_7551,N_2928,N_4843);
nand U7552 (N_7552,N_1687,N_2810);
or U7553 (N_7553,N_4042,N_1758);
nor U7554 (N_7554,N_1866,N_4483);
nor U7555 (N_7555,N_1772,N_2942);
and U7556 (N_7556,N_4986,N_612);
nor U7557 (N_7557,N_4286,N_239);
and U7558 (N_7558,N_2436,N_132);
and U7559 (N_7559,N_4727,N_27);
xnor U7560 (N_7560,N_1796,N_4407);
nor U7561 (N_7561,N_3146,N_4445);
or U7562 (N_7562,N_2374,N_2944);
or U7563 (N_7563,N_1677,N_2100);
or U7564 (N_7564,N_970,N_3272);
nand U7565 (N_7565,N_4081,N_1949);
xor U7566 (N_7566,N_650,N_3683);
or U7567 (N_7567,N_4473,N_226);
and U7568 (N_7568,N_2786,N_775);
xor U7569 (N_7569,N_4874,N_1976);
xor U7570 (N_7570,N_2241,N_2506);
and U7571 (N_7571,N_1746,N_2314);
nand U7572 (N_7572,N_15,N_589);
or U7573 (N_7573,N_4028,N_3195);
nor U7574 (N_7574,N_2642,N_3231);
nand U7575 (N_7575,N_3373,N_1892);
xnor U7576 (N_7576,N_2966,N_1724);
xnor U7577 (N_7577,N_1969,N_2677);
nand U7578 (N_7578,N_4367,N_31);
nor U7579 (N_7579,N_4109,N_2082);
nor U7580 (N_7580,N_359,N_3137);
xnor U7581 (N_7581,N_186,N_48);
nor U7582 (N_7582,N_4217,N_912);
or U7583 (N_7583,N_1134,N_1811);
nand U7584 (N_7584,N_2840,N_1911);
xnor U7585 (N_7585,N_3391,N_326);
nand U7586 (N_7586,N_2305,N_1919);
nand U7587 (N_7587,N_4012,N_3952);
nor U7588 (N_7588,N_1933,N_593);
nor U7589 (N_7589,N_2021,N_1745);
and U7590 (N_7590,N_4550,N_2286);
and U7591 (N_7591,N_353,N_3068);
nand U7592 (N_7592,N_4394,N_2299);
nor U7593 (N_7593,N_4978,N_4266);
nor U7594 (N_7594,N_4611,N_2439);
nor U7595 (N_7595,N_2926,N_2064);
and U7596 (N_7596,N_3297,N_349);
nand U7597 (N_7597,N_2685,N_3870);
xor U7598 (N_7598,N_1776,N_1788);
or U7599 (N_7599,N_1519,N_2869);
nor U7600 (N_7600,N_385,N_325);
nor U7601 (N_7601,N_933,N_1932);
or U7602 (N_7602,N_4789,N_1228);
or U7603 (N_7603,N_56,N_1994);
nor U7604 (N_7604,N_4028,N_2124);
and U7605 (N_7605,N_3532,N_3056);
and U7606 (N_7606,N_149,N_1063);
xnor U7607 (N_7607,N_4048,N_2770);
or U7608 (N_7608,N_4312,N_3383);
or U7609 (N_7609,N_290,N_4589);
or U7610 (N_7610,N_197,N_4320);
or U7611 (N_7611,N_4344,N_3055);
nor U7612 (N_7612,N_1291,N_305);
or U7613 (N_7613,N_2279,N_205);
and U7614 (N_7614,N_3531,N_3890);
xor U7615 (N_7615,N_1174,N_3299);
nor U7616 (N_7616,N_2569,N_3563);
or U7617 (N_7617,N_3624,N_3100);
or U7618 (N_7618,N_3901,N_1505);
xnor U7619 (N_7619,N_2201,N_4348);
xnor U7620 (N_7620,N_3244,N_4525);
nor U7621 (N_7621,N_687,N_666);
nor U7622 (N_7622,N_4149,N_3754);
nand U7623 (N_7623,N_813,N_3725);
nor U7624 (N_7624,N_3956,N_3411);
or U7625 (N_7625,N_2019,N_2980);
nor U7626 (N_7626,N_3810,N_3697);
nand U7627 (N_7627,N_3441,N_3551);
nand U7628 (N_7628,N_1083,N_3270);
nor U7629 (N_7629,N_27,N_37);
nor U7630 (N_7630,N_2231,N_1134);
nand U7631 (N_7631,N_1917,N_2782);
or U7632 (N_7632,N_2602,N_2723);
and U7633 (N_7633,N_1234,N_4532);
or U7634 (N_7634,N_250,N_3587);
and U7635 (N_7635,N_2094,N_3140);
nand U7636 (N_7636,N_3955,N_286);
or U7637 (N_7637,N_1647,N_1182);
and U7638 (N_7638,N_2167,N_1759);
nand U7639 (N_7639,N_3359,N_501);
nor U7640 (N_7640,N_4435,N_946);
xor U7641 (N_7641,N_573,N_4441);
xor U7642 (N_7642,N_455,N_4203);
nor U7643 (N_7643,N_2472,N_4959);
or U7644 (N_7644,N_1888,N_2710);
nand U7645 (N_7645,N_1035,N_2636);
nand U7646 (N_7646,N_2603,N_2768);
or U7647 (N_7647,N_2153,N_4841);
xnor U7648 (N_7648,N_3805,N_1547);
nand U7649 (N_7649,N_3580,N_1896);
or U7650 (N_7650,N_10,N_1048);
or U7651 (N_7651,N_1620,N_3251);
and U7652 (N_7652,N_4407,N_3664);
nor U7653 (N_7653,N_2365,N_1521);
nor U7654 (N_7654,N_1908,N_4037);
xor U7655 (N_7655,N_2072,N_2937);
nor U7656 (N_7656,N_4762,N_1816);
xnor U7657 (N_7657,N_3903,N_3163);
xnor U7658 (N_7658,N_3724,N_3576);
nand U7659 (N_7659,N_2817,N_460);
xnor U7660 (N_7660,N_67,N_3315);
nand U7661 (N_7661,N_3023,N_4426);
or U7662 (N_7662,N_3631,N_743);
xor U7663 (N_7663,N_4163,N_104);
xor U7664 (N_7664,N_628,N_3921);
nand U7665 (N_7665,N_943,N_1871);
xnor U7666 (N_7666,N_779,N_2703);
xor U7667 (N_7667,N_551,N_2709);
or U7668 (N_7668,N_1210,N_3249);
xnor U7669 (N_7669,N_4922,N_1366);
and U7670 (N_7670,N_121,N_3406);
nand U7671 (N_7671,N_915,N_2152);
or U7672 (N_7672,N_3612,N_4782);
and U7673 (N_7673,N_1230,N_3029);
and U7674 (N_7674,N_443,N_1024);
or U7675 (N_7675,N_3458,N_2563);
nand U7676 (N_7676,N_1899,N_3127);
or U7677 (N_7677,N_295,N_152);
nand U7678 (N_7678,N_2138,N_468);
and U7679 (N_7679,N_1431,N_398);
and U7680 (N_7680,N_1186,N_2036);
or U7681 (N_7681,N_1831,N_1588);
xor U7682 (N_7682,N_1946,N_944);
and U7683 (N_7683,N_699,N_3572);
xor U7684 (N_7684,N_965,N_2899);
nor U7685 (N_7685,N_1741,N_3475);
and U7686 (N_7686,N_2034,N_4988);
nor U7687 (N_7687,N_823,N_4299);
nand U7688 (N_7688,N_2210,N_2056);
xnor U7689 (N_7689,N_2494,N_2379);
nor U7690 (N_7690,N_276,N_329);
xnor U7691 (N_7691,N_1105,N_2650);
nand U7692 (N_7692,N_4907,N_46);
and U7693 (N_7693,N_1180,N_1125);
nand U7694 (N_7694,N_2582,N_919);
xor U7695 (N_7695,N_1923,N_2537);
nor U7696 (N_7696,N_4179,N_4889);
xor U7697 (N_7697,N_4535,N_3661);
nor U7698 (N_7698,N_4606,N_3368);
and U7699 (N_7699,N_3899,N_1458);
nor U7700 (N_7700,N_2543,N_2459);
or U7701 (N_7701,N_652,N_3617);
nand U7702 (N_7702,N_4267,N_932);
or U7703 (N_7703,N_3644,N_2643);
nand U7704 (N_7704,N_2436,N_257);
or U7705 (N_7705,N_1300,N_3303);
or U7706 (N_7706,N_3641,N_858);
nand U7707 (N_7707,N_1303,N_1814);
nor U7708 (N_7708,N_4190,N_4315);
and U7709 (N_7709,N_268,N_687);
and U7710 (N_7710,N_1718,N_4829);
or U7711 (N_7711,N_321,N_1410);
and U7712 (N_7712,N_951,N_2256);
nor U7713 (N_7713,N_1346,N_1620);
and U7714 (N_7714,N_2224,N_4931);
xnor U7715 (N_7715,N_3886,N_1854);
or U7716 (N_7716,N_66,N_2687);
nor U7717 (N_7717,N_3322,N_4957);
xnor U7718 (N_7718,N_2649,N_69);
or U7719 (N_7719,N_4653,N_1219);
or U7720 (N_7720,N_1836,N_1793);
and U7721 (N_7721,N_2647,N_70);
and U7722 (N_7722,N_4071,N_1001);
or U7723 (N_7723,N_2859,N_4027);
xnor U7724 (N_7724,N_3395,N_4346);
nand U7725 (N_7725,N_4812,N_1060);
nor U7726 (N_7726,N_3559,N_4734);
and U7727 (N_7727,N_3180,N_37);
or U7728 (N_7728,N_1276,N_4254);
nand U7729 (N_7729,N_1961,N_1428);
and U7730 (N_7730,N_4113,N_4663);
and U7731 (N_7731,N_388,N_3308);
nand U7732 (N_7732,N_2849,N_3198);
nand U7733 (N_7733,N_3870,N_1604);
xor U7734 (N_7734,N_536,N_1729);
nand U7735 (N_7735,N_2770,N_317);
nor U7736 (N_7736,N_1720,N_2656);
or U7737 (N_7737,N_1683,N_695);
nand U7738 (N_7738,N_1341,N_1623);
and U7739 (N_7739,N_3755,N_2176);
and U7740 (N_7740,N_3094,N_3912);
nand U7741 (N_7741,N_4167,N_1910);
and U7742 (N_7742,N_1104,N_4345);
nor U7743 (N_7743,N_3064,N_4812);
nor U7744 (N_7744,N_3213,N_3504);
nor U7745 (N_7745,N_838,N_4818);
nand U7746 (N_7746,N_4070,N_1330);
nand U7747 (N_7747,N_1058,N_633);
or U7748 (N_7748,N_564,N_309);
xnor U7749 (N_7749,N_3953,N_1807);
xnor U7750 (N_7750,N_1086,N_4549);
nor U7751 (N_7751,N_4120,N_4008);
nand U7752 (N_7752,N_1756,N_3091);
nor U7753 (N_7753,N_230,N_2792);
or U7754 (N_7754,N_1758,N_3065);
or U7755 (N_7755,N_1999,N_810);
nor U7756 (N_7756,N_4799,N_1315);
and U7757 (N_7757,N_3567,N_3290);
nand U7758 (N_7758,N_3613,N_4975);
nand U7759 (N_7759,N_4208,N_2953);
nand U7760 (N_7760,N_2352,N_3217);
xnor U7761 (N_7761,N_3103,N_2475);
nand U7762 (N_7762,N_2101,N_3499);
or U7763 (N_7763,N_740,N_1678);
nor U7764 (N_7764,N_1276,N_4779);
nand U7765 (N_7765,N_3282,N_4287);
nand U7766 (N_7766,N_3230,N_2334);
or U7767 (N_7767,N_2317,N_1263);
nor U7768 (N_7768,N_3362,N_3897);
and U7769 (N_7769,N_2411,N_4428);
xnor U7770 (N_7770,N_184,N_3215);
nor U7771 (N_7771,N_765,N_3544);
or U7772 (N_7772,N_1348,N_3986);
nand U7773 (N_7773,N_3355,N_213);
or U7774 (N_7774,N_2316,N_422);
and U7775 (N_7775,N_1696,N_992);
or U7776 (N_7776,N_3555,N_972);
and U7777 (N_7777,N_3319,N_1359);
or U7778 (N_7778,N_4532,N_1871);
nor U7779 (N_7779,N_1373,N_2177);
nor U7780 (N_7780,N_3869,N_3644);
or U7781 (N_7781,N_321,N_1110);
nor U7782 (N_7782,N_2851,N_4160);
or U7783 (N_7783,N_1116,N_4513);
and U7784 (N_7784,N_27,N_4993);
and U7785 (N_7785,N_3318,N_4070);
or U7786 (N_7786,N_4514,N_3605);
and U7787 (N_7787,N_517,N_4030);
or U7788 (N_7788,N_3673,N_947);
xor U7789 (N_7789,N_4063,N_1067);
nand U7790 (N_7790,N_4779,N_3260);
nand U7791 (N_7791,N_2901,N_2282);
or U7792 (N_7792,N_2163,N_998);
xnor U7793 (N_7793,N_1052,N_149);
nor U7794 (N_7794,N_4605,N_901);
or U7795 (N_7795,N_4547,N_206);
nand U7796 (N_7796,N_450,N_731);
nand U7797 (N_7797,N_1054,N_1068);
and U7798 (N_7798,N_1132,N_2446);
nand U7799 (N_7799,N_4418,N_3792);
and U7800 (N_7800,N_247,N_2032);
and U7801 (N_7801,N_4463,N_2097);
nand U7802 (N_7802,N_3877,N_2777);
xor U7803 (N_7803,N_4634,N_156);
nand U7804 (N_7804,N_4376,N_2201);
nand U7805 (N_7805,N_4207,N_995);
xor U7806 (N_7806,N_2730,N_826);
and U7807 (N_7807,N_4245,N_994);
or U7808 (N_7808,N_292,N_1597);
or U7809 (N_7809,N_1926,N_1822);
or U7810 (N_7810,N_1213,N_2491);
xor U7811 (N_7811,N_3045,N_1911);
nor U7812 (N_7812,N_884,N_324);
nor U7813 (N_7813,N_3420,N_2770);
xor U7814 (N_7814,N_3971,N_861);
or U7815 (N_7815,N_3578,N_1973);
and U7816 (N_7816,N_3089,N_1298);
nor U7817 (N_7817,N_1964,N_993);
nor U7818 (N_7818,N_4004,N_240);
or U7819 (N_7819,N_3457,N_777);
nand U7820 (N_7820,N_4434,N_3970);
xor U7821 (N_7821,N_2382,N_3009);
and U7822 (N_7822,N_4597,N_1393);
xor U7823 (N_7823,N_280,N_496);
and U7824 (N_7824,N_3433,N_71);
nand U7825 (N_7825,N_3629,N_1310);
nor U7826 (N_7826,N_3379,N_713);
and U7827 (N_7827,N_2475,N_3796);
or U7828 (N_7828,N_3797,N_3845);
nor U7829 (N_7829,N_302,N_1082);
and U7830 (N_7830,N_2057,N_3422);
or U7831 (N_7831,N_96,N_1099);
nand U7832 (N_7832,N_1243,N_2984);
and U7833 (N_7833,N_4289,N_425);
nand U7834 (N_7834,N_374,N_3828);
and U7835 (N_7835,N_1694,N_3413);
and U7836 (N_7836,N_2802,N_3784);
and U7837 (N_7837,N_553,N_2119);
nand U7838 (N_7838,N_122,N_3744);
and U7839 (N_7839,N_2606,N_2874);
nand U7840 (N_7840,N_3225,N_97);
or U7841 (N_7841,N_3671,N_806);
and U7842 (N_7842,N_699,N_3437);
nor U7843 (N_7843,N_2279,N_2735);
or U7844 (N_7844,N_2019,N_3799);
nor U7845 (N_7845,N_3700,N_3819);
nor U7846 (N_7846,N_1385,N_4777);
nor U7847 (N_7847,N_4106,N_3293);
xor U7848 (N_7848,N_4151,N_4316);
xor U7849 (N_7849,N_3807,N_321);
or U7850 (N_7850,N_2811,N_609);
xor U7851 (N_7851,N_1635,N_3119);
xor U7852 (N_7852,N_2317,N_1153);
nand U7853 (N_7853,N_3247,N_2721);
nand U7854 (N_7854,N_2587,N_4566);
and U7855 (N_7855,N_4551,N_4616);
nor U7856 (N_7856,N_2979,N_4946);
and U7857 (N_7857,N_1164,N_3487);
nand U7858 (N_7858,N_4073,N_2494);
or U7859 (N_7859,N_3946,N_2716);
or U7860 (N_7860,N_2183,N_2023);
or U7861 (N_7861,N_4046,N_3040);
xor U7862 (N_7862,N_497,N_3792);
xnor U7863 (N_7863,N_357,N_1682);
or U7864 (N_7864,N_1431,N_2296);
and U7865 (N_7865,N_4782,N_4852);
xor U7866 (N_7866,N_2212,N_961);
nor U7867 (N_7867,N_3390,N_607);
nand U7868 (N_7868,N_3464,N_3611);
xor U7869 (N_7869,N_4809,N_3143);
xor U7870 (N_7870,N_4348,N_896);
xnor U7871 (N_7871,N_1146,N_2505);
nor U7872 (N_7872,N_3132,N_2322);
nor U7873 (N_7873,N_246,N_1211);
xnor U7874 (N_7874,N_1842,N_4898);
nand U7875 (N_7875,N_1614,N_588);
nor U7876 (N_7876,N_4920,N_2128);
and U7877 (N_7877,N_1740,N_4170);
or U7878 (N_7878,N_2052,N_3742);
and U7879 (N_7879,N_4016,N_3361);
nor U7880 (N_7880,N_138,N_778);
and U7881 (N_7881,N_3845,N_3068);
nor U7882 (N_7882,N_4411,N_3662);
nor U7883 (N_7883,N_2761,N_829);
or U7884 (N_7884,N_3287,N_4230);
xor U7885 (N_7885,N_3939,N_4690);
nand U7886 (N_7886,N_274,N_855);
xnor U7887 (N_7887,N_4353,N_2621);
and U7888 (N_7888,N_3576,N_4340);
nor U7889 (N_7889,N_2512,N_3382);
and U7890 (N_7890,N_4964,N_4710);
nand U7891 (N_7891,N_408,N_1226);
nand U7892 (N_7892,N_3072,N_3018);
or U7893 (N_7893,N_1687,N_4969);
nor U7894 (N_7894,N_2868,N_3477);
nand U7895 (N_7895,N_1824,N_1451);
nor U7896 (N_7896,N_891,N_119);
or U7897 (N_7897,N_2827,N_4760);
and U7898 (N_7898,N_2731,N_4856);
nand U7899 (N_7899,N_602,N_4799);
and U7900 (N_7900,N_2766,N_4344);
and U7901 (N_7901,N_4231,N_631);
and U7902 (N_7902,N_4355,N_325);
xnor U7903 (N_7903,N_3681,N_2839);
xnor U7904 (N_7904,N_1999,N_3481);
xnor U7905 (N_7905,N_4342,N_3756);
xor U7906 (N_7906,N_1333,N_4772);
nand U7907 (N_7907,N_2267,N_2045);
nor U7908 (N_7908,N_3320,N_1762);
nor U7909 (N_7909,N_3707,N_1570);
nand U7910 (N_7910,N_4871,N_2182);
nand U7911 (N_7911,N_138,N_4631);
or U7912 (N_7912,N_4433,N_1137);
or U7913 (N_7913,N_1375,N_2445);
nor U7914 (N_7914,N_1845,N_4982);
or U7915 (N_7915,N_3799,N_3990);
and U7916 (N_7916,N_3044,N_621);
and U7917 (N_7917,N_2720,N_2865);
nor U7918 (N_7918,N_37,N_4768);
nor U7919 (N_7919,N_2336,N_4937);
or U7920 (N_7920,N_3125,N_3720);
nor U7921 (N_7921,N_4868,N_3501);
nor U7922 (N_7922,N_1559,N_4483);
and U7923 (N_7923,N_2767,N_4224);
and U7924 (N_7924,N_1479,N_4969);
nand U7925 (N_7925,N_3136,N_1690);
and U7926 (N_7926,N_247,N_1353);
nand U7927 (N_7927,N_178,N_3560);
nand U7928 (N_7928,N_428,N_4640);
nand U7929 (N_7929,N_1176,N_2483);
and U7930 (N_7930,N_3865,N_3302);
and U7931 (N_7931,N_3667,N_3693);
nand U7932 (N_7932,N_541,N_2429);
nand U7933 (N_7933,N_302,N_243);
nand U7934 (N_7934,N_3093,N_4806);
nor U7935 (N_7935,N_1726,N_2798);
or U7936 (N_7936,N_115,N_776);
or U7937 (N_7937,N_680,N_1585);
or U7938 (N_7938,N_383,N_4040);
xor U7939 (N_7939,N_2625,N_2339);
or U7940 (N_7940,N_2267,N_248);
or U7941 (N_7941,N_3378,N_2981);
or U7942 (N_7942,N_2135,N_3999);
and U7943 (N_7943,N_1623,N_2260);
nand U7944 (N_7944,N_4950,N_676);
or U7945 (N_7945,N_998,N_4902);
nand U7946 (N_7946,N_1136,N_2299);
or U7947 (N_7947,N_128,N_1624);
nand U7948 (N_7948,N_656,N_3060);
xnor U7949 (N_7949,N_4540,N_2376);
nand U7950 (N_7950,N_419,N_3076);
xnor U7951 (N_7951,N_840,N_396);
or U7952 (N_7952,N_3780,N_4563);
or U7953 (N_7953,N_91,N_1493);
nor U7954 (N_7954,N_1601,N_1141);
xnor U7955 (N_7955,N_2069,N_878);
and U7956 (N_7956,N_4283,N_3204);
xnor U7957 (N_7957,N_650,N_1132);
and U7958 (N_7958,N_2576,N_2043);
nor U7959 (N_7959,N_1627,N_3830);
nand U7960 (N_7960,N_2744,N_3894);
and U7961 (N_7961,N_523,N_412);
nor U7962 (N_7962,N_3322,N_4844);
nor U7963 (N_7963,N_4683,N_104);
xor U7964 (N_7964,N_4074,N_4997);
nor U7965 (N_7965,N_1677,N_1163);
or U7966 (N_7966,N_3942,N_2706);
nand U7967 (N_7967,N_1124,N_349);
xnor U7968 (N_7968,N_2473,N_4833);
nor U7969 (N_7969,N_2789,N_4639);
and U7970 (N_7970,N_4400,N_350);
or U7971 (N_7971,N_574,N_1832);
nor U7972 (N_7972,N_4764,N_3330);
nor U7973 (N_7973,N_845,N_3440);
xor U7974 (N_7974,N_2234,N_1085);
and U7975 (N_7975,N_22,N_656);
nor U7976 (N_7976,N_4002,N_4728);
nand U7977 (N_7977,N_3617,N_2159);
or U7978 (N_7978,N_1663,N_2712);
or U7979 (N_7979,N_863,N_1979);
nor U7980 (N_7980,N_4247,N_3551);
nor U7981 (N_7981,N_3820,N_4068);
or U7982 (N_7982,N_2952,N_1545);
xor U7983 (N_7983,N_4214,N_1476);
and U7984 (N_7984,N_1302,N_343);
nor U7985 (N_7985,N_4298,N_3767);
nor U7986 (N_7986,N_4823,N_3355);
nor U7987 (N_7987,N_2862,N_4880);
or U7988 (N_7988,N_4931,N_450);
nor U7989 (N_7989,N_2044,N_2043);
nand U7990 (N_7990,N_2649,N_4072);
or U7991 (N_7991,N_133,N_38);
xnor U7992 (N_7992,N_4127,N_1581);
and U7993 (N_7993,N_4657,N_238);
and U7994 (N_7994,N_2917,N_2359);
and U7995 (N_7995,N_4835,N_1593);
and U7996 (N_7996,N_681,N_2357);
or U7997 (N_7997,N_1814,N_4101);
nand U7998 (N_7998,N_4285,N_1740);
xnor U7999 (N_7999,N_546,N_94);
and U8000 (N_8000,N_1278,N_4657);
nor U8001 (N_8001,N_1707,N_4856);
and U8002 (N_8002,N_2630,N_589);
nand U8003 (N_8003,N_119,N_1937);
or U8004 (N_8004,N_2716,N_114);
nor U8005 (N_8005,N_3245,N_3267);
xor U8006 (N_8006,N_2197,N_2858);
or U8007 (N_8007,N_4355,N_3812);
and U8008 (N_8008,N_3367,N_3115);
nand U8009 (N_8009,N_2208,N_3829);
nand U8010 (N_8010,N_932,N_3418);
or U8011 (N_8011,N_3301,N_3400);
and U8012 (N_8012,N_1055,N_1433);
nor U8013 (N_8013,N_1682,N_3123);
or U8014 (N_8014,N_4647,N_3169);
nor U8015 (N_8015,N_4287,N_4547);
and U8016 (N_8016,N_1778,N_985);
nor U8017 (N_8017,N_1751,N_1160);
nand U8018 (N_8018,N_1632,N_873);
nand U8019 (N_8019,N_1627,N_3872);
nand U8020 (N_8020,N_3055,N_3397);
and U8021 (N_8021,N_4179,N_1000);
xnor U8022 (N_8022,N_343,N_1685);
or U8023 (N_8023,N_1137,N_2059);
nand U8024 (N_8024,N_961,N_3539);
nand U8025 (N_8025,N_3535,N_1554);
xnor U8026 (N_8026,N_3003,N_2083);
or U8027 (N_8027,N_4906,N_1725);
and U8028 (N_8028,N_4724,N_996);
xnor U8029 (N_8029,N_414,N_4312);
nor U8030 (N_8030,N_2800,N_757);
xor U8031 (N_8031,N_4519,N_661);
nand U8032 (N_8032,N_1016,N_1701);
and U8033 (N_8033,N_1329,N_4857);
xor U8034 (N_8034,N_2124,N_3909);
or U8035 (N_8035,N_3825,N_2365);
and U8036 (N_8036,N_2483,N_970);
xor U8037 (N_8037,N_4533,N_1443);
xnor U8038 (N_8038,N_1827,N_3504);
xor U8039 (N_8039,N_2324,N_532);
or U8040 (N_8040,N_502,N_1800);
nor U8041 (N_8041,N_3181,N_616);
or U8042 (N_8042,N_2788,N_1294);
xnor U8043 (N_8043,N_358,N_1702);
nand U8044 (N_8044,N_3375,N_36);
and U8045 (N_8045,N_4441,N_1462);
nand U8046 (N_8046,N_935,N_1592);
xnor U8047 (N_8047,N_447,N_3604);
or U8048 (N_8048,N_1920,N_1236);
and U8049 (N_8049,N_3402,N_90);
xor U8050 (N_8050,N_1913,N_2530);
or U8051 (N_8051,N_2900,N_2493);
nor U8052 (N_8052,N_124,N_4156);
and U8053 (N_8053,N_3985,N_4576);
xor U8054 (N_8054,N_1820,N_4535);
nand U8055 (N_8055,N_3485,N_230);
xor U8056 (N_8056,N_3559,N_2614);
xnor U8057 (N_8057,N_760,N_4192);
xnor U8058 (N_8058,N_2159,N_1288);
or U8059 (N_8059,N_3170,N_125);
nand U8060 (N_8060,N_985,N_1126);
nand U8061 (N_8061,N_4692,N_4031);
and U8062 (N_8062,N_444,N_3857);
xnor U8063 (N_8063,N_3145,N_1766);
and U8064 (N_8064,N_1683,N_3791);
and U8065 (N_8065,N_4267,N_3593);
nor U8066 (N_8066,N_4593,N_737);
nor U8067 (N_8067,N_1238,N_1709);
or U8068 (N_8068,N_648,N_1245);
or U8069 (N_8069,N_1819,N_3485);
or U8070 (N_8070,N_4088,N_1961);
nor U8071 (N_8071,N_4989,N_4791);
nor U8072 (N_8072,N_4911,N_4028);
xor U8073 (N_8073,N_1394,N_1537);
and U8074 (N_8074,N_1676,N_2496);
xor U8075 (N_8075,N_2350,N_4347);
or U8076 (N_8076,N_3457,N_4942);
and U8077 (N_8077,N_925,N_4625);
and U8078 (N_8078,N_2686,N_4454);
or U8079 (N_8079,N_3136,N_363);
and U8080 (N_8080,N_4978,N_1797);
and U8081 (N_8081,N_2082,N_4871);
or U8082 (N_8082,N_1262,N_226);
xnor U8083 (N_8083,N_4678,N_2035);
nor U8084 (N_8084,N_96,N_4202);
or U8085 (N_8085,N_1767,N_4545);
or U8086 (N_8086,N_3684,N_2648);
and U8087 (N_8087,N_1307,N_4946);
nor U8088 (N_8088,N_4589,N_205);
nor U8089 (N_8089,N_4110,N_4700);
xor U8090 (N_8090,N_2220,N_3095);
nand U8091 (N_8091,N_4745,N_4806);
or U8092 (N_8092,N_2459,N_4369);
nand U8093 (N_8093,N_429,N_484);
xor U8094 (N_8094,N_2709,N_2378);
nand U8095 (N_8095,N_3662,N_1714);
and U8096 (N_8096,N_4210,N_2671);
nand U8097 (N_8097,N_974,N_4661);
xnor U8098 (N_8098,N_73,N_2424);
or U8099 (N_8099,N_3951,N_1100);
or U8100 (N_8100,N_2879,N_4185);
nor U8101 (N_8101,N_742,N_1093);
xnor U8102 (N_8102,N_4801,N_2552);
and U8103 (N_8103,N_1425,N_3229);
xnor U8104 (N_8104,N_3958,N_147);
nor U8105 (N_8105,N_4735,N_2209);
xor U8106 (N_8106,N_1832,N_4971);
xnor U8107 (N_8107,N_4303,N_1611);
nand U8108 (N_8108,N_2704,N_3978);
or U8109 (N_8109,N_2355,N_1393);
nor U8110 (N_8110,N_1047,N_3166);
nand U8111 (N_8111,N_540,N_3840);
nand U8112 (N_8112,N_2037,N_171);
xnor U8113 (N_8113,N_4317,N_1324);
nand U8114 (N_8114,N_866,N_4814);
or U8115 (N_8115,N_1826,N_4863);
and U8116 (N_8116,N_2916,N_1704);
nand U8117 (N_8117,N_1973,N_1785);
xnor U8118 (N_8118,N_1541,N_602);
and U8119 (N_8119,N_3151,N_4399);
xnor U8120 (N_8120,N_510,N_1875);
and U8121 (N_8121,N_476,N_4681);
and U8122 (N_8122,N_9,N_2656);
and U8123 (N_8123,N_4045,N_579);
nor U8124 (N_8124,N_1952,N_4923);
nand U8125 (N_8125,N_287,N_1427);
nor U8126 (N_8126,N_4399,N_2023);
xor U8127 (N_8127,N_4211,N_1549);
or U8128 (N_8128,N_1774,N_3902);
and U8129 (N_8129,N_4172,N_2878);
nor U8130 (N_8130,N_2942,N_1100);
or U8131 (N_8131,N_3019,N_4687);
or U8132 (N_8132,N_1004,N_1885);
nand U8133 (N_8133,N_510,N_3973);
nand U8134 (N_8134,N_4544,N_4091);
nand U8135 (N_8135,N_2475,N_2780);
nand U8136 (N_8136,N_3039,N_2197);
and U8137 (N_8137,N_3292,N_4104);
nor U8138 (N_8138,N_4262,N_1142);
and U8139 (N_8139,N_2002,N_4023);
nand U8140 (N_8140,N_1848,N_1846);
xnor U8141 (N_8141,N_3180,N_1928);
nor U8142 (N_8142,N_4216,N_3672);
nor U8143 (N_8143,N_4438,N_2262);
and U8144 (N_8144,N_2195,N_3308);
nor U8145 (N_8145,N_3462,N_4918);
or U8146 (N_8146,N_111,N_3490);
or U8147 (N_8147,N_3034,N_4420);
nand U8148 (N_8148,N_1189,N_1146);
nand U8149 (N_8149,N_3051,N_2967);
nor U8150 (N_8150,N_3228,N_3262);
nor U8151 (N_8151,N_1276,N_2278);
xnor U8152 (N_8152,N_2398,N_4725);
and U8153 (N_8153,N_236,N_4196);
nand U8154 (N_8154,N_3613,N_1169);
and U8155 (N_8155,N_775,N_86);
and U8156 (N_8156,N_2270,N_2932);
nand U8157 (N_8157,N_120,N_915);
nor U8158 (N_8158,N_2806,N_2214);
and U8159 (N_8159,N_825,N_3239);
and U8160 (N_8160,N_4405,N_3126);
xnor U8161 (N_8161,N_37,N_4510);
nand U8162 (N_8162,N_4593,N_1137);
nor U8163 (N_8163,N_2071,N_435);
nand U8164 (N_8164,N_3646,N_4096);
nand U8165 (N_8165,N_1436,N_4998);
xor U8166 (N_8166,N_4659,N_1573);
and U8167 (N_8167,N_143,N_654);
or U8168 (N_8168,N_1292,N_1241);
nand U8169 (N_8169,N_2234,N_2332);
and U8170 (N_8170,N_3569,N_896);
and U8171 (N_8171,N_3355,N_1196);
or U8172 (N_8172,N_3727,N_4659);
and U8173 (N_8173,N_912,N_3301);
and U8174 (N_8174,N_923,N_3867);
and U8175 (N_8175,N_990,N_210);
or U8176 (N_8176,N_4248,N_2851);
nor U8177 (N_8177,N_4266,N_1757);
nand U8178 (N_8178,N_1767,N_3904);
nor U8179 (N_8179,N_77,N_921);
xor U8180 (N_8180,N_775,N_1577);
xnor U8181 (N_8181,N_274,N_3370);
or U8182 (N_8182,N_163,N_1292);
xor U8183 (N_8183,N_1214,N_4734);
nand U8184 (N_8184,N_3596,N_4933);
xnor U8185 (N_8185,N_4184,N_10);
or U8186 (N_8186,N_654,N_0);
xnor U8187 (N_8187,N_4351,N_2149);
nand U8188 (N_8188,N_288,N_2227);
xnor U8189 (N_8189,N_3612,N_1672);
or U8190 (N_8190,N_3047,N_479);
and U8191 (N_8191,N_336,N_1721);
nand U8192 (N_8192,N_3605,N_4671);
and U8193 (N_8193,N_2027,N_3843);
and U8194 (N_8194,N_4965,N_4425);
xnor U8195 (N_8195,N_2082,N_2397);
xnor U8196 (N_8196,N_1808,N_4371);
and U8197 (N_8197,N_1044,N_4211);
xor U8198 (N_8198,N_1962,N_1556);
xor U8199 (N_8199,N_2087,N_3274);
or U8200 (N_8200,N_3071,N_4902);
nand U8201 (N_8201,N_4237,N_1512);
and U8202 (N_8202,N_3279,N_1366);
xnor U8203 (N_8203,N_4378,N_3146);
nand U8204 (N_8204,N_1700,N_813);
nand U8205 (N_8205,N_4722,N_24);
or U8206 (N_8206,N_4901,N_1397);
nor U8207 (N_8207,N_4390,N_1457);
nand U8208 (N_8208,N_2945,N_3398);
nor U8209 (N_8209,N_2063,N_4617);
and U8210 (N_8210,N_4269,N_782);
xnor U8211 (N_8211,N_1897,N_793);
nor U8212 (N_8212,N_403,N_3651);
or U8213 (N_8213,N_3376,N_3703);
nand U8214 (N_8214,N_283,N_488);
and U8215 (N_8215,N_281,N_1346);
xnor U8216 (N_8216,N_194,N_69);
or U8217 (N_8217,N_350,N_2936);
and U8218 (N_8218,N_4848,N_4567);
or U8219 (N_8219,N_840,N_3418);
nor U8220 (N_8220,N_3680,N_3475);
xor U8221 (N_8221,N_849,N_4782);
nand U8222 (N_8222,N_3485,N_2111);
or U8223 (N_8223,N_4247,N_3810);
nand U8224 (N_8224,N_3554,N_2860);
nand U8225 (N_8225,N_4792,N_1732);
or U8226 (N_8226,N_282,N_967);
nor U8227 (N_8227,N_279,N_1214);
and U8228 (N_8228,N_2189,N_1849);
or U8229 (N_8229,N_4537,N_4701);
nor U8230 (N_8230,N_2790,N_1443);
nor U8231 (N_8231,N_3458,N_1661);
nor U8232 (N_8232,N_2907,N_3789);
nand U8233 (N_8233,N_4144,N_3638);
and U8234 (N_8234,N_2309,N_4741);
or U8235 (N_8235,N_4684,N_260);
nor U8236 (N_8236,N_3684,N_865);
or U8237 (N_8237,N_1682,N_4171);
xor U8238 (N_8238,N_261,N_250);
xor U8239 (N_8239,N_439,N_3756);
nor U8240 (N_8240,N_1021,N_3881);
and U8241 (N_8241,N_1450,N_2512);
nand U8242 (N_8242,N_3820,N_4748);
nor U8243 (N_8243,N_898,N_2100);
or U8244 (N_8244,N_726,N_4249);
nand U8245 (N_8245,N_567,N_733);
or U8246 (N_8246,N_3481,N_1422);
and U8247 (N_8247,N_3876,N_4592);
and U8248 (N_8248,N_4776,N_460);
and U8249 (N_8249,N_3240,N_2874);
nand U8250 (N_8250,N_1738,N_4402);
nand U8251 (N_8251,N_2637,N_1574);
nand U8252 (N_8252,N_4806,N_123);
or U8253 (N_8253,N_831,N_1854);
xor U8254 (N_8254,N_3387,N_2245);
xor U8255 (N_8255,N_1963,N_1341);
nand U8256 (N_8256,N_1224,N_2768);
nor U8257 (N_8257,N_4378,N_2287);
or U8258 (N_8258,N_2604,N_720);
nor U8259 (N_8259,N_185,N_4015);
or U8260 (N_8260,N_1935,N_1217);
and U8261 (N_8261,N_2539,N_4346);
xnor U8262 (N_8262,N_1800,N_853);
xor U8263 (N_8263,N_1104,N_2437);
and U8264 (N_8264,N_939,N_3941);
xor U8265 (N_8265,N_493,N_905);
xnor U8266 (N_8266,N_1158,N_3524);
xnor U8267 (N_8267,N_1146,N_2958);
xor U8268 (N_8268,N_3710,N_2193);
and U8269 (N_8269,N_4115,N_1856);
or U8270 (N_8270,N_1527,N_2799);
nor U8271 (N_8271,N_3743,N_4237);
or U8272 (N_8272,N_4473,N_2008);
nor U8273 (N_8273,N_1380,N_303);
and U8274 (N_8274,N_4103,N_3540);
xnor U8275 (N_8275,N_4064,N_2412);
nand U8276 (N_8276,N_2326,N_186);
and U8277 (N_8277,N_1898,N_3764);
and U8278 (N_8278,N_2303,N_2096);
or U8279 (N_8279,N_3847,N_459);
or U8280 (N_8280,N_273,N_2213);
xor U8281 (N_8281,N_4110,N_4785);
nand U8282 (N_8282,N_1989,N_1096);
nor U8283 (N_8283,N_1890,N_102);
nand U8284 (N_8284,N_2529,N_1485);
xnor U8285 (N_8285,N_3241,N_4929);
nor U8286 (N_8286,N_4870,N_100);
and U8287 (N_8287,N_1164,N_3298);
and U8288 (N_8288,N_4043,N_595);
xnor U8289 (N_8289,N_1306,N_151);
xnor U8290 (N_8290,N_2179,N_4670);
nor U8291 (N_8291,N_3410,N_1771);
or U8292 (N_8292,N_4123,N_4393);
nor U8293 (N_8293,N_4062,N_4718);
nor U8294 (N_8294,N_2451,N_1293);
and U8295 (N_8295,N_1743,N_3489);
xor U8296 (N_8296,N_98,N_2681);
or U8297 (N_8297,N_2997,N_2597);
and U8298 (N_8298,N_1995,N_1970);
or U8299 (N_8299,N_973,N_2109);
xor U8300 (N_8300,N_1838,N_2560);
nand U8301 (N_8301,N_4996,N_3802);
and U8302 (N_8302,N_2505,N_1156);
or U8303 (N_8303,N_3139,N_2910);
and U8304 (N_8304,N_1952,N_29);
nand U8305 (N_8305,N_2127,N_2813);
and U8306 (N_8306,N_3434,N_2709);
xor U8307 (N_8307,N_1594,N_2681);
xor U8308 (N_8308,N_2667,N_2397);
or U8309 (N_8309,N_1384,N_430);
or U8310 (N_8310,N_1882,N_1782);
nand U8311 (N_8311,N_2674,N_3522);
nand U8312 (N_8312,N_768,N_3627);
nor U8313 (N_8313,N_4582,N_2141);
or U8314 (N_8314,N_271,N_4516);
nor U8315 (N_8315,N_49,N_307);
xnor U8316 (N_8316,N_1199,N_1711);
or U8317 (N_8317,N_146,N_3711);
or U8318 (N_8318,N_1233,N_4542);
nor U8319 (N_8319,N_1559,N_1673);
nor U8320 (N_8320,N_4795,N_3139);
or U8321 (N_8321,N_3843,N_3862);
nand U8322 (N_8322,N_3145,N_4567);
or U8323 (N_8323,N_2084,N_375);
xnor U8324 (N_8324,N_597,N_807);
nand U8325 (N_8325,N_478,N_1017);
nor U8326 (N_8326,N_3672,N_4637);
or U8327 (N_8327,N_179,N_285);
or U8328 (N_8328,N_3036,N_4622);
and U8329 (N_8329,N_2177,N_2357);
or U8330 (N_8330,N_1053,N_4411);
xor U8331 (N_8331,N_1458,N_4286);
nand U8332 (N_8332,N_4382,N_2922);
or U8333 (N_8333,N_1677,N_2645);
or U8334 (N_8334,N_4513,N_1278);
or U8335 (N_8335,N_4005,N_3843);
nand U8336 (N_8336,N_227,N_1342);
and U8337 (N_8337,N_2626,N_2839);
xnor U8338 (N_8338,N_3348,N_1768);
nor U8339 (N_8339,N_304,N_3106);
nand U8340 (N_8340,N_2198,N_3027);
nor U8341 (N_8341,N_4073,N_2691);
or U8342 (N_8342,N_4815,N_3186);
or U8343 (N_8343,N_3415,N_3816);
nand U8344 (N_8344,N_4447,N_4101);
nand U8345 (N_8345,N_2956,N_1877);
nand U8346 (N_8346,N_2241,N_2264);
xor U8347 (N_8347,N_1149,N_654);
nor U8348 (N_8348,N_4468,N_1657);
or U8349 (N_8349,N_417,N_1910);
nor U8350 (N_8350,N_1651,N_2206);
nor U8351 (N_8351,N_2378,N_2332);
xor U8352 (N_8352,N_4766,N_3908);
and U8353 (N_8353,N_3260,N_214);
and U8354 (N_8354,N_2232,N_272);
and U8355 (N_8355,N_1502,N_1872);
nand U8356 (N_8356,N_3022,N_1810);
nor U8357 (N_8357,N_3083,N_4330);
nor U8358 (N_8358,N_3343,N_3707);
xor U8359 (N_8359,N_3422,N_1459);
nand U8360 (N_8360,N_2488,N_2692);
xor U8361 (N_8361,N_4110,N_2018);
xnor U8362 (N_8362,N_774,N_1108);
nand U8363 (N_8363,N_2803,N_998);
xor U8364 (N_8364,N_369,N_1531);
nand U8365 (N_8365,N_782,N_2235);
or U8366 (N_8366,N_208,N_1880);
or U8367 (N_8367,N_3365,N_3335);
xor U8368 (N_8368,N_3319,N_3583);
or U8369 (N_8369,N_734,N_4948);
nor U8370 (N_8370,N_1231,N_2054);
nor U8371 (N_8371,N_3992,N_4387);
nand U8372 (N_8372,N_835,N_3836);
nand U8373 (N_8373,N_1738,N_99);
xnor U8374 (N_8374,N_3162,N_2441);
nor U8375 (N_8375,N_3626,N_184);
xor U8376 (N_8376,N_2848,N_4828);
or U8377 (N_8377,N_1731,N_2295);
xor U8378 (N_8378,N_2379,N_1795);
xor U8379 (N_8379,N_676,N_3108);
or U8380 (N_8380,N_4317,N_2145);
or U8381 (N_8381,N_452,N_3661);
xor U8382 (N_8382,N_326,N_1542);
or U8383 (N_8383,N_2664,N_4324);
nor U8384 (N_8384,N_2414,N_1607);
nand U8385 (N_8385,N_2962,N_2760);
nand U8386 (N_8386,N_2450,N_531);
nand U8387 (N_8387,N_3825,N_2792);
or U8388 (N_8388,N_1063,N_1869);
xnor U8389 (N_8389,N_550,N_3475);
nand U8390 (N_8390,N_4983,N_2497);
nand U8391 (N_8391,N_2977,N_2720);
xor U8392 (N_8392,N_3651,N_4887);
xor U8393 (N_8393,N_2655,N_1913);
or U8394 (N_8394,N_324,N_3215);
xor U8395 (N_8395,N_1254,N_608);
nor U8396 (N_8396,N_59,N_3944);
nor U8397 (N_8397,N_4600,N_4233);
nor U8398 (N_8398,N_2655,N_2018);
or U8399 (N_8399,N_3812,N_998);
xnor U8400 (N_8400,N_1872,N_2174);
and U8401 (N_8401,N_1611,N_3036);
and U8402 (N_8402,N_437,N_654);
nand U8403 (N_8403,N_1919,N_1490);
or U8404 (N_8404,N_542,N_3740);
nor U8405 (N_8405,N_856,N_4130);
nor U8406 (N_8406,N_2994,N_4581);
nor U8407 (N_8407,N_1915,N_4564);
xor U8408 (N_8408,N_1460,N_2999);
and U8409 (N_8409,N_429,N_502);
xor U8410 (N_8410,N_903,N_4390);
xor U8411 (N_8411,N_1810,N_4745);
nand U8412 (N_8412,N_1292,N_769);
xor U8413 (N_8413,N_3708,N_1615);
nand U8414 (N_8414,N_4198,N_1815);
or U8415 (N_8415,N_2976,N_4562);
and U8416 (N_8416,N_410,N_1415);
nor U8417 (N_8417,N_577,N_2321);
nor U8418 (N_8418,N_4617,N_1102);
and U8419 (N_8419,N_3000,N_3998);
and U8420 (N_8420,N_805,N_4885);
xor U8421 (N_8421,N_353,N_1959);
nand U8422 (N_8422,N_4358,N_693);
or U8423 (N_8423,N_2157,N_2256);
nor U8424 (N_8424,N_2530,N_59);
xor U8425 (N_8425,N_2412,N_1517);
xnor U8426 (N_8426,N_1959,N_2927);
nand U8427 (N_8427,N_140,N_956);
nand U8428 (N_8428,N_4087,N_1460);
or U8429 (N_8429,N_1489,N_2968);
nor U8430 (N_8430,N_539,N_4641);
nand U8431 (N_8431,N_3860,N_1937);
xor U8432 (N_8432,N_4946,N_2634);
nand U8433 (N_8433,N_3415,N_2558);
or U8434 (N_8434,N_3374,N_3342);
xnor U8435 (N_8435,N_4470,N_4145);
or U8436 (N_8436,N_4718,N_1730);
and U8437 (N_8437,N_2463,N_4806);
nor U8438 (N_8438,N_3867,N_1352);
xor U8439 (N_8439,N_4272,N_4636);
nor U8440 (N_8440,N_1988,N_4413);
xnor U8441 (N_8441,N_4981,N_1055);
nand U8442 (N_8442,N_1181,N_4393);
nand U8443 (N_8443,N_4786,N_958);
nand U8444 (N_8444,N_3993,N_4513);
and U8445 (N_8445,N_3873,N_568);
nor U8446 (N_8446,N_3299,N_2430);
nand U8447 (N_8447,N_2032,N_3234);
nand U8448 (N_8448,N_2841,N_3803);
and U8449 (N_8449,N_1794,N_3716);
xor U8450 (N_8450,N_2380,N_335);
or U8451 (N_8451,N_1108,N_4330);
nor U8452 (N_8452,N_1290,N_1634);
and U8453 (N_8453,N_2546,N_1196);
nor U8454 (N_8454,N_184,N_3982);
nand U8455 (N_8455,N_2039,N_1918);
or U8456 (N_8456,N_2041,N_2316);
nor U8457 (N_8457,N_990,N_916);
or U8458 (N_8458,N_432,N_2050);
or U8459 (N_8459,N_451,N_4166);
xor U8460 (N_8460,N_2760,N_4349);
and U8461 (N_8461,N_1680,N_2231);
or U8462 (N_8462,N_1115,N_2758);
or U8463 (N_8463,N_455,N_1690);
xor U8464 (N_8464,N_4163,N_1352);
xnor U8465 (N_8465,N_4695,N_925);
or U8466 (N_8466,N_2464,N_4120);
xnor U8467 (N_8467,N_4214,N_3218);
nand U8468 (N_8468,N_808,N_1914);
nand U8469 (N_8469,N_1751,N_3528);
nand U8470 (N_8470,N_4682,N_1278);
and U8471 (N_8471,N_651,N_3011);
and U8472 (N_8472,N_1829,N_1949);
nor U8473 (N_8473,N_2516,N_2677);
nand U8474 (N_8474,N_1827,N_3619);
nor U8475 (N_8475,N_2814,N_2495);
and U8476 (N_8476,N_1970,N_2582);
and U8477 (N_8477,N_2184,N_1400);
and U8478 (N_8478,N_2579,N_4729);
nand U8479 (N_8479,N_757,N_1830);
nor U8480 (N_8480,N_2514,N_1204);
or U8481 (N_8481,N_1773,N_1007);
or U8482 (N_8482,N_2794,N_1336);
xnor U8483 (N_8483,N_1382,N_2169);
nor U8484 (N_8484,N_4504,N_1636);
nand U8485 (N_8485,N_4828,N_1537);
or U8486 (N_8486,N_4430,N_3418);
or U8487 (N_8487,N_3430,N_4347);
nor U8488 (N_8488,N_3027,N_1783);
xnor U8489 (N_8489,N_2817,N_816);
and U8490 (N_8490,N_760,N_2420);
xor U8491 (N_8491,N_2288,N_3263);
and U8492 (N_8492,N_122,N_1508);
nand U8493 (N_8493,N_2181,N_2825);
and U8494 (N_8494,N_4552,N_4542);
and U8495 (N_8495,N_2681,N_1077);
xnor U8496 (N_8496,N_2009,N_298);
and U8497 (N_8497,N_2495,N_2370);
or U8498 (N_8498,N_832,N_1014);
xor U8499 (N_8499,N_290,N_3821);
and U8500 (N_8500,N_2426,N_1270);
nor U8501 (N_8501,N_3899,N_4740);
nand U8502 (N_8502,N_541,N_2699);
nand U8503 (N_8503,N_874,N_3917);
xor U8504 (N_8504,N_2378,N_3931);
nor U8505 (N_8505,N_4370,N_3496);
or U8506 (N_8506,N_2357,N_1774);
and U8507 (N_8507,N_863,N_340);
or U8508 (N_8508,N_73,N_3394);
nand U8509 (N_8509,N_995,N_3480);
nor U8510 (N_8510,N_4318,N_2045);
xnor U8511 (N_8511,N_1355,N_2483);
and U8512 (N_8512,N_989,N_4659);
nor U8513 (N_8513,N_4130,N_3488);
or U8514 (N_8514,N_4126,N_1054);
nand U8515 (N_8515,N_751,N_54);
xnor U8516 (N_8516,N_27,N_4287);
nand U8517 (N_8517,N_3844,N_4069);
nand U8518 (N_8518,N_1915,N_1766);
or U8519 (N_8519,N_28,N_207);
xnor U8520 (N_8520,N_1525,N_302);
nand U8521 (N_8521,N_4868,N_2866);
xor U8522 (N_8522,N_3505,N_1928);
or U8523 (N_8523,N_1612,N_4552);
xor U8524 (N_8524,N_1012,N_1595);
and U8525 (N_8525,N_3331,N_2480);
xor U8526 (N_8526,N_2214,N_1885);
nand U8527 (N_8527,N_1915,N_2037);
or U8528 (N_8528,N_4055,N_1859);
nand U8529 (N_8529,N_4357,N_641);
nand U8530 (N_8530,N_3488,N_4883);
xor U8531 (N_8531,N_1811,N_1980);
and U8532 (N_8532,N_3482,N_4760);
nor U8533 (N_8533,N_3273,N_4203);
and U8534 (N_8534,N_4507,N_1608);
nor U8535 (N_8535,N_80,N_1463);
nand U8536 (N_8536,N_3537,N_2349);
nand U8537 (N_8537,N_3817,N_4863);
and U8538 (N_8538,N_355,N_4659);
xor U8539 (N_8539,N_2732,N_4926);
xnor U8540 (N_8540,N_2478,N_3143);
xnor U8541 (N_8541,N_3125,N_660);
or U8542 (N_8542,N_2124,N_2902);
nor U8543 (N_8543,N_4174,N_936);
nand U8544 (N_8544,N_2485,N_1549);
and U8545 (N_8545,N_1895,N_570);
and U8546 (N_8546,N_3512,N_4943);
or U8547 (N_8547,N_4571,N_4795);
xnor U8548 (N_8548,N_4743,N_4049);
xor U8549 (N_8549,N_2712,N_3106);
xnor U8550 (N_8550,N_1904,N_2380);
nor U8551 (N_8551,N_3715,N_3540);
nand U8552 (N_8552,N_2147,N_263);
nand U8553 (N_8553,N_2706,N_3478);
and U8554 (N_8554,N_834,N_400);
nor U8555 (N_8555,N_4489,N_3001);
nand U8556 (N_8556,N_1034,N_2031);
or U8557 (N_8557,N_1921,N_1426);
or U8558 (N_8558,N_1959,N_4858);
or U8559 (N_8559,N_2209,N_1697);
and U8560 (N_8560,N_2607,N_957);
and U8561 (N_8561,N_1056,N_2539);
nor U8562 (N_8562,N_506,N_337);
or U8563 (N_8563,N_1839,N_3733);
and U8564 (N_8564,N_981,N_2779);
or U8565 (N_8565,N_3538,N_996);
or U8566 (N_8566,N_1691,N_4048);
nor U8567 (N_8567,N_1831,N_3359);
nand U8568 (N_8568,N_2941,N_579);
xor U8569 (N_8569,N_2818,N_335);
and U8570 (N_8570,N_4805,N_392);
xnor U8571 (N_8571,N_1787,N_4437);
and U8572 (N_8572,N_3001,N_695);
and U8573 (N_8573,N_2741,N_2708);
and U8574 (N_8574,N_4615,N_1370);
xnor U8575 (N_8575,N_1127,N_3618);
xor U8576 (N_8576,N_2062,N_4145);
or U8577 (N_8577,N_1116,N_2958);
nor U8578 (N_8578,N_3376,N_3660);
and U8579 (N_8579,N_215,N_814);
nand U8580 (N_8580,N_1476,N_1168);
or U8581 (N_8581,N_4987,N_4668);
or U8582 (N_8582,N_492,N_1626);
xor U8583 (N_8583,N_2019,N_2375);
nand U8584 (N_8584,N_3288,N_985);
xnor U8585 (N_8585,N_2073,N_481);
nor U8586 (N_8586,N_3342,N_1131);
nand U8587 (N_8587,N_1760,N_3404);
xnor U8588 (N_8588,N_1037,N_3501);
or U8589 (N_8589,N_1807,N_4434);
and U8590 (N_8590,N_4700,N_316);
xnor U8591 (N_8591,N_2141,N_1240);
xnor U8592 (N_8592,N_3558,N_996);
and U8593 (N_8593,N_1036,N_3103);
nor U8594 (N_8594,N_3050,N_3105);
or U8595 (N_8595,N_1820,N_4490);
xnor U8596 (N_8596,N_459,N_1494);
nand U8597 (N_8597,N_1163,N_3430);
or U8598 (N_8598,N_297,N_4355);
nor U8599 (N_8599,N_178,N_3907);
nand U8600 (N_8600,N_528,N_2629);
and U8601 (N_8601,N_1483,N_4855);
and U8602 (N_8602,N_1410,N_4016);
and U8603 (N_8603,N_3227,N_3628);
nand U8604 (N_8604,N_403,N_3771);
nor U8605 (N_8605,N_1169,N_3545);
xor U8606 (N_8606,N_4829,N_1771);
and U8607 (N_8607,N_274,N_987);
and U8608 (N_8608,N_1671,N_2447);
nor U8609 (N_8609,N_2736,N_2448);
xor U8610 (N_8610,N_3334,N_267);
nor U8611 (N_8611,N_225,N_1091);
nand U8612 (N_8612,N_3309,N_4463);
xor U8613 (N_8613,N_1735,N_4605);
and U8614 (N_8614,N_1058,N_1548);
xnor U8615 (N_8615,N_2441,N_4152);
and U8616 (N_8616,N_3668,N_3897);
nand U8617 (N_8617,N_3520,N_2285);
nor U8618 (N_8618,N_3659,N_4723);
nand U8619 (N_8619,N_2636,N_1865);
and U8620 (N_8620,N_4372,N_4436);
nor U8621 (N_8621,N_3958,N_1295);
xor U8622 (N_8622,N_1668,N_763);
or U8623 (N_8623,N_182,N_947);
or U8624 (N_8624,N_979,N_3074);
and U8625 (N_8625,N_534,N_4133);
nor U8626 (N_8626,N_1460,N_3934);
and U8627 (N_8627,N_4297,N_21);
or U8628 (N_8628,N_1863,N_554);
and U8629 (N_8629,N_1153,N_166);
and U8630 (N_8630,N_2339,N_2068);
nand U8631 (N_8631,N_3383,N_1296);
xor U8632 (N_8632,N_2855,N_4602);
xor U8633 (N_8633,N_3399,N_1230);
xor U8634 (N_8634,N_2211,N_444);
nand U8635 (N_8635,N_2481,N_3242);
nor U8636 (N_8636,N_2963,N_2493);
nand U8637 (N_8637,N_3120,N_839);
xor U8638 (N_8638,N_104,N_485);
nor U8639 (N_8639,N_4839,N_691);
xnor U8640 (N_8640,N_4226,N_2713);
xnor U8641 (N_8641,N_522,N_3139);
nand U8642 (N_8642,N_626,N_1014);
and U8643 (N_8643,N_2803,N_4377);
xor U8644 (N_8644,N_4927,N_836);
nor U8645 (N_8645,N_1748,N_3650);
xor U8646 (N_8646,N_2693,N_3844);
nand U8647 (N_8647,N_857,N_454);
or U8648 (N_8648,N_1971,N_2484);
nand U8649 (N_8649,N_487,N_1471);
nor U8650 (N_8650,N_1735,N_4410);
nor U8651 (N_8651,N_4742,N_2159);
or U8652 (N_8652,N_540,N_4128);
and U8653 (N_8653,N_3579,N_4722);
nor U8654 (N_8654,N_66,N_2811);
and U8655 (N_8655,N_1899,N_2101);
and U8656 (N_8656,N_996,N_2651);
nor U8657 (N_8657,N_64,N_2104);
nand U8658 (N_8658,N_711,N_406);
xnor U8659 (N_8659,N_1080,N_2157);
nand U8660 (N_8660,N_2704,N_4247);
nand U8661 (N_8661,N_533,N_4191);
and U8662 (N_8662,N_213,N_1246);
or U8663 (N_8663,N_1665,N_1266);
nor U8664 (N_8664,N_4534,N_2216);
xnor U8665 (N_8665,N_1324,N_1778);
or U8666 (N_8666,N_3668,N_1620);
xnor U8667 (N_8667,N_680,N_2372);
and U8668 (N_8668,N_3203,N_114);
nand U8669 (N_8669,N_2266,N_81);
or U8670 (N_8670,N_1735,N_2342);
nand U8671 (N_8671,N_2769,N_2200);
and U8672 (N_8672,N_3425,N_4169);
nand U8673 (N_8673,N_1044,N_747);
and U8674 (N_8674,N_636,N_4198);
or U8675 (N_8675,N_89,N_4899);
xor U8676 (N_8676,N_20,N_64);
nor U8677 (N_8677,N_4719,N_4876);
nor U8678 (N_8678,N_2108,N_2014);
and U8679 (N_8679,N_2800,N_2906);
nand U8680 (N_8680,N_3393,N_2704);
or U8681 (N_8681,N_393,N_1813);
and U8682 (N_8682,N_1866,N_120);
and U8683 (N_8683,N_1309,N_3758);
nand U8684 (N_8684,N_2646,N_3355);
nand U8685 (N_8685,N_3614,N_3548);
and U8686 (N_8686,N_4096,N_1208);
xnor U8687 (N_8687,N_187,N_1768);
or U8688 (N_8688,N_1702,N_4686);
and U8689 (N_8689,N_1091,N_1896);
nor U8690 (N_8690,N_904,N_1544);
and U8691 (N_8691,N_2492,N_4707);
xor U8692 (N_8692,N_974,N_1524);
and U8693 (N_8693,N_4772,N_3585);
nand U8694 (N_8694,N_4899,N_3100);
and U8695 (N_8695,N_4256,N_3237);
nand U8696 (N_8696,N_834,N_4062);
xor U8697 (N_8697,N_767,N_2148);
nand U8698 (N_8698,N_1342,N_4343);
xor U8699 (N_8699,N_3131,N_799);
or U8700 (N_8700,N_2233,N_3697);
nor U8701 (N_8701,N_1872,N_2330);
and U8702 (N_8702,N_1202,N_1354);
nor U8703 (N_8703,N_1814,N_833);
nor U8704 (N_8704,N_4319,N_2191);
and U8705 (N_8705,N_3491,N_978);
xor U8706 (N_8706,N_4713,N_4749);
and U8707 (N_8707,N_3171,N_2047);
nand U8708 (N_8708,N_1295,N_897);
nor U8709 (N_8709,N_2975,N_1019);
xnor U8710 (N_8710,N_2740,N_3321);
xnor U8711 (N_8711,N_4390,N_3277);
or U8712 (N_8712,N_1504,N_4009);
xnor U8713 (N_8713,N_2944,N_4306);
and U8714 (N_8714,N_3796,N_4688);
nand U8715 (N_8715,N_618,N_253);
nand U8716 (N_8716,N_4837,N_2714);
and U8717 (N_8717,N_3433,N_245);
nand U8718 (N_8718,N_1284,N_3032);
nand U8719 (N_8719,N_3923,N_4502);
or U8720 (N_8720,N_3186,N_1307);
xor U8721 (N_8721,N_388,N_3872);
nand U8722 (N_8722,N_3467,N_4291);
xor U8723 (N_8723,N_2412,N_3818);
nor U8724 (N_8724,N_2361,N_4610);
xor U8725 (N_8725,N_529,N_1131);
xnor U8726 (N_8726,N_3437,N_2339);
xnor U8727 (N_8727,N_2752,N_2395);
nand U8728 (N_8728,N_3866,N_3267);
and U8729 (N_8729,N_4415,N_2746);
nor U8730 (N_8730,N_832,N_2876);
nand U8731 (N_8731,N_3659,N_3257);
nor U8732 (N_8732,N_226,N_2877);
and U8733 (N_8733,N_242,N_3943);
nand U8734 (N_8734,N_1940,N_1641);
nor U8735 (N_8735,N_1508,N_4540);
and U8736 (N_8736,N_4561,N_4525);
and U8737 (N_8737,N_3596,N_486);
nand U8738 (N_8738,N_3180,N_2835);
xor U8739 (N_8739,N_4294,N_4745);
or U8740 (N_8740,N_381,N_303);
nand U8741 (N_8741,N_1409,N_4356);
or U8742 (N_8742,N_563,N_3118);
nor U8743 (N_8743,N_3727,N_3921);
and U8744 (N_8744,N_3158,N_2151);
or U8745 (N_8745,N_4399,N_1322);
and U8746 (N_8746,N_1975,N_1403);
and U8747 (N_8747,N_3183,N_3252);
nor U8748 (N_8748,N_1585,N_2708);
xor U8749 (N_8749,N_4825,N_380);
or U8750 (N_8750,N_4910,N_2097);
and U8751 (N_8751,N_4432,N_2583);
and U8752 (N_8752,N_1671,N_4536);
nand U8753 (N_8753,N_2659,N_2465);
xnor U8754 (N_8754,N_1103,N_107);
or U8755 (N_8755,N_756,N_3687);
nor U8756 (N_8756,N_233,N_2867);
nor U8757 (N_8757,N_1714,N_1639);
and U8758 (N_8758,N_919,N_3375);
and U8759 (N_8759,N_1735,N_4473);
xnor U8760 (N_8760,N_2688,N_4711);
or U8761 (N_8761,N_2349,N_4743);
and U8762 (N_8762,N_1822,N_133);
nor U8763 (N_8763,N_4136,N_2626);
xor U8764 (N_8764,N_1277,N_1891);
and U8765 (N_8765,N_689,N_2669);
and U8766 (N_8766,N_1557,N_3923);
and U8767 (N_8767,N_842,N_4830);
or U8768 (N_8768,N_4956,N_1419);
nor U8769 (N_8769,N_794,N_932);
nand U8770 (N_8770,N_4933,N_4639);
or U8771 (N_8771,N_2029,N_272);
and U8772 (N_8772,N_930,N_266);
nor U8773 (N_8773,N_781,N_1320);
or U8774 (N_8774,N_4502,N_164);
nand U8775 (N_8775,N_3010,N_3539);
nand U8776 (N_8776,N_897,N_3360);
and U8777 (N_8777,N_859,N_2202);
nor U8778 (N_8778,N_3041,N_2370);
or U8779 (N_8779,N_2089,N_1151);
xor U8780 (N_8780,N_1537,N_4086);
or U8781 (N_8781,N_4473,N_2260);
nor U8782 (N_8782,N_3137,N_4616);
and U8783 (N_8783,N_105,N_3114);
xnor U8784 (N_8784,N_2833,N_1126);
or U8785 (N_8785,N_2082,N_844);
and U8786 (N_8786,N_4153,N_3773);
nor U8787 (N_8787,N_2764,N_4008);
nor U8788 (N_8788,N_1780,N_3966);
and U8789 (N_8789,N_4007,N_958);
nor U8790 (N_8790,N_1467,N_2038);
nor U8791 (N_8791,N_1541,N_1308);
or U8792 (N_8792,N_798,N_986);
or U8793 (N_8793,N_812,N_804);
nand U8794 (N_8794,N_1386,N_4351);
nand U8795 (N_8795,N_568,N_4931);
and U8796 (N_8796,N_1161,N_4736);
nor U8797 (N_8797,N_3650,N_4921);
nor U8798 (N_8798,N_4196,N_1035);
nor U8799 (N_8799,N_1203,N_182);
xnor U8800 (N_8800,N_4286,N_4259);
or U8801 (N_8801,N_73,N_4501);
and U8802 (N_8802,N_4310,N_869);
xnor U8803 (N_8803,N_4754,N_4404);
nor U8804 (N_8804,N_1663,N_694);
nand U8805 (N_8805,N_2131,N_3621);
and U8806 (N_8806,N_1885,N_1787);
nand U8807 (N_8807,N_4548,N_1634);
or U8808 (N_8808,N_3872,N_2009);
xor U8809 (N_8809,N_103,N_995);
nor U8810 (N_8810,N_146,N_0);
or U8811 (N_8811,N_3646,N_3951);
or U8812 (N_8812,N_4103,N_1932);
or U8813 (N_8813,N_3808,N_3224);
and U8814 (N_8814,N_3292,N_1723);
xor U8815 (N_8815,N_4161,N_1480);
xor U8816 (N_8816,N_3306,N_4229);
or U8817 (N_8817,N_1570,N_2884);
xor U8818 (N_8818,N_2917,N_2661);
and U8819 (N_8819,N_4949,N_1324);
nor U8820 (N_8820,N_1912,N_38);
or U8821 (N_8821,N_1758,N_3428);
or U8822 (N_8822,N_3687,N_1092);
nor U8823 (N_8823,N_789,N_3752);
or U8824 (N_8824,N_1983,N_1796);
nand U8825 (N_8825,N_1344,N_2936);
xnor U8826 (N_8826,N_3377,N_4936);
nor U8827 (N_8827,N_4881,N_3929);
or U8828 (N_8828,N_1982,N_4034);
xnor U8829 (N_8829,N_556,N_2400);
and U8830 (N_8830,N_385,N_4277);
and U8831 (N_8831,N_369,N_2217);
nor U8832 (N_8832,N_4670,N_3565);
and U8833 (N_8833,N_3809,N_3040);
nand U8834 (N_8834,N_1493,N_3560);
xor U8835 (N_8835,N_1429,N_2663);
or U8836 (N_8836,N_248,N_4002);
and U8837 (N_8837,N_35,N_2198);
nand U8838 (N_8838,N_3760,N_1242);
nand U8839 (N_8839,N_4651,N_2588);
nor U8840 (N_8840,N_3242,N_3989);
and U8841 (N_8841,N_917,N_2987);
xnor U8842 (N_8842,N_717,N_83);
and U8843 (N_8843,N_2352,N_4724);
nor U8844 (N_8844,N_4628,N_3158);
or U8845 (N_8845,N_3907,N_1585);
nand U8846 (N_8846,N_84,N_1987);
nand U8847 (N_8847,N_1061,N_3505);
or U8848 (N_8848,N_1479,N_3660);
nand U8849 (N_8849,N_1085,N_4317);
nor U8850 (N_8850,N_2222,N_1280);
nor U8851 (N_8851,N_755,N_456);
nor U8852 (N_8852,N_1162,N_3353);
xnor U8853 (N_8853,N_2325,N_3911);
and U8854 (N_8854,N_4888,N_2191);
nor U8855 (N_8855,N_3659,N_3837);
or U8856 (N_8856,N_4697,N_2836);
or U8857 (N_8857,N_3335,N_3043);
nand U8858 (N_8858,N_3046,N_3217);
nand U8859 (N_8859,N_1575,N_4243);
nand U8860 (N_8860,N_4315,N_3842);
nor U8861 (N_8861,N_4480,N_3091);
nand U8862 (N_8862,N_2335,N_2446);
and U8863 (N_8863,N_3076,N_1395);
nor U8864 (N_8864,N_2294,N_4365);
nand U8865 (N_8865,N_1492,N_662);
xnor U8866 (N_8866,N_1802,N_3109);
nand U8867 (N_8867,N_2535,N_4192);
and U8868 (N_8868,N_895,N_790);
nand U8869 (N_8869,N_3551,N_3475);
or U8870 (N_8870,N_1948,N_3680);
xnor U8871 (N_8871,N_4722,N_1717);
nand U8872 (N_8872,N_4485,N_116);
or U8873 (N_8873,N_1696,N_4971);
nand U8874 (N_8874,N_237,N_1998);
or U8875 (N_8875,N_3773,N_3508);
nand U8876 (N_8876,N_675,N_4607);
and U8877 (N_8877,N_279,N_4897);
nor U8878 (N_8878,N_3136,N_3071);
xor U8879 (N_8879,N_2411,N_2856);
xor U8880 (N_8880,N_3780,N_1228);
nor U8881 (N_8881,N_1607,N_1398);
nand U8882 (N_8882,N_2464,N_1881);
and U8883 (N_8883,N_3991,N_4987);
and U8884 (N_8884,N_4365,N_1165);
and U8885 (N_8885,N_4504,N_4106);
or U8886 (N_8886,N_4055,N_1985);
nor U8887 (N_8887,N_1136,N_4418);
or U8888 (N_8888,N_2659,N_4987);
nor U8889 (N_8889,N_4825,N_3650);
nor U8890 (N_8890,N_897,N_4344);
or U8891 (N_8891,N_1969,N_1110);
xnor U8892 (N_8892,N_4461,N_1143);
or U8893 (N_8893,N_3725,N_4931);
and U8894 (N_8894,N_2109,N_3290);
or U8895 (N_8895,N_3588,N_1313);
and U8896 (N_8896,N_3520,N_975);
and U8897 (N_8897,N_4953,N_329);
and U8898 (N_8898,N_4207,N_4417);
xnor U8899 (N_8899,N_4627,N_2063);
nor U8900 (N_8900,N_3326,N_1894);
nand U8901 (N_8901,N_3743,N_728);
and U8902 (N_8902,N_2167,N_2170);
and U8903 (N_8903,N_1684,N_3673);
nand U8904 (N_8904,N_3777,N_2366);
xor U8905 (N_8905,N_4302,N_4049);
nor U8906 (N_8906,N_4782,N_3363);
nand U8907 (N_8907,N_2621,N_4468);
nand U8908 (N_8908,N_4641,N_4984);
or U8909 (N_8909,N_3245,N_2522);
nor U8910 (N_8910,N_16,N_4818);
nor U8911 (N_8911,N_4579,N_509);
nor U8912 (N_8912,N_4061,N_3492);
xor U8913 (N_8913,N_1789,N_2784);
nand U8914 (N_8914,N_3225,N_3280);
nor U8915 (N_8915,N_3988,N_4270);
xnor U8916 (N_8916,N_2131,N_4619);
and U8917 (N_8917,N_4322,N_4711);
and U8918 (N_8918,N_4996,N_4876);
xor U8919 (N_8919,N_2443,N_185);
or U8920 (N_8920,N_4857,N_4680);
or U8921 (N_8921,N_64,N_557);
xor U8922 (N_8922,N_4249,N_2350);
nor U8923 (N_8923,N_3896,N_1384);
nor U8924 (N_8924,N_3340,N_1533);
nand U8925 (N_8925,N_2742,N_2074);
nor U8926 (N_8926,N_2286,N_4368);
nor U8927 (N_8927,N_4619,N_2021);
nor U8928 (N_8928,N_802,N_4805);
xor U8929 (N_8929,N_2917,N_315);
and U8930 (N_8930,N_4387,N_383);
or U8931 (N_8931,N_1878,N_3360);
nor U8932 (N_8932,N_3959,N_4174);
nor U8933 (N_8933,N_274,N_3973);
xor U8934 (N_8934,N_4892,N_3921);
nand U8935 (N_8935,N_1158,N_4772);
and U8936 (N_8936,N_2352,N_1395);
and U8937 (N_8937,N_2572,N_3031);
nor U8938 (N_8938,N_396,N_1738);
xnor U8939 (N_8939,N_4074,N_4829);
and U8940 (N_8940,N_1311,N_2684);
and U8941 (N_8941,N_1130,N_4832);
and U8942 (N_8942,N_4506,N_835);
and U8943 (N_8943,N_2230,N_4212);
or U8944 (N_8944,N_3853,N_2909);
or U8945 (N_8945,N_2564,N_4594);
and U8946 (N_8946,N_1966,N_3805);
xor U8947 (N_8947,N_1914,N_855);
xor U8948 (N_8948,N_126,N_3132);
or U8949 (N_8949,N_4318,N_4333);
xnor U8950 (N_8950,N_3852,N_2508);
and U8951 (N_8951,N_1497,N_4559);
nor U8952 (N_8952,N_2482,N_1657);
nor U8953 (N_8953,N_3543,N_1005);
and U8954 (N_8954,N_2233,N_2091);
xnor U8955 (N_8955,N_1889,N_3072);
nand U8956 (N_8956,N_4693,N_4334);
xnor U8957 (N_8957,N_4432,N_2238);
nor U8958 (N_8958,N_930,N_1240);
nand U8959 (N_8959,N_64,N_335);
xnor U8960 (N_8960,N_2701,N_1683);
xor U8961 (N_8961,N_3354,N_102);
or U8962 (N_8962,N_2738,N_2305);
xor U8963 (N_8963,N_85,N_1328);
and U8964 (N_8964,N_4031,N_2919);
xnor U8965 (N_8965,N_4571,N_4993);
nor U8966 (N_8966,N_1976,N_4602);
nor U8967 (N_8967,N_88,N_1699);
or U8968 (N_8968,N_258,N_3289);
or U8969 (N_8969,N_37,N_669);
xnor U8970 (N_8970,N_2419,N_671);
or U8971 (N_8971,N_2083,N_1998);
or U8972 (N_8972,N_4629,N_1825);
xor U8973 (N_8973,N_690,N_3228);
xor U8974 (N_8974,N_2605,N_3213);
nand U8975 (N_8975,N_4885,N_2902);
or U8976 (N_8976,N_2384,N_3666);
xnor U8977 (N_8977,N_3420,N_4352);
or U8978 (N_8978,N_3834,N_770);
xor U8979 (N_8979,N_3586,N_3218);
nand U8980 (N_8980,N_71,N_2895);
nand U8981 (N_8981,N_4102,N_4898);
and U8982 (N_8982,N_2972,N_1397);
xnor U8983 (N_8983,N_2560,N_399);
nand U8984 (N_8984,N_525,N_1373);
xor U8985 (N_8985,N_272,N_3510);
xor U8986 (N_8986,N_2747,N_1618);
nor U8987 (N_8987,N_2581,N_2013);
and U8988 (N_8988,N_3287,N_3218);
xnor U8989 (N_8989,N_3332,N_3381);
xnor U8990 (N_8990,N_1827,N_2668);
or U8991 (N_8991,N_2795,N_2624);
or U8992 (N_8992,N_355,N_4554);
or U8993 (N_8993,N_2072,N_4956);
nand U8994 (N_8994,N_4823,N_2953);
nor U8995 (N_8995,N_198,N_1551);
nor U8996 (N_8996,N_1528,N_2485);
nand U8997 (N_8997,N_1693,N_45);
xnor U8998 (N_8998,N_2493,N_853);
nor U8999 (N_8999,N_299,N_719);
or U9000 (N_9000,N_2963,N_4127);
and U9001 (N_9001,N_1929,N_2583);
nor U9002 (N_9002,N_4194,N_1345);
or U9003 (N_9003,N_1112,N_3409);
or U9004 (N_9004,N_1874,N_962);
xnor U9005 (N_9005,N_155,N_4982);
nand U9006 (N_9006,N_4442,N_2161);
or U9007 (N_9007,N_675,N_531);
nand U9008 (N_9008,N_204,N_4405);
xor U9009 (N_9009,N_54,N_1140);
nand U9010 (N_9010,N_3298,N_3039);
nor U9011 (N_9011,N_3131,N_1862);
xor U9012 (N_9012,N_4060,N_4399);
nor U9013 (N_9013,N_3624,N_1206);
nor U9014 (N_9014,N_4903,N_4293);
or U9015 (N_9015,N_2950,N_4175);
nor U9016 (N_9016,N_2950,N_3939);
and U9017 (N_9017,N_3895,N_1853);
nand U9018 (N_9018,N_307,N_1793);
nand U9019 (N_9019,N_852,N_4011);
nor U9020 (N_9020,N_350,N_3040);
nor U9021 (N_9021,N_2691,N_4681);
nand U9022 (N_9022,N_1870,N_19);
or U9023 (N_9023,N_4081,N_879);
xor U9024 (N_9024,N_3011,N_2539);
nand U9025 (N_9025,N_2056,N_3782);
or U9026 (N_9026,N_3955,N_4988);
xnor U9027 (N_9027,N_2377,N_2385);
xor U9028 (N_9028,N_3376,N_2306);
and U9029 (N_9029,N_1506,N_2867);
and U9030 (N_9030,N_4381,N_4962);
and U9031 (N_9031,N_373,N_1141);
xnor U9032 (N_9032,N_3343,N_4492);
nor U9033 (N_9033,N_1095,N_3468);
xnor U9034 (N_9034,N_3049,N_4319);
nor U9035 (N_9035,N_2270,N_11);
nor U9036 (N_9036,N_3423,N_66);
nand U9037 (N_9037,N_3414,N_4963);
and U9038 (N_9038,N_619,N_891);
nor U9039 (N_9039,N_2542,N_3482);
or U9040 (N_9040,N_4182,N_1328);
and U9041 (N_9041,N_1474,N_1179);
xnor U9042 (N_9042,N_194,N_4272);
or U9043 (N_9043,N_2848,N_1365);
or U9044 (N_9044,N_4262,N_4482);
xor U9045 (N_9045,N_2432,N_3861);
xnor U9046 (N_9046,N_1225,N_4646);
nand U9047 (N_9047,N_3863,N_1319);
xor U9048 (N_9048,N_194,N_4554);
nand U9049 (N_9049,N_1848,N_4767);
xor U9050 (N_9050,N_1286,N_4779);
nand U9051 (N_9051,N_203,N_260);
or U9052 (N_9052,N_316,N_1378);
nor U9053 (N_9053,N_2593,N_4652);
nor U9054 (N_9054,N_1468,N_1889);
nand U9055 (N_9055,N_3210,N_2665);
or U9056 (N_9056,N_2837,N_4603);
or U9057 (N_9057,N_383,N_33);
xor U9058 (N_9058,N_176,N_4494);
nand U9059 (N_9059,N_4539,N_4504);
and U9060 (N_9060,N_799,N_3100);
or U9061 (N_9061,N_228,N_2259);
or U9062 (N_9062,N_2337,N_3065);
nor U9063 (N_9063,N_3857,N_3952);
or U9064 (N_9064,N_2904,N_1180);
xnor U9065 (N_9065,N_4470,N_3000);
or U9066 (N_9066,N_4791,N_3011);
or U9067 (N_9067,N_2522,N_1511);
nand U9068 (N_9068,N_1907,N_3278);
nand U9069 (N_9069,N_2036,N_1587);
nand U9070 (N_9070,N_1695,N_4339);
xor U9071 (N_9071,N_278,N_4498);
xnor U9072 (N_9072,N_4039,N_1776);
or U9073 (N_9073,N_76,N_458);
xor U9074 (N_9074,N_1705,N_1122);
or U9075 (N_9075,N_2948,N_631);
nand U9076 (N_9076,N_267,N_2901);
or U9077 (N_9077,N_3780,N_1705);
xor U9078 (N_9078,N_3243,N_1248);
or U9079 (N_9079,N_635,N_4137);
xnor U9080 (N_9080,N_552,N_4273);
nor U9081 (N_9081,N_3415,N_4367);
nand U9082 (N_9082,N_4761,N_89);
xor U9083 (N_9083,N_848,N_1122);
and U9084 (N_9084,N_3730,N_705);
nor U9085 (N_9085,N_233,N_4556);
xnor U9086 (N_9086,N_1107,N_658);
nand U9087 (N_9087,N_3727,N_109);
and U9088 (N_9088,N_4166,N_1331);
xor U9089 (N_9089,N_4066,N_2777);
nor U9090 (N_9090,N_1666,N_1920);
or U9091 (N_9091,N_2574,N_1075);
nand U9092 (N_9092,N_882,N_543);
nor U9093 (N_9093,N_753,N_4489);
xnor U9094 (N_9094,N_3371,N_4512);
and U9095 (N_9095,N_615,N_4809);
nand U9096 (N_9096,N_1793,N_2401);
xor U9097 (N_9097,N_2121,N_4183);
or U9098 (N_9098,N_1320,N_2639);
and U9099 (N_9099,N_1036,N_567);
and U9100 (N_9100,N_4435,N_1442);
and U9101 (N_9101,N_614,N_3225);
xor U9102 (N_9102,N_3156,N_3146);
nand U9103 (N_9103,N_3550,N_4541);
nor U9104 (N_9104,N_133,N_1276);
xnor U9105 (N_9105,N_1915,N_3116);
or U9106 (N_9106,N_4891,N_140);
nand U9107 (N_9107,N_342,N_2554);
xor U9108 (N_9108,N_2011,N_98);
nor U9109 (N_9109,N_4933,N_3572);
and U9110 (N_9110,N_440,N_2028);
xnor U9111 (N_9111,N_192,N_4701);
xor U9112 (N_9112,N_970,N_2790);
and U9113 (N_9113,N_2309,N_3303);
nand U9114 (N_9114,N_3344,N_436);
xor U9115 (N_9115,N_2586,N_2285);
nor U9116 (N_9116,N_1681,N_2776);
nor U9117 (N_9117,N_2893,N_913);
xnor U9118 (N_9118,N_3496,N_2501);
and U9119 (N_9119,N_3402,N_4030);
and U9120 (N_9120,N_1202,N_3389);
nor U9121 (N_9121,N_3025,N_705);
and U9122 (N_9122,N_2703,N_3673);
nor U9123 (N_9123,N_4476,N_1499);
nor U9124 (N_9124,N_3341,N_4848);
and U9125 (N_9125,N_1537,N_1824);
nor U9126 (N_9126,N_4130,N_4965);
xnor U9127 (N_9127,N_1893,N_3932);
or U9128 (N_9128,N_4103,N_2810);
and U9129 (N_9129,N_4412,N_1105);
nor U9130 (N_9130,N_1512,N_1280);
and U9131 (N_9131,N_2742,N_3032);
and U9132 (N_9132,N_4589,N_3059);
nand U9133 (N_9133,N_3063,N_4335);
xnor U9134 (N_9134,N_536,N_4773);
and U9135 (N_9135,N_3897,N_359);
nand U9136 (N_9136,N_1211,N_894);
nor U9137 (N_9137,N_3982,N_3744);
and U9138 (N_9138,N_237,N_4762);
nor U9139 (N_9139,N_2409,N_4023);
nor U9140 (N_9140,N_4926,N_367);
xnor U9141 (N_9141,N_3302,N_455);
or U9142 (N_9142,N_3861,N_488);
nand U9143 (N_9143,N_3283,N_4816);
and U9144 (N_9144,N_2725,N_2902);
nor U9145 (N_9145,N_4334,N_3189);
or U9146 (N_9146,N_1083,N_3953);
xor U9147 (N_9147,N_4437,N_1206);
nand U9148 (N_9148,N_4942,N_921);
nor U9149 (N_9149,N_669,N_1959);
xnor U9150 (N_9150,N_2523,N_125);
nand U9151 (N_9151,N_4874,N_1986);
nand U9152 (N_9152,N_3633,N_2314);
xor U9153 (N_9153,N_2309,N_1514);
and U9154 (N_9154,N_1699,N_1819);
nor U9155 (N_9155,N_3172,N_2373);
and U9156 (N_9156,N_3470,N_2056);
xnor U9157 (N_9157,N_602,N_1466);
or U9158 (N_9158,N_2383,N_4387);
xor U9159 (N_9159,N_1880,N_4017);
and U9160 (N_9160,N_3143,N_185);
xor U9161 (N_9161,N_2158,N_409);
xor U9162 (N_9162,N_3273,N_3470);
nor U9163 (N_9163,N_3861,N_2091);
nand U9164 (N_9164,N_1108,N_1607);
or U9165 (N_9165,N_576,N_4850);
and U9166 (N_9166,N_305,N_4398);
xnor U9167 (N_9167,N_3797,N_2036);
nand U9168 (N_9168,N_1075,N_1713);
or U9169 (N_9169,N_4969,N_2871);
nor U9170 (N_9170,N_2063,N_3126);
xnor U9171 (N_9171,N_3596,N_714);
nor U9172 (N_9172,N_2264,N_3838);
or U9173 (N_9173,N_2469,N_3772);
nand U9174 (N_9174,N_3947,N_2399);
or U9175 (N_9175,N_2042,N_141);
xor U9176 (N_9176,N_111,N_3119);
and U9177 (N_9177,N_3916,N_4808);
xnor U9178 (N_9178,N_2354,N_4833);
xor U9179 (N_9179,N_1731,N_2303);
and U9180 (N_9180,N_1022,N_153);
nor U9181 (N_9181,N_391,N_2487);
and U9182 (N_9182,N_4252,N_3961);
nand U9183 (N_9183,N_1231,N_947);
and U9184 (N_9184,N_4365,N_1944);
and U9185 (N_9185,N_3543,N_1427);
nand U9186 (N_9186,N_343,N_975);
nor U9187 (N_9187,N_386,N_2634);
nand U9188 (N_9188,N_3116,N_3263);
and U9189 (N_9189,N_4557,N_922);
nor U9190 (N_9190,N_208,N_980);
nand U9191 (N_9191,N_2353,N_561);
nand U9192 (N_9192,N_4651,N_472);
nand U9193 (N_9193,N_3745,N_4519);
nand U9194 (N_9194,N_4286,N_4599);
or U9195 (N_9195,N_714,N_889);
or U9196 (N_9196,N_1623,N_2359);
and U9197 (N_9197,N_4938,N_251);
nor U9198 (N_9198,N_4988,N_4703);
and U9199 (N_9199,N_1102,N_1874);
nor U9200 (N_9200,N_3392,N_780);
and U9201 (N_9201,N_1880,N_3329);
or U9202 (N_9202,N_4690,N_1207);
nand U9203 (N_9203,N_3751,N_3110);
nor U9204 (N_9204,N_858,N_4650);
xnor U9205 (N_9205,N_4077,N_1775);
nor U9206 (N_9206,N_203,N_1532);
xnor U9207 (N_9207,N_1669,N_3866);
nand U9208 (N_9208,N_4936,N_620);
nand U9209 (N_9209,N_4413,N_708);
xor U9210 (N_9210,N_3704,N_4321);
nor U9211 (N_9211,N_2040,N_4212);
nand U9212 (N_9212,N_4227,N_3341);
or U9213 (N_9213,N_2470,N_2312);
nor U9214 (N_9214,N_1128,N_4220);
nand U9215 (N_9215,N_1742,N_1287);
and U9216 (N_9216,N_3262,N_4677);
nor U9217 (N_9217,N_4946,N_442);
or U9218 (N_9218,N_4926,N_2311);
or U9219 (N_9219,N_4688,N_3836);
xor U9220 (N_9220,N_4850,N_1743);
and U9221 (N_9221,N_3731,N_948);
nand U9222 (N_9222,N_3448,N_3017);
nand U9223 (N_9223,N_2811,N_1673);
or U9224 (N_9224,N_2387,N_1871);
nand U9225 (N_9225,N_2806,N_4192);
and U9226 (N_9226,N_2736,N_926);
and U9227 (N_9227,N_3219,N_4728);
nor U9228 (N_9228,N_1013,N_104);
nor U9229 (N_9229,N_4578,N_3316);
and U9230 (N_9230,N_4410,N_2223);
or U9231 (N_9231,N_753,N_3180);
nand U9232 (N_9232,N_1190,N_3624);
or U9233 (N_9233,N_3758,N_2256);
nand U9234 (N_9234,N_3170,N_3638);
xor U9235 (N_9235,N_1401,N_2513);
or U9236 (N_9236,N_3760,N_4314);
and U9237 (N_9237,N_4576,N_539);
and U9238 (N_9238,N_2758,N_2705);
or U9239 (N_9239,N_2473,N_521);
xnor U9240 (N_9240,N_1160,N_3069);
nor U9241 (N_9241,N_1379,N_3577);
xor U9242 (N_9242,N_2343,N_3628);
xnor U9243 (N_9243,N_70,N_2534);
nand U9244 (N_9244,N_4237,N_3313);
and U9245 (N_9245,N_2865,N_136);
nor U9246 (N_9246,N_3975,N_2599);
nand U9247 (N_9247,N_2882,N_4823);
nor U9248 (N_9248,N_1268,N_4555);
nor U9249 (N_9249,N_1276,N_958);
xor U9250 (N_9250,N_3408,N_4069);
and U9251 (N_9251,N_1702,N_1669);
xor U9252 (N_9252,N_2131,N_3265);
nor U9253 (N_9253,N_2805,N_3607);
and U9254 (N_9254,N_4791,N_4644);
and U9255 (N_9255,N_2003,N_3525);
xor U9256 (N_9256,N_1457,N_3787);
xor U9257 (N_9257,N_2560,N_1643);
nand U9258 (N_9258,N_3737,N_4010);
nor U9259 (N_9259,N_3585,N_1116);
and U9260 (N_9260,N_2652,N_798);
xnor U9261 (N_9261,N_2875,N_2016);
nor U9262 (N_9262,N_4285,N_2994);
and U9263 (N_9263,N_3440,N_1432);
or U9264 (N_9264,N_2529,N_1809);
or U9265 (N_9265,N_3134,N_4139);
nor U9266 (N_9266,N_4671,N_1652);
nor U9267 (N_9267,N_3086,N_3197);
nor U9268 (N_9268,N_4101,N_633);
nand U9269 (N_9269,N_3659,N_2184);
nor U9270 (N_9270,N_105,N_824);
or U9271 (N_9271,N_1524,N_1746);
nand U9272 (N_9272,N_4062,N_1996);
and U9273 (N_9273,N_1337,N_189);
nand U9274 (N_9274,N_4937,N_671);
nor U9275 (N_9275,N_4420,N_2907);
and U9276 (N_9276,N_4661,N_2147);
nor U9277 (N_9277,N_941,N_2861);
nand U9278 (N_9278,N_3259,N_980);
nand U9279 (N_9279,N_615,N_1601);
or U9280 (N_9280,N_1481,N_2402);
nor U9281 (N_9281,N_46,N_953);
nor U9282 (N_9282,N_2917,N_3751);
nand U9283 (N_9283,N_2931,N_4486);
and U9284 (N_9284,N_3617,N_4049);
or U9285 (N_9285,N_3415,N_69);
nor U9286 (N_9286,N_778,N_3946);
or U9287 (N_9287,N_2513,N_2301);
or U9288 (N_9288,N_3626,N_3291);
or U9289 (N_9289,N_2225,N_914);
nand U9290 (N_9290,N_3549,N_2809);
nand U9291 (N_9291,N_782,N_4051);
and U9292 (N_9292,N_879,N_2175);
nand U9293 (N_9293,N_3077,N_4771);
or U9294 (N_9294,N_1031,N_534);
nand U9295 (N_9295,N_1176,N_2807);
nor U9296 (N_9296,N_3222,N_4010);
and U9297 (N_9297,N_2678,N_2003);
and U9298 (N_9298,N_1297,N_4722);
xor U9299 (N_9299,N_629,N_2608);
or U9300 (N_9300,N_204,N_3984);
or U9301 (N_9301,N_259,N_3905);
and U9302 (N_9302,N_4071,N_1535);
nand U9303 (N_9303,N_3775,N_896);
xor U9304 (N_9304,N_2004,N_4088);
and U9305 (N_9305,N_1188,N_4902);
and U9306 (N_9306,N_3191,N_1336);
nand U9307 (N_9307,N_290,N_1275);
nor U9308 (N_9308,N_3782,N_1480);
nand U9309 (N_9309,N_3026,N_3931);
and U9310 (N_9310,N_582,N_3747);
nand U9311 (N_9311,N_3278,N_1553);
nand U9312 (N_9312,N_4370,N_2500);
and U9313 (N_9313,N_1338,N_4726);
or U9314 (N_9314,N_4147,N_4428);
nand U9315 (N_9315,N_549,N_262);
nand U9316 (N_9316,N_1716,N_3919);
or U9317 (N_9317,N_2097,N_331);
or U9318 (N_9318,N_4198,N_1633);
and U9319 (N_9319,N_2468,N_3684);
or U9320 (N_9320,N_1032,N_3420);
nor U9321 (N_9321,N_4719,N_4441);
or U9322 (N_9322,N_2618,N_2416);
and U9323 (N_9323,N_3457,N_4420);
nand U9324 (N_9324,N_4023,N_3840);
or U9325 (N_9325,N_1819,N_212);
nand U9326 (N_9326,N_3998,N_2334);
and U9327 (N_9327,N_379,N_4782);
or U9328 (N_9328,N_3037,N_1104);
nand U9329 (N_9329,N_4719,N_1483);
or U9330 (N_9330,N_2130,N_1437);
xnor U9331 (N_9331,N_507,N_2389);
nor U9332 (N_9332,N_2194,N_121);
xnor U9333 (N_9333,N_3380,N_652);
nor U9334 (N_9334,N_2547,N_2927);
xor U9335 (N_9335,N_1911,N_2180);
nand U9336 (N_9336,N_1679,N_4002);
nor U9337 (N_9337,N_895,N_4683);
xnor U9338 (N_9338,N_4588,N_1604);
nor U9339 (N_9339,N_377,N_1301);
nand U9340 (N_9340,N_1729,N_1543);
and U9341 (N_9341,N_198,N_1986);
or U9342 (N_9342,N_406,N_3812);
nand U9343 (N_9343,N_1148,N_1283);
or U9344 (N_9344,N_444,N_275);
nor U9345 (N_9345,N_3288,N_1262);
xnor U9346 (N_9346,N_4300,N_3559);
and U9347 (N_9347,N_86,N_2707);
and U9348 (N_9348,N_665,N_4986);
nand U9349 (N_9349,N_729,N_174);
xor U9350 (N_9350,N_2985,N_4037);
and U9351 (N_9351,N_4463,N_3745);
and U9352 (N_9352,N_741,N_2655);
xor U9353 (N_9353,N_2005,N_3497);
or U9354 (N_9354,N_3669,N_2198);
nand U9355 (N_9355,N_203,N_2427);
xor U9356 (N_9356,N_3084,N_2735);
nor U9357 (N_9357,N_4545,N_4565);
and U9358 (N_9358,N_490,N_810);
nor U9359 (N_9359,N_412,N_136);
or U9360 (N_9360,N_1399,N_549);
and U9361 (N_9361,N_4024,N_2668);
xor U9362 (N_9362,N_3384,N_3165);
nor U9363 (N_9363,N_1081,N_3408);
and U9364 (N_9364,N_1221,N_4196);
and U9365 (N_9365,N_4478,N_3103);
and U9366 (N_9366,N_716,N_4635);
or U9367 (N_9367,N_3464,N_4971);
xor U9368 (N_9368,N_3597,N_3703);
nand U9369 (N_9369,N_4370,N_731);
or U9370 (N_9370,N_4257,N_585);
nand U9371 (N_9371,N_1576,N_1633);
xor U9372 (N_9372,N_3337,N_3662);
nand U9373 (N_9373,N_4204,N_2606);
nand U9374 (N_9374,N_4968,N_3952);
xor U9375 (N_9375,N_2701,N_1441);
nand U9376 (N_9376,N_4456,N_543);
and U9377 (N_9377,N_914,N_4110);
nor U9378 (N_9378,N_3660,N_3821);
nor U9379 (N_9379,N_2501,N_2990);
or U9380 (N_9380,N_3209,N_1491);
or U9381 (N_9381,N_426,N_4833);
nor U9382 (N_9382,N_3593,N_4382);
and U9383 (N_9383,N_1972,N_1207);
xor U9384 (N_9384,N_2967,N_713);
nor U9385 (N_9385,N_89,N_3845);
and U9386 (N_9386,N_4397,N_4863);
xnor U9387 (N_9387,N_2596,N_2220);
nor U9388 (N_9388,N_732,N_4819);
nand U9389 (N_9389,N_3216,N_4646);
xor U9390 (N_9390,N_3241,N_822);
or U9391 (N_9391,N_4634,N_3665);
xor U9392 (N_9392,N_1871,N_2690);
xnor U9393 (N_9393,N_2482,N_2641);
xor U9394 (N_9394,N_4061,N_871);
nand U9395 (N_9395,N_3428,N_3485);
nand U9396 (N_9396,N_4328,N_4590);
xor U9397 (N_9397,N_4809,N_2344);
nand U9398 (N_9398,N_4496,N_159);
nand U9399 (N_9399,N_437,N_4735);
xor U9400 (N_9400,N_3158,N_4232);
or U9401 (N_9401,N_1326,N_1756);
or U9402 (N_9402,N_1049,N_2563);
nand U9403 (N_9403,N_3285,N_1823);
nand U9404 (N_9404,N_2394,N_2466);
and U9405 (N_9405,N_4357,N_4020);
xnor U9406 (N_9406,N_4448,N_567);
and U9407 (N_9407,N_2653,N_2875);
xor U9408 (N_9408,N_3413,N_4245);
or U9409 (N_9409,N_1451,N_3858);
and U9410 (N_9410,N_4591,N_3627);
xnor U9411 (N_9411,N_2294,N_2048);
and U9412 (N_9412,N_1437,N_3503);
nand U9413 (N_9413,N_631,N_1949);
nand U9414 (N_9414,N_202,N_1767);
nand U9415 (N_9415,N_2651,N_4331);
nand U9416 (N_9416,N_1176,N_4580);
xor U9417 (N_9417,N_3062,N_561);
nand U9418 (N_9418,N_4608,N_3462);
nand U9419 (N_9419,N_4133,N_4522);
xor U9420 (N_9420,N_780,N_2451);
and U9421 (N_9421,N_2921,N_3016);
or U9422 (N_9422,N_1052,N_844);
or U9423 (N_9423,N_1330,N_2534);
nor U9424 (N_9424,N_4538,N_373);
or U9425 (N_9425,N_2142,N_2389);
and U9426 (N_9426,N_4751,N_2138);
and U9427 (N_9427,N_1104,N_1059);
or U9428 (N_9428,N_1574,N_2543);
or U9429 (N_9429,N_205,N_2957);
nand U9430 (N_9430,N_2892,N_4170);
and U9431 (N_9431,N_2791,N_2815);
or U9432 (N_9432,N_4958,N_2468);
nor U9433 (N_9433,N_2990,N_787);
or U9434 (N_9434,N_49,N_949);
xnor U9435 (N_9435,N_3078,N_456);
xor U9436 (N_9436,N_2533,N_4526);
xnor U9437 (N_9437,N_3278,N_1270);
or U9438 (N_9438,N_740,N_764);
nand U9439 (N_9439,N_1688,N_2065);
xnor U9440 (N_9440,N_2775,N_3027);
and U9441 (N_9441,N_2846,N_4207);
or U9442 (N_9442,N_1766,N_365);
xor U9443 (N_9443,N_1207,N_2780);
nor U9444 (N_9444,N_290,N_4853);
and U9445 (N_9445,N_2694,N_1145);
or U9446 (N_9446,N_2450,N_1491);
xnor U9447 (N_9447,N_3056,N_4307);
or U9448 (N_9448,N_2453,N_2289);
nand U9449 (N_9449,N_637,N_3217);
or U9450 (N_9450,N_691,N_4389);
xnor U9451 (N_9451,N_1979,N_1616);
or U9452 (N_9452,N_4411,N_1319);
and U9453 (N_9453,N_352,N_4381);
and U9454 (N_9454,N_1659,N_2620);
and U9455 (N_9455,N_4681,N_610);
or U9456 (N_9456,N_341,N_85);
nand U9457 (N_9457,N_86,N_1106);
and U9458 (N_9458,N_2945,N_3803);
nand U9459 (N_9459,N_4056,N_1093);
or U9460 (N_9460,N_3975,N_2863);
and U9461 (N_9461,N_462,N_2557);
xor U9462 (N_9462,N_2141,N_1505);
xnor U9463 (N_9463,N_407,N_2363);
xnor U9464 (N_9464,N_926,N_4706);
nand U9465 (N_9465,N_1722,N_2223);
or U9466 (N_9466,N_104,N_4729);
xor U9467 (N_9467,N_1764,N_4751);
and U9468 (N_9468,N_3846,N_390);
and U9469 (N_9469,N_3202,N_566);
or U9470 (N_9470,N_1470,N_3963);
or U9471 (N_9471,N_4198,N_3854);
or U9472 (N_9472,N_4633,N_2613);
or U9473 (N_9473,N_3278,N_2633);
nand U9474 (N_9474,N_1420,N_849);
xor U9475 (N_9475,N_1231,N_1700);
nand U9476 (N_9476,N_29,N_3505);
and U9477 (N_9477,N_681,N_1729);
nor U9478 (N_9478,N_1203,N_4606);
or U9479 (N_9479,N_2651,N_3262);
nor U9480 (N_9480,N_774,N_3743);
xor U9481 (N_9481,N_3871,N_1371);
and U9482 (N_9482,N_4092,N_4306);
or U9483 (N_9483,N_4753,N_1761);
xor U9484 (N_9484,N_4102,N_1684);
nor U9485 (N_9485,N_4498,N_575);
xnor U9486 (N_9486,N_4047,N_2349);
nand U9487 (N_9487,N_445,N_3655);
nand U9488 (N_9488,N_503,N_1605);
or U9489 (N_9489,N_3983,N_4483);
nand U9490 (N_9490,N_4250,N_4533);
nand U9491 (N_9491,N_2200,N_3726);
and U9492 (N_9492,N_1164,N_1497);
nor U9493 (N_9493,N_3682,N_2103);
nand U9494 (N_9494,N_1417,N_4006);
nand U9495 (N_9495,N_2276,N_3042);
nand U9496 (N_9496,N_409,N_1263);
nand U9497 (N_9497,N_4298,N_136);
or U9498 (N_9498,N_3018,N_1636);
xnor U9499 (N_9499,N_2312,N_2428);
nor U9500 (N_9500,N_2496,N_1689);
and U9501 (N_9501,N_2706,N_809);
xnor U9502 (N_9502,N_1089,N_2397);
nand U9503 (N_9503,N_847,N_3784);
or U9504 (N_9504,N_1284,N_1640);
and U9505 (N_9505,N_1617,N_1306);
and U9506 (N_9506,N_4647,N_796);
xnor U9507 (N_9507,N_1430,N_4485);
or U9508 (N_9508,N_3254,N_2040);
nor U9509 (N_9509,N_3421,N_4322);
or U9510 (N_9510,N_536,N_2752);
nor U9511 (N_9511,N_2436,N_708);
and U9512 (N_9512,N_2389,N_2110);
nand U9513 (N_9513,N_4010,N_3624);
nand U9514 (N_9514,N_345,N_2955);
nor U9515 (N_9515,N_1490,N_4912);
xor U9516 (N_9516,N_93,N_4480);
xnor U9517 (N_9517,N_187,N_3230);
or U9518 (N_9518,N_2189,N_1520);
nand U9519 (N_9519,N_4249,N_473);
xnor U9520 (N_9520,N_920,N_3515);
nand U9521 (N_9521,N_3150,N_3868);
nand U9522 (N_9522,N_885,N_3604);
xnor U9523 (N_9523,N_2729,N_2032);
xor U9524 (N_9524,N_3726,N_1412);
xnor U9525 (N_9525,N_950,N_4403);
or U9526 (N_9526,N_560,N_1041);
or U9527 (N_9527,N_3728,N_1889);
xor U9528 (N_9528,N_2174,N_3588);
nand U9529 (N_9529,N_176,N_1608);
nor U9530 (N_9530,N_536,N_3309);
or U9531 (N_9531,N_1479,N_506);
xor U9532 (N_9532,N_1777,N_3180);
xor U9533 (N_9533,N_150,N_2695);
nand U9534 (N_9534,N_3365,N_3548);
nor U9535 (N_9535,N_2773,N_2277);
nand U9536 (N_9536,N_2405,N_4736);
xor U9537 (N_9537,N_283,N_123);
or U9538 (N_9538,N_2693,N_3314);
and U9539 (N_9539,N_903,N_1031);
nand U9540 (N_9540,N_2719,N_1798);
xnor U9541 (N_9541,N_4853,N_1520);
and U9542 (N_9542,N_1530,N_585);
nand U9543 (N_9543,N_2965,N_1752);
xor U9544 (N_9544,N_3958,N_3873);
xor U9545 (N_9545,N_4779,N_2830);
nor U9546 (N_9546,N_2947,N_3434);
xnor U9547 (N_9547,N_2461,N_3488);
and U9548 (N_9548,N_714,N_3575);
nor U9549 (N_9549,N_1503,N_3261);
nand U9550 (N_9550,N_1889,N_2167);
and U9551 (N_9551,N_260,N_522);
or U9552 (N_9552,N_4915,N_912);
nand U9553 (N_9553,N_2209,N_4626);
nand U9554 (N_9554,N_1614,N_442);
nand U9555 (N_9555,N_529,N_4345);
nand U9556 (N_9556,N_2879,N_2357);
or U9557 (N_9557,N_720,N_1980);
nand U9558 (N_9558,N_3775,N_744);
or U9559 (N_9559,N_1439,N_3344);
or U9560 (N_9560,N_1998,N_1828);
nand U9561 (N_9561,N_1715,N_4006);
and U9562 (N_9562,N_3149,N_4910);
nor U9563 (N_9563,N_3081,N_2434);
or U9564 (N_9564,N_3651,N_3263);
or U9565 (N_9565,N_998,N_3950);
nor U9566 (N_9566,N_3410,N_424);
nor U9567 (N_9567,N_2045,N_190);
and U9568 (N_9568,N_2096,N_408);
nor U9569 (N_9569,N_1547,N_4085);
or U9570 (N_9570,N_1848,N_606);
or U9571 (N_9571,N_4732,N_1716);
and U9572 (N_9572,N_1910,N_4809);
or U9573 (N_9573,N_2959,N_4361);
nor U9574 (N_9574,N_1391,N_311);
xor U9575 (N_9575,N_1756,N_3585);
or U9576 (N_9576,N_4217,N_4824);
nand U9577 (N_9577,N_99,N_1297);
and U9578 (N_9578,N_3711,N_11);
or U9579 (N_9579,N_3050,N_3020);
or U9580 (N_9580,N_1126,N_1531);
or U9581 (N_9581,N_1733,N_2095);
and U9582 (N_9582,N_1686,N_2422);
nand U9583 (N_9583,N_2277,N_1096);
nor U9584 (N_9584,N_3156,N_588);
nand U9585 (N_9585,N_686,N_2539);
and U9586 (N_9586,N_2490,N_1705);
nor U9587 (N_9587,N_2274,N_3652);
xor U9588 (N_9588,N_4762,N_2540);
nor U9589 (N_9589,N_2079,N_579);
nor U9590 (N_9590,N_4042,N_3838);
xnor U9591 (N_9591,N_1807,N_2315);
and U9592 (N_9592,N_4745,N_2901);
or U9593 (N_9593,N_4424,N_3969);
xnor U9594 (N_9594,N_3203,N_3797);
and U9595 (N_9595,N_4298,N_515);
or U9596 (N_9596,N_2510,N_3173);
xnor U9597 (N_9597,N_506,N_3699);
or U9598 (N_9598,N_3427,N_2348);
and U9599 (N_9599,N_2235,N_2887);
nand U9600 (N_9600,N_1507,N_1290);
or U9601 (N_9601,N_3164,N_4649);
and U9602 (N_9602,N_997,N_1291);
nand U9603 (N_9603,N_3264,N_651);
xor U9604 (N_9604,N_1526,N_1599);
xor U9605 (N_9605,N_2115,N_2924);
nand U9606 (N_9606,N_4220,N_3901);
and U9607 (N_9607,N_527,N_253);
and U9608 (N_9608,N_4901,N_4545);
xnor U9609 (N_9609,N_4195,N_833);
xnor U9610 (N_9610,N_3817,N_710);
and U9611 (N_9611,N_2755,N_867);
nor U9612 (N_9612,N_4128,N_1633);
nand U9613 (N_9613,N_4377,N_4554);
or U9614 (N_9614,N_4232,N_4520);
nand U9615 (N_9615,N_3484,N_2240);
nand U9616 (N_9616,N_3971,N_762);
xnor U9617 (N_9617,N_4796,N_3723);
nand U9618 (N_9618,N_2797,N_1297);
nand U9619 (N_9619,N_2447,N_2278);
and U9620 (N_9620,N_4219,N_747);
and U9621 (N_9621,N_3930,N_1904);
xnor U9622 (N_9622,N_3761,N_412);
or U9623 (N_9623,N_4445,N_1227);
nor U9624 (N_9624,N_4429,N_3903);
nor U9625 (N_9625,N_2965,N_3880);
and U9626 (N_9626,N_1855,N_4710);
nor U9627 (N_9627,N_4697,N_2498);
nor U9628 (N_9628,N_1612,N_1314);
or U9629 (N_9629,N_702,N_3712);
and U9630 (N_9630,N_4204,N_2304);
or U9631 (N_9631,N_3088,N_2500);
nor U9632 (N_9632,N_2100,N_4871);
nand U9633 (N_9633,N_3969,N_992);
nor U9634 (N_9634,N_316,N_1388);
nor U9635 (N_9635,N_2156,N_20);
nor U9636 (N_9636,N_2095,N_4032);
or U9637 (N_9637,N_511,N_4660);
xor U9638 (N_9638,N_2112,N_3499);
nand U9639 (N_9639,N_373,N_3723);
xor U9640 (N_9640,N_1109,N_3235);
and U9641 (N_9641,N_128,N_587);
and U9642 (N_9642,N_468,N_3185);
or U9643 (N_9643,N_1040,N_954);
nand U9644 (N_9644,N_2649,N_137);
or U9645 (N_9645,N_1717,N_8);
xor U9646 (N_9646,N_4107,N_3316);
or U9647 (N_9647,N_1516,N_3183);
nor U9648 (N_9648,N_612,N_591);
and U9649 (N_9649,N_3828,N_2452);
or U9650 (N_9650,N_614,N_2953);
nand U9651 (N_9651,N_1864,N_843);
nand U9652 (N_9652,N_3685,N_1019);
nor U9653 (N_9653,N_2859,N_2019);
or U9654 (N_9654,N_4388,N_3411);
xnor U9655 (N_9655,N_3135,N_2881);
and U9656 (N_9656,N_3548,N_841);
and U9657 (N_9657,N_4996,N_63);
xor U9658 (N_9658,N_518,N_2865);
nand U9659 (N_9659,N_1091,N_677);
xor U9660 (N_9660,N_2718,N_4087);
and U9661 (N_9661,N_1074,N_4840);
or U9662 (N_9662,N_423,N_4550);
nor U9663 (N_9663,N_2970,N_2131);
and U9664 (N_9664,N_4136,N_1957);
and U9665 (N_9665,N_1510,N_2773);
and U9666 (N_9666,N_249,N_3575);
nand U9667 (N_9667,N_785,N_3201);
and U9668 (N_9668,N_4493,N_2286);
or U9669 (N_9669,N_1748,N_3403);
nand U9670 (N_9670,N_3098,N_2080);
or U9671 (N_9671,N_2094,N_3880);
nor U9672 (N_9672,N_3367,N_790);
or U9673 (N_9673,N_306,N_592);
and U9674 (N_9674,N_3726,N_2635);
xnor U9675 (N_9675,N_1740,N_134);
nand U9676 (N_9676,N_1432,N_1260);
nand U9677 (N_9677,N_3964,N_2599);
or U9678 (N_9678,N_2785,N_2273);
xor U9679 (N_9679,N_4306,N_1589);
nand U9680 (N_9680,N_947,N_3525);
and U9681 (N_9681,N_3531,N_2088);
and U9682 (N_9682,N_267,N_1183);
nand U9683 (N_9683,N_1132,N_1624);
xnor U9684 (N_9684,N_4456,N_1549);
and U9685 (N_9685,N_2489,N_3231);
nand U9686 (N_9686,N_349,N_1069);
and U9687 (N_9687,N_581,N_4190);
or U9688 (N_9688,N_4929,N_4128);
nor U9689 (N_9689,N_3609,N_1506);
and U9690 (N_9690,N_4631,N_1667);
nor U9691 (N_9691,N_706,N_3373);
nor U9692 (N_9692,N_3401,N_2685);
and U9693 (N_9693,N_4778,N_3304);
and U9694 (N_9694,N_3371,N_1579);
nor U9695 (N_9695,N_4994,N_1863);
nor U9696 (N_9696,N_3949,N_3808);
nor U9697 (N_9697,N_1014,N_4821);
nand U9698 (N_9698,N_2113,N_2577);
nor U9699 (N_9699,N_719,N_3267);
nand U9700 (N_9700,N_4680,N_2605);
xnor U9701 (N_9701,N_3104,N_4933);
nor U9702 (N_9702,N_2284,N_3305);
or U9703 (N_9703,N_3215,N_1365);
or U9704 (N_9704,N_2032,N_182);
or U9705 (N_9705,N_2913,N_12);
xnor U9706 (N_9706,N_4076,N_3202);
nand U9707 (N_9707,N_1041,N_4098);
nor U9708 (N_9708,N_4075,N_4573);
and U9709 (N_9709,N_3250,N_3849);
xor U9710 (N_9710,N_978,N_416);
and U9711 (N_9711,N_3447,N_3841);
nand U9712 (N_9712,N_334,N_1499);
xor U9713 (N_9713,N_1945,N_4858);
nor U9714 (N_9714,N_223,N_968);
and U9715 (N_9715,N_1594,N_894);
and U9716 (N_9716,N_2416,N_3763);
nor U9717 (N_9717,N_2778,N_489);
and U9718 (N_9718,N_4422,N_3638);
nand U9719 (N_9719,N_2910,N_4408);
or U9720 (N_9720,N_3469,N_2550);
or U9721 (N_9721,N_462,N_1605);
nand U9722 (N_9722,N_3660,N_2799);
nand U9723 (N_9723,N_3791,N_4134);
nor U9724 (N_9724,N_2777,N_1242);
and U9725 (N_9725,N_3095,N_2807);
and U9726 (N_9726,N_4274,N_759);
nor U9727 (N_9727,N_1779,N_4922);
or U9728 (N_9728,N_2353,N_4557);
and U9729 (N_9729,N_3948,N_3534);
and U9730 (N_9730,N_374,N_3704);
or U9731 (N_9731,N_2399,N_2796);
or U9732 (N_9732,N_4212,N_4535);
or U9733 (N_9733,N_1226,N_999);
nor U9734 (N_9734,N_3175,N_2436);
nand U9735 (N_9735,N_960,N_290);
nand U9736 (N_9736,N_4555,N_7);
xor U9737 (N_9737,N_2378,N_981);
and U9738 (N_9738,N_657,N_1742);
xor U9739 (N_9739,N_2027,N_194);
or U9740 (N_9740,N_285,N_4244);
or U9741 (N_9741,N_3563,N_2690);
xnor U9742 (N_9742,N_1353,N_2201);
nand U9743 (N_9743,N_4960,N_3466);
or U9744 (N_9744,N_509,N_732);
and U9745 (N_9745,N_3333,N_360);
nand U9746 (N_9746,N_2099,N_3322);
and U9747 (N_9747,N_3849,N_3876);
xor U9748 (N_9748,N_3620,N_3774);
xor U9749 (N_9749,N_953,N_2425);
nor U9750 (N_9750,N_3131,N_4798);
nand U9751 (N_9751,N_3879,N_2042);
or U9752 (N_9752,N_1827,N_124);
or U9753 (N_9753,N_2483,N_2358);
or U9754 (N_9754,N_3654,N_925);
nand U9755 (N_9755,N_1479,N_4571);
or U9756 (N_9756,N_1832,N_1456);
and U9757 (N_9757,N_3632,N_1849);
and U9758 (N_9758,N_1239,N_4638);
or U9759 (N_9759,N_1257,N_1417);
and U9760 (N_9760,N_3375,N_322);
and U9761 (N_9761,N_1530,N_2448);
and U9762 (N_9762,N_3486,N_3229);
xnor U9763 (N_9763,N_3220,N_2545);
nor U9764 (N_9764,N_4851,N_2317);
and U9765 (N_9765,N_1759,N_3231);
nand U9766 (N_9766,N_3288,N_552);
and U9767 (N_9767,N_2508,N_4887);
nor U9768 (N_9768,N_491,N_1953);
or U9769 (N_9769,N_3977,N_2318);
and U9770 (N_9770,N_1699,N_655);
xnor U9771 (N_9771,N_524,N_659);
nand U9772 (N_9772,N_4573,N_3740);
and U9773 (N_9773,N_1438,N_3642);
xor U9774 (N_9774,N_388,N_2949);
nor U9775 (N_9775,N_2436,N_4475);
or U9776 (N_9776,N_924,N_2598);
nand U9777 (N_9777,N_3366,N_882);
nor U9778 (N_9778,N_1621,N_831);
or U9779 (N_9779,N_270,N_2016);
or U9780 (N_9780,N_4278,N_1442);
nor U9781 (N_9781,N_1527,N_3790);
xor U9782 (N_9782,N_1588,N_4565);
and U9783 (N_9783,N_722,N_824);
xor U9784 (N_9784,N_1682,N_1039);
nand U9785 (N_9785,N_3786,N_1611);
nand U9786 (N_9786,N_1211,N_4108);
xnor U9787 (N_9787,N_1554,N_2071);
or U9788 (N_9788,N_4,N_4947);
or U9789 (N_9789,N_659,N_3291);
xnor U9790 (N_9790,N_3344,N_4551);
or U9791 (N_9791,N_2696,N_3168);
xor U9792 (N_9792,N_1411,N_3589);
xor U9793 (N_9793,N_1232,N_1415);
xor U9794 (N_9794,N_3582,N_1337);
nor U9795 (N_9795,N_2386,N_669);
nor U9796 (N_9796,N_868,N_2552);
or U9797 (N_9797,N_2338,N_2792);
xor U9798 (N_9798,N_906,N_2423);
xnor U9799 (N_9799,N_160,N_1702);
nor U9800 (N_9800,N_4448,N_1978);
and U9801 (N_9801,N_2466,N_2271);
and U9802 (N_9802,N_3633,N_3991);
and U9803 (N_9803,N_2190,N_3278);
nor U9804 (N_9804,N_1971,N_4433);
and U9805 (N_9805,N_2892,N_1831);
and U9806 (N_9806,N_4369,N_4513);
nor U9807 (N_9807,N_2535,N_2475);
nor U9808 (N_9808,N_1186,N_960);
or U9809 (N_9809,N_2201,N_3270);
or U9810 (N_9810,N_4457,N_4340);
and U9811 (N_9811,N_4614,N_1824);
nor U9812 (N_9812,N_30,N_2553);
xor U9813 (N_9813,N_1383,N_817);
xnor U9814 (N_9814,N_4567,N_2587);
nor U9815 (N_9815,N_1542,N_2228);
or U9816 (N_9816,N_3463,N_366);
and U9817 (N_9817,N_2922,N_215);
xnor U9818 (N_9818,N_4448,N_859);
xor U9819 (N_9819,N_1921,N_344);
xnor U9820 (N_9820,N_3259,N_2446);
xor U9821 (N_9821,N_2272,N_119);
and U9822 (N_9822,N_1729,N_2778);
nand U9823 (N_9823,N_4684,N_907);
and U9824 (N_9824,N_77,N_3567);
nand U9825 (N_9825,N_2649,N_4772);
nand U9826 (N_9826,N_4515,N_1564);
nand U9827 (N_9827,N_3753,N_1984);
and U9828 (N_9828,N_1540,N_3797);
nor U9829 (N_9829,N_3733,N_1557);
or U9830 (N_9830,N_2949,N_522);
or U9831 (N_9831,N_4906,N_2427);
xnor U9832 (N_9832,N_3966,N_1346);
xnor U9833 (N_9833,N_2875,N_336);
or U9834 (N_9834,N_245,N_2230);
and U9835 (N_9835,N_2747,N_2188);
and U9836 (N_9836,N_55,N_3345);
and U9837 (N_9837,N_1789,N_4937);
nor U9838 (N_9838,N_2935,N_3512);
nand U9839 (N_9839,N_2348,N_2998);
nand U9840 (N_9840,N_319,N_1336);
or U9841 (N_9841,N_1971,N_3263);
xnor U9842 (N_9842,N_1281,N_4215);
and U9843 (N_9843,N_2056,N_2526);
or U9844 (N_9844,N_4752,N_954);
nor U9845 (N_9845,N_1987,N_2026);
xnor U9846 (N_9846,N_4408,N_25);
nor U9847 (N_9847,N_1599,N_1968);
nor U9848 (N_9848,N_4696,N_2419);
nand U9849 (N_9849,N_4323,N_4625);
nand U9850 (N_9850,N_4038,N_2358);
or U9851 (N_9851,N_3479,N_3607);
or U9852 (N_9852,N_4636,N_3831);
or U9853 (N_9853,N_96,N_1091);
nand U9854 (N_9854,N_1340,N_3313);
xnor U9855 (N_9855,N_1563,N_1854);
and U9856 (N_9856,N_2058,N_1639);
or U9857 (N_9857,N_4651,N_3786);
and U9858 (N_9858,N_3629,N_4999);
or U9859 (N_9859,N_190,N_3885);
or U9860 (N_9860,N_353,N_2388);
and U9861 (N_9861,N_4076,N_4663);
xnor U9862 (N_9862,N_3921,N_4594);
nor U9863 (N_9863,N_382,N_4052);
nor U9864 (N_9864,N_3131,N_591);
and U9865 (N_9865,N_1008,N_2197);
xor U9866 (N_9866,N_2799,N_4990);
nand U9867 (N_9867,N_919,N_4529);
or U9868 (N_9868,N_3028,N_4861);
xnor U9869 (N_9869,N_1425,N_4522);
nand U9870 (N_9870,N_3518,N_4352);
nor U9871 (N_9871,N_184,N_4541);
and U9872 (N_9872,N_3154,N_4399);
nand U9873 (N_9873,N_4010,N_2614);
or U9874 (N_9874,N_2994,N_4630);
xnor U9875 (N_9875,N_2948,N_933);
nor U9876 (N_9876,N_4030,N_3585);
and U9877 (N_9877,N_1998,N_1660);
xor U9878 (N_9878,N_1926,N_1416);
or U9879 (N_9879,N_3410,N_1341);
or U9880 (N_9880,N_2181,N_214);
or U9881 (N_9881,N_2265,N_643);
nor U9882 (N_9882,N_2874,N_2818);
nor U9883 (N_9883,N_3605,N_3436);
xor U9884 (N_9884,N_3350,N_4489);
nand U9885 (N_9885,N_4455,N_1063);
or U9886 (N_9886,N_931,N_4437);
nor U9887 (N_9887,N_2095,N_2569);
and U9888 (N_9888,N_4255,N_4453);
and U9889 (N_9889,N_4830,N_2199);
nor U9890 (N_9890,N_998,N_4581);
or U9891 (N_9891,N_1462,N_1686);
nor U9892 (N_9892,N_3275,N_15);
nand U9893 (N_9893,N_1355,N_45);
xnor U9894 (N_9894,N_4109,N_4799);
or U9895 (N_9895,N_2768,N_2634);
xnor U9896 (N_9896,N_3764,N_4576);
nor U9897 (N_9897,N_4756,N_3063);
nand U9898 (N_9898,N_3596,N_789);
nor U9899 (N_9899,N_3592,N_3199);
or U9900 (N_9900,N_903,N_549);
xor U9901 (N_9901,N_3992,N_276);
xor U9902 (N_9902,N_1324,N_2428);
and U9903 (N_9903,N_4630,N_3745);
or U9904 (N_9904,N_3761,N_1479);
nor U9905 (N_9905,N_2255,N_3336);
xor U9906 (N_9906,N_1931,N_4965);
or U9907 (N_9907,N_2249,N_2861);
or U9908 (N_9908,N_1532,N_740);
xnor U9909 (N_9909,N_4983,N_433);
xnor U9910 (N_9910,N_430,N_1003);
xnor U9911 (N_9911,N_1879,N_1615);
xor U9912 (N_9912,N_1500,N_2107);
xor U9913 (N_9913,N_3442,N_2201);
and U9914 (N_9914,N_2717,N_3077);
or U9915 (N_9915,N_3896,N_1809);
and U9916 (N_9916,N_2397,N_4673);
xor U9917 (N_9917,N_4412,N_4703);
or U9918 (N_9918,N_1257,N_395);
xor U9919 (N_9919,N_2309,N_3662);
or U9920 (N_9920,N_2842,N_3820);
xor U9921 (N_9921,N_2409,N_664);
xnor U9922 (N_9922,N_564,N_3754);
xor U9923 (N_9923,N_646,N_4532);
nor U9924 (N_9924,N_3619,N_3914);
nand U9925 (N_9925,N_2210,N_1088);
nand U9926 (N_9926,N_3310,N_919);
nor U9927 (N_9927,N_545,N_4766);
xnor U9928 (N_9928,N_4170,N_2969);
nand U9929 (N_9929,N_2829,N_539);
or U9930 (N_9930,N_4507,N_623);
nand U9931 (N_9931,N_1774,N_1423);
nor U9932 (N_9932,N_1458,N_2697);
nor U9933 (N_9933,N_4312,N_659);
or U9934 (N_9934,N_491,N_3739);
xnor U9935 (N_9935,N_2818,N_3434);
nor U9936 (N_9936,N_2526,N_4882);
and U9937 (N_9937,N_2944,N_3028);
or U9938 (N_9938,N_305,N_4105);
xor U9939 (N_9939,N_1380,N_3512);
nand U9940 (N_9940,N_3996,N_2619);
xor U9941 (N_9941,N_572,N_2182);
and U9942 (N_9942,N_1506,N_2495);
nor U9943 (N_9943,N_724,N_1528);
nand U9944 (N_9944,N_2157,N_799);
nand U9945 (N_9945,N_772,N_2353);
nand U9946 (N_9946,N_3458,N_3932);
and U9947 (N_9947,N_4910,N_3953);
or U9948 (N_9948,N_1160,N_1479);
or U9949 (N_9949,N_4475,N_3046);
or U9950 (N_9950,N_4001,N_3174);
xor U9951 (N_9951,N_4118,N_3411);
or U9952 (N_9952,N_4232,N_536);
and U9953 (N_9953,N_2289,N_2003);
nor U9954 (N_9954,N_136,N_4342);
nand U9955 (N_9955,N_1573,N_3586);
nand U9956 (N_9956,N_1721,N_4602);
xor U9957 (N_9957,N_4098,N_4091);
and U9958 (N_9958,N_2803,N_3219);
and U9959 (N_9959,N_2144,N_1877);
and U9960 (N_9960,N_1825,N_1081);
nand U9961 (N_9961,N_2279,N_1106);
or U9962 (N_9962,N_4818,N_3899);
xor U9963 (N_9963,N_2710,N_2226);
nor U9964 (N_9964,N_2635,N_4671);
xor U9965 (N_9965,N_3233,N_889);
or U9966 (N_9966,N_3375,N_1961);
or U9967 (N_9967,N_4790,N_1212);
nand U9968 (N_9968,N_892,N_594);
or U9969 (N_9969,N_2393,N_1696);
nand U9970 (N_9970,N_1979,N_4758);
or U9971 (N_9971,N_2432,N_4633);
or U9972 (N_9972,N_3009,N_3738);
xor U9973 (N_9973,N_4190,N_2628);
nand U9974 (N_9974,N_1638,N_94);
nand U9975 (N_9975,N_2815,N_2351);
and U9976 (N_9976,N_2946,N_95);
and U9977 (N_9977,N_4798,N_4206);
or U9978 (N_9978,N_4477,N_3898);
nor U9979 (N_9979,N_1121,N_3861);
nor U9980 (N_9980,N_1481,N_1944);
and U9981 (N_9981,N_4060,N_1751);
nor U9982 (N_9982,N_4540,N_4681);
xor U9983 (N_9983,N_3510,N_4397);
and U9984 (N_9984,N_3581,N_717);
nand U9985 (N_9985,N_3704,N_3077);
xor U9986 (N_9986,N_4175,N_2045);
nor U9987 (N_9987,N_3759,N_2155);
xor U9988 (N_9988,N_2123,N_2929);
and U9989 (N_9989,N_2729,N_793);
or U9990 (N_9990,N_1692,N_2683);
nand U9991 (N_9991,N_3,N_988);
xnor U9992 (N_9992,N_3218,N_105);
nand U9993 (N_9993,N_498,N_2874);
and U9994 (N_9994,N_53,N_914);
nor U9995 (N_9995,N_1994,N_1918);
and U9996 (N_9996,N_629,N_4964);
xor U9997 (N_9997,N_1759,N_936);
nand U9998 (N_9998,N_877,N_4640);
and U9999 (N_9999,N_2784,N_4955);
nand U10000 (N_10000,N_5539,N_6638);
nor U10001 (N_10001,N_7201,N_9168);
and U10002 (N_10002,N_5963,N_5485);
and U10003 (N_10003,N_6853,N_5528);
and U10004 (N_10004,N_6558,N_9154);
xnor U10005 (N_10005,N_9803,N_9821);
nand U10006 (N_10006,N_9028,N_6186);
nor U10007 (N_10007,N_8917,N_8997);
nor U10008 (N_10008,N_6532,N_5697);
nor U10009 (N_10009,N_5933,N_6528);
or U10010 (N_10010,N_9605,N_9954);
nor U10011 (N_10011,N_7145,N_8724);
or U10012 (N_10012,N_8849,N_6876);
nor U10013 (N_10013,N_7687,N_7511);
nor U10014 (N_10014,N_9575,N_7611);
nand U10015 (N_10015,N_8144,N_9628);
nor U10016 (N_10016,N_8830,N_7872);
or U10017 (N_10017,N_5052,N_5257);
or U10018 (N_10018,N_5405,N_5364);
nand U10019 (N_10019,N_9325,N_5049);
xnor U10020 (N_10020,N_7799,N_8592);
nand U10021 (N_10021,N_7616,N_9226);
or U10022 (N_10022,N_6652,N_6172);
nor U10023 (N_10023,N_7630,N_8384);
and U10024 (N_10024,N_9093,N_8395);
or U10025 (N_10025,N_6438,N_9912);
nor U10026 (N_10026,N_6810,N_9430);
xor U10027 (N_10027,N_7798,N_6405);
xnor U10028 (N_10028,N_5242,N_8879);
xnor U10029 (N_10029,N_8749,N_8921);
nand U10030 (N_10030,N_5321,N_5526);
xor U10031 (N_10031,N_8211,N_6150);
nand U10032 (N_10032,N_9561,N_8140);
and U10033 (N_10033,N_5846,N_7628);
nand U10034 (N_10034,N_5320,N_6848);
nand U10035 (N_10035,N_5538,N_6597);
and U10036 (N_10036,N_8782,N_7476);
and U10037 (N_10037,N_6279,N_5802);
or U10038 (N_10038,N_5647,N_9651);
xnor U10039 (N_10039,N_6934,N_5984);
xor U10040 (N_10040,N_9685,N_5236);
nor U10041 (N_10041,N_5724,N_6308);
or U10042 (N_10042,N_7512,N_8359);
and U10043 (N_10043,N_6696,N_5830);
nand U10044 (N_10044,N_6072,N_7463);
nor U10045 (N_10045,N_9566,N_8662);
nor U10046 (N_10046,N_5200,N_6453);
and U10047 (N_10047,N_9948,N_5627);
nand U10048 (N_10048,N_6512,N_6859);
xor U10049 (N_10049,N_9852,N_7956);
nor U10050 (N_10050,N_7744,N_6775);
or U10051 (N_10051,N_5029,N_5165);
xnor U10052 (N_10052,N_9621,N_9815);
or U10053 (N_10053,N_5918,N_6651);
or U10054 (N_10054,N_8496,N_6871);
and U10055 (N_10055,N_6141,N_8486);
nor U10056 (N_10056,N_7438,N_8363);
or U10057 (N_10057,N_6268,N_9393);
and U10058 (N_10058,N_9564,N_8223);
xor U10059 (N_10059,N_5305,N_5121);
nand U10060 (N_10060,N_9778,N_9938);
or U10061 (N_10061,N_8641,N_7778);
or U10062 (N_10062,N_9887,N_6857);
nand U10063 (N_10063,N_7711,N_5151);
xnor U10064 (N_10064,N_5383,N_9704);
and U10065 (N_10065,N_7980,N_6081);
nor U10066 (N_10066,N_7229,N_7312);
or U10067 (N_10067,N_8827,N_8970);
or U10068 (N_10068,N_9634,N_7268);
nor U10069 (N_10069,N_6395,N_8817);
and U10070 (N_10070,N_6443,N_6855);
nor U10071 (N_10071,N_8050,N_9919);
xor U10072 (N_10072,N_5138,N_5637);
nand U10073 (N_10073,N_5490,N_9654);
and U10074 (N_10074,N_7447,N_5112);
or U10075 (N_10075,N_5212,N_7501);
nand U10076 (N_10076,N_5074,N_8784);
or U10077 (N_10077,N_6388,N_5433);
nor U10078 (N_10078,N_9280,N_7454);
and U10079 (N_10079,N_5949,N_9565);
nand U10080 (N_10080,N_8658,N_6232);
xor U10081 (N_10081,N_5421,N_9313);
or U10082 (N_10082,N_6290,N_5615);
nor U10083 (N_10083,N_7164,N_6970);
nand U10084 (N_10084,N_5294,N_6974);
or U10085 (N_10085,N_8113,N_9265);
or U10086 (N_10086,N_7964,N_6258);
or U10087 (N_10087,N_5658,N_5593);
and U10088 (N_10088,N_6989,N_9023);
nor U10089 (N_10089,N_9013,N_8736);
or U10090 (N_10090,N_5071,N_5501);
xor U10091 (N_10091,N_7242,N_7063);
and U10092 (N_10092,N_6152,N_6682);
xor U10093 (N_10093,N_8112,N_5811);
nor U10094 (N_10094,N_5887,N_5907);
xnor U10095 (N_10095,N_7364,N_8543);
nor U10096 (N_10096,N_5763,N_7523);
nor U10097 (N_10097,N_9335,N_9553);
or U10098 (N_10098,N_9688,N_6215);
and U10099 (N_10099,N_7252,N_7198);
or U10100 (N_10100,N_6497,N_7383);
xnor U10101 (N_10101,N_6101,N_5894);
xnor U10102 (N_10102,N_5347,N_7689);
xor U10103 (N_10103,N_9472,N_7489);
nand U10104 (N_10104,N_5643,N_5234);
xnor U10105 (N_10105,N_5829,N_8005);
or U10106 (N_10106,N_8468,N_5155);
and U10107 (N_10107,N_6997,N_5446);
xor U10108 (N_10108,N_7434,N_5101);
or U10109 (N_10109,N_8504,N_9059);
and U10110 (N_10110,N_6433,N_7772);
nor U10111 (N_10111,N_5263,N_5036);
nor U10112 (N_10112,N_6389,N_8924);
xor U10113 (N_10113,N_9513,N_8520);
nor U10114 (N_10114,N_6650,N_6729);
and U10115 (N_10115,N_9806,N_7070);
or U10116 (N_10116,N_8435,N_9407);
or U10117 (N_10117,N_6017,N_7975);
and U10118 (N_10118,N_8816,N_8730);
nor U10119 (N_10119,N_9632,N_7251);
and U10120 (N_10120,N_7688,N_7718);
xor U10121 (N_10121,N_5319,N_6129);
or U10122 (N_10122,N_6767,N_9310);
nand U10123 (N_10123,N_8769,N_8820);
nand U10124 (N_10124,N_5472,N_7542);
xor U10125 (N_10125,N_6280,N_5605);
nand U10126 (N_10126,N_8625,N_5955);
nand U10127 (N_10127,N_9087,N_9579);
and U10128 (N_10128,N_5299,N_9252);
nor U10129 (N_10129,N_6070,N_6107);
nor U10130 (N_10130,N_8860,N_6121);
or U10131 (N_10131,N_9996,N_6694);
xnor U10132 (N_10132,N_5799,N_7901);
xor U10133 (N_10133,N_8835,N_6078);
xor U10134 (N_10134,N_7836,N_6439);
nor U10135 (N_10135,N_9989,N_6282);
or U10136 (N_10136,N_6408,N_7045);
or U10137 (N_10137,N_6190,N_8758);
or U10138 (N_10138,N_8811,N_6688);
nor U10139 (N_10139,N_6628,N_7931);
or U10140 (N_10140,N_7617,N_5468);
xnor U10141 (N_10141,N_7203,N_6448);
nand U10142 (N_10142,N_7482,N_5042);
nand U10143 (N_10143,N_5199,N_9135);
nand U10144 (N_10144,N_6985,N_8834);
nor U10145 (N_10145,N_7776,N_6194);
xor U10146 (N_10146,N_6449,N_7710);
or U10147 (N_10147,N_6541,N_9677);
nand U10148 (N_10148,N_8068,N_5149);
nand U10149 (N_10149,N_9365,N_6836);
or U10150 (N_10150,N_5358,N_5389);
xor U10151 (N_10151,N_9164,N_8652);
or U10152 (N_10152,N_8532,N_5237);
nand U10153 (N_10153,N_7792,N_5513);
and U10154 (N_10154,N_7825,N_5926);
and U10155 (N_10155,N_6745,N_8360);
xnor U10156 (N_10156,N_8407,N_6206);
or U10157 (N_10157,N_7178,N_7235);
or U10158 (N_10158,N_6302,N_7297);
xor U10159 (N_10159,N_8019,N_8974);
nand U10160 (N_10160,N_9589,N_7466);
or U10161 (N_10161,N_7076,N_9437);
xor U10162 (N_10162,N_6478,N_8557);
xor U10163 (N_10163,N_5194,N_5486);
nor U10164 (N_10164,N_9511,N_8577);
xor U10165 (N_10165,N_6851,N_7957);
nand U10166 (N_10166,N_5790,N_6227);
or U10167 (N_10167,N_8150,N_8097);
nor U10168 (N_10168,N_5185,N_9452);
nand U10169 (N_10169,N_5938,N_8372);
xor U10170 (N_10170,N_6106,N_7195);
nand U10171 (N_10171,N_9411,N_5686);
xor U10172 (N_10172,N_9999,N_5027);
and U10173 (N_10173,N_8147,N_8611);
nor U10174 (N_10174,N_7245,N_9991);
nor U10175 (N_10175,N_7499,N_9895);
nand U10176 (N_10176,N_7994,N_8159);
xor U10177 (N_10177,N_7459,N_5759);
nand U10178 (N_10178,N_7111,N_9030);
and U10179 (N_10179,N_7638,N_7594);
and U10180 (N_10180,N_6151,N_8871);
or U10181 (N_10181,N_6033,N_6169);
nor U10182 (N_10182,N_8710,N_7884);
xor U10183 (N_10183,N_5009,N_5323);
xnor U10184 (N_10184,N_6752,N_6642);
nand U10185 (N_10185,N_6707,N_8690);
or U10186 (N_10186,N_6444,N_5307);
or U10187 (N_10187,N_6915,N_9540);
or U10188 (N_10188,N_7845,N_5552);
and U10189 (N_10189,N_6637,N_8403);
and U10190 (N_10190,N_9233,N_8181);
nor U10191 (N_10191,N_7952,N_7899);
or U10192 (N_10192,N_5688,N_5306);
and U10193 (N_10193,N_7046,N_5571);
and U10194 (N_10194,N_9378,N_5904);
nor U10195 (N_10195,N_9470,N_9921);
nor U10196 (N_10196,N_7951,N_5505);
and U10197 (N_10197,N_9101,N_8206);
xnor U10198 (N_10198,N_7030,N_9084);
or U10199 (N_10199,N_8594,N_7143);
xor U10200 (N_10200,N_9717,N_9570);
nand U10201 (N_10201,N_9219,N_7129);
nand U10202 (N_10202,N_5303,N_6063);
nor U10203 (N_10203,N_7025,N_9067);
and U10204 (N_10204,N_5426,N_6056);
nor U10205 (N_10205,N_8900,N_8312);
and U10206 (N_10206,N_6464,N_8729);
xnor U10207 (N_10207,N_8261,N_7519);
nand U10208 (N_10208,N_5633,N_6509);
and U10209 (N_10209,N_7414,N_5120);
or U10210 (N_10210,N_7486,N_6479);
and U10211 (N_10211,N_8476,N_6248);
or U10212 (N_10212,N_6678,N_9548);
nand U10213 (N_10213,N_7552,N_9758);
xor U10214 (N_10214,N_6401,N_7780);
nor U10215 (N_10215,N_5300,N_6483);
nor U10216 (N_10216,N_5317,N_6817);
nor U10217 (N_10217,N_9952,N_5709);
or U10218 (N_10218,N_7054,N_7323);
or U10219 (N_10219,N_8684,N_8963);
or U10220 (N_10220,N_6935,N_6153);
and U10221 (N_10221,N_9997,N_9930);
or U10222 (N_10222,N_8057,N_9406);
nor U10223 (N_10223,N_7914,N_9495);
nor U10224 (N_10224,N_7878,N_9746);
nand U10225 (N_10225,N_5664,N_9681);
or U10226 (N_10226,N_7289,N_9200);
nand U10227 (N_10227,N_5708,N_7576);
nand U10228 (N_10228,N_5924,N_9480);
xor U10229 (N_10229,N_5466,N_7044);
nor U10230 (N_10230,N_9780,N_5506);
and U10231 (N_10231,N_9834,N_9196);
and U10232 (N_10232,N_6199,N_5013);
and U10233 (N_10233,N_7284,N_9061);
xor U10234 (N_10234,N_5570,N_7859);
nand U10235 (N_10235,N_9960,N_6491);
or U10236 (N_10236,N_9530,N_6096);
and U10237 (N_10237,N_8017,N_5797);
xor U10238 (N_10238,N_8512,N_8876);
nand U10239 (N_10239,N_7181,N_6109);
nor U10240 (N_10240,N_8034,N_7303);
and U10241 (N_10241,N_6122,N_7574);
nor U10242 (N_10242,N_6815,N_9745);
xor U10243 (N_10243,N_8009,N_9959);
and U10244 (N_10244,N_6288,N_5026);
or U10245 (N_10245,N_7422,N_7308);
xor U10246 (N_10246,N_5959,N_5469);
and U10247 (N_10247,N_6045,N_5249);
and U10248 (N_10248,N_7255,N_7266);
xor U10249 (N_10249,N_6559,N_8825);
or U10250 (N_10250,N_8258,N_7742);
xor U10251 (N_10251,N_6736,N_9272);
xnor U10252 (N_10252,N_5621,N_7029);
and U10253 (N_10253,N_5183,N_5967);
or U10254 (N_10254,N_5649,N_9064);
nand U10255 (N_10255,N_6837,N_6536);
xor U10256 (N_10256,N_9870,N_9418);
or U10257 (N_10257,N_8174,N_9016);
and U10258 (N_10258,N_8288,N_9772);
and U10259 (N_10259,N_9877,N_8627);
or U10260 (N_10260,N_7442,N_6455);
or U10261 (N_10261,N_9390,N_5872);
xnor U10262 (N_10262,N_9885,N_7564);
xnor U10263 (N_10263,N_9062,N_6486);
nor U10264 (N_10264,N_9615,N_6346);
and U10265 (N_10265,N_8638,N_6720);
nor U10266 (N_10266,N_6051,N_5073);
xor U10267 (N_10267,N_7568,N_9420);
and U10268 (N_10268,N_9805,N_5198);
xor U10269 (N_10269,N_7468,N_7259);
xor U10270 (N_10270,N_5162,N_9661);
nand U10271 (N_10271,N_8184,N_6420);
nand U10272 (N_10272,N_8481,N_8912);
or U10273 (N_10273,N_5292,N_6012);
and U10274 (N_10274,N_9309,N_5197);
xor U10275 (N_10275,N_8252,N_6368);
and U10276 (N_10276,N_9337,N_7374);
xnor U10277 (N_10277,N_8374,N_6432);
nand U10278 (N_10278,N_7522,N_6948);
and U10279 (N_10279,N_6235,N_9032);
nor U10280 (N_10280,N_6270,N_7356);
xor U10281 (N_10281,N_8482,N_6896);
nand U10282 (N_10282,N_8254,N_7079);
nor U10283 (N_10283,N_5577,N_8420);
nand U10284 (N_10284,N_5262,N_5998);
and U10285 (N_10285,N_9800,N_8348);
xor U10286 (N_10286,N_6730,N_5330);
nand U10287 (N_10287,N_9118,N_6703);
or U10288 (N_10288,N_7987,N_9881);
xor U10289 (N_10289,N_5931,N_7332);
nand U10290 (N_10290,N_8693,N_9240);
xor U10291 (N_10291,N_8785,N_5956);
or U10292 (N_10292,N_6862,N_9024);
nand U10293 (N_10293,N_6972,N_7413);
nor U10294 (N_10294,N_7902,N_9002);
or U10295 (N_10295,N_9205,N_9665);
nor U10296 (N_10296,N_9146,N_8882);
and U10297 (N_10297,N_9449,N_8895);
nor U10298 (N_10298,N_6252,N_9929);
nand U10299 (N_10299,N_8561,N_6306);
or U10300 (N_10300,N_9576,N_8660);
and U10301 (N_10301,N_5588,N_9379);
and U10302 (N_10302,N_5333,N_5619);
xnor U10303 (N_10303,N_9730,N_8665);
and U10304 (N_10304,N_7701,N_9319);
xnor U10305 (N_10305,N_6276,N_7661);
xnor U10306 (N_10306,N_7812,N_9010);
nor U10307 (N_10307,N_6905,N_9491);
and U10308 (N_10308,N_8193,N_7763);
nor U10309 (N_10309,N_7717,N_6445);
nand U10310 (N_10310,N_8191,N_8927);
or U10311 (N_10311,N_5224,N_6293);
nand U10312 (N_10312,N_7550,N_5130);
and U10313 (N_10313,N_8283,N_8326);
or U10314 (N_10314,N_6787,N_9211);
nand U10315 (N_10315,N_7598,N_7092);
and U10316 (N_10316,N_9713,N_8722);
and U10317 (N_10317,N_6971,N_6452);
and U10318 (N_10318,N_7094,N_8219);
and U10319 (N_10319,N_9645,N_8337);
nand U10320 (N_10320,N_7065,N_7493);
xor U10321 (N_10321,N_9558,N_9445);
or U10322 (N_10322,N_8383,N_8197);
or U10323 (N_10323,N_7134,N_9964);
xor U10324 (N_10324,N_6038,N_9250);
or U10325 (N_10325,N_6034,N_6892);
or U10326 (N_10326,N_8687,N_5676);
nor U10327 (N_10327,N_9435,N_7754);
nor U10328 (N_10328,N_5328,N_9297);
and U10329 (N_10329,N_9180,N_8657);
or U10330 (N_10330,N_7648,N_8302);
or U10331 (N_10331,N_6487,N_8189);
nand U10332 (N_10332,N_9988,N_6554);
nor U10333 (N_10333,N_8382,N_6534);
xor U10334 (N_10334,N_5774,N_7163);
or U10335 (N_10335,N_8418,N_9759);
nor U10336 (N_10336,N_9535,N_5308);
nor U10337 (N_10337,N_5082,N_6672);
and U10338 (N_10338,N_9199,N_8727);
or U10339 (N_10339,N_8506,N_6986);
nand U10340 (N_10340,N_9550,N_8479);
xor U10341 (N_10341,N_6612,N_9409);
nand U10342 (N_10342,N_8414,N_5772);
or U10343 (N_10343,N_7965,N_9096);
or U10344 (N_10344,N_9722,N_5831);
nor U10345 (N_10345,N_8537,N_6867);
nand U10346 (N_10346,N_8572,N_5509);
nor U10347 (N_10347,N_9275,N_8129);
or U10348 (N_10348,N_7927,N_5527);
xnor U10349 (N_10349,N_9892,N_6230);
nand U10350 (N_10350,N_7894,N_5815);
nor U10351 (N_10351,N_6006,N_9732);
nand U10352 (N_10352,N_5804,N_5144);
nor U10353 (N_10353,N_5873,N_8308);
xnor U10354 (N_10354,N_8031,N_7887);
nand U10355 (N_10355,N_5034,N_9539);
nand U10356 (N_10356,N_8851,N_8704);
xnor U10357 (N_10357,N_7386,N_9245);
nor U10358 (N_10358,N_9691,N_6819);
xnor U10359 (N_10359,N_8616,N_7378);
xor U10360 (N_10360,N_8004,N_9242);
nand U10361 (N_10361,N_8919,N_6947);
nand U10362 (N_10362,N_6372,N_8433);
nand U10363 (N_10363,N_8554,N_5534);
xor U10364 (N_10364,N_5845,N_5271);
and U10365 (N_10365,N_5483,N_6358);
nand U10366 (N_10366,N_6383,N_9126);
and U10367 (N_10367,N_9288,N_9674);
nor U10368 (N_10368,N_7254,N_5739);
and U10369 (N_10369,N_9440,N_7880);
or U10370 (N_10370,N_6626,N_9973);
or U10371 (N_10371,N_8668,N_7566);
xnor U10372 (N_10372,N_9157,N_9474);
or U10373 (N_10373,N_9484,N_9367);
and U10374 (N_10374,N_9022,N_7755);
nand U10375 (N_10375,N_6609,N_8455);
or U10376 (N_10376,N_9637,N_9939);
xor U10377 (N_10377,N_9764,N_9998);
xnor U10378 (N_10378,N_6116,N_5522);
nand U10379 (N_10379,N_5078,N_7806);
nor U10380 (N_10380,N_8651,N_5640);
or U10381 (N_10381,N_7504,N_7043);
nand U10382 (N_10382,N_6976,N_5394);
nand U10383 (N_10383,N_5022,N_7651);
nor U10384 (N_10384,N_6126,N_7498);
or U10385 (N_10385,N_8056,N_7008);
and U10386 (N_10386,N_6506,N_9496);
and U10387 (N_10387,N_9372,N_7815);
nand U10388 (N_10388,N_8939,N_5598);
or U10389 (N_10389,N_9695,N_5978);
xor U10390 (N_10390,N_6812,N_5752);
or U10391 (N_10391,N_9458,N_9342);
xnor U10392 (N_10392,N_5944,N_5470);
nand U10393 (N_10393,N_5208,N_7457);
nor U10394 (N_10394,N_5126,N_9676);
and U10395 (N_10395,N_9940,N_7290);
or U10396 (N_10396,N_5946,N_7371);
xor U10397 (N_10397,N_6669,N_7695);
nor U10398 (N_10398,N_9107,N_7607);
or U10399 (N_10399,N_6908,N_8063);
xnor U10400 (N_10400,N_7857,N_7496);
nor U10401 (N_10401,N_6391,N_7456);
xor U10402 (N_10402,N_9385,N_5182);
or U10403 (N_10403,N_7404,N_8256);
nand U10404 (N_10404,N_7591,N_6317);
and U10405 (N_10405,N_8702,N_5717);
nor U10406 (N_10406,N_7627,N_6663);
xor U10407 (N_10407,N_5267,N_9413);
and U10408 (N_10408,N_8599,N_7021);
or U10409 (N_10409,N_9597,N_7270);
nand U10410 (N_10410,N_7061,N_9562);
xor U10411 (N_10411,N_8138,N_5813);
xor U10412 (N_10412,N_5157,N_5391);
or U10413 (N_10413,N_5561,N_8319);
xor U10414 (N_10414,N_6042,N_6182);
nor U10415 (N_10415,N_8001,N_7977);
or U10416 (N_10416,N_7601,N_5154);
nand U10417 (N_10417,N_9784,N_6300);
nor U10418 (N_10418,N_6762,N_9403);
and U10419 (N_10419,N_5278,N_7177);
or U10420 (N_10420,N_9398,N_6243);
nand U10421 (N_10421,N_8737,N_7423);
nor U10422 (N_10422,N_5402,N_9050);
nand U10423 (N_10423,N_9427,N_8523);
or U10424 (N_10424,N_9209,N_8406);
xor U10425 (N_10425,N_9049,N_5217);
nor U10426 (N_10426,N_7668,N_7882);
or U10427 (N_10427,N_9015,N_6339);
nand U10428 (N_10428,N_9492,N_6573);
or U10429 (N_10429,N_9065,N_5738);
xor U10430 (N_10430,N_8224,N_8462);
nand U10431 (N_10431,N_8584,N_5861);
or U10432 (N_10432,N_9174,N_5106);
or U10433 (N_10433,N_8578,N_5438);
nand U10434 (N_10434,N_8458,N_8438);
nand U10435 (N_10435,N_9898,N_8325);
nand U10436 (N_10436,N_8813,N_8440);
or U10437 (N_10437,N_6158,N_9011);
nor U10438 (N_10438,N_6591,N_5675);
xor U10439 (N_10439,N_8327,N_8719);
nand U10440 (N_10440,N_9468,N_6835);
and U10441 (N_10441,N_6114,N_7309);
xor U10442 (N_10442,N_6510,N_9903);
or U10443 (N_10443,N_8808,N_8400);
nand U10444 (N_10444,N_8913,N_8942);
or U10445 (N_10445,N_7770,N_5566);
xnor U10446 (N_10446,N_9020,N_5479);
xor U10447 (N_10447,N_5840,N_5196);
xor U10448 (N_10448,N_5612,N_9499);
nor U10449 (N_10449,N_7157,N_9963);
nor U10450 (N_10450,N_5094,N_6823);
nor U10451 (N_10451,N_5791,N_9757);
nor U10452 (N_10452,N_5742,N_8214);
and U10453 (N_10453,N_9286,N_5608);
nor U10454 (N_10454,N_9195,N_5460);
nand U10455 (N_10455,N_9009,N_8647);
and U10456 (N_10456,N_9906,N_8216);
and U10457 (N_10457,N_7988,N_6690);
nor U10458 (N_10458,N_5443,N_7310);
nor U10459 (N_10459,N_5171,N_8257);
nand U10460 (N_10460,N_8992,N_6797);
or U10461 (N_10461,N_9257,N_7835);
or U10462 (N_10462,N_7828,N_7804);
xnor U10463 (N_10463,N_8077,N_8279);
xor U10464 (N_10464,N_7474,N_9813);
nor U10465 (N_10465,N_9640,N_8016);
nor U10466 (N_10466,N_7612,N_9160);
and U10467 (N_10467,N_8802,N_8116);
nor U10468 (N_10468,N_7118,N_5090);
or U10469 (N_10469,N_7161,N_7805);
or U10470 (N_10470,N_8300,N_7603);
xor U10471 (N_10471,N_5281,N_8725);
xnor U10472 (N_10472,N_7889,N_9488);
xnor U10473 (N_10473,N_9983,N_9833);
nor U10474 (N_10474,N_9871,N_5504);
xnor U10475 (N_10475,N_5775,N_8809);
nand U10476 (N_10476,N_8480,N_7774);
or U10477 (N_10477,N_9979,N_9254);
nor U10478 (N_10478,N_7059,N_6340);
nor U10479 (N_10479,N_5565,N_6607);
or U10480 (N_10480,N_6304,N_8186);
nand U10481 (N_10481,N_5229,N_5007);
nor U10482 (N_10482,N_7257,N_8078);
xor U10483 (N_10483,N_8923,N_6785);
nor U10484 (N_10484,N_6477,N_8329);
nand U10485 (N_10485,N_6667,N_8741);
xnor U10486 (N_10486,N_5673,N_5329);
or U10487 (N_10487,N_6356,N_8015);
or U10488 (N_10488,N_8541,N_7866);
xor U10489 (N_10489,N_7097,N_5080);
or U10490 (N_10490,N_9142,N_7822);
nand U10491 (N_10491,N_9760,N_9075);
nor U10492 (N_10492,N_6965,N_5368);
xor U10493 (N_10493,N_6640,N_6394);
and U10494 (N_10494,N_5595,N_9971);
and U10495 (N_10495,N_9453,N_9400);
nor U10496 (N_10496,N_5140,N_9781);
nand U10497 (N_10497,N_8379,N_5692);
nand U10498 (N_10498,N_8201,N_6701);
nand U10499 (N_10499,N_6733,N_6705);
nand U10500 (N_10500,N_7974,N_8441);
nand U10501 (N_10501,N_5800,N_5064);
xor U10502 (N_10502,N_6221,N_7821);
xnor U10503 (N_10503,N_8463,N_9875);
and U10504 (N_10504,N_5514,N_5950);
nor U10505 (N_10505,N_9134,N_9666);
nor U10506 (N_10506,N_7949,N_7004);
xor U10507 (N_10507,N_8993,N_8229);
and U10508 (N_10508,N_8635,N_7944);
or U10509 (N_10509,N_9958,N_6283);
or U10510 (N_10510,N_8049,N_6933);
nor U10511 (N_10511,N_7620,N_8751);
nor U10512 (N_10512,N_5367,N_8213);
xor U10513 (N_10513,N_9082,N_5545);
xor U10514 (N_10514,N_7636,N_8101);
xor U10515 (N_10515,N_8046,N_8274);
xor U10516 (N_10516,N_5985,N_5387);
xnor U10517 (N_10517,N_6155,N_9192);
nor U10518 (N_10518,N_6914,N_8220);
xnor U10519 (N_10519,N_9876,N_8894);
xnor U10520 (N_10520,N_6173,N_7524);
xor U10521 (N_10521,N_5351,N_5525);
xor U10522 (N_10522,N_8985,N_9439);
nor U10523 (N_10523,N_8999,N_9503);
and U10524 (N_10524,N_6267,N_9516);
xnor U10525 (N_10525,N_6465,N_5805);
xnor U10526 (N_10526,N_9543,N_9487);
nand U10527 (N_10527,N_6832,N_6061);
nand U10528 (N_10528,N_9684,N_8806);
nor U10529 (N_10529,N_8944,N_6769);
nand U10530 (N_10530,N_5502,N_9846);
nand U10531 (N_10531,N_7441,N_7359);
nor U10532 (N_10532,N_5256,N_6024);
and U10533 (N_10533,N_7895,N_7096);
nor U10534 (N_10534,N_8585,N_6735);
nor U10535 (N_10535,N_6217,N_8347);
nand U10536 (N_10536,N_6749,N_6943);
nand U10537 (N_10537,N_5109,N_6856);
or U10538 (N_10538,N_7225,N_9698);
nand U10539 (N_10539,N_8222,N_5350);
nand U10540 (N_10540,N_6621,N_7657);
and U10541 (N_10541,N_8528,N_6315);
nand U10542 (N_10542,N_5986,N_5980);
nor U10543 (N_10543,N_8413,N_7304);
or U10544 (N_10544,N_8795,N_6668);
nor U10545 (N_10545,N_5169,N_8425);
nor U10546 (N_10546,N_8582,N_6952);
and U10547 (N_10547,N_7911,N_7064);
or U10548 (N_10548,N_7995,N_7009);
nand U10549 (N_10549,N_6689,N_8152);
nand U10550 (N_10550,N_7996,N_6020);
nand U10551 (N_10551,N_5835,N_9076);
or U10552 (N_10552,N_9063,N_9305);
or U10553 (N_10553,N_5365,N_6105);
nand U10554 (N_10554,N_7216,N_8552);
or U10555 (N_10555,N_7810,N_7231);
xor U10556 (N_10556,N_8509,N_9019);
xor U10557 (N_10557,N_8073,N_9682);
or U10558 (N_10558,N_8766,N_7513);
or U10559 (N_10559,N_6312,N_7743);
and U10560 (N_10560,N_5793,N_8877);
nand U10561 (N_10561,N_6613,N_6784);
nor U10562 (N_10562,N_5035,N_7834);
and U10563 (N_10563,N_6687,N_6224);
nand U10564 (N_10564,N_7106,N_8284);
nand U10565 (N_10565,N_8531,N_5767);
or U10566 (N_10566,N_5760,N_9629);
nand U10567 (N_10567,N_8856,N_7132);
xnor U10568 (N_10568,N_7572,N_9114);
nor U10569 (N_10569,N_8094,N_9529);
and U10570 (N_10570,N_6494,N_9447);
and U10571 (N_10571,N_7168,N_5293);
nor U10572 (N_10572,N_6098,N_7274);
nand U10573 (N_10573,N_6828,N_7739);
xnor U10574 (N_10574,N_5761,N_9375);
or U10575 (N_10575,N_7146,N_9036);
and U10576 (N_10576,N_5902,N_6692);
and U10577 (N_10577,N_7535,N_7013);
nand U10578 (N_10578,N_8916,N_8255);
or U10579 (N_10579,N_7069,N_8601);
xor U10580 (N_10580,N_6811,N_6163);
and U10581 (N_10581,N_5718,N_9494);
nor U10582 (N_10582,N_6392,N_9504);
and U10583 (N_10583,N_8234,N_9317);
xor U10584 (N_10584,N_7392,N_5086);
nand U10585 (N_10585,N_7232,N_6629);
xor U10586 (N_10586,N_8037,N_6260);
or U10587 (N_10587,N_8909,N_7172);
and U10588 (N_10588,N_5927,N_8434);
nor U10589 (N_10589,N_5436,N_5936);
or U10590 (N_10590,N_6052,N_8431);
and U10591 (N_10591,N_9601,N_7098);
xnor U10592 (N_10592,N_9949,N_7105);
or U10593 (N_10593,N_9460,N_8654);
xnor U10594 (N_10594,N_7311,N_5932);
nand U10595 (N_10595,N_9344,N_5275);
nor U10596 (N_10596,N_7324,N_9739);
or U10597 (N_10597,N_6417,N_5749);
or U10598 (N_10598,N_9423,N_6387);
or U10599 (N_10599,N_5853,N_8059);
nand U10600 (N_10600,N_5569,N_9177);
xnor U10601 (N_10601,N_6702,N_9264);
nor U10602 (N_10602,N_5520,N_9515);
xnor U10603 (N_10603,N_6148,N_5482);
xnor U10604 (N_10604,N_7465,N_9961);
or U10605 (N_10605,N_6463,N_8464);
nand U10606 (N_10606,N_8792,N_6543);
and U10607 (N_10607,N_5150,N_6369);
and U10608 (N_10608,N_8376,N_8362);
or U10609 (N_10609,N_8718,N_9771);
nand U10610 (N_10610,N_6805,N_7903);
and U10611 (N_10611,N_8911,N_6087);
or U10612 (N_10612,N_5105,N_7516);
and U10613 (N_10613,N_7101,N_8814);
or U10614 (N_10614,N_5445,N_7220);
and U10615 (N_10615,N_5883,N_9942);
xor U10616 (N_10616,N_7771,N_8842);
xor U10617 (N_10617,N_5231,N_8930);
xnor U10618 (N_10618,N_6482,N_5758);
nor U10619 (N_10619,N_6723,N_5316);
nand U10620 (N_10620,N_5123,N_5607);
nor U10621 (N_10621,N_9914,N_5594);
xnor U10622 (N_10622,N_5476,N_5578);
nand U10623 (N_10623,N_7035,N_7015);
nor U10624 (N_10624,N_5576,N_8961);
and U10625 (N_10625,N_7686,N_9891);
and U10626 (N_10626,N_9249,N_7224);
or U10627 (N_10627,N_7071,N_7999);
xnor U10628 (N_10628,N_9255,N_5818);
nor U10629 (N_10629,N_6567,N_6225);
or U10630 (N_10630,N_7756,N_6334);
or U10631 (N_10631,N_5972,N_9261);
nor U10632 (N_10632,N_8208,N_9568);
and U10633 (N_10633,N_7208,N_6608);
or U10634 (N_10634,N_8295,N_5191);
and U10635 (N_10635,N_8778,N_7002);
and U10636 (N_10636,N_6980,N_8810);
xnor U10637 (N_10637,N_7728,N_8024);
and U10638 (N_10638,N_5651,N_6354);
nor U10639 (N_10639,N_9551,N_6095);
or U10640 (N_10640,N_9387,N_9383);
nor U10641 (N_10641,N_7831,N_9557);
and U10642 (N_10642,N_8120,N_6374);
nor U10643 (N_10643,N_9974,N_9386);
xnor U10644 (N_10644,N_7823,N_9755);
and U10645 (N_10645,N_6873,N_7122);
xnor U10646 (N_10646,N_7734,N_8949);
nand U10647 (N_10647,N_8081,N_9191);
xor U10648 (N_10648,N_9039,N_7349);
xnor U10649 (N_10649,N_8489,N_8282);
or U10650 (N_10650,N_6750,N_6829);
and U10651 (N_10651,N_5396,N_7426);
or U10652 (N_10652,N_6695,N_8429);
and U10653 (N_10653,N_8010,N_6593);
xnor U10654 (N_10654,N_9572,N_6803);
nor U10655 (N_10655,N_8385,N_6115);
or U10656 (N_10656,N_7745,N_5424);
and U10657 (N_10657,N_8217,N_5395);
nor U10658 (N_10658,N_6531,N_6874);
and U10659 (N_10659,N_7946,N_6331);
nand U10660 (N_10660,N_7779,N_8952);
nand U10661 (N_10661,N_7124,N_5725);
or U10662 (N_10662,N_9148,N_5046);
nand U10663 (N_10663,N_7322,N_6342);
xnor U10664 (N_10664,N_7275,N_8620);
xnor U10665 (N_10665,N_5099,N_8733);
or U10666 (N_10666,N_8764,N_9098);
nand U10667 (N_10667,N_8218,N_8176);
nand U10668 (N_10668,N_8984,N_6363);
and U10669 (N_10669,N_8090,N_6906);
or U10670 (N_10670,N_8158,N_9399);
and U10671 (N_10671,N_5253,N_9357);
or U10672 (N_10672,N_9426,N_9175);
nand U10673 (N_10673,N_6108,N_6639);
nor U10674 (N_10674,N_7588,N_5240);
and U10675 (N_10675,N_8607,N_6201);
xnor U10676 (N_10676,N_6530,N_8897);
nor U10677 (N_10677,N_7545,N_8676);
nand U10678 (N_10678,N_5721,N_9941);
nand U10679 (N_10679,N_9222,N_8483);
and U10680 (N_10680,N_7869,N_6824);
or U10681 (N_10681,N_6119,N_6019);
nand U10682 (N_10682,N_7407,N_6661);
nand U10683 (N_10683,N_6133,N_9542);
xor U10684 (N_10684,N_5659,N_7387);
or U10685 (N_10685,N_6845,N_6526);
xor U10686 (N_10686,N_8439,N_7490);
and U10687 (N_10687,N_9186,N_7960);
xnor U10688 (N_10688,N_9294,N_8069);
nor U10689 (N_10689,N_6954,N_5954);
nand U10690 (N_10690,N_5063,N_8287);
or U10691 (N_10691,N_9649,N_6301);
nor U10692 (N_10692,N_7372,N_8783);
xor U10693 (N_10693,N_8270,N_9296);
and U10694 (N_10694,N_8210,N_9792);
and U10695 (N_10695,N_9657,N_9106);
or U10696 (N_10696,N_8307,N_7425);
or U10697 (N_10697,N_8247,N_6085);
nand U10698 (N_10698,N_5854,N_6813);
or U10699 (N_10699,N_8745,N_7078);
or U10700 (N_10700,N_9326,N_6588);
or U10701 (N_10701,N_5713,N_5494);
nor U10702 (N_10702,N_7452,N_9775);
or U10703 (N_10703,N_5137,N_6743);
nor U10704 (N_10704,N_8497,N_6165);
nor U10705 (N_10705,N_6546,N_5159);
xnor U10706 (N_10706,N_8818,N_8227);
nor U10707 (N_10707,N_7072,N_9531);
xnor U10708 (N_10708,N_5784,N_5441);
or U10709 (N_10709,N_7583,N_5678);
or U10710 (N_10710,N_5459,N_6447);
nor U10711 (N_10711,N_9823,N_9856);
and U10712 (N_10712,N_9408,N_9776);
and U10713 (N_10713,N_5409,N_8891);
and U10714 (N_10714,N_9841,N_6715);
or U10715 (N_10715,N_8790,N_5702);
or U10716 (N_10716,N_8890,N_6825);
xor U10717 (N_10717,N_6021,N_8313);
nor U10718 (N_10718,N_8470,N_6292);
or U10719 (N_10719,N_6441,N_8093);
nor U10720 (N_10720,N_8576,N_7840);
nor U10721 (N_10721,N_6058,N_8109);
xnor U10722 (N_10722,N_5694,N_5601);
nor U10723 (N_10723,N_8242,N_5771);
and U10724 (N_10724,N_5929,N_8603);
xor U10725 (N_10725,N_8102,N_5820);
and U10726 (N_10726,N_8478,N_6581);
and U10727 (N_10727,N_9907,N_9622);
nand U10728 (N_10728,N_5397,N_5745);
nand U10729 (N_10729,N_7991,N_5628);
nor U10730 (N_10730,N_5687,N_8349);
nand U10731 (N_10731,N_5575,N_6009);
nand U10732 (N_10732,N_6804,N_5735);
nor U10733 (N_10733,N_6575,N_5039);
and U10734 (N_10734,N_9489,N_6879);
or U10735 (N_10735,N_6424,N_7204);
or U10736 (N_10736,N_9889,N_9648);
nand U10737 (N_10737,N_6467,N_6488);
xor U10738 (N_10738,N_9915,N_8351);
nand U10739 (N_10739,N_7850,N_6036);
nor U10740 (N_10740,N_8038,N_5188);
nor U10741 (N_10741,N_5597,N_6590);
and U10742 (N_10742,N_6209,N_7777);
nand U10743 (N_10743,N_6594,N_5005);
nor U10744 (N_10744,N_8354,N_5404);
or U10745 (N_10745,N_9262,N_6307);
nand U10746 (N_10746,N_5399,N_6184);
xor U10747 (N_10747,N_9603,N_5529);
nand U10748 (N_10748,N_8335,N_5327);
and U10749 (N_10749,N_9302,N_8996);
and U10750 (N_10750,N_7243,N_6039);
or U10751 (N_10751,N_6380,N_6205);
or U10752 (N_10752,N_8278,N_8881);
xor U10753 (N_10753,N_6323,N_7481);
nor U10754 (N_10754,N_9179,N_8002);
and U10755 (N_10755,N_8233,N_9618);
nand U10756 (N_10756,N_6513,N_8143);
xor U10757 (N_10757,N_5363,N_5720);
nand U10758 (N_10758,N_9451,N_9725);
nand U10759 (N_10759,N_8051,N_7816);
nor U10760 (N_10760,N_8573,N_8110);
nand U10761 (N_10761,N_8862,N_7958);
or U10762 (N_10762,N_9247,N_6571);
xor U10763 (N_10763,N_9214,N_7282);
nor U10764 (N_10764,N_7112,N_9985);
xnor U10765 (N_10765,N_7842,N_7199);
xnor U10766 (N_10766,N_6517,N_7336);
xor U10767 (N_10767,N_7147,N_5266);
and U10768 (N_10768,N_5500,N_5091);
xnor U10769 (N_10769,N_6237,N_8065);
or U10770 (N_10770,N_6332,N_6489);
and U10771 (N_10771,N_9718,N_6658);
nand U10772 (N_10772,N_9055,N_5497);
xor U10773 (N_10773,N_5801,N_7354);
and U10774 (N_10774,N_9647,N_7813);
and U10775 (N_10775,N_7475,N_8029);
or U10776 (N_10776,N_6361,N_8389);
xnor U10777 (N_10777,N_5683,N_7185);
nand U10778 (N_10778,N_8600,N_9465);
nand U10779 (N_10779,N_8203,N_9785);
nor U10780 (N_10780,N_5622,N_6984);
nor U10781 (N_10781,N_8511,N_8023);
xnor U10782 (N_10782,N_8791,N_5269);
and U10783 (N_10783,N_7409,N_5499);
and U10784 (N_10784,N_7608,N_8987);
or U10785 (N_10785,N_9592,N_8717);
nor U10786 (N_10786,N_9818,N_9817);
nand U10787 (N_10787,N_7876,N_5516);
xnor U10788 (N_10788,N_8020,N_9268);
nand U10789 (N_10789,N_5238,N_6570);
nor U10790 (N_10790,N_5284,N_8488);
nand U10791 (N_10791,N_8765,N_5075);
or U10792 (N_10792,N_7389,N_6566);
nand U10793 (N_10793,N_7554,N_9599);
nor U10794 (N_10794,N_6903,N_8968);
xnor U10795 (N_10795,N_8241,N_7807);
nor U10796 (N_10796,N_7528,N_6328);
nand U10797 (N_10797,N_7320,N_6602);
xor U10798 (N_10798,N_8199,N_8340);
and U10799 (N_10799,N_5332,N_8940);
or U10800 (N_10800,N_9128,N_5746);
xor U10801 (N_10801,N_9935,N_8753);
nor U10802 (N_10802,N_6294,N_5059);
xor U10803 (N_10803,N_7058,N_7085);
and U10804 (N_10804,N_8000,N_5430);
nor U10805 (N_10805,N_8378,N_9838);
xnor U10806 (N_10806,N_7183,N_6630);
and U10807 (N_10807,N_5828,N_8872);
or U10808 (N_10808,N_9664,N_9580);
and U10809 (N_10809,N_6159,N_5190);
nand U10810 (N_10810,N_6233,N_5061);
or U10811 (N_10811,N_8175,N_7676);
xnor U10812 (N_10812,N_7451,N_9402);
xnor U10813 (N_10813,N_5114,N_5376);
or U10814 (N_10814,N_9396,N_5244);
nor U10815 (N_10815,N_9731,N_7192);
nor U10816 (N_10816,N_7327,N_6870);
nor U10817 (N_10817,N_8346,N_5870);
xnor U10818 (N_10818,N_8865,N_6916);
nor U10819 (N_10819,N_8868,N_9475);
nor U10820 (N_10820,N_8602,N_6207);
and U10821 (N_10821,N_5947,N_9549);
nand U10822 (N_10822,N_6795,N_7624);
nor U10823 (N_10823,N_6345,N_7095);
nand U10824 (N_10824,N_7694,N_8293);
nor U10825 (N_10825,N_8167,N_9980);
xor U10826 (N_10826,N_7126,N_7047);
or U10827 (N_10827,N_5085,N_9441);
or U10828 (N_10828,N_6636,N_7945);
xor U10829 (N_10829,N_8863,N_5769);
nand U10830 (N_10830,N_6093,N_7942);
and U10831 (N_10831,N_8276,N_7941);
xor U10832 (N_10832,N_6427,N_6548);
or U10833 (N_10833,N_9671,N_9239);
or U10834 (N_10834,N_7912,N_7215);
nand U10835 (N_10835,N_6698,N_8269);
nor U10836 (N_10836,N_6820,N_6940);
nor U10837 (N_10837,N_9110,N_6274);
and U10838 (N_10838,N_8098,N_6711);
or U10839 (N_10839,N_6944,N_9054);
or U10840 (N_10840,N_9505,N_6347);
nand U10841 (N_10841,N_9165,N_5104);
nand U10842 (N_10842,N_5903,N_7705);
and U10843 (N_10843,N_8266,N_8317);
and U10844 (N_10844,N_8365,N_6418);
nor U10845 (N_10845,N_8986,N_5264);
nor U10846 (N_10846,N_9913,N_8744);
and U10847 (N_10847,N_6726,N_5180);
or U10848 (N_10848,N_9519,N_7180);
xnor U10849 (N_10849,N_9810,N_7130);
xor U10850 (N_10850,N_8301,N_6665);
nand U10851 (N_10851,N_5875,N_5096);
or U10852 (N_10852,N_9158,N_6926);
nor U10853 (N_10853,N_9552,N_8883);
xnor U10854 (N_10854,N_9349,N_7644);
xor U10855 (N_10855,N_8886,N_6990);
xor U10856 (N_10856,N_6863,N_7547);
or U10857 (N_10857,N_7843,N_5920);
xor U10858 (N_10858,N_9450,N_6343);
nand U10859 (N_10859,N_8712,N_9922);
nor U10860 (N_10860,N_5309,N_5921);
nand U10861 (N_10861,N_9520,N_7947);
nor U10862 (N_10862,N_5380,N_6234);
nor U10863 (N_10863,N_6877,N_6407);
or U10864 (N_10864,N_5925,N_8843);
nand U10865 (N_10865,N_7765,N_9721);
nor U10866 (N_10866,N_5016,N_8852);
xnor U10867 (N_10867,N_7596,N_6261);
nor U10868 (N_10868,N_8639,N_9183);
nand U10869 (N_10869,N_8671,N_5221);
or U10870 (N_10870,N_5458,N_9533);
xnor U10871 (N_10871,N_5556,N_7174);
nand U10872 (N_10872,N_7019,N_5741);
nand U10873 (N_10873,N_9072,N_6552);
and U10874 (N_10874,N_6844,N_9238);
nand U10875 (N_10875,N_5279,N_8950);
nor U10876 (N_10876,N_8396,N_5969);
xor U10877 (N_10877,N_5295,N_6007);
nor U10878 (N_10878,N_9256,N_7250);
nor U10879 (N_10879,N_6616,N_9920);
nand U10880 (N_10880,N_9987,N_7530);
xnor U10881 (N_10881,N_5650,N_9703);
nand U10882 (N_10882,N_9314,N_7748);
and U10883 (N_10883,N_6547,N_6617);
or U10884 (N_10884,N_9352,N_9613);
or U10885 (N_10885,N_5492,N_7824);
nand U10886 (N_10886,N_9125,N_6922);
nand U10887 (N_10887,N_9373,N_6239);
xnor U10888 (N_10888,N_6434,N_5937);
nand U10889 (N_10889,N_5025,N_5161);
xor U10890 (N_10890,N_6041,N_6909);
nand U10891 (N_10891,N_6067,N_7573);
or U10892 (N_10892,N_7347,N_5881);
nor U10893 (N_10893,N_8723,N_5648);
xor U10894 (N_10894,N_7348,N_5939);
nor U10895 (N_10895,N_7419,N_9865);
or U10896 (N_10896,N_5070,N_8493);
or U10897 (N_10897,N_5076,N_7652);
xnor U10898 (N_10898,N_9476,N_7160);
or U10899 (N_10899,N_8524,N_5945);
and U10900 (N_10900,N_7241,N_6808);
and U10901 (N_10901,N_6898,N_5652);
nor U10902 (N_10902,N_5773,N_5289);
or U10903 (N_10903,N_9769,N_8453);
and U10904 (N_10904,N_8035,N_6135);
and U10905 (N_10905,N_9270,N_5863);
nand U10906 (N_10906,N_5301,N_6378);
and U10907 (N_10907,N_8350,N_9794);
and U10908 (N_10908,N_8290,N_8661);
nor U10909 (N_10909,N_9812,N_7206);
and U10910 (N_10910,N_8082,N_9006);
xnor U10911 (N_10911,N_7153,N_6450);
nor U10912 (N_10912,N_8517,N_6961);
nand U10913 (N_10913,N_5177,N_8975);
nor U10914 (N_10914,N_7890,N_5789);
or U10915 (N_10915,N_6550,N_8409);
nand U10916 (N_10916,N_6244,N_9113);
nor U10917 (N_10917,N_7193,N_6102);
xnor U10918 (N_10918,N_6753,N_7793);
and U10919 (N_10919,N_9936,N_9131);
or U10920 (N_10920,N_5890,N_8544);
and U10921 (N_10921,N_8789,N_7221);
nor U10922 (N_10922,N_9136,N_5068);
xor U10923 (N_10923,N_7622,N_5260);
and U10924 (N_10924,N_7081,N_8253);
nand U10925 (N_10925,N_9321,N_5635);
xor U10926 (N_10926,N_5783,N_5354);
and U10927 (N_10927,N_9616,N_6064);
nor U10928 (N_10928,N_6490,N_6131);
nor U10929 (N_10929,N_9320,N_9438);
and U10930 (N_10930,N_9700,N_7640);
or U10931 (N_10931,N_8500,N_8180);
or U10932 (N_10932,N_9144,N_5273);
nand U10933 (N_10933,N_5661,N_9060);
nor U10934 (N_10934,N_5239,N_6911);
nor U10935 (N_10935,N_5342,N_9692);
or U10936 (N_10936,N_5344,N_5535);
xnor U10937 (N_10937,N_5693,N_5193);
xnor U10938 (N_10938,N_7131,N_9594);
nor U10939 (N_10939,N_7558,N_9127);
nand U10940 (N_10940,N_8779,N_9716);
or U10941 (N_10941,N_8264,N_6605);
xor U10942 (N_10942,N_6606,N_6080);
nand U10943 (N_10943,N_6144,N_5414);
xor U10944 (N_10944,N_8084,N_5765);
or U10945 (N_10945,N_7795,N_6250);
xor U10946 (N_10946,N_5871,N_8505);
nor U10947 (N_10947,N_6794,N_8892);
or U10948 (N_10948,N_9733,N_8204);
or U10949 (N_10949,N_7794,N_8688);
or U10950 (N_10950,N_9585,N_6132);
xnor U10951 (N_10951,N_9206,N_6263);
nand U10952 (N_10952,N_7334,N_7827);
nand U10953 (N_10953,N_5172,N_6484);
or U10954 (N_10954,N_9743,N_8352);
xor U10955 (N_10955,N_6710,N_9003);
nor U10956 (N_10956,N_8165,N_6686);
nand U10957 (N_10957,N_9442,N_5590);
and U10958 (N_10958,N_5047,N_9787);
xnor U10959 (N_10959,N_8104,N_9267);
nor U10960 (N_10960,N_7614,N_9853);
nor U10961 (N_10961,N_6744,N_9184);
or U10962 (N_10962,N_7117,N_5930);
nor U10963 (N_10963,N_7565,N_6284);
nand U10964 (N_10964,N_6998,N_8320);
nand U10965 (N_10965,N_8387,N_5503);
nand U10966 (N_10966,N_6627,N_9341);
nor U10967 (N_10967,N_7350,N_8760);
and U10968 (N_10968,N_5699,N_9752);
nand U10969 (N_10969,N_6635,N_7345);
and U10970 (N_10970,N_5655,N_5226);
and U10971 (N_10971,N_7090,N_9546);
and U10972 (N_10972,N_6223,N_5370);
or U10973 (N_10973,N_8936,N_5743);
and U10974 (N_10974,N_9048,N_9678);
nor U10975 (N_10975,N_7802,N_6322);
nor U10976 (N_10976,N_7680,N_6987);
xor U10977 (N_10977,N_9130,N_6318);
and U10978 (N_10978,N_5916,N_5953);
nand U10979 (N_10979,N_5254,N_6218);
or U10980 (N_10980,N_6195,N_5753);
nor U10981 (N_10981,N_7609,N_7277);
xnor U10982 (N_10982,N_9151,N_7502);
nand U10983 (N_10983,N_6788,N_6964);
nand U10984 (N_10984,N_9972,N_9071);
nor U10985 (N_10985,N_6458,N_8099);
nor U10986 (N_10986,N_8388,N_6674);
or U10987 (N_10987,N_8454,N_8934);
nor U10988 (N_10988,N_5919,N_5014);
nor U10989 (N_10989,N_8032,N_7954);
and U10990 (N_10990,N_7182,N_6583);
xor U10991 (N_10991,N_8011,N_9619);
nand U10992 (N_10992,N_5119,N_7142);
nor U10993 (N_10993,N_6029,N_7784);
nand U10994 (N_10994,N_7760,N_8731);
nand U10995 (N_10995,N_5961,N_9029);
nand U10996 (N_10996,N_6178,N_9773);
nand U10997 (N_10997,N_7696,N_5072);
nor U10998 (N_10998,N_9545,N_9611);
and U10999 (N_10999,N_7769,N_9831);
nor U11000 (N_11000,N_8071,N_6511);
and U11001 (N_11001,N_8529,N_5519);
nor U11002 (N_11002,N_9461,N_7301);
nor U11003 (N_11003,N_8358,N_8969);
nor U11004 (N_11004,N_7602,N_6281);
xor U11005 (N_11005,N_9181,N_8776);
nand U11006 (N_11006,N_5842,N_5125);
or U11007 (N_11007,N_7679,N_9804);
and U11008 (N_11008,N_8867,N_6203);
xor U11009 (N_11009,N_6561,N_6187);
and U11010 (N_11010,N_5174,N_9953);
or U11011 (N_11011,N_8248,N_9446);
nor U11012 (N_11012,N_5055,N_9469);
and U11013 (N_11013,N_8928,N_9203);
xor U11014 (N_11014,N_9701,N_9207);
or U11015 (N_11015,N_8774,N_5733);
xor U11016 (N_11016,N_7593,N_6188);
or U11017 (N_11017,N_7462,N_5833);
or U11018 (N_11018,N_5657,N_5089);
and U11019 (N_11019,N_6953,N_8589);
xnor U11020 (N_11020,N_6742,N_8981);
or U11021 (N_11021,N_7955,N_6568);
nor U11022 (N_11022,N_7388,N_9807);
or U11023 (N_11023,N_5403,N_6978);
and U11024 (N_11024,N_9863,N_7361);
nor U11025 (N_11025,N_6875,N_5400);
nor U11026 (N_11026,N_7757,N_5568);
nand U11027 (N_11027,N_9522,N_8633);
xnor U11028 (N_11028,N_7540,N_8915);
xor U11029 (N_11029,N_8514,N_7148);
nand U11030 (N_11030,N_6939,N_5646);
or U11031 (N_11031,N_7660,N_7753);
and U11032 (N_11032,N_9869,N_6551);
or U11033 (N_11033,N_8162,N_8331);
nand U11034 (N_11034,N_7370,N_6049);
nand U11035 (N_11035,N_5906,N_6246);
or U11036 (N_11036,N_8231,N_8832);
and U11037 (N_11037,N_5855,N_9237);
nand U11038 (N_11038,N_7736,N_8617);
xnor U11039 (N_11039,N_5747,N_5286);
nand U11040 (N_11040,N_7291,N_8106);
nand U11041 (N_11041,N_9673,N_7119);
xnor U11042 (N_11042,N_6737,N_5866);
nand U11043 (N_11043,N_9510,N_6198);
nand U11044 (N_11044,N_7102,N_7515);
or U11045 (N_11045,N_6889,N_5762);
nor U11046 (N_11046,N_9719,N_8858);
xor U11047 (N_11047,N_9897,N_8926);
and U11048 (N_11048,N_6724,N_9777);
xor U11049 (N_11049,N_9602,N_6923);
and U11050 (N_11050,N_9679,N_7979);
and U11051 (N_11051,N_9353,N_5156);
xor U11052 (N_11052,N_9119,N_8726);
nand U11053 (N_11053,N_8824,N_5685);
nor U11054 (N_11054,N_9728,N_5756);
xor U11055 (N_11055,N_9464,N_9281);
and U11056 (N_11056,N_5792,N_6066);
nor U11057 (N_11057,N_6699,N_7285);
nor U11058 (N_11058,N_6834,N_9829);
nor U11059 (N_11059,N_7093,N_5987);
or U11060 (N_11060,N_8465,N_8836);
xnor U11061 (N_11061,N_8026,N_5095);
or U11062 (N_11062,N_5379,N_9726);
and U11063 (N_11063,N_9218,N_6791);
nor U11064 (N_11064,N_6242,N_7750);
or U11065 (N_11065,N_6910,N_5195);
nor U11066 (N_11066,N_9851,N_8137);
xnor U11067 (N_11067,N_5324,N_9284);
nor U11068 (N_11068,N_8160,N_9843);
xnor U11069 (N_11069,N_7900,N_8402);
and U11070 (N_11070,N_8139,N_6035);
and U11071 (N_11071,N_5423,N_5359);
nor U11072 (N_11072,N_8271,N_8938);
or U11073 (N_11073,N_9156,N_7416);
xor U11074 (N_11074,N_7934,N_8540);
or U11075 (N_11075,N_8321,N_5203);
and U11076 (N_11076,N_8324,N_7508);
nor U11077 (N_11077,N_6498,N_8833);
or U11078 (N_11078,N_7440,N_5065);
xor U11079 (N_11079,N_8135,N_7152);
nor U11080 (N_11080,N_5415,N_5146);
nand U11081 (N_11081,N_9235,N_7543);
nor U11082 (N_11082,N_5732,N_6937);
or U11083 (N_11083,N_7091,N_6393);
or U11084 (N_11084,N_6525,N_5166);
xor U11085 (N_11085,N_5302,N_5766);
or U11086 (N_11086,N_7673,N_5970);
xnor U11087 (N_11087,N_9962,N_9643);
nand U11088 (N_11088,N_5757,N_7248);
and U11089 (N_11089,N_6537,N_8182);
xor U11090 (N_11090,N_8922,N_5807);
or U11091 (N_11091,N_9662,N_7684);
and U11092 (N_11092,N_7262,N_9436);
xor U11093 (N_11093,N_5864,N_7639);
xor U11094 (N_11094,N_7186,N_5979);
or U11095 (N_11095,N_6846,N_5318);
or U11096 (N_11096,N_6761,N_7051);
and U11097 (N_11097,N_6770,N_7212);
nor U11098 (N_11098,N_7621,N_9141);
xnor U11099 (N_11099,N_7115,N_6679);
and U11100 (N_11100,N_8538,N_8142);
and U11101 (N_11101,N_7406,N_6309);
or U11102 (N_11102,N_9371,N_5495);
or U11103 (N_11103,N_5876,N_7967);
nand U11104 (N_11104,N_7940,N_7272);
or U11105 (N_11105,N_9588,N_9042);
and U11106 (N_11106,N_7518,N_5898);
or U11107 (N_11107,N_9041,N_7541);
or U11108 (N_11108,N_6082,N_7580);
nand U11109 (N_11109,N_6754,N_8460);
nand U11110 (N_11110,N_5037,N_8275);
nand U11111 (N_11111,N_8355,N_5951);
nor U11112 (N_11112,N_7237,N_6134);
xor U11113 (N_11113,N_8674,N_5209);
nand U11114 (N_11114,N_8706,N_6431);
xor U11115 (N_11115,N_6295,N_8920);
and U11116 (N_11116,N_9300,N_8796);
xnor U11117 (N_11117,N_9178,N_8306);
or U11118 (N_11118,N_9593,N_9947);
nor U11119 (N_11119,N_8391,N_8079);
and U11120 (N_11120,N_6880,N_9824);
and U11121 (N_11121,N_6247,N_6579);
and U11122 (N_11122,N_9230,N_9811);
nor U11123 (N_11123,N_8025,N_6174);
or U11124 (N_11124,N_6852,N_9053);
nor U11125 (N_11125,N_9038,N_5834);
or U11126 (N_11126,N_8061,N_6068);
nand U11127 (N_11127,N_9525,N_9358);
or U11128 (N_11128,N_6983,N_7520);
nor U11129 (N_11129,N_5481,N_9007);
xnor U11130 (N_11130,N_8522,N_5609);
xnor U11131 (N_11131,N_6366,N_8134);
nand U11132 (N_11132,N_8597,N_7381);
nand U11133 (N_11133,N_8131,N_8471);
xor U11134 (N_11134,N_8957,N_6214);
or U11135 (N_11135,N_8958,N_6254);
xor U11136 (N_11136,N_8788,N_9879);
nand U11137 (N_11137,N_5473,N_6337);
or U11138 (N_11138,N_7897,N_5054);
xor U11139 (N_11139,N_5338,N_6562);
xnor U11140 (N_11140,N_7658,N_9115);
xnor U11141 (N_11141,N_6582,N_9660);
nor U11142 (N_11142,N_7725,N_7582);
xnor U11143 (N_11143,N_5355,N_8798);
nand U11144 (N_11144,N_6177,N_9123);
nand U11145 (N_11145,N_5689,N_9957);
xor U11146 (N_11146,N_6386,N_8398);
xor U11147 (N_11147,N_8410,N_6015);
nand U11148 (N_11148,N_7233,N_9376);
nand U11149 (N_11149,N_6885,N_8262);
nor U11150 (N_11150,N_5398,N_9534);
nor U11151 (N_11151,N_8628,N_7700);
nor U11152 (N_11152,N_9609,N_9324);
nor U11153 (N_11153,N_7238,N_7128);
xor U11154 (N_11154,N_9538,N_5796);
nand U11155 (N_11155,N_8447,N_5117);
nand U11156 (N_11156,N_8805,N_9401);
and U11157 (N_11157,N_7073,N_5884);
or U11158 (N_11158,N_7218,N_6644);
and U11159 (N_11159,N_8672,N_8508);
and U11160 (N_11160,N_8953,N_7278);
nor U11161 (N_11161,N_9163,N_6503);
and U11162 (N_11162,N_9750,N_7037);
nor U11163 (N_11163,N_9845,N_9934);
xnor U11164 (N_11164,N_9849,N_7075);
xor U11165 (N_11165,N_6228,N_8437);
nand U11166 (N_11166,N_5511,N_6904);
nand U11167 (N_11167,N_7970,N_5823);
or U11168 (N_11168,N_9137,N_5667);
nand U11169 (N_11169,N_7749,N_8121);
and U11170 (N_11170,N_8720,N_8007);
nor U11171 (N_11171,N_6505,N_9738);
nor U11172 (N_11172,N_9058,N_6240);
xor U11173 (N_11173,N_5814,N_5862);
and U11174 (N_11174,N_8967,N_6200);
and U11175 (N_11175,N_9574,N_8132);
and U11176 (N_11176,N_8149,N_8838);
or U11177 (N_11177,N_9644,N_5222);
and U11178 (N_11178,N_6907,N_9425);
and U11179 (N_11179,N_7948,N_7400);
xnor U11180 (N_11180,N_5464,N_5110);
and U11181 (N_11181,N_9734,N_7615);
and U11182 (N_11182,N_8443,N_5737);
and U11183 (N_11183,N_5228,N_5274);
or U11184 (N_11184,N_7662,N_9888);
nand U11185 (N_11185,N_9108,N_6376);
nand U11186 (N_11186,N_8333,N_7133);
or U11187 (N_11187,N_7893,N_8485);
xnor U11188 (N_11188,N_8427,N_7507);
nand U11189 (N_11189,N_7732,N_7149);
nand U11190 (N_11190,N_8853,N_5480);
nand U11191 (N_11191,N_8156,N_6895);
or U11192 (N_11192,N_8067,N_6516);
nand U11193 (N_11193,N_7553,N_9018);
and U11194 (N_11194,N_5779,N_5192);
nand U11195 (N_11195,N_9600,N_5960);
or U11196 (N_11196,N_5084,N_7138);
and U11197 (N_11197,N_7619,N_6137);
and U11198 (N_11198,N_7200,N_5780);
nand U11199 (N_11199,N_7319,N_8373);
nor U11200 (N_11200,N_9266,N_5020);
or U11201 (N_11201,N_7039,N_8356);
or U11202 (N_11202,N_8357,N_8925);
nand U11203 (N_11203,N_7099,N_7683);
nand U11204 (N_11204,N_9636,N_7196);
nor U11205 (N_11205,N_5434,N_9825);
nand U11206 (N_11206,N_8679,N_7189);
xor U11207 (N_11207,N_5326,N_8304);
and U11208 (N_11208,N_5069,N_9332);
nand U11209 (N_11209,N_7194,N_9518);
or U11210 (N_11210,N_8580,N_5006);
nor U11211 (N_11211,N_9292,N_5942);
or U11212 (N_11212,N_6572,N_8245);
nor U11213 (N_11213,N_6062,N_8192);
xnor U11214 (N_11214,N_7026,N_9653);
and U11215 (N_11215,N_7123,N_9668);
and U11216 (N_11216,N_9537,N_7411);
xnor U11217 (N_11217,N_6286,N_7222);
and U11218 (N_11218,N_6789,N_6496);
nor U11219 (N_11219,N_8472,N_8446);
and U11220 (N_11220,N_5477,N_9956);
or U11221 (N_11221,N_7435,N_9786);
nor U11222 (N_11222,N_9244,N_5223);
nor U11223 (N_11223,N_9744,N_9658);
nor U11224 (N_11224,N_8559,N_6040);
or U11225 (N_11225,N_7892,N_5465);
nand U11226 (N_11226,N_8244,N_8631);
nand U11227 (N_11227,N_8370,N_7424);
nand U11228 (N_11228,N_9697,N_5113);
or U11229 (N_11229,N_9112,N_7338);
nor U11230 (N_11230,N_9056,N_6167);
nand U11231 (N_11231,N_6772,N_8228);
nor U11232 (N_11232,N_8759,N_6774);
xor U11233 (N_11233,N_7228,N_9536);
or U11234 (N_11234,N_5341,N_7391);
or U11235 (N_11235,N_5669,N_7546);
nor U11236 (N_11236,N_7715,N_5343);
nor U11237 (N_11237,N_8546,N_5087);
nor U11238 (N_11238,N_8232,N_6222);
and U11239 (N_11239,N_6968,N_6927);
nand U11240 (N_11240,N_7169,N_5167);
nand U11241 (N_11241,N_9176,N_5454);
nand U11242 (N_11242,N_9554,N_6924);
xor U11243 (N_11243,N_7548,N_9874);
and U11244 (N_11244,N_9187,N_7393);
or U11245 (N_11245,N_6786,N_9384);
or U11246 (N_11246,N_9111,N_5056);
and U11247 (N_11247,N_6967,N_9581);
or U11248 (N_11248,N_8964,N_9316);
and U11249 (N_11249,N_6764,N_7862);
xor U11250 (N_11250,N_7517,N_7395);
xnor U11251 (N_11251,N_5533,N_5439);
xnor U11252 (N_11252,N_7641,N_9788);
xor U11253 (N_11253,N_8870,N_7001);
xor U11254 (N_11254,N_7509,N_7767);
and U11255 (N_11255,N_7534,N_5388);
nor U11256 (N_11256,N_6938,N_7826);
xor U11257 (N_11257,N_9740,N_5736);
xnor U11258 (N_11258,N_8342,N_7563);
nand U11259 (N_11259,N_9901,N_5826);
xnor U11260 (N_11260,N_6843,N_5551);
and U11261 (N_11261,N_9369,N_9481);
nor U11262 (N_11262,N_6759,N_6110);
nor U11263 (N_11263,N_8328,N_7068);
or U11264 (N_11264,N_6847,N_9070);
and U11265 (N_11265,N_5618,N_7343);
nor U11266 (N_11266,N_8845,N_9978);
nand U11267 (N_11267,N_5008,N_8168);
or U11268 (N_11268,N_6018,N_8124);
nand U11269 (N_11269,N_7962,N_7510);
nand U11270 (N_11270,N_5122,N_5325);
nand U11271 (N_11271,N_7136,N_7761);
or U11272 (N_11272,N_5164,N_7341);
nor U11273 (N_11273,N_6145,N_8972);
or U11274 (N_11274,N_9995,N_7560);
xor U11275 (N_11275,N_6050,N_6492);
or U11276 (N_11276,N_5369,N_9590);
nand U11277 (N_11277,N_8459,N_7396);
or U11278 (N_11278,N_6092,N_9559);
or U11279 (N_11279,N_5705,N_7848);
nor U11280 (N_11280,N_7678,N_6451);
or U11281 (N_11281,N_5067,N_5893);
xnor U11282 (N_11282,N_8341,N_5002);
and U11283 (N_11283,N_7555,N_8709);
or U11284 (N_11284,N_8606,N_8977);
xor U11285 (N_11285,N_6790,N_5311);
nand U11286 (N_11286,N_8770,N_5726);
nand U11287 (N_11287,N_9269,N_5727);
and U11288 (N_11288,N_7398,N_5339);
nand U11289 (N_11289,N_8994,N_8491);
or U11290 (N_11290,N_8401,N_6481);
or U11291 (N_11291,N_8467,N_6403);
and U11292 (N_11292,N_9624,N_9783);
nand U11293 (N_11293,N_9872,N_5213);
nor U11294 (N_11294,N_8022,N_7863);
nor U11295 (N_11295,N_8941,N_8415);
or U11296 (N_11296,N_6521,N_6176);
nand U11297 (N_11297,N_5729,N_6364);
nand U11298 (N_11298,N_5496,N_9931);
nor U11299 (N_11299,N_8545,N_9500);
xnor U11300 (N_11300,N_9099,N_6973);
nor U11301 (N_11301,N_7450,N_7599);
nor U11302 (N_11302,N_7494,N_7790);
nand U11303 (N_11303,N_5051,N_9631);
nand U11304 (N_11304,N_8405,N_5596);
or U11305 (N_11305,N_5507,N_5334);
xor U11306 (N_11306,N_7797,N_7315);
nand U11307 (N_11307,N_9293,N_8797);
nor U11308 (N_11308,N_9188,N_9443);
nand U11309 (N_11309,N_5406,N_9820);
xor U11310 (N_11310,N_5670,N_6046);
nand U11311 (N_11311,N_7373,N_8122);
and U11312 (N_11312,N_6057,N_5915);
nand U11313 (N_11313,N_8587,N_6691);
nor U11314 (N_11314,N_8100,N_7167);
nand U11315 (N_11315,N_8353,N_6124);
nand U11316 (N_11316,N_9944,N_5062);
or U11317 (N_11317,N_8119,N_8153);
nand U11318 (N_11318,N_6941,N_6713);
xnor U11319 (N_11319,N_7041,N_9139);
and U11320 (N_11320,N_8136,N_7211);
nand U11321 (N_11321,N_6768,N_6266);
and U11322 (N_11322,N_6091,N_6780);
nand U11323 (N_11323,N_5900,N_7571);
and U11324 (N_11324,N_5021,N_9236);
nand U11325 (N_11325,N_7783,N_5132);
and U11326 (N_11326,N_7645,N_5564);
or U11327 (N_11327,N_9232,N_6249);
or U11328 (N_11328,N_9133,N_5922);
nor U11329 (N_11329,N_9274,N_9092);
xor U11330 (N_11330,N_8743,N_8450);
nand U11331 (N_11331,N_6928,N_6936);
and U11332 (N_11332,N_7067,N_5536);
or U11333 (N_11333,N_9308,N_7670);
nor U11334 (N_11334,N_7926,N_7050);
or U11335 (N_11335,N_6603,N_9635);
nor U11336 (N_11336,N_8989,N_6883);
xnor U11337 (N_11337,N_9992,N_9659);
and U11338 (N_11338,N_7712,N_6975);
xnor U11339 (N_11339,N_7521,N_5869);
or U11340 (N_11340,N_8169,N_9212);
or U11341 (N_11341,N_6352,N_9523);
xor U11342 (N_11342,N_7796,N_8265);
or U11343 (N_11343,N_5639,N_9336);
xor U11344 (N_11344,N_5181,N_7300);
nor U11345 (N_11345,N_7150,N_5202);
nand U11346 (N_11346,N_9150,N_5674);
nor U11347 (N_11347,N_5610,N_5935);
or U11348 (N_11348,N_6599,N_6472);
or U11349 (N_11349,N_8656,N_5730);
nor U11350 (N_11350,N_9937,N_7775);
and U11351 (N_11351,N_8750,N_9197);
nand U11352 (N_11352,N_5983,N_8692);
and U11353 (N_11353,N_7156,N_5728);
nand U11354 (N_11354,N_9984,N_9793);
and U11355 (N_11355,N_6671,N_7861);
nand U11356 (N_11356,N_9343,N_5620);
xor U11357 (N_11357,N_6262,N_5679);
and U11358 (N_11358,N_9454,N_5654);
nand U11359 (N_11359,N_7589,N_5160);
xnor U11360 (N_11360,N_6333,N_7127);
or U11361 (N_11361,N_6643,N_8292);
and U11362 (N_11362,N_9569,N_5889);
xnor U11363 (N_11363,N_7265,N_5187);
xor U11364 (N_11364,N_5798,N_6760);
nand U11365 (N_11365,N_6584,N_7764);
and U11366 (N_11366,N_5997,N_8044);
and U11367 (N_11367,N_5848,N_9339);
and U11368 (N_11368,N_6589,N_8239);
nand U11369 (N_11369,N_5077,N_6709);
xor U11370 (N_11370,N_9578,N_5560);
nor U11371 (N_11371,N_6359,N_8664);
xnor U11372 (N_11372,N_8604,N_7538);
xnor U11373 (N_11373,N_7629,N_8567);
nand U11374 (N_11374,N_5923,N_7104);
nand U11375 (N_11375,N_9737,N_5976);
nand U11376 (N_11376,N_5092,N_8296);
nand U11377 (N_11377,N_7432,N_7027);
or U11378 (N_11378,N_9004,N_9289);
nand U11379 (N_11379,N_7249,N_7369);
nand U11380 (N_11380,N_9121,N_6154);
or U11381 (N_11381,N_6740,N_8553);
and U11382 (N_11382,N_6899,N_9567);
and U11383 (N_11383,N_5489,N_6887);
and U11384 (N_11384,N_6142,N_7049);
nand U11385 (N_11385,N_5819,N_6275);
or U11386 (N_11386,N_5282,N_6816);
or U11387 (N_11387,N_6094,N_5604);
nor U11388 (N_11388,N_6355,N_6540);
nor U11389 (N_11389,N_6783,N_7317);
nor U11390 (N_11390,N_5417,N_8721);
xnor U11391 (N_11391,N_5865,N_8503);
nor U11392 (N_11392,N_8991,N_7239);
nor U11393 (N_11393,N_8146,N_7655);
nand U11394 (N_11394,N_6982,N_8310);
and U11395 (N_11395,N_8701,N_7151);
nand U11396 (N_11396,N_7048,N_9751);
nand U11397 (N_11397,N_5541,N_5653);
and U11398 (N_11398,N_5549,N_5366);
and U11399 (N_11399,N_7847,N_9638);
or U11400 (N_11400,N_8366,N_8494);
xnor U11401 (N_11401,N_7217,N_8955);
and U11402 (N_11402,N_7852,N_6897);
xor U11403 (N_11403,N_7727,N_8773);
and U11404 (N_11404,N_8931,N_7610);
and U11405 (N_11405,N_6814,N_9303);
or U11406 (N_11406,N_6365,N_8521);
or U11407 (N_11407,N_7108,N_7898);
and U11408 (N_11408,N_8965,N_9395);
and U11409 (N_11409,N_6586,N_7473);
or U11410 (N_11410,N_9909,N_5205);
or U11411 (N_11411,N_5247,N_5478);
xor U11412 (N_11412,N_7646,N_9623);
and U11413 (N_11413,N_6600,N_8933);
xnor U11414 (N_11414,N_7881,N_7738);
and U11415 (N_11415,N_9933,N_9221);
xor U11416 (N_11416,N_8190,N_7033);
and U11417 (N_11417,N_5429,N_7038);
nand U11418 (N_11418,N_5057,N_8899);
and U11419 (N_11419,N_7040,N_6831);
xnor U11420 (N_11420,N_8575,N_9301);
nand U11421 (N_11421,N_8563,N_8062);
nand U11422 (N_11422,N_9389,N_7746);
and U11423 (N_11423,N_8547,N_9797);
xor U11424 (N_11424,N_9017,N_9976);
and U11425 (N_11425,N_8484,N_5625);
xnor U11426 (N_11426,N_8669,N_9724);
nor U11427 (N_11427,N_7613,N_9547);
xor U11428 (N_11428,N_6325,N_5982);
nor U11429 (N_11429,N_9428,N_6912);
nor U11430 (N_11430,N_6656,N_7643);
nor U11431 (N_11431,N_5487,N_6348);
and U11432 (N_11432,N_7469,N_9854);
or U11433 (N_11433,N_6166,N_8850);
or U11434 (N_11434,N_9422,N_8377);
nor U11435 (N_11435,N_7005,N_8294);
and U11436 (N_11436,N_9502,N_8565);
xnor U11437 (N_11437,N_7871,N_9591);
and U11438 (N_11438,N_5456,N_6776);
nand U11439 (N_11439,N_7246,N_5147);
nor U11440 (N_11440,N_7730,N_5908);
and U11441 (N_11441,N_8118,N_7981);
or U11442 (N_11442,N_5373,N_6507);
xnor U11443 (N_11443,N_7179,N_8103);
xor U11444 (N_11444,N_9946,N_8533);
xnor U11445 (N_11445,N_7858,N_6404);
nor U11446 (N_11446,N_8829,N_8889);
nand U11447 (N_11447,N_8202,N_5897);
nor U11448 (N_11448,N_8408,N_6164);
nand U11449 (N_11449,N_7906,N_6127);
nor U11450 (N_11450,N_5313,N_9340);
nand U11451 (N_11451,N_6216,N_5782);
nand U11452 (N_11452,N_5832,N_6826);
and U11453 (N_11453,N_6822,N_6112);
or U11454 (N_11454,N_7197,N_9000);
or U11455 (N_11455,N_7483,N_9532);
nand U11456 (N_11456,N_6456,N_6185);
nor U11457 (N_11457,N_8502,N_9541);
nor U11458 (N_11458,N_7570,N_7056);
or U11459 (N_11459,N_5251,N_6801);
or U11460 (N_11460,N_7427,N_6022);
and U11461 (N_11461,N_8534,N_8694);
or U11462 (N_11462,N_6004,N_5630);
nor U11463 (N_11463,N_9455,N_9431);
or U11464 (N_11464,N_6564,N_9858);
nor U11465 (N_11465,N_5134,N_7366);
nor U11466 (N_11466,N_8848,N_8734);
xor U11467 (N_11467,N_5614,N_9663);
xnor U11468 (N_11468,N_6269,N_5410);
and U11469 (N_11469,N_6104,N_7856);
xnor U11470 (N_11470,N_9444,N_7088);
nor U11471 (N_11471,N_9577,N_7841);
or U11472 (N_11472,N_6469,N_8457);
or U11473 (N_11473,N_8375,N_5444);
or U11474 (N_11474,N_7891,N_9977);
and U11475 (N_11475,N_8107,N_8330);
or U11476 (N_11476,N_9094,N_8322);
nor U11477 (N_11477,N_9448,N_9190);
or U11478 (N_11478,N_7747,N_8703);
or U11479 (N_11479,N_8623,N_9282);
nor U11480 (N_11480,N_7140,N_5453);
nor U11481 (N_11481,N_6259,N_6800);
and U11482 (N_11482,N_8763,N_9045);
nor U11483 (N_11483,N_6758,N_9708);
and U11484 (N_11484,N_6390,N_5335);
nand U11485 (N_11485,N_8133,N_6557);
xor U11486 (N_11486,N_5810,N_8526);
nand U11487 (N_11487,N_5542,N_5754);
and U11488 (N_11488,N_5599,N_7716);
and U11489 (N_11489,N_8681,N_8905);
and U11490 (N_11490,N_5372,N_9902);
nor U11491 (N_11491,N_8990,N_5968);
nand U11492 (N_11492,N_9227,N_5852);
nor U11493 (N_11493,N_6475,N_6499);
xor U11494 (N_11494,N_6027,N_6716);
and U11495 (N_11495,N_6219,N_8424);
xor U11496 (N_11496,N_8048,N_9867);
xor U11497 (N_11497,N_8861,N_6156);
or U11498 (N_11498,N_8527,N_8237);
nor U11499 (N_11499,N_5914,N_6065);
or U11500 (N_11500,N_5232,N_7429);
nand U11501 (N_11501,N_5314,N_5656);
nand U11502 (N_11502,N_5616,N_6793);
or U11503 (N_11503,N_8583,N_6125);
or U11504 (N_11504,N_6728,N_6428);
nor U11505 (N_11505,N_7983,N_9868);
or U11506 (N_11506,N_9122,N_6088);
xor U11507 (N_11507,N_7210,N_8875);
or U11508 (N_11508,N_7380,N_5880);
or U11509 (N_11509,N_6470,N_7578);
xor U11510 (N_11510,N_7159,N_7184);
nand U11511 (N_11511,N_6076,N_6272);
and U11512 (N_11512,N_7377,N_8945);
nor U11513 (N_11513,N_5348,N_9916);
and U11514 (N_11514,N_7175,N_5768);
and U11515 (N_11515,N_9899,N_8711);
and U11516 (N_11516,N_7226,N_7287);
xnor U11517 (N_11517,N_5579,N_7293);
xnor U11518 (N_11518,N_8707,N_7961);
or U11519 (N_11519,N_5672,N_5554);
or U11520 (N_11520,N_6442,N_6662);
nor U11521 (N_11521,N_6160,N_7060);
xnor U11522 (N_11522,N_7820,N_6440);
and U11523 (N_11523,N_8914,N_6796);
xnor U11524 (N_11524,N_8752,N_6833);
nor U11525 (N_11525,N_5584,N_7933);
nand U11526 (N_11526,N_5178,N_8495);
xnor U11527 (N_11527,N_7922,N_5431);
or U11528 (N_11528,N_8828,N_9043);
and U11529 (N_11529,N_6538,N_7915);
or U11530 (N_11530,N_9485,N_8677);
nand U11531 (N_11531,N_9686,N_6676);
nor U11532 (N_11532,N_6620,N_6446);
or U11533 (N_11533,N_6360,N_5794);
nand U11534 (N_11534,N_8629,N_8183);
xor U11535 (N_11535,N_7787,N_7449);
nor U11536 (N_11536,N_8309,N_5012);
nor U11537 (N_11537,N_9706,N_9918);
nor U11538 (N_11538,N_7532,N_7851);
nor U11539 (N_11539,N_5148,N_7080);
nand U11540 (N_11540,N_8343,N_9808);
nand U11541 (N_11541,N_9193,N_7969);
and U11542 (N_11542,N_8929,N_7006);
xnor U11543 (N_11543,N_5128,N_8626);
or U11544 (N_11544,N_7973,N_7559);
nor U11545 (N_11545,N_6988,N_6396);
nand U11546 (N_11546,N_9840,N_6991);
nor U11547 (N_11547,N_9556,N_6257);
nor U11548 (N_11548,N_7531,N_7503);
xnor U11549 (N_11549,N_7666,N_6979);
xnor U11550 (N_11550,N_9528,N_8951);
xor U11551 (N_11551,N_8205,N_6919);
and U11552 (N_11552,N_6055,N_6850);
or U11553 (N_11553,N_8072,N_7631);
or U11554 (N_11554,N_9334,N_7492);
nand U11555 (N_11555,N_7292,N_8884);
nand U11556 (N_11556,N_6841,N_5700);
nand U11557 (N_11557,N_6422,N_6942);
or U11558 (N_11558,N_7663,N_6721);
nor U11559 (N_11559,N_6037,N_8052);
and U11560 (N_11560,N_5644,N_8756);
or U11561 (N_11561,N_8086,N_7114);
xnor U11562 (N_11562,N_5288,N_5785);
nor U11563 (N_11563,N_5031,N_8695);
xor U11564 (N_11564,N_6075,N_8298);
or U11565 (N_11565,N_5378,N_8416);
or U11566 (N_11566,N_9331,N_8047);
xor U11567 (N_11567,N_7412,N_6929);
and U11568 (N_11568,N_6367,N_6623);
and U11569 (N_11569,N_5392,N_9167);
xnor U11570 (N_11570,N_7077,N_9276);
nor U11571 (N_11571,N_5452,N_5510);
and U11572 (N_11572,N_8188,N_8780);
or U11573 (N_11573,N_7997,N_9968);
and U11574 (N_11574,N_8954,N_9608);
nor U11575 (N_11575,N_8442,N_5993);
or U11576 (N_11576,N_6932,N_8498);
nand U11577 (N_11577,N_5776,N_6518);
xor U11578 (N_11578,N_9707,N_7529);
nor U11579 (N_11579,N_8935,N_9463);
nand U11580 (N_11580,N_6864,N_5210);
nand U11581 (N_11581,N_8646,N_7443);
nor U11582 (N_11582,N_9844,N_6647);
nand U11583 (N_11583,N_7258,N_5973);
or U11584 (N_11584,N_8251,N_5204);
and U11585 (N_11585,N_6955,N_6891);
nor U11586 (N_11586,N_7497,N_5777);
nor U11587 (N_11587,N_7271,N_6327);
and U11588 (N_11588,N_6918,N_7405);
xor U11589 (N_11589,N_8006,N_7650);
or U11590 (N_11590,N_9225,N_6090);
nor U11591 (N_11591,N_9159,N_7675);
nand U11592 (N_11592,N_5995,N_6708);
xor U11593 (N_11593,N_8289,N_6574);
nor U11594 (N_11594,N_5461,N_8039);
and U11595 (N_11595,N_6175,N_7083);
nand U11596 (N_11596,N_8141,N_5948);
xor U11597 (N_11597,N_9675,N_8194);
or U11598 (N_11598,N_7219,N_7448);
nor U11599 (N_11599,N_7107,N_8821);
nor U11600 (N_11600,N_6083,N_7759);
or U11601 (N_11601,N_7536,N_6071);
nand U11602 (N_11602,N_5888,N_5457);
or U11603 (N_11603,N_7417,N_8786);
nor U11604 (N_11604,N_6059,N_7283);
xor U11605 (N_11605,N_5353,N_9251);
and U11606 (N_11606,N_9905,N_7288);
and U11607 (N_11607,N_9842,N_5632);
nand U11608 (N_11608,N_6717,N_6913);
nor U11609 (N_11609,N_8117,N_6560);
nor U11610 (N_11610,N_8649,N_8888);
xnor U11611 (N_11611,N_7883,N_5340);
nand U11612 (N_11612,N_5041,N_6074);
or U11613 (N_11613,N_6459,N_9886);
nor U11614 (N_11614,N_5124,N_6994);
nand U11615 (N_11615,N_9315,N_8874);
nor U11616 (N_11616,N_6500,N_5413);
and U11617 (N_11617,N_8030,N_9478);
nor U11618 (N_11618,N_9208,N_7625);
or U11619 (N_11619,N_8683,N_8844);
xnor U11620 (N_11620,N_6349,N_8574);
nor U11621 (N_11621,N_8960,N_6700);
and U11622 (N_11622,N_6043,N_9394);
xor U11623 (N_11623,N_8636,N_8761);
xor U11624 (N_11624,N_9753,N_7514);
or U11625 (N_11625,N_7014,N_5040);
xor U11626 (N_11626,N_5032,N_7864);
xor U11627 (N_11627,N_6060,N_5310);
and U11628 (N_11628,N_6278,N_7690);
or U11629 (N_11629,N_9655,N_6818);
and U11630 (N_11630,N_9204,N_5418);
nor U11631 (N_11631,N_6462,N_6659);
or U11632 (N_11632,N_8060,N_8742);
xnor U11633 (N_11633,N_5017,N_5698);
xor U11634 (N_11634,N_7408,N_9104);
or U11635 (N_11635,N_7633,N_8536);
and U11636 (N_11636,N_7139,N_7032);
and U11637 (N_11637,N_6025,N_9563);
nor U11638 (N_11638,N_8151,N_6047);
xnor U11639 (N_11639,N_8896,N_9917);
and U11640 (N_11640,N_6316,N_5201);
nor U11641 (N_11641,N_8161,N_6840);
and U11642 (N_11642,N_6226,N_9291);
or U11643 (N_11643,N_5131,N_8477);
or U11644 (N_11644,N_8128,N_7762);
and U11645 (N_11645,N_8854,N_5821);
and U11646 (N_11646,N_9670,N_9754);
nor U11647 (N_11647,N_6890,N_6807);
and U11648 (N_11648,N_8645,N_6468);
and U11649 (N_11649,N_8249,N_8643);
or U11650 (N_11650,N_8907,N_8822);
nor U11651 (N_11651,N_7984,N_6128);
and U11652 (N_11652,N_5755,N_8705);
xnor U11653 (N_11653,N_9086,N_6614);
nor U11654 (N_11654,N_9506,N_6704);
nor U11655 (N_11655,N_7205,N_8064);
xnor U11656 (N_11656,N_8880,N_9279);
xor U11657 (N_11657,N_9587,N_9381);
nor U11658 (N_11658,N_7544,N_7141);
nor U11659 (N_11659,N_8170,N_5681);
nand U11660 (N_11660,N_7737,N_7653);
or U11661 (N_11661,N_5216,N_5540);
nand U11662 (N_11662,N_9583,N_6992);
or U11663 (N_11663,N_5100,N_9217);
and U11664 (N_11664,N_6320,N_8154);
and U11665 (N_11665,N_7868,N_5624);
or U11666 (N_11666,N_6712,N_9273);
nor U11667 (N_11667,N_5230,N_7166);
xor U11668 (N_11668,N_6161,N_8859);
nor U11669 (N_11669,N_7280,N_5331);
nor U11670 (N_11670,N_7340,N_9354);
nor U11671 (N_11671,N_9928,N_5714);
or U11672 (N_11672,N_8404,N_5048);
nand U11673 (N_11673,N_9945,N_6830);
or U11674 (N_11674,N_6436,N_9950);
nor U11675 (N_11675,N_8272,N_8092);
and U11676 (N_11676,N_8423,N_9741);
nand U11677 (N_11677,N_6008,N_7740);
nand U11678 (N_11678,N_9046,N_6181);
or U11679 (N_11679,N_9419,N_7294);
xor U11680 (N_11680,N_9185,N_5701);
or U11681 (N_11681,N_7723,N_7418);
and U11682 (N_11682,N_9415,N_7214);
xnor U11683 (N_11683,N_5715,N_5312);
and U11684 (N_11684,N_5129,N_5992);
or U11685 (N_11685,N_8195,N_7154);
nand U11686 (N_11686,N_9714,N_9610);
and U11687 (N_11687,N_8303,N_8558);
and U11688 (N_11688,N_7626,N_8225);
xor U11689 (N_11689,N_7634,N_9900);
nand U11690 (N_11690,N_8644,N_8390);
and U11691 (N_11691,N_6522,N_5498);
and U11692 (N_11692,N_7074,N_9117);
and U11693 (N_11693,N_6519,N_6957);
and U11694 (N_11694,N_8336,N_7296);
nand U11695 (N_11695,N_8501,N_6162);
nor U11696 (N_11696,N_9189,N_7720);
nand U11697 (N_11697,N_5345,N_5543);
nor U11698 (N_11698,N_9709,N_5965);
nand U11699 (N_11699,N_9260,N_6585);
nand U11700 (N_11700,N_5966,N_5098);
nor U11701 (N_11701,N_9392,N_8361);
xor U11702 (N_11702,N_7191,N_8177);
or U11703 (N_11703,N_9890,N_8212);
nor U11704 (N_11704,N_8619,N_7819);
nor U11705 (N_11705,N_6993,N_6861);
xnor U11706 (N_11706,N_7003,N_9370);
and U11707 (N_11707,N_7692,N_5867);
and U11708 (N_11708,N_5562,N_9271);
nand U11709 (N_11709,N_8794,N_8185);
nand U11710 (N_11710,N_7467,N_9573);
xor U11711 (N_11711,N_8297,N_5261);
nand U11712 (N_11712,N_9347,N_9414);
and U11713 (N_11713,N_7034,N_5521);
and U11714 (N_11714,N_5432,N_9765);
nor U11715 (N_11715,N_7365,N_6329);
and U11716 (N_11716,N_5856,N_5088);
or U11717 (N_11717,N_5812,N_6524);
or U11718 (N_11718,N_9620,N_5928);
nand U11719 (N_11719,N_7667,N_9085);
and U11720 (N_11720,N_9943,N_5626);
and U11721 (N_11721,N_7575,N_9105);
nor U11722 (N_11722,N_5879,N_9924);
or U11723 (N_11723,N_6171,N_8956);
nor U11724 (N_11724,N_5974,N_9880);
or U11725 (N_11725,N_9712,N_6718);
xor U11726 (N_11726,N_7213,N_6598);
nand U11727 (N_11727,N_8430,N_7480);
xnor U11728 (N_11728,N_8114,N_9229);
or U11729 (N_11729,N_8008,N_5878);
or U11730 (N_11730,N_5385,N_5547);
nand U11731 (N_11731,N_9299,N_8250);
and U11732 (N_11732,N_7943,N_6596);
xor U11733 (N_11733,N_6031,N_5567);
nand U11734 (N_11734,N_9350,N_6084);
nand U11735 (N_11735,N_8230,N_7818);
nand U11736 (N_11736,N_7854,N_9951);
nor U11737 (N_11737,N_5371,N_9742);
xor U11738 (N_11738,N_6888,N_7247);
or U11739 (N_11739,N_7295,N_5682);
and U11740 (N_11740,N_7190,N_7632);
or U11741 (N_11741,N_7264,N_7709);
or U11742 (N_11742,N_5838,N_9926);
xor U11743 (N_11743,N_6681,N_6069);
or U11744 (N_11744,N_7654,N_6950);
and U11745 (N_11745,N_8535,N_5837);
nand U11746 (N_11746,N_9966,N_7837);
xnor U11747 (N_11747,N_7234,N_5703);
nor U11748 (N_11748,N_6779,N_9514);
and U11749 (N_11749,N_5859,N_8428);
xnor U11750 (N_11750,N_7921,N_6005);
or U11751 (N_11751,N_8564,N_5118);
and U11752 (N_11752,N_6238,N_8277);
xor U11753 (N_11753,N_7121,N_8397);
nor U11754 (N_11754,N_6400,N_6917);
or U11755 (N_11755,N_8445,N_6338);
and U11756 (N_11756,N_8598,N_8670);
or U11757 (N_11757,N_6515,N_5512);
or U11758 (N_11758,N_9497,N_6030);
nor U11759 (N_11759,N_8973,N_6781);
or U11760 (N_11760,N_5555,N_7886);
nor U11761 (N_11761,N_8708,N_6959);
xnor U11762 (N_11762,N_8339,N_9295);
and U11763 (N_11763,N_5265,N_9652);
and U11764 (N_11764,N_9756,N_5751);
and U11765 (N_11765,N_5645,N_9582);
nand U11766 (N_11766,N_7669,N_5530);
nor U11767 (N_11767,N_8713,N_9894);
nor U11768 (N_11768,N_7800,N_5606);
nand U11769 (N_11769,N_5901,N_5015);
nand U11770 (N_11770,N_5786,N_5255);
xnor U11771 (N_11771,N_8893,N_7642);
nor U11772 (N_11772,N_5695,N_7561);
nand U11773 (N_11773,N_7604,N_9253);
xnor U11774 (N_11774,N_6576,N_8432);
xnor U11775 (N_11775,N_7209,N_8054);
and U11776 (N_11776,N_9614,N_6398);
or U11777 (N_11777,N_7445,N_8596);
nand U11778 (N_11778,N_5168,N_7236);
nor U11779 (N_11779,N_5152,N_9694);
xnor U11780 (N_11780,N_9904,N_7355);
nor U11781 (N_11781,N_6256,N_9090);
or U11782 (N_11782,N_8323,N_7562);
and U11783 (N_11783,N_6675,N_5248);
nand U11784 (N_11784,N_8878,N_7928);
xor U11785 (N_11785,N_5994,N_5233);
nor U11786 (N_11786,N_6170,N_6504);
nor U11787 (N_11787,N_8637,N_7007);
or U11788 (N_11788,N_5860,N_5449);
nor U11789 (N_11789,N_5252,N_7351);
and U11790 (N_11790,N_9462,N_9986);
nand U11791 (N_11791,N_8448,N_7664);
xnor U11792 (N_11792,N_6725,N_7299);
nand U11793 (N_11793,N_5740,N_7385);
nand U11794 (N_11794,N_7089,N_7649);
and U11795 (N_11795,N_9359,N_8675);
and U11796 (N_11796,N_8947,N_7993);
xnor U11797 (N_11797,N_5962,N_7768);
and U11798 (N_11798,N_9215,N_8367);
nor U11799 (N_11799,N_9416,N_6849);
nand U11800 (N_11800,N_6430,N_7733);
nand U11801 (N_11801,N_9782,N_5975);
xnor U11802 (N_11802,N_9182,N_8281);
xor U11803 (N_11803,N_6117,N_5420);
nand U11804 (N_11804,N_7328,N_9198);
xor U11805 (N_11805,N_5788,N_9606);
nor U11806 (N_11806,N_8033,N_5532);
or U11807 (N_11807,N_5642,N_5550);
and U11808 (N_11808,N_5911,N_9228);
xnor U11809 (N_11809,N_8815,N_7368);
and U11810 (N_11810,N_7586,N_7137);
and U11811 (N_11811,N_7230,N_6969);
or U11812 (N_11812,N_6755,N_8173);
xor U11813 (N_11813,N_8571,N_8904);
or U11814 (N_11814,N_6265,N_5999);
and U11815 (N_11815,N_5710,N_6884);
and U11816 (N_11816,N_9102,N_8045);
xnor U11817 (N_11817,N_9116,N_6746);
or U11818 (N_11818,N_6751,N_5660);
nand U11819 (N_11819,N_5053,N_5272);
xnor U11820 (N_11820,N_8422,N_7022);
nand U11821 (N_11821,N_8732,N_6495);
nor U11822 (N_11822,N_7966,N_5435);
nand U11823 (N_11823,N_7587,N_9097);
and U11824 (N_11824,N_5803,N_6748);
xnor U11825 (N_11825,N_8085,N_9360);
and U11826 (N_11826,N_8013,N_9626);
or U11827 (N_11827,N_7478,N_5591);
nor U11828 (N_11828,N_7786,N_6866);
nand U11829 (N_11829,N_9391,N_5484);
nand U11830 (N_11830,N_9216,N_6411);
nand U11831 (N_11831,N_5028,N_6556);
or U11832 (N_11832,N_9884,N_7533);
nor U11833 (N_11833,N_6299,N_9702);
nand U11834 (N_11834,N_5304,N_8903);
nand U11835 (N_11835,N_6229,N_5136);
nand U11836 (N_11836,N_7306,N_6130);
nand U11837 (N_11837,N_6680,N_8667);
nand U11838 (N_11838,N_5905,N_8490);
xor U11839 (N_11839,N_5083,N_8799);
xnor U11840 (N_11840,N_9224,N_8747);
or U11841 (N_11841,N_9456,N_6633);
nor U11842 (N_11842,N_9095,N_7382);
and U11843 (N_11843,N_8624,N_5184);
nor U11844 (N_11844,N_6821,N_5079);
or U11845 (N_11845,N_5638,N_9667);
xor U11846 (N_11846,N_6719,N_5524);
nor U11847 (N_11847,N_7976,N_6419);
and U11848 (N_11848,N_9364,N_9766);
xor U11849 (N_11849,N_5662,N_5145);
or U11850 (N_11850,N_6397,N_9690);
and U11851 (N_11851,N_6949,N_5641);
or U11852 (N_11852,N_9630,N_9153);
nor U11853 (N_11853,N_7402,N_6426);
nand U11854 (N_11854,N_6931,N_6619);
xor U11855 (N_11855,N_8157,N_8525);
or U11856 (N_11856,N_9970,N_9604);
and U11857 (N_11857,N_8196,N_7087);
xnor U11858 (N_11858,N_7782,N_5868);
and U11859 (N_11859,N_6901,N_7908);
xor U11860 (N_11860,N_8735,N_8108);
nor U11861 (N_11861,N_7735,N_6771);
and U11862 (N_11862,N_5808,N_7464);
and U11863 (N_11863,N_5246,N_6473);
or U11864 (N_11864,N_6731,N_8444);
and U11865 (N_11865,N_5892,N_8285);
or U11866 (N_11866,N_8775,N_5629);
or U11867 (N_11867,N_6673,N_8650);
nor U11868 (N_11868,N_9612,N_7244);
and U11869 (N_11869,N_9847,N_6657);
or U11870 (N_11870,N_7202,N_6471);
nor U11871 (N_11871,N_9527,N_5592);
or U11872 (N_11872,N_8556,N_8680);
nor U11873 (N_11873,N_9927,N_5173);
xnor U11874 (N_11874,N_6139,N_5107);
nand U11875 (N_11875,N_8539,N_5518);
xor U11876 (N_11876,N_6143,N_5691);
and U11877 (N_11877,N_7120,N_7919);
or U11878 (N_11878,N_9768,N_7446);
nor U11879 (N_11879,N_7963,N_5066);
nor U11880 (N_11880,N_5666,N_6604);
and U11881 (N_11881,N_9068,N_6204);
and U11882 (N_11882,N_5135,N_7273);
and U11883 (N_11883,N_7907,N_9656);
or U11884 (N_11884,N_9120,N_7924);
or U11885 (N_11885,N_5419,N_8411);
nand U11886 (N_11886,N_5407,N_6869);
nor U11887 (N_11887,N_6421,N_6632);
and U11888 (N_11888,N_9882,N_9014);
and U11889 (N_11889,N_5668,N_8074);
or U11890 (N_11890,N_7989,N_9498);
and U11891 (N_11891,N_7125,N_5677);
xor U11892 (N_11892,N_9727,N_9311);
nand U11893 (N_11893,N_6625,N_9356);
or U11894 (N_11894,N_7867,N_8226);
nand U11895 (N_11895,N_8076,N_6350);
nor U11896 (N_11896,N_5111,N_9994);
or U11897 (N_11897,N_8053,N_6287);
nor U11898 (N_11898,N_7488,N_7326);
xnor U11899 (N_11899,N_9544,N_7731);
nand U11900 (N_11900,N_7605,N_6654);
and U11901 (N_11901,N_6798,N_8012);
and U11902 (N_11902,N_6697,N_9862);
nand U11903 (N_11903,N_8655,N_8028);
or U11904 (N_11904,N_9982,N_8280);
xnor U11905 (N_11905,N_8569,N_8971);
or U11906 (N_11906,N_5750,N_6189);
xor U11907 (N_11907,N_7376,N_7333);
and U11908 (N_11908,N_8716,N_9348);
nor U11909 (N_11909,N_6765,N_8215);
nor U11910 (N_11910,N_6429,N_6677);
or U11911 (N_11911,N_7000,N_5764);
nor U11912 (N_11912,N_8469,N_8246);
or U11913 (N_11913,N_9417,N_6577);
and U11914 (N_11914,N_8740,N_8392);
xor U11915 (N_11915,N_5613,N_6028);
xor U11916 (N_11916,N_9517,N_7714);
nor U11917 (N_11917,N_6330,N_5493);
nand U11918 (N_11918,N_7053,N_7207);
xor U11919 (N_11919,N_8399,N_5989);
xnor U11920 (N_11920,N_8864,N_5844);
nor U11921 (N_11921,N_9770,N_9259);
xor U11922 (N_11922,N_9693,N_5425);
or U11923 (N_11923,N_5003,N_5517);
xnor U11924 (N_11924,N_6341,N_8659);
xor U11925 (N_11925,N_5585,N_5045);
or U11926 (N_11926,N_7100,N_8748);
nand U11927 (N_11927,N_7551,N_6212);
nor U11928 (N_11928,N_7318,N_9361);
nor U11929 (N_11929,N_7472,N_8640);
xor U11930 (N_11930,N_6706,N_7109);
and U11931 (N_11931,N_5600,N_6963);
nor U11932 (N_11932,N_9051,N_6493);
or U11933 (N_11933,N_7592,N_7062);
xnor U11934 (N_11934,N_6649,N_8492);
or U11935 (N_11935,N_8419,N_9231);
or U11936 (N_11936,N_5822,N_7342);
or U11937 (N_11937,N_6872,N_9747);
and U11938 (N_11938,N_8959,N_7176);
nand U11939 (N_11939,N_6839,N_8682);
xnor U11940 (N_11940,N_7539,N_5544);
xnor U11941 (N_11941,N_5943,N_8334);
and U11942 (N_11942,N_7353,N_6615);
nor U11943 (N_11943,N_8595,N_6179);
nand U11944 (N_11944,N_7066,N_7916);
and U11945 (N_11945,N_5207,N_9925);
and U11946 (N_11946,N_7344,N_7791);
xor U11947 (N_11947,N_7853,N_7362);
nand U11948 (N_11948,N_8040,N_5617);
nor U11949 (N_11949,N_7665,N_6377);
or U11950 (N_11950,N_6894,N_9040);
or U11951 (N_11951,N_9981,N_9434);
nor U11952 (N_11952,N_5891,N_6113);
or U11953 (N_11953,N_8088,N_7103);
xor U11954 (N_11954,N_7367,N_8548);
nor U11955 (N_11955,N_8027,N_9091);
xnor U11956 (N_11956,N_5427,N_7703);
nor U11957 (N_11957,N_5582,N_6220);
or U11958 (N_11958,N_9080,N_5043);
nor U11959 (N_11959,N_5235,N_6502);
nor U11960 (N_11960,N_8823,N_8344);
or U11961 (N_11961,N_6533,N_9306);
nand U11962 (N_11962,N_5001,N_5381);
or U11963 (N_11963,N_7579,N_7722);
and U11964 (N_11964,N_8978,N_7888);
nand U11965 (N_11965,N_5215,N_9304);
or U11966 (N_11966,N_9078,N_7024);
and U11967 (N_11967,N_6296,N_9035);
or U11968 (N_11968,N_8837,N_8449);
or U11969 (N_11969,N_8696,N_9241);
nand U11970 (N_11970,N_7358,N_6520);
nor U11971 (N_11971,N_6842,N_6739);
nor U11972 (N_11972,N_6371,N_8263);
or U11973 (N_11973,N_9073,N_7860);
nor U11974 (N_11974,N_9861,N_6693);
nand U11975 (N_11975,N_6336,N_7801);
nor U11976 (N_11976,N_9850,N_6999);
xor U11977 (N_11977,N_5108,N_7155);
or U11978 (N_11978,N_6077,N_7875);
xnor U11979 (N_11979,N_5127,N_8932);
xnor U11980 (N_11980,N_7428,N_8115);
xnor U11981 (N_11981,N_7811,N_9374);
or U11982 (N_11982,N_9595,N_8164);
or U11983 (N_11983,N_7031,N_8826);
xnor U11984 (N_11984,N_7479,N_5227);
or U11985 (N_11985,N_6858,N_5455);
or U11986 (N_11986,N_9258,N_9816);
or U11987 (N_11987,N_5631,N_7260);
xnor U11988 (N_11988,N_7384,N_8560);
nor U11989 (N_11989,N_7752,N_6196);
nand U11990 (N_11990,N_6303,N_9351);
or U11991 (N_11991,N_5474,N_5401);
nand U11992 (N_11992,N_9213,N_6089);
and U11993 (N_11993,N_8728,N_5475);
and U11994 (N_11994,N_7325,N_7276);
or U11995 (N_11995,N_7849,N_8043);
nand U11996 (N_11996,N_6565,N_6660);
nor U11997 (N_11997,N_7597,N_5004);
and U11998 (N_11998,N_7187,N_5731);
and U11999 (N_11999,N_7267,N_7012);
or U12000 (N_12000,N_5356,N_8055);
xnor U12001 (N_12001,N_5211,N_8087);
xor U12002 (N_12002,N_8562,N_7158);
nor U12003 (N_12003,N_9642,N_5018);
xnor U12004 (N_12004,N_6410,N_6402);
or U12005 (N_12005,N_7936,N_5322);
xor U12006 (N_12006,N_5179,N_9835);
and U12007 (N_12007,N_7729,N_7036);
xor U12008 (N_12008,N_9404,N_8091);
or U12009 (N_12009,N_9346,N_6921);
nand U12010 (N_12010,N_9412,N_8612);
xor U12011 (N_12011,N_7781,N_7766);
nor U12012 (N_12012,N_8530,N_6601);
nand U12013 (N_12013,N_8801,N_6399);
and U12014 (N_12014,N_8386,N_8793);
xor U12015 (N_12015,N_9081,N_5416);
nor U12016 (N_12016,N_6773,N_6782);
xor U12017 (N_12017,N_8846,N_9377);
nor U12018 (N_12018,N_7330,N_7436);
or U12019 (N_12019,N_6958,N_9508);
xnor U12020 (N_12020,N_6624,N_5816);
or U12021 (N_12021,N_5558,N_7713);
and U12022 (N_12022,N_9748,N_6747);
nor U12023 (N_12023,N_7704,N_5847);
nor U12024 (N_12024,N_7809,N_6231);
nand U12025 (N_12025,N_8976,N_5357);
xor U12026 (N_12026,N_5806,N_5038);
nor U12027 (N_12027,N_7042,N_9327);
and U12028 (N_12028,N_9723,N_8126);
nor U12029 (N_12029,N_6357,N_7281);
nand U12030 (N_12030,N_9828,N_7279);
nor U12031 (N_12031,N_6412,N_5580);
and U12032 (N_12032,N_6099,N_9368);
and U12033 (N_12033,N_5081,N_6353);
xor U12034 (N_12034,N_8042,N_8426);
or U12035 (N_12035,N_9796,N_8474);
nor U12036 (N_12036,N_8948,N_7116);
or U12037 (N_12037,N_8648,N_7110);
nand U12038 (N_12038,N_9338,N_8738);
nand U12039 (N_12039,N_5141,N_9234);
and U12040 (N_12040,N_5553,N_7910);
nor U12041 (N_12041,N_5315,N_5849);
nand U12042 (N_12042,N_8839,N_6618);
nand U12043 (N_12043,N_9762,N_6264);
or U12044 (N_12044,N_6655,N_7909);
and U12045 (N_12045,N_5176,N_7788);
or U12046 (N_12046,N_8555,N_8318);
xor U12047 (N_12047,N_8209,N_9380);
nor U12048 (N_12048,N_6684,N_8962);
xor U12049 (N_12049,N_8642,N_6136);
or U12050 (N_12050,N_7314,N_6634);
xnor U12051 (N_12051,N_6001,N_8260);
nor U12052 (N_12052,N_8686,N_9819);
xnor U12053 (N_12053,N_7677,N_5408);
nor U12054 (N_12054,N_9145,N_8179);
xnor U12055 (N_12055,N_9586,N_5563);
nor U12056 (N_12056,N_7789,N_9795);
xor U12057 (N_12057,N_5296,N_8568);
and U12058 (N_12058,N_7885,N_6799);
and U12059 (N_12059,N_7590,N_9967);
or U12060 (N_12060,N_6714,N_9466);
nand U12061 (N_12061,N_7549,N_5910);
or U12062 (N_12062,N_8998,N_6645);
nor U12063 (N_12063,N_5158,N_5964);
xnor U12064 (N_12064,N_5874,N_5971);
nand U12065 (N_12065,N_5684,N_8634);
xnor U12066 (N_12066,N_8316,N_8369);
or U12067 (N_12067,N_9077,N_9172);
or U12068 (N_12068,N_6622,N_8593);
nand U12069 (N_12069,N_6193,N_8590);
or U12070 (N_12070,N_7170,N_8111);
xnor U12071 (N_12071,N_8381,N_6555);
and U12072 (N_12072,N_5277,N_5843);
nand U12073 (N_12073,N_6197,N_9627);
and U12074 (N_12074,N_7390,N_9975);
xnor U12075 (N_12075,N_9138,N_5603);
nand U12076 (N_12076,N_8542,N_6241);
and U12077 (N_12077,N_7577,N_6149);
and U12078 (N_12078,N_8983,N_6011);
nor U12079 (N_12079,N_6213,N_6580);
xnor U12080 (N_12080,N_5546,N_8807);
or U12081 (N_12081,N_5857,N_7403);
xnor U12082 (N_12082,N_6882,N_9526);
xor U12083 (N_12083,N_5706,N_9908);
or U12084 (N_12084,N_6379,N_5258);
xor U12085 (N_12085,N_5885,N_6245);
or U12086 (N_12086,N_6138,N_8221);
nor U12087 (N_12087,N_7671,N_8268);
and U12088 (N_12088,N_5153,N_9711);
xnor U12089 (N_12089,N_9598,N_5463);
nand U12090 (N_12090,N_7477,N_8673);
nand U12091 (N_12091,N_9790,N_7930);
xor U12092 (N_12092,N_8123,N_8207);
nor U12093 (N_12093,N_5023,N_8857);
nand U12094 (N_12094,N_8685,N_8127);
and U12095 (N_12095,N_9715,N_8036);
and U12096 (N_12096,N_9005,N_9990);
xor U12097 (N_12097,N_7352,N_7838);
nand U12098 (N_12098,N_7685,N_8518);
nand U12099 (N_12099,N_8887,N_9100);
xor U12100 (N_12100,N_9459,N_6180);
and U12101 (N_12101,N_8982,N_6271);
nor U12102 (N_12102,N_9878,N_7261);
nand U12103 (N_12103,N_5011,N_9689);
or U12104 (N_12104,N_6756,N_7527);
nand U12105 (N_12105,N_7470,N_8800);
xor U12106 (N_12106,N_8777,N_6648);
and U12107 (N_12107,N_5707,N_6413);
and U12108 (N_12108,N_6809,N_6461);
or U12109 (N_12109,N_5116,N_7953);
or U12110 (N_12110,N_9855,N_9672);
xnor U12111 (N_12111,N_7918,N_9830);
nand U12112 (N_12112,N_7415,N_8618);
xnor U12113 (N_12113,N_8172,N_7011);
or U12114 (N_12114,N_9473,N_6893);
or U12115 (N_12115,N_6016,N_9893);
or U12116 (N_12116,N_8918,N_5352);
nor U12117 (N_12117,N_5690,N_6946);
or U12118 (N_12118,N_5895,N_6523);
xor U12119 (N_12119,N_5722,N_5851);
nor U12120 (N_12120,N_8622,N_6311);
nand U12121 (N_12121,N_9720,N_9584);
nand U12122 (N_12122,N_7978,N_7433);
nand U12123 (N_12123,N_9467,N_7394);
and U12124 (N_12124,N_8436,N_8273);
and U12125 (N_12125,N_7581,N_6321);
nor U12126 (N_12126,N_6319,N_8417);
and U12127 (N_12127,N_9802,N_8666);
xnor U12128 (N_12128,N_8163,N_9410);
and U12129 (N_12129,N_9873,N_5636);
nand U12130 (N_12130,N_8754,N_5375);
and U12131 (N_12131,N_8698,N_7363);
xor U12132 (N_12132,N_6631,N_6610);
nor U12133 (N_12133,N_8714,N_6960);
nor U12134 (N_12134,N_6956,N_7505);
and U12135 (N_12135,N_5097,N_7896);
nand U12136 (N_12136,N_5623,N_6514);
nor U12137 (N_12137,N_5133,N_8507);
xor U12138 (N_12138,N_5019,N_9779);
nor U12139 (N_12139,N_9405,N_7263);
and U12140 (N_12140,N_6763,N_5050);
nand U12141 (N_12141,N_7431,N_7785);
nand U12142 (N_12142,N_7173,N_6920);
and U12143 (N_12143,N_5093,N_9132);
and U12144 (N_12144,N_9329,N_7656);
nand U12145 (N_12145,N_9008,N_9814);
nor U12146 (N_12146,N_7682,N_5913);
xor U12147 (N_12147,N_7595,N_6995);
xor U12148 (N_12148,N_7420,N_6406);
or U12149 (N_12149,N_8678,N_9388);
xnor U12150 (N_12150,N_9170,N_7460);
or U12151 (N_12151,N_6277,N_9355);
nor U12152 (N_12152,N_6370,N_7339);
and U12153 (N_12153,N_5858,N_9026);
and U12154 (N_12154,N_7113,N_6044);
and U12155 (N_12155,N_9037,N_9312);
nand U12156 (N_12156,N_6977,N_7929);
and U12157 (N_12157,N_6945,N_5744);
nand U12158 (N_12158,N_7430,N_5770);
nor U12159 (N_12159,N_6416,N_9483);
or U12160 (N_12160,N_8299,N_7495);
or U12161 (N_12161,N_9079,N_7256);
and U12162 (N_12162,N_8966,N_9883);
nand U12163 (N_12163,N_6930,N_8608);
and U12164 (N_12164,N_9433,N_5586);
xnor U12165 (N_12165,N_8080,N_7925);
nand U12166 (N_12166,N_5218,N_5298);
nor U12167 (N_12167,N_5390,N_7485);
or U12168 (N_12168,N_5778,N_9911);
and U12169 (N_12169,N_9832,N_8515);
nand U12170 (N_12170,N_5245,N_8475);
and U12171 (N_12171,N_7223,N_8995);
nand U12172 (N_12172,N_5912,N_5573);
nand U12173 (N_12173,N_7171,N_5437);
or U12174 (N_12174,N_9283,N_7814);
xnor U12175 (N_12175,N_6460,N_7023);
xor U12176 (N_12176,N_6476,N_9173);
xnor U12177 (N_12177,N_5361,N_7950);
and U12178 (N_12178,N_6802,N_5285);
xor U12179 (N_12179,N_9791,N_6592);
nand U12180 (N_12180,N_8200,N_9798);
nor U12181 (N_12181,N_9705,N_9617);
nand U12182 (N_12182,N_8873,N_6653);
nand U12183 (N_12183,N_6211,N_8243);
and U12184 (N_12184,N_5952,N_7316);
xor U12185 (N_12185,N_7986,N_8345);
nor U12186 (N_12186,N_8075,N_7968);
xor U12187 (N_12187,N_8145,N_9560);
or U12188 (N_12188,N_5280,N_6326);
nand U12189 (N_12189,N_7331,N_9363);
or U12190 (N_12190,N_8187,N_8901);
nand U12191 (N_12191,N_7082,N_9074);
xnor U12192 (N_12192,N_6563,N_8238);
nand U12193 (N_12193,N_5447,N_6026);
and U12194 (N_12194,N_9194,N_7484);
xor U12195 (N_12195,N_7697,N_8804);
xnor U12196 (N_12196,N_9639,N_7028);
nor U12197 (N_12197,N_7346,N_6685);
xnor U12198 (N_12198,N_9287,N_7830);
or U12199 (N_12199,N_6553,N_9507);
nor U12200 (N_12200,N_6324,N_7832);
and U12201 (N_12201,N_9345,N_7020);
xnor U12202 (N_12202,N_5882,N_8614);
xor U12203 (N_12203,N_7839,N_9044);
or U12204 (N_12204,N_9521,N_6373);
and U12205 (N_12205,N_6881,N_9923);
nor U12206 (N_12206,N_6886,N_6251);
nor U12207 (N_12207,N_7691,N_8910);
xnor U12208 (N_12208,N_9512,N_6191);
or U12209 (N_12209,N_7321,N_8371);
nand U12210 (N_12210,N_5877,N_9330);
xor U12211 (N_12211,N_6375,N_6010);
and U12212 (N_12212,N_5712,N_6079);
nor U12213 (N_12213,N_6297,N_7286);
nand U12214 (N_12214,N_9607,N_6454);
nor U12215 (N_12215,N_5440,N_8235);
nor U12216 (N_12216,N_6425,N_5186);
xor U12217 (N_12217,N_7567,N_9201);
or U12218 (N_12218,N_5382,N_6474);
or U12219 (N_12219,N_5206,N_6168);
and U12220 (N_12220,N_7833,N_6734);
nand U12221 (N_12221,N_5163,N_5491);
nand U12222 (N_12222,N_6578,N_9646);
nand U12223 (N_12223,N_7162,N_9432);
nor U12224 (N_12224,N_8259,N_6722);
nor U12225 (N_12225,N_9246,N_7188);
or U12226 (N_12226,N_7635,N_5448);
xnor U12227 (N_12227,N_7506,N_8840);
nand U12228 (N_12228,N_7698,N_9822);
and U12229 (N_12229,N_5189,N_8018);
or U12230 (N_12230,N_9836,N_6611);
xor U12231 (N_12231,N_6120,N_7935);
and U12232 (N_12232,N_5934,N_5250);
nor U12233 (N_12233,N_8105,N_9486);
and U12234 (N_12234,N_5010,N_6981);
nand U12235 (N_12235,N_6683,N_6053);
or U12236 (N_12236,N_7086,N_7010);
xnor U12237 (N_12237,N_7537,N_8812);
or U12238 (N_12238,N_6670,N_9429);
xnor U12239 (N_12239,N_8332,N_7758);
or U12240 (N_12240,N_5270,N_9210);
nor U12241 (N_12241,N_9860,N_7829);
nand U12242 (N_12242,N_5102,N_9323);
nand U12243 (N_12243,N_8315,N_9736);
nand U12244 (N_12244,N_5103,N_6641);
or U12245 (N_12245,N_8691,N_9089);
nand U12246 (N_12246,N_5723,N_7803);
xor U12247 (N_12247,N_8041,N_5384);
or U12248 (N_12248,N_8787,N_8715);
and U12249 (N_12249,N_5611,N_9839);
or U12250 (N_12250,N_9220,N_5990);
and U12251 (N_12251,N_8566,N_8855);
and U12252 (N_12252,N_6362,N_7606);
nor U12253 (N_12253,N_7672,N_7972);
xnor U12254 (N_12254,N_9774,N_6384);
xor U12255 (N_12255,N_8095,N_5991);
nor U12256 (N_12256,N_5899,N_7461);
xor U12257 (N_12257,N_9490,N_9799);
or U12258 (N_12258,N_6146,N_7018);
and U12259 (N_12259,N_7647,N_8908);
and U12260 (N_12260,N_5290,N_7721);
xor U12261 (N_12261,N_8613,N_7707);
and U12262 (N_12262,N_5515,N_8902);
and U12263 (N_12263,N_8551,N_5557);
nor U12264 (N_12264,N_7865,N_6054);
nand U12265 (N_12265,N_5589,N_9683);
nor U12266 (N_12266,N_8581,N_9278);
or U12267 (N_12267,N_8610,N_9735);
xnor U12268 (N_12268,N_6310,N_7600);
and U12269 (N_12269,N_5827,N_6409);
xnor U12270 (N_12270,N_6535,N_5471);
nand U12271 (N_12271,N_9052,N_9479);
and U12272 (N_12272,N_6298,N_5988);
or U12273 (N_12273,N_5411,N_5000);
nor U12274 (N_12274,N_8513,N_5346);
nand U12275 (N_12275,N_7985,N_9057);
and U12276 (N_12276,N_7699,N_7618);
xor U12277 (N_12277,N_8070,N_8586);
nand U12278 (N_12278,N_9421,N_9027);
nand U12279 (N_12279,N_9140,N_7357);
and U12280 (N_12280,N_5024,N_5817);
and U12281 (N_12281,N_5462,N_9263);
nand U12282 (N_12282,N_7681,N_8866);
and U12283 (N_12283,N_8198,N_9955);
and U12284 (N_12284,N_9161,N_9509);
and U12285 (N_12285,N_8236,N_7055);
or U12286 (N_12286,N_6000,N_5896);
or U12287 (N_12287,N_7846,N_7870);
or U12288 (N_12288,N_7471,N_5214);
nor U12289 (N_12289,N_8314,N_8456);
and U12290 (N_12290,N_5523,N_6996);
nor U12291 (N_12291,N_5734,N_7329);
nand U12292 (N_12292,N_7959,N_5349);
xnor U12293 (N_12293,N_5393,N_6255);
xor U12294 (N_12294,N_6962,N_7556);
and U12295 (N_12295,N_7439,N_5033);
nand U12296 (N_12296,N_6385,N_9066);
xor U12297 (N_12297,N_7375,N_8550);
nor U12298 (N_12298,N_6542,N_6285);
nor U12299 (N_12299,N_9650,N_9290);
xor U12300 (N_12300,N_6951,N_5143);
xnor U12301 (N_12301,N_5531,N_8615);
or U12302 (N_12302,N_5836,N_5602);
nand U12303 (N_12303,N_8364,N_9382);
xor U12304 (N_12304,N_7584,N_7913);
nor U12305 (N_12305,N_9083,N_7302);
and U12306 (N_12306,N_7873,N_6253);
nor U12307 (N_12307,N_9012,N_8267);
xnor U12308 (N_12308,N_5839,N_6086);
or U12309 (N_12309,N_7240,N_9001);
or U12310 (N_12310,N_8831,N_5060);
nor U12311 (N_12311,N_8746,N_5671);
or U12312 (N_12312,N_6147,N_7724);
nand U12313 (N_12313,N_8819,N_9699);
xor U12314 (N_12314,N_7808,N_5374);
nand U12315 (N_12315,N_8393,N_8781);
nand U12316 (N_12316,N_8697,N_7920);
nand U12317 (N_12317,N_6902,N_8178);
xor U12318 (N_12318,N_8937,N_7305);
nor U12319 (N_12319,N_5451,N_7990);
xnor U12320 (N_12320,N_7491,N_9482);
nor U12321 (N_12321,N_6435,N_8148);
xnor U12322 (N_12322,N_7165,N_9555);
or U12323 (N_12323,N_8510,N_6806);
and U12324 (N_12324,N_9457,N_7932);
nor U12325 (N_12325,N_7253,N_8451);
nor U12326 (N_12326,N_6314,N_6466);
and U12327 (N_12327,N_8632,N_5377);
and U12328 (N_12328,N_6100,N_8412);
and U12329 (N_12329,N_8380,N_7877);
nand U12330 (N_12330,N_9857,N_5467);
xnor U12331 (N_12331,N_6527,N_7379);
nor U12332 (N_12332,N_7557,N_5219);
or U12333 (N_12333,N_6344,N_5297);
or U12334 (N_12334,N_6838,N_5716);
or U12335 (N_12335,N_7455,N_5170);
nand U12336 (N_12336,N_8739,N_8368);
nor U12337 (N_12337,N_9827,N_9362);
nor U12338 (N_12338,N_7693,N_6966);
or U12339 (N_12339,N_8421,N_9993);
nor U12340 (N_12340,N_8768,N_7337);
nor U12341 (N_12341,N_6048,N_8898);
or U12342 (N_12342,N_7982,N_6273);
nand U12343 (N_12343,N_6123,N_7917);
nand U12344 (N_12344,N_8757,N_9149);
nand U12345 (N_12345,N_6097,N_9397);
nor U12346 (N_12346,N_5841,N_6925);
and U12347 (N_12347,N_6900,N_5825);
or U12348 (N_12348,N_8979,N_5587);
nor U12349 (N_12349,N_8021,N_5268);
or U12350 (N_12350,N_6878,N_6023);
or U12351 (N_12351,N_8755,N_8869);
nor U12352 (N_12352,N_8591,N_9285);
xnor U12353 (N_12353,N_9729,N_7659);
and U12354 (N_12354,N_8772,N_9124);
nand U12355 (N_12355,N_6381,N_6860);
nor U12356 (N_12356,N_6414,N_6539);
xor U12357 (N_12357,N_9749,N_9641);
nor U12358 (N_12358,N_9809,N_6738);
xor U12359 (N_12359,N_5787,N_9969);
or U12360 (N_12360,N_8003,N_9333);
nor U12361 (N_12361,N_9307,N_6457);
or U12362 (N_12362,N_9088,N_7751);
nor U12363 (N_12363,N_8847,N_7135);
xor U12364 (N_12364,N_9763,N_8653);
xor U12365 (N_12365,N_7623,N_5958);
nor U12366 (N_12366,N_7569,N_8980);
nand U12367 (N_12367,N_8689,N_5241);
and U12368 (N_12368,N_8125,N_8663);
xor U12369 (N_12369,N_7971,N_8762);
nand U12370 (N_12370,N_5634,N_9143);
or U12371 (N_12371,N_7453,N_5360);
or U12372 (N_12372,N_5225,N_9680);
or U12373 (N_12373,N_9826,N_8549);
xnor U12374 (N_12374,N_9166,N_6202);
xor U12375 (N_12375,N_5665,N_5508);
nor U12376 (N_12376,N_8943,N_7874);
nor U12377 (N_12377,N_9171,N_5711);
nand U12378 (N_12378,N_7437,N_6423);
and U12379 (N_12379,N_6545,N_7500);
and U12380 (N_12380,N_9625,N_8767);
nor U12381 (N_12381,N_6183,N_7401);
xor U12382 (N_12382,N_6757,N_6508);
xnor U12383 (N_12383,N_7879,N_7937);
or U12384 (N_12384,N_5719,N_8473);
nand U12385 (N_12385,N_5442,N_8305);
nor U12386 (N_12386,N_6236,N_9859);
nor U12387 (N_12387,N_8841,N_9471);
nor U12388 (N_12388,N_7052,N_5142);
and U12389 (N_12389,N_5030,N_5175);
nor U12390 (N_12390,N_5574,N_7298);
nor U12391 (N_12391,N_9761,N_7708);
and U12392 (N_12392,N_8988,N_9866);
and U12393 (N_12393,N_6032,N_7938);
nand U12394 (N_12394,N_7410,N_6415);
and U12395 (N_12395,N_7307,N_5850);
nand U12396 (N_12396,N_8630,N_9424);
nand U12397 (N_12397,N_9524,N_6646);
nor U12398 (N_12398,N_6587,N_5781);
nor U12399 (N_12399,N_7992,N_8605);
and U12400 (N_12400,N_8171,N_7905);
xor U12401 (N_12401,N_7487,N_9965);
xnor U12402 (N_12402,N_5291,N_6854);
or U12403 (N_12403,N_6501,N_8394);
and U12404 (N_12404,N_6741,N_5981);
xnor U12405 (N_12405,N_6003,N_8570);
nor U12406 (N_12406,N_5809,N_9169);
nor U12407 (N_12407,N_9896,N_5259);
or U12408 (N_12408,N_7525,N_9710);
nor U12409 (N_12409,N_7817,N_8885);
nor U12410 (N_12410,N_6335,N_6192);
nand U12411 (N_12411,N_9162,N_8803);
nor U12412 (N_12412,N_5362,N_9493);
and U12413 (N_12413,N_8096,N_5336);
nor U12414 (N_12414,N_7674,N_5583);
nand U12415 (N_12415,N_6313,N_8452);
xor U12416 (N_12416,N_5058,N_7637);
and U12417 (N_12417,N_5909,N_5276);
or U12418 (N_12418,N_5115,N_9223);
and U12419 (N_12419,N_7397,N_6014);
nor U12420 (N_12420,N_9033,N_8130);
nand U12421 (N_12421,N_5139,N_9103);
or U12422 (N_12422,N_5917,N_9322);
or U12423 (N_12423,N_7585,N_5572);
nor U12424 (N_12424,N_6073,N_8089);
xnor U12425 (N_12425,N_8579,N_7399);
or U12426 (N_12426,N_6013,N_6732);
xnor U12427 (N_12427,N_7939,N_5386);
nand U12428 (N_12428,N_6351,N_9910);
xor U12429 (N_12429,N_9696,N_9202);
xor U12430 (N_12430,N_7998,N_6827);
or U12431 (N_12431,N_9596,N_6549);
nand U12432 (N_12432,N_7923,N_6103);
nand U12433 (N_12433,N_7269,N_5450);
or U12434 (N_12434,N_5422,N_9129);
or U12435 (N_12435,N_8621,N_9047);
or U12436 (N_12436,N_6544,N_7016);
nor U12437 (N_12437,N_6485,N_6157);
and U12438 (N_12438,N_6664,N_9687);
or U12439 (N_12439,N_5663,N_8286);
and U12440 (N_12440,N_5220,N_5548);
and U12441 (N_12441,N_7360,N_5704);
xnor U12442 (N_12442,N_9669,N_9864);
nand U12443 (N_12443,N_6118,N_9837);
or U12444 (N_12444,N_9571,N_6289);
nand U12445 (N_12445,N_9155,N_8014);
and U12446 (N_12446,N_6140,N_8058);
and U12447 (N_12447,N_9025,N_5559);
nor U12448 (N_12448,N_5996,N_6777);
nand U12449 (N_12449,N_7458,N_5243);
nand U12450 (N_12450,N_9243,N_8609);
and U12451 (N_12451,N_5044,N_7702);
xnor U12452 (N_12452,N_7773,N_7741);
xor U12453 (N_12453,N_9366,N_5680);
and U12454 (N_12454,N_7144,N_5795);
and U12455 (N_12455,N_5428,N_9932);
xnor U12456 (N_12456,N_6727,N_6666);
nor U12457 (N_12457,N_7726,N_6111);
or U12458 (N_12458,N_6480,N_7057);
nor U12459 (N_12459,N_6792,N_5748);
and U12460 (N_12460,N_6865,N_5941);
nand U12461 (N_12461,N_5537,N_8906);
nor U12462 (N_12462,N_9069,N_6529);
or U12463 (N_12463,N_7706,N_9789);
nor U12464 (N_12464,N_5977,N_7335);
nor U12465 (N_12465,N_8291,N_8699);
nor U12466 (N_12466,N_7719,N_9767);
xnor U12467 (N_12467,N_6208,N_6569);
or U12468 (N_12468,N_6437,N_6382);
xor U12469 (N_12469,N_8487,N_8519);
and U12470 (N_12470,N_5940,N_6766);
or U12471 (N_12471,N_5581,N_8311);
nand U12472 (N_12472,N_9248,N_8499);
or U12473 (N_12473,N_8700,N_8771);
and U12474 (N_12474,N_7844,N_5488);
or U12475 (N_12475,N_8338,N_9328);
or U12476 (N_12476,N_8946,N_5337);
and U12477 (N_12477,N_6002,N_6778);
and U12478 (N_12478,N_7855,N_8466);
nand U12479 (N_12479,N_9152,N_9277);
nand U12480 (N_12480,N_6210,N_7904);
or U12481 (N_12481,N_8240,N_9021);
xnor U12482 (N_12482,N_8166,N_5824);
and U12483 (N_12483,N_5696,N_8588);
nand U12484 (N_12484,N_9633,N_7526);
nand U12485 (N_12485,N_9298,N_8516);
nand U12486 (N_12486,N_5283,N_8155);
or U12487 (N_12487,N_7313,N_9318);
nand U12488 (N_12488,N_6291,N_9477);
nand U12489 (N_12489,N_8083,N_5886);
or U12490 (N_12490,N_7444,N_8461);
nor U12491 (N_12491,N_9031,N_9034);
xor U12492 (N_12492,N_9848,N_5412);
xnor U12493 (N_12493,N_5957,N_7421);
nand U12494 (N_12494,N_6595,N_5287);
nand U12495 (N_12495,N_9109,N_8066);
xnor U12496 (N_12496,N_9801,N_6305);
and U12497 (N_12497,N_7084,N_6868);
xor U12498 (N_12498,N_9147,N_7227);
nor U12499 (N_12499,N_7017,N_9501);
xnor U12500 (N_12500,N_7666,N_6949);
xor U12501 (N_12501,N_5643,N_6538);
or U12502 (N_12502,N_5194,N_7189);
xor U12503 (N_12503,N_5159,N_5880);
nand U12504 (N_12504,N_8825,N_6467);
nor U12505 (N_12505,N_5588,N_7930);
or U12506 (N_12506,N_9239,N_8123);
xor U12507 (N_12507,N_7043,N_5794);
nand U12508 (N_12508,N_7758,N_9843);
nor U12509 (N_12509,N_8740,N_9150);
nor U12510 (N_12510,N_9581,N_7695);
nor U12511 (N_12511,N_9132,N_9392);
or U12512 (N_12512,N_9043,N_5467);
and U12513 (N_12513,N_7694,N_9911);
nor U12514 (N_12514,N_6055,N_7943);
nand U12515 (N_12515,N_8056,N_5432);
xor U12516 (N_12516,N_9188,N_6085);
nand U12517 (N_12517,N_8019,N_5030);
nor U12518 (N_12518,N_8192,N_8507);
nor U12519 (N_12519,N_8755,N_7982);
xnor U12520 (N_12520,N_9664,N_7622);
and U12521 (N_12521,N_9247,N_8469);
and U12522 (N_12522,N_6922,N_7832);
xnor U12523 (N_12523,N_6425,N_7475);
nand U12524 (N_12524,N_6226,N_9926);
or U12525 (N_12525,N_5886,N_9127);
nor U12526 (N_12526,N_6355,N_6109);
nor U12527 (N_12527,N_8051,N_8956);
xnor U12528 (N_12528,N_9314,N_5313);
nand U12529 (N_12529,N_9766,N_7256);
nor U12530 (N_12530,N_7351,N_5376);
or U12531 (N_12531,N_5430,N_7648);
xnor U12532 (N_12532,N_8647,N_6004);
nand U12533 (N_12533,N_6090,N_7343);
or U12534 (N_12534,N_5194,N_9479);
nand U12535 (N_12535,N_7593,N_6805);
xnor U12536 (N_12536,N_7553,N_6630);
or U12537 (N_12537,N_6052,N_5833);
nor U12538 (N_12538,N_7266,N_6626);
or U12539 (N_12539,N_6632,N_8818);
nor U12540 (N_12540,N_7656,N_6073);
nor U12541 (N_12541,N_7096,N_6481);
xor U12542 (N_12542,N_7158,N_6259);
nand U12543 (N_12543,N_7992,N_7629);
nand U12544 (N_12544,N_5128,N_7653);
nand U12545 (N_12545,N_6758,N_5051);
nand U12546 (N_12546,N_7951,N_8887);
xor U12547 (N_12547,N_7207,N_7658);
and U12548 (N_12548,N_9532,N_9061);
nor U12549 (N_12549,N_7231,N_6932);
nand U12550 (N_12550,N_9530,N_5195);
and U12551 (N_12551,N_7055,N_6817);
nand U12552 (N_12552,N_9961,N_7238);
and U12553 (N_12553,N_7012,N_8892);
xnor U12554 (N_12554,N_5945,N_6430);
nor U12555 (N_12555,N_7878,N_8378);
nor U12556 (N_12556,N_5733,N_8479);
xor U12557 (N_12557,N_8431,N_7194);
nor U12558 (N_12558,N_6915,N_6134);
nor U12559 (N_12559,N_6492,N_6655);
and U12560 (N_12560,N_7139,N_9606);
xnor U12561 (N_12561,N_8287,N_9083);
nand U12562 (N_12562,N_9092,N_7621);
xnor U12563 (N_12563,N_9864,N_7620);
xor U12564 (N_12564,N_5856,N_6827);
nor U12565 (N_12565,N_7054,N_7070);
or U12566 (N_12566,N_7194,N_7615);
or U12567 (N_12567,N_6175,N_5294);
xnor U12568 (N_12568,N_6966,N_7341);
and U12569 (N_12569,N_9789,N_8941);
nand U12570 (N_12570,N_6876,N_9026);
nand U12571 (N_12571,N_5410,N_6402);
nand U12572 (N_12572,N_9886,N_8790);
and U12573 (N_12573,N_6915,N_7940);
nor U12574 (N_12574,N_5473,N_7960);
and U12575 (N_12575,N_8333,N_7692);
nand U12576 (N_12576,N_8177,N_9310);
xnor U12577 (N_12577,N_6540,N_6350);
xnor U12578 (N_12578,N_6774,N_6964);
or U12579 (N_12579,N_6185,N_7385);
or U12580 (N_12580,N_5016,N_6476);
nor U12581 (N_12581,N_5298,N_5612);
nand U12582 (N_12582,N_5391,N_9407);
and U12583 (N_12583,N_5090,N_5726);
xor U12584 (N_12584,N_9207,N_5429);
nand U12585 (N_12585,N_8897,N_8422);
nor U12586 (N_12586,N_6308,N_9556);
or U12587 (N_12587,N_9174,N_8663);
and U12588 (N_12588,N_6308,N_9632);
and U12589 (N_12589,N_9435,N_9498);
nor U12590 (N_12590,N_8283,N_9675);
xnor U12591 (N_12591,N_7485,N_6000);
or U12592 (N_12592,N_6358,N_7996);
and U12593 (N_12593,N_5719,N_9107);
nand U12594 (N_12594,N_5007,N_9832);
xor U12595 (N_12595,N_9548,N_8344);
and U12596 (N_12596,N_7664,N_8274);
nor U12597 (N_12597,N_6377,N_8339);
or U12598 (N_12598,N_9454,N_8438);
and U12599 (N_12599,N_8605,N_7938);
or U12600 (N_12600,N_8697,N_7418);
xnor U12601 (N_12601,N_7120,N_5086);
nor U12602 (N_12602,N_5221,N_7133);
nand U12603 (N_12603,N_5879,N_9344);
or U12604 (N_12604,N_5587,N_8754);
or U12605 (N_12605,N_5263,N_8473);
xor U12606 (N_12606,N_8176,N_5830);
and U12607 (N_12607,N_7715,N_9649);
and U12608 (N_12608,N_8623,N_9613);
and U12609 (N_12609,N_7030,N_9009);
and U12610 (N_12610,N_7988,N_8401);
nand U12611 (N_12611,N_5420,N_5049);
xor U12612 (N_12612,N_5331,N_7043);
nand U12613 (N_12613,N_7677,N_5739);
xor U12614 (N_12614,N_8990,N_8888);
nor U12615 (N_12615,N_7862,N_9407);
nor U12616 (N_12616,N_8009,N_7648);
xnor U12617 (N_12617,N_7531,N_8125);
xnor U12618 (N_12618,N_6372,N_8584);
nor U12619 (N_12619,N_5371,N_9260);
nand U12620 (N_12620,N_7971,N_5389);
xnor U12621 (N_12621,N_7730,N_8714);
nor U12622 (N_12622,N_5072,N_6939);
and U12623 (N_12623,N_7721,N_8624);
nand U12624 (N_12624,N_5127,N_8072);
and U12625 (N_12625,N_5874,N_7528);
nand U12626 (N_12626,N_7204,N_9699);
nand U12627 (N_12627,N_8617,N_7658);
nor U12628 (N_12628,N_6870,N_5007);
nor U12629 (N_12629,N_7408,N_7584);
and U12630 (N_12630,N_6877,N_5210);
xnor U12631 (N_12631,N_8251,N_9035);
nor U12632 (N_12632,N_8757,N_7034);
or U12633 (N_12633,N_8827,N_7173);
and U12634 (N_12634,N_9397,N_8969);
or U12635 (N_12635,N_8672,N_7987);
or U12636 (N_12636,N_9633,N_8170);
or U12637 (N_12637,N_7361,N_5710);
and U12638 (N_12638,N_8020,N_6223);
and U12639 (N_12639,N_5380,N_7952);
and U12640 (N_12640,N_9774,N_6349);
nor U12641 (N_12641,N_8286,N_5725);
nand U12642 (N_12642,N_9054,N_5115);
nor U12643 (N_12643,N_6215,N_6692);
nand U12644 (N_12644,N_6587,N_6135);
or U12645 (N_12645,N_7633,N_7374);
xor U12646 (N_12646,N_9788,N_8580);
xor U12647 (N_12647,N_9968,N_6321);
nor U12648 (N_12648,N_6640,N_9363);
and U12649 (N_12649,N_9177,N_8272);
or U12650 (N_12650,N_5185,N_6131);
nand U12651 (N_12651,N_8452,N_8585);
nor U12652 (N_12652,N_7235,N_5166);
xor U12653 (N_12653,N_8569,N_9238);
nor U12654 (N_12654,N_7987,N_5655);
xor U12655 (N_12655,N_7466,N_9362);
xor U12656 (N_12656,N_6208,N_5312);
or U12657 (N_12657,N_5450,N_5661);
or U12658 (N_12658,N_8489,N_8890);
nor U12659 (N_12659,N_5410,N_6792);
or U12660 (N_12660,N_7411,N_6927);
nand U12661 (N_12661,N_5097,N_7550);
xor U12662 (N_12662,N_8164,N_9642);
nand U12663 (N_12663,N_9346,N_5967);
nand U12664 (N_12664,N_8823,N_8939);
nand U12665 (N_12665,N_8376,N_9827);
or U12666 (N_12666,N_7573,N_8615);
xor U12667 (N_12667,N_8657,N_8263);
nor U12668 (N_12668,N_9591,N_5609);
nor U12669 (N_12669,N_6561,N_8938);
or U12670 (N_12670,N_5052,N_7808);
xnor U12671 (N_12671,N_8119,N_6569);
xor U12672 (N_12672,N_5486,N_5613);
nand U12673 (N_12673,N_7031,N_6659);
and U12674 (N_12674,N_5904,N_9511);
or U12675 (N_12675,N_6930,N_8171);
and U12676 (N_12676,N_6443,N_7334);
and U12677 (N_12677,N_5750,N_8891);
nand U12678 (N_12678,N_7228,N_5469);
and U12679 (N_12679,N_7571,N_5012);
xor U12680 (N_12680,N_6999,N_7628);
and U12681 (N_12681,N_9089,N_5879);
or U12682 (N_12682,N_9225,N_6352);
nand U12683 (N_12683,N_6079,N_9891);
nor U12684 (N_12684,N_9129,N_8873);
xnor U12685 (N_12685,N_8448,N_7522);
nor U12686 (N_12686,N_6203,N_5093);
and U12687 (N_12687,N_7403,N_9018);
or U12688 (N_12688,N_8300,N_7309);
nand U12689 (N_12689,N_6946,N_6056);
or U12690 (N_12690,N_5853,N_8816);
nand U12691 (N_12691,N_6029,N_9963);
xor U12692 (N_12692,N_7485,N_5254);
nand U12693 (N_12693,N_7955,N_5436);
or U12694 (N_12694,N_5327,N_6600);
and U12695 (N_12695,N_9349,N_9007);
nand U12696 (N_12696,N_7602,N_7751);
or U12697 (N_12697,N_7577,N_8474);
nor U12698 (N_12698,N_6739,N_8195);
nor U12699 (N_12699,N_6667,N_7901);
or U12700 (N_12700,N_5484,N_8527);
xor U12701 (N_12701,N_5978,N_6633);
xor U12702 (N_12702,N_9065,N_9931);
nor U12703 (N_12703,N_7629,N_6817);
and U12704 (N_12704,N_7484,N_5311);
or U12705 (N_12705,N_9423,N_5752);
and U12706 (N_12706,N_5702,N_6536);
or U12707 (N_12707,N_8354,N_6233);
or U12708 (N_12708,N_5337,N_8751);
nand U12709 (N_12709,N_8868,N_9874);
nand U12710 (N_12710,N_7359,N_8385);
nor U12711 (N_12711,N_6574,N_7635);
or U12712 (N_12712,N_8436,N_5952);
nor U12713 (N_12713,N_7052,N_5409);
and U12714 (N_12714,N_9446,N_7968);
and U12715 (N_12715,N_5635,N_9039);
nand U12716 (N_12716,N_5424,N_5923);
and U12717 (N_12717,N_9435,N_6744);
or U12718 (N_12718,N_6992,N_6982);
or U12719 (N_12719,N_7778,N_7013);
and U12720 (N_12720,N_7664,N_5597);
and U12721 (N_12721,N_6614,N_8441);
nand U12722 (N_12722,N_7348,N_7208);
nand U12723 (N_12723,N_7479,N_5523);
xor U12724 (N_12724,N_6745,N_6735);
nand U12725 (N_12725,N_8602,N_8383);
xor U12726 (N_12726,N_9021,N_6981);
nor U12727 (N_12727,N_7509,N_5210);
nand U12728 (N_12728,N_8594,N_8988);
xor U12729 (N_12729,N_9084,N_9048);
or U12730 (N_12730,N_5651,N_7545);
or U12731 (N_12731,N_7565,N_9305);
xnor U12732 (N_12732,N_7154,N_6935);
and U12733 (N_12733,N_9663,N_7695);
xor U12734 (N_12734,N_5643,N_7733);
nand U12735 (N_12735,N_6046,N_9899);
nand U12736 (N_12736,N_9174,N_7794);
and U12737 (N_12737,N_6212,N_8028);
nor U12738 (N_12738,N_7635,N_7636);
xor U12739 (N_12739,N_9009,N_5350);
xnor U12740 (N_12740,N_5719,N_5631);
xor U12741 (N_12741,N_5416,N_8569);
and U12742 (N_12742,N_6376,N_7649);
and U12743 (N_12743,N_5650,N_9457);
and U12744 (N_12744,N_8382,N_6619);
nor U12745 (N_12745,N_8374,N_7008);
nand U12746 (N_12746,N_6185,N_9159);
nor U12747 (N_12747,N_8171,N_6762);
nand U12748 (N_12748,N_9197,N_6666);
or U12749 (N_12749,N_7501,N_9977);
nor U12750 (N_12750,N_6722,N_7019);
and U12751 (N_12751,N_5382,N_7206);
nand U12752 (N_12752,N_5763,N_5785);
nand U12753 (N_12753,N_5725,N_5796);
nor U12754 (N_12754,N_8671,N_5117);
or U12755 (N_12755,N_9018,N_6721);
xnor U12756 (N_12756,N_6816,N_7833);
nand U12757 (N_12757,N_7978,N_8294);
or U12758 (N_12758,N_8265,N_8359);
nor U12759 (N_12759,N_7291,N_7027);
nand U12760 (N_12760,N_9633,N_6895);
nor U12761 (N_12761,N_5505,N_9389);
nand U12762 (N_12762,N_8132,N_6939);
or U12763 (N_12763,N_5863,N_5434);
nor U12764 (N_12764,N_8045,N_9416);
nor U12765 (N_12765,N_8130,N_5262);
nand U12766 (N_12766,N_7578,N_5523);
nand U12767 (N_12767,N_9324,N_9419);
xor U12768 (N_12768,N_9566,N_9966);
xnor U12769 (N_12769,N_6989,N_6602);
xor U12770 (N_12770,N_5890,N_9474);
or U12771 (N_12771,N_5970,N_9563);
or U12772 (N_12772,N_8872,N_6526);
or U12773 (N_12773,N_9111,N_6884);
nor U12774 (N_12774,N_6242,N_8394);
xnor U12775 (N_12775,N_5165,N_5727);
nor U12776 (N_12776,N_5227,N_8809);
nand U12777 (N_12777,N_8624,N_8786);
nand U12778 (N_12778,N_6742,N_6724);
nand U12779 (N_12779,N_5523,N_7507);
nand U12780 (N_12780,N_6468,N_8224);
and U12781 (N_12781,N_7705,N_5692);
nand U12782 (N_12782,N_6809,N_8012);
nor U12783 (N_12783,N_5086,N_8950);
and U12784 (N_12784,N_9591,N_9484);
and U12785 (N_12785,N_7275,N_8060);
nand U12786 (N_12786,N_7037,N_5370);
nor U12787 (N_12787,N_9297,N_8282);
and U12788 (N_12788,N_5439,N_6185);
or U12789 (N_12789,N_9038,N_8888);
nor U12790 (N_12790,N_9390,N_7162);
nor U12791 (N_12791,N_9783,N_7580);
and U12792 (N_12792,N_5957,N_5404);
nor U12793 (N_12793,N_9323,N_9015);
or U12794 (N_12794,N_6237,N_7602);
nand U12795 (N_12795,N_8100,N_8811);
and U12796 (N_12796,N_6481,N_6147);
xor U12797 (N_12797,N_8616,N_5348);
and U12798 (N_12798,N_9704,N_6403);
xor U12799 (N_12799,N_9217,N_8964);
xnor U12800 (N_12800,N_6382,N_6991);
or U12801 (N_12801,N_5780,N_7400);
xor U12802 (N_12802,N_7639,N_8461);
and U12803 (N_12803,N_8531,N_9676);
nand U12804 (N_12804,N_9470,N_7918);
xor U12805 (N_12805,N_8222,N_5669);
or U12806 (N_12806,N_5066,N_6731);
nor U12807 (N_12807,N_5217,N_6780);
or U12808 (N_12808,N_5183,N_7367);
or U12809 (N_12809,N_9172,N_5187);
nand U12810 (N_12810,N_6198,N_6410);
nand U12811 (N_12811,N_7508,N_9714);
nand U12812 (N_12812,N_5022,N_9168);
and U12813 (N_12813,N_9656,N_6689);
xnor U12814 (N_12814,N_8218,N_6679);
or U12815 (N_12815,N_5583,N_8562);
and U12816 (N_12816,N_5703,N_5158);
xor U12817 (N_12817,N_8485,N_5685);
and U12818 (N_12818,N_5124,N_9207);
and U12819 (N_12819,N_6489,N_6833);
nor U12820 (N_12820,N_6602,N_7406);
or U12821 (N_12821,N_5143,N_7713);
xor U12822 (N_12822,N_7078,N_8703);
nor U12823 (N_12823,N_6942,N_7407);
xor U12824 (N_12824,N_9522,N_6294);
and U12825 (N_12825,N_7852,N_6915);
and U12826 (N_12826,N_6488,N_7813);
or U12827 (N_12827,N_9644,N_9614);
nand U12828 (N_12828,N_6566,N_9555);
nor U12829 (N_12829,N_7978,N_6457);
or U12830 (N_12830,N_9599,N_8825);
or U12831 (N_12831,N_6014,N_6765);
xnor U12832 (N_12832,N_7335,N_6820);
nand U12833 (N_12833,N_5425,N_8691);
nand U12834 (N_12834,N_8627,N_5274);
and U12835 (N_12835,N_6260,N_7907);
nand U12836 (N_12836,N_9790,N_6959);
and U12837 (N_12837,N_8020,N_8412);
and U12838 (N_12838,N_8187,N_9468);
nor U12839 (N_12839,N_8496,N_6172);
nand U12840 (N_12840,N_9797,N_9722);
nand U12841 (N_12841,N_6041,N_8890);
or U12842 (N_12842,N_9886,N_7203);
xor U12843 (N_12843,N_7326,N_7904);
and U12844 (N_12844,N_8255,N_9123);
or U12845 (N_12845,N_8966,N_9538);
xor U12846 (N_12846,N_5488,N_6529);
nand U12847 (N_12847,N_5676,N_8324);
or U12848 (N_12848,N_5733,N_5998);
nor U12849 (N_12849,N_6307,N_7128);
and U12850 (N_12850,N_8243,N_8823);
nor U12851 (N_12851,N_5577,N_9730);
nor U12852 (N_12852,N_6935,N_9494);
and U12853 (N_12853,N_9986,N_8068);
and U12854 (N_12854,N_9130,N_9743);
nor U12855 (N_12855,N_7835,N_8958);
nor U12856 (N_12856,N_7901,N_9497);
and U12857 (N_12857,N_9621,N_9432);
nand U12858 (N_12858,N_5592,N_6687);
and U12859 (N_12859,N_8996,N_9115);
and U12860 (N_12860,N_9703,N_5438);
nand U12861 (N_12861,N_8734,N_7584);
nor U12862 (N_12862,N_9921,N_6137);
nand U12863 (N_12863,N_7042,N_9951);
or U12864 (N_12864,N_7732,N_8383);
nor U12865 (N_12865,N_8856,N_7934);
nor U12866 (N_12866,N_8993,N_6157);
nand U12867 (N_12867,N_8949,N_6087);
and U12868 (N_12868,N_5171,N_9482);
or U12869 (N_12869,N_8076,N_6895);
or U12870 (N_12870,N_7606,N_9592);
and U12871 (N_12871,N_5675,N_7374);
or U12872 (N_12872,N_8231,N_5367);
or U12873 (N_12873,N_9185,N_5189);
nor U12874 (N_12874,N_5849,N_8840);
nand U12875 (N_12875,N_7036,N_7268);
or U12876 (N_12876,N_6735,N_7526);
xnor U12877 (N_12877,N_5144,N_8234);
xor U12878 (N_12878,N_7803,N_8583);
xor U12879 (N_12879,N_9627,N_9830);
or U12880 (N_12880,N_6048,N_7739);
or U12881 (N_12881,N_6754,N_7920);
nor U12882 (N_12882,N_9944,N_9631);
or U12883 (N_12883,N_8121,N_8153);
and U12884 (N_12884,N_6598,N_9935);
nand U12885 (N_12885,N_9631,N_5863);
nor U12886 (N_12886,N_9224,N_6111);
nand U12887 (N_12887,N_5375,N_8794);
nand U12888 (N_12888,N_8529,N_5568);
nor U12889 (N_12889,N_7586,N_6721);
xnor U12890 (N_12890,N_5045,N_7974);
xor U12891 (N_12891,N_7364,N_8629);
or U12892 (N_12892,N_6289,N_9314);
and U12893 (N_12893,N_6323,N_6081);
nor U12894 (N_12894,N_5025,N_8054);
or U12895 (N_12895,N_9510,N_7979);
nor U12896 (N_12896,N_5030,N_6074);
and U12897 (N_12897,N_8438,N_8717);
nand U12898 (N_12898,N_5895,N_9295);
or U12899 (N_12899,N_5213,N_9524);
nor U12900 (N_12900,N_5405,N_5240);
xor U12901 (N_12901,N_8652,N_9186);
nand U12902 (N_12902,N_7027,N_7920);
nor U12903 (N_12903,N_8564,N_7697);
or U12904 (N_12904,N_7113,N_5411);
or U12905 (N_12905,N_6460,N_8803);
and U12906 (N_12906,N_7777,N_6279);
xnor U12907 (N_12907,N_8990,N_7636);
and U12908 (N_12908,N_8695,N_8100);
nand U12909 (N_12909,N_7390,N_7836);
nand U12910 (N_12910,N_5667,N_6481);
nor U12911 (N_12911,N_8529,N_8768);
nor U12912 (N_12912,N_7719,N_9293);
and U12913 (N_12913,N_5673,N_7123);
xnor U12914 (N_12914,N_9901,N_9204);
xor U12915 (N_12915,N_6189,N_7753);
xnor U12916 (N_12916,N_7102,N_5862);
nand U12917 (N_12917,N_7432,N_8531);
nand U12918 (N_12918,N_9810,N_6891);
and U12919 (N_12919,N_7280,N_7028);
nor U12920 (N_12920,N_8555,N_5088);
or U12921 (N_12921,N_9969,N_8685);
xnor U12922 (N_12922,N_5789,N_7918);
or U12923 (N_12923,N_5915,N_6991);
and U12924 (N_12924,N_7880,N_8230);
nor U12925 (N_12925,N_7867,N_5233);
nand U12926 (N_12926,N_8663,N_8673);
nor U12927 (N_12927,N_9143,N_5688);
nor U12928 (N_12928,N_7327,N_5406);
nand U12929 (N_12929,N_9304,N_5776);
or U12930 (N_12930,N_8645,N_9678);
or U12931 (N_12931,N_6649,N_9606);
xor U12932 (N_12932,N_7513,N_9452);
or U12933 (N_12933,N_8591,N_6113);
xor U12934 (N_12934,N_9620,N_7989);
nor U12935 (N_12935,N_5098,N_8800);
nand U12936 (N_12936,N_8186,N_8125);
nand U12937 (N_12937,N_9961,N_7943);
nand U12938 (N_12938,N_7213,N_9648);
or U12939 (N_12939,N_5269,N_9209);
and U12940 (N_12940,N_6295,N_9985);
nor U12941 (N_12941,N_6907,N_5996);
xor U12942 (N_12942,N_9057,N_9465);
nand U12943 (N_12943,N_8995,N_6663);
nor U12944 (N_12944,N_5471,N_7692);
nor U12945 (N_12945,N_5553,N_7010);
nand U12946 (N_12946,N_8242,N_6085);
xnor U12947 (N_12947,N_7327,N_8990);
and U12948 (N_12948,N_8396,N_5418);
nor U12949 (N_12949,N_8148,N_8769);
xnor U12950 (N_12950,N_5094,N_7008);
xor U12951 (N_12951,N_9827,N_7408);
nor U12952 (N_12952,N_6592,N_5331);
xnor U12953 (N_12953,N_9316,N_6034);
nand U12954 (N_12954,N_5290,N_5086);
nor U12955 (N_12955,N_9946,N_7297);
or U12956 (N_12956,N_5311,N_8098);
xor U12957 (N_12957,N_6868,N_6130);
and U12958 (N_12958,N_5041,N_8662);
or U12959 (N_12959,N_7547,N_5239);
xnor U12960 (N_12960,N_6566,N_8022);
and U12961 (N_12961,N_6659,N_6346);
xnor U12962 (N_12962,N_5477,N_7345);
xnor U12963 (N_12963,N_8282,N_6700);
and U12964 (N_12964,N_5182,N_5540);
or U12965 (N_12965,N_6646,N_8044);
and U12966 (N_12966,N_6456,N_7526);
xnor U12967 (N_12967,N_7071,N_9879);
and U12968 (N_12968,N_7946,N_9133);
and U12969 (N_12969,N_8737,N_5300);
or U12970 (N_12970,N_9914,N_8399);
nand U12971 (N_12971,N_5949,N_7480);
xnor U12972 (N_12972,N_8982,N_8736);
xor U12973 (N_12973,N_6829,N_5192);
or U12974 (N_12974,N_7167,N_5870);
xor U12975 (N_12975,N_6912,N_7435);
and U12976 (N_12976,N_8152,N_5140);
nor U12977 (N_12977,N_6749,N_6131);
and U12978 (N_12978,N_7609,N_5624);
nor U12979 (N_12979,N_6533,N_5599);
xnor U12980 (N_12980,N_9372,N_6537);
or U12981 (N_12981,N_6374,N_5348);
and U12982 (N_12982,N_9991,N_7858);
or U12983 (N_12983,N_9829,N_6570);
xor U12984 (N_12984,N_8271,N_5352);
or U12985 (N_12985,N_7602,N_7929);
nand U12986 (N_12986,N_7105,N_9600);
and U12987 (N_12987,N_5227,N_7870);
xnor U12988 (N_12988,N_6429,N_8895);
and U12989 (N_12989,N_9475,N_7276);
and U12990 (N_12990,N_9772,N_9126);
xor U12991 (N_12991,N_5521,N_9623);
and U12992 (N_12992,N_9403,N_8561);
or U12993 (N_12993,N_9670,N_8755);
and U12994 (N_12994,N_7328,N_5753);
nor U12995 (N_12995,N_7138,N_6528);
nand U12996 (N_12996,N_7885,N_7173);
xor U12997 (N_12997,N_7712,N_9780);
and U12998 (N_12998,N_7957,N_9867);
nor U12999 (N_12999,N_9793,N_6557);
and U13000 (N_13000,N_9407,N_8572);
and U13001 (N_13001,N_8859,N_7355);
xnor U13002 (N_13002,N_7859,N_7492);
or U13003 (N_13003,N_5871,N_8445);
or U13004 (N_13004,N_8025,N_9820);
or U13005 (N_13005,N_7024,N_5438);
xor U13006 (N_13006,N_7712,N_7460);
xor U13007 (N_13007,N_6417,N_6539);
nor U13008 (N_13008,N_6900,N_9803);
nand U13009 (N_13009,N_8586,N_8883);
and U13010 (N_13010,N_5591,N_7364);
nand U13011 (N_13011,N_6163,N_8598);
xor U13012 (N_13012,N_7797,N_5408);
or U13013 (N_13013,N_5557,N_8695);
and U13014 (N_13014,N_7974,N_9888);
and U13015 (N_13015,N_5293,N_7312);
or U13016 (N_13016,N_8297,N_6438);
and U13017 (N_13017,N_8689,N_6600);
or U13018 (N_13018,N_8504,N_5561);
xor U13019 (N_13019,N_8876,N_5676);
xnor U13020 (N_13020,N_9168,N_9198);
xnor U13021 (N_13021,N_5016,N_5067);
xor U13022 (N_13022,N_8563,N_6457);
nor U13023 (N_13023,N_6177,N_8735);
nand U13024 (N_13024,N_7424,N_6054);
nand U13025 (N_13025,N_6523,N_8332);
and U13026 (N_13026,N_5241,N_5686);
and U13027 (N_13027,N_5025,N_5548);
xor U13028 (N_13028,N_8375,N_5871);
nand U13029 (N_13029,N_6280,N_6588);
nor U13030 (N_13030,N_6689,N_9610);
xor U13031 (N_13031,N_8257,N_5015);
nor U13032 (N_13032,N_9365,N_5714);
xor U13033 (N_13033,N_9252,N_5653);
nor U13034 (N_13034,N_8687,N_5863);
nor U13035 (N_13035,N_9944,N_5796);
and U13036 (N_13036,N_9213,N_8500);
xnor U13037 (N_13037,N_8220,N_6434);
and U13038 (N_13038,N_9599,N_7543);
or U13039 (N_13039,N_8402,N_7786);
or U13040 (N_13040,N_5865,N_8760);
nand U13041 (N_13041,N_6778,N_9296);
nor U13042 (N_13042,N_5175,N_6964);
or U13043 (N_13043,N_7024,N_9035);
xnor U13044 (N_13044,N_6050,N_5262);
nor U13045 (N_13045,N_6469,N_8819);
or U13046 (N_13046,N_8817,N_6691);
nand U13047 (N_13047,N_6026,N_5505);
or U13048 (N_13048,N_8187,N_5982);
and U13049 (N_13049,N_9703,N_5236);
xnor U13050 (N_13050,N_6247,N_8798);
nand U13051 (N_13051,N_9238,N_8392);
and U13052 (N_13052,N_8674,N_7722);
nor U13053 (N_13053,N_7122,N_7807);
nor U13054 (N_13054,N_7476,N_9370);
and U13055 (N_13055,N_8353,N_5178);
and U13056 (N_13056,N_9698,N_9725);
nor U13057 (N_13057,N_5135,N_8609);
nor U13058 (N_13058,N_6644,N_7193);
xnor U13059 (N_13059,N_5465,N_9839);
nand U13060 (N_13060,N_5634,N_8376);
or U13061 (N_13061,N_5452,N_6960);
nand U13062 (N_13062,N_5196,N_8598);
or U13063 (N_13063,N_5210,N_7277);
xnor U13064 (N_13064,N_8097,N_5759);
nand U13065 (N_13065,N_5215,N_7243);
and U13066 (N_13066,N_5326,N_7578);
xnor U13067 (N_13067,N_5283,N_9497);
xnor U13068 (N_13068,N_8719,N_7470);
nand U13069 (N_13069,N_6364,N_8507);
xnor U13070 (N_13070,N_6209,N_9854);
or U13071 (N_13071,N_5624,N_9085);
and U13072 (N_13072,N_5876,N_9536);
xnor U13073 (N_13073,N_5503,N_8966);
nor U13074 (N_13074,N_8419,N_6104);
or U13075 (N_13075,N_9757,N_8190);
nor U13076 (N_13076,N_7570,N_7142);
and U13077 (N_13077,N_6735,N_6992);
nor U13078 (N_13078,N_6248,N_7185);
xnor U13079 (N_13079,N_8420,N_9526);
xor U13080 (N_13080,N_5372,N_5414);
and U13081 (N_13081,N_8276,N_7510);
or U13082 (N_13082,N_9368,N_9389);
and U13083 (N_13083,N_5514,N_7148);
or U13084 (N_13084,N_7591,N_9305);
nor U13085 (N_13085,N_5563,N_7106);
nand U13086 (N_13086,N_8051,N_5518);
nand U13087 (N_13087,N_5395,N_7268);
or U13088 (N_13088,N_9781,N_6638);
nor U13089 (N_13089,N_9057,N_7244);
or U13090 (N_13090,N_8391,N_8196);
xnor U13091 (N_13091,N_7371,N_8003);
nor U13092 (N_13092,N_6243,N_5317);
nand U13093 (N_13093,N_9992,N_7899);
nand U13094 (N_13094,N_6399,N_6928);
xnor U13095 (N_13095,N_7848,N_8269);
nand U13096 (N_13096,N_6591,N_8151);
nand U13097 (N_13097,N_5934,N_8872);
nand U13098 (N_13098,N_6951,N_8334);
nand U13099 (N_13099,N_9651,N_9595);
and U13100 (N_13100,N_7533,N_9447);
nor U13101 (N_13101,N_9703,N_9062);
nor U13102 (N_13102,N_8667,N_9508);
or U13103 (N_13103,N_9920,N_9402);
xor U13104 (N_13104,N_6203,N_8574);
or U13105 (N_13105,N_8331,N_8443);
nand U13106 (N_13106,N_8827,N_8920);
and U13107 (N_13107,N_8533,N_5811);
nor U13108 (N_13108,N_6350,N_9679);
xnor U13109 (N_13109,N_7100,N_6574);
nor U13110 (N_13110,N_6581,N_5378);
nand U13111 (N_13111,N_5642,N_7612);
or U13112 (N_13112,N_9219,N_5121);
or U13113 (N_13113,N_9346,N_7906);
nand U13114 (N_13114,N_7191,N_9619);
xor U13115 (N_13115,N_5739,N_7363);
nand U13116 (N_13116,N_9365,N_8394);
or U13117 (N_13117,N_9075,N_5612);
and U13118 (N_13118,N_5260,N_9136);
and U13119 (N_13119,N_9535,N_8473);
or U13120 (N_13120,N_5072,N_5023);
xor U13121 (N_13121,N_7375,N_7957);
xnor U13122 (N_13122,N_9402,N_9407);
or U13123 (N_13123,N_9597,N_8273);
nand U13124 (N_13124,N_6764,N_7329);
nand U13125 (N_13125,N_9178,N_7798);
xor U13126 (N_13126,N_9030,N_9727);
and U13127 (N_13127,N_5882,N_5782);
xor U13128 (N_13128,N_6738,N_6119);
nand U13129 (N_13129,N_8059,N_6862);
and U13130 (N_13130,N_5276,N_9681);
nand U13131 (N_13131,N_9462,N_8825);
and U13132 (N_13132,N_6040,N_6209);
or U13133 (N_13133,N_8174,N_5304);
xnor U13134 (N_13134,N_9405,N_9960);
or U13135 (N_13135,N_7995,N_8260);
xnor U13136 (N_13136,N_9045,N_8073);
or U13137 (N_13137,N_9574,N_7316);
xor U13138 (N_13138,N_5435,N_8009);
nor U13139 (N_13139,N_9050,N_5076);
nand U13140 (N_13140,N_5570,N_8422);
xnor U13141 (N_13141,N_6592,N_6377);
nand U13142 (N_13142,N_6227,N_5850);
or U13143 (N_13143,N_9393,N_8885);
or U13144 (N_13144,N_7533,N_8993);
or U13145 (N_13145,N_5826,N_8918);
nor U13146 (N_13146,N_9469,N_9429);
or U13147 (N_13147,N_5601,N_7905);
and U13148 (N_13148,N_7420,N_5756);
and U13149 (N_13149,N_8780,N_6412);
xnor U13150 (N_13150,N_9097,N_7351);
and U13151 (N_13151,N_5681,N_5667);
xor U13152 (N_13152,N_8929,N_6913);
nor U13153 (N_13153,N_8062,N_5475);
nor U13154 (N_13154,N_8013,N_5013);
and U13155 (N_13155,N_5045,N_6692);
xor U13156 (N_13156,N_9317,N_6374);
and U13157 (N_13157,N_9083,N_9217);
xnor U13158 (N_13158,N_5081,N_7156);
nand U13159 (N_13159,N_9741,N_7992);
nor U13160 (N_13160,N_7205,N_5290);
nand U13161 (N_13161,N_9792,N_7699);
xnor U13162 (N_13162,N_5065,N_5385);
or U13163 (N_13163,N_6421,N_5350);
xnor U13164 (N_13164,N_9005,N_6008);
nor U13165 (N_13165,N_9800,N_5173);
nor U13166 (N_13166,N_7579,N_9718);
and U13167 (N_13167,N_7159,N_7602);
nand U13168 (N_13168,N_5471,N_9566);
xnor U13169 (N_13169,N_5637,N_7580);
xor U13170 (N_13170,N_7087,N_6965);
or U13171 (N_13171,N_8391,N_6758);
or U13172 (N_13172,N_5498,N_9837);
nand U13173 (N_13173,N_8879,N_8860);
xnor U13174 (N_13174,N_9991,N_8202);
xor U13175 (N_13175,N_5954,N_7542);
xor U13176 (N_13176,N_8568,N_8653);
xor U13177 (N_13177,N_6562,N_7719);
xor U13178 (N_13178,N_6154,N_8428);
xor U13179 (N_13179,N_6136,N_6894);
nand U13180 (N_13180,N_5869,N_7292);
xnor U13181 (N_13181,N_7368,N_7773);
nand U13182 (N_13182,N_5133,N_6202);
or U13183 (N_13183,N_8581,N_7786);
nand U13184 (N_13184,N_8422,N_5519);
or U13185 (N_13185,N_6280,N_5407);
or U13186 (N_13186,N_8384,N_5425);
or U13187 (N_13187,N_6223,N_8532);
and U13188 (N_13188,N_5657,N_6034);
nand U13189 (N_13189,N_5974,N_8015);
xor U13190 (N_13190,N_7482,N_8783);
nand U13191 (N_13191,N_7683,N_6016);
nor U13192 (N_13192,N_7245,N_5007);
and U13193 (N_13193,N_9439,N_9384);
and U13194 (N_13194,N_6857,N_6883);
nand U13195 (N_13195,N_9833,N_6824);
or U13196 (N_13196,N_6890,N_7794);
nand U13197 (N_13197,N_9393,N_5471);
and U13198 (N_13198,N_7203,N_9515);
or U13199 (N_13199,N_7246,N_5569);
nand U13200 (N_13200,N_5853,N_6593);
nor U13201 (N_13201,N_8442,N_7805);
and U13202 (N_13202,N_8837,N_5613);
nand U13203 (N_13203,N_8815,N_6426);
xnor U13204 (N_13204,N_8996,N_8328);
nor U13205 (N_13205,N_7642,N_5766);
nand U13206 (N_13206,N_6356,N_5616);
nor U13207 (N_13207,N_6232,N_5657);
nor U13208 (N_13208,N_7059,N_7542);
or U13209 (N_13209,N_7616,N_8811);
or U13210 (N_13210,N_6351,N_7970);
nand U13211 (N_13211,N_9723,N_5870);
nand U13212 (N_13212,N_9305,N_6435);
nor U13213 (N_13213,N_6291,N_9126);
xor U13214 (N_13214,N_8527,N_6274);
or U13215 (N_13215,N_6035,N_7406);
nor U13216 (N_13216,N_7107,N_6148);
or U13217 (N_13217,N_6373,N_7922);
nand U13218 (N_13218,N_9461,N_6825);
xor U13219 (N_13219,N_6549,N_9498);
nand U13220 (N_13220,N_8132,N_6416);
nor U13221 (N_13221,N_5045,N_7112);
xor U13222 (N_13222,N_8988,N_7910);
xor U13223 (N_13223,N_9626,N_5732);
and U13224 (N_13224,N_8163,N_5574);
nand U13225 (N_13225,N_5259,N_8068);
nand U13226 (N_13226,N_6553,N_6060);
nor U13227 (N_13227,N_8836,N_9892);
xor U13228 (N_13228,N_9663,N_6763);
nand U13229 (N_13229,N_9153,N_8721);
nor U13230 (N_13230,N_9223,N_5843);
or U13231 (N_13231,N_7940,N_9781);
or U13232 (N_13232,N_7404,N_8764);
and U13233 (N_13233,N_5342,N_7187);
and U13234 (N_13234,N_8686,N_6748);
nand U13235 (N_13235,N_5109,N_5996);
and U13236 (N_13236,N_6133,N_6039);
nand U13237 (N_13237,N_9297,N_9084);
nand U13238 (N_13238,N_9852,N_8443);
nand U13239 (N_13239,N_7992,N_6664);
or U13240 (N_13240,N_7763,N_6494);
nand U13241 (N_13241,N_5241,N_6958);
and U13242 (N_13242,N_8376,N_5259);
nand U13243 (N_13243,N_5406,N_7599);
or U13244 (N_13244,N_9240,N_5234);
and U13245 (N_13245,N_6212,N_7336);
xor U13246 (N_13246,N_6733,N_6828);
or U13247 (N_13247,N_6738,N_7892);
xnor U13248 (N_13248,N_9046,N_8059);
and U13249 (N_13249,N_5871,N_7522);
or U13250 (N_13250,N_7687,N_8393);
xor U13251 (N_13251,N_8153,N_8722);
and U13252 (N_13252,N_8725,N_9440);
nand U13253 (N_13253,N_7695,N_7826);
or U13254 (N_13254,N_5758,N_6537);
nor U13255 (N_13255,N_8829,N_9041);
xnor U13256 (N_13256,N_5712,N_7140);
and U13257 (N_13257,N_6340,N_7264);
xor U13258 (N_13258,N_5636,N_6658);
and U13259 (N_13259,N_8652,N_9281);
or U13260 (N_13260,N_9986,N_7760);
or U13261 (N_13261,N_5600,N_5983);
nor U13262 (N_13262,N_8882,N_7287);
xor U13263 (N_13263,N_7950,N_9400);
nor U13264 (N_13264,N_9181,N_9645);
nor U13265 (N_13265,N_9818,N_5206);
and U13266 (N_13266,N_8561,N_9432);
nor U13267 (N_13267,N_8604,N_8406);
and U13268 (N_13268,N_6126,N_7327);
xor U13269 (N_13269,N_7006,N_8357);
nor U13270 (N_13270,N_8081,N_6954);
and U13271 (N_13271,N_7780,N_7093);
nor U13272 (N_13272,N_8263,N_6808);
or U13273 (N_13273,N_7026,N_5277);
and U13274 (N_13274,N_9852,N_8527);
or U13275 (N_13275,N_7678,N_9709);
and U13276 (N_13276,N_6381,N_6988);
or U13277 (N_13277,N_7625,N_9463);
nand U13278 (N_13278,N_6678,N_8161);
or U13279 (N_13279,N_5700,N_5541);
or U13280 (N_13280,N_9120,N_5242);
or U13281 (N_13281,N_8565,N_6969);
or U13282 (N_13282,N_9163,N_8748);
nor U13283 (N_13283,N_6562,N_8795);
or U13284 (N_13284,N_8181,N_7884);
or U13285 (N_13285,N_8166,N_5726);
or U13286 (N_13286,N_7056,N_7780);
or U13287 (N_13287,N_8786,N_8319);
and U13288 (N_13288,N_6993,N_9441);
or U13289 (N_13289,N_7524,N_6027);
nand U13290 (N_13290,N_7189,N_6723);
nand U13291 (N_13291,N_9399,N_6067);
nand U13292 (N_13292,N_8367,N_9113);
and U13293 (N_13293,N_8061,N_9999);
nor U13294 (N_13294,N_6461,N_9664);
nor U13295 (N_13295,N_6470,N_7901);
and U13296 (N_13296,N_7954,N_6429);
nand U13297 (N_13297,N_5353,N_6470);
nor U13298 (N_13298,N_9086,N_9765);
nand U13299 (N_13299,N_5562,N_9368);
xnor U13300 (N_13300,N_6462,N_6883);
xnor U13301 (N_13301,N_9971,N_9456);
nor U13302 (N_13302,N_8384,N_5454);
nor U13303 (N_13303,N_8591,N_5112);
nor U13304 (N_13304,N_9700,N_6842);
nor U13305 (N_13305,N_7939,N_8762);
or U13306 (N_13306,N_6706,N_5436);
nand U13307 (N_13307,N_8695,N_6079);
xnor U13308 (N_13308,N_8694,N_6561);
and U13309 (N_13309,N_6326,N_8922);
xor U13310 (N_13310,N_5475,N_6864);
and U13311 (N_13311,N_7039,N_8713);
or U13312 (N_13312,N_6211,N_5194);
xnor U13313 (N_13313,N_9935,N_7730);
nand U13314 (N_13314,N_5715,N_9675);
nand U13315 (N_13315,N_8509,N_5550);
nor U13316 (N_13316,N_5059,N_5347);
nand U13317 (N_13317,N_5246,N_8196);
or U13318 (N_13318,N_5924,N_9042);
xnor U13319 (N_13319,N_7674,N_6139);
nor U13320 (N_13320,N_6771,N_8630);
nand U13321 (N_13321,N_6717,N_8750);
nand U13322 (N_13322,N_7197,N_9364);
nor U13323 (N_13323,N_7813,N_5601);
xnor U13324 (N_13324,N_5009,N_5579);
nand U13325 (N_13325,N_7875,N_8349);
nand U13326 (N_13326,N_9939,N_6639);
xor U13327 (N_13327,N_9590,N_9397);
nor U13328 (N_13328,N_6449,N_6309);
and U13329 (N_13329,N_8084,N_5782);
or U13330 (N_13330,N_6438,N_9167);
nor U13331 (N_13331,N_5456,N_9298);
nor U13332 (N_13332,N_9022,N_7933);
nor U13333 (N_13333,N_7842,N_8337);
nor U13334 (N_13334,N_7979,N_9100);
and U13335 (N_13335,N_7942,N_5525);
and U13336 (N_13336,N_8745,N_5447);
nand U13337 (N_13337,N_5029,N_9295);
xnor U13338 (N_13338,N_8166,N_7407);
or U13339 (N_13339,N_5083,N_5817);
xnor U13340 (N_13340,N_6301,N_5969);
nor U13341 (N_13341,N_9817,N_8837);
nor U13342 (N_13342,N_6646,N_8233);
nand U13343 (N_13343,N_6066,N_6084);
nor U13344 (N_13344,N_5286,N_9751);
and U13345 (N_13345,N_8272,N_6349);
xor U13346 (N_13346,N_5839,N_5206);
and U13347 (N_13347,N_5525,N_9614);
and U13348 (N_13348,N_6565,N_9938);
xor U13349 (N_13349,N_7012,N_9577);
and U13350 (N_13350,N_5016,N_7379);
or U13351 (N_13351,N_8818,N_7185);
and U13352 (N_13352,N_9502,N_8574);
and U13353 (N_13353,N_5806,N_5997);
nor U13354 (N_13354,N_5034,N_5282);
nand U13355 (N_13355,N_9948,N_8940);
xnor U13356 (N_13356,N_5734,N_5324);
or U13357 (N_13357,N_7892,N_5024);
nor U13358 (N_13358,N_8171,N_5956);
or U13359 (N_13359,N_5218,N_7365);
nor U13360 (N_13360,N_7572,N_8161);
and U13361 (N_13361,N_7110,N_7615);
and U13362 (N_13362,N_8295,N_6841);
xnor U13363 (N_13363,N_7333,N_7027);
or U13364 (N_13364,N_9392,N_6684);
nor U13365 (N_13365,N_9898,N_5800);
xor U13366 (N_13366,N_9478,N_5595);
xor U13367 (N_13367,N_5104,N_7050);
xor U13368 (N_13368,N_6124,N_9157);
or U13369 (N_13369,N_6891,N_7173);
xnor U13370 (N_13370,N_6115,N_7704);
and U13371 (N_13371,N_7525,N_5134);
and U13372 (N_13372,N_5131,N_6890);
xnor U13373 (N_13373,N_5463,N_5895);
nand U13374 (N_13374,N_7120,N_7148);
xnor U13375 (N_13375,N_8063,N_8378);
nand U13376 (N_13376,N_5922,N_6707);
or U13377 (N_13377,N_9137,N_7914);
and U13378 (N_13378,N_5883,N_9028);
nor U13379 (N_13379,N_9403,N_8917);
or U13380 (N_13380,N_5780,N_6671);
xnor U13381 (N_13381,N_6237,N_9281);
and U13382 (N_13382,N_8079,N_6234);
xor U13383 (N_13383,N_5852,N_9802);
nor U13384 (N_13384,N_7194,N_9054);
and U13385 (N_13385,N_9674,N_9355);
and U13386 (N_13386,N_5782,N_5436);
or U13387 (N_13387,N_5235,N_6003);
xnor U13388 (N_13388,N_7391,N_5461);
or U13389 (N_13389,N_5238,N_5596);
or U13390 (N_13390,N_8890,N_7591);
and U13391 (N_13391,N_7663,N_9058);
nand U13392 (N_13392,N_8423,N_8851);
nor U13393 (N_13393,N_6365,N_9718);
nor U13394 (N_13394,N_6890,N_5398);
nand U13395 (N_13395,N_7059,N_5617);
nor U13396 (N_13396,N_8698,N_6122);
or U13397 (N_13397,N_8072,N_6791);
or U13398 (N_13398,N_7553,N_6664);
and U13399 (N_13399,N_9108,N_7660);
and U13400 (N_13400,N_7469,N_6123);
nand U13401 (N_13401,N_7769,N_9540);
xor U13402 (N_13402,N_6793,N_7222);
nand U13403 (N_13403,N_9617,N_9100);
nor U13404 (N_13404,N_9494,N_9506);
nand U13405 (N_13405,N_9519,N_9759);
xnor U13406 (N_13406,N_7110,N_9981);
and U13407 (N_13407,N_8199,N_6332);
nand U13408 (N_13408,N_6603,N_5779);
or U13409 (N_13409,N_6450,N_9164);
nor U13410 (N_13410,N_6751,N_6382);
xnor U13411 (N_13411,N_6404,N_7291);
nand U13412 (N_13412,N_5339,N_8366);
and U13413 (N_13413,N_7555,N_9096);
nor U13414 (N_13414,N_5913,N_8781);
xor U13415 (N_13415,N_8663,N_8304);
nor U13416 (N_13416,N_5751,N_9604);
xor U13417 (N_13417,N_9129,N_6499);
and U13418 (N_13418,N_9665,N_8226);
nor U13419 (N_13419,N_7570,N_5026);
or U13420 (N_13420,N_6296,N_5129);
nor U13421 (N_13421,N_5502,N_8517);
and U13422 (N_13422,N_5441,N_7262);
and U13423 (N_13423,N_5214,N_7024);
or U13424 (N_13424,N_5452,N_7823);
nor U13425 (N_13425,N_8480,N_7850);
nor U13426 (N_13426,N_7371,N_5995);
nand U13427 (N_13427,N_5565,N_7593);
xnor U13428 (N_13428,N_8890,N_6997);
or U13429 (N_13429,N_5767,N_9929);
nor U13430 (N_13430,N_9424,N_5081);
or U13431 (N_13431,N_7678,N_7113);
nor U13432 (N_13432,N_7802,N_5174);
and U13433 (N_13433,N_7305,N_6121);
nor U13434 (N_13434,N_9080,N_9947);
nor U13435 (N_13435,N_8824,N_9307);
and U13436 (N_13436,N_9386,N_6984);
nor U13437 (N_13437,N_7380,N_6522);
xnor U13438 (N_13438,N_7256,N_5630);
and U13439 (N_13439,N_6202,N_6325);
xor U13440 (N_13440,N_6737,N_7088);
nor U13441 (N_13441,N_7077,N_8605);
xor U13442 (N_13442,N_5701,N_5629);
and U13443 (N_13443,N_9894,N_6675);
nor U13444 (N_13444,N_8581,N_7448);
nor U13445 (N_13445,N_5202,N_6894);
nand U13446 (N_13446,N_9477,N_5492);
nor U13447 (N_13447,N_6242,N_5382);
or U13448 (N_13448,N_7480,N_5830);
xor U13449 (N_13449,N_6028,N_5561);
and U13450 (N_13450,N_8791,N_5942);
and U13451 (N_13451,N_8303,N_9121);
nand U13452 (N_13452,N_6365,N_6488);
and U13453 (N_13453,N_7729,N_6820);
nand U13454 (N_13454,N_5203,N_6598);
and U13455 (N_13455,N_7059,N_9853);
nor U13456 (N_13456,N_9563,N_5258);
or U13457 (N_13457,N_8167,N_8929);
and U13458 (N_13458,N_9878,N_8001);
xor U13459 (N_13459,N_7635,N_9582);
nor U13460 (N_13460,N_7137,N_6734);
nand U13461 (N_13461,N_9128,N_9197);
or U13462 (N_13462,N_8685,N_5419);
or U13463 (N_13463,N_9602,N_9937);
xnor U13464 (N_13464,N_7260,N_8851);
xor U13465 (N_13465,N_8575,N_6409);
nor U13466 (N_13466,N_8891,N_6423);
and U13467 (N_13467,N_6241,N_6849);
nand U13468 (N_13468,N_5204,N_6755);
xor U13469 (N_13469,N_6825,N_7828);
and U13470 (N_13470,N_8915,N_6201);
nor U13471 (N_13471,N_6272,N_5499);
nor U13472 (N_13472,N_8884,N_6305);
or U13473 (N_13473,N_7350,N_5702);
xnor U13474 (N_13474,N_7053,N_9500);
and U13475 (N_13475,N_8580,N_8281);
or U13476 (N_13476,N_7920,N_9686);
nor U13477 (N_13477,N_5667,N_6001);
xor U13478 (N_13478,N_8263,N_7027);
nand U13479 (N_13479,N_6704,N_6070);
and U13480 (N_13480,N_8023,N_8267);
xnor U13481 (N_13481,N_7453,N_8363);
or U13482 (N_13482,N_5838,N_7857);
or U13483 (N_13483,N_8393,N_6722);
xor U13484 (N_13484,N_7431,N_9226);
nand U13485 (N_13485,N_7195,N_9106);
nor U13486 (N_13486,N_7030,N_9109);
nand U13487 (N_13487,N_7517,N_6154);
nor U13488 (N_13488,N_9504,N_6065);
and U13489 (N_13489,N_9534,N_8226);
nor U13490 (N_13490,N_9635,N_8319);
nand U13491 (N_13491,N_6663,N_9159);
xnor U13492 (N_13492,N_9097,N_6683);
and U13493 (N_13493,N_6208,N_7454);
and U13494 (N_13494,N_5983,N_5808);
or U13495 (N_13495,N_8145,N_7377);
nand U13496 (N_13496,N_9733,N_9814);
nand U13497 (N_13497,N_9185,N_6979);
nor U13498 (N_13498,N_7307,N_9093);
or U13499 (N_13499,N_6288,N_6577);
and U13500 (N_13500,N_5206,N_7382);
nand U13501 (N_13501,N_7057,N_7621);
or U13502 (N_13502,N_7074,N_9298);
or U13503 (N_13503,N_8291,N_9076);
or U13504 (N_13504,N_7840,N_8012);
or U13505 (N_13505,N_8635,N_7245);
and U13506 (N_13506,N_9170,N_6093);
or U13507 (N_13507,N_7606,N_8791);
nor U13508 (N_13508,N_6242,N_5985);
nor U13509 (N_13509,N_7944,N_7775);
and U13510 (N_13510,N_9085,N_8134);
nand U13511 (N_13511,N_8833,N_5750);
and U13512 (N_13512,N_8106,N_8358);
nor U13513 (N_13513,N_9067,N_7225);
xor U13514 (N_13514,N_6465,N_7240);
xor U13515 (N_13515,N_5638,N_9193);
nor U13516 (N_13516,N_5948,N_7585);
and U13517 (N_13517,N_7358,N_6936);
and U13518 (N_13518,N_7242,N_6224);
xor U13519 (N_13519,N_5243,N_7165);
nand U13520 (N_13520,N_9929,N_7697);
nand U13521 (N_13521,N_8975,N_7945);
nand U13522 (N_13522,N_9837,N_7624);
nor U13523 (N_13523,N_7890,N_5523);
xor U13524 (N_13524,N_8419,N_8354);
or U13525 (N_13525,N_6027,N_5757);
nor U13526 (N_13526,N_9151,N_9858);
xnor U13527 (N_13527,N_9773,N_5744);
nand U13528 (N_13528,N_9425,N_8387);
nor U13529 (N_13529,N_5418,N_8336);
or U13530 (N_13530,N_9619,N_7490);
xnor U13531 (N_13531,N_6480,N_9745);
nand U13532 (N_13532,N_5314,N_5801);
xor U13533 (N_13533,N_7989,N_8732);
nand U13534 (N_13534,N_5554,N_6124);
xor U13535 (N_13535,N_7077,N_7353);
nand U13536 (N_13536,N_9774,N_8265);
and U13537 (N_13537,N_7893,N_9271);
or U13538 (N_13538,N_7229,N_8894);
nand U13539 (N_13539,N_9849,N_5052);
nor U13540 (N_13540,N_8083,N_5279);
xor U13541 (N_13541,N_8657,N_9081);
nor U13542 (N_13542,N_8353,N_9413);
nand U13543 (N_13543,N_7303,N_5422);
or U13544 (N_13544,N_7171,N_6900);
nor U13545 (N_13545,N_6762,N_6319);
and U13546 (N_13546,N_5115,N_9851);
nor U13547 (N_13547,N_7256,N_7299);
nor U13548 (N_13548,N_6450,N_6336);
nand U13549 (N_13549,N_8228,N_7213);
xor U13550 (N_13550,N_8666,N_9438);
nand U13551 (N_13551,N_5810,N_9755);
xnor U13552 (N_13552,N_9311,N_8788);
nand U13553 (N_13553,N_9515,N_5125);
nor U13554 (N_13554,N_7876,N_9375);
or U13555 (N_13555,N_9208,N_6710);
nand U13556 (N_13556,N_5588,N_7587);
nor U13557 (N_13557,N_9928,N_6338);
and U13558 (N_13558,N_5908,N_8081);
xnor U13559 (N_13559,N_7763,N_6363);
nand U13560 (N_13560,N_9725,N_8668);
nor U13561 (N_13561,N_6500,N_6741);
and U13562 (N_13562,N_5662,N_8184);
nand U13563 (N_13563,N_6229,N_9447);
or U13564 (N_13564,N_9075,N_6235);
xnor U13565 (N_13565,N_8363,N_5900);
or U13566 (N_13566,N_5684,N_7716);
and U13567 (N_13567,N_7740,N_6059);
xnor U13568 (N_13568,N_9935,N_7731);
nor U13569 (N_13569,N_9614,N_5318);
and U13570 (N_13570,N_8373,N_5403);
or U13571 (N_13571,N_7697,N_8906);
and U13572 (N_13572,N_6193,N_8736);
or U13573 (N_13573,N_9989,N_5432);
xor U13574 (N_13574,N_6632,N_5809);
nor U13575 (N_13575,N_6324,N_5909);
xnor U13576 (N_13576,N_5183,N_9571);
xor U13577 (N_13577,N_6239,N_6148);
nand U13578 (N_13578,N_8364,N_7439);
nor U13579 (N_13579,N_6828,N_9716);
nand U13580 (N_13580,N_9587,N_6679);
or U13581 (N_13581,N_5013,N_7563);
or U13582 (N_13582,N_8768,N_7119);
nand U13583 (N_13583,N_5478,N_6514);
and U13584 (N_13584,N_9689,N_7179);
nor U13585 (N_13585,N_6943,N_5805);
or U13586 (N_13586,N_7140,N_5949);
or U13587 (N_13587,N_5859,N_8381);
nor U13588 (N_13588,N_9989,N_5820);
or U13589 (N_13589,N_7131,N_6227);
nor U13590 (N_13590,N_5342,N_9246);
and U13591 (N_13591,N_9514,N_8426);
and U13592 (N_13592,N_5339,N_8635);
or U13593 (N_13593,N_7117,N_8710);
nor U13594 (N_13594,N_5755,N_9443);
or U13595 (N_13595,N_8930,N_6641);
nor U13596 (N_13596,N_5876,N_7443);
and U13597 (N_13597,N_9100,N_8489);
nand U13598 (N_13598,N_9647,N_5657);
nand U13599 (N_13599,N_5534,N_6887);
or U13600 (N_13600,N_9786,N_9514);
nand U13601 (N_13601,N_5752,N_7746);
and U13602 (N_13602,N_5317,N_7018);
nor U13603 (N_13603,N_7862,N_8976);
and U13604 (N_13604,N_9999,N_9748);
nor U13605 (N_13605,N_8079,N_7268);
nand U13606 (N_13606,N_5928,N_7829);
nand U13607 (N_13607,N_7798,N_9616);
or U13608 (N_13608,N_5516,N_6499);
nor U13609 (N_13609,N_5919,N_9567);
nor U13610 (N_13610,N_7095,N_9032);
nand U13611 (N_13611,N_9902,N_7812);
or U13612 (N_13612,N_9494,N_6465);
and U13613 (N_13613,N_9244,N_8812);
or U13614 (N_13614,N_9123,N_9483);
nand U13615 (N_13615,N_5427,N_9646);
nand U13616 (N_13616,N_8621,N_7099);
xor U13617 (N_13617,N_8836,N_6953);
nor U13618 (N_13618,N_5774,N_9745);
and U13619 (N_13619,N_6710,N_7110);
nor U13620 (N_13620,N_6548,N_7113);
nor U13621 (N_13621,N_7794,N_6748);
or U13622 (N_13622,N_7986,N_8661);
or U13623 (N_13623,N_5159,N_7232);
nand U13624 (N_13624,N_7564,N_6988);
nand U13625 (N_13625,N_6620,N_5419);
nor U13626 (N_13626,N_5461,N_5426);
nand U13627 (N_13627,N_5365,N_9005);
nand U13628 (N_13628,N_7282,N_8951);
xnor U13629 (N_13629,N_7514,N_8182);
and U13630 (N_13630,N_7613,N_8593);
or U13631 (N_13631,N_8840,N_5981);
nor U13632 (N_13632,N_8715,N_5406);
nand U13633 (N_13633,N_7090,N_5133);
and U13634 (N_13634,N_7653,N_8201);
and U13635 (N_13635,N_9536,N_5543);
nor U13636 (N_13636,N_7823,N_6460);
and U13637 (N_13637,N_9519,N_5689);
xnor U13638 (N_13638,N_9905,N_9812);
and U13639 (N_13639,N_8615,N_8705);
nor U13640 (N_13640,N_8738,N_5412);
nor U13641 (N_13641,N_7857,N_7620);
nand U13642 (N_13642,N_5577,N_8581);
nand U13643 (N_13643,N_7353,N_5431);
or U13644 (N_13644,N_5172,N_7333);
and U13645 (N_13645,N_9228,N_9715);
or U13646 (N_13646,N_5278,N_8929);
xnor U13647 (N_13647,N_6501,N_7576);
or U13648 (N_13648,N_5238,N_9383);
xnor U13649 (N_13649,N_9558,N_6685);
nand U13650 (N_13650,N_8723,N_9131);
or U13651 (N_13651,N_7320,N_5625);
nor U13652 (N_13652,N_5734,N_5234);
xor U13653 (N_13653,N_7703,N_7081);
and U13654 (N_13654,N_9217,N_6088);
xor U13655 (N_13655,N_5312,N_6241);
nand U13656 (N_13656,N_7988,N_8900);
nor U13657 (N_13657,N_6180,N_7518);
nor U13658 (N_13658,N_8828,N_6872);
nand U13659 (N_13659,N_9752,N_9331);
nand U13660 (N_13660,N_8175,N_8775);
nor U13661 (N_13661,N_7452,N_5796);
xnor U13662 (N_13662,N_9876,N_7642);
nor U13663 (N_13663,N_8104,N_9469);
xor U13664 (N_13664,N_5082,N_9052);
or U13665 (N_13665,N_7968,N_8987);
and U13666 (N_13666,N_7034,N_8405);
or U13667 (N_13667,N_7114,N_5312);
or U13668 (N_13668,N_9377,N_5141);
xor U13669 (N_13669,N_9308,N_8515);
or U13670 (N_13670,N_9097,N_9377);
or U13671 (N_13671,N_6094,N_6823);
or U13672 (N_13672,N_7376,N_5928);
or U13673 (N_13673,N_6337,N_5752);
or U13674 (N_13674,N_6015,N_6831);
or U13675 (N_13675,N_6765,N_6718);
xor U13676 (N_13676,N_7677,N_7955);
and U13677 (N_13677,N_8629,N_6053);
or U13678 (N_13678,N_7193,N_6576);
nand U13679 (N_13679,N_7964,N_8873);
nand U13680 (N_13680,N_7291,N_7990);
or U13681 (N_13681,N_9523,N_9029);
nand U13682 (N_13682,N_5878,N_5359);
and U13683 (N_13683,N_6180,N_7394);
and U13684 (N_13684,N_7154,N_6276);
nor U13685 (N_13685,N_7096,N_6658);
nor U13686 (N_13686,N_9897,N_6894);
and U13687 (N_13687,N_9393,N_6817);
or U13688 (N_13688,N_7010,N_9169);
or U13689 (N_13689,N_6621,N_5065);
xnor U13690 (N_13690,N_5132,N_5727);
xnor U13691 (N_13691,N_9308,N_9281);
nand U13692 (N_13692,N_5448,N_9172);
nor U13693 (N_13693,N_8307,N_5470);
nand U13694 (N_13694,N_9066,N_8254);
nand U13695 (N_13695,N_9560,N_5148);
nor U13696 (N_13696,N_8836,N_6942);
and U13697 (N_13697,N_6794,N_5466);
nor U13698 (N_13698,N_7306,N_6238);
nand U13699 (N_13699,N_9316,N_5904);
or U13700 (N_13700,N_7354,N_5873);
or U13701 (N_13701,N_6725,N_7979);
xor U13702 (N_13702,N_7617,N_6294);
nor U13703 (N_13703,N_9197,N_6345);
and U13704 (N_13704,N_6820,N_7765);
nor U13705 (N_13705,N_5666,N_5561);
and U13706 (N_13706,N_5133,N_5142);
or U13707 (N_13707,N_7373,N_7203);
and U13708 (N_13708,N_6563,N_8932);
xnor U13709 (N_13709,N_8619,N_7603);
xnor U13710 (N_13710,N_9085,N_6518);
xor U13711 (N_13711,N_7088,N_8446);
nor U13712 (N_13712,N_8926,N_5423);
xnor U13713 (N_13713,N_8260,N_7485);
or U13714 (N_13714,N_5738,N_6770);
nor U13715 (N_13715,N_7045,N_7572);
and U13716 (N_13716,N_6839,N_7275);
xnor U13717 (N_13717,N_8578,N_5678);
and U13718 (N_13718,N_7995,N_8706);
nor U13719 (N_13719,N_8369,N_8902);
and U13720 (N_13720,N_6304,N_8468);
xor U13721 (N_13721,N_8933,N_6355);
xor U13722 (N_13722,N_7142,N_7669);
and U13723 (N_13723,N_7400,N_6197);
nor U13724 (N_13724,N_7207,N_5550);
nor U13725 (N_13725,N_8332,N_5814);
nor U13726 (N_13726,N_8897,N_6533);
or U13727 (N_13727,N_6983,N_8876);
nor U13728 (N_13728,N_7574,N_9079);
or U13729 (N_13729,N_9291,N_9668);
nand U13730 (N_13730,N_9574,N_9127);
nand U13731 (N_13731,N_5167,N_5020);
xnor U13732 (N_13732,N_7276,N_9078);
nor U13733 (N_13733,N_5025,N_9260);
and U13734 (N_13734,N_7577,N_7297);
nand U13735 (N_13735,N_7890,N_9080);
or U13736 (N_13736,N_7552,N_6897);
or U13737 (N_13737,N_6382,N_9886);
or U13738 (N_13738,N_6459,N_7134);
or U13739 (N_13739,N_8496,N_6976);
or U13740 (N_13740,N_9695,N_8504);
nor U13741 (N_13741,N_6842,N_7357);
nand U13742 (N_13742,N_7116,N_8903);
or U13743 (N_13743,N_6778,N_6783);
nand U13744 (N_13744,N_9465,N_6217);
or U13745 (N_13745,N_7193,N_8341);
nand U13746 (N_13746,N_5701,N_5585);
and U13747 (N_13747,N_9177,N_5037);
and U13748 (N_13748,N_9870,N_7452);
xor U13749 (N_13749,N_6031,N_9984);
nand U13750 (N_13750,N_5865,N_5795);
nand U13751 (N_13751,N_7618,N_8880);
nor U13752 (N_13752,N_5223,N_7398);
and U13753 (N_13753,N_6119,N_5164);
or U13754 (N_13754,N_5547,N_7444);
nor U13755 (N_13755,N_7689,N_6418);
and U13756 (N_13756,N_5787,N_5201);
or U13757 (N_13757,N_9809,N_8771);
or U13758 (N_13758,N_5528,N_6905);
or U13759 (N_13759,N_7672,N_9587);
nand U13760 (N_13760,N_5039,N_8682);
or U13761 (N_13761,N_6721,N_5402);
xnor U13762 (N_13762,N_5922,N_8590);
or U13763 (N_13763,N_9128,N_8165);
nand U13764 (N_13764,N_5411,N_6515);
and U13765 (N_13765,N_7339,N_6259);
nor U13766 (N_13766,N_9847,N_9867);
or U13767 (N_13767,N_6427,N_8317);
or U13768 (N_13768,N_7919,N_7191);
or U13769 (N_13769,N_7911,N_6891);
xor U13770 (N_13770,N_8604,N_8974);
or U13771 (N_13771,N_5572,N_8956);
and U13772 (N_13772,N_6483,N_9548);
nand U13773 (N_13773,N_5052,N_5842);
and U13774 (N_13774,N_8965,N_9295);
or U13775 (N_13775,N_8641,N_5769);
xor U13776 (N_13776,N_5971,N_8177);
or U13777 (N_13777,N_6152,N_9505);
xnor U13778 (N_13778,N_7797,N_6015);
and U13779 (N_13779,N_9706,N_5298);
nor U13780 (N_13780,N_8450,N_7977);
and U13781 (N_13781,N_8810,N_6287);
nor U13782 (N_13782,N_9928,N_5484);
and U13783 (N_13783,N_8173,N_9947);
and U13784 (N_13784,N_9854,N_7088);
or U13785 (N_13785,N_7218,N_6565);
and U13786 (N_13786,N_7334,N_7623);
nand U13787 (N_13787,N_8793,N_7256);
or U13788 (N_13788,N_9741,N_8799);
nand U13789 (N_13789,N_8629,N_9529);
nor U13790 (N_13790,N_8684,N_8081);
or U13791 (N_13791,N_6740,N_9561);
nand U13792 (N_13792,N_7396,N_6922);
xnor U13793 (N_13793,N_5365,N_8088);
or U13794 (N_13794,N_8394,N_7647);
xnor U13795 (N_13795,N_6511,N_5164);
or U13796 (N_13796,N_7937,N_5565);
nand U13797 (N_13797,N_6485,N_6339);
nand U13798 (N_13798,N_9897,N_7821);
nand U13799 (N_13799,N_8975,N_7450);
and U13800 (N_13800,N_7834,N_6415);
and U13801 (N_13801,N_5534,N_8994);
nand U13802 (N_13802,N_8621,N_5329);
xnor U13803 (N_13803,N_5085,N_9028);
xnor U13804 (N_13804,N_6161,N_8626);
xnor U13805 (N_13805,N_8171,N_7256);
xor U13806 (N_13806,N_9637,N_5818);
and U13807 (N_13807,N_7621,N_9738);
xnor U13808 (N_13808,N_8406,N_8817);
or U13809 (N_13809,N_9774,N_7764);
xnor U13810 (N_13810,N_8530,N_7828);
nand U13811 (N_13811,N_5376,N_7205);
nor U13812 (N_13812,N_5026,N_7425);
and U13813 (N_13813,N_6274,N_5839);
or U13814 (N_13814,N_9994,N_6331);
nor U13815 (N_13815,N_6365,N_5203);
nor U13816 (N_13816,N_8396,N_5521);
xor U13817 (N_13817,N_8017,N_8319);
xor U13818 (N_13818,N_7876,N_7197);
xnor U13819 (N_13819,N_5093,N_8192);
and U13820 (N_13820,N_7815,N_5106);
nor U13821 (N_13821,N_6027,N_5539);
and U13822 (N_13822,N_8315,N_5575);
and U13823 (N_13823,N_6446,N_9879);
xnor U13824 (N_13824,N_5308,N_8020);
nor U13825 (N_13825,N_9084,N_8011);
nor U13826 (N_13826,N_7873,N_5190);
and U13827 (N_13827,N_7211,N_5966);
nand U13828 (N_13828,N_5005,N_8013);
or U13829 (N_13829,N_8116,N_6389);
or U13830 (N_13830,N_5614,N_7089);
or U13831 (N_13831,N_6678,N_6277);
nor U13832 (N_13832,N_7427,N_5920);
xnor U13833 (N_13833,N_9699,N_8033);
xor U13834 (N_13834,N_8325,N_9074);
or U13835 (N_13835,N_7892,N_5906);
or U13836 (N_13836,N_6596,N_9691);
xor U13837 (N_13837,N_5565,N_7521);
and U13838 (N_13838,N_6369,N_8596);
nand U13839 (N_13839,N_6000,N_7113);
or U13840 (N_13840,N_6735,N_9191);
or U13841 (N_13841,N_5292,N_8783);
or U13842 (N_13842,N_8816,N_7067);
nor U13843 (N_13843,N_5359,N_7935);
nand U13844 (N_13844,N_9483,N_7187);
and U13845 (N_13845,N_7354,N_7185);
or U13846 (N_13846,N_6307,N_7368);
and U13847 (N_13847,N_5226,N_5768);
nand U13848 (N_13848,N_7104,N_7785);
and U13849 (N_13849,N_8913,N_9450);
nor U13850 (N_13850,N_8641,N_5820);
xor U13851 (N_13851,N_6191,N_6430);
nor U13852 (N_13852,N_5607,N_7897);
nor U13853 (N_13853,N_5740,N_7848);
or U13854 (N_13854,N_9130,N_9568);
and U13855 (N_13855,N_9719,N_5560);
and U13856 (N_13856,N_9960,N_7651);
xor U13857 (N_13857,N_7682,N_6146);
xor U13858 (N_13858,N_9770,N_6975);
and U13859 (N_13859,N_7464,N_9359);
nand U13860 (N_13860,N_9410,N_7441);
or U13861 (N_13861,N_6085,N_8938);
or U13862 (N_13862,N_6578,N_9827);
or U13863 (N_13863,N_7562,N_6337);
or U13864 (N_13864,N_5408,N_7778);
and U13865 (N_13865,N_8022,N_9208);
xnor U13866 (N_13866,N_7045,N_8115);
nor U13867 (N_13867,N_8950,N_7018);
or U13868 (N_13868,N_7556,N_7325);
xnor U13869 (N_13869,N_9195,N_6934);
nand U13870 (N_13870,N_7299,N_8330);
nor U13871 (N_13871,N_8542,N_5546);
or U13872 (N_13872,N_5886,N_5985);
and U13873 (N_13873,N_7521,N_5451);
or U13874 (N_13874,N_6423,N_6222);
and U13875 (N_13875,N_5201,N_6258);
nand U13876 (N_13876,N_5543,N_5057);
or U13877 (N_13877,N_8452,N_7270);
or U13878 (N_13878,N_9569,N_9131);
nand U13879 (N_13879,N_5394,N_8251);
and U13880 (N_13880,N_5640,N_8039);
or U13881 (N_13881,N_6772,N_8128);
or U13882 (N_13882,N_8168,N_5246);
nand U13883 (N_13883,N_9392,N_8987);
and U13884 (N_13884,N_9561,N_8651);
and U13885 (N_13885,N_7045,N_6883);
nor U13886 (N_13886,N_7058,N_9493);
and U13887 (N_13887,N_8393,N_6836);
nand U13888 (N_13888,N_9456,N_8712);
or U13889 (N_13889,N_8532,N_6520);
or U13890 (N_13890,N_9954,N_9749);
xor U13891 (N_13891,N_6870,N_9427);
xnor U13892 (N_13892,N_7211,N_8929);
nor U13893 (N_13893,N_9508,N_6185);
and U13894 (N_13894,N_6288,N_5743);
nor U13895 (N_13895,N_5337,N_9413);
or U13896 (N_13896,N_8396,N_5616);
and U13897 (N_13897,N_9620,N_7455);
and U13898 (N_13898,N_6315,N_8947);
or U13899 (N_13899,N_7518,N_8687);
or U13900 (N_13900,N_8641,N_5910);
nand U13901 (N_13901,N_8430,N_9586);
nand U13902 (N_13902,N_6441,N_8719);
and U13903 (N_13903,N_9670,N_9455);
xnor U13904 (N_13904,N_9808,N_5824);
nand U13905 (N_13905,N_6469,N_5532);
nand U13906 (N_13906,N_8862,N_9865);
or U13907 (N_13907,N_7164,N_9018);
and U13908 (N_13908,N_5046,N_6630);
nand U13909 (N_13909,N_8540,N_9583);
xor U13910 (N_13910,N_8160,N_7286);
nor U13911 (N_13911,N_5282,N_7826);
xnor U13912 (N_13912,N_5779,N_9509);
and U13913 (N_13913,N_5489,N_8302);
and U13914 (N_13914,N_6652,N_9522);
or U13915 (N_13915,N_8388,N_6559);
nand U13916 (N_13916,N_6673,N_5943);
xor U13917 (N_13917,N_9669,N_7503);
and U13918 (N_13918,N_9464,N_9285);
xor U13919 (N_13919,N_7761,N_6539);
or U13920 (N_13920,N_8747,N_5066);
nor U13921 (N_13921,N_8605,N_6345);
xnor U13922 (N_13922,N_8340,N_6970);
nor U13923 (N_13923,N_9646,N_5088);
and U13924 (N_13924,N_7514,N_8255);
xor U13925 (N_13925,N_9437,N_8444);
or U13926 (N_13926,N_5972,N_9429);
and U13927 (N_13927,N_9863,N_5028);
and U13928 (N_13928,N_5188,N_9349);
nand U13929 (N_13929,N_6549,N_6594);
nor U13930 (N_13930,N_5508,N_9844);
and U13931 (N_13931,N_6866,N_5740);
xnor U13932 (N_13932,N_7629,N_8782);
or U13933 (N_13933,N_6262,N_7893);
or U13934 (N_13934,N_5127,N_6186);
nand U13935 (N_13935,N_9238,N_6054);
and U13936 (N_13936,N_9561,N_6378);
or U13937 (N_13937,N_8484,N_5220);
xnor U13938 (N_13938,N_8657,N_5236);
nand U13939 (N_13939,N_5926,N_6100);
or U13940 (N_13940,N_9153,N_8676);
nand U13941 (N_13941,N_7387,N_7647);
and U13942 (N_13942,N_9217,N_9179);
nor U13943 (N_13943,N_5436,N_6245);
or U13944 (N_13944,N_8530,N_6580);
nand U13945 (N_13945,N_6675,N_7785);
or U13946 (N_13946,N_8561,N_6387);
nor U13947 (N_13947,N_6692,N_8544);
nand U13948 (N_13948,N_8180,N_5501);
nor U13949 (N_13949,N_7692,N_7833);
nor U13950 (N_13950,N_5071,N_6848);
and U13951 (N_13951,N_8240,N_7764);
xnor U13952 (N_13952,N_8033,N_9396);
xnor U13953 (N_13953,N_9308,N_5955);
and U13954 (N_13954,N_5546,N_9708);
or U13955 (N_13955,N_6118,N_6751);
or U13956 (N_13956,N_8138,N_9015);
nand U13957 (N_13957,N_5825,N_7530);
nand U13958 (N_13958,N_9170,N_9422);
or U13959 (N_13959,N_9147,N_9808);
xor U13960 (N_13960,N_8615,N_5486);
and U13961 (N_13961,N_8499,N_5994);
xnor U13962 (N_13962,N_8213,N_9957);
nand U13963 (N_13963,N_7837,N_7897);
or U13964 (N_13964,N_7164,N_7544);
nand U13965 (N_13965,N_9109,N_6651);
or U13966 (N_13966,N_8152,N_8762);
xor U13967 (N_13967,N_6626,N_5141);
xor U13968 (N_13968,N_7626,N_9604);
or U13969 (N_13969,N_8853,N_5265);
xor U13970 (N_13970,N_5038,N_9673);
or U13971 (N_13971,N_5664,N_8607);
nand U13972 (N_13972,N_5924,N_8080);
xnor U13973 (N_13973,N_7373,N_8906);
nor U13974 (N_13974,N_9113,N_8684);
and U13975 (N_13975,N_7912,N_5794);
nand U13976 (N_13976,N_5332,N_5315);
xor U13977 (N_13977,N_8979,N_7262);
nor U13978 (N_13978,N_5736,N_5818);
nand U13979 (N_13979,N_7848,N_7093);
or U13980 (N_13980,N_8659,N_7367);
xnor U13981 (N_13981,N_7619,N_7183);
or U13982 (N_13982,N_7887,N_9123);
xor U13983 (N_13983,N_8294,N_8193);
xor U13984 (N_13984,N_7142,N_7048);
nor U13985 (N_13985,N_8763,N_8111);
or U13986 (N_13986,N_7700,N_9876);
and U13987 (N_13987,N_7584,N_6939);
xor U13988 (N_13988,N_9049,N_8785);
nand U13989 (N_13989,N_6143,N_9435);
nor U13990 (N_13990,N_5252,N_7310);
xor U13991 (N_13991,N_9127,N_6589);
xnor U13992 (N_13992,N_7486,N_8827);
xor U13993 (N_13993,N_9396,N_5393);
nor U13994 (N_13994,N_9164,N_9245);
nand U13995 (N_13995,N_6816,N_5647);
nand U13996 (N_13996,N_7273,N_6536);
or U13997 (N_13997,N_9164,N_8867);
xor U13998 (N_13998,N_7984,N_5341);
or U13999 (N_13999,N_7492,N_5223);
or U14000 (N_14000,N_8376,N_7024);
nor U14001 (N_14001,N_8205,N_8133);
xnor U14002 (N_14002,N_8116,N_7492);
nor U14003 (N_14003,N_8753,N_5365);
and U14004 (N_14004,N_7611,N_8082);
xor U14005 (N_14005,N_5557,N_5463);
nor U14006 (N_14006,N_7581,N_9245);
nand U14007 (N_14007,N_9104,N_5171);
xor U14008 (N_14008,N_5090,N_9434);
or U14009 (N_14009,N_8238,N_8724);
or U14010 (N_14010,N_6268,N_6441);
nand U14011 (N_14011,N_7805,N_8477);
nor U14012 (N_14012,N_7631,N_5431);
and U14013 (N_14013,N_5375,N_7367);
nand U14014 (N_14014,N_9822,N_6698);
xnor U14015 (N_14015,N_5037,N_9850);
xor U14016 (N_14016,N_6603,N_7200);
nand U14017 (N_14017,N_7531,N_8259);
xnor U14018 (N_14018,N_6761,N_8022);
nor U14019 (N_14019,N_5500,N_7876);
nor U14020 (N_14020,N_6706,N_6000);
or U14021 (N_14021,N_8816,N_9231);
or U14022 (N_14022,N_5587,N_8414);
xor U14023 (N_14023,N_7632,N_7184);
nand U14024 (N_14024,N_5972,N_7807);
xnor U14025 (N_14025,N_5095,N_5433);
and U14026 (N_14026,N_5890,N_5611);
nor U14027 (N_14027,N_7239,N_6657);
nor U14028 (N_14028,N_6233,N_9014);
and U14029 (N_14029,N_9701,N_9641);
or U14030 (N_14030,N_9090,N_7814);
or U14031 (N_14031,N_9090,N_5949);
or U14032 (N_14032,N_7167,N_9946);
xnor U14033 (N_14033,N_9387,N_7785);
xor U14034 (N_14034,N_5170,N_8033);
xnor U14035 (N_14035,N_7081,N_9019);
and U14036 (N_14036,N_6955,N_8586);
xnor U14037 (N_14037,N_7255,N_8645);
or U14038 (N_14038,N_7819,N_9572);
nor U14039 (N_14039,N_6715,N_7758);
nand U14040 (N_14040,N_9455,N_9954);
xnor U14041 (N_14041,N_5722,N_8457);
or U14042 (N_14042,N_8516,N_5899);
or U14043 (N_14043,N_9305,N_7227);
nand U14044 (N_14044,N_9598,N_7901);
nor U14045 (N_14045,N_8799,N_8350);
or U14046 (N_14046,N_9449,N_6748);
or U14047 (N_14047,N_9264,N_6500);
nand U14048 (N_14048,N_5029,N_7216);
xnor U14049 (N_14049,N_8724,N_6421);
xnor U14050 (N_14050,N_5206,N_8974);
and U14051 (N_14051,N_9807,N_9766);
and U14052 (N_14052,N_6211,N_6767);
and U14053 (N_14053,N_9304,N_8946);
and U14054 (N_14054,N_8912,N_6207);
nand U14055 (N_14055,N_7297,N_6310);
nand U14056 (N_14056,N_5981,N_6527);
xor U14057 (N_14057,N_8055,N_9652);
or U14058 (N_14058,N_8390,N_7452);
or U14059 (N_14059,N_5232,N_5506);
or U14060 (N_14060,N_9387,N_7446);
nor U14061 (N_14061,N_6626,N_9640);
nand U14062 (N_14062,N_7117,N_5687);
or U14063 (N_14063,N_5325,N_8734);
and U14064 (N_14064,N_8894,N_9496);
xor U14065 (N_14065,N_6039,N_6529);
and U14066 (N_14066,N_6312,N_5058);
and U14067 (N_14067,N_8582,N_9204);
or U14068 (N_14068,N_9826,N_6052);
or U14069 (N_14069,N_9414,N_7629);
and U14070 (N_14070,N_9043,N_8785);
or U14071 (N_14071,N_9790,N_6655);
nor U14072 (N_14072,N_8753,N_9323);
and U14073 (N_14073,N_6058,N_8475);
nand U14074 (N_14074,N_5942,N_6472);
nand U14075 (N_14075,N_9045,N_9177);
or U14076 (N_14076,N_9892,N_7643);
or U14077 (N_14077,N_6925,N_7259);
nand U14078 (N_14078,N_8241,N_5309);
xnor U14079 (N_14079,N_7912,N_7692);
nand U14080 (N_14080,N_8425,N_9077);
nand U14081 (N_14081,N_7691,N_7627);
and U14082 (N_14082,N_5355,N_5635);
nor U14083 (N_14083,N_7227,N_8633);
and U14084 (N_14084,N_7416,N_7857);
nor U14085 (N_14085,N_5405,N_5029);
or U14086 (N_14086,N_8584,N_8145);
nand U14087 (N_14087,N_6242,N_7711);
and U14088 (N_14088,N_8338,N_7572);
nor U14089 (N_14089,N_5856,N_7196);
nand U14090 (N_14090,N_5336,N_8836);
or U14091 (N_14091,N_6494,N_9579);
xnor U14092 (N_14092,N_8561,N_8609);
or U14093 (N_14093,N_7710,N_9921);
or U14094 (N_14094,N_9310,N_6922);
xnor U14095 (N_14095,N_9793,N_7687);
nand U14096 (N_14096,N_7832,N_5752);
nor U14097 (N_14097,N_7476,N_5946);
and U14098 (N_14098,N_9738,N_6705);
and U14099 (N_14099,N_9103,N_8014);
and U14100 (N_14100,N_8166,N_9116);
xnor U14101 (N_14101,N_6046,N_6165);
or U14102 (N_14102,N_8790,N_6429);
xnor U14103 (N_14103,N_8885,N_9584);
and U14104 (N_14104,N_9513,N_9735);
xor U14105 (N_14105,N_7909,N_7068);
nor U14106 (N_14106,N_7473,N_7149);
xor U14107 (N_14107,N_6256,N_7848);
nor U14108 (N_14108,N_5148,N_7950);
or U14109 (N_14109,N_6866,N_9430);
xnor U14110 (N_14110,N_9687,N_6760);
or U14111 (N_14111,N_9096,N_9052);
or U14112 (N_14112,N_7630,N_6394);
nand U14113 (N_14113,N_7441,N_7609);
nor U14114 (N_14114,N_5277,N_5888);
nor U14115 (N_14115,N_5883,N_7455);
nor U14116 (N_14116,N_7623,N_8642);
or U14117 (N_14117,N_7903,N_9054);
xnor U14118 (N_14118,N_5423,N_7291);
xnor U14119 (N_14119,N_6404,N_9767);
nand U14120 (N_14120,N_6882,N_8458);
nor U14121 (N_14121,N_7573,N_6319);
or U14122 (N_14122,N_5805,N_5445);
nand U14123 (N_14123,N_5852,N_8721);
or U14124 (N_14124,N_6312,N_9307);
nor U14125 (N_14125,N_5951,N_8378);
xnor U14126 (N_14126,N_7582,N_7935);
nand U14127 (N_14127,N_5728,N_5554);
nand U14128 (N_14128,N_5247,N_9697);
xnor U14129 (N_14129,N_9626,N_8558);
nor U14130 (N_14130,N_8248,N_8512);
xnor U14131 (N_14131,N_8719,N_8226);
nand U14132 (N_14132,N_5794,N_7335);
or U14133 (N_14133,N_5129,N_5735);
or U14134 (N_14134,N_7151,N_6976);
nor U14135 (N_14135,N_5463,N_7314);
or U14136 (N_14136,N_9339,N_5760);
and U14137 (N_14137,N_8843,N_5783);
or U14138 (N_14138,N_7382,N_6826);
xor U14139 (N_14139,N_9302,N_7331);
or U14140 (N_14140,N_8362,N_5573);
or U14141 (N_14141,N_9014,N_8829);
and U14142 (N_14142,N_5104,N_6913);
and U14143 (N_14143,N_6785,N_8245);
xnor U14144 (N_14144,N_8314,N_7719);
nand U14145 (N_14145,N_6283,N_8327);
and U14146 (N_14146,N_8047,N_9708);
and U14147 (N_14147,N_6359,N_9812);
xor U14148 (N_14148,N_8951,N_9646);
nor U14149 (N_14149,N_5711,N_5747);
nor U14150 (N_14150,N_8418,N_5483);
and U14151 (N_14151,N_7809,N_6275);
and U14152 (N_14152,N_7475,N_9740);
nor U14153 (N_14153,N_8055,N_6678);
xor U14154 (N_14154,N_5669,N_9051);
nand U14155 (N_14155,N_5556,N_8593);
nor U14156 (N_14156,N_9987,N_5123);
or U14157 (N_14157,N_6844,N_7415);
and U14158 (N_14158,N_5327,N_9344);
nor U14159 (N_14159,N_7026,N_8845);
xor U14160 (N_14160,N_5601,N_6540);
nor U14161 (N_14161,N_9885,N_5303);
nand U14162 (N_14162,N_7513,N_6049);
nand U14163 (N_14163,N_8665,N_6837);
nor U14164 (N_14164,N_7269,N_6635);
nor U14165 (N_14165,N_6127,N_7156);
or U14166 (N_14166,N_7646,N_7559);
nand U14167 (N_14167,N_8079,N_9914);
xnor U14168 (N_14168,N_5774,N_9965);
nand U14169 (N_14169,N_8814,N_8715);
nor U14170 (N_14170,N_6487,N_7208);
and U14171 (N_14171,N_9157,N_5650);
nand U14172 (N_14172,N_5951,N_9532);
nor U14173 (N_14173,N_9237,N_6812);
xor U14174 (N_14174,N_8179,N_7399);
nand U14175 (N_14175,N_7453,N_6099);
nand U14176 (N_14176,N_9132,N_7608);
nand U14177 (N_14177,N_6997,N_5001);
nor U14178 (N_14178,N_5845,N_9659);
xnor U14179 (N_14179,N_8029,N_5410);
xor U14180 (N_14180,N_8836,N_7993);
nand U14181 (N_14181,N_5507,N_6721);
nor U14182 (N_14182,N_6356,N_6721);
nand U14183 (N_14183,N_9796,N_7973);
nand U14184 (N_14184,N_8274,N_6577);
and U14185 (N_14185,N_8043,N_7499);
nand U14186 (N_14186,N_8056,N_6510);
nand U14187 (N_14187,N_5369,N_5149);
or U14188 (N_14188,N_6876,N_9625);
nand U14189 (N_14189,N_7589,N_7624);
nand U14190 (N_14190,N_6133,N_5997);
and U14191 (N_14191,N_9776,N_6701);
xnor U14192 (N_14192,N_5563,N_8909);
nand U14193 (N_14193,N_8453,N_8092);
xnor U14194 (N_14194,N_7440,N_9868);
xnor U14195 (N_14195,N_6040,N_7353);
xor U14196 (N_14196,N_5823,N_5528);
or U14197 (N_14197,N_7989,N_6904);
or U14198 (N_14198,N_8712,N_8236);
xor U14199 (N_14199,N_7957,N_8004);
and U14200 (N_14200,N_7328,N_6564);
nor U14201 (N_14201,N_9741,N_5077);
nor U14202 (N_14202,N_5875,N_5624);
xnor U14203 (N_14203,N_6450,N_7029);
and U14204 (N_14204,N_5892,N_6151);
nand U14205 (N_14205,N_6443,N_9637);
nor U14206 (N_14206,N_6423,N_6025);
nand U14207 (N_14207,N_5465,N_9370);
xor U14208 (N_14208,N_5104,N_8006);
and U14209 (N_14209,N_8086,N_5192);
and U14210 (N_14210,N_9921,N_7771);
and U14211 (N_14211,N_6791,N_6053);
nand U14212 (N_14212,N_6885,N_8814);
or U14213 (N_14213,N_5178,N_7761);
nand U14214 (N_14214,N_7063,N_6321);
and U14215 (N_14215,N_6117,N_6749);
and U14216 (N_14216,N_7215,N_9008);
xnor U14217 (N_14217,N_7557,N_9129);
nand U14218 (N_14218,N_5000,N_9450);
nand U14219 (N_14219,N_9302,N_9628);
or U14220 (N_14220,N_9910,N_7314);
and U14221 (N_14221,N_9660,N_6186);
and U14222 (N_14222,N_6110,N_9032);
and U14223 (N_14223,N_5021,N_8880);
nor U14224 (N_14224,N_5585,N_5794);
nand U14225 (N_14225,N_6207,N_8655);
nor U14226 (N_14226,N_9326,N_5680);
xnor U14227 (N_14227,N_7253,N_7682);
and U14228 (N_14228,N_7217,N_9806);
or U14229 (N_14229,N_9852,N_5547);
nand U14230 (N_14230,N_8616,N_9707);
nand U14231 (N_14231,N_8073,N_6660);
xor U14232 (N_14232,N_9433,N_5191);
and U14233 (N_14233,N_9757,N_6807);
nor U14234 (N_14234,N_5764,N_9369);
or U14235 (N_14235,N_5670,N_5875);
nor U14236 (N_14236,N_9352,N_6796);
nor U14237 (N_14237,N_8897,N_9354);
and U14238 (N_14238,N_5069,N_6415);
xor U14239 (N_14239,N_8375,N_5384);
and U14240 (N_14240,N_9665,N_9230);
and U14241 (N_14241,N_9403,N_8761);
xor U14242 (N_14242,N_5409,N_6254);
xor U14243 (N_14243,N_7879,N_9648);
or U14244 (N_14244,N_8170,N_8216);
nand U14245 (N_14245,N_8855,N_9893);
and U14246 (N_14246,N_5701,N_5752);
or U14247 (N_14247,N_5116,N_7955);
xor U14248 (N_14248,N_6558,N_7843);
and U14249 (N_14249,N_7777,N_5174);
or U14250 (N_14250,N_9545,N_9439);
nand U14251 (N_14251,N_7384,N_8173);
nand U14252 (N_14252,N_6432,N_9144);
or U14253 (N_14253,N_5860,N_6140);
and U14254 (N_14254,N_5029,N_9956);
xor U14255 (N_14255,N_5807,N_9940);
nor U14256 (N_14256,N_7168,N_9297);
and U14257 (N_14257,N_5359,N_9898);
and U14258 (N_14258,N_5633,N_6598);
xnor U14259 (N_14259,N_5057,N_5090);
nor U14260 (N_14260,N_7943,N_8453);
nor U14261 (N_14261,N_8690,N_7923);
nand U14262 (N_14262,N_8000,N_7196);
nand U14263 (N_14263,N_9524,N_8063);
and U14264 (N_14264,N_9270,N_5996);
nand U14265 (N_14265,N_7008,N_9241);
and U14266 (N_14266,N_7779,N_6148);
nor U14267 (N_14267,N_9613,N_5368);
or U14268 (N_14268,N_9369,N_6760);
nor U14269 (N_14269,N_7838,N_7129);
and U14270 (N_14270,N_8458,N_5605);
nor U14271 (N_14271,N_8070,N_7313);
xnor U14272 (N_14272,N_7845,N_8108);
xnor U14273 (N_14273,N_8580,N_7271);
and U14274 (N_14274,N_5323,N_9922);
xor U14275 (N_14275,N_9903,N_8360);
xnor U14276 (N_14276,N_9966,N_8820);
nand U14277 (N_14277,N_7474,N_5597);
and U14278 (N_14278,N_6558,N_7239);
and U14279 (N_14279,N_7933,N_5421);
xor U14280 (N_14280,N_5518,N_6479);
nor U14281 (N_14281,N_7097,N_6993);
nand U14282 (N_14282,N_6698,N_7340);
nor U14283 (N_14283,N_5090,N_9444);
or U14284 (N_14284,N_7985,N_9884);
or U14285 (N_14285,N_5572,N_8856);
or U14286 (N_14286,N_5092,N_5213);
nand U14287 (N_14287,N_5506,N_8192);
xor U14288 (N_14288,N_8356,N_9877);
nor U14289 (N_14289,N_9077,N_5938);
or U14290 (N_14290,N_5057,N_7424);
and U14291 (N_14291,N_7549,N_6222);
xor U14292 (N_14292,N_6089,N_7135);
nor U14293 (N_14293,N_6927,N_9371);
and U14294 (N_14294,N_6299,N_8326);
and U14295 (N_14295,N_8935,N_7135);
or U14296 (N_14296,N_7239,N_7021);
xnor U14297 (N_14297,N_9533,N_9475);
nand U14298 (N_14298,N_6843,N_6122);
xnor U14299 (N_14299,N_6478,N_8186);
xnor U14300 (N_14300,N_5292,N_5873);
and U14301 (N_14301,N_6283,N_8733);
nand U14302 (N_14302,N_7759,N_7984);
and U14303 (N_14303,N_8651,N_7419);
xor U14304 (N_14304,N_8394,N_7759);
and U14305 (N_14305,N_5632,N_5199);
xor U14306 (N_14306,N_6383,N_8960);
or U14307 (N_14307,N_6913,N_8245);
nand U14308 (N_14308,N_8810,N_7573);
nor U14309 (N_14309,N_5839,N_9282);
or U14310 (N_14310,N_5258,N_7840);
nor U14311 (N_14311,N_9224,N_7419);
and U14312 (N_14312,N_8400,N_6190);
and U14313 (N_14313,N_5405,N_8238);
xnor U14314 (N_14314,N_6744,N_7299);
nor U14315 (N_14315,N_7424,N_6911);
nor U14316 (N_14316,N_9424,N_5521);
xor U14317 (N_14317,N_6101,N_5272);
xnor U14318 (N_14318,N_7842,N_8872);
xor U14319 (N_14319,N_7110,N_7765);
nor U14320 (N_14320,N_7259,N_5605);
and U14321 (N_14321,N_5389,N_8350);
and U14322 (N_14322,N_8500,N_9990);
or U14323 (N_14323,N_9389,N_6368);
and U14324 (N_14324,N_6167,N_5073);
xnor U14325 (N_14325,N_7633,N_9907);
and U14326 (N_14326,N_9173,N_8709);
nor U14327 (N_14327,N_5047,N_9278);
or U14328 (N_14328,N_8752,N_7520);
and U14329 (N_14329,N_9476,N_8097);
xor U14330 (N_14330,N_9502,N_5614);
xor U14331 (N_14331,N_6831,N_9372);
nand U14332 (N_14332,N_9944,N_9663);
xnor U14333 (N_14333,N_8352,N_5341);
xnor U14334 (N_14334,N_9013,N_8053);
nor U14335 (N_14335,N_6470,N_9236);
nor U14336 (N_14336,N_7804,N_5758);
and U14337 (N_14337,N_6083,N_8638);
xor U14338 (N_14338,N_7131,N_7639);
nand U14339 (N_14339,N_6836,N_5886);
xnor U14340 (N_14340,N_8122,N_5109);
xnor U14341 (N_14341,N_6698,N_8390);
or U14342 (N_14342,N_5573,N_8305);
nand U14343 (N_14343,N_7035,N_6789);
nand U14344 (N_14344,N_6930,N_8797);
xor U14345 (N_14345,N_7283,N_8751);
nand U14346 (N_14346,N_6779,N_6008);
and U14347 (N_14347,N_8332,N_7158);
xnor U14348 (N_14348,N_8441,N_8848);
xnor U14349 (N_14349,N_6218,N_6530);
or U14350 (N_14350,N_9654,N_7930);
and U14351 (N_14351,N_8830,N_7336);
or U14352 (N_14352,N_8969,N_9825);
or U14353 (N_14353,N_6503,N_7658);
xor U14354 (N_14354,N_8938,N_9979);
and U14355 (N_14355,N_8635,N_5506);
and U14356 (N_14356,N_7878,N_6921);
nand U14357 (N_14357,N_8688,N_7227);
xor U14358 (N_14358,N_5835,N_7453);
or U14359 (N_14359,N_8925,N_7546);
nor U14360 (N_14360,N_9610,N_8107);
nor U14361 (N_14361,N_8104,N_6186);
nor U14362 (N_14362,N_8654,N_9459);
or U14363 (N_14363,N_7755,N_5414);
and U14364 (N_14364,N_6315,N_6209);
and U14365 (N_14365,N_5011,N_8772);
xnor U14366 (N_14366,N_9688,N_8396);
or U14367 (N_14367,N_5114,N_7170);
nand U14368 (N_14368,N_9292,N_8140);
and U14369 (N_14369,N_5074,N_9528);
or U14370 (N_14370,N_6737,N_9131);
xnor U14371 (N_14371,N_7518,N_9339);
and U14372 (N_14372,N_7049,N_9070);
nor U14373 (N_14373,N_9764,N_5051);
or U14374 (N_14374,N_7738,N_7130);
nor U14375 (N_14375,N_6291,N_5946);
nand U14376 (N_14376,N_7162,N_5161);
or U14377 (N_14377,N_8997,N_5155);
nand U14378 (N_14378,N_8120,N_8753);
or U14379 (N_14379,N_7471,N_7289);
nand U14380 (N_14380,N_7905,N_6866);
nand U14381 (N_14381,N_9069,N_5169);
nor U14382 (N_14382,N_8970,N_6079);
and U14383 (N_14383,N_6268,N_7588);
nand U14384 (N_14384,N_7013,N_7526);
nor U14385 (N_14385,N_6444,N_9578);
nand U14386 (N_14386,N_5136,N_7421);
xor U14387 (N_14387,N_6080,N_9102);
nor U14388 (N_14388,N_5372,N_7834);
nand U14389 (N_14389,N_7217,N_6917);
and U14390 (N_14390,N_9167,N_5753);
or U14391 (N_14391,N_8722,N_9160);
and U14392 (N_14392,N_5512,N_8313);
and U14393 (N_14393,N_5971,N_8943);
or U14394 (N_14394,N_6146,N_7322);
nor U14395 (N_14395,N_7793,N_9448);
and U14396 (N_14396,N_9266,N_8449);
or U14397 (N_14397,N_5987,N_9698);
nand U14398 (N_14398,N_5894,N_7932);
and U14399 (N_14399,N_8371,N_9332);
and U14400 (N_14400,N_6183,N_7323);
xnor U14401 (N_14401,N_9176,N_7811);
or U14402 (N_14402,N_9478,N_9598);
and U14403 (N_14403,N_8560,N_6355);
or U14404 (N_14404,N_7189,N_6439);
nand U14405 (N_14405,N_8630,N_5792);
or U14406 (N_14406,N_6949,N_8833);
nor U14407 (N_14407,N_9600,N_5029);
or U14408 (N_14408,N_7227,N_5776);
nand U14409 (N_14409,N_7955,N_8852);
and U14410 (N_14410,N_7498,N_6479);
and U14411 (N_14411,N_6791,N_9034);
or U14412 (N_14412,N_7190,N_7372);
nand U14413 (N_14413,N_7044,N_9291);
nor U14414 (N_14414,N_5602,N_5450);
nor U14415 (N_14415,N_8130,N_5750);
nor U14416 (N_14416,N_9859,N_6879);
nand U14417 (N_14417,N_5451,N_9077);
xnor U14418 (N_14418,N_9239,N_7147);
and U14419 (N_14419,N_6635,N_6715);
or U14420 (N_14420,N_5223,N_8941);
nor U14421 (N_14421,N_5015,N_6467);
xnor U14422 (N_14422,N_5652,N_5774);
nand U14423 (N_14423,N_7871,N_6654);
xor U14424 (N_14424,N_7395,N_6556);
or U14425 (N_14425,N_8259,N_7629);
or U14426 (N_14426,N_9271,N_6379);
nand U14427 (N_14427,N_5202,N_8587);
or U14428 (N_14428,N_8751,N_6046);
nand U14429 (N_14429,N_8548,N_7016);
xnor U14430 (N_14430,N_7844,N_5957);
xor U14431 (N_14431,N_6558,N_9080);
xor U14432 (N_14432,N_6988,N_9888);
nand U14433 (N_14433,N_5700,N_8404);
nand U14434 (N_14434,N_7033,N_6254);
nor U14435 (N_14435,N_9803,N_7909);
and U14436 (N_14436,N_7034,N_9498);
or U14437 (N_14437,N_8495,N_8914);
or U14438 (N_14438,N_8186,N_8347);
or U14439 (N_14439,N_6833,N_7288);
xor U14440 (N_14440,N_9153,N_5305);
nand U14441 (N_14441,N_8865,N_8707);
nor U14442 (N_14442,N_6111,N_7603);
and U14443 (N_14443,N_7579,N_6428);
and U14444 (N_14444,N_7058,N_9518);
nor U14445 (N_14445,N_7688,N_9136);
nand U14446 (N_14446,N_6212,N_7070);
or U14447 (N_14447,N_9209,N_7779);
and U14448 (N_14448,N_7090,N_7759);
xor U14449 (N_14449,N_9340,N_5196);
nand U14450 (N_14450,N_6359,N_7998);
nand U14451 (N_14451,N_7995,N_5049);
nand U14452 (N_14452,N_9998,N_6841);
and U14453 (N_14453,N_8799,N_8542);
or U14454 (N_14454,N_7450,N_8650);
or U14455 (N_14455,N_9674,N_9716);
nor U14456 (N_14456,N_6776,N_5860);
nand U14457 (N_14457,N_6691,N_6208);
nand U14458 (N_14458,N_5352,N_5635);
and U14459 (N_14459,N_7512,N_6793);
xnor U14460 (N_14460,N_8643,N_8818);
nand U14461 (N_14461,N_5914,N_6830);
xor U14462 (N_14462,N_9062,N_7564);
nand U14463 (N_14463,N_5632,N_5451);
xor U14464 (N_14464,N_9859,N_7767);
nor U14465 (N_14465,N_5629,N_5287);
nor U14466 (N_14466,N_8874,N_8983);
xnor U14467 (N_14467,N_8669,N_8691);
xor U14468 (N_14468,N_5773,N_5888);
xnor U14469 (N_14469,N_9658,N_6613);
and U14470 (N_14470,N_8658,N_8265);
nand U14471 (N_14471,N_5730,N_6269);
or U14472 (N_14472,N_5504,N_9303);
and U14473 (N_14473,N_6415,N_7050);
or U14474 (N_14474,N_7653,N_7387);
or U14475 (N_14475,N_5659,N_7162);
xnor U14476 (N_14476,N_5351,N_5092);
nand U14477 (N_14477,N_6992,N_8627);
and U14478 (N_14478,N_8853,N_9764);
nor U14479 (N_14479,N_5019,N_8798);
nand U14480 (N_14480,N_8915,N_9968);
nor U14481 (N_14481,N_9916,N_6143);
xnor U14482 (N_14482,N_9917,N_8027);
or U14483 (N_14483,N_9147,N_6925);
nor U14484 (N_14484,N_6319,N_6079);
nor U14485 (N_14485,N_7754,N_7877);
and U14486 (N_14486,N_8161,N_6909);
nor U14487 (N_14487,N_9336,N_7978);
nor U14488 (N_14488,N_8860,N_6387);
and U14489 (N_14489,N_6512,N_6197);
nand U14490 (N_14490,N_6966,N_6257);
or U14491 (N_14491,N_7044,N_6013);
or U14492 (N_14492,N_6936,N_7732);
and U14493 (N_14493,N_5734,N_6141);
nor U14494 (N_14494,N_5882,N_9604);
and U14495 (N_14495,N_5246,N_9736);
and U14496 (N_14496,N_9426,N_6433);
nand U14497 (N_14497,N_9808,N_9836);
or U14498 (N_14498,N_8694,N_7053);
or U14499 (N_14499,N_5660,N_6284);
nor U14500 (N_14500,N_7895,N_8292);
and U14501 (N_14501,N_8479,N_9545);
xor U14502 (N_14502,N_7136,N_5099);
and U14503 (N_14503,N_8802,N_6925);
nand U14504 (N_14504,N_5497,N_5956);
xor U14505 (N_14505,N_6798,N_8677);
nor U14506 (N_14506,N_6257,N_9852);
nand U14507 (N_14507,N_7281,N_7875);
xnor U14508 (N_14508,N_5461,N_6228);
xor U14509 (N_14509,N_6261,N_5517);
nand U14510 (N_14510,N_7665,N_5042);
or U14511 (N_14511,N_5025,N_7586);
and U14512 (N_14512,N_8622,N_7121);
xnor U14513 (N_14513,N_5669,N_6717);
nand U14514 (N_14514,N_8020,N_6081);
xor U14515 (N_14515,N_9344,N_8757);
nand U14516 (N_14516,N_8309,N_9535);
or U14517 (N_14517,N_5666,N_6966);
xnor U14518 (N_14518,N_6861,N_6581);
nor U14519 (N_14519,N_9165,N_5980);
or U14520 (N_14520,N_6938,N_7102);
nand U14521 (N_14521,N_5420,N_8684);
nor U14522 (N_14522,N_7503,N_6190);
xnor U14523 (N_14523,N_9857,N_9514);
nand U14524 (N_14524,N_5681,N_9761);
nor U14525 (N_14525,N_7585,N_9333);
nand U14526 (N_14526,N_5296,N_5064);
nor U14527 (N_14527,N_7586,N_5559);
xnor U14528 (N_14528,N_6425,N_9652);
and U14529 (N_14529,N_6995,N_5113);
xnor U14530 (N_14530,N_9196,N_8579);
and U14531 (N_14531,N_5884,N_8960);
nor U14532 (N_14532,N_7223,N_8906);
nand U14533 (N_14533,N_6575,N_7431);
nor U14534 (N_14534,N_6787,N_5987);
xor U14535 (N_14535,N_6672,N_6075);
nand U14536 (N_14536,N_7160,N_9161);
or U14537 (N_14537,N_7534,N_9560);
nand U14538 (N_14538,N_8416,N_8078);
xnor U14539 (N_14539,N_5550,N_9132);
nor U14540 (N_14540,N_7403,N_8709);
or U14541 (N_14541,N_9471,N_9586);
xnor U14542 (N_14542,N_9242,N_5910);
or U14543 (N_14543,N_6798,N_9323);
xnor U14544 (N_14544,N_9030,N_9748);
xor U14545 (N_14545,N_9905,N_5295);
nand U14546 (N_14546,N_8010,N_8050);
nor U14547 (N_14547,N_9487,N_6011);
or U14548 (N_14548,N_7492,N_8211);
and U14549 (N_14549,N_8123,N_5269);
xnor U14550 (N_14550,N_6117,N_8895);
or U14551 (N_14551,N_5682,N_8829);
nor U14552 (N_14552,N_9778,N_5747);
or U14553 (N_14553,N_5970,N_9736);
or U14554 (N_14554,N_6734,N_5827);
or U14555 (N_14555,N_7148,N_6604);
xnor U14556 (N_14556,N_5756,N_8781);
nand U14557 (N_14557,N_8167,N_8352);
or U14558 (N_14558,N_7172,N_7795);
xnor U14559 (N_14559,N_8963,N_8624);
nor U14560 (N_14560,N_5131,N_6062);
or U14561 (N_14561,N_8556,N_9210);
nand U14562 (N_14562,N_9865,N_7835);
xnor U14563 (N_14563,N_5025,N_5542);
xnor U14564 (N_14564,N_8256,N_9864);
or U14565 (N_14565,N_5904,N_5031);
and U14566 (N_14566,N_8152,N_7988);
xnor U14567 (N_14567,N_6820,N_7280);
nand U14568 (N_14568,N_6553,N_5472);
and U14569 (N_14569,N_9730,N_9253);
nand U14570 (N_14570,N_5352,N_9164);
or U14571 (N_14571,N_9576,N_5924);
nor U14572 (N_14572,N_9935,N_5004);
and U14573 (N_14573,N_9976,N_6248);
or U14574 (N_14574,N_9386,N_7914);
nand U14575 (N_14575,N_6803,N_5996);
and U14576 (N_14576,N_6628,N_5351);
xor U14577 (N_14577,N_9497,N_8698);
or U14578 (N_14578,N_5561,N_5470);
nor U14579 (N_14579,N_8070,N_6499);
xnor U14580 (N_14580,N_5931,N_6541);
nor U14581 (N_14581,N_9598,N_9117);
xnor U14582 (N_14582,N_9692,N_7638);
and U14583 (N_14583,N_8878,N_8176);
nor U14584 (N_14584,N_7648,N_7678);
nor U14585 (N_14585,N_8744,N_6023);
and U14586 (N_14586,N_7117,N_6426);
nor U14587 (N_14587,N_9235,N_5056);
nand U14588 (N_14588,N_9043,N_7291);
nand U14589 (N_14589,N_5095,N_6448);
or U14590 (N_14590,N_9922,N_8348);
nor U14591 (N_14591,N_8721,N_9050);
xor U14592 (N_14592,N_6986,N_8385);
and U14593 (N_14593,N_6534,N_7974);
xnor U14594 (N_14594,N_9112,N_7111);
nor U14595 (N_14595,N_6282,N_9053);
nor U14596 (N_14596,N_5423,N_8748);
or U14597 (N_14597,N_5131,N_7373);
and U14598 (N_14598,N_9073,N_8849);
nand U14599 (N_14599,N_8521,N_5905);
or U14600 (N_14600,N_8699,N_8849);
nand U14601 (N_14601,N_6186,N_8833);
nor U14602 (N_14602,N_5751,N_7087);
nand U14603 (N_14603,N_8060,N_6064);
or U14604 (N_14604,N_6144,N_5396);
and U14605 (N_14605,N_9679,N_9290);
nor U14606 (N_14606,N_9921,N_7466);
or U14607 (N_14607,N_9764,N_9625);
and U14608 (N_14608,N_6937,N_8059);
or U14609 (N_14609,N_7160,N_9734);
xnor U14610 (N_14610,N_6285,N_7624);
or U14611 (N_14611,N_9955,N_6101);
and U14612 (N_14612,N_9353,N_8084);
nor U14613 (N_14613,N_7899,N_5023);
or U14614 (N_14614,N_6077,N_7284);
and U14615 (N_14615,N_9472,N_8649);
or U14616 (N_14616,N_9696,N_7271);
nand U14617 (N_14617,N_5183,N_5085);
xor U14618 (N_14618,N_9457,N_5644);
xor U14619 (N_14619,N_5224,N_6869);
xor U14620 (N_14620,N_7883,N_9515);
nand U14621 (N_14621,N_5951,N_7002);
xnor U14622 (N_14622,N_6388,N_9041);
nand U14623 (N_14623,N_8519,N_5607);
or U14624 (N_14624,N_8236,N_7342);
nor U14625 (N_14625,N_9418,N_7391);
xnor U14626 (N_14626,N_5289,N_6782);
nand U14627 (N_14627,N_5587,N_9497);
and U14628 (N_14628,N_5424,N_6355);
nand U14629 (N_14629,N_5673,N_7165);
and U14630 (N_14630,N_8637,N_5371);
or U14631 (N_14631,N_8365,N_5989);
and U14632 (N_14632,N_5976,N_5497);
and U14633 (N_14633,N_9985,N_9624);
or U14634 (N_14634,N_7997,N_7657);
nand U14635 (N_14635,N_5075,N_9652);
xnor U14636 (N_14636,N_9985,N_9242);
nor U14637 (N_14637,N_7619,N_6583);
nor U14638 (N_14638,N_7383,N_5804);
and U14639 (N_14639,N_9660,N_8376);
nand U14640 (N_14640,N_6735,N_9141);
and U14641 (N_14641,N_5879,N_6571);
xor U14642 (N_14642,N_5841,N_7445);
xor U14643 (N_14643,N_7736,N_6299);
or U14644 (N_14644,N_9652,N_5329);
nand U14645 (N_14645,N_8231,N_9064);
nand U14646 (N_14646,N_9917,N_9265);
nand U14647 (N_14647,N_9921,N_6886);
xnor U14648 (N_14648,N_6598,N_7911);
or U14649 (N_14649,N_5794,N_5922);
nand U14650 (N_14650,N_9633,N_6532);
nor U14651 (N_14651,N_5907,N_5244);
or U14652 (N_14652,N_9120,N_6528);
and U14653 (N_14653,N_7114,N_8942);
nor U14654 (N_14654,N_7997,N_6327);
nand U14655 (N_14655,N_9230,N_9827);
nor U14656 (N_14656,N_6105,N_6548);
or U14657 (N_14657,N_5918,N_6890);
xor U14658 (N_14658,N_8546,N_9945);
xor U14659 (N_14659,N_6246,N_8700);
nand U14660 (N_14660,N_9300,N_7058);
or U14661 (N_14661,N_7465,N_7871);
and U14662 (N_14662,N_9635,N_7148);
or U14663 (N_14663,N_8243,N_5184);
or U14664 (N_14664,N_9876,N_7328);
nor U14665 (N_14665,N_6894,N_5541);
nand U14666 (N_14666,N_6872,N_5431);
or U14667 (N_14667,N_7239,N_6123);
nand U14668 (N_14668,N_5535,N_5071);
and U14669 (N_14669,N_5857,N_8697);
and U14670 (N_14670,N_5531,N_6536);
nor U14671 (N_14671,N_6325,N_6366);
nand U14672 (N_14672,N_8517,N_8341);
or U14673 (N_14673,N_5227,N_8637);
nor U14674 (N_14674,N_9878,N_8244);
nand U14675 (N_14675,N_6139,N_5093);
nor U14676 (N_14676,N_8540,N_5034);
xnor U14677 (N_14677,N_5891,N_7448);
nand U14678 (N_14678,N_7568,N_8642);
nand U14679 (N_14679,N_6897,N_9894);
or U14680 (N_14680,N_7322,N_6429);
or U14681 (N_14681,N_6412,N_8192);
xor U14682 (N_14682,N_9588,N_8781);
nand U14683 (N_14683,N_6523,N_7521);
nor U14684 (N_14684,N_5796,N_9962);
xnor U14685 (N_14685,N_8494,N_5763);
or U14686 (N_14686,N_8575,N_6930);
xnor U14687 (N_14687,N_8312,N_7205);
or U14688 (N_14688,N_6843,N_5268);
nor U14689 (N_14689,N_9116,N_7903);
or U14690 (N_14690,N_6777,N_5489);
xor U14691 (N_14691,N_5742,N_7991);
or U14692 (N_14692,N_6822,N_5602);
nand U14693 (N_14693,N_7960,N_8624);
nand U14694 (N_14694,N_8112,N_7919);
xnor U14695 (N_14695,N_6242,N_5654);
and U14696 (N_14696,N_9162,N_8351);
nand U14697 (N_14697,N_8423,N_6489);
xor U14698 (N_14698,N_6416,N_7892);
or U14699 (N_14699,N_8444,N_7666);
nor U14700 (N_14700,N_6177,N_5153);
or U14701 (N_14701,N_5988,N_5608);
xor U14702 (N_14702,N_6832,N_8881);
or U14703 (N_14703,N_6162,N_5094);
nand U14704 (N_14704,N_6724,N_9301);
nand U14705 (N_14705,N_6400,N_5199);
nand U14706 (N_14706,N_6858,N_5217);
nor U14707 (N_14707,N_7193,N_9380);
nor U14708 (N_14708,N_7755,N_9464);
or U14709 (N_14709,N_7355,N_9627);
nand U14710 (N_14710,N_6368,N_5998);
and U14711 (N_14711,N_8265,N_5383);
xor U14712 (N_14712,N_9252,N_7127);
xnor U14713 (N_14713,N_8752,N_7489);
xnor U14714 (N_14714,N_5061,N_9977);
and U14715 (N_14715,N_7512,N_6389);
or U14716 (N_14716,N_7757,N_5949);
or U14717 (N_14717,N_6665,N_6191);
nor U14718 (N_14718,N_9852,N_7685);
nand U14719 (N_14719,N_7977,N_7683);
nor U14720 (N_14720,N_9795,N_5024);
nor U14721 (N_14721,N_9013,N_6646);
or U14722 (N_14722,N_5867,N_8064);
nor U14723 (N_14723,N_7663,N_8601);
nand U14724 (N_14724,N_9337,N_6718);
nand U14725 (N_14725,N_7586,N_5276);
nor U14726 (N_14726,N_7144,N_8973);
and U14727 (N_14727,N_9023,N_8317);
nor U14728 (N_14728,N_7482,N_9297);
or U14729 (N_14729,N_7437,N_7528);
nand U14730 (N_14730,N_9192,N_9324);
xor U14731 (N_14731,N_5679,N_8493);
xor U14732 (N_14732,N_9370,N_7312);
nand U14733 (N_14733,N_9874,N_5326);
or U14734 (N_14734,N_9832,N_7244);
or U14735 (N_14735,N_7817,N_8954);
nor U14736 (N_14736,N_5865,N_9547);
or U14737 (N_14737,N_6871,N_9292);
and U14738 (N_14738,N_6252,N_8801);
nand U14739 (N_14739,N_5365,N_6773);
and U14740 (N_14740,N_6026,N_9671);
nand U14741 (N_14741,N_9079,N_8624);
nor U14742 (N_14742,N_8086,N_7648);
nor U14743 (N_14743,N_8136,N_5476);
and U14744 (N_14744,N_9873,N_5802);
nand U14745 (N_14745,N_5443,N_6484);
nand U14746 (N_14746,N_5490,N_8023);
and U14747 (N_14747,N_9309,N_6165);
nor U14748 (N_14748,N_5856,N_5317);
nand U14749 (N_14749,N_5778,N_8915);
nor U14750 (N_14750,N_9488,N_5223);
or U14751 (N_14751,N_7297,N_7348);
and U14752 (N_14752,N_6572,N_8096);
xor U14753 (N_14753,N_8278,N_9268);
xor U14754 (N_14754,N_5960,N_7821);
nor U14755 (N_14755,N_9339,N_9598);
and U14756 (N_14756,N_6676,N_5904);
or U14757 (N_14757,N_9953,N_6085);
nand U14758 (N_14758,N_8819,N_5641);
or U14759 (N_14759,N_7198,N_8957);
or U14760 (N_14760,N_9868,N_8885);
nand U14761 (N_14761,N_7511,N_9389);
and U14762 (N_14762,N_6165,N_7513);
and U14763 (N_14763,N_6195,N_5106);
or U14764 (N_14764,N_6047,N_7159);
and U14765 (N_14765,N_7024,N_6147);
or U14766 (N_14766,N_5112,N_6431);
and U14767 (N_14767,N_7456,N_9272);
nand U14768 (N_14768,N_9018,N_5457);
and U14769 (N_14769,N_7760,N_6869);
nor U14770 (N_14770,N_7503,N_9922);
or U14771 (N_14771,N_9426,N_9183);
and U14772 (N_14772,N_8382,N_8204);
and U14773 (N_14773,N_8901,N_9666);
nor U14774 (N_14774,N_7701,N_8079);
nand U14775 (N_14775,N_9552,N_7664);
or U14776 (N_14776,N_7133,N_5919);
or U14777 (N_14777,N_9185,N_8493);
xor U14778 (N_14778,N_7830,N_9044);
or U14779 (N_14779,N_6029,N_9087);
xor U14780 (N_14780,N_8882,N_8580);
nand U14781 (N_14781,N_8802,N_5027);
or U14782 (N_14782,N_8829,N_9230);
nand U14783 (N_14783,N_6842,N_6148);
xor U14784 (N_14784,N_5932,N_8656);
or U14785 (N_14785,N_8651,N_9781);
nand U14786 (N_14786,N_5193,N_5052);
or U14787 (N_14787,N_7481,N_8398);
and U14788 (N_14788,N_9505,N_6802);
and U14789 (N_14789,N_6743,N_6749);
xnor U14790 (N_14790,N_5404,N_9078);
nand U14791 (N_14791,N_5459,N_7881);
xnor U14792 (N_14792,N_5172,N_5279);
nor U14793 (N_14793,N_6070,N_6615);
and U14794 (N_14794,N_5609,N_5534);
or U14795 (N_14795,N_5439,N_5077);
or U14796 (N_14796,N_5292,N_8276);
and U14797 (N_14797,N_9205,N_5497);
nor U14798 (N_14798,N_5905,N_7300);
nand U14799 (N_14799,N_6777,N_8107);
nor U14800 (N_14800,N_7176,N_5025);
nand U14801 (N_14801,N_8139,N_5180);
xor U14802 (N_14802,N_8794,N_9454);
xor U14803 (N_14803,N_8520,N_6766);
xor U14804 (N_14804,N_8131,N_5941);
and U14805 (N_14805,N_6164,N_8515);
nor U14806 (N_14806,N_7329,N_8294);
or U14807 (N_14807,N_5062,N_8001);
and U14808 (N_14808,N_9271,N_5092);
nand U14809 (N_14809,N_6456,N_8612);
xor U14810 (N_14810,N_6829,N_7891);
and U14811 (N_14811,N_9093,N_6427);
and U14812 (N_14812,N_8577,N_7078);
and U14813 (N_14813,N_8080,N_5415);
nor U14814 (N_14814,N_6208,N_7039);
nor U14815 (N_14815,N_8939,N_6679);
nand U14816 (N_14816,N_5624,N_6802);
and U14817 (N_14817,N_7372,N_9530);
and U14818 (N_14818,N_5488,N_6217);
xor U14819 (N_14819,N_9318,N_6819);
nand U14820 (N_14820,N_6460,N_5728);
or U14821 (N_14821,N_9240,N_9238);
and U14822 (N_14822,N_5392,N_7416);
nand U14823 (N_14823,N_7277,N_5514);
nand U14824 (N_14824,N_6868,N_5317);
nor U14825 (N_14825,N_7944,N_7226);
nor U14826 (N_14826,N_8032,N_6793);
xor U14827 (N_14827,N_6379,N_8800);
nand U14828 (N_14828,N_7990,N_7771);
nand U14829 (N_14829,N_7875,N_8972);
xor U14830 (N_14830,N_7073,N_5526);
xor U14831 (N_14831,N_8400,N_7419);
or U14832 (N_14832,N_5383,N_5002);
or U14833 (N_14833,N_8038,N_8753);
xor U14834 (N_14834,N_9025,N_6696);
or U14835 (N_14835,N_7580,N_6195);
nor U14836 (N_14836,N_7635,N_9472);
nor U14837 (N_14837,N_5771,N_6262);
nor U14838 (N_14838,N_5174,N_8214);
or U14839 (N_14839,N_8033,N_9978);
nor U14840 (N_14840,N_7931,N_6171);
nand U14841 (N_14841,N_6507,N_6454);
xnor U14842 (N_14842,N_9562,N_9481);
nor U14843 (N_14843,N_7230,N_5699);
xnor U14844 (N_14844,N_9263,N_6410);
or U14845 (N_14845,N_7169,N_7378);
nor U14846 (N_14846,N_8393,N_5934);
and U14847 (N_14847,N_9111,N_5547);
xnor U14848 (N_14848,N_8224,N_5460);
and U14849 (N_14849,N_6723,N_7855);
or U14850 (N_14850,N_6335,N_9670);
xor U14851 (N_14851,N_6064,N_7998);
and U14852 (N_14852,N_7893,N_9776);
nor U14853 (N_14853,N_7198,N_6602);
nand U14854 (N_14854,N_6786,N_5355);
nor U14855 (N_14855,N_5300,N_7640);
and U14856 (N_14856,N_5312,N_9204);
or U14857 (N_14857,N_8900,N_6588);
and U14858 (N_14858,N_7900,N_7578);
nor U14859 (N_14859,N_9046,N_6949);
or U14860 (N_14860,N_6015,N_6886);
or U14861 (N_14861,N_8603,N_7165);
or U14862 (N_14862,N_6662,N_7281);
and U14863 (N_14863,N_5374,N_5243);
nor U14864 (N_14864,N_9845,N_5175);
nand U14865 (N_14865,N_8998,N_6251);
or U14866 (N_14866,N_5031,N_9896);
nor U14867 (N_14867,N_8287,N_6052);
and U14868 (N_14868,N_6839,N_7502);
or U14869 (N_14869,N_8287,N_9293);
nand U14870 (N_14870,N_8917,N_8799);
or U14871 (N_14871,N_9291,N_5559);
nor U14872 (N_14872,N_8663,N_9763);
nor U14873 (N_14873,N_8600,N_5908);
or U14874 (N_14874,N_5905,N_5404);
nand U14875 (N_14875,N_5103,N_5969);
or U14876 (N_14876,N_9207,N_9443);
xnor U14877 (N_14877,N_7093,N_6906);
xnor U14878 (N_14878,N_9197,N_6865);
nor U14879 (N_14879,N_5888,N_5027);
nor U14880 (N_14880,N_6109,N_7202);
xnor U14881 (N_14881,N_8230,N_8610);
nor U14882 (N_14882,N_7319,N_7139);
nor U14883 (N_14883,N_8313,N_9785);
nor U14884 (N_14884,N_9071,N_8425);
or U14885 (N_14885,N_5152,N_8193);
nand U14886 (N_14886,N_5808,N_5669);
and U14887 (N_14887,N_7433,N_7059);
and U14888 (N_14888,N_6191,N_7788);
nand U14889 (N_14889,N_9889,N_8588);
xor U14890 (N_14890,N_6057,N_9924);
nor U14891 (N_14891,N_9634,N_8560);
nand U14892 (N_14892,N_8620,N_9244);
and U14893 (N_14893,N_7522,N_8960);
nor U14894 (N_14894,N_8879,N_6281);
nor U14895 (N_14895,N_5970,N_9448);
or U14896 (N_14896,N_6413,N_8243);
nor U14897 (N_14897,N_7488,N_5500);
nor U14898 (N_14898,N_5554,N_7878);
and U14899 (N_14899,N_7000,N_8955);
xor U14900 (N_14900,N_9125,N_6120);
xor U14901 (N_14901,N_5239,N_6052);
or U14902 (N_14902,N_8869,N_5843);
or U14903 (N_14903,N_7728,N_7554);
or U14904 (N_14904,N_5199,N_8257);
nand U14905 (N_14905,N_8533,N_9187);
or U14906 (N_14906,N_8191,N_5754);
nor U14907 (N_14907,N_7176,N_7942);
xnor U14908 (N_14908,N_8544,N_9969);
and U14909 (N_14909,N_9379,N_6717);
xnor U14910 (N_14910,N_7213,N_6311);
or U14911 (N_14911,N_9290,N_5657);
and U14912 (N_14912,N_8213,N_9933);
and U14913 (N_14913,N_9894,N_8553);
nand U14914 (N_14914,N_8325,N_7189);
nor U14915 (N_14915,N_8556,N_6214);
and U14916 (N_14916,N_9995,N_6164);
nand U14917 (N_14917,N_7581,N_7985);
xor U14918 (N_14918,N_8009,N_6132);
or U14919 (N_14919,N_7120,N_6579);
and U14920 (N_14920,N_9924,N_6040);
nor U14921 (N_14921,N_5701,N_9310);
nor U14922 (N_14922,N_6452,N_8766);
and U14923 (N_14923,N_8753,N_6602);
xor U14924 (N_14924,N_9350,N_8241);
nor U14925 (N_14925,N_6885,N_8687);
or U14926 (N_14926,N_6298,N_9932);
or U14927 (N_14927,N_9595,N_8720);
nor U14928 (N_14928,N_6290,N_6269);
xor U14929 (N_14929,N_6435,N_8921);
nand U14930 (N_14930,N_5628,N_5825);
and U14931 (N_14931,N_9791,N_5249);
xor U14932 (N_14932,N_5639,N_7149);
nor U14933 (N_14933,N_5609,N_5629);
nor U14934 (N_14934,N_5350,N_6674);
xor U14935 (N_14935,N_6550,N_7792);
xor U14936 (N_14936,N_9229,N_9315);
and U14937 (N_14937,N_8027,N_8552);
and U14938 (N_14938,N_6105,N_6055);
or U14939 (N_14939,N_6169,N_9609);
nor U14940 (N_14940,N_8028,N_6438);
nor U14941 (N_14941,N_6988,N_5066);
xor U14942 (N_14942,N_7929,N_8257);
or U14943 (N_14943,N_7992,N_9577);
nor U14944 (N_14944,N_6515,N_9870);
nor U14945 (N_14945,N_9845,N_6363);
nor U14946 (N_14946,N_7160,N_8429);
and U14947 (N_14947,N_5918,N_7848);
xor U14948 (N_14948,N_7235,N_7831);
and U14949 (N_14949,N_5868,N_6221);
nor U14950 (N_14950,N_9530,N_8749);
or U14951 (N_14951,N_6479,N_8648);
nor U14952 (N_14952,N_9012,N_6074);
xor U14953 (N_14953,N_7648,N_5871);
or U14954 (N_14954,N_5210,N_5576);
nor U14955 (N_14955,N_9497,N_9191);
nor U14956 (N_14956,N_7840,N_5647);
nand U14957 (N_14957,N_9777,N_6255);
nor U14958 (N_14958,N_6890,N_5599);
and U14959 (N_14959,N_8589,N_5375);
xor U14960 (N_14960,N_9935,N_7800);
nor U14961 (N_14961,N_7992,N_8150);
and U14962 (N_14962,N_7815,N_8125);
nand U14963 (N_14963,N_5526,N_7925);
nor U14964 (N_14964,N_6815,N_7106);
nand U14965 (N_14965,N_8788,N_7532);
or U14966 (N_14966,N_8823,N_5691);
and U14967 (N_14967,N_8697,N_8490);
nand U14968 (N_14968,N_6682,N_6663);
nand U14969 (N_14969,N_5360,N_7381);
nor U14970 (N_14970,N_9377,N_5831);
xor U14971 (N_14971,N_5824,N_8630);
nor U14972 (N_14972,N_7340,N_8416);
nor U14973 (N_14973,N_5407,N_7343);
nor U14974 (N_14974,N_8804,N_5213);
xnor U14975 (N_14975,N_8195,N_7676);
and U14976 (N_14976,N_8913,N_7513);
nor U14977 (N_14977,N_8106,N_8589);
or U14978 (N_14978,N_9209,N_7757);
nor U14979 (N_14979,N_9622,N_6682);
and U14980 (N_14980,N_7815,N_7034);
nor U14981 (N_14981,N_8730,N_6925);
and U14982 (N_14982,N_7410,N_6702);
and U14983 (N_14983,N_6126,N_9789);
xnor U14984 (N_14984,N_8198,N_7076);
and U14985 (N_14985,N_5339,N_7211);
nand U14986 (N_14986,N_7757,N_9067);
nor U14987 (N_14987,N_8780,N_7301);
xor U14988 (N_14988,N_9338,N_6396);
nand U14989 (N_14989,N_8406,N_9751);
or U14990 (N_14990,N_6498,N_6258);
or U14991 (N_14991,N_6050,N_6591);
and U14992 (N_14992,N_9185,N_8287);
nor U14993 (N_14993,N_9660,N_8272);
nor U14994 (N_14994,N_9836,N_5766);
or U14995 (N_14995,N_6653,N_5401);
nand U14996 (N_14996,N_6135,N_9426);
or U14997 (N_14997,N_6171,N_5595);
nor U14998 (N_14998,N_6946,N_7911);
and U14999 (N_14999,N_5846,N_5405);
nand U15000 (N_15000,N_12008,N_12237);
or U15001 (N_15001,N_13281,N_14065);
nor U15002 (N_15002,N_12478,N_12160);
and U15003 (N_15003,N_12889,N_13125);
nand U15004 (N_15004,N_12029,N_11850);
nand U15005 (N_15005,N_14300,N_14247);
nand U15006 (N_15006,N_14912,N_11098);
nand U15007 (N_15007,N_14558,N_10009);
or U15008 (N_15008,N_11639,N_13935);
and U15009 (N_15009,N_10429,N_11315);
xnor U15010 (N_15010,N_14739,N_13058);
xnor U15011 (N_15011,N_10182,N_13398);
nor U15012 (N_15012,N_14480,N_12632);
nand U15013 (N_15013,N_13893,N_11249);
nand U15014 (N_15014,N_12261,N_14210);
nor U15015 (N_15015,N_11414,N_14914);
and U15016 (N_15016,N_10595,N_11829);
xnor U15017 (N_15017,N_13662,N_14053);
nand U15018 (N_15018,N_11378,N_10589);
nand U15019 (N_15019,N_11805,N_14905);
or U15020 (N_15020,N_12064,N_12580);
xor U15021 (N_15021,N_13897,N_11761);
and U15022 (N_15022,N_11867,N_10486);
and U15023 (N_15023,N_14773,N_11253);
and U15024 (N_15024,N_11248,N_10105);
nor U15025 (N_15025,N_13369,N_13599);
xor U15026 (N_15026,N_12334,N_13700);
and U15027 (N_15027,N_14978,N_14075);
nor U15028 (N_15028,N_11105,N_12525);
and U15029 (N_15029,N_11936,N_13002);
xor U15030 (N_15030,N_12773,N_11721);
or U15031 (N_15031,N_11183,N_10163);
xnor U15032 (N_15032,N_13324,N_14462);
xor U15033 (N_15033,N_10336,N_11088);
nor U15034 (N_15034,N_10296,N_12583);
nand U15035 (N_15035,N_12420,N_14740);
xor U15036 (N_15036,N_10558,N_14568);
or U15037 (N_15037,N_13245,N_13944);
or U15038 (N_15038,N_14800,N_14158);
xnor U15039 (N_15039,N_14636,N_12318);
or U15040 (N_15040,N_14996,N_10270);
nor U15041 (N_15041,N_10534,N_13078);
nand U15042 (N_15042,N_13653,N_10667);
nor U15043 (N_15043,N_12876,N_11050);
nor U15044 (N_15044,N_11444,N_14391);
nor U15045 (N_15045,N_14529,N_13129);
nor U15046 (N_15046,N_13259,N_13060);
and U15047 (N_15047,N_13684,N_11106);
and U15048 (N_15048,N_14502,N_12852);
nand U15049 (N_15049,N_14850,N_12354);
nor U15050 (N_15050,N_10921,N_10982);
or U15051 (N_15051,N_10700,N_10398);
xnor U15052 (N_15052,N_11785,N_12813);
nor U15053 (N_15053,N_14389,N_10642);
nand U15054 (N_15054,N_11541,N_12652);
nor U15055 (N_15055,N_10627,N_10751);
xnor U15056 (N_15056,N_10251,N_14325);
nor U15057 (N_15057,N_12799,N_14493);
and U15058 (N_15058,N_10658,N_13524);
nor U15059 (N_15059,N_11672,N_13422);
nor U15060 (N_15060,N_11907,N_14433);
and U15061 (N_15061,N_10690,N_10613);
nor U15062 (N_15062,N_14876,N_12836);
nor U15063 (N_15063,N_12833,N_10086);
and U15064 (N_15064,N_12188,N_13400);
and U15065 (N_15065,N_11468,N_12447);
nand U15066 (N_15066,N_10910,N_13996);
nor U15067 (N_15067,N_14828,N_13315);
and U15068 (N_15068,N_13555,N_14018);
xnor U15069 (N_15069,N_10616,N_11154);
and U15070 (N_15070,N_14199,N_10634);
nand U15071 (N_15071,N_12186,N_13101);
nand U15072 (N_15072,N_14193,N_10779);
nor U15073 (N_15073,N_10004,N_14814);
xnor U15074 (N_15074,N_13337,N_10447);
or U15075 (N_15075,N_11202,N_10278);
and U15076 (N_15076,N_14104,N_13968);
nand U15077 (N_15077,N_12722,N_11512);
nand U15078 (N_15078,N_13900,N_14342);
nor U15079 (N_15079,N_11087,N_12646);
or U15080 (N_15080,N_10238,N_12359);
xnor U15081 (N_15081,N_10005,N_11518);
nor U15082 (N_15082,N_13250,N_10942);
or U15083 (N_15083,N_11575,N_13881);
or U15084 (N_15084,N_10783,N_14795);
nor U15085 (N_15085,N_10331,N_10709);
nor U15086 (N_15086,N_13045,N_14947);
nor U15087 (N_15087,N_11270,N_12746);
or U15088 (N_15088,N_10601,N_14805);
xor U15089 (N_15089,N_13163,N_12111);
and U15090 (N_15090,N_11796,N_12004);
or U15091 (N_15091,N_10615,N_13931);
and U15092 (N_15092,N_10473,N_11382);
nor U15093 (N_15093,N_13283,N_13044);
xnor U15094 (N_15094,N_14810,N_13674);
or U15095 (N_15095,N_14402,N_14553);
nor U15096 (N_15096,N_14596,N_14126);
nand U15097 (N_15097,N_11044,N_12647);
xnor U15098 (N_15098,N_10552,N_14903);
and U15099 (N_15099,N_13278,N_13956);
nor U15100 (N_15100,N_11727,N_13456);
or U15101 (N_15101,N_10402,N_12503);
nand U15102 (N_15102,N_12568,N_12310);
and U15103 (N_15103,N_12912,N_12792);
xnor U15104 (N_15104,N_11993,N_13731);
xnor U15105 (N_15105,N_13092,N_10519);
nand U15106 (N_15106,N_10040,N_12247);
and U15107 (N_15107,N_13572,N_12462);
nand U15108 (N_15108,N_14677,N_12806);
xnor U15109 (N_15109,N_12596,N_12293);
nand U15110 (N_15110,N_10323,N_10264);
or U15111 (N_15111,N_13114,N_14772);
and U15112 (N_15112,N_10769,N_11973);
or U15113 (N_15113,N_12013,N_11827);
nor U15114 (N_15114,N_11307,N_11905);
and U15115 (N_15115,N_11257,N_14484);
xor U15116 (N_15116,N_10316,N_14497);
nand U15117 (N_15117,N_14139,N_13710);
nor U15118 (N_15118,N_10633,N_14920);
or U15119 (N_15119,N_10015,N_12952);
or U15120 (N_15120,N_11640,N_12490);
and U15121 (N_15121,N_13067,N_11121);
nand U15122 (N_15122,N_13701,N_11464);
nand U15123 (N_15123,N_11294,N_10970);
or U15124 (N_15124,N_14608,N_11846);
nor U15125 (N_15125,N_13170,N_12241);
xnor U15126 (N_15126,N_14984,N_12951);
or U15127 (N_15127,N_13513,N_13272);
nand U15128 (N_15128,N_13759,N_11880);
or U15129 (N_15129,N_14085,N_12549);
nand U15130 (N_15130,N_10366,N_11886);
nand U15131 (N_15131,N_10891,N_14913);
or U15132 (N_15132,N_12970,N_10506);
and U15133 (N_15133,N_10889,N_13853);
nand U15134 (N_15134,N_11092,N_11400);
nand U15135 (N_15135,N_13074,N_13924);
xor U15136 (N_15136,N_10020,N_10137);
or U15137 (N_15137,N_11794,N_14244);
or U15138 (N_15138,N_11372,N_11490);
and U15139 (N_15139,N_11434,N_10666);
xnor U15140 (N_15140,N_11084,N_11064);
nand U15141 (N_15141,N_10508,N_13730);
or U15142 (N_15142,N_12655,N_11140);
xnor U15143 (N_15143,N_11412,N_12974);
xor U15144 (N_15144,N_10021,N_13346);
and U15145 (N_15145,N_12193,N_12692);
and U15146 (N_15146,N_10496,N_12807);
nand U15147 (N_15147,N_13015,N_14446);
or U15148 (N_15148,N_11071,N_14485);
nand U15149 (N_15149,N_11941,N_13951);
nor U15150 (N_15150,N_10051,N_11157);
nand U15151 (N_15151,N_11230,N_10579);
and U15152 (N_15152,N_14916,N_10947);
and U15153 (N_15153,N_11932,N_12963);
nand U15154 (N_15154,N_12663,N_11255);
nand U15155 (N_15155,N_10090,N_12234);
xnor U15156 (N_15156,N_11839,N_10155);
nor U15157 (N_15157,N_11531,N_10883);
xnor U15158 (N_15158,N_14915,N_10975);
or U15159 (N_15159,N_14812,N_13929);
xor U15160 (N_15160,N_13809,N_12515);
xor U15161 (N_15161,N_14892,N_10441);
or U15162 (N_15162,N_14015,N_14603);
and U15163 (N_15163,N_13589,N_14673);
xnor U15164 (N_15164,N_12971,N_13005);
or U15165 (N_15165,N_10629,N_10925);
xor U15166 (N_15166,N_14624,N_14815);
xor U15167 (N_15167,N_11356,N_10459);
nor U15168 (N_15168,N_10135,N_14404);
nor U15169 (N_15169,N_14185,N_13762);
or U15170 (N_15170,N_13692,N_14487);
and U15171 (N_15171,N_13746,N_14450);
xor U15172 (N_15172,N_13781,N_14243);
xnor U15173 (N_15173,N_10056,N_10263);
and U15174 (N_15174,N_10242,N_10121);
and U15175 (N_15175,N_13038,N_11842);
nand U15176 (N_15176,N_14718,N_13357);
xor U15177 (N_15177,N_13852,N_13468);
nand U15178 (N_15178,N_10950,N_14051);
xnor U15179 (N_15179,N_13778,N_10686);
nor U15180 (N_15180,N_13171,N_10810);
nand U15181 (N_15181,N_12638,N_10442);
xor U15182 (N_15182,N_13327,N_13506);
xnor U15183 (N_15183,N_14380,N_11415);
or U15184 (N_15184,N_13073,N_11738);
nand U15185 (N_15185,N_13528,N_10806);
nor U15186 (N_15186,N_14216,N_11890);
and U15187 (N_15187,N_13391,N_11205);
xor U15188 (N_15188,N_12795,N_10730);
nand U15189 (N_15189,N_13821,N_13247);
and U15190 (N_15190,N_10661,N_10913);
nor U15191 (N_15191,N_14349,N_11368);
nor U15192 (N_15192,N_10738,N_10964);
nor U15193 (N_15193,N_10591,N_12601);
xnor U15194 (N_15194,N_12244,N_11511);
and U15195 (N_15195,N_10837,N_14527);
nor U15196 (N_15196,N_13543,N_11859);
or U15197 (N_15197,N_11254,N_10969);
and U15198 (N_15198,N_11705,N_14198);
xor U15199 (N_15199,N_12329,N_12651);
xnor U15200 (N_15200,N_13796,N_13179);
or U15201 (N_15201,N_14960,N_13514);
nor U15202 (N_15202,N_12706,N_12623);
nand U15203 (N_15203,N_14521,N_11942);
nand U15204 (N_15204,N_10179,N_11013);
and U15205 (N_15205,N_13783,N_10100);
nor U15206 (N_15206,N_10070,N_11929);
or U15207 (N_15207,N_12194,N_14021);
or U15208 (N_15208,N_14345,N_11605);
nand U15209 (N_15209,N_12664,N_10292);
nand U15210 (N_15210,N_10432,N_11686);
nor U15211 (N_15211,N_10003,N_13289);
nor U15212 (N_15212,N_10492,N_14843);
xor U15213 (N_15213,N_12164,N_11323);
nand U15214 (N_15214,N_14834,N_11814);
nor U15215 (N_15215,N_13539,N_10032);
xnor U15216 (N_15216,N_11655,N_14826);
and U15217 (N_15217,N_10220,N_14897);
nand U15218 (N_15218,N_13494,N_11999);
nand U15219 (N_15219,N_10156,N_10229);
xor U15220 (N_15220,N_13891,N_11542);
xnor U15221 (N_15221,N_13342,N_10458);
and U15222 (N_15222,N_10113,N_13303);
or U15223 (N_15223,N_12180,N_12454);
nor U15224 (N_15224,N_10226,N_11723);
nor U15225 (N_15225,N_11118,N_13901);
and U15226 (N_15226,N_14797,N_13048);
xor U15227 (N_15227,N_14144,N_13379);
or U15228 (N_15228,N_14879,N_13328);
nor U15229 (N_15229,N_13030,N_13202);
nor U15230 (N_15230,N_13325,N_12408);
and U15231 (N_15231,N_12383,N_14824);
or U15232 (N_15232,N_11800,N_10415);
xnor U15233 (N_15233,N_13523,N_13651);
nand U15234 (N_15234,N_13595,N_14482);
nor U15235 (N_15235,N_10280,N_13384);
nor U15236 (N_15236,N_11070,N_12299);
or U15237 (N_15237,N_12994,N_13645);
nand U15238 (N_15238,N_12765,N_11494);
nor U15239 (N_15239,N_10048,N_14310);
xor U15240 (N_15240,N_13847,N_10770);
and U15241 (N_15241,N_11914,N_13641);
nand U15242 (N_15242,N_12197,N_14442);
or U15243 (N_15243,N_13209,N_10830);
nor U15244 (N_15244,N_10903,N_10944);
or U15245 (N_15245,N_10218,N_14518);
or U15246 (N_15246,N_12691,N_10499);
nand U15247 (N_15247,N_14143,N_10710);
xor U15248 (N_15248,N_12783,N_10013);
and U15249 (N_15249,N_11950,N_12223);
nor U15250 (N_15250,N_11495,N_10896);
xor U15251 (N_15251,N_14534,N_10685);
xnor U15252 (N_15252,N_10598,N_14398);
nand U15253 (N_15253,N_14737,N_12283);
and U15254 (N_15254,N_11446,N_14113);
nor U15255 (N_15255,N_12053,N_14930);
nand U15256 (N_15256,N_13949,N_14103);
and U15257 (N_15257,N_11110,N_12409);
xor U15258 (N_15258,N_12091,N_14659);
or U15259 (N_15259,N_10140,N_10334);
or U15260 (N_15260,N_14956,N_10592);
xor U15261 (N_15261,N_11038,N_12001);
or U15262 (N_15262,N_12217,N_12155);
xnor U15263 (N_15263,N_14069,N_12564);
and U15264 (N_15264,N_11833,N_11178);
xor U15265 (N_15265,N_11990,N_10481);
or U15266 (N_15266,N_14384,N_12399);
nor U15267 (N_15267,N_10721,N_11613);
nand U15268 (N_15268,N_10472,N_13848);
and U15269 (N_15269,N_11791,N_10082);
nor U15270 (N_15270,N_13512,N_10396);
xnor U15271 (N_15271,N_10553,N_13119);
xor U15272 (N_15272,N_13608,N_14291);
nand U15273 (N_15273,N_11740,N_11571);
and U15274 (N_15274,N_10906,N_12007);
xnor U15275 (N_15275,N_13583,N_14615);
xor U15276 (N_15276,N_11015,N_11685);
and U15277 (N_15277,N_14919,N_10528);
and U15278 (N_15278,N_13664,N_11832);
xnor U15279 (N_15279,N_13288,N_13688);
or U15280 (N_15280,N_14640,N_14159);
or U15281 (N_15281,N_10077,N_10389);
and U15282 (N_15282,N_13254,N_13139);
nor U15283 (N_15283,N_11055,N_12770);
nand U15284 (N_15284,N_14064,N_13872);
nor U15285 (N_15285,N_12395,N_10216);
xnor U15286 (N_15286,N_14288,N_12881);
and U15287 (N_15287,N_10992,N_10231);
and U15288 (N_15288,N_11526,N_11689);
or U15289 (N_15289,N_14286,N_11865);
xor U15290 (N_15290,N_11674,N_13909);
nor U15291 (N_15291,N_11696,N_11530);
nand U15292 (N_15292,N_11172,N_13994);
nand U15293 (N_15293,N_14767,N_10007);
and U15294 (N_15294,N_14923,N_14670);
nor U15295 (N_15295,N_10490,N_11312);
and U15296 (N_15296,N_10060,N_12469);
or U15297 (N_15297,N_11213,N_12088);
xor U15298 (N_15298,N_11609,N_11008);
and U15299 (N_15299,N_12452,N_14691);
or U15300 (N_15300,N_12352,N_11483);
or U15301 (N_15301,N_10711,N_10548);
nor U15302 (N_15302,N_10018,N_14076);
xor U15303 (N_15303,N_12896,N_10780);
xnor U15304 (N_15304,N_14801,N_14437);
nand U15305 (N_15305,N_13727,N_11091);
xor U15306 (N_15306,N_14990,N_14492);
xnor U15307 (N_15307,N_13983,N_12914);
xor U15308 (N_15308,N_11673,N_12927);
nand U15309 (N_15309,N_13823,N_12901);
xor U15310 (N_15310,N_13458,N_10976);
and U15311 (N_15311,N_11195,N_12514);
nand U15312 (N_15312,N_11974,N_11401);
nor U15313 (N_15313,N_10914,N_12906);
or U15314 (N_15314,N_10219,N_13370);
and U15315 (N_15315,N_11308,N_11864);
nand U15316 (N_15316,N_11365,N_10973);
and U15317 (N_15317,N_14412,N_11653);
xnor U15318 (N_15318,N_11036,N_11704);
xnor U15319 (N_15319,N_10495,N_14170);
nand U15320 (N_15320,N_13740,N_13266);
nor U15321 (N_15321,N_13803,N_13070);
nor U15322 (N_15322,N_10412,N_14741);
nor U15323 (N_15323,N_13226,N_11559);
nor U15324 (N_15324,N_13009,N_10045);
nand U15325 (N_15325,N_13818,N_12398);
or U15326 (N_15326,N_13162,N_14871);
nor U15327 (N_15327,N_12553,N_11767);
or U15328 (N_15328,N_12205,N_11712);
nand U15329 (N_15329,N_14593,N_12100);
and U15330 (N_15330,N_11471,N_13987);
xnor U15331 (N_15331,N_12280,N_13261);
nor U15332 (N_15332,N_12089,N_10536);
xor U15333 (N_15333,N_11159,N_13175);
xor U15334 (N_15334,N_12769,N_10234);
or U15335 (N_15335,N_14292,N_13576);
nand U15336 (N_15336,N_11759,N_11169);
xnor U15337 (N_15337,N_12500,N_14887);
and U15338 (N_15338,N_10407,N_12232);
nand U15339 (N_15339,N_11340,N_11185);
or U15340 (N_15340,N_12995,N_13188);
nand U15341 (N_15341,N_12911,N_12338);
nor U15342 (N_15342,N_10697,N_11977);
and U15343 (N_15343,N_14410,N_11131);
nor U15344 (N_15344,N_13100,N_13023);
or U15345 (N_15345,N_14403,N_11247);
nand U15346 (N_15346,N_14804,N_11509);
or U15347 (N_15347,N_13947,N_13981);
nor U15348 (N_15348,N_13186,N_12885);
and U15349 (N_15349,N_11028,N_12364);
nand U15350 (N_15350,N_11196,N_13560);
nor U15351 (N_15351,N_12708,N_13934);
or U15352 (N_15352,N_12882,N_14878);
xnor U15353 (N_15353,N_11928,N_13992);
nor U15354 (N_15354,N_10380,N_13211);
or U15355 (N_15355,N_10621,N_12723);
xor U15356 (N_15356,N_13414,N_13066);
nor U15357 (N_15357,N_14322,N_13098);
and U15358 (N_15358,N_13428,N_13239);
nor U15359 (N_15359,N_11775,N_12046);
nand U15360 (N_15360,N_10109,N_10993);
nor U15361 (N_15361,N_13235,N_14661);
and U15362 (N_15362,N_11289,N_13349);
nor U15363 (N_15363,N_10813,N_10924);
and U15364 (N_15364,N_13362,N_13197);
nor U15365 (N_15365,N_13671,N_12909);
xnor U15366 (N_15366,N_11465,N_11297);
nor U15367 (N_15367,N_10868,N_14283);
nand U15368 (N_15368,N_10243,N_13216);
nand U15369 (N_15369,N_10504,N_10375);
and U15370 (N_15370,N_11717,N_11399);
or U15371 (N_15371,N_12033,N_11458);
and U15372 (N_15372,N_10204,N_12864);
nand U15373 (N_15373,N_10230,N_12919);
xor U15374 (N_15374,N_12548,N_13902);
nor U15375 (N_15375,N_10359,N_14809);
nand U15376 (N_15376,N_13627,N_11987);
xor U15377 (N_15377,N_12316,N_14898);
and U15378 (N_15378,N_11228,N_10773);
nand U15379 (N_15379,N_10450,N_10577);
or U15380 (N_15380,N_14995,N_11947);
nand U15381 (N_15381,N_12529,N_14825);
and U15382 (N_15382,N_12934,N_13718);
or U15383 (N_15383,N_10554,N_11888);
xor U15384 (N_15384,N_14362,N_10948);
xor U15385 (N_15385,N_14970,N_12533);
nor U15386 (N_15386,N_10724,N_14277);
nor U15387 (N_15387,N_11630,N_14318);
nand U15388 (N_15388,N_13178,N_14893);
or U15389 (N_15389,N_13722,N_14265);
xor U15390 (N_15390,N_12169,N_14336);
nand U15391 (N_15391,N_12945,N_11459);
nand U15392 (N_15392,N_11077,N_14116);
nand U15393 (N_15393,N_12973,N_14394);
and U15394 (N_15394,N_11500,N_14551);
nand U15395 (N_15395,N_13433,N_14846);
and U15396 (N_15396,N_14781,N_11309);
nor U15397 (N_15397,N_12410,N_13658);
nor U15398 (N_15398,N_12323,N_11810);
nor U15399 (N_15399,N_12425,N_13850);
and U15400 (N_15400,N_11144,N_10146);
xnor U15401 (N_15401,N_10475,N_13293);
or U15402 (N_15402,N_13372,N_13252);
and U15403 (N_15403,N_12543,N_13166);
nand U15404 (N_15404,N_10171,N_12895);
and U15405 (N_15405,N_13427,N_11758);
xnor U15406 (N_15406,N_10625,N_14606);
nor U15407 (N_15407,N_14862,N_10319);
or U15408 (N_15408,N_10831,N_10571);
nand U15409 (N_15409,N_13308,N_12279);
and U15410 (N_15410,N_12242,N_11944);
or U15411 (N_15411,N_13380,N_13046);
or U15412 (N_15412,N_14589,N_13227);
and U15413 (N_15413,N_12070,N_14419);
xor U15414 (N_15414,N_12841,N_13610);
or U15415 (N_15415,N_13706,N_11748);
and U15416 (N_15416,N_13165,N_13383);
and U15417 (N_15417,N_12118,N_14604);
nand U15418 (N_15418,N_12146,N_12278);
nor U15419 (N_15419,N_12892,N_13320);
and U15420 (N_15420,N_11838,N_14307);
nor U15421 (N_15421,N_14082,N_10977);
nor U15422 (N_15422,N_14109,N_14189);
and U15423 (N_15423,N_11584,N_14359);
or U15424 (N_15424,N_12745,N_12311);
nand U15425 (N_15425,N_12137,N_14114);
and U15426 (N_15426,N_10332,N_12270);
or U15427 (N_15427,N_11007,N_12990);
nand U15428 (N_15428,N_12439,N_10130);
or U15429 (N_15429,N_12397,N_13057);
or U15430 (N_15430,N_11124,N_11732);
nand U15431 (N_15431,N_11787,N_14863);
or U15432 (N_15432,N_13779,N_13142);
xnor U15433 (N_15433,N_13302,N_11508);
nand U15434 (N_15434,N_12024,N_10606);
and U15435 (N_15435,N_12041,N_10527);
nor U15436 (N_15436,N_14561,N_11894);
or U15437 (N_15437,N_12050,N_13221);
nor U15438 (N_15438,N_13151,N_14983);
and U15439 (N_15439,N_12742,N_11598);
xor U15440 (N_15440,N_12348,N_11646);
nor U15441 (N_15441,N_12018,N_11388);
and U15442 (N_15442,N_13973,N_12516);
and U15443 (N_15443,N_13242,N_10755);
nor U15444 (N_15444,N_11349,N_10956);
and U15445 (N_15445,N_12363,N_10289);
nor U15446 (N_15446,N_14697,N_14790);
nand U15447 (N_15447,N_12558,N_10065);
nand U15448 (N_15448,N_12459,N_14117);
or U15449 (N_15449,N_10016,N_10797);
xor U15450 (N_15450,N_12600,N_13036);
xnor U15451 (N_15451,N_12255,N_11343);
and U15452 (N_15452,N_11879,N_13265);
and U15453 (N_15453,N_11707,N_14874);
or U15454 (N_15454,N_13336,N_11428);
xnor U15455 (N_15455,N_14488,N_13262);
nor U15456 (N_15456,N_11352,N_14902);
or U15457 (N_15457,N_10605,N_10767);
xor U15458 (N_15458,N_12757,N_10960);
nor U15459 (N_15459,N_12052,N_11029);
or U15460 (N_15460,N_13210,N_11777);
nand U15461 (N_15461,N_11854,N_11171);
nand U15462 (N_15462,N_10559,N_11432);
nand U15463 (N_15463,N_13084,N_11953);
xnor U15464 (N_15464,N_12267,N_12435);
and U15465 (N_15465,N_11250,N_10456);
and U15466 (N_15466,N_11636,N_14866);
nor U15467 (N_15467,N_13780,N_13896);
and U15468 (N_15468,N_10731,N_14141);
or U15469 (N_15469,N_14260,N_10035);
nand U15470 (N_15470,N_14782,N_10215);
or U15471 (N_15471,N_12767,N_12532);
or U15472 (N_15472,N_10849,N_14569);
nand U15473 (N_15473,N_10543,N_14386);
xor U15474 (N_15474,N_14855,N_11109);
or U15475 (N_15475,N_14026,N_12289);
and U15476 (N_15476,N_13373,N_11650);
xor U15477 (N_15477,N_12755,N_10378);
xnor U15478 (N_15478,N_11398,N_14233);
nor U15479 (N_15479,N_12659,N_10134);
nand U15480 (N_15480,N_10097,N_13003);
xor U15481 (N_15481,N_14148,N_12204);
nand U15482 (N_15482,N_14627,N_12626);
or U15483 (N_15483,N_14279,N_14547);
xnor U15484 (N_15484,N_10454,N_13564);
xnor U15485 (N_15485,N_14885,N_13785);
nand U15486 (N_15486,N_13614,N_11687);
nand U15487 (N_15487,N_14516,N_10712);
nand U15488 (N_15488,N_13470,N_11090);
and U15489 (N_15489,N_14702,N_12263);
and U15490 (N_15490,N_10256,N_10699);
nor U15491 (N_15491,N_10392,N_11397);
nor U15492 (N_15492,N_14102,N_13864);
and U15493 (N_15493,N_12291,N_13215);
nand U15494 (N_15494,N_10855,N_12654);
xor U15495 (N_15495,N_10940,N_10981);
and U15496 (N_15496,N_12272,N_11628);
and U15497 (N_15497,N_13980,N_10271);
nand U15498 (N_15498,N_10728,N_11692);
nand U15499 (N_15499,N_12473,N_11460);
xor U15500 (N_15500,N_11203,N_11709);
xnor U15501 (N_15501,N_14925,N_12181);
or U15502 (N_15502,N_12026,N_13425);
and U15503 (N_15503,N_13953,N_12750);
or U15504 (N_15504,N_14329,N_10514);
or U15505 (N_15505,N_10714,N_10503);
xnor U15506 (N_15506,N_12358,N_12872);
and U15507 (N_15507,N_11778,N_14038);
nor U15508 (N_15508,N_12861,N_10560);
nand U15509 (N_15509,N_11688,N_11235);
nor U15510 (N_15510,N_11361,N_10647);
nand U15511 (N_15511,N_14605,N_12677);
nor U15512 (N_15512,N_12547,N_12844);
nor U15513 (N_15513,N_14723,N_14316);
and U15514 (N_15514,N_13797,N_14417);
nand U15515 (N_15515,N_11793,N_13829);
or U15516 (N_15516,N_13519,N_13150);
and U15517 (N_15517,N_12159,N_10335);
nand U15518 (N_15518,N_12382,N_10012);
nor U15519 (N_15519,N_10946,N_13812);
xor U15520 (N_15520,N_13537,N_11986);
xnor U15521 (N_15521,N_11593,N_10261);
xor U15522 (N_15522,N_11431,N_11411);
xor U15523 (N_15523,N_10972,N_13366);
or U15524 (N_15524,N_11946,N_12006);
nor U15525 (N_15525,N_13007,N_12812);
xnor U15526 (N_15526,N_11348,N_10079);
or U15527 (N_15527,N_10143,N_14583);
nor U15528 (N_15528,N_13620,N_14352);
xnor U15529 (N_15529,N_10118,N_10817);
or U15530 (N_15530,N_10870,N_11893);
nor U15531 (N_15531,N_10632,N_11616);
or U15532 (N_15532,N_14963,N_11935);
and U15533 (N_15533,N_10812,N_10428);
or U15534 (N_15534,N_13566,N_13657);
nor U15535 (N_15535,N_11417,N_10224);
xnor U15536 (N_15536,N_12305,N_14177);
nand U15537 (N_15537,N_11219,N_14676);
xnor U15538 (N_15538,N_13134,N_10857);
xor U15539 (N_15539,N_10909,N_14333);
or U15540 (N_15540,N_12377,N_12555);
or U15541 (N_15541,N_13360,N_12847);
or U15542 (N_15542,N_10808,N_12612);
or U15543 (N_15543,N_13683,N_14302);
nand U15544 (N_15544,N_10725,N_14149);
and U15545 (N_15545,N_11871,N_13606);
xnor U15546 (N_15546,N_12522,N_13086);
and U15547 (N_15547,N_14848,N_14669);
nor U15548 (N_15548,N_14927,N_13693);
xor U15549 (N_15549,N_14759,N_11006);
or U15550 (N_15550,N_10083,N_11525);
or U15551 (N_15551,N_14201,N_14592);
or U15552 (N_15552,N_14634,N_12068);
xnor U15553 (N_15553,N_10794,N_10547);
nor U15554 (N_15554,N_14167,N_11966);
nand U15555 (N_15555,N_10600,N_13721);
xor U15556 (N_15556,N_13410,N_14136);
or U15557 (N_15557,N_11849,N_12258);
nor U15558 (N_15558,N_10892,N_11299);
or U15559 (N_15559,N_11117,N_10381);
nand U15560 (N_15560,N_11698,N_10662);
nor U15561 (N_15561,N_13787,N_12226);
xor U15562 (N_15562,N_11702,N_11964);
xor U15563 (N_15563,N_10672,N_12456);
and U15564 (N_15564,N_13922,N_10825);
xor U15565 (N_15565,N_10068,N_11802);
and U15566 (N_15566,N_10153,N_10011);
nor U15567 (N_15567,N_11912,N_10568);
and U15568 (N_15568,N_13766,N_14839);
and U15569 (N_15569,N_13619,N_14582);
and U15570 (N_15570,N_14436,N_14917);
or U15571 (N_15571,N_12821,N_10067);
or U15572 (N_15572,N_13085,N_13348);
xnor U15573 (N_15573,N_12665,N_14266);
or U15574 (N_15574,N_12154,N_11057);
nand U15575 (N_15575,N_12787,N_14533);
nand U15576 (N_15576,N_10607,N_12959);
or U15577 (N_15577,N_13013,N_13600);
and U15578 (N_15578,N_10599,N_13103);
or U15579 (N_15579,N_14474,N_10421);
nor U15580 (N_15580,N_14667,N_13670);
xor U15581 (N_15581,N_14409,N_11831);
nand U15582 (N_15582,N_10037,N_12421);
xor U15583 (N_15583,N_10920,N_13364);
and U15584 (N_15584,N_11735,N_13088);
xor U15585 (N_15585,N_12304,N_11279);
xnor U15586 (N_15586,N_12002,N_13313);
nor U15587 (N_15587,N_11667,N_13412);
xnor U15588 (N_15588,N_10217,N_14572);
nand U15589 (N_15589,N_11173,N_13811);
and U15590 (N_15590,N_12360,N_12749);
or U15591 (N_15591,N_14774,N_10643);
or U15592 (N_15592,N_13229,N_10430);
and U15593 (N_15593,N_10784,N_11965);
nand U15594 (N_15594,N_12309,N_13546);
and U15595 (N_15595,N_13748,N_11755);
and U15596 (N_15596,N_12135,N_14305);
nor U15597 (N_15597,N_10128,N_11313);
nor U15598 (N_15598,N_13984,N_11770);
nor U15599 (N_15599,N_10756,N_11874);
nand U15600 (N_15600,N_11059,N_11291);
nand U15601 (N_15601,N_14675,N_13948);
xnor U15602 (N_15602,N_12130,N_10576);
nand U15603 (N_15603,N_12401,N_13873);
xnor U15604 (N_15604,N_10901,N_11782);
nor U15605 (N_15605,N_10286,N_12565);
and U15606 (N_15606,N_14657,N_10122);
or U15607 (N_15607,N_13611,N_10638);
nand U15608 (N_15608,N_14563,N_12489);
xor U15609 (N_15609,N_12740,N_13813);
nor U15610 (N_15610,N_12729,N_12766);
nand U15611 (N_15611,N_10227,N_14508);
and U15612 (N_15612,N_13716,N_14628);
and U15613 (N_15613,N_10085,N_13886);
and U15614 (N_15614,N_13267,N_14466);
nor U15615 (N_15615,N_11961,N_14382);
and U15616 (N_15616,N_12947,N_14165);
or U15617 (N_15617,N_11737,N_11125);
or U15618 (N_15618,N_11258,N_14153);
nor U15619 (N_15619,N_10801,N_10740);
xor U15620 (N_15620,N_13689,N_13257);
and U15621 (N_15621,N_11537,N_13039);
xnor U15622 (N_15622,N_14899,N_14770);
xor U15623 (N_15623,N_11165,N_14859);
nor U15624 (N_15624,N_11823,N_12481);
nand U15625 (N_15625,N_10139,N_12736);
nor U15626 (N_15626,N_13361,N_14997);
nand U15627 (N_15627,N_11407,N_10990);
nor U15628 (N_15628,N_10183,N_11877);
xnor U15629 (N_15629,N_10517,N_14035);
nand U15630 (N_15630,N_13094,N_14837);
and U15631 (N_15631,N_10006,N_12458);
nor U15632 (N_15632,N_13581,N_13063);
or U15633 (N_15633,N_10066,N_10790);
and U15634 (N_15634,N_11572,N_11350);
nor U15635 (N_15635,N_12402,N_11336);
nor U15636 (N_15636,N_11046,N_10161);
and U15637 (N_15637,N_14094,N_13939);
and U15638 (N_15638,N_14687,N_10312);
nor U15639 (N_15639,N_12785,N_12403);
nor U15640 (N_15640,N_14602,N_12675);
nand U15641 (N_15641,N_11678,N_10322);
nand U15642 (N_15642,N_13578,N_11396);
xor U15643 (N_15643,N_14010,N_11037);
and U15644 (N_15644,N_11076,N_12907);
and U15645 (N_15645,N_13580,N_11021);
nor U15646 (N_15646,N_14212,N_12545);
or U15647 (N_15647,N_12185,N_10114);
xnor U15648 (N_15648,N_13501,N_11099);
nand U15649 (N_15649,N_10943,N_12980);
nor U15650 (N_15650,N_12030,N_13451);
and U15651 (N_15651,N_13915,N_11744);
or U15652 (N_15652,N_10356,N_10419);
nand U15653 (N_15653,N_13478,N_13885);
nor U15654 (N_15654,N_14453,N_10582);
and U15655 (N_15655,N_11532,N_14385);
and U15656 (N_15656,N_10551,N_13660);
or U15657 (N_15657,N_10505,N_10513);
and U15658 (N_15658,N_11741,N_10368);
or U15659 (N_15659,N_13930,N_14183);
nand U15660 (N_15660,N_11281,N_10639);
nor U15661 (N_15661,N_14794,N_10440);
or U15662 (N_15662,N_10819,N_12619);
nor U15663 (N_15663,N_10955,N_11014);
nor U15664 (N_15664,N_11634,N_14526);
or U15665 (N_15665,N_11011,N_14922);
xnor U15666 (N_15666,N_12000,N_10650);
and U15667 (N_15667,N_10520,N_10445);
or U15668 (N_15668,N_10031,N_14660);
or U15669 (N_15669,N_12987,N_13686);
xnor U15670 (N_15670,N_12170,N_13777);
or U15671 (N_15671,N_10994,N_11353);
xnor U15672 (N_15672,N_11366,N_10357);
and U15673 (N_15673,N_10235,N_14957);
xor U15674 (N_15674,N_11423,N_13936);
nand U15675 (N_15675,N_10737,N_14748);
and U15676 (N_15676,N_14796,N_14730);
or U15677 (N_15677,N_14469,N_11660);
nand U15678 (N_15678,N_11816,N_13876);
nand U15679 (N_15679,N_13715,N_14296);
or U15680 (N_15680,N_13582,N_14037);
and U15681 (N_15681,N_10583,N_13429);
or U15682 (N_15682,N_10030,N_14190);
and U15683 (N_15683,N_12732,N_13687);
and U15684 (N_15684,N_12333,N_10715);
nor U15685 (N_15685,N_13107,N_13263);
xnor U15686 (N_15686,N_13967,N_13329);
or U15687 (N_15687,N_12349,N_13164);
nor U15688 (N_15688,N_14254,N_10168);
or U15689 (N_15689,N_12519,N_10383);
xnor U15690 (N_15690,N_13894,N_11546);
nand U15691 (N_15691,N_12560,N_14686);
and U15692 (N_15692,N_14744,N_13858);
or U15693 (N_15693,N_12637,N_14931);
nand U15694 (N_15694,N_14418,N_11133);
xor U15695 (N_15695,N_11844,N_11019);
and U15696 (N_15696,N_13482,N_10170);
nor U15697 (N_15697,N_12697,N_11504);
xnor U15698 (N_15698,N_14750,N_12288);
or U15699 (N_15699,N_12801,N_11241);
nor U15700 (N_15700,N_13368,N_14680);
nand U15701 (N_15701,N_11948,N_14991);
nand U15702 (N_15702,N_10745,N_14219);
nor U15703 (N_15703,N_13041,N_12989);
or U15704 (N_15704,N_10815,N_10034);
nand U15705 (N_15705,N_10689,N_11420);
nand U15706 (N_15706,N_14560,N_13786);
nand U15707 (N_15707,N_12282,N_12225);
nor U15708 (N_15708,N_13958,N_13841);
and U15709 (N_15709,N_13676,N_11756);
and U15710 (N_15710,N_14778,N_11904);
and U15711 (N_15711,N_12230,N_14643);
or U15712 (N_15712,N_14769,N_12385);
and U15713 (N_15713,N_12233,N_10966);
or U15714 (N_15714,N_10562,N_14032);
and U15715 (N_15715,N_11733,N_14475);
and U15716 (N_15716,N_10330,N_12804);
xnor U15717 (N_15717,N_10811,N_13594);
nand U15718 (N_15718,N_10269,N_14465);
nand U15719 (N_15719,N_13377,N_10954);
xor U15720 (N_15720,N_14784,N_10327);
nor U15721 (N_15721,N_12948,N_13499);
nor U15722 (N_15722,N_13908,N_14588);
or U15723 (N_15723,N_13401,N_14431);
nor U15724 (N_15724,N_10501,N_14789);
or U15725 (N_15725,N_10640,N_13472);
nor U15726 (N_15726,N_11768,N_12798);
nand U15727 (N_15727,N_13810,N_11403);
nor U15728 (N_15728,N_14369,N_14022);
nor U15729 (N_15729,N_10320,N_10774);
and U15730 (N_15730,N_14538,N_13149);
or U15731 (N_15731,N_12012,N_12405);
nor U15732 (N_15732,N_13075,N_11405);
or U15733 (N_15733,N_11215,N_13156);
nor U15734 (N_15734,N_14043,N_10361);
nor U15735 (N_15735,N_13794,N_12407);
or U15736 (N_15736,N_13999,N_14423);
nand U15737 (N_15737,N_13898,N_12958);
xnor U15738 (N_15738,N_14847,N_14424);
nand U15739 (N_15739,N_12455,N_10371);
xnor U15740 (N_15740,N_14982,N_12893);
or U15741 (N_15741,N_14227,N_14591);
or U15742 (N_15742,N_11424,N_10406);
nand U15743 (N_15743,N_13489,N_11031);
nor U15744 (N_15744,N_13995,N_14505);
and U15745 (N_15745,N_13446,N_10985);
nor U15746 (N_15746,N_10986,N_12062);
and U15747 (N_15747,N_11311,N_10028);
nor U15748 (N_15748,N_12502,N_14335);
or U15749 (N_15749,N_11439,N_12028);
nand U15750 (N_15750,N_13024,N_13626);
xnor U15751 (N_15751,N_10148,N_13940);
xor U15752 (N_15752,N_13228,N_10002);
xnor U15753 (N_15753,N_13301,N_11135);
nor U15754 (N_15754,N_11493,N_14162);
or U15755 (N_15755,N_13174,N_14191);
nor U15756 (N_15756,N_10963,N_12540);
and U15757 (N_15757,N_14347,N_13256);
and U15758 (N_15758,N_12944,N_13678);
xnor U15759 (N_15759,N_11684,N_12521);
and U15760 (N_15760,N_13828,N_12903);
nand U15761 (N_15761,N_10228,N_13681);
and U15762 (N_15762,N_14057,N_10252);
or U15763 (N_15763,N_14061,N_13111);
xnor U15764 (N_15764,N_13128,N_13264);
or U15765 (N_15765,N_10435,N_10660);
xor U15766 (N_15766,N_12035,N_10485);
nor U15767 (N_15767,N_12176,N_14060);
nor U15768 (N_15768,N_13443,N_11119);
and U15769 (N_15769,N_11080,N_13407);
or U15770 (N_15770,N_14392,N_13826);
xnor U15771 (N_15771,N_14452,N_12346);
nor U15772 (N_15772,N_13394,N_13431);
xnor U15773 (N_15773,N_13473,N_10154);
nor U15774 (N_15774,N_14157,N_10590);
nand U15775 (N_15775,N_11317,N_10565);
nand U15776 (N_15776,N_11583,N_12823);
nor U15777 (N_15777,N_10507,N_12709);
nor U15778 (N_15778,N_14429,N_13061);
nor U15779 (N_15779,N_14974,N_14268);
nor U15780 (N_15780,N_13833,N_11664);
and U15781 (N_15781,N_10515,N_10567);
and U15782 (N_15782,N_10791,N_14792);
xor U15783 (N_15783,N_14000,N_10782);
and U15784 (N_15784,N_10203,N_13304);
and U15785 (N_15785,N_10865,N_11322);
nand U15786 (N_15786,N_12495,N_13287);
nor U15787 (N_15787,N_10836,N_14120);
and U15788 (N_15788,N_12542,N_14539);
nor U15789 (N_15789,N_13331,N_14028);
or U15790 (N_15790,N_13351,N_10748);
xnor U15791 (N_15791,N_14584,N_13271);
nor U15792 (N_15792,N_13381,N_13405);
and U15793 (N_15793,N_13732,N_12714);
nand U15794 (N_15794,N_11949,N_11209);
and U15795 (N_15795,N_14528,N_12136);
or U15796 (N_15796,N_10372,N_11962);
nand U15797 (N_15797,N_11150,N_11883);
nor U15798 (N_15798,N_12222,N_13510);
nand U15799 (N_15799,N_12929,N_11058);
nor U15800 (N_15800,N_10908,N_14363);
xor U15801 (N_15801,N_14644,N_14752);
xnor U15802 (N_15802,N_10123,N_11697);
or U15803 (N_15803,N_12686,N_12734);
nor U15804 (N_15804,N_13464,N_12081);
nand U15805 (N_15805,N_11543,N_11657);
xnor U15806 (N_15806,N_11720,N_10190);
xnor U15807 (N_15807,N_11392,N_13274);
and U15808 (N_15808,N_10893,N_13363);
xnor U15809 (N_15809,N_13839,N_12695);
or U15810 (N_15810,N_11980,N_10705);
and U15811 (N_15811,N_11455,N_10025);
or U15812 (N_15812,N_11766,N_10047);
or U15813 (N_15813,N_12719,N_13093);
nor U15814 (N_15814,N_14111,N_13863);
and U15815 (N_15815,N_14091,N_12537);
nor U15816 (N_15816,N_12950,N_14900);
nand U15817 (N_15817,N_14443,N_14119);
nand U15818 (N_15818,N_14554,N_12015);
nor U15819 (N_15819,N_11430,N_10678);
or U15820 (N_15820,N_12888,N_14567);
nor U15821 (N_15821,N_10719,N_13712);
nor U15822 (N_15822,N_14315,N_11573);
or U15823 (N_15823,N_10848,N_10523);
and U15824 (N_15824,N_13492,N_10355);
xor U15825 (N_15825,N_14852,N_13444);
nand U15826 (N_15826,N_14454,N_13634);
and U15827 (N_15827,N_10403,N_12344);
xor U15828 (N_15828,N_13053,N_10116);
or U15829 (N_15829,N_14638,N_12819);
nand U15830 (N_15830,N_12977,N_11093);
nand U15831 (N_15831,N_12760,N_13733);
nor U15832 (N_15832,N_14445,N_11222);
and U15833 (N_15833,N_10311,N_12440);
nand U15834 (N_15834,N_11959,N_12192);
xor U15835 (N_15835,N_10934,N_14617);
xor U15836 (N_15836,N_10839,N_12577);
and U15837 (N_15837,N_12961,N_10349);
or U15838 (N_15838,N_12641,N_13652);
nand U15839 (N_15839,N_10126,N_10493);
or U15840 (N_15840,N_12618,N_12744);
xnor U15841 (N_15841,N_11237,N_14263);
nor U15842 (N_15842,N_11561,N_10405);
or U15843 (N_15843,N_14304,N_14535);
xor U15844 (N_15844,N_12925,N_10706);
and U15845 (N_15845,N_10641,N_11752);
nand U15846 (N_15846,N_10274,N_13776);
nor U15847 (N_15847,N_14164,N_10911);
and U15848 (N_15848,N_14749,N_12590);
nand U15849 (N_15849,N_12631,N_11835);
xnor U15850 (N_15850,N_13844,N_12758);
xnor U15851 (N_15851,N_12999,N_12488);
xnor U15852 (N_15852,N_12576,N_13051);
nor U15853 (N_15853,N_11586,N_12862);
xnor U15854 (N_15854,N_10930,N_10957);
nand U15855 (N_15855,N_10483,N_11069);
nand U15856 (N_15856,N_13851,N_10423);
xnor U15857 (N_15857,N_13734,N_14935);
and U15858 (N_15858,N_12979,N_14712);
nand U15859 (N_15859,N_10014,N_12115);
or U15860 (N_15860,N_12084,N_10895);
or U15861 (N_15861,N_14868,N_13081);
or U15862 (N_15862,N_13889,N_11700);
nand U15863 (N_15863,N_14448,N_12754);
xnor U15864 (N_15864,N_10747,N_12144);
or U15865 (N_15865,N_13775,N_12245);
nand U15866 (N_15866,N_11669,N_12325);
nand U15867 (N_15867,N_10022,N_14985);
nand U15868 (N_15868,N_12800,N_11469);
and U15869 (N_15869,N_10258,N_10597);
xnor U15870 (N_15870,N_10879,N_14351);
or U15871 (N_15871,N_12032,N_12069);
nand U15872 (N_15872,N_14470,N_12866);
or U15873 (N_15873,N_14695,N_13837);
nor U15874 (N_15874,N_12132,N_10098);
nor U15875 (N_15875,N_14328,N_12879);
xor U15876 (N_15876,N_12842,N_13234);
nor U15877 (N_15877,N_11619,N_12669);
nor U15878 (N_15878,N_10828,N_14343);
nand U15879 (N_15879,N_13253,N_13424);
nor U15880 (N_15880,N_12157,N_10129);
and U15881 (N_15881,N_13068,N_12436);
and U15882 (N_15882,N_13913,N_10847);
and U15883 (N_15883,N_11830,N_10604);
nand U15884 (N_15884,N_13630,N_11454);
xor U15885 (N_15885,N_11743,N_10851);
and U15886 (N_15886,N_13806,N_11989);
or U15887 (N_15887,N_13880,N_12775);
and U15888 (N_15888,N_11956,N_10859);
nor U15889 (N_15889,N_12450,N_13644);
or U15890 (N_15890,N_12427,N_13577);
and U15891 (N_15891,N_10470,N_12827);
xor U15892 (N_15892,N_10469,N_13867);
nand U15893 (N_15893,N_13957,N_11018);
xnor U15894 (N_15894,N_14703,N_10133);
nor U15895 (N_15895,N_10619,N_13617);
and U15896 (N_15896,N_14215,N_10418);
and U15897 (N_15897,N_11642,N_10433);
or U15898 (N_15898,N_11143,N_10631);
xor U15899 (N_15899,N_12962,N_10017);
nand U15900 (N_15900,N_14971,N_13140);
nand U15901 (N_15901,N_13974,N_11954);
nor U15902 (N_15902,N_13836,N_12759);
and U15903 (N_15903,N_11482,N_10905);
or U15904 (N_15904,N_10237,N_14147);
and U15905 (N_15905,N_11034,N_14714);
nor U15906 (N_15906,N_12182,N_11338);
or U15907 (N_15907,N_12998,N_12090);
nor U15908 (N_15908,N_12913,N_12867);
nor U15909 (N_15909,N_13062,N_12964);
xor U15910 (N_15910,N_12725,N_10257);
or U15911 (N_15911,N_11332,N_10890);
nand U15912 (N_15912,N_12116,N_12884);
nor U15913 (N_15913,N_14998,N_11882);
nor U15914 (N_15914,N_11538,N_12541);
or U15915 (N_15915,N_11022,N_11916);
nor U15916 (N_15916,N_10814,N_13238);
or U15917 (N_15917,N_14753,N_13770);
xnor U15918 (N_15918,N_10795,N_10820);
nand U15919 (N_15919,N_11513,N_10185);
or U15920 (N_15920,N_12284,N_13804);
and U15921 (N_15921,N_12196,N_11265);
and U15922 (N_15922,N_10904,N_13986);
nor U15923 (N_15923,N_13126,N_11895);
and U15924 (N_15924,N_11734,N_13049);
nand U15925 (N_15925,N_13454,N_11901);
nor U15926 (N_15926,N_13338,N_11288);
and U15927 (N_15927,N_14393,N_10965);
or U15928 (N_15928,N_12367,N_13725);
and U15929 (N_15929,N_12203,N_12924);
xnor U15930 (N_15930,N_14217,N_12887);
or U15931 (N_15931,N_13830,N_10733);
nand U15932 (N_15932,N_10807,N_12392);
nand U15933 (N_15933,N_11271,N_11120);
xnor U15934 (N_15934,N_11497,N_11360);
nor U15935 (N_15935,N_11701,N_11967);
nand U15936 (N_15936,N_13065,N_11301);
nand U15937 (N_15937,N_13542,N_11244);
nor U15938 (N_15938,N_14756,N_11462);
xor U15939 (N_15939,N_13601,N_11718);
and U15940 (N_15940,N_12449,N_11739);
nor U15941 (N_15941,N_14729,N_12935);
or U15942 (N_15942,N_13172,N_10046);
xor U15943 (N_15943,N_11342,N_10894);
or U15944 (N_15944,N_12830,N_12530);
nand U15945 (N_15945,N_13022,N_14907);
nor U15946 (N_15946,N_12504,N_10826);
xor U15947 (N_15947,N_11590,N_12699);
and U15948 (N_15948,N_11781,N_11671);
xnor U15949 (N_15949,N_12832,N_12221);
nor U15950 (N_15950,N_14918,N_10058);
nor U15951 (N_15951,N_10410,N_14736);
nor U15952 (N_15952,N_14115,N_12301);
nor U15953 (N_15953,N_13534,N_11607);
xnor U15954 (N_15954,N_12843,N_14587);
nand U15955 (N_15955,N_12614,N_11193);
nand U15956 (N_15956,N_11528,N_12138);
and U15957 (N_15957,N_11303,N_11010);
nand U15958 (N_15958,N_14964,N_12808);
nor U15959 (N_15959,N_12212,N_12674);
or U15960 (N_15960,N_13933,N_12264);
xnor U15961 (N_15961,N_13792,N_11751);
nor U15962 (N_15962,N_11376,N_11229);
nor U15963 (N_15963,N_13760,N_10187);
and U15964 (N_15964,N_10675,N_11218);
and U15965 (N_15965,N_11729,N_14576);
nand U15966 (N_15966,N_13144,N_11992);
xor U15967 (N_15967,N_13102,N_13497);
nor U15968 (N_15968,N_11045,N_13793);
nor U15969 (N_15969,N_11413,N_11114);
nor U15970 (N_15970,N_10832,N_10382);
xor U15971 (N_15971,N_12321,N_14231);
xnor U15972 (N_15972,N_11602,N_12793);
and U15973 (N_15973,N_11370,N_12776);
or U15974 (N_15974,N_10850,N_14775);
xor U15975 (N_15975,N_11274,N_12593);
nor U15976 (N_15976,N_14168,N_12351);
xor U15977 (N_15977,N_14207,N_12639);
nor U15978 (N_15978,N_13054,N_12905);
and U15979 (N_15979,N_10900,N_11515);
xnor U15980 (N_15980,N_14821,N_14285);
nor U15981 (N_15981,N_12595,N_12575);
xnor U15982 (N_15982,N_11535,N_14506);
xnor U15983 (N_15983,N_11385,N_11002);
xor U15984 (N_15984,N_10671,N_11860);
and U15985 (N_15985,N_13764,N_10680);
or U15986 (N_15986,N_10339,N_11618);
and U15987 (N_15987,N_12434,N_13219);
nor U15988 (N_15988,N_10347,N_13386);
xnor U15989 (N_15989,N_11680,N_13371);
nor U15990 (N_15990,N_10928,N_13511);
xnor U15991 (N_15991,N_11763,N_13017);
or U15992 (N_15992,N_14665,N_12134);
nand U15993 (N_15993,N_13493,N_12139);
and U15994 (N_15994,N_13773,N_14955);
nor U15995 (N_15995,N_13323,N_10399);
and U15996 (N_15996,N_10306,N_10147);
or U15997 (N_15997,N_14169,N_12253);
xor U15998 (N_15998,N_11547,N_13800);
nand U15999 (N_15999,N_12531,N_12101);
and U16000 (N_16000,N_12712,N_12058);
nand U16001 (N_16001,N_12786,N_11523);
nand U16002 (N_16002,N_14999,N_10462);
nand U16003 (N_16003,N_12127,N_11190);
nand U16004 (N_16004,N_14353,N_10345);
and U16005 (N_16005,N_13435,N_13033);
nand U16006 (N_16006,N_13176,N_12563);
and U16007 (N_16007,N_14123,N_10293);
nand U16008 (N_16008,N_10151,N_13541);
nor U16009 (N_16009,N_11435,N_12748);
xnor U16010 (N_16010,N_12501,N_14586);
nand U16011 (N_16011,N_13815,N_11083);
nor U16012 (N_16012,N_13032,N_13319);
xor U16013 (N_16013,N_14545,N_11210);
and U16014 (N_16014,N_14357,N_14099);
nor U16015 (N_16015,N_12324,N_13525);
nand U16016 (N_16016,N_12551,N_11005);
or U16017 (N_16017,N_13439,N_10838);
and U16018 (N_16018,N_12431,N_13476);
and U16019 (N_16019,N_10983,N_10884);
xnor U16020 (N_16020,N_11473,N_14738);
or U16021 (N_16021,N_14287,N_12873);
xor U16022 (N_16022,N_11009,N_12751);
nor U16023 (N_16023,N_13280,N_10474);
xor U16024 (N_16024,N_14705,N_10630);
or U16025 (N_16025,N_11820,N_14334);
xor U16026 (N_16026,N_14127,N_11772);
nor U16027 (N_16027,N_11395,N_14299);
nand U16028 (N_16028,N_11576,N_14574);
nand U16029 (N_16029,N_13498,N_10844);
and U16030 (N_16030,N_11452,N_12578);
and U16031 (N_16031,N_14838,N_10262);
and U16032 (N_16032,N_12371,N_10537);
and U16033 (N_16033,N_14760,N_10735);
xor U16034 (N_16034,N_12366,N_11869);
xor U16035 (N_16035,N_13612,N_12661);
xor U16036 (N_16036,N_11184,N_13618);
xor U16037 (N_16037,N_13735,N_12150);
and U16038 (N_16038,N_14662,N_14229);
or U16039 (N_16039,N_14213,N_12556);
nor U16040 (N_16040,N_12331,N_14245);
nor U16041 (N_16041,N_11030,N_14590);
and U16042 (N_16042,N_12140,N_13993);
xnor U16043 (N_16043,N_10169,N_12648);
and U16044 (N_16044,N_13952,N_11485);
and U16045 (N_16045,N_12528,N_13286);
nand U16046 (N_16046,N_13237,N_11466);
xor U16047 (N_16047,N_11945,N_12335);
or U16048 (N_16048,N_12273,N_14030);
nor U16049 (N_16049,N_12051,N_12174);
xnor U16050 (N_16050,N_12124,N_11402);
nor U16051 (N_16051,N_11138,N_13173);
nor U16052 (N_16052,N_12636,N_10693);
nor U16053 (N_16053,N_14441,N_12523);
nand U16054 (N_16054,N_11127,N_14205);
nor U16055 (N_16055,N_10365,N_14829);
xnor U16056 (N_16056,N_10823,N_12298);
xor U16057 (N_16057,N_13533,N_10677);
nand U16058 (N_16058,N_13292,N_13113);
and U16059 (N_16059,N_11001,N_13521);
or U16060 (N_16060,N_12968,N_12165);
nand U16061 (N_16061,N_14645,N_12014);
and U16062 (N_16062,N_12622,N_13353);
nand U16063 (N_16063,N_11548,N_13457);
nand U16064 (N_16064,N_14074,N_14014);
and U16065 (N_16065,N_10027,N_12839);
or U16066 (N_16066,N_14253,N_13399);
or U16067 (N_16067,N_12043,N_13719);
nor U16068 (N_16068,N_12768,N_14802);
or U16069 (N_16069,N_13605,N_12546);
and U16070 (N_16070,N_13198,N_11156);
nand U16071 (N_16071,N_12559,N_12942);
nand U16072 (N_16072,N_10388,N_14860);
xnor U16073 (N_16073,N_14882,N_11910);
nor U16074 (N_16074,N_12086,N_10736);
nor U16075 (N_16075,N_10075,N_12413);
and U16076 (N_16076,N_13339,N_11256);
or U16077 (N_16077,N_13868,N_11656);
xor U16078 (N_16078,N_10991,N_12259);
xor U16079 (N_16079,N_13807,N_13403);
and U16080 (N_16080,N_12591,N_12306);
or U16081 (N_16081,N_13801,N_10716);
xor U16082 (N_16082,N_10239,N_12199);
nor U16083 (N_16083,N_14639,N_13522);
or U16084 (N_16084,N_11757,N_12805);
nor U16085 (N_16085,N_12161,N_10212);
nor U16086 (N_16086,N_12448,N_13460);
or U16087 (N_16087,N_11522,N_14098);
and U16088 (N_16088,N_12191,N_12173);
or U16089 (N_16089,N_13535,N_12327);
or U16090 (N_16090,N_13469,N_14537);
xnor U16091 (N_16091,N_12055,N_10749);
nor U16092 (N_16092,N_11625,N_14954);
and U16093 (N_16093,N_10255,N_11463);
nand U16094 (N_16094,N_14459,N_10958);
nor U16095 (N_16095,N_13964,N_13491);
nand U16096 (N_16096,N_12009,N_11600);
or U16097 (N_16097,N_10288,N_11346);
nor U16098 (N_16098,N_14130,N_14808);
xor U16099 (N_16099,N_14658,N_13668);
xnor U16100 (N_16100,N_13040,N_13859);
nand U16101 (N_16101,N_14224,N_11457);
or U16102 (N_16102,N_14510,N_10024);
nand U16103 (N_16103,N_10044,N_12561);
or U16104 (N_16104,N_12109,N_10804);
nand U16105 (N_16105,N_14180,N_10809);
or U16106 (N_16106,N_13184,N_13680);
xnor U16107 (N_16107,N_11527,N_14672);
nor U16108 (N_16108,N_13465,N_14755);
or U16109 (N_16109,N_11958,N_10691);
xnor U16110 (N_16110,N_13069,N_13574);
nor U16111 (N_16111,N_11539,N_13515);
and U16112 (N_16112,N_13453,N_14237);
nor U16113 (N_16113,N_10464,N_14531);
xor U16114 (N_16114,N_13376,N_14251);
or U16115 (N_16115,N_11503,N_13350);
nor U16116 (N_16116,N_11889,N_10785);
nor U16117 (N_16117,N_14467,N_13923);
or U16118 (N_16118,N_12728,N_12328);
and U16119 (N_16119,N_10240,N_13545);
nand U16120 (N_16120,N_14951,N_11911);
nand U16121 (N_16121,N_13123,N_10757);
nor U16122 (N_16122,N_11226,N_12172);
or U16123 (N_16123,N_11565,N_11148);
xnor U16124 (N_16124,N_10933,N_10142);
and U16125 (N_16125,N_10967,N_11367);
or U16126 (N_16126,N_11779,N_13761);
nand U16127 (N_16127,N_13737,N_14786);
nor U16128 (N_16128,N_13463,N_13131);
and U16129 (N_16129,N_13782,N_12189);
nor U16130 (N_16130,N_14058,N_12021);
xor U16131 (N_16131,N_14735,N_11979);
nand U16132 (N_16132,N_14430,N_14544);
or U16133 (N_16133,N_14949,N_14211);
nor U16134 (N_16134,N_14671,N_14009);
or U16135 (N_16135,N_10704,N_12771);
nor U16136 (N_16136,N_13690,N_10535);
nand U16137 (N_16137,N_14888,N_10041);
nand U16138 (N_16138,N_11876,N_13072);
and U16139 (N_16139,N_10937,N_13720);
nand U16140 (N_16140,N_12218,N_12849);
and U16141 (N_16141,N_13946,N_11305);
nand U16142 (N_16142,N_13314,N_10696);
and U16143 (N_16143,N_14841,N_14308);
or U16144 (N_16144,N_13225,N_10789);
nor U16145 (N_16145,N_11703,N_13059);
and U16146 (N_16146,N_11197,N_11824);
nor U16147 (N_16147,N_11909,N_10912);
xor U16148 (N_16148,N_13146,N_10120);
and U16149 (N_16149,N_12249,N_14373);
xnor U16150 (N_16150,N_14520,N_14468);
xor U16151 (N_16151,N_12082,N_11448);
nand U16152 (N_16152,N_10679,N_11433);
and U16153 (N_16153,N_10866,N_10115);
nor U16154 (N_16154,N_14220,N_13321);
nand U16155 (N_16155,N_13154,N_10961);
nand U16156 (N_16156,N_13496,N_11477);
xor U16157 (N_16157,N_13004,N_14642);
xnor U16158 (N_16158,N_10225,N_14683);
and U16159 (N_16159,N_12780,N_13487);
xnor U16160 (N_16160,N_12739,N_11094);
and U16161 (N_16161,N_11217,N_10196);
or U16162 (N_16162,N_14239,N_13270);
xor U16163 (N_16163,N_14324,N_12391);
nor U16164 (N_16164,N_13665,N_14062);
xor U16165 (N_16165,N_10664,N_10718);
nor U16166 (N_16166,N_10039,N_13385);
xor U16167 (N_16167,N_12922,N_14089);
nor U16168 (N_16168,N_14152,N_14339);
nor U16169 (N_16169,N_14282,N_11521);
nand U16170 (N_16170,N_11708,N_14613);
xnor U16171 (N_16171,N_12838,N_13663);
or U16172 (N_16172,N_12678,N_13448);
nor U16173 (N_16173,N_12057,N_12077);
nand U16174 (N_16174,N_14851,N_13832);
xnor U16175 (N_16175,N_13108,N_13471);
xnor U16176 (N_16176,N_14652,N_10308);
or U16177 (N_16177,N_12362,N_12653);
nand U16178 (N_16178,N_11771,N_10917);
nand U16179 (N_16179,N_12715,N_11817);
xnor U16180 (N_16180,N_12941,N_10489);
xor U16181 (N_16181,N_12790,N_10094);
and U16182 (N_16182,N_11931,N_11130);
xor U16183 (N_16183,N_13479,N_14566);
xor U16184 (N_16184,N_14763,N_13136);
or U16185 (N_16185,N_12243,N_14101);
nor U16186 (N_16186,N_13928,N_13695);
or U16187 (N_16187,N_14002,N_12588);
xnor U16188 (N_16188,N_13001,N_12538);
and U16189 (N_16189,N_14174,N_11875);
nor U16190 (N_16190,N_13402,N_10061);
or U16191 (N_16191,N_11736,N_10214);
nor U16192 (N_16192,N_11795,N_11621);
nand U16193 (N_16193,N_13426,N_10471);
and U16194 (N_16194,N_11610,N_10325);
nor U16195 (N_16195,N_13333,N_10455);
nand U16196 (N_16196,N_12404,N_11111);
or U16197 (N_16197,N_11676,N_14494);
or U16198 (N_16198,N_13666,N_10887);
xnor U16199 (N_16199,N_14543,N_14052);
xor U16200 (N_16200,N_11581,N_13406);
xnor U16201 (N_16201,N_12477,N_14451);
nor U16202 (N_16202,N_12552,N_10862);
nor U16203 (N_16203,N_11919,N_14631);
or U16204 (N_16204,N_11577,N_13236);
xnor U16205 (N_16205,N_13845,N_13095);
or U16206 (N_16206,N_10119,N_14776);
nand U16207 (N_16207,N_10324,N_13861);
and U16208 (N_16208,N_12307,N_11053);
nor U16209 (N_16209,N_11730,N_13788);
xor U16210 (N_16210,N_14066,N_10352);
or U16211 (N_16211,N_12662,N_14238);
nand U16212 (N_16212,N_14909,N_13284);
nand U16213 (N_16213,N_11115,N_12509);
nor U16214 (N_16214,N_13442,N_11128);
xnor U16215 (N_16215,N_13192,N_13874);
nor U16216 (N_16216,N_14623,N_11510);
or U16217 (N_16217,N_13441,N_14942);
xor U16218 (N_16218,N_10413,N_12206);
or U16219 (N_16219,N_13214,N_10344);
and U16220 (N_16220,N_11383,N_10348);
or U16221 (N_16221,N_12589,N_10502);
nand U16222 (N_16222,N_11287,N_11578);
nor U16223 (N_16223,N_14565,N_11004);
and U16224 (N_16224,N_11491,N_13971);
xnor U16225 (N_16225,N_11540,N_12296);
and U16226 (N_16226,N_14788,N_14731);
nand U16227 (N_16227,N_12379,N_12871);
nand U16228 (N_16228,N_10222,N_14405);
xnor U16229 (N_16229,N_12630,N_11555);
xnor U16230 (N_16230,N_10164,N_10099);
and U16231 (N_16231,N_11663,N_14601);
or U16232 (N_16232,N_11223,N_11714);
xor U16233 (N_16233,N_13026,N_10144);
nand U16234 (N_16234,N_11591,N_11926);
and U16235 (N_16235,N_11164,N_10309);
and U16236 (N_16236,N_12730,N_11813);
xnor U16237 (N_16237,N_14936,N_14525);
nand U16238 (N_16238,N_13708,N_12219);
or U16239 (N_16239,N_13104,N_12417);
nor U16240 (N_16240,N_13153,N_12315);
xor U16241 (N_16241,N_10845,N_10302);
xor U16242 (N_16242,N_10437,N_11566);
and U16243 (N_16243,N_14455,N_12920);
nor U16244 (N_16244,N_14105,N_12753);
nand U16245 (N_16245,N_10778,N_14059);
or U16246 (N_16246,N_11821,N_11073);
xnor U16247 (N_16247,N_14259,N_13276);
and U16248 (N_16248,N_11644,N_10223);
nand U16249 (N_16249,N_14503,N_11903);
nor U16250 (N_16250,N_10453,N_14258);
or U16251 (N_16251,N_13109,N_13316);
and U16252 (N_16252,N_13490,N_10771);
nor U16253 (N_16253,N_13392,N_10042);
or U16254 (N_16254,N_13569,N_14311);
and U16255 (N_16255,N_12356,N_12389);
or U16256 (N_16256,N_14223,N_10676);
xnor U16257 (N_16257,N_12926,N_11097);
or U16258 (N_16258,N_13418,N_12645);
and U16259 (N_16259,N_13805,N_13042);
or U16260 (N_16260,N_14685,N_10563);
and U16261 (N_16261,N_12045,N_14414);
or U16262 (N_16262,N_14320,N_12597);
and U16263 (N_16263,N_11017,N_10180);
or U16264 (N_16264,N_10764,N_14941);
or U16265 (N_16265,N_11048,N_13682);
and U16266 (N_16266,N_13691,N_10054);
nand U16267 (N_16267,N_10283,N_10313);
or U16268 (N_16268,N_11635,N_12534);
nor U16269 (N_16269,N_13318,N_11262);
nand U16270 (N_16270,N_10328,N_14515);
or U16271 (N_16271,N_14621,N_13505);
and U16272 (N_16272,N_14881,N_10055);
nor U16273 (N_16273,N_12373,N_12513);
or U16274 (N_16274,N_13090,N_13099);
or U16275 (N_16275,N_14570,N_12486);
and U16276 (N_16276,N_13430,N_12883);
or U16277 (N_16277,N_10654,N_11808);
nand U16278 (N_16278,N_12396,N_14765);
nand U16279 (N_16279,N_11467,N_12326);
xor U16280 (N_16280,N_14071,N_11161);
or U16281 (N_16281,N_14046,N_14987);
or U16282 (N_16282,N_10923,N_11479);
nor U16283 (N_16283,N_14597,N_12067);
or U16284 (N_16284,N_12341,N_11819);
nor U16285 (N_16285,N_12096,N_14321);
xor U16286 (N_16286,N_13588,N_14249);
nor U16287 (N_16287,N_14042,N_14594);
and U16288 (N_16288,N_11275,N_11878);
xnor U16289 (N_16289,N_12216,N_12092);
nor U16290 (N_16290,N_10636,N_11180);
nor U16291 (N_16291,N_11060,N_12526);
xor U16292 (N_16292,N_10460,N_11716);
xor U16293 (N_16293,N_13639,N_14641);
and U16294 (N_16294,N_10360,N_10136);
and U16295 (N_16295,N_10194,N_11693);
nor U16296 (N_16296,N_10670,N_10602);
and U16297 (N_16297,N_11331,N_11243);
and U16298 (N_16298,N_10213,N_10979);
and U16299 (N_16299,N_14440,N_12153);
nand U16300 (N_16300,N_11104,N_14135);
and U16301 (N_16301,N_14696,N_14420);
and U16302 (N_16302,N_14161,N_13127);
and U16303 (N_16303,N_13739,N_14289);
nor U16304 (N_16304,N_12465,N_11344);
or U16305 (N_16305,N_14364,N_10096);
xnor U16306 (N_16306,N_13918,N_13255);
or U16307 (N_16307,N_13365,N_12418);
nor U16308 (N_16308,N_13685,N_13260);
nor U16309 (N_16309,N_11476,N_12290);
nand U16310 (N_16310,N_10907,N_12195);
xor U16311 (N_16311,N_10996,N_12202);
or U16312 (N_16312,N_13621,N_12956);
or U16313 (N_16313,N_12162,N_11815);
or U16314 (N_16314,N_11750,N_11359);
nand U16315 (N_16315,N_14270,N_12381);
nand U16316 (N_16316,N_10610,N_11622);
or U16317 (N_16317,N_14854,N_12374);
or U16318 (N_16318,N_10744,N_14086);
or U16319 (N_16319,N_13246,N_10342);
xnor U16320 (N_16320,N_13483,N_10645);
or U16321 (N_16321,N_10713,N_13802);
or U16322 (N_16322,N_12438,N_14378);
xor U16323 (N_16323,N_14853,N_10902);
xor U16324 (N_16324,N_12498,N_11812);
or U16325 (N_16325,N_13557,N_12025);
nand U16326 (N_16326,N_10422,N_14742);
nor U16327 (N_16327,N_12487,N_13825);
nor U16328 (N_16328,N_10949,N_12112);
or U16329 (N_16329,N_10668,N_14681);
and U16330 (N_16330,N_10867,N_12772);
xnor U16331 (N_16331,N_12063,N_13884);
and U16332 (N_16332,N_11214,N_11421);
or U16333 (N_16333,N_12860,N_14840);
xnor U16334 (N_16334,N_13115,N_13205);
xor U16335 (N_16335,N_11529,N_13404);
or U16336 (N_16336,N_13177,N_13118);
xor U16337 (N_16337,N_11749,N_12536);
xnor U16338 (N_16338,N_14976,N_11699);
and U16339 (N_16339,N_14458,N_11769);
or U16340 (N_16340,N_11204,N_14734);
or U16341 (N_16341,N_11872,N_12294);
xor U16342 (N_16342,N_14764,N_14131);
and U16343 (N_16343,N_14491,N_12262);
nand U16344 (N_16344,N_12076,N_12658);
and U16345 (N_16345,N_13477,N_14056);
nor U16346 (N_16346,N_13268,N_11524);
nand U16347 (N_16347,N_11981,N_14407);
nand U16348 (N_16348,N_11670,N_14609);
nand U16349 (N_16349,N_14350,N_11386);
nor U16350 (N_16350,N_12148,N_13616);
or U16351 (N_16351,N_14206,N_13707);
and U16352 (N_16352,N_14428,N_10500);
or U16353 (N_16353,N_11924,N_11170);
and U16354 (N_16354,N_14361,N_13419);
and U16355 (N_16355,N_11474,N_12343);
or U16356 (N_16356,N_12582,N_14280);
or U16357 (N_16357,N_12236,N_11836);
nor U16358 (N_16358,N_13540,N_12428);
or U16359 (N_16359,N_13677,N_12764);
or U16360 (N_16360,N_11416,N_14365);
and U16361 (N_16361,N_11774,N_12938);
and U16362 (N_16362,N_13757,N_11102);
nand U16363 (N_16363,N_12668,N_13921);
nand U16364 (N_16364,N_13480,N_11374);
xor U16365 (N_16365,N_10273,N_13352);
nor U16366 (N_16366,N_14622,N_12083);
or U16367 (N_16367,N_10580,N_13750);
xnor U16368 (N_16368,N_11939,N_10053);
and U16369 (N_16369,N_10846,N_11507);
nor U16370 (N_16370,N_10084,N_10584);
and U16371 (N_16371,N_12976,N_14067);
nand U16372 (N_16372,N_14573,N_10127);
or U16373 (N_16373,N_14323,N_11327);
or U16374 (N_16374,N_14004,N_14700);
nor U16375 (N_16375,N_12693,N_11728);
and U16376 (N_16376,N_13016,N_12313);
xor U16377 (N_16377,N_10426,N_14989);
nor U16378 (N_16378,N_14699,N_14872);
xor U16379 (N_16379,N_14301,N_14827);
nand U16380 (N_16380,N_11341,N_10209);
or U16381 (N_16381,N_12295,N_11267);
and U16382 (N_16382,N_11260,N_12074);
nand U16383 (N_16383,N_14399,N_12370);
or U16384 (N_16384,N_11711,N_11379);
and U16385 (N_16385,N_11450,N_13375);
nand U16386 (N_16386,N_14371,N_13082);
or U16387 (N_16387,N_10929,N_10175);
nand U16388 (N_16388,N_14625,N_12604);
xor U16389 (N_16389,N_12716,N_13206);
nor U16390 (N_16390,N_13389,N_11760);
nor U16391 (N_16391,N_14490,N_11568);
xnor U16392 (N_16392,N_14416,N_12642);
and U16393 (N_16393,N_12900,N_12445);
or U16394 (N_16394,N_10358,N_12126);
or U16395 (N_16395,N_12687,N_12865);
or U16396 (N_16396,N_14595,N_11690);
and U16397 (N_16397,N_14648,N_10159);
nor U16398 (N_16398,N_13814,N_10516);
or U16399 (N_16399,N_11394,N_11570);
or U16400 (N_16400,N_10401,N_10093);
xnor U16401 (N_16401,N_12156,N_13347);
and U16402 (N_16402,N_11567,N_12705);
nand U16403 (N_16403,N_10541,N_14579);
nor U16404 (N_16404,N_14690,N_14298);
xnor U16405 (N_16405,N_12511,N_10157);
xor U16406 (N_16406,N_12571,N_12491);
or U16407 (N_16407,N_10540,N_11362);
nor U16408 (N_16408,N_11408,N_10315);
and U16409 (N_16409,N_11442,N_12023);
or U16410 (N_16410,N_10919,N_12468);
or U16411 (N_16411,N_11938,N_14908);
nor U16412 (N_16412,N_10221,N_10149);
nand U16413 (N_16413,N_11224,N_10297);
and U16414 (N_16414,N_10824,N_12954);
or U16415 (N_16415,N_12087,N_12003);
nand U16416 (N_16416,N_14830,N_12265);
and U16417 (N_16417,N_11283,N_10694);
nor U16418 (N_16418,N_13475,N_13145);
and U16419 (N_16419,N_10391,N_13882);
nor U16420 (N_16420,N_10072,N_13772);
or U16421 (N_16421,N_11764,N_14293);
or U16422 (N_16422,N_12794,N_12085);
xor U16423 (N_16423,N_14121,N_13416);
or U16424 (N_16424,N_13547,N_11633);
nand U16425 (N_16425,N_14408,N_11418);
and U16426 (N_16426,N_10408,N_12863);
or U16427 (N_16427,N_11968,N_13155);
and U16428 (N_16428,N_11182,N_10538);
xor U16429 (N_16429,N_10935,N_10787);
nand U16430 (N_16430,N_13020,N_13516);
nor U16431 (N_16431,N_10260,N_14877);
and U16432 (N_16432,N_11470,N_11492);
and U16433 (N_16433,N_14262,N_13586);
nand U16434 (N_16434,N_11234,N_11020);
or U16435 (N_16435,N_12815,N_13532);
nand U16436 (N_16436,N_12897,N_13018);
nor U16437 (N_16437,N_10069,N_11648);
xor U16438 (N_16438,N_11351,N_13941);
or U16439 (N_16439,N_10303,N_13503);
nor U16440 (N_16440,N_12544,N_12566);
nand U16441 (N_16441,N_13089,N_13213);
and U16442 (N_16442,N_14720,N_13713);
xor U16443 (N_16443,N_11056,N_11649);
nand U16444 (N_16444,N_12617,N_10276);
and U16445 (N_16445,N_14861,N_12224);
and U16446 (N_16446,N_10587,N_14449);
nor U16447 (N_16447,N_12437,N_10110);
nor U16448 (N_16448,N_10202,N_14456);
nand U16449 (N_16449,N_10842,N_10556);
nand U16450 (N_16450,N_13183,N_12312);
and U16451 (N_16451,N_12075,N_10518);
or U16452 (N_16452,N_13311,N_14073);
nor U16453 (N_16453,N_13434,N_10438);
nand U16454 (N_16454,N_14294,N_14924);
or U16455 (N_16455,N_10393,N_13856);
nand U16456 (N_16456,N_14108,N_14374);
and U16457 (N_16457,N_12868,N_11100);
xor U16458 (N_16458,N_12446,N_12778);
nand U16459 (N_16459,N_13726,N_13241);
nor U16460 (N_16460,N_11475,N_13910);
xnor U16461 (N_16461,N_11742,N_12904);
xnor U16462 (N_16462,N_14432,N_11579);
xnor U16463 (N_16463,N_10307,N_14275);
and U16464 (N_16464,N_13334,N_11637);
or U16465 (N_16465,N_11194,N_14156);
nor U16466 (N_16466,N_11427,N_12036);
xor U16467 (N_16467,N_10649,N_11074);
xnor U16468 (N_16468,N_10722,N_10885);
or U16469 (N_16469,N_10387,N_10272);
xor U16470 (N_16470,N_12365,N_12049);
nor U16471 (N_16471,N_14559,N_12635);
or U16472 (N_16472,N_13526,N_14684);
and U16473 (N_16473,N_12079,N_10107);
xor U16474 (N_16474,N_11501,N_11604);
xor U16475 (N_16475,N_10370,N_10310);
nand U16476 (N_16476,N_10466,N_13137);
nand U16477 (N_16477,N_10431,N_13966);
nor U16478 (N_16478,N_10443,N_10818);
xor U16479 (N_16479,N_11599,N_13203);
or U16480 (N_16480,N_13925,N_14202);
nor U16481 (N_16481,N_11375,N_10653);
xor U16482 (N_16482,N_11047,N_13028);
nand U16483 (N_16483,N_14001,N_13034);
xnor U16484 (N_16484,N_11240,N_10295);
xnor U16485 (N_16485,N_11003,N_11175);
nor U16486 (N_16486,N_13382,N_10480);
nand U16487 (N_16487,N_10444,N_10298);
xor U16488 (N_16488,N_10236,N_11496);
nor U16489 (N_16489,N_13536,N_11694);
nand U16490 (N_16490,N_11146,N_14196);
or U16491 (N_16491,N_13704,N_10076);
or U16492 (N_16492,N_13661,N_11134);
xnor U16493 (N_16493,N_14707,N_11245);
or U16494 (N_16494,N_10628,N_10593);
nor U16495 (N_16495,N_12095,N_14650);
or U16496 (N_16496,N_13187,N_10329);
and U16497 (N_16497,N_11389,N_11033);
xnor U16498 (N_16498,N_14745,N_12967);
nand U16499 (N_16499,N_12851,N_14317);
xnor U16500 (N_16500,N_12143,N_12955);
nand U16501 (N_16501,N_14724,N_13180);
or U16502 (N_16502,N_12908,N_14271);
xnor U16503 (N_16503,N_14019,N_11612);
nor U16504 (N_16504,N_12476,N_14713);
and U16505 (N_16505,N_12916,N_14095);
and U16506 (N_16506,N_12281,N_13531);
xnor U16507 (N_16507,N_11851,N_12496);
and U16508 (N_16508,N_12949,N_12345);
nand U16509 (N_16509,N_11201,N_14096);
and U16510 (N_16510,N_10816,N_11153);
and U16511 (N_16511,N_13388,N_11574);
and U16512 (N_16512,N_10763,N_10898);
xnor U16513 (N_16513,N_14651,N_13697);
or U16514 (N_16514,N_14630,N_13518);
nor U16515 (N_16515,N_14757,N_13997);
nor U16516 (N_16516,N_14571,N_12579);
nand U16517 (N_16517,N_13450,N_12960);
and U16518 (N_16518,N_11601,N_11066);
and U16519 (N_16519,N_11278,N_13201);
or U16520 (N_16520,N_10620,N_14655);
or U16521 (N_16521,N_10425,N_13417);
nand U16522 (N_16522,N_11429,N_10498);
xor U16523 (N_16523,N_14806,N_12178);
or U16524 (N_16524,N_13152,N_14679);
nand U16525 (N_16525,N_10189,N_12107);
xor U16526 (N_16526,N_10409,N_10124);
nor U16527 (N_16527,N_14532,N_12975);
nor U16528 (N_16528,N_10173,N_11972);
and U16529 (N_16529,N_13527,N_11449);
xnor U16530 (N_16530,N_14580,N_13307);
nand U16531 (N_16531,N_13191,N_11329);
or U16532 (N_16532,N_10246,N_10754);
xor U16533 (N_16533,N_13919,N_10974);
nand U16534 (N_16534,N_10915,N_10052);
nor U16535 (N_16535,N_13305,N_13887);
nand U16536 (N_16536,N_14472,N_14549);
or U16537 (N_16537,N_13656,N_12747);
nand U16538 (N_16538,N_14733,N_13130);
xor U16539 (N_16539,N_12840,N_10510);
or U16540 (N_16540,N_10549,N_13709);
and U16541 (N_16541,N_11594,N_14269);
xor U16542 (N_16542,N_10539,N_10768);
or U16543 (N_16543,N_11934,N_11754);
nand U16544 (N_16544,N_10971,N_14507);
nand U16545 (N_16545,N_12376,N_10081);
and U16546 (N_16546,N_13991,N_11645);
and U16547 (N_16547,N_12453,N_10457);
or U16548 (N_16548,N_14653,N_13598);
and U16549 (N_16549,N_10614,N_13552);
nand U16550 (N_16550,N_12789,N_13597);
and U16551 (N_16551,N_13083,N_10092);
and U16552 (N_16552,N_12246,N_12210);
or U16553 (N_16553,N_14222,N_13096);
or U16554 (N_16554,N_14938,N_12016);
nor U16555 (N_16555,N_12809,N_11390);
or U16556 (N_16556,N_13753,N_10112);
and U16557 (N_16557,N_12802,N_14771);
or U16558 (N_16558,N_10673,N_13650);
xor U16559 (N_16559,N_11221,N_10166);
and U16560 (N_16560,N_12110,N_14780);
nand U16561 (N_16561,N_10792,N_12248);
xor U16562 (N_16562,N_14719,N_13279);
and U16563 (N_16563,N_10125,N_13738);
nor U16564 (N_16564,N_12822,N_10101);
or U16565 (N_16565,N_14937,N_12741);
xor U16566 (N_16566,N_12254,N_13502);
xnor U16567 (N_16567,N_11502,N_13249);
xnor U16568 (N_16568,N_12634,N_13355);
or U16569 (N_16569,N_14422,N_12019);
xor U16570 (N_16570,N_12460,N_10250);
and U16571 (N_16571,N_13728,N_10688);
and U16572 (N_16572,N_10876,N_11828);
nor U16573 (N_16573,N_13567,N_11661);
nand U16574 (N_16574,N_13326,N_13575);
or U16575 (N_16575,N_12479,N_14118);
xnor U16576 (N_16576,N_10478,N_13138);
or U16577 (N_16577,N_12738,N_12198);
and U16578 (N_16578,N_10341,N_10138);
nor U16579 (N_16579,N_13631,N_10318);
nand U16580 (N_16580,N_14647,N_10997);
and U16581 (N_16581,N_13411,N_11488);
xor U16582 (N_16582,N_13077,N_14008);
xnor U16583 (N_16583,N_11290,N_14721);
or U16584 (N_16584,N_14341,N_14831);
xor U16585 (N_16585,N_14093,N_13636);
nor U16586 (N_16586,N_10275,N_14355);
nor U16587 (N_16587,N_12275,N_11481);
nor U16588 (N_16588,N_12414,N_14844);
xnor U16589 (N_16589,N_14649,N_12899);
and U16590 (N_16590,N_10698,N_10612);
xnor U16591 (N_16591,N_13698,N_13559);
or U16592 (N_16592,N_10532,N_12042);
nor U16593 (N_16593,N_11955,N_12878);
and U16594 (N_16594,N_10043,N_10572);
or U16595 (N_16595,N_12378,N_11108);
or U16596 (N_16596,N_13998,N_14977);
nor U16597 (N_16597,N_10835,N_11132);
and U16598 (N_16598,N_10198,N_14106);
xnor U16599 (N_16599,N_12602,N_11167);
xor U16600 (N_16600,N_10395,N_14218);
xnor U16601 (N_16601,N_12657,N_10581);
nand U16602 (N_16602,N_13052,N_12946);
nand U16603 (N_16603,N_11347,N_14489);
and U16604 (N_16604,N_11995,N_13926);
and U16605 (N_16605,N_13975,N_10557);
xor U16606 (N_16606,N_14024,N_14088);
nand U16607 (N_16607,N_11963,N_13857);
nor U16608 (N_16608,N_14793,N_11606);
and U16609 (N_16609,N_12585,N_14688);
xor U16610 (N_16610,N_13169,N_11627);
and U16611 (N_16611,N_14178,N_12507);
and U16612 (N_16612,N_10279,N_13504);
nor U16613 (N_16613,N_14087,N_12149);
or U16614 (N_16614,N_11426,N_11273);
xnor U16615 (N_16615,N_12788,N_12608);
nor U16616 (N_16616,N_13193,N_14461);
or U16617 (N_16617,N_10059,N_11176);
and U16618 (N_16618,N_11345,N_10019);
nand U16619 (N_16619,N_12044,N_10988);
nor U16620 (N_16620,N_14003,N_13031);
or U16621 (N_16621,N_10184,N_11155);
nor U16622 (N_16622,N_10899,N_13232);
nor U16623 (N_16623,N_11320,N_10266);
or U16624 (N_16624,N_13711,N_11393);
or U16625 (N_16625,N_11545,N_10829);
nand U16626 (N_16626,N_13584,N_13840);
nand U16627 (N_16627,N_12133,N_13960);
or U16628 (N_16628,N_12721,N_11726);
nand U16629 (N_16629,N_13055,N_11638);
nor U16630 (N_16630,N_13300,N_13790);
or U16631 (N_16631,N_13702,N_14785);
xnor U16632 (N_16632,N_11923,N_11266);
and U16633 (N_16633,N_12034,N_10617);
or U16634 (N_16634,N_10822,N_11614);
xor U16635 (N_16635,N_13920,N_12108);
nor U16636 (N_16636,N_13356,N_10452);
nor U16637 (N_16637,N_11806,N_14303);
or U16638 (N_16638,N_10741,N_12762);
or U16639 (N_16639,N_12820,N_14255);
nor U16640 (N_16640,N_13696,N_12554);
and U16641 (N_16641,N_14184,N_12685);
nand U16642 (N_16642,N_13344,N_11318);
xnor U16643 (N_16643,N_14726,N_14610);
and U16644 (N_16644,N_10253,N_14689);
or U16645 (N_16645,N_10781,N_13269);
and U16646 (N_16646,N_10927,N_13064);
or U16647 (N_16647,N_12380,N_13295);
nor U16648 (N_16648,N_14290,N_12774);
nand U16649 (N_16649,N_12613,N_12097);
nand U16650 (N_16650,N_14581,N_11913);
nor U16651 (N_16651,N_12690,N_12129);
nor U16652 (N_16652,N_11137,N_12818);
and U16653 (N_16653,N_10411,N_13784);
nor U16654 (N_16654,N_14400,N_12054);
and U16655 (N_16655,N_11597,N_14519);
or U16656 (N_16656,N_10326,N_13789);
nand U16657 (N_16657,N_13010,N_13819);
nand U16658 (N_16658,N_10287,N_14986);
nor U16659 (N_16659,N_10277,N_10594);
nor U16660 (N_16660,N_14235,N_12683);
nor U16661 (N_16661,N_11075,N_14100);
xor U16662 (N_16662,N_14256,N_11984);
and U16663 (N_16663,N_13091,N_11233);
xor U16664 (N_16664,N_11472,N_10980);
xnor U16665 (N_16665,N_13240,N_11101);
or U16666 (N_16666,N_14426,N_11900);
nand U16667 (N_16667,N_12810,N_11629);
nand U16668 (N_16668,N_10995,N_11659);
and U16669 (N_16669,N_14072,N_14348);
nor U16670 (N_16670,N_14154,N_14754);
nand U16671 (N_16671,N_12869,N_11652);
and U16672 (N_16672,N_12996,N_14716);
nor U16673 (N_16673,N_14081,N_10162);
or U16674 (N_16674,N_10317,N_13437);
nand U16675 (N_16675,N_10254,N_11626);
nand U16676 (N_16676,N_13294,N_14179);
nand U16677 (N_16677,N_11662,N_10379);
and U16678 (N_16678,N_13669,N_14959);
xor U16679 (N_16679,N_11438,N_10703);
nor U16680 (N_16680,N_11719,N_13592);
xnor U16681 (N_16681,N_13799,N_10759);
or U16682 (N_16682,N_12724,N_13635);
nor U16683 (N_16683,N_12017,N_10436);
nor U16684 (N_16684,N_10494,N_11380);
nor U16685 (N_16685,N_12122,N_11334);
or U16686 (N_16686,N_14708,N_14029);
nor U16687 (N_16687,N_12594,N_11988);
or U16688 (N_16688,N_10141,N_10843);
and U16689 (N_16689,N_12424,N_12777);
nand U16690 (N_16690,N_13467,N_14811);
nor U16691 (N_16691,N_14988,N_13632);
nand U16692 (N_16692,N_11025,N_11799);
or U16693 (N_16693,N_11994,N_14948);
nand U16694 (N_16694,N_11149,N_12387);
nor U16695 (N_16695,N_12616,N_10695);
or U16696 (N_16696,N_10777,N_10404);
nand U16697 (N_16697,N_11136,N_14036);
or U16698 (N_16698,N_12679,N_12972);
or U16699 (N_16699,N_11922,N_12039);
nand U16700 (N_16700,N_13736,N_10522);
nor U16701 (N_16701,N_10087,N_10939);
and U16702 (N_16702,N_13508,N_14890);
or U16703 (N_16703,N_10659,N_13285);
nand U16704 (N_16704,N_11206,N_12535);
xnor U16705 (N_16705,N_13854,N_14953);
or U16706 (N_16706,N_14666,N_13869);
nor U16707 (N_16707,N_14693,N_10877);
or U16708 (N_16708,N_11587,N_14966);
or U16709 (N_16709,N_13899,N_10743);
nand U16710 (N_16710,N_14822,N_13207);
nor U16711 (N_16711,N_11857,N_12072);
and U16712 (N_16712,N_10211,N_13189);
nand U16713 (N_16713,N_12933,N_12718);
nor U16714 (N_16714,N_13233,N_11902);
xnor U16715 (N_16715,N_12983,N_11855);
xnor U16716 (N_16716,N_14463,N_13959);
or U16717 (N_16717,N_14438,N_12520);
nand U16718 (N_16718,N_14297,N_11304);
nor U16719 (N_16719,N_13282,N_12711);
xnor U16720 (N_16720,N_14536,N_11550);
and U16721 (N_16721,N_12898,N_14962);
nand U16722 (N_16722,N_14820,N_14932);
nand U16723 (N_16723,N_12939,N_10449);
and U16724 (N_16724,N_14635,N_14904);
nand U16725 (N_16725,N_11499,N_14619);
nor U16726 (N_16726,N_12285,N_12681);
and U16727 (N_16727,N_11358,N_11706);
or U16728 (N_16728,N_11174,N_11852);
nand U16729 (N_16729,N_10897,N_11284);
xor U16730 (N_16730,N_12080,N_12093);
or U16731 (N_16731,N_10987,N_14758);
nand U16732 (N_16732,N_14928,N_10861);
nor U16733 (N_16733,N_11951,N_11651);
nor U16734 (N_16734,N_12227,N_14836);
nor U16735 (N_16735,N_13954,N_12880);
xnor U16736 (N_16736,N_13461,N_14706);
nor U16737 (N_16737,N_13397,N_13679);
xor U16738 (N_16738,N_10390,N_12628);
or U16739 (N_16739,N_12574,N_10569);
or U16740 (N_16740,N_10268,N_11603);
nand U16741 (N_16741,N_11163,N_10561);
or U16742 (N_16742,N_11983,N_10439);
nor U16743 (N_16743,N_10739,N_12940);
nand U16744 (N_16744,N_13905,N_11811);
nand U16745 (N_16745,N_10416,N_13866);
nor U16746 (N_16746,N_12720,N_13243);
and U16747 (N_16747,N_14372,N_10750);
nor U16748 (N_16748,N_10734,N_13298);
nand U16749 (N_16749,N_11298,N_14578);
and U16750 (N_16750,N_13585,N_13613);
or U16751 (N_16751,N_11641,N_10918);
and U16752 (N_16752,N_12059,N_13883);
xor U16753 (N_16753,N_11292,N_12859);
and U16754 (N_16754,N_12423,N_11122);
nor U16755 (N_16755,N_12499,N_13989);
xnor U16756 (N_16756,N_12400,N_11310);
nand U16757 (N_16757,N_14128,N_10872);
nand U16758 (N_16758,N_13945,N_11631);
nand U16759 (N_16759,N_11051,N_12856);
xor U16760 (N_16760,N_10886,N_10078);
nand U16761 (N_16761,N_11780,N_11624);
and U16762 (N_16762,N_12817,N_11441);
or U16763 (N_16763,N_14376,N_13297);
and U16764 (N_16764,N_12855,N_11162);
xor U16765 (N_16765,N_12027,N_10968);
and U16766 (N_16766,N_13988,N_11826);
xor U16767 (N_16767,N_12183,N_14327);
nor U16768 (N_16768,N_13990,N_14306);
xnor U16769 (N_16769,N_13638,N_11181);
nor U16770 (N_16770,N_13021,N_11809);
or U16771 (N_16771,N_13080,N_13538);
or U16772 (N_16772,N_13196,N_10916);
nand U16773 (N_16773,N_14346,N_13415);
xor U16774 (N_16774,N_11776,N_12816);
nor U16775 (N_16775,N_14208,N_10669);
and U16776 (N_16776,N_13332,N_10385);
xnor U16777 (N_16777,N_10945,N_14523);
nor U16778 (N_16778,N_12518,N_13795);
or U16779 (N_16779,N_10882,N_10720);
or U16780 (N_16780,N_13299,N_10574);
nor U16781 (N_16781,N_14562,N_10663);
nand U16782 (N_16782,N_14727,N_10881);
xor U16783 (N_16783,N_10732,N_13673);
nand U16784 (N_16784,N_14994,N_12303);
and U16785 (N_16785,N_14173,N_12031);
nor U16786 (N_16786,N_10989,N_10962);
nor U16787 (N_16787,N_14599,N_12966);
nor U16788 (N_16788,N_13291,N_13296);
xnor U16789 (N_16789,N_11620,N_14980);
nor U16790 (N_16790,N_13624,N_11868);
and U16791 (N_16791,N_11837,N_11746);
or U16792 (N_16792,N_12105,N_13306);
and U16793 (N_16793,N_12257,N_12314);
nand U16794 (N_16794,N_14175,N_10821);
and U16795 (N_16795,N_13012,N_13961);
and U16796 (N_16796,N_12412,N_11489);
xnor U16797 (N_16797,N_12587,N_12779);
and U16798 (N_16798,N_13877,N_13587);
nand U16799 (N_16799,N_10265,N_12229);
nand U16800 (N_16800,N_12147,N_14711);
xnor U16801 (N_16801,N_13835,N_13817);
and U16802 (N_16802,N_12643,N_11179);
and U16803 (N_16803,N_10578,N_12163);
nand U16804 (N_16804,N_14476,N_14577);
or U16805 (N_16805,N_10186,N_10033);
and U16806 (N_16806,N_14396,N_10049);
or U16807 (N_16807,N_13112,N_11498);
and U16808 (N_16808,N_13485,N_11200);
xnor U16809 (N_16809,N_10158,N_12339);
nand U16810 (N_16810,N_10521,N_13754);
nor U16811 (N_16811,N_11306,N_14138);
or U16812 (N_16812,N_13105,N_12676);
nand U16813 (N_16813,N_11976,N_14047);
or U16814 (N_16814,N_11065,N_12485);
xnor U16815 (N_16815,N_13374,N_14968);
nor U16816 (N_16816,N_10023,N_10106);
xor U16817 (N_16817,N_12390,N_14889);
and U16818 (N_16818,N_11998,N_12510);
and U16819 (N_16819,N_10953,N_12411);
and U16820 (N_16820,N_12965,N_11445);
or U16821 (N_16821,N_10803,N_11191);
xor U16822 (N_16822,N_14728,N_14481);
nand U16823 (N_16823,N_13110,N_13358);
xnor U16824 (N_16824,N_12493,N_14145);
or U16825 (N_16825,N_13117,N_12689);
nor U16826 (N_16826,N_11326,N_10772);
or U16827 (N_16827,N_12701,N_10192);
nand U16828 (N_16828,N_14039,N_10038);
xor U16829 (N_16829,N_14278,N_14564);
nand U16830 (N_16830,N_13395,N_13943);
or U16831 (N_16831,N_12355,N_13637);
and U16832 (N_16832,N_12368,N_11647);
xor U16833 (N_16833,N_14818,N_13157);
and U16834 (N_16834,N_10871,N_11286);
xnor U16835 (N_16835,N_10998,N_14395);
nor U16836 (N_16836,N_13756,N_14236);
and U16837 (N_16837,N_13699,N_11026);
or U16838 (N_16838,N_11062,N_11654);
xor U16839 (N_16839,N_12828,N_10573);
or U16840 (N_16840,N_11818,N_12606);
or U16841 (N_16841,N_12347,N_13050);
nand U16842 (N_16842,N_10802,N_12444);
nand U16843 (N_16843,N_14946,N_10936);
or U16844 (N_16844,N_14150,N_11357);
nor U16845 (N_16845,N_14427,N_14961);
xnor U16846 (N_16846,N_13440,N_11085);
nand U16847 (N_16847,N_14542,N_12512);
and U16848 (N_16848,N_12384,N_14743);
nand U16849 (N_16849,N_11534,N_12957);
or U16850 (N_16850,N_11677,N_13758);
and U16851 (N_16851,N_11422,N_12505);
or U16852 (N_16852,N_10746,N_12710);
xnor U16853 (N_16853,N_11925,N_12937);
or U16854 (N_16854,N_13413,N_11384);
xor U16855 (N_16855,N_12443,N_13509);
nor U16856 (N_16856,N_13455,N_10657);
nor U16857 (N_16857,N_11558,N_10869);
nand U16858 (N_16858,N_10467,N_11713);
nor U16859 (N_16859,N_14952,N_13484);
nor U16860 (N_16860,N_10245,N_10427);
xnor U16861 (N_16861,N_11242,N_11896);
and U16862 (N_16862,N_14598,N_11536);
xnor U16863 (N_16863,N_12214,N_14865);
nand U16864 (N_16864,N_13181,N_14204);
xor U16865 (N_16865,N_14746,N_13649);
xor U16866 (N_16866,N_14633,N_11325);
or U16867 (N_16867,N_12846,N_10036);
and U16868 (N_16868,N_10512,N_13978);
and U16869 (N_16869,N_14777,N_10131);
nor U16870 (N_16870,N_14319,N_10207);
nand U16871 (N_16871,N_13025,N_12763);
nand U16872 (N_16872,N_11887,N_10723);
xnor U16873 (N_16873,N_13769,N_12463);
xor U16874 (N_16874,N_14993,N_12569);
nor U16875 (N_16875,N_12113,N_14125);
nand U16876 (N_16876,N_14511,N_11227);
xnor U16877 (N_16877,N_10111,N_11908);
or U16878 (N_16878,N_10786,N_13888);
and U16879 (N_16879,N_13551,N_10931);
or U16880 (N_16880,N_11103,N_13972);
or U16881 (N_16881,N_11971,N_14548);
or U16882 (N_16882,N_13590,N_10117);
xor U16883 (N_16883,N_13965,N_13520);
or U16884 (N_16884,N_14620,N_14498);
or U16885 (N_16885,N_14314,N_14514);
nor U16886 (N_16886,N_12187,N_14969);
or U16887 (N_16887,N_12981,N_10073);
and U16888 (N_16888,N_11052,N_12572);
or U16889 (N_16889,N_12426,N_11484);
xnor U16890 (N_16890,N_11505,N_12179);
nor U16891 (N_16891,N_13258,N_10343);
or U16892 (N_16892,N_11480,N_11487);
nand U16893 (N_16893,N_14783,N_10417);
or U16894 (N_16894,N_13217,N_10199);
nor U16895 (N_16895,N_11725,N_13820);
and U16896 (N_16896,N_10461,N_14933);
nand U16897 (N_16897,N_11282,N_11623);
nor U16898 (N_16898,N_13640,N_12743);
xnor U16899 (N_16899,N_13904,N_14083);
nand U16900 (N_16900,N_12020,N_14979);
nand U16901 (N_16901,N_14232,N_10397);
or U16902 (N_16902,N_11027,N_10800);
or U16903 (N_16903,N_12508,N_14124);
nor U16904 (N_16904,N_14732,N_12251);
and U16905 (N_16905,N_12277,N_13340);
xnor U16906 (N_16906,N_11239,N_13672);
nand U16907 (N_16907,N_10301,N_10999);
xnor U16908 (N_16908,N_14313,N_12369);
nand U16909 (N_16909,N_13879,N_11595);
nor U16910 (N_16910,N_12986,N_14366);
nor U16911 (N_16911,N_13571,N_10374);
and U16912 (N_16912,N_11762,N_10497);
nor U16913 (N_16913,N_12357,N_11724);
or U16914 (N_16914,N_10858,N_14632);
xnor U16915 (N_16915,N_11845,N_13120);
and U16916 (N_16916,N_12953,N_12752);
xnor U16917 (N_16917,N_11632,N_13628);
or U16918 (N_16918,N_10542,N_11617);
nor U16919 (N_16919,N_10259,N_11324);
or U16920 (N_16920,N_14068,N_10291);
or U16921 (N_16921,N_12527,N_12441);
and U16922 (N_16922,N_12011,N_11141);
nand U16923 (N_16923,N_10346,N_13745);
nor U16924 (N_16924,N_13222,N_12803);
nand U16925 (N_16925,N_12467,N_10377);
and U16926 (N_16926,N_14483,N_14054);
and U16927 (N_16927,N_13459,N_10247);
xor U16928 (N_16928,N_11940,N_10029);
nor U16929 (N_16929,N_12910,N_11354);
xor U16930 (N_16930,N_10160,N_14787);
nand U16931 (N_16931,N_12997,N_12048);
nand U16932 (N_16932,N_11991,N_13481);
nor U16933 (N_16933,N_12451,N_10062);
or U16934 (N_16934,N_12702,N_10095);
nand U16935 (N_16935,N_13147,N_12761);
and U16936 (N_16936,N_10856,N_14715);
xor U16937 (N_16937,N_10314,N_11783);
nor U16938 (N_16938,N_10181,N_11681);
nand U16939 (N_16939,N_13932,N_12620);
nand U16940 (N_16940,N_12471,N_13185);
nor U16941 (N_16941,N_11691,N_12142);
or U16942 (N_16942,N_13220,N_14230);
or U16943 (N_16943,N_11683,N_11943);
nor U16944 (N_16944,N_14250,N_11369);
or U16945 (N_16945,N_11765,N_13838);
nor U16946 (N_16946,N_13647,N_14496);
nand U16947 (N_16947,N_11316,N_12837);
nand U16948 (N_16948,N_11937,N_14875);
nand U16949 (N_16949,N_14155,N_12737);
and U16950 (N_16950,N_10089,N_10350);
nand U16951 (N_16951,N_14934,N_12350);
xor U16952 (N_16952,N_12845,N_12375);
or U16953 (N_16953,N_10001,N_12874);
or U16954 (N_16954,N_14228,N_11041);
xor U16955 (N_16955,N_13985,N_13168);
nor U16956 (N_16956,N_10284,N_11166);
or U16957 (N_16957,N_11187,N_13143);
nor U16958 (N_16958,N_11451,N_10674);
nand U16959 (N_16959,N_14910,N_12660);
and U16960 (N_16960,N_14284,N_13862);
nand U16961 (N_16961,N_14869,N_10176);
and U16962 (N_16962,N_11177,N_13729);
or U16963 (N_16963,N_14710,N_14807);
or U16964 (N_16964,N_14248,N_11186);
nor U16965 (N_16965,N_11192,N_12621);
or U16966 (N_16966,N_11236,N_10635);
or U16967 (N_16967,N_12482,N_13603);
or U16968 (N_16968,N_11885,N_14654);
nand U16969 (N_16969,N_11486,N_10108);
and U16970 (N_16970,N_11856,N_14891);
and U16971 (N_16971,N_13447,N_10637);
xor U16972 (N_16972,N_10367,N_10708);
xor U16973 (N_16973,N_14477,N_14762);
and U16974 (N_16974,N_10545,N_11293);
or U16975 (N_16975,N_11560,N_11067);
nand U16976 (N_16976,N_12915,N_12388);
nand U16977 (N_16977,N_10701,N_14129);
nand U16978 (N_16978,N_11049,N_13654);
nand U16979 (N_16979,N_10533,N_10854);
or U16980 (N_16980,N_11551,N_11419);
and U16981 (N_16981,N_12297,N_14055);
nand U16982 (N_16982,N_14246,N_11784);
and U16983 (N_16983,N_13562,N_11199);
nand U16984 (N_16984,N_10400,N_12707);
xnor U16985 (N_16985,N_10477,N_11321);
xor U16986 (N_16986,N_13741,N_11211);
or U16987 (N_16987,N_14943,N_12213);
xnor U16988 (N_16988,N_13462,N_13390);
nand U16989 (N_16989,N_11695,N_14444);
nor U16990 (N_16990,N_13622,N_13950);
and U16991 (N_16991,N_13914,N_13724);
xor U16992 (N_16992,N_13248,N_14798);
and U16993 (N_16993,N_10305,N_10191);
and U16994 (N_16994,N_14194,N_10150);
nor U16995 (N_16995,N_11081,N_14945);
nor U16996 (N_16996,N_10793,N_10294);
xnor U16997 (N_16997,N_13182,N_11679);
or U16998 (N_16998,N_10338,N_12834);
xor U16999 (N_16999,N_12131,N_12152);
nor U17000 (N_17000,N_10000,N_14084);
xor U17001 (N_17001,N_12633,N_14181);
nand U17002 (N_17002,N_13043,N_11319);
or U17003 (N_17003,N_11437,N_13436);
nor U17004 (N_17004,N_14823,N_11263);
and U17005 (N_17005,N_12269,N_12717);
and U17006 (N_17006,N_14137,N_11238);
xnor U17007 (N_17007,N_13056,N_14025);
or U17008 (N_17008,N_10526,N_12603);
or U17009 (N_17009,N_10509,N_10468);
nand U17010 (N_17010,N_12666,N_14842);
nand U17011 (N_17011,N_12171,N_12010);
nand U17012 (N_17012,N_12167,N_14276);
xnor U17013 (N_17013,N_14612,N_11152);
nor U17014 (N_17014,N_12667,N_10351);
xnor U17015 (N_17015,N_13079,N_14146);
nor U17016 (N_17016,N_14530,N_14495);
xnor U17017 (N_17017,N_14011,N_11858);
nor U17018 (N_17018,N_14274,N_12474);
and U17019 (N_17019,N_14112,N_12969);
nor U17020 (N_17020,N_13846,N_14939);
xor U17021 (N_17021,N_11970,N_11129);
nand U17022 (N_17022,N_11302,N_11891);
and U17023 (N_17023,N_12128,N_11533);
and U17024 (N_17024,N_11436,N_10249);
or U17025 (N_17025,N_14387,N_13014);
or U17026 (N_17026,N_14944,N_11519);
nor U17027 (N_17027,N_10233,N_10376);
xnor U17028 (N_17028,N_14281,N_12151);
and U17029 (N_17029,N_12250,N_12117);
nand U17030 (N_17030,N_13970,N_11792);
nand U17031 (N_17031,N_10796,N_14895);
and U17032 (N_17032,N_11960,N_14425);
and U17033 (N_17033,N_12492,N_13449);
and U17034 (N_17034,N_12644,N_13855);
xnor U17035 (N_17035,N_12078,N_14209);
or U17036 (N_17036,N_10941,N_10145);
nand U17037 (N_17037,N_12853,N_11554);
nor U17038 (N_17038,N_10938,N_12756);
or U17039 (N_17039,N_12696,N_12894);
nand U17040 (N_17040,N_14234,N_12524);
nand U17041 (N_17041,N_10624,N_13831);
or U17042 (N_17042,N_12517,N_11285);
and U17043 (N_17043,N_13642,N_12570);
xnor U17044 (N_17044,N_13977,N_13667);
nor U17045 (N_17045,N_12991,N_14921);
nor U17046 (N_17046,N_12727,N_11232);
nor U17047 (N_17047,N_13006,N_13148);
or U17048 (N_17048,N_10206,N_12483);
xnor U17049 (N_17049,N_13359,N_12550);
and U17050 (N_17050,N_12848,N_14016);
and U17051 (N_17051,N_10760,N_14747);
nand U17052 (N_17052,N_10840,N_11078);
nor U17053 (N_17053,N_11068,N_10682);
nor U17054 (N_17054,N_12302,N_14858);
nand U17055 (N_17055,N_11848,N_14171);
or U17056 (N_17056,N_11280,N_11841);
nor U17057 (N_17057,N_11822,N_10210);
and U17058 (N_17058,N_13849,N_13231);
nand U17059 (N_17059,N_13717,N_12640);
nor U17060 (N_17060,N_12539,N_14813);
nand U17061 (N_17061,N_14134,N_12104);
or U17062 (N_17062,N_12292,N_13675);
nand U17063 (N_17063,N_13751,N_13563);
or U17064 (N_17064,N_11834,N_11807);
and U17065 (N_17065,N_12287,N_12682);
nand U17066 (N_17066,N_11252,N_10080);
and U17067 (N_17067,N_14132,N_12037);
nand U17068 (N_17068,N_11082,N_13593);
xnor U17069 (N_17069,N_10299,N_13517);
or U17070 (N_17070,N_13367,N_11790);
xnor U17071 (N_17071,N_14626,N_13133);
xnor U17072 (N_17072,N_14092,N_14240);
or U17073 (N_17073,N_14401,N_10841);
xor U17074 (N_17074,N_12332,N_10626);
xnor U17075 (N_17075,N_10026,N_12592);
nand U17076 (N_17076,N_13755,N_13212);
and U17077 (N_17077,N_12557,N_10984);
nand U17078 (N_17078,N_13744,N_13160);
xnor U17079 (N_17079,N_14338,N_14614);
nand U17080 (N_17080,N_14447,N_13604);
nand U17081 (N_17081,N_13625,N_12931);
and U17082 (N_17082,N_11168,N_12342);
xnor U17083 (N_17083,N_12238,N_12831);
nor U17084 (N_17084,N_10853,N_12308);
and U17085 (N_17085,N_11116,N_14663);
nand U17086 (N_17086,N_12857,N_12276);
nand U17087 (N_17087,N_11107,N_12573);
xor U17088 (N_17088,N_12073,N_11453);
and U17089 (N_17089,N_11363,N_14833);
xnor U17090 (N_17090,N_13911,N_14005);
nand U17091 (N_17091,N_12158,N_11212);
xnor U17092 (N_17092,N_11314,N_12581);
nand U17093 (N_17093,N_10197,N_10208);
and U17094 (N_17094,N_11355,N_14434);
or U17095 (N_17095,N_14078,N_11032);
or U17096 (N_17096,N_12300,N_10588);
xnor U17097 (N_17097,N_11985,N_11054);
or U17098 (N_17098,N_14486,N_13834);
and U17099 (N_17099,N_14926,N_10232);
and U17100 (N_17100,N_12066,N_12713);
or U17101 (N_17101,N_10267,N_13558);
and U17102 (N_17102,N_12317,N_13912);
nor U17103 (N_17103,N_14045,N_10104);
nor U17104 (N_17104,N_13565,N_10152);
or U17105 (N_17105,N_10742,N_12835);
xnor U17106 (N_17106,N_14023,N_13568);
or U17107 (N_17107,N_14133,N_14901);
or U17108 (N_17108,N_13409,N_10707);
nor U17109 (N_17109,N_13892,N_12703);
xnor U17110 (N_17110,N_10178,N_14555);
and U17111 (N_17111,N_12065,N_12782);
or U17112 (N_17112,N_13623,N_12615);
nor U17113 (N_17113,N_13310,N_12209);
and U17114 (N_17114,N_13591,N_10304);
nor U17115 (N_17115,N_11259,N_12584);
or U17116 (N_17116,N_11801,N_14415);
nor U17117 (N_17117,N_14390,N_13860);
nor U17118 (N_17118,N_10761,N_10484);
or U17119 (N_17119,N_14709,N_13749);
xnor U17120 (N_17120,N_10586,N_12656);
and U17121 (N_17121,N_13161,N_10479);
nor U17122 (N_17122,N_12361,N_13705);
nor U17123 (N_17123,N_10414,N_13955);
xor U17124 (N_17124,N_13530,N_13071);
nor U17125 (N_17125,N_14252,N_11404);
xnor U17126 (N_17126,N_12457,N_10926);
and U17127 (N_17127,N_11276,N_12824);
and U17128 (N_17128,N_11786,N_10932);
or U17129 (N_17129,N_12698,N_14226);
xor U17130 (N_17130,N_14044,N_10833);
or U17131 (N_17131,N_13438,N_12177);
or U17132 (N_17132,N_13330,N_10195);
or U17133 (N_17133,N_11803,N_11043);
xnor U17134 (N_17134,N_13937,N_14200);
and U17135 (N_17135,N_14522,N_13474);
nand U17136 (N_17136,N_14575,N_10064);
and U17137 (N_17137,N_13548,N_10860);
and U17138 (N_17138,N_11722,N_14894);
nor U17139 (N_17139,N_10655,N_11921);
or U17140 (N_17140,N_14766,N_12201);
nor U17141 (N_17141,N_12605,N_10063);
and U17142 (N_17142,N_11863,N_11873);
nor U17143 (N_17143,N_14884,N_13423);
xnor U17144 (N_17144,N_13969,N_14090);
or U17145 (N_17145,N_14040,N_13714);
and U17146 (N_17146,N_12207,N_12650);
or U17147 (N_17147,N_10798,N_10752);
nand U17148 (N_17148,N_13124,N_14856);
nand U17149 (N_17149,N_13602,N_13122);
nand U17150 (N_17150,N_10644,N_14501);
nand U17151 (N_17151,N_13199,N_13190);
xnor U17152 (N_17152,N_13159,N_13230);
nor U17153 (N_17153,N_12497,N_14107);
nor U17154 (N_17154,N_11556,N_10805);
xor U17155 (N_17155,N_13903,N_14354);
nor U17156 (N_17156,N_14379,N_10511);
and U17157 (N_17157,N_14883,N_12422);
and U17158 (N_17158,N_11682,N_10726);
nor U17159 (N_17159,N_10652,N_14048);
nor U17160 (N_17160,N_14682,N_14668);
and U17161 (N_17161,N_10530,N_13141);
or U17162 (N_17162,N_13742,N_10201);
nand U17163 (N_17163,N_11096,N_13208);
xor U17164 (N_17164,N_11151,N_12610);
nor U17165 (N_17165,N_11012,N_11147);
nor U17166 (N_17166,N_10775,N_13507);
nor U17167 (N_17167,N_10451,N_13962);
xor U17168 (N_17168,N_13116,N_11978);
nand U17169 (N_17169,N_12870,N_11112);
xnor U17170 (N_17170,N_11335,N_11514);
nor U17171 (N_17171,N_14356,N_13767);
nor U17172 (N_17172,N_13486,N_11063);
nand U17173 (N_17173,N_12190,N_11588);
or U17174 (N_17174,N_13723,N_12353);
nor U17175 (N_17175,N_12586,N_14160);
xnor U17176 (N_17176,N_14906,N_10174);
nor U17177 (N_17177,N_14500,N_12215);
nand U17178 (N_17178,N_11898,N_12125);
nand U17179 (N_17179,N_14080,N_13488);
or U17180 (N_17180,N_14473,N_10165);
xor U17181 (N_17181,N_11251,N_12330);
nand U17182 (N_17182,N_13387,N_11933);
or U17183 (N_17183,N_14857,N_11440);
or U17184 (N_17184,N_11268,N_13561);
nor U17185 (N_17185,N_11747,N_14411);
nor U17186 (N_17186,N_11569,N_13194);
nor U17187 (N_17187,N_10570,N_14832);
xnor U17188 (N_17188,N_13019,N_10873);
and U17189 (N_17189,N_12985,N_13822);
nor U17190 (N_17190,N_14479,N_10766);
xnor U17191 (N_17191,N_10167,N_13871);
xor U17192 (N_17192,N_12472,N_10241);
or U17193 (N_17193,N_12120,N_10487);
and U17194 (N_17194,N_14017,N_11665);
and U17195 (N_17195,N_13132,N_12286);
nand U17196 (N_17196,N_12609,N_11589);
and U17197 (N_17197,N_10386,N_11461);
or U17198 (N_17198,N_10491,N_12252);
xor U17199 (N_17199,N_11296,N_12984);
nand U17200 (N_17200,N_12814,N_14880);
nand U17201 (N_17201,N_14540,N_14616);
or U17202 (N_17202,N_10394,N_14186);
or U17203 (N_17203,N_13273,N_12461);
nor U17204 (N_17204,N_10951,N_13106);
and U17205 (N_17205,N_10646,N_10282);
nor U17206 (N_17206,N_12220,N_10656);
xnor U17207 (N_17207,N_12598,N_12239);
and U17208 (N_17208,N_12797,N_11373);
and U17209 (N_17209,N_11804,N_12268);
nand U17210 (N_17210,N_13942,N_12372);
and U17211 (N_17211,N_12731,N_13895);
xnor U17212 (N_17212,N_12858,N_12005);
xnor U17213 (N_17213,N_14406,N_12200);
and U17214 (N_17214,N_14779,N_14499);
nand U17215 (N_17215,N_12796,N_11447);
or U17216 (N_17216,N_11920,N_11975);
or U17217 (N_17217,N_14950,N_14524);
xor U17218 (N_17218,N_12235,N_12231);
xor U17219 (N_17219,N_10683,N_13290);
nand U17220 (N_17220,N_13752,N_13008);
or U17221 (N_17221,N_10333,N_11862);
or U17222 (N_17222,N_10369,N_14845);
nor U17223 (N_17223,N_14471,N_14027);
and U17224 (N_17224,N_10762,N_10765);
nand U17225 (N_17225,N_10103,N_14694);
or U17226 (N_17226,N_11897,N_11337);
nor U17227 (N_17227,N_12607,N_14607);
nand U17228 (N_17228,N_10596,N_14460);
xnor U17229 (N_17229,N_13556,N_11089);
or U17230 (N_17230,N_12694,N_11917);
or U17231 (N_17231,N_12240,N_13553);
nor U17232 (N_17232,N_11840,N_10525);
or U17233 (N_17233,N_13917,N_13167);
nor U17234 (N_17234,N_12928,N_13648);
and U17235 (N_17235,N_11552,N_13223);
xor U17236 (N_17236,N_12322,N_10340);
xnor U17237 (N_17237,N_12094,N_11339);
or U17238 (N_17238,N_12274,N_14312);
nand U17239 (N_17239,N_11996,N_14007);
nor U17240 (N_17240,N_14761,N_14873);
and U17241 (N_17241,N_11261,N_14330);
nor U17242 (N_17242,N_10687,N_10566);
and U17243 (N_17243,N_10354,N_14656);
or U17244 (N_17244,N_10476,N_10188);
nor U17245 (N_17245,N_11145,N_12168);
xnor U17246 (N_17246,N_14070,N_11952);
nand U17247 (N_17247,N_11884,N_10524);
or U17248 (N_17248,N_13000,N_13251);
nor U17249 (N_17249,N_12680,N_11016);
nor U17250 (N_17250,N_12040,N_13335);
xnor U17251 (N_17251,N_12271,N_10618);
nand U17252 (N_17252,N_13629,N_13768);
nor U17253 (N_17253,N_12993,N_14791);
or U17254 (N_17254,N_11745,N_10300);
nand U17255 (N_17255,N_10531,N_12921);
or U17256 (N_17256,N_11246,N_11881);
xnor U17257 (N_17257,N_11866,N_14267);
nor U17258 (N_17258,N_13345,N_14097);
nor U17259 (N_17259,N_12599,N_14629);
nand U17260 (N_17260,N_12700,N_14360);
or U17261 (N_17261,N_11564,N_13843);
or U17262 (N_17262,N_11364,N_12464);
or U17263 (N_17263,N_14886,N_10285);
and U17264 (N_17264,N_12791,N_12494);
xor U17265 (N_17265,N_11892,N_12891);
xnor U17266 (N_17266,N_10864,N_12056);
nor U17267 (N_17267,N_13579,N_11039);
nor U17268 (N_17268,N_11000,N_12886);
nor U17269 (N_17269,N_11797,N_11580);
or U17270 (N_17270,N_13076,N_13029);
nor U17271 (N_17271,N_12930,N_14166);
or U17272 (N_17272,N_14358,N_11410);
xnor U17273 (N_17273,N_13824,N_14646);
and U17274 (N_17274,N_14911,N_12319);
or U17275 (N_17275,N_12936,N_10717);
xor U17276 (N_17276,N_13393,N_13529);
and U17277 (N_17277,N_12121,N_14257);
nor U17278 (N_17278,N_14367,N_10874);
xnor U17279 (N_17279,N_14992,N_10488);
nor U17280 (N_17280,N_13938,N_11666);
nand U17281 (N_17281,N_14203,N_13097);
or U17282 (N_17282,N_11957,N_12419);
and U17283 (N_17283,N_11160,N_13354);
and U17284 (N_17284,N_14835,N_13659);
and U17285 (N_17285,N_10622,N_11333);
and U17286 (N_17286,N_12826,N_11870);
or U17287 (N_17287,N_13875,N_10875);
or U17288 (N_17288,N_11225,N_12978);
nor U17289 (N_17289,N_11371,N_12673);
and U17290 (N_17290,N_10575,N_10248);
or U17291 (N_17291,N_14332,N_11079);
and U17292 (N_17292,N_11300,N_14326);
nand U17293 (N_17293,N_10776,N_11409);
nand U17294 (N_17294,N_10585,N_12022);
xor U17295 (N_17295,N_11544,N_14457);
nor U17296 (N_17296,N_13878,N_14692);
nand U17297 (N_17297,N_14421,N_12649);
nor U17298 (N_17298,N_10364,N_14063);
or U17299 (N_17299,N_13309,N_10434);
or U17300 (N_17300,N_14331,N_10050);
nor U17301 (N_17301,N_10281,N_13798);
nor U17302 (N_17302,N_14140,N_13646);
xor U17303 (N_17303,N_14967,N_12902);
xor U17304 (N_17304,N_12406,N_10648);
nor U17305 (N_17305,N_12811,N_10623);
or U17306 (N_17306,N_13341,N_12829);
nor U17307 (N_17307,N_14264,N_12688);
xor U17308 (N_17308,N_13703,N_10564);
or U17309 (N_17309,N_13609,N_10880);
or U17310 (N_17310,N_12061,N_12416);
and U17311 (N_17311,N_14197,N_11042);
or U17312 (N_17312,N_14512,N_10888);
nor U17313 (N_17313,N_14552,N_14803);
xor U17314 (N_17314,N_11264,N_11207);
and U17315 (N_17315,N_14929,N_10205);
nand U17316 (N_17316,N_13791,N_14701);
and U17317 (N_17317,N_11773,N_11997);
and U17318 (N_17318,N_14413,N_12484);
or U17319 (N_17319,N_14192,N_13643);
or U17320 (N_17320,N_12060,N_14273);
xnor U17321 (N_17321,N_14439,N_11553);
xnor U17322 (N_17322,N_14896,N_13432);
nor U17323 (N_17323,N_11126,N_14698);
nand U17324 (N_17324,N_12256,N_10463);
xor U17325 (N_17325,N_13275,N_11035);
and U17326 (N_17326,N_14272,N_13158);
xnor U17327 (N_17327,N_14295,N_11158);
nand U17328 (N_17328,N_11208,N_13135);
xnor U17329 (N_17329,N_11478,N_13765);
nand U17330 (N_17330,N_12208,N_12038);
xor U17331 (N_17331,N_13927,N_10665);
and U17332 (N_17332,N_14867,N_10702);
and U17333 (N_17333,N_11789,N_12890);
or U17334 (N_17334,N_11024,N_12071);
nand U17335 (N_17335,N_10684,N_12266);
nand U17336 (N_17336,N_12854,N_11381);
nand U17337 (N_17337,N_13452,N_11517);
or U17338 (N_17338,N_10753,N_12733);
or U17339 (N_17339,N_10555,N_10611);
or U17340 (N_17340,N_10177,N_11520);
and U17341 (N_17341,N_11377,N_11982);
xnor U17342 (N_17342,N_14033,N_11798);
nand U17343 (N_17343,N_11330,N_12684);
xor U17344 (N_17344,N_14600,N_11615);
and U17345 (N_17345,N_10878,N_11927);
nor U17346 (N_17346,N_11861,N_12475);
and U17347 (N_17347,N_12430,N_12099);
nand U17348 (N_17348,N_13277,N_11391);
or U17349 (N_17349,N_11443,N_10603);
xor U17350 (N_17350,N_13035,N_12672);
and U17351 (N_17351,N_11061,N_11072);
nand U17352 (N_17352,N_14664,N_11930);
or U17353 (N_17353,N_13743,N_14006);
xor U17354 (N_17354,N_10922,N_10008);
or U17355 (N_17355,N_14182,N_12625);
xnor U17356 (N_17356,N_13204,N_13655);
nor U17357 (N_17357,N_14241,N_11269);
nor U17358 (N_17358,N_14377,N_13027);
xnor U17359 (N_17359,N_12336,N_11710);
nand U17360 (N_17360,N_14012,N_11277);
or U17361 (N_17361,N_10482,N_12166);
or U17362 (N_17362,N_14585,N_11456);
xnor U17363 (N_17363,N_13615,N_10337);
nand U17364 (N_17364,N_14768,N_10952);
nor U17365 (N_17365,N_14541,N_10362);
or U17366 (N_17366,N_10071,N_14725);
and U17367 (N_17367,N_11189,N_14013);
or U17368 (N_17368,N_13916,N_14041);
nor U17369 (N_17369,N_10529,N_12784);
and U17370 (N_17370,N_10363,N_12433);
and U17371 (N_17371,N_11231,N_14975);
and U17372 (N_17372,N_13466,N_13544);
nor U17373 (N_17373,N_10852,N_12260);
nor U17374 (N_17374,N_12726,N_13607);
or U17375 (N_17375,N_14972,N_12442);
nor U17376 (N_17376,N_14513,N_11406);
nand U17377 (N_17377,N_14172,N_10681);
nor U17378 (N_17378,N_14383,N_14309);
nand U17379 (N_17379,N_13906,N_11095);
xnor U17380 (N_17380,N_14435,N_12735);
or U17381 (N_17381,N_12337,N_10074);
nor U17382 (N_17382,N_11516,N_14050);
xnor U17383 (N_17383,N_11853,N_10799);
nor U17384 (N_17384,N_13445,N_12988);
or U17385 (N_17385,N_10420,N_13037);
nor U17386 (N_17386,N_10544,N_11899);
or U17387 (N_17387,N_11387,N_11915);
nand U17388 (N_17388,N_14020,N_11142);
or U17389 (N_17389,N_13747,N_11918);
xnor U17390 (N_17390,N_13573,N_12145);
xnor U17391 (N_17391,N_13976,N_14110);
xnor U17392 (N_17392,N_14637,N_12175);
nor U17393 (N_17393,N_12394,N_10608);
nand U17394 (N_17394,N_14031,N_12141);
nor U17395 (N_17395,N_14176,N_10290);
xnor U17396 (N_17396,N_12340,N_12567);
nor U17397 (N_17397,N_11086,N_10193);
or U17398 (N_17398,N_11753,N_13982);
xor U17399 (N_17399,N_13317,N_14557);
xnor U17400 (N_17400,N_12704,N_11220);
nor U17401 (N_17401,N_13011,N_13378);
xnor U17402 (N_17402,N_12386,N_12184);
xnor U17403 (N_17403,N_13816,N_13420);
and U17404 (N_17404,N_10244,N_14163);
and U17405 (N_17405,N_12611,N_14973);
and U17406 (N_17406,N_13865,N_14618);
xnor U17407 (N_17407,N_11675,N_14242);
xor U17408 (N_17408,N_11328,N_14864);
nor U17409 (N_17409,N_14819,N_10200);
and U17410 (N_17410,N_13570,N_13694);
nor U17411 (N_17411,N_13907,N_10446);
or U17412 (N_17412,N_14344,N_12429);
nor U17413 (N_17413,N_11295,N_12320);
or U17414 (N_17414,N_11825,N_12228);
or U17415 (N_17415,N_11139,N_13195);
xnor U17416 (N_17416,N_10010,N_14504);
nor U17417 (N_17417,N_13121,N_11023);
and U17418 (N_17418,N_11557,N_10057);
or U17419 (N_17419,N_11040,N_10863);
or U17420 (N_17420,N_14849,N_14187);
xor U17421 (N_17421,N_12123,N_13312);
nor U17422 (N_17422,N_13771,N_13396);
and U17423 (N_17423,N_11788,N_11562);
and U17424 (N_17424,N_12781,N_11969);
nand U17425 (N_17425,N_11596,N_12102);
or U17426 (N_17426,N_14368,N_14611);
or U17427 (N_17427,N_14704,N_11123);
nand U17428 (N_17428,N_12470,N_14214);
and U17429 (N_17429,N_13549,N_12480);
nor U17430 (N_17430,N_12114,N_14388);
nor U17431 (N_17431,N_12393,N_12627);
nand U17432 (N_17432,N_11582,N_13218);
or U17433 (N_17433,N_11563,N_14397);
or U17434 (N_17434,N_14722,N_10834);
and U17435 (N_17435,N_13322,N_12466);
or U17436 (N_17436,N_10321,N_11608);
nor U17437 (N_17437,N_12918,N_10758);
or U17438 (N_17438,N_12098,N_14049);
nor U17439 (N_17439,N_10373,N_14034);
nor U17440 (N_17440,N_12506,N_10172);
and U17441 (N_17441,N_13774,N_13200);
and U17442 (N_17442,N_14381,N_14478);
or U17443 (N_17443,N_12624,N_14816);
and U17444 (N_17444,N_12992,N_13890);
nand U17445 (N_17445,N_11658,N_12670);
nor U17446 (N_17446,N_11425,N_11611);
nand U17447 (N_17447,N_10827,N_10353);
nor U17448 (N_17448,N_14221,N_11549);
nand U17449 (N_17449,N_13550,N_13633);
nand U17450 (N_17450,N_14225,N_14151);
xnor U17451 (N_17451,N_12877,N_14517);
nand U17452 (N_17452,N_13224,N_14375);
or U17453 (N_17453,N_14079,N_12671);
and U17454 (N_17454,N_12629,N_14077);
or U17455 (N_17455,N_11731,N_10727);
and U17456 (N_17456,N_14370,N_14674);
nor U17457 (N_17457,N_14546,N_10102);
or U17458 (N_17458,N_12923,N_11506);
xnor U17459 (N_17459,N_10729,N_14337);
and U17460 (N_17460,N_11198,N_14188);
and U17461 (N_17461,N_12103,N_10384);
xnor U17462 (N_17462,N_13554,N_13842);
xor U17463 (N_17463,N_11643,N_11272);
or U17464 (N_17464,N_10546,N_11906);
or U17465 (N_17465,N_14550,N_13870);
nand U17466 (N_17466,N_13421,N_13808);
and U17467 (N_17467,N_13408,N_10424);
nor U17468 (N_17468,N_11188,N_10448);
nand U17469 (N_17469,N_14799,N_12982);
and U17470 (N_17470,N_12917,N_14142);
nand U17471 (N_17471,N_13047,N_14340);
nor U17472 (N_17472,N_14965,N_10465);
xor U17473 (N_17473,N_13495,N_11715);
xor U17474 (N_17474,N_13963,N_11668);
xor U17475 (N_17475,N_14261,N_12415);
and U17476 (N_17476,N_12932,N_12562);
nor U17477 (N_17477,N_12119,N_13827);
or U17478 (N_17478,N_13979,N_11847);
and U17479 (N_17479,N_14509,N_12047);
nor U17480 (N_17480,N_14556,N_11216);
nand U17481 (N_17481,N_13087,N_11843);
nand U17482 (N_17482,N_14817,N_12211);
and U17483 (N_17483,N_10651,N_11585);
xor U17484 (N_17484,N_14940,N_11592);
xor U17485 (N_17485,N_14958,N_10132);
xnor U17486 (N_17486,N_12943,N_13244);
xnor U17487 (N_17487,N_10959,N_13500);
xor U17488 (N_17488,N_13763,N_12825);
xnor U17489 (N_17489,N_12875,N_13596);
or U17490 (N_17490,N_10609,N_12106);
nand U17491 (N_17491,N_14195,N_14981);
and U17492 (N_17492,N_14122,N_10978);
and U17493 (N_17493,N_14717,N_13343);
nand U17494 (N_17494,N_10550,N_10091);
nand U17495 (N_17495,N_10788,N_12850);
and U17496 (N_17496,N_14464,N_12432);
nand U17497 (N_17497,N_14751,N_14870);
xor U17498 (N_17498,N_11113,N_10088);
xnor U17499 (N_17499,N_10692,N_14678);
and U17500 (N_17500,N_10744,N_11336);
nor U17501 (N_17501,N_12858,N_14227);
nand U17502 (N_17502,N_10714,N_11299);
nand U17503 (N_17503,N_12121,N_14108);
xnor U17504 (N_17504,N_11008,N_10236);
and U17505 (N_17505,N_13430,N_10485);
nand U17506 (N_17506,N_13713,N_14115);
or U17507 (N_17507,N_11372,N_10525);
xor U17508 (N_17508,N_10242,N_11159);
nor U17509 (N_17509,N_12638,N_12269);
xnor U17510 (N_17510,N_10726,N_12256);
or U17511 (N_17511,N_10976,N_13606);
and U17512 (N_17512,N_14780,N_14448);
xor U17513 (N_17513,N_10115,N_13042);
xor U17514 (N_17514,N_14551,N_13123);
and U17515 (N_17515,N_12387,N_11466);
and U17516 (N_17516,N_13364,N_13124);
or U17517 (N_17517,N_10653,N_11908);
and U17518 (N_17518,N_11118,N_10064);
nand U17519 (N_17519,N_10950,N_13203);
or U17520 (N_17520,N_12754,N_14223);
or U17521 (N_17521,N_11814,N_11151);
xnor U17522 (N_17522,N_12144,N_10899);
nor U17523 (N_17523,N_12247,N_12551);
xor U17524 (N_17524,N_12100,N_11522);
and U17525 (N_17525,N_13481,N_13110);
xnor U17526 (N_17526,N_11075,N_14596);
xnor U17527 (N_17527,N_11081,N_10830);
nor U17528 (N_17528,N_12738,N_12551);
and U17529 (N_17529,N_14690,N_12788);
nor U17530 (N_17530,N_11507,N_10324);
xnor U17531 (N_17531,N_13360,N_14328);
xnor U17532 (N_17532,N_11776,N_13046);
or U17533 (N_17533,N_12413,N_14040);
xor U17534 (N_17534,N_10313,N_13347);
nand U17535 (N_17535,N_13341,N_14193);
nor U17536 (N_17536,N_11631,N_10914);
xor U17537 (N_17537,N_12069,N_11790);
or U17538 (N_17538,N_14092,N_10652);
xnor U17539 (N_17539,N_14362,N_11788);
nor U17540 (N_17540,N_13104,N_10967);
or U17541 (N_17541,N_14664,N_14109);
nor U17542 (N_17542,N_10784,N_13034);
or U17543 (N_17543,N_13374,N_11306);
nor U17544 (N_17544,N_12832,N_11760);
and U17545 (N_17545,N_11729,N_10888);
nand U17546 (N_17546,N_13329,N_11133);
nor U17547 (N_17547,N_14461,N_13449);
nor U17548 (N_17548,N_10097,N_13169);
or U17549 (N_17549,N_10538,N_10338);
or U17550 (N_17550,N_12139,N_13421);
and U17551 (N_17551,N_11940,N_12488);
or U17552 (N_17552,N_12791,N_13314);
or U17553 (N_17553,N_13806,N_10215);
or U17554 (N_17554,N_13855,N_10901);
xnor U17555 (N_17555,N_10928,N_11796);
nor U17556 (N_17556,N_11718,N_14584);
or U17557 (N_17557,N_10971,N_10751);
nor U17558 (N_17558,N_13255,N_12806);
or U17559 (N_17559,N_13871,N_10592);
xor U17560 (N_17560,N_14007,N_11217);
nand U17561 (N_17561,N_14386,N_14261);
or U17562 (N_17562,N_10860,N_12014);
or U17563 (N_17563,N_13700,N_14631);
xor U17564 (N_17564,N_10551,N_11217);
or U17565 (N_17565,N_14534,N_12962);
xor U17566 (N_17566,N_13211,N_14699);
nor U17567 (N_17567,N_10926,N_10543);
nand U17568 (N_17568,N_11656,N_11071);
and U17569 (N_17569,N_14271,N_12177);
nor U17570 (N_17570,N_10833,N_10121);
nor U17571 (N_17571,N_10553,N_11494);
nand U17572 (N_17572,N_13682,N_10431);
xnor U17573 (N_17573,N_13710,N_14607);
nand U17574 (N_17574,N_13034,N_11131);
and U17575 (N_17575,N_11707,N_13404);
nor U17576 (N_17576,N_13903,N_11149);
or U17577 (N_17577,N_11912,N_12311);
or U17578 (N_17578,N_12108,N_12484);
or U17579 (N_17579,N_13828,N_12323);
xnor U17580 (N_17580,N_10044,N_11367);
nand U17581 (N_17581,N_10300,N_14281);
nor U17582 (N_17582,N_12236,N_11877);
nand U17583 (N_17583,N_14576,N_11081);
nand U17584 (N_17584,N_14038,N_11225);
nor U17585 (N_17585,N_10911,N_11597);
nor U17586 (N_17586,N_13876,N_14829);
nand U17587 (N_17587,N_14123,N_14144);
or U17588 (N_17588,N_12506,N_13848);
and U17589 (N_17589,N_14801,N_11251);
and U17590 (N_17590,N_13821,N_11381);
nand U17591 (N_17591,N_11632,N_13132);
or U17592 (N_17592,N_13485,N_12254);
xor U17593 (N_17593,N_13072,N_13373);
and U17594 (N_17594,N_12899,N_13635);
and U17595 (N_17595,N_11349,N_13513);
or U17596 (N_17596,N_13071,N_13763);
xor U17597 (N_17597,N_10419,N_12899);
nand U17598 (N_17598,N_10084,N_10895);
or U17599 (N_17599,N_10289,N_14378);
or U17600 (N_17600,N_10431,N_10156);
nor U17601 (N_17601,N_10885,N_14659);
nand U17602 (N_17602,N_14456,N_10278);
nand U17603 (N_17603,N_12510,N_11975);
xnor U17604 (N_17604,N_14664,N_11264);
and U17605 (N_17605,N_10074,N_11928);
or U17606 (N_17606,N_13987,N_13370);
xor U17607 (N_17607,N_10439,N_10168);
xor U17608 (N_17608,N_13107,N_11161);
nand U17609 (N_17609,N_11197,N_10127);
xnor U17610 (N_17610,N_14855,N_14767);
or U17611 (N_17611,N_13455,N_13539);
or U17612 (N_17612,N_14284,N_13094);
and U17613 (N_17613,N_13703,N_14314);
xor U17614 (N_17614,N_14221,N_13319);
xnor U17615 (N_17615,N_12583,N_13994);
nor U17616 (N_17616,N_10581,N_12035);
and U17617 (N_17617,N_14873,N_14586);
and U17618 (N_17618,N_13413,N_13340);
and U17619 (N_17619,N_10794,N_13404);
nor U17620 (N_17620,N_14471,N_12486);
or U17621 (N_17621,N_12802,N_10983);
nor U17622 (N_17622,N_14164,N_13827);
and U17623 (N_17623,N_14971,N_13127);
or U17624 (N_17624,N_13002,N_11237);
and U17625 (N_17625,N_12096,N_10279);
or U17626 (N_17626,N_12343,N_11364);
nand U17627 (N_17627,N_12111,N_10890);
nor U17628 (N_17628,N_11455,N_14329);
nor U17629 (N_17629,N_10291,N_12739);
or U17630 (N_17630,N_14672,N_14997);
or U17631 (N_17631,N_13963,N_12671);
nand U17632 (N_17632,N_14235,N_13143);
xor U17633 (N_17633,N_14855,N_12949);
nand U17634 (N_17634,N_12233,N_11182);
or U17635 (N_17635,N_11397,N_13533);
xor U17636 (N_17636,N_10022,N_10406);
and U17637 (N_17637,N_11996,N_11876);
or U17638 (N_17638,N_10980,N_11515);
and U17639 (N_17639,N_11930,N_13908);
nor U17640 (N_17640,N_14934,N_13028);
xor U17641 (N_17641,N_13814,N_14348);
or U17642 (N_17642,N_10869,N_12569);
nand U17643 (N_17643,N_12792,N_14328);
and U17644 (N_17644,N_12756,N_13481);
or U17645 (N_17645,N_14240,N_11479);
xor U17646 (N_17646,N_14821,N_14094);
xor U17647 (N_17647,N_12738,N_11929);
xor U17648 (N_17648,N_10660,N_12123);
or U17649 (N_17649,N_14712,N_13123);
xor U17650 (N_17650,N_12845,N_10544);
nand U17651 (N_17651,N_13648,N_12247);
and U17652 (N_17652,N_10351,N_13227);
nor U17653 (N_17653,N_12744,N_10372);
xor U17654 (N_17654,N_12516,N_12846);
and U17655 (N_17655,N_11875,N_11244);
and U17656 (N_17656,N_11304,N_12884);
nor U17657 (N_17657,N_12976,N_12390);
xor U17658 (N_17658,N_14810,N_11973);
and U17659 (N_17659,N_13217,N_11861);
nor U17660 (N_17660,N_11957,N_11904);
or U17661 (N_17661,N_10161,N_10252);
nor U17662 (N_17662,N_13245,N_12559);
or U17663 (N_17663,N_14456,N_10346);
nor U17664 (N_17664,N_10753,N_14364);
xor U17665 (N_17665,N_13811,N_14828);
nand U17666 (N_17666,N_13620,N_11020);
xor U17667 (N_17667,N_11237,N_12538);
xor U17668 (N_17668,N_12625,N_14377);
and U17669 (N_17669,N_10200,N_13303);
or U17670 (N_17670,N_13044,N_12128);
or U17671 (N_17671,N_11729,N_10409);
and U17672 (N_17672,N_14507,N_13518);
xor U17673 (N_17673,N_10679,N_10983);
and U17674 (N_17674,N_10837,N_14494);
nand U17675 (N_17675,N_11016,N_12257);
or U17676 (N_17676,N_12827,N_10054);
nand U17677 (N_17677,N_13476,N_14259);
nor U17678 (N_17678,N_10321,N_14502);
or U17679 (N_17679,N_14501,N_13746);
or U17680 (N_17680,N_11019,N_10128);
or U17681 (N_17681,N_14649,N_10534);
nor U17682 (N_17682,N_11615,N_11319);
nor U17683 (N_17683,N_14394,N_13754);
xor U17684 (N_17684,N_12518,N_10248);
xor U17685 (N_17685,N_12017,N_10495);
nand U17686 (N_17686,N_13157,N_13105);
or U17687 (N_17687,N_12253,N_11949);
nor U17688 (N_17688,N_12379,N_12704);
nor U17689 (N_17689,N_14300,N_12033);
or U17690 (N_17690,N_10367,N_11486);
or U17691 (N_17691,N_11881,N_12824);
nand U17692 (N_17692,N_12681,N_13276);
xnor U17693 (N_17693,N_11243,N_13372);
or U17694 (N_17694,N_10053,N_10248);
and U17695 (N_17695,N_14177,N_14517);
xnor U17696 (N_17696,N_13894,N_14355);
nand U17697 (N_17697,N_11200,N_11435);
xnor U17698 (N_17698,N_11801,N_12212);
or U17699 (N_17699,N_14525,N_11179);
xor U17700 (N_17700,N_12165,N_11087);
xnor U17701 (N_17701,N_11790,N_13671);
nor U17702 (N_17702,N_14309,N_14632);
nor U17703 (N_17703,N_14122,N_13420);
xnor U17704 (N_17704,N_10049,N_12798);
and U17705 (N_17705,N_12958,N_14056);
xnor U17706 (N_17706,N_12832,N_12797);
or U17707 (N_17707,N_12171,N_11625);
xor U17708 (N_17708,N_11208,N_10307);
nand U17709 (N_17709,N_11608,N_13639);
nand U17710 (N_17710,N_10434,N_11817);
xor U17711 (N_17711,N_12948,N_14887);
or U17712 (N_17712,N_14815,N_11402);
or U17713 (N_17713,N_12701,N_10591);
nor U17714 (N_17714,N_10806,N_14348);
and U17715 (N_17715,N_12229,N_10988);
nand U17716 (N_17716,N_11561,N_13294);
nor U17717 (N_17717,N_13207,N_12802);
and U17718 (N_17718,N_10314,N_11865);
nor U17719 (N_17719,N_12856,N_11082);
nand U17720 (N_17720,N_14305,N_11971);
and U17721 (N_17721,N_14534,N_13073);
or U17722 (N_17722,N_14662,N_12397);
xnor U17723 (N_17723,N_13217,N_14758);
nand U17724 (N_17724,N_13484,N_11002);
or U17725 (N_17725,N_11740,N_10455);
and U17726 (N_17726,N_13981,N_14583);
and U17727 (N_17727,N_13489,N_13194);
nand U17728 (N_17728,N_11533,N_14520);
or U17729 (N_17729,N_11296,N_11813);
nor U17730 (N_17730,N_13723,N_11386);
xnor U17731 (N_17731,N_11671,N_11611);
nor U17732 (N_17732,N_10475,N_14892);
nand U17733 (N_17733,N_13392,N_10271);
nand U17734 (N_17734,N_10784,N_12654);
or U17735 (N_17735,N_13368,N_12351);
and U17736 (N_17736,N_11813,N_11137);
and U17737 (N_17737,N_10995,N_10997);
nand U17738 (N_17738,N_14064,N_11103);
and U17739 (N_17739,N_13737,N_11720);
and U17740 (N_17740,N_14989,N_10559);
nand U17741 (N_17741,N_10039,N_13317);
xor U17742 (N_17742,N_11972,N_10786);
and U17743 (N_17743,N_11522,N_12512);
nand U17744 (N_17744,N_11621,N_10296);
or U17745 (N_17745,N_14650,N_13882);
nor U17746 (N_17746,N_12297,N_11768);
nor U17747 (N_17747,N_10431,N_14615);
nand U17748 (N_17748,N_14998,N_10626);
nor U17749 (N_17749,N_10863,N_12316);
nand U17750 (N_17750,N_10813,N_14601);
and U17751 (N_17751,N_13531,N_10131);
or U17752 (N_17752,N_11370,N_12954);
and U17753 (N_17753,N_14681,N_12677);
nand U17754 (N_17754,N_13811,N_13438);
and U17755 (N_17755,N_10998,N_14096);
nor U17756 (N_17756,N_13594,N_11367);
or U17757 (N_17757,N_10973,N_11628);
nand U17758 (N_17758,N_14430,N_14704);
and U17759 (N_17759,N_12089,N_14959);
xor U17760 (N_17760,N_10874,N_13546);
nand U17761 (N_17761,N_12923,N_14361);
and U17762 (N_17762,N_10175,N_12635);
xor U17763 (N_17763,N_11794,N_11712);
and U17764 (N_17764,N_10436,N_12970);
xnor U17765 (N_17765,N_14799,N_11841);
or U17766 (N_17766,N_13946,N_10361);
and U17767 (N_17767,N_12080,N_10487);
nor U17768 (N_17768,N_13071,N_14189);
or U17769 (N_17769,N_10427,N_12275);
nand U17770 (N_17770,N_13321,N_14284);
and U17771 (N_17771,N_10572,N_14474);
nand U17772 (N_17772,N_10618,N_11029);
or U17773 (N_17773,N_14069,N_12047);
xnor U17774 (N_17774,N_10255,N_10699);
nor U17775 (N_17775,N_13923,N_11629);
nand U17776 (N_17776,N_13274,N_12169);
xnor U17777 (N_17777,N_10979,N_12653);
or U17778 (N_17778,N_13175,N_12113);
or U17779 (N_17779,N_10369,N_12041);
or U17780 (N_17780,N_14508,N_12542);
xnor U17781 (N_17781,N_14403,N_12352);
xor U17782 (N_17782,N_14793,N_10559);
or U17783 (N_17783,N_13480,N_11566);
nor U17784 (N_17784,N_14346,N_11430);
nand U17785 (N_17785,N_11174,N_12469);
xor U17786 (N_17786,N_13543,N_12061);
and U17787 (N_17787,N_12179,N_11682);
nor U17788 (N_17788,N_11850,N_10171);
xnor U17789 (N_17789,N_12255,N_12937);
nor U17790 (N_17790,N_11708,N_12421);
nand U17791 (N_17791,N_10854,N_14196);
nor U17792 (N_17792,N_10027,N_11860);
or U17793 (N_17793,N_13210,N_11685);
or U17794 (N_17794,N_12473,N_14926);
xor U17795 (N_17795,N_10564,N_11383);
nand U17796 (N_17796,N_13971,N_14818);
and U17797 (N_17797,N_13822,N_11664);
or U17798 (N_17798,N_14540,N_12032);
and U17799 (N_17799,N_12986,N_12316);
and U17800 (N_17800,N_12959,N_11774);
nand U17801 (N_17801,N_10487,N_14063);
or U17802 (N_17802,N_11816,N_12940);
nand U17803 (N_17803,N_10395,N_14933);
and U17804 (N_17804,N_12262,N_13627);
and U17805 (N_17805,N_13536,N_10758);
and U17806 (N_17806,N_14588,N_13448);
and U17807 (N_17807,N_13089,N_11656);
nor U17808 (N_17808,N_11803,N_10352);
nor U17809 (N_17809,N_11576,N_14707);
and U17810 (N_17810,N_14509,N_11054);
nand U17811 (N_17811,N_10978,N_13723);
nor U17812 (N_17812,N_10292,N_11482);
nand U17813 (N_17813,N_14813,N_10295);
and U17814 (N_17814,N_14496,N_11084);
xor U17815 (N_17815,N_12236,N_13144);
xor U17816 (N_17816,N_14385,N_14889);
nand U17817 (N_17817,N_13888,N_13798);
and U17818 (N_17818,N_12865,N_10075);
xor U17819 (N_17819,N_12753,N_10113);
xor U17820 (N_17820,N_14125,N_11141);
and U17821 (N_17821,N_14168,N_10688);
and U17822 (N_17822,N_12260,N_14394);
xnor U17823 (N_17823,N_13650,N_10934);
nor U17824 (N_17824,N_13399,N_14304);
and U17825 (N_17825,N_10711,N_14594);
nand U17826 (N_17826,N_14540,N_12439);
nand U17827 (N_17827,N_11114,N_11754);
and U17828 (N_17828,N_11770,N_13268);
and U17829 (N_17829,N_11370,N_11462);
or U17830 (N_17830,N_12738,N_12258);
or U17831 (N_17831,N_12629,N_11290);
or U17832 (N_17832,N_14119,N_13410);
nand U17833 (N_17833,N_13400,N_10851);
nand U17834 (N_17834,N_11450,N_10664);
and U17835 (N_17835,N_14260,N_11576);
xnor U17836 (N_17836,N_11458,N_10141);
nor U17837 (N_17837,N_12551,N_14890);
nor U17838 (N_17838,N_10192,N_14105);
xor U17839 (N_17839,N_12398,N_14405);
or U17840 (N_17840,N_14851,N_12299);
nor U17841 (N_17841,N_12625,N_10946);
or U17842 (N_17842,N_14098,N_10847);
xor U17843 (N_17843,N_11784,N_11987);
and U17844 (N_17844,N_10546,N_10915);
nor U17845 (N_17845,N_12642,N_13075);
nor U17846 (N_17846,N_13246,N_11321);
or U17847 (N_17847,N_14769,N_11879);
or U17848 (N_17848,N_13018,N_14544);
or U17849 (N_17849,N_12140,N_13784);
or U17850 (N_17850,N_11241,N_10941);
xnor U17851 (N_17851,N_14619,N_13239);
and U17852 (N_17852,N_10831,N_12131);
or U17853 (N_17853,N_14100,N_12536);
xnor U17854 (N_17854,N_11133,N_11952);
and U17855 (N_17855,N_11227,N_14491);
nor U17856 (N_17856,N_10891,N_12754);
or U17857 (N_17857,N_13888,N_10338);
or U17858 (N_17858,N_11189,N_11689);
and U17859 (N_17859,N_11017,N_10999);
xor U17860 (N_17860,N_11948,N_13311);
nand U17861 (N_17861,N_13220,N_11130);
xor U17862 (N_17862,N_14441,N_10692);
xnor U17863 (N_17863,N_11554,N_11600);
xnor U17864 (N_17864,N_13825,N_13625);
nor U17865 (N_17865,N_14576,N_14369);
nand U17866 (N_17866,N_13427,N_13560);
xnor U17867 (N_17867,N_13165,N_12365);
nand U17868 (N_17868,N_10441,N_14753);
xor U17869 (N_17869,N_11664,N_12665);
nand U17870 (N_17870,N_10869,N_14253);
or U17871 (N_17871,N_14212,N_14021);
nor U17872 (N_17872,N_14299,N_13970);
or U17873 (N_17873,N_12690,N_12079);
and U17874 (N_17874,N_11459,N_10729);
or U17875 (N_17875,N_14526,N_14746);
xnor U17876 (N_17876,N_12818,N_14574);
or U17877 (N_17877,N_13399,N_13140);
xor U17878 (N_17878,N_13463,N_12622);
nor U17879 (N_17879,N_14098,N_13652);
nand U17880 (N_17880,N_13185,N_13871);
or U17881 (N_17881,N_10896,N_13393);
xor U17882 (N_17882,N_10739,N_12874);
xor U17883 (N_17883,N_13865,N_14863);
and U17884 (N_17884,N_12639,N_13666);
or U17885 (N_17885,N_11808,N_10673);
nand U17886 (N_17886,N_14598,N_12931);
or U17887 (N_17887,N_12109,N_14650);
nor U17888 (N_17888,N_11983,N_14728);
nor U17889 (N_17889,N_11702,N_14405);
or U17890 (N_17890,N_11087,N_14928);
nand U17891 (N_17891,N_14293,N_13633);
xor U17892 (N_17892,N_10853,N_12026);
nand U17893 (N_17893,N_11302,N_11242);
xnor U17894 (N_17894,N_14716,N_13627);
nand U17895 (N_17895,N_11514,N_13318);
xnor U17896 (N_17896,N_14961,N_11252);
nor U17897 (N_17897,N_12678,N_10746);
nor U17898 (N_17898,N_12385,N_13391);
xnor U17899 (N_17899,N_14333,N_12650);
nand U17900 (N_17900,N_10649,N_14363);
nand U17901 (N_17901,N_13424,N_14084);
xnor U17902 (N_17902,N_11315,N_12205);
nor U17903 (N_17903,N_13775,N_12276);
and U17904 (N_17904,N_13731,N_11662);
and U17905 (N_17905,N_14367,N_12165);
nor U17906 (N_17906,N_11049,N_11821);
nand U17907 (N_17907,N_10767,N_13532);
xnor U17908 (N_17908,N_12155,N_12519);
nand U17909 (N_17909,N_12732,N_12908);
nor U17910 (N_17910,N_12394,N_11896);
nor U17911 (N_17911,N_13607,N_11270);
or U17912 (N_17912,N_11067,N_12593);
and U17913 (N_17913,N_10880,N_13483);
xor U17914 (N_17914,N_12283,N_11871);
xor U17915 (N_17915,N_14573,N_10610);
and U17916 (N_17916,N_13156,N_11968);
or U17917 (N_17917,N_12718,N_10594);
and U17918 (N_17918,N_13194,N_12794);
nand U17919 (N_17919,N_13599,N_12288);
and U17920 (N_17920,N_11058,N_14999);
nor U17921 (N_17921,N_12939,N_10456);
and U17922 (N_17922,N_13604,N_11591);
xnor U17923 (N_17923,N_12083,N_12799);
nand U17924 (N_17924,N_14141,N_10489);
xnor U17925 (N_17925,N_14903,N_10107);
xor U17926 (N_17926,N_12186,N_10796);
or U17927 (N_17927,N_13890,N_11395);
nand U17928 (N_17928,N_12223,N_12404);
nand U17929 (N_17929,N_13802,N_12629);
nor U17930 (N_17930,N_11814,N_11132);
and U17931 (N_17931,N_12116,N_13748);
and U17932 (N_17932,N_13099,N_10583);
nand U17933 (N_17933,N_11138,N_13492);
nand U17934 (N_17934,N_13374,N_13340);
nand U17935 (N_17935,N_10530,N_12924);
and U17936 (N_17936,N_14903,N_14996);
xor U17937 (N_17937,N_14407,N_10021);
and U17938 (N_17938,N_13190,N_11871);
xnor U17939 (N_17939,N_14566,N_10630);
nor U17940 (N_17940,N_10441,N_10234);
xnor U17941 (N_17941,N_13929,N_14584);
and U17942 (N_17942,N_14796,N_12527);
or U17943 (N_17943,N_11094,N_13959);
or U17944 (N_17944,N_11836,N_12484);
nor U17945 (N_17945,N_12309,N_14603);
nor U17946 (N_17946,N_10789,N_13422);
nor U17947 (N_17947,N_13628,N_10808);
or U17948 (N_17948,N_13947,N_12298);
or U17949 (N_17949,N_14898,N_14731);
and U17950 (N_17950,N_14897,N_14939);
nor U17951 (N_17951,N_10891,N_12661);
and U17952 (N_17952,N_10951,N_10397);
nor U17953 (N_17953,N_13370,N_14279);
or U17954 (N_17954,N_14895,N_13543);
and U17955 (N_17955,N_11564,N_14215);
nor U17956 (N_17956,N_10313,N_10890);
or U17957 (N_17957,N_12143,N_10661);
and U17958 (N_17958,N_14162,N_12667);
nand U17959 (N_17959,N_10058,N_11912);
nor U17960 (N_17960,N_10615,N_13910);
or U17961 (N_17961,N_11911,N_12081);
nand U17962 (N_17962,N_11509,N_10651);
nor U17963 (N_17963,N_14976,N_12329);
or U17964 (N_17964,N_10204,N_12749);
nor U17965 (N_17965,N_12414,N_13491);
or U17966 (N_17966,N_12568,N_13394);
or U17967 (N_17967,N_10337,N_11160);
and U17968 (N_17968,N_10683,N_12614);
or U17969 (N_17969,N_12282,N_12634);
nand U17970 (N_17970,N_10386,N_12091);
xnor U17971 (N_17971,N_14382,N_10027);
nand U17972 (N_17972,N_11442,N_11340);
nand U17973 (N_17973,N_12474,N_11281);
xnor U17974 (N_17974,N_12640,N_14413);
nor U17975 (N_17975,N_13099,N_10451);
xnor U17976 (N_17976,N_11153,N_11597);
nand U17977 (N_17977,N_12475,N_14378);
or U17978 (N_17978,N_12431,N_11275);
nor U17979 (N_17979,N_13644,N_14843);
nand U17980 (N_17980,N_13977,N_13498);
and U17981 (N_17981,N_10646,N_14205);
or U17982 (N_17982,N_14902,N_12578);
nor U17983 (N_17983,N_12428,N_10737);
nand U17984 (N_17984,N_14284,N_14950);
nand U17985 (N_17985,N_12276,N_13263);
and U17986 (N_17986,N_10568,N_13330);
or U17987 (N_17987,N_11405,N_10590);
nor U17988 (N_17988,N_10690,N_12364);
nor U17989 (N_17989,N_13641,N_10715);
xnor U17990 (N_17990,N_11563,N_11011);
nor U17991 (N_17991,N_14139,N_13828);
or U17992 (N_17992,N_11047,N_11592);
and U17993 (N_17993,N_11376,N_10438);
xor U17994 (N_17994,N_11066,N_13144);
and U17995 (N_17995,N_14071,N_13822);
xor U17996 (N_17996,N_14411,N_14568);
and U17997 (N_17997,N_10075,N_10845);
and U17998 (N_17998,N_10098,N_11224);
and U17999 (N_17999,N_10873,N_11013);
nor U18000 (N_18000,N_12843,N_11974);
and U18001 (N_18001,N_10753,N_12886);
and U18002 (N_18002,N_11701,N_14372);
xor U18003 (N_18003,N_13273,N_14646);
nand U18004 (N_18004,N_11514,N_14787);
nand U18005 (N_18005,N_11638,N_12812);
or U18006 (N_18006,N_13075,N_12676);
and U18007 (N_18007,N_10276,N_14386);
xor U18008 (N_18008,N_11744,N_10021);
xnor U18009 (N_18009,N_10705,N_13533);
nor U18010 (N_18010,N_14963,N_12317);
and U18011 (N_18011,N_10787,N_12591);
xor U18012 (N_18012,N_13210,N_10481);
or U18013 (N_18013,N_10619,N_13990);
nand U18014 (N_18014,N_10379,N_11827);
nor U18015 (N_18015,N_10981,N_14666);
xnor U18016 (N_18016,N_14818,N_10144);
nor U18017 (N_18017,N_14138,N_11959);
and U18018 (N_18018,N_10825,N_12611);
and U18019 (N_18019,N_14364,N_10490);
xor U18020 (N_18020,N_12418,N_11806);
nand U18021 (N_18021,N_13474,N_12229);
nand U18022 (N_18022,N_10176,N_14718);
nand U18023 (N_18023,N_14482,N_14324);
nand U18024 (N_18024,N_10722,N_10489);
and U18025 (N_18025,N_13371,N_14602);
nor U18026 (N_18026,N_13884,N_13227);
nor U18027 (N_18027,N_12193,N_11756);
nand U18028 (N_18028,N_14071,N_11422);
xnor U18029 (N_18029,N_14487,N_14515);
nor U18030 (N_18030,N_11628,N_13781);
nor U18031 (N_18031,N_13908,N_11824);
xor U18032 (N_18032,N_10859,N_12989);
xor U18033 (N_18033,N_10897,N_14423);
xor U18034 (N_18034,N_11298,N_11021);
xor U18035 (N_18035,N_11523,N_11030);
nor U18036 (N_18036,N_12415,N_12380);
or U18037 (N_18037,N_14823,N_14372);
nor U18038 (N_18038,N_11681,N_14382);
and U18039 (N_18039,N_11288,N_13144);
or U18040 (N_18040,N_14613,N_14464);
or U18041 (N_18041,N_14241,N_10073);
nor U18042 (N_18042,N_12855,N_10837);
or U18043 (N_18043,N_12845,N_10407);
and U18044 (N_18044,N_14659,N_11000);
and U18045 (N_18045,N_14709,N_14078);
or U18046 (N_18046,N_12613,N_11191);
or U18047 (N_18047,N_11195,N_12582);
or U18048 (N_18048,N_11096,N_12140);
nand U18049 (N_18049,N_13935,N_10389);
nand U18050 (N_18050,N_14801,N_14866);
nand U18051 (N_18051,N_11143,N_14010);
nand U18052 (N_18052,N_12959,N_13776);
xor U18053 (N_18053,N_11657,N_11257);
or U18054 (N_18054,N_10810,N_11845);
nand U18055 (N_18055,N_13142,N_10787);
and U18056 (N_18056,N_13341,N_13910);
xor U18057 (N_18057,N_11289,N_11677);
xnor U18058 (N_18058,N_14289,N_12046);
xor U18059 (N_18059,N_12161,N_10130);
nand U18060 (N_18060,N_14622,N_10019);
nand U18061 (N_18061,N_13424,N_12076);
and U18062 (N_18062,N_10924,N_14934);
nor U18063 (N_18063,N_12070,N_13010);
nand U18064 (N_18064,N_11131,N_14555);
and U18065 (N_18065,N_11097,N_13817);
xnor U18066 (N_18066,N_10418,N_11574);
xor U18067 (N_18067,N_10759,N_12808);
xnor U18068 (N_18068,N_12772,N_13009);
nor U18069 (N_18069,N_13350,N_12009);
nor U18070 (N_18070,N_12955,N_11371);
or U18071 (N_18071,N_11149,N_12570);
nand U18072 (N_18072,N_10375,N_12817);
or U18073 (N_18073,N_14960,N_12843);
nand U18074 (N_18074,N_13051,N_11645);
or U18075 (N_18075,N_12356,N_13270);
xnor U18076 (N_18076,N_14996,N_10049);
nor U18077 (N_18077,N_14193,N_13414);
nand U18078 (N_18078,N_12432,N_11224);
and U18079 (N_18079,N_12718,N_14575);
and U18080 (N_18080,N_12424,N_13557);
and U18081 (N_18081,N_13124,N_14977);
or U18082 (N_18082,N_12482,N_13285);
and U18083 (N_18083,N_13471,N_13152);
and U18084 (N_18084,N_14178,N_12819);
nand U18085 (N_18085,N_11674,N_11188);
or U18086 (N_18086,N_10522,N_10711);
and U18087 (N_18087,N_14113,N_13890);
xnor U18088 (N_18088,N_10013,N_11337);
and U18089 (N_18089,N_13244,N_12680);
or U18090 (N_18090,N_12056,N_14603);
or U18091 (N_18091,N_13332,N_14431);
or U18092 (N_18092,N_10700,N_14868);
nor U18093 (N_18093,N_14216,N_12044);
and U18094 (N_18094,N_12193,N_10584);
nand U18095 (N_18095,N_10788,N_13565);
and U18096 (N_18096,N_13574,N_12700);
nor U18097 (N_18097,N_10446,N_11335);
nand U18098 (N_18098,N_14711,N_12976);
or U18099 (N_18099,N_11878,N_10580);
nor U18100 (N_18100,N_10145,N_14259);
nor U18101 (N_18101,N_11359,N_10956);
xnor U18102 (N_18102,N_13744,N_13371);
or U18103 (N_18103,N_11712,N_14331);
or U18104 (N_18104,N_11164,N_10999);
or U18105 (N_18105,N_11626,N_13232);
nand U18106 (N_18106,N_11192,N_10171);
xor U18107 (N_18107,N_13433,N_13355);
xor U18108 (N_18108,N_12986,N_14725);
and U18109 (N_18109,N_11341,N_11124);
and U18110 (N_18110,N_12680,N_13279);
xor U18111 (N_18111,N_13675,N_12820);
and U18112 (N_18112,N_12800,N_12733);
nor U18113 (N_18113,N_14069,N_13246);
nand U18114 (N_18114,N_12773,N_11020);
xor U18115 (N_18115,N_12185,N_11134);
and U18116 (N_18116,N_11838,N_12714);
and U18117 (N_18117,N_14906,N_11626);
xnor U18118 (N_18118,N_13584,N_10089);
and U18119 (N_18119,N_12576,N_12222);
and U18120 (N_18120,N_14851,N_11276);
nor U18121 (N_18121,N_13744,N_10719);
xor U18122 (N_18122,N_14941,N_13452);
nor U18123 (N_18123,N_10262,N_14060);
nor U18124 (N_18124,N_10213,N_13369);
and U18125 (N_18125,N_12482,N_14442);
nor U18126 (N_18126,N_12665,N_12725);
nor U18127 (N_18127,N_14225,N_14360);
or U18128 (N_18128,N_14813,N_13524);
or U18129 (N_18129,N_14936,N_10722);
xor U18130 (N_18130,N_14462,N_13462);
nand U18131 (N_18131,N_11888,N_13969);
nor U18132 (N_18132,N_10341,N_14884);
nor U18133 (N_18133,N_12483,N_13496);
and U18134 (N_18134,N_11953,N_12240);
and U18135 (N_18135,N_10224,N_11892);
or U18136 (N_18136,N_12277,N_12536);
or U18137 (N_18137,N_10718,N_13172);
or U18138 (N_18138,N_10881,N_10646);
xor U18139 (N_18139,N_12528,N_12935);
nor U18140 (N_18140,N_10555,N_12797);
nand U18141 (N_18141,N_13915,N_10116);
nand U18142 (N_18142,N_14642,N_11452);
nand U18143 (N_18143,N_13073,N_10575);
nor U18144 (N_18144,N_10482,N_10921);
nand U18145 (N_18145,N_14583,N_10623);
xor U18146 (N_18146,N_14094,N_14272);
and U18147 (N_18147,N_12741,N_12926);
nand U18148 (N_18148,N_12538,N_10120);
and U18149 (N_18149,N_10486,N_14021);
nor U18150 (N_18150,N_14511,N_10144);
or U18151 (N_18151,N_10889,N_11263);
xnor U18152 (N_18152,N_14228,N_10421);
nor U18153 (N_18153,N_14910,N_14382);
or U18154 (N_18154,N_11864,N_13999);
and U18155 (N_18155,N_12816,N_14460);
or U18156 (N_18156,N_14337,N_13900);
or U18157 (N_18157,N_11569,N_11545);
xnor U18158 (N_18158,N_10712,N_14141);
nand U18159 (N_18159,N_14548,N_10849);
or U18160 (N_18160,N_11873,N_14909);
and U18161 (N_18161,N_10646,N_12206);
xnor U18162 (N_18162,N_10018,N_13155);
or U18163 (N_18163,N_14205,N_10315);
xor U18164 (N_18164,N_12943,N_10864);
xor U18165 (N_18165,N_11134,N_14570);
or U18166 (N_18166,N_11966,N_10342);
nand U18167 (N_18167,N_10762,N_14217);
or U18168 (N_18168,N_12106,N_12716);
xnor U18169 (N_18169,N_10243,N_12528);
and U18170 (N_18170,N_11621,N_10639);
or U18171 (N_18171,N_13867,N_13785);
nand U18172 (N_18172,N_14204,N_10413);
xor U18173 (N_18173,N_12516,N_14133);
xnor U18174 (N_18174,N_11644,N_11321);
and U18175 (N_18175,N_14698,N_11936);
or U18176 (N_18176,N_10495,N_12469);
xor U18177 (N_18177,N_14884,N_12760);
xnor U18178 (N_18178,N_13155,N_10492);
and U18179 (N_18179,N_11127,N_14611);
xnor U18180 (N_18180,N_14095,N_13870);
or U18181 (N_18181,N_11127,N_12354);
xnor U18182 (N_18182,N_12320,N_13578);
and U18183 (N_18183,N_11337,N_11868);
nor U18184 (N_18184,N_10830,N_14113);
nor U18185 (N_18185,N_12205,N_12422);
nand U18186 (N_18186,N_12857,N_10739);
or U18187 (N_18187,N_14128,N_10352);
and U18188 (N_18188,N_13157,N_13441);
nor U18189 (N_18189,N_13922,N_14923);
nor U18190 (N_18190,N_12239,N_12887);
nand U18191 (N_18191,N_12058,N_13651);
nor U18192 (N_18192,N_10696,N_14200);
or U18193 (N_18193,N_11858,N_12897);
xnor U18194 (N_18194,N_12372,N_13514);
and U18195 (N_18195,N_10925,N_11161);
nor U18196 (N_18196,N_13970,N_14122);
or U18197 (N_18197,N_13256,N_14378);
and U18198 (N_18198,N_14767,N_10922);
xnor U18199 (N_18199,N_13621,N_12983);
and U18200 (N_18200,N_12805,N_10205);
nor U18201 (N_18201,N_12258,N_14730);
xnor U18202 (N_18202,N_11556,N_10395);
nor U18203 (N_18203,N_14730,N_10287);
or U18204 (N_18204,N_13997,N_12004);
and U18205 (N_18205,N_13330,N_13366);
or U18206 (N_18206,N_12472,N_13978);
nor U18207 (N_18207,N_12400,N_12591);
nor U18208 (N_18208,N_11387,N_13423);
nand U18209 (N_18209,N_11360,N_13930);
nor U18210 (N_18210,N_13686,N_13438);
nor U18211 (N_18211,N_14226,N_10445);
and U18212 (N_18212,N_10222,N_14077);
nand U18213 (N_18213,N_14695,N_10158);
xor U18214 (N_18214,N_11413,N_10151);
and U18215 (N_18215,N_14832,N_10067);
and U18216 (N_18216,N_14007,N_12850);
xor U18217 (N_18217,N_10483,N_10355);
or U18218 (N_18218,N_14583,N_11367);
xnor U18219 (N_18219,N_13540,N_14825);
and U18220 (N_18220,N_12698,N_12783);
and U18221 (N_18221,N_13367,N_13249);
xor U18222 (N_18222,N_11434,N_11382);
nor U18223 (N_18223,N_14946,N_14398);
and U18224 (N_18224,N_14987,N_14921);
nand U18225 (N_18225,N_13630,N_14686);
xnor U18226 (N_18226,N_13569,N_11397);
xnor U18227 (N_18227,N_10583,N_12157);
nor U18228 (N_18228,N_14168,N_12493);
xnor U18229 (N_18229,N_11457,N_13443);
nand U18230 (N_18230,N_13782,N_11395);
xnor U18231 (N_18231,N_12478,N_13386);
and U18232 (N_18232,N_13763,N_13218);
nor U18233 (N_18233,N_11862,N_10726);
nor U18234 (N_18234,N_13989,N_11327);
xnor U18235 (N_18235,N_13807,N_12612);
and U18236 (N_18236,N_13847,N_12311);
and U18237 (N_18237,N_13994,N_12361);
and U18238 (N_18238,N_14020,N_10374);
xnor U18239 (N_18239,N_12015,N_12641);
xnor U18240 (N_18240,N_11515,N_14865);
and U18241 (N_18241,N_14251,N_11524);
or U18242 (N_18242,N_13735,N_12389);
and U18243 (N_18243,N_10577,N_10988);
or U18244 (N_18244,N_10434,N_12590);
nand U18245 (N_18245,N_14665,N_12468);
nand U18246 (N_18246,N_14671,N_11763);
and U18247 (N_18247,N_13503,N_12177);
or U18248 (N_18248,N_12867,N_13792);
xor U18249 (N_18249,N_13516,N_11358);
and U18250 (N_18250,N_14872,N_13714);
or U18251 (N_18251,N_13597,N_12840);
nand U18252 (N_18252,N_12533,N_11469);
or U18253 (N_18253,N_10704,N_14666);
or U18254 (N_18254,N_11195,N_13493);
xor U18255 (N_18255,N_12941,N_10523);
xor U18256 (N_18256,N_10160,N_11510);
and U18257 (N_18257,N_13879,N_14959);
nand U18258 (N_18258,N_13760,N_14988);
and U18259 (N_18259,N_13197,N_13576);
nor U18260 (N_18260,N_14980,N_14658);
xnor U18261 (N_18261,N_12116,N_14613);
or U18262 (N_18262,N_14363,N_14114);
nand U18263 (N_18263,N_12134,N_10972);
nand U18264 (N_18264,N_11255,N_14996);
nor U18265 (N_18265,N_12708,N_13976);
or U18266 (N_18266,N_11394,N_13798);
xor U18267 (N_18267,N_10437,N_12490);
nor U18268 (N_18268,N_13210,N_10807);
xnor U18269 (N_18269,N_14438,N_10738);
or U18270 (N_18270,N_10062,N_11005);
or U18271 (N_18271,N_14348,N_13745);
nand U18272 (N_18272,N_12594,N_14853);
and U18273 (N_18273,N_12511,N_13153);
or U18274 (N_18274,N_12278,N_14712);
nand U18275 (N_18275,N_11043,N_10542);
nand U18276 (N_18276,N_10537,N_13228);
nand U18277 (N_18277,N_14580,N_10464);
nor U18278 (N_18278,N_14201,N_12401);
nand U18279 (N_18279,N_13634,N_13847);
and U18280 (N_18280,N_14945,N_11834);
and U18281 (N_18281,N_10438,N_11505);
xor U18282 (N_18282,N_10897,N_14171);
nand U18283 (N_18283,N_12596,N_13535);
nor U18284 (N_18284,N_14048,N_13572);
xnor U18285 (N_18285,N_12281,N_14918);
or U18286 (N_18286,N_12154,N_14368);
xnor U18287 (N_18287,N_11840,N_14552);
and U18288 (N_18288,N_13828,N_12467);
or U18289 (N_18289,N_11170,N_10384);
nand U18290 (N_18290,N_11118,N_14199);
xnor U18291 (N_18291,N_10096,N_12669);
or U18292 (N_18292,N_12478,N_13519);
nand U18293 (N_18293,N_11878,N_11284);
and U18294 (N_18294,N_13550,N_14275);
xnor U18295 (N_18295,N_14310,N_10699);
or U18296 (N_18296,N_13803,N_10393);
and U18297 (N_18297,N_13097,N_13478);
and U18298 (N_18298,N_13444,N_10149);
or U18299 (N_18299,N_12722,N_11172);
or U18300 (N_18300,N_14092,N_13923);
nor U18301 (N_18301,N_11689,N_13145);
nand U18302 (N_18302,N_11453,N_14616);
nand U18303 (N_18303,N_10900,N_14405);
nand U18304 (N_18304,N_13301,N_14646);
xnor U18305 (N_18305,N_11483,N_12343);
and U18306 (N_18306,N_13448,N_13676);
nor U18307 (N_18307,N_11486,N_12990);
nor U18308 (N_18308,N_14105,N_11964);
xnor U18309 (N_18309,N_10770,N_11765);
xnor U18310 (N_18310,N_11582,N_11193);
xor U18311 (N_18311,N_12579,N_13503);
nand U18312 (N_18312,N_12269,N_14935);
xor U18313 (N_18313,N_11407,N_13753);
xnor U18314 (N_18314,N_11052,N_13021);
or U18315 (N_18315,N_10287,N_13791);
and U18316 (N_18316,N_11451,N_13485);
nor U18317 (N_18317,N_11638,N_12850);
nor U18318 (N_18318,N_13824,N_11354);
nand U18319 (N_18319,N_12198,N_14034);
xnor U18320 (N_18320,N_12303,N_13688);
and U18321 (N_18321,N_11101,N_13458);
and U18322 (N_18322,N_12261,N_11479);
or U18323 (N_18323,N_12147,N_11106);
or U18324 (N_18324,N_13362,N_10357);
nand U18325 (N_18325,N_12029,N_14932);
or U18326 (N_18326,N_11959,N_12720);
and U18327 (N_18327,N_14692,N_11377);
and U18328 (N_18328,N_12423,N_12792);
and U18329 (N_18329,N_10713,N_10206);
nand U18330 (N_18330,N_13292,N_13421);
nand U18331 (N_18331,N_11741,N_14055);
nor U18332 (N_18332,N_13724,N_12609);
nand U18333 (N_18333,N_11785,N_14821);
nor U18334 (N_18334,N_11185,N_12680);
nor U18335 (N_18335,N_11658,N_14709);
or U18336 (N_18336,N_14921,N_10776);
and U18337 (N_18337,N_12259,N_12305);
or U18338 (N_18338,N_10415,N_12308);
nor U18339 (N_18339,N_14490,N_12426);
xor U18340 (N_18340,N_11488,N_14555);
nor U18341 (N_18341,N_10833,N_12510);
or U18342 (N_18342,N_12407,N_14542);
nand U18343 (N_18343,N_12555,N_13260);
or U18344 (N_18344,N_10731,N_10628);
nand U18345 (N_18345,N_13380,N_13294);
and U18346 (N_18346,N_11561,N_14936);
or U18347 (N_18347,N_14675,N_12602);
xor U18348 (N_18348,N_14404,N_10708);
or U18349 (N_18349,N_13112,N_12663);
and U18350 (N_18350,N_13597,N_11616);
nand U18351 (N_18351,N_14604,N_10939);
and U18352 (N_18352,N_10629,N_13426);
nor U18353 (N_18353,N_12695,N_12530);
xnor U18354 (N_18354,N_13066,N_13658);
nand U18355 (N_18355,N_11628,N_10469);
nand U18356 (N_18356,N_14142,N_11533);
nand U18357 (N_18357,N_11834,N_14434);
and U18358 (N_18358,N_13687,N_10654);
xnor U18359 (N_18359,N_11104,N_12867);
nor U18360 (N_18360,N_14559,N_11053);
xnor U18361 (N_18361,N_13539,N_10161);
nor U18362 (N_18362,N_14854,N_10227);
nor U18363 (N_18363,N_14790,N_10783);
and U18364 (N_18364,N_12408,N_14058);
xor U18365 (N_18365,N_11115,N_12491);
and U18366 (N_18366,N_10341,N_14065);
or U18367 (N_18367,N_12310,N_10901);
nor U18368 (N_18368,N_11588,N_12778);
or U18369 (N_18369,N_11085,N_12529);
and U18370 (N_18370,N_11334,N_14797);
xor U18371 (N_18371,N_11327,N_12405);
or U18372 (N_18372,N_13978,N_10749);
nor U18373 (N_18373,N_13897,N_13586);
nor U18374 (N_18374,N_11639,N_13151);
or U18375 (N_18375,N_14465,N_13709);
or U18376 (N_18376,N_12285,N_12623);
xor U18377 (N_18377,N_11387,N_11342);
xnor U18378 (N_18378,N_10384,N_11312);
nor U18379 (N_18379,N_11973,N_11301);
and U18380 (N_18380,N_10261,N_11344);
or U18381 (N_18381,N_13848,N_10815);
nor U18382 (N_18382,N_10548,N_10646);
and U18383 (N_18383,N_10444,N_10333);
nand U18384 (N_18384,N_13820,N_12886);
or U18385 (N_18385,N_13672,N_14353);
and U18386 (N_18386,N_14395,N_12116);
nand U18387 (N_18387,N_12433,N_13118);
and U18388 (N_18388,N_13416,N_10617);
and U18389 (N_18389,N_14031,N_13745);
xor U18390 (N_18390,N_13592,N_13062);
nor U18391 (N_18391,N_11856,N_12321);
nand U18392 (N_18392,N_10155,N_12914);
and U18393 (N_18393,N_14527,N_13155);
xor U18394 (N_18394,N_14912,N_13987);
and U18395 (N_18395,N_13163,N_13066);
nand U18396 (N_18396,N_12417,N_14028);
or U18397 (N_18397,N_12570,N_10963);
xor U18398 (N_18398,N_10841,N_10336);
nor U18399 (N_18399,N_12192,N_13565);
or U18400 (N_18400,N_10483,N_13333);
xor U18401 (N_18401,N_11783,N_11968);
nor U18402 (N_18402,N_12450,N_10277);
nor U18403 (N_18403,N_14092,N_10615);
xor U18404 (N_18404,N_10999,N_10679);
or U18405 (N_18405,N_12077,N_14400);
nor U18406 (N_18406,N_13233,N_14966);
nand U18407 (N_18407,N_11039,N_12428);
xor U18408 (N_18408,N_13808,N_12941);
or U18409 (N_18409,N_13206,N_12589);
and U18410 (N_18410,N_13701,N_13059);
and U18411 (N_18411,N_11924,N_12294);
xnor U18412 (N_18412,N_13237,N_10119);
or U18413 (N_18413,N_13737,N_12301);
and U18414 (N_18414,N_14543,N_12600);
and U18415 (N_18415,N_11928,N_13917);
nor U18416 (N_18416,N_11542,N_14428);
nor U18417 (N_18417,N_10567,N_11168);
or U18418 (N_18418,N_14937,N_13201);
or U18419 (N_18419,N_10186,N_10330);
or U18420 (N_18420,N_13312,N_11470);
nor U18421 (N_18421,N_11842,N_11800);
nand U18422 (N_18422,N_14455,N_14272);
and U18423 (N_18423,N_13415,N_14391);
xor U18424 (N_18424,N_12229,N_13884);
nor U18425 (N_18425,N_10949,N_13598);
nor U18426 (N_18426,N_13086,N_10148);
xor U18427 (N_18427,N_11709,N_14794);
xor U18428 (N_18428,N_13002,N_12718);
or U18429 (N_18429,N_14371,N_13297);
xor U18430 (N_18430,N_11284,N_12524);
xnor U18431 (N_18431,N_14326,N_12255);
nand U18432 (N_18432,N_10428,N_14005);
and U18433 (N_18433,N_10933,N_11335);
or U18434 (N_18434,N_13104,N_10241);
nor U18435 (N_18435,N_13245,N_14682);
xnor U18436 (N_18436,N_11931,N_12068);
or U18437 (N_18437,N_10333,N_13050);
nor U18438 (N_18438,N_12998,N_12027);
and U18439 (N_18439,N_11250,N_14735);
xor U18440 (N_18440,N_12328,N_12366);
and U18441 (N_18441,N_11591,N_10973);
and U18442 (N_18442,N_10429,N_12799);
nand U18443 (N_18443,N_13620,N_11929);
nand U18444 (N_18444,N_14850,N_13726);
xnor U18445 (N_18445,N_14347,N_11802);
and U18446 (N_18446,N_12980,N_10436);
or U18447 (N_18447,N_12224,N_10336);
nand U18448 (N_18448,N_14193,N_14833);
or U18449 (N_18449,N_14683,N_14769);
or U18450 (N_18450,N_11269,N_11360);
nor U18451 (N_18451,N_11547,N_13525);
or U18452 (N_18452,N_12475,N_10865);
and U18453 (N_18453,N_10975,N_11724);
nand U18454 (N_18454,N_14414,N_10641);
xor U18455 (N_18455,N_14171,N_11505);
nand U18456 (N_18456,N_11330,N_10271);
nor U18457 (N_18457,N_12660,N_12700);
nor U18458 (N_18458,N_10629,N_12444);
nand U18459 (N_18459,N_14320,N_12697);
and U18460 (N_18460,N_10696,N_14379);
or U18461 (N_18461,N_13662,N_12516);
or U18462 (N_18462,N_14441,N_13159);
and U18463 (N_18463,N_14150,N_11302);
nor U18464 (N_18464,N_12295,N_14946);
nor U18465 (N_18465,N_13546,N_11775);
nand U18466 (N_18466,N_13219,N_11330);
nor U18467 (N_18467,N_13056,N_14810);
and U18468 (N_18468,N_11962,N_13676);
nor U18469 (N_18469,N_12390,N_14212);
or U18470 (N_18470,N_10428,N_13773);
nand U18471 (N_18471,N_10856,N_14061);
nor U18472 (N_18472,N_10235,N_10182);
and U18473 (N_18473,N_13677,N_10300);
nand U18474 (N_18474,N_12086,N_10668);
or U18475 (N_18475,N_12007,N_13362);
xor U18476 (N_18476,N_10995,N_14359);
xor U18477 (N_18477,N_11172,N_12797);
or U18478 (N_18478,N_14428,N_11306);
or U18479 (N_18479,N_13956,N_10655);
or U18480 (N_18480,N_10185,N_11213);
nor U18481 (N_18481,N_12975,N_14837);
nor U18482 (N_18482,N_10728,N_13793);
and U18483 (N_18483,N_12617,N_11590);
xnor U18484 (N_18484,N_12833,N_13996);
nand U18485 (N_18485,N_14201,N_12164);
xor U18486 (N_18486,N_13984,N_11397);
nor U18487 (N_18487,N_11658,N_12928);
nand U18488 (N_18488,N_14429,N_10592);
nand U18489 (N_18489,N_10032,N_12751);
and U18490 (N_18490,N_12280,N_13968);
and U18491 (N_18491,N_10489,N_14331);
and U18492 (N_18492,N_12196,N_14490);
nand U18493 (N_18493,N_14456,N_14758);
or U18494 (N_18494,N_14694,N_10511);
and U18495 (N_18495,N_14639,N_14905);
nor U18496 (N_18496,N_14455,N_13539);
or U18497 (N_18497,N_10822,N_13003);
xnor U18498 (N_18498,N_11005,N_13387);
and U18499 (N_18499,N_10794,N_14567);
nor U18500 (N_18500,N_14481,N_14510);
and U18501 (N_18501,N_14947,N_10048);
or U18502 (N_18502,N_13033,N_13586);
and U18503 (N_18503,N_11996,N_13332);
and U18504 (N_18504,N_12097,N_12425);
and U18505 (N_18505,N_10840,N_11079);
xor U18506 (N_18506,N_12179,N_14951);
nor U18507 (N_18507,N_12009,N_11282);
nor U18508 (N_18508,N_11068,N_11402);
xor U18509 (N_18509,N_12007,N_10122);
and U18510 (N_18510,N_11455,N_12452);
and U18511 (N_18511,N_10019,N_10501);
nand U18512 (N_18512,N_10504,N_11285);
and U18513 (N_18513,N_14694,N_11713);
nand U18514 (N_18514,N_11041,N_10915);
nor U18515 (N_18515,N_13611,N_13736);
or U18516 (N_18516,N_14253,N_11254);
or U18517 (N_18517,N_11320,N_14521);
nand U18518 (N_18518,N_10829,N_12831);
nand U18519 (N_18519,N_14291,N_13363);
or U18520 (N_18520,N_14673,N_10568);
nor U18521 (N_18521,N_10820,N_14434);
and U18522 (N_18522,N_11440,N_11643);
or U18523 (N_18523,N_13188,N_10905);
nor U18524 (N_18524,N_13898,N_10575);
xor U18525 (N_18525,N_11320,N_14306);
nand U18526 (N_18526,N_12393,N_14419);
and U18527 (N_18527,N_12437,N_11429);
nor U18528 (N_18528,N_13961,N_14814);
nor U18529 (N_18529,N_13543,N_14307);
or U18530 (N_18530,N_13405,N_14282);
nor U18531 (N_18531,N_11643,N_13299);
xnor U18532 (N_18532,N_12044,N_14893);
nor U18533 (N_18533,N_12426,N_14866);
nor U18534 (N_18534,N_13567,N_10121);
or U18535 (N_18535,N_10109,N_11840);
and U18536 (N_18536,N_14339,N_13301);
nand U18537 (N_18537,N_12700,N_14824);
xnor U18538 (N_18538,N_14190,N_11261);
and U18539 (N_18539,N_12676,N_13663);
or U18540 (N_18540,N_12069,N_10790);
or U18541 (N_18541,N_10171,N_11996);
nand U18542 (N_18542,N_10292,N_14846);
nand U18543 (N_18543,N_12838,N_10831);
or U18544 (N_18544,N_11669,N_10766);
or U18545 (N_18545,N_10089,N_11519);
and U18546 (N_18546,N_12289,N_13350);
xnor U18547 (N_18547,N_12697,N_12098);
nand U18548 (N_18548,N_12638,N_14146);
nand U18549 (N_18549,N_12381,N_11988);
xnor U18550 (N_18550,N_13873,N_14556);
and U18551 (N_18551,N_13675,N_11128);
nand U18552 (N_18552,N_12154,N_10908);
nor U18553 (N_18553,N_14190,N_10399);
nor U18554 (N_18554,N_13368,N_12786);
nand U18555 (N_18555,N_11790,N_11107);
nand U18556 (N_18556,N_12235,N_12089);
nor U18557 (N_18557,N_11604,N_11123);
and U18558 (N_18558,N_12356,N_14976);
nor U18559 (N_18559,N_13972,N_13177);
nand U18560 (N_18560,N_14779,N_10011);
xor U18561 (N_18561,N_11643,N_14886);
or U18562 (N_18562,N_13981,N_10215);
and U18563 (N_18563,N_13713,N_12664);
or U18564 (N_18564,N_10771,N_13630);
xnor U18565 (N_18565,N_14647,N_13363);
nor U18566 (N_18566,N_14028,N_14519);
and U18567 (N_18567,N_12316,N_12324);
xnor U18568 (N_18568,N_14783,N_12154);
or U18569 (N_18569,N_11630,N_11260);
xor U18570 (N_18570,N_13903,N_11332);
nor U18571 (N_18571,N_13171,N_12082);
and U18572 (N_18572,N_14439,N_11958);
and U18573 (N_18573,N_11054,N_10690);
xor U18574 (N_18574,N_11205,N_13321);
nor U18575 (N_18575,N_11774,N_11449);
nand U18576 (N_18576,N_12709,N_12333);
and U18577 (N_18577,N_10837,N_11380);
or U18578 (N_18578,N_13157,N_14235);
nand U18579 (N_18579,N_12133,N_14751);
xor U18580 (N_18580,N_11522,N_14013);
xnor U18581 (N_18581,N_11720,N_14501);
and U18582 (N_18582,N_12250,N_14484);
and U18583 (N_18583,N_13313,N_10085);
or U18584 (N_18584,N_10027,N_13281);
or U18585 (N_18585,N_14048,N_11835);
xor U18586 (N_18586,N_14989,N_13166);
or U18587 (N_18587,N_14475,N_14138);
nor U18588 (N_18588,N_12722,N_12118);
and U18589 (N_18589,N_14842,N_11394);
and U18590 (N_18590,N_13809,N_12293);
and U18591 (N_18591,N_13715,N_14298);
or U18592 (N_18592,N_10217,N_13751);
nor U18593 (N_18593,N_11640,N_13923);
nor U18594 (N_18594,N_12686,N_11188);
nor U18595 (N_18595,N_10695,N_14445);
or U18596 (N_18596,N_11137,N_11829);
or U18597 (N_18597,N_13227,N_13713);
nor U18598 (N_18598,N_13407,N_14964);
xnor U18599 (N_18599,N_11665,N_13191);
xor U18600 (N_18600,N_13824,N_14578);
and U18601 (N_18601,N_11627,N_14882);
or U18602 (N_18602,N_11776,N_11637);
nor U18603 (N_18603,N_11136,N_12259);
nand U18604 (N_18604,N_14216,N_11188);
and U18605 (N_18605,N_12784,N_13025);
and U18606 (N_18606,N_11640,N_12593);
xor U18607 (N_18607,N_12378,N_11575);
or U18608 (N_18608,N_12992,N_14730);
and U18609 (N_18609,N_14312,N_13685);
or U18610 (N_18610,N_13869,N_13929);
xnor U18611 (N_18611,N_12565,N_13027);
and U18612 (N_18612,N_14592,N_11228);
xor U18613 (N_18613,N_13614,N_10059);
nand U18614 (N_18614,N_11486,N_11025);
nor U18615 (N_18615,N_14832,N_11639);
nor U18616 (N_18616,N_12274,N_14950);
nor U18617 (N_18617,N_12421,N_11736);
xor U18618 (N_18618,N_14050,N_11223);
nor U18619 (N_18619,N_14376,N_12003);
or U18620 (N_18620,N_11245,N_10904);
and U18621 (N_18621,N_14878,N_14165);
and U18622 (N_18622,N_12643,N_13273);
or U18623 (N_18623,N_13366,N_14203);
xnor U18624 (N_18624,N_12931,N_11661);
or U18625 (N_18625,N_11851,N_14480);
or U18626 (N_18626,N_14971,N_11878);
nor U18627 (N_18627,N_14916,N_12912);
or U18628 (N_18628,N_12495,N_10918);
or U18629 (N_18629,N_14386,N_12305);
nand U18630 (N_18630,N_13766,N_11132);
nand U18631 (N_18631,N_12207,N_11718);
and U18632 (N_18632,N_12881,N_10898);
xor U18633 (N_18633,N_11370,N_13742);
nand U18634 (N_18634,N_12493,N_14373);
xnor U18635 (N_18635,N_10192,N_13010);
nand U18636 (N_18636,N_13050,N_12047);
nand U18637 (N_18637,N_12566,N_11006);
and U18638 (N_18638,N_14896,N_12603);
nor U18639 (N_18639,N_12032,N_14734);
xor U18640 (N_18640,N_12893,N_13342);
xor U18641 (N_18641,N_10943,N_10535);
or U18642 (N_18642,N_11046,N_10753);
nand U18643 (N_18643,N_13435,N_12206);
or U18644 (N_18644,N_11181,N_14870);
or U18645 (N_18645,N_14045,N_11116);
nor U18646 (N_18646,N_11501,N_11961);
nor U18647 (N_18647,N_10339,N_10870);
nand U18648 (N_18648,N_14788,N_14993);
and U18649 (N_18649,N_13323,N_14374);
nand U18650 (N_18650,N_10708,N_10601);
nor U18651 (N_18651,N_12643,N_13005);
nor U18652 (N_18652,N_13265,N_12888);
nand U18653 (N_18653,N_12072,N_10275);
nor U18654 (N_18654,N_12225,N_14090);
nor U18655 (N_18655,N_10248,N_13884);
nand U18656 (N_18656,N_11348,N_12083);
or U18657 (N_18657,N_12897,N_14812);
nor U18658 (N_18658,N_14995,N_10627);
nand U18659 (N_18659,N_13285,N_10247);
nor U18660 (N_18660,N_13691,N_14211);
or U18661 (N_18661,N_13074,N_10391);
nor U18662 (N_18662,N_14799,N_14552);
or U18663 (N_18663,N_10238,N_13190);
xor U18664 (N_18664,N_10158,N_14076);
or U18665 (N_18665,N_12645,N_10142);
nor U18666 (N_18666,N_10692,N_11909);
nor U18667 (N_18667,N_13646,N_14975);
and U18668 (N_18668,N_10543,N_11704);
nor U18669 (N_18669,N_12888,N_10637);
nand U18670 (N_18670,N_12820,N_14479);
xnor U18671 (N_18671,N_11479,N_11515);
and U18672 (N_18672,N_14543,N_14477);
or U18673 (N_18673,N_13741,N_14410);
or U18674 (N_18674,N_14619,N_11522);
and U18675 (N_18675,N_10537,N_14215);
nand U18676 (N_18676,N_12595,N_12888);
and U18677 (N_18677,N_13195,N_12088);
and U18678 (N_18678,N_11176,N_11210);
and U18679 (N_18679,N_11095,N_14768);
or U18680 (N_18680,N_10848,N_12818);
or U18681 (N_18681,N_13743,N_14933);
nand U18682 (N_18682,N_14841,N_11204);
or U18683 (N_18683,N_10045,N_13131);
and U18684 (N_18684,N_14330,N_11482);
nor U18685 (N_18685,N_14766,N_14818);
and U18686 (N_18686,N_13055,N_12226);
nand U18687 (N_18687,N_10325,N_14809);
nand U18688 (N_18688,N_13479,N_11277);
nor U18689 (N_18689,N_13245,N_13163);
and U18690 (N_18690,N_10119,N_13618);
nand U18691 (N_18691,N_11781,N_13016);
xor U18692 (N_18692,N_12732,N_13613);
nor U18693 (N_18693,N_13288,N_10492);
xnor U18694 (N_18694,N_10207,N_13222);
nand U18695 (N_18695,N_11465,N_12424);
or U18696 (N_18696,N_14469,N_11120);
xor U18697 (N_18697,N_13336,N_10727);
nor U18698 (N_18698,N_13160,N_14635);
xor U18699 (N_18699,N_10301,N_12806);
and U18700 (N_18700,N_14004,N_10693);
xnor U18701 (N_18701,N_11223,N_12305);
xnor U18702 (N_18702,N_14417,N_11657);
nor U18703 (N_18703,N_14095,N_11852);
nor U18704 (N_18704,N_12372,N_14781);
nor U18705 (N_18705,N_11171,N_12519);
xnor U18706 (N_18706,N_11138,N_11646);
nand U18707 (N_18707,N_10806,N_10427);
nand U18708 (N_18708,N_11672,N_11522);
nand U18709 (N_18709,N_14281,N_10629);
nor U18710 (N_18710,N_10965,N_11951);
or U18711 (N_18711,N_11926,N_12291);
nand U18712 (N_18712,N_13619,N_13050);
or U18713 (N_18713,N_14856,N_14445);
nor U18714 (N_18714,N_12424,N_13379);
nor U18715 (N_18715,N_14485,N_12525);
nand U18716 (N_18716,N_10383,N_13221);
nor U18717 (N_18717,N_14288,N_14917);
nand U18718 (N_18718,N_14673,N_12740);
xnor U18719 (N_18719,N_12381,N_11996);
nand U18720 (N_18720,N_11980,N_10972);
nor U18721 (N_18721,N_11860,N_12880);
and U18722 (N_18722,N_14269,N_14317);
nand U18723 (N_18723,N_11068,N_11635);
and U18724 (N_18724,N_12090,N_14291);
nor U18725 (N_18725,N_11592,N_13753);
and U18726 (N_18726,N_14738,N_10480);
nor U18727 (N_18727,N_10350,N_14487);
and U18728 (N_18728,N_14390,N_13472);
nor U18729 (N_18729,N_10299,N_11158);
nor U18730 (N_18730,N_13146,N_11887);
nand U18731 (N_18731,N_10734,N_13810);
xnor U18732 (N_18732,N_14878,N_13280);
and U18733 (N_18733,N_11705,N_14547);
nor U18734 (N_18734,N_12190,N_13247);
xnor U18735 (N_18735,N_13569,N_14996);
xor U18736 (N_18736,N_11996,N_12529);
and U18737 (N_18737,N_11200,N_10799);
nand U18738 (N_18738,N_14884,N_10011);
or U18739 (N_18739,N_10751,N_14537);
or U18740 (N_18740,N_13741,N_11614);
nand U18741 (N_18741,N_11622,N_13461);
and U18742 (N_18742,N_11918,N_13955);
xnor U18743 (N_18743,N_10547,N_12112);
nor U18744 (N_18744,N_14768,N_11600);
and U18745 (N_18745,N_14467,N_11367);
nor U18746 (N_18746,N_14826,N_11467);
or U18747 (N_18747,N_12597,N_10807);
nor U18748 (N_18748,N_12148,N_10280);
and U18749 (N_18749,N_11568,N_13733);
and U18750 (N_18750,N_14239,N_10580);
or U18751 (N_18751,N_14130,N_14408);
or U18752 (N_18752,N_10884,N_13881);
xor U18753 (N_18753,N_12342,N_14446);
nor U18754 (N_18754,N_13115,N_11095);
or U18755 (N_18755,N_14427,N_13593);
nand U18756 (N_18756,N_12647,N_11395);
nor U18757 (N_18757,N_10373,N_13363);
nor U18758 (N_18758,N_12413,N_12985);
nand U18759 (N_18759,N_10874,N_12459);
and U18760 (N_18760,N_14914,N_10016);
xor U18761 (N_18761,N_10063,N_12623);
xnor U18762 (N_18762,N_14494,N_14196);
xnor U18763 (N_18763,N_13692,N_10687);
nand U18764 (N_18764,N_12989,N_10068);
and U18765 (N_18765,N_14576,N_11350);
nor U18766 (N_18766,N_14408,N_13045);
xor U18767 (N_18767,N_10403,N_13263);
or U18768 (N_18768,N_13886,N_13467);
or U18769 (N_18769,N_14481,N_13064);
nand U18770 (N_18770,N_11643,N_10479);
and U18771 (N_18771,N_13007,N_14472);
and U18772 (N_18772,N_10356,N_11826);
or U18773 (N_18773,N_10550,N_10631);
and U18774 (N_18774,N_10469,N_12696);
xor U18775 (N_18775,N_13757,N_12625);
or U18776 (N_18776,N_12966,N_14012);
nand U18777 (N_18777,N_12713,N_13277);
and U18778 (N_18778,N_13859,N_14483);
nand U18779 (N_18779,N_11580,N_10282);
nand U18780 (N_18780,N_13864,N_13038);
xor U18781 (N_18781,N_14822,N_11476);
and U18782 (N_18782,N_14766,N_10939);
xnor U18783 (N_18783,N_10337,N_10492);
nand U18784 (N_18784,N_11996,N_10070);
nor U18785 (N_18785,N_12190,N_14974);
xnor U18786 (N_18786,N_13101,N_14987);
or U18787 (N_18787,N_14710,N_10533);
or U18788 (N_18788,N_14125,N_11849);
nand U18789 (N_18789,N_10836,N_10773);
xor U18790 (N_18790,N_11100,N_12872);
nand U18791 (N_18791,N_11111,N_12983);
or U18792 (N_18792,N_14251,N_13078);
nand U18793 (N_18793,N_14368,N_13835);
and U18794 (N_18794,N_13638,N_14561);
and U18795 (N_18795,N_12794,N_12150);
xor U18796 (N_18796,N_12498,N_10559);
and U18797 (N_18797,N_10914,N_13811);
nor U18798 (N_18798,N_10385,N_11912);
nor U18799 (N_18799,N_11833,N_11235);
nand U18800 (N_18800,N_14217,N_13409);
and U18801 (N_18801,N_13407,N_13449);
nand U18802 (N_18802,N_10386,N_14022);
nor U18803 (N_18803,N_12173,N_12775);
and U18804 (N_18804,N_11742,N_12909);
or U18805 (N_18805,N_11729,N_10049);
xnor U18806 (N_18806,N_11355,N_10268);
xnor U18807 (N_18807,N_13488,N_13400);
xnor U18808 (N_18808,N_13515,N_14686);
nor U18809 (N_18809,N_14259,N_13680);
nand U18810 (N_18810,N_13116,N_11083);
xnor U18811 (N_18811,N_11709,N_14670);
nor U18812 (N_18812,N_13411,N_11520);
nand U18813 (N_18813,N_12130,N_10031);
or U18814 (N_18814,N_14346,N_11884);
or U18815 (N_18815,N_10338,N_10474);
xor U18816 (N_18816,N_11116,N_13257);
or U18817 (N_18817,N_13711,N_10663);
nor U18818 (N_18818,N_12801,N_14582);
and U18819 (N_18819,N_11136,N_11244);
nand U18820 (N_18820,N_14651,N_13587);
or U18821 (N_18821,N_14387,N_11905);
nand U18822 (N_18822,N_14123,N_13302);
nand U18823 (N_18823,N_12582,N_14361);
or U18824 (N_18824,N_10154,N_10239);
or U18825 (N_18825,N_10684,N_13407);
xor U18826 (N_18826,N_13413,N_10795);
or U18827 (N_18827,N_10507,N_10842);
nor U18828 (N_18828,N_11109,N_12184);
nor U18829 (N_18829,N_12944,N_14331);
nor U18830 (N_18830,N_14931,N_13141);
nand U18831 (N_18831,N_13903,N_14730);
nor U18832 (N_18832,N_10320,N_12471);
nor U18833 (N_18833,N_13584,N_12677);
nand U18834 (N_18834,N_10459,N_10947);
xor U18835 (N_18835,N_14254,N_11284);
nor U18836 (N_18836,N_11313,N_14754);
or U18837 (N_18837,N_13640,N_10115);
nand U18838 (N_18838,N_11814,N_12509);
nor U18839 (N_18839,N_10025,N_13013);
nor U18840 (N_18840,N_10148,N_11159);
xor U18841 (N_18841,N_10527,N_11121);
and U18842 (N_18842,N_11740,N_11515);
and U18843 (N_18843,N_14142,N_10619);
or U18844 (N_18844,N_13207,N_11625);
nand U18845 (N_18845,N_12982,N_12227);
or U18846 (N_18846,N_12124,N_10936);
nor U18847 (N_18847,N_13462,N_14519);
nand U18848 (N_18848,N_11191,N_10317);
nor U18849 (N_18849,N_14983,N_12773);
or U18850 (N_18850,N_14608,N_12300);
nand U18851 (N_18851,N_12804,N_11521);
or U18852 (N_18852,N_10728,N_10791);
and U18853 (N_18853,N_12913,N_14386);
nand U18854 (N_18854,N_10737,N_10139);
and U18855 (N_18855,N_12622,N_12170);
nor U18856 (N_18856,N_14092,N_11276);
nand U18857 (N_18857,N_14947,N_14145);
or U18858 (N_18858,N_10372,N_14696);
and U18859 (N_18859,N_12776,N_11373);
nor U18860 (N_18860,N_10188,N_12806);
and U18861 (N_18861,N_13189,N_10443);
nand U18862 (N_18862,N_14957,N_10156);
nor U18863 (N_18863,N_13813,N_11269);
xor U18864 (N_18864,N_12584,N_12889);
nand U18865 (N_18865,N_12590,N_13897);
or U18866 (N_18866,N_14064,N_12557);
or U18867 (N_18867,N_14203,N_11878);
nand U18868 (N_18868,N_12447,N_10867);
nand U18869 (N_18869,N_14458,N_10133);
or U18870 (N_18870,N_10652,N_13367);
nand U18871 (N_18871,N_12661,N_11111);
nor U18872 (N_18872,N_10727,N_13178);
xor U18873 (N_18873,N_11857,N_10650);
or U18874 (N_18874,N_10581,N_11710);
and U18875 (N_18875,N_12558,N_12539);
xnor U18876 (N_18876,N_14453,N_10093);
or U18877 (N_18877,N_10567,N_14882);
or U18878 (N_18878,N_13362,N_14468);
nand U18879 (N_18879,N_14019,N_10497);
or U18880 (N_18880,N_14888,N_10984);
xor U18881 (N_18881,N_12841,N_14732);
xnor U18882 (N_18882,N_10827,N_11173);
nand U18883 (N_18883,N_11282,N_14409);
nand U18884 (N_18884,N_14065,N_10758);
nor U18885 (N_18885,N_10275,N_14659);
and U18886 (N_18886,N_11176,N_13495);
xnor U18887 (N_18887,N_11432,N_14978);
and U18888 (N_18888,N_11912,N_14860);
nand U18889 (N_18889,N_12499,N_13646);
and U18890 (N_18890,N_13221,N_13124);
nor U18891 (N_18891,N_10023,N_13212);
xnor U18892 (N_18892,N_14769,N_13951);
nor U18893 (N_18893,N_10333,N_13046);
and U18894 (N_18894,N_14765,N_14481);
nor U18895 (N_18895,N_10203,N_13892);
and U18896 (N_18896,N_14912,N_10816);
and U18897 (N_18897,N_13102,N_10815);
nand U18898 (N_18898,N_13201,N_12666);
nor U18899 (N_18899,N_10650,N_13751);
nor U18900 (N_18900,N_10210,N_10856);
xor U18901 (N_18901,N_13660,N_11674);
xor U18902 (N_18902,N_13599,N_10065);
nand U18903 (N_18903,N_12432,N_11384);
nor U18904 (N_18904,N_13907,N_13306);
nand U18905 (N_18905,N_10088,N_10869);
xnor U18906 (N_18906,N_10365,N_13447);
nand U18907 (N_18907,N_14279,N_11601);
and U18908 (N_18908,N_10205,N_14677);
or U18909 (N_18909,N_14363,N_12147);
or U18910 (N_18910,N_11415,N_12061);
or U18911 (N_18911,N_10543,N_10513);
nand U18912 (N_18912,N_13424,N_11608);
or U18913 (N_18913,N_14954,N_10466);
xnor U18914 (N_18914,N_10682,N_11588);
and U18915 (N_18915,N_13897,N_13686);
and U18916 (N_18916,N_11192,N_13401);
xnor U18917 (N_18917,N_10230,N_12430);
xor U18918 (N_18918,N_13033,N_13467);
nor U18919 (N_18919,N_12438,N_13816);
xnor U18920 (N_18920,N_14491,N_10973);
nand U18921 (N_18921,N_10261,N_10123);
or U18922 (N_18922,N_13225,N_10557);
nand U18923 (N_18923,N_13668,N_12499);
nand U18924 (N_18924,N_13430,N_12271);
and U18925 (N_18925,N_10076,N_12076);
or U18926 (N_18926,N_14425,N_13639);
or U18927 (N_18927,N_14239,N_11722);
or U18928 (N_18928,N_10458,N_13061);
nand U18929 (N_18929,N_13195,N_11909);
nor U18930 (N_18930,N_10026,N_10920);
and U18931 (N_18931,N_14597,N_10365);
xnor U18932 (N_18932,N_10028,N_13986);
and U18933 (N_18933,N_14029,N_12010);
xor U18934 (N_18934,N_10935,N_11552);
or U18935 (N_18935,N_12849,N_13989);
and U18936 (N_18936,N_14018,N_13810);
xor U18937 (N_18937,N_12177,N_12156);
nand U18938 (N_18938,N_12331,N_14496);
or U18939 (N_18939,N_13872,N_10522);
nor U18940 (N_18940,N_12461,N_14978);
and U18941 (N_18941,N_14114,N_12692);
or U18942 (N_18942,N_13199,N_12413);
and U18943 (N_18943,N_12131,N_14870);
nor U18944 (N_18944,N_12324,N_10221);
nor U18945 (N_18945,N_11598,N_14336);
or U18946 (N_18946,N_13086,N_12514);
nand U18947 (N_18947,N_11537,N_11794);
xor U18948 (N_18948,N_10725,N_14017);
or U18949 (N_18949,N_14956,N_13180);
xor U18950 (N_18950,N_13056,N_14225);
nor U18951 (N_18951,N_14907,N_13768);
nand U18952 (N_18952,N_13678,N_12918);
and U18953 (N_18953,N_13883,N_11395);
or U18954 (N_18954,N_13325,N_11708);
xor U18955 (N_18955,N_13400,N_13023);
or U18956 (N_18956,N_14460,N_14314);
nand U18957 (N_18957,N_12178,N_10230);
nor U18958 (N_18958,N_10908,N_11880);
xor U18959 (N_18959,N_11198,N_12605);
and U18960 (N_18960,N_12365,N_13537);
nor U18961 (N_18961,N_11336,N_13523);
xor U18962 (N_18962,N_11827,N_12287);
nor U18963 (N_18963,N_10714,N_12659);
nand U18964 (N_18964,N_13525,N_10889);
nand U18965 (N_18965,N_14639,N_12262);
or U18966 (N_18966,N_11558,N_13654);
nor U18967 (N_18967,N_11059,N_12732);
nor U18968 (N_18968,N_13215,N_14560);
and U18969 (N_18969,N_14028,N_12136);
and U18970 (N_18970,N_13862,N_10053);
or U18971 (N_18971,N_11400,N_13365);
and U18972 (N_18972,N_10796,N_14656);
nor U18973 (N_18973,N_11295,N_11006);
nand U18974 (N_18974,N_14226,N_13023);
nor U18975 (N_18975,N_12796,N_10276);
and U18976 (N_18976,N_14905,N_13299);
nand U18977 (N_18977,N_11857,N_11410);
and U18978 (N_18978,N_13261,N_10541);
nor U18979 (N_18979,N_14515,N_13413);
and U18980 (N_18980,N_11606,N_12773);
or U18981 (N_18981,N_12135,N_13110);
xnor U18982 (N_18982,N_14707,N_11580);
nor U18983 (N_18983,N_14762,N_12781);
xor U18984 (N_18984,N_13585,N_10953);
xnor U18985 (N_18985,N_14672,N_11528);
nand U18986 (N_18986,N_11999,N_11599);
and U18987 (N_18987,N_10785,N_11551);
nor U18988 (N_18988,N_12168,N_13891);
nand U18989 (N_18989,N_14373,N_11596);
nor U18990 (N_18990,N_11824,N_14799);
nor U18991 (N_18991,N_12311,N_14593);
xor U18992 (N_18992,N_12556,N_13857);
or U18993 (N_18993,N_13244,N_12728);
and U18994 (N_18994,N_13759,N_11189);
or U18995 (N_18995,N_10363,N_13564);
xor U18996 (N_18996,N_10492,N_11898);
or U18997 (N_18997,N_11456,N_10214);
nand U18998 (N_18998,N_10785,N_14401);
or U18999 (N_18999,N_13306,N_11787);
nand U19000 (N_19000,N_10611,N_14760);
nor U19001 (N_19001,N_12054,N_10788);
nand U19002 (N_19002,N_14692,N_13971);
and U19003 (N_19003,N_11825,N_11359);
or U19004 (N_19004,N_11487,N_14524);
xnor U19005 (N_19005,N_13798,N_11786);
nor U19006 (N_19006,N_13222,N_12420);
nand U19007 (N_19007,N_13828,N_11827);
nand U19008 (N_19008,N_10742,N_10682);
or U19009 (N_19009,N_11283,N_14393);
xor U19010 (N_19010,N_13778,N_13026);
xor U19011 (N_19011,N_14480,N_14229);
or U19012 (N_19012,N_14795,N_10265);
or U19013 (N_19013,N_11212,N_11734);
or U19014 (N_19014,N_10934,N_14595);
nor U19015 (N_19015,N_10809,N_11674);
or U19016 (N_19016,N_10924,N_12604);
nand U19017 (N_19017,N_10580,N_14594);
nand U19018 (N_19018,N_10133,N_13854);
or U19019 (N_19019,N_10912,N_12269);
or U19020 (N_19020,N_13206,N_10306);
nor U19021 (N_19021,N_11137,N_13022);
nand U19022 (N_19022,N_14836,N_11057);
nand U19023 (N_19023,N_14826,N_14563);
and U19024 (N_19024,N_13094,N_10689);
and U19025 (N_19025,N_14847,N_11947);
nor U19026 (N_19026,N_10470,N_12377);
nor U19027 (N_19027,N_14272,N_12841);
and U19028 (N_19028,N_11089,N_12738);
xnor U19029 (N_19029,N_10336,N_11857);
or U19030 (N_19030,N_14878,N_14193);
nor U19031 (N_19031,N_14026,N_14630);
xor U19032 (N_19032,N_12031,N_13152);
xor U19033 (N_19033,N_10327,N_13040);
nand U19034 (N_19034,N_12385,N_10425);
xnor U19035 (N_19035,N_12979,N_14430);
and U19036 (N_19036,N_14046,N_10747);
nand U19037 (N_19037,N_13073,N_13664);
nor U19038 (N_19038,N_13546,N_12258);
xor U19039 (N_19039,N_14887,N_10179);
nor U19040 (N_19040,N_12361,N_13952);
nand U19041 (N_19041,N_10562,N_10621);
and U19042 (N_19042,N_12240,N_10841);
nor U19043 (N_19043,N_13570,N_13526);
nand U19044 (N_19044,N_11130,N_11811);
or U19045 (N_19045,N_12413,N_13668);
nand U19046 (N_19046,N_10164,N_14637);
and U19047 (N_19047,N_10213,N_12962);
or U19048 (N_19048,N_12937,N_10636);
nor U19049 (N_19049,N_11607,N_10801);
nor U19050 (N_19050,N_13065,N_12015);
and U19051 (N_19051,N_11900,N_11029);
nor U19052 (N_19052,N_13339,N_10187);
nor U19053 (N_19053,N_14382,N_14086);
xor U19054 (N_19054,N_10252,N_11018);
xor U19055 (N_19055,N_11662,N_11739);
or U19056 (N_19056,N_12325,N_14126);
nor U19057 (N_19057,N_12712,N_13810);
nor U19058 (N_19058,N_13695,N_12383);
xnor U19059 (N_19059,N_14244,N_10177);
nor U19060 (N_19060,N_14519,N_12573);
nor U19061 (N_19061,N_14378,N_10873);
nor U19062 (N_19062,N_12370,N_11148);
and U19063 (N_19063,N_11028,N_14813);
and U19064 (N_19064,N_12721,N_10869);
nand U19065 (N_19065,N_12976,N_12205);
and U19066 (N_19066,N_10868,N_13337);
nor U19067 (N_19067,N_12006,N_12320);
nand U19068 (N_19068,N_13965,N_11559);
or U19069 (N_19069,N_12413,N_14312);
xnor U19070 (N_19070,N_11998,N_13848);
or U19071 (N_19071,N_12627,N_14271);
xnor U19072 (N_19072,N_13327,N_14735);
and U19073 (N_19073,N_14482,N_10012);
nor U19074 (N_19074,N_12732,N_11039);
nand U19075 (N_19075,N_11736,N_10145);
or U19076 (N_19076,N_13311,N_14156);
xor U19077 (N_19077,N_12786,N_13704);
nor U19078 (N_19078,N_12250,N_12400);
or U19079 (N_19079,N_13135,N_14944);
nor U19080 (N_19080,N_11657,N_10347);
and U19081 (N_19081,N_12323,N_11332);
nor U19082 (N_19082,N_12978,N_14272);
or U19083 (N_19083,N_11076,N_11498);
or U19084 (N_19084,N_13140,N_13340);
nor U19085 (N_19085,N_11995,N_14026);
nand U19086 (N_19086,N_11357,N_13451);
nor U19087 (N_19087,N_14633,N_11344);
nand U19088 (N_19088,N_12252,N_13549);
and U19089 (N_19089,N_13562,N_12558);
nand U19090 (N_19090,N_14521,N_11348);
and U19091 (N_19091,N_13717,N_11752);
nor U19092 (N_19092,N_10393,N_13622);
nand U19093 (N_19093,N_12858,N_10971);
nor U19094 (N_19094,N_12546,N_14838);
nor U19095 (N_19095,N_14825,N_14173);
or U19096 (N_19096,N_10438,N_12155);
and U19097 (N_19097,N_14907,N_10447);
and U19098 (N_19098,N_11962,N_12781);
nor U19099 (N_19099,N_13834,N_13706);
nor U19100 (N_19100,N_11963,N_12151);
nand U19101 (N_19101,N_13947,N_13234);
nor U19102 (N_19102,N_12252,N_11835);
or U19103 (N_19103,N_10571,N_10520);
and U19104 (N_19104,N_13483,N_11606);
nand U19105 (N_19105,N_10226,N_11373);
or U19106 (N_19106,N_11964,N_14370);
and U19107 (N_19107,N_10230,N_11257);
nor U19108 (N_19108,N_12176,N_12074);
xor U19109 (N_19109,N_10517,N_11661);
xnor U19110 (N_19110,N_10189,N_14870);
xor U19111 (N_19111,N_11278,N_12113);
or U19112 (N_19112,N_11025,N_10907);
xnor U19113 (N_19113,N_11165,N_14329);
and U19114 (N_19114,N_13394,N_10705);
and U19115 (N_19115,N_11062,N_12529);
nor U19116 (N_19116,N_12246,N_11739);
and U19117 (N_19117,N_12664,N_13754);
nor U19118 (N_19118,N_14970,N_14996);
or U19119 (N_19119,N_14155,N_11095);
xor U19120 (N_19120,N_11679,N_12395);
and U19121 (N_19121,N_11507,N_10748);
nor U19122 (N_19122,N_11869,N_12573);
or U19123 (N_19123,N_12406,N_10425);
xor U19124 (N_19124,N_12421,N_14327);
xor U19125 (N_19125,N_13562,N_11168);
xnor U19126 (N_19126,N_13742,N_10226);
and U19127 (N_19127,N_13727,N_11431);
or U19128 (N_19128,N_12489,N_11368);
and U19129 (N_19129,N_10808,N_14763);
xnor U19130 (N_19130,N_10021,N_12545);
nand U19131 (N_19131,N_11395,N_11343);
nand U19132 (N_19132,N_10004,N_11458);
xor U19133 (N_19133,N_14217,N_10229);
xor U19134 (N_19134,N_14713,N_11551);
xnor U19135 (N_19135,N_12007,N_12457);
nand U19136 (N_19136,N_14630,N_12818);
nand U19137 (N_19137,N_14022,N_13395);
xor U19138 (N_19138,N_13975,N_13865);
xor U19139 (N_19139,N_11854,N_13827);
nor U19140 (N_19140,N_13748,N_14522);
xnor U19141 (N_19141,N_13805,N_12739);
nand U19142 (N_19142,N_14757,N_12969);
nor U19143 (N_19143,N_13731,N_14372);
or U19144 (N_19144,N_12736,N_14187);
xor U19145 (N_19145,N_14429,N_13415);
nand U19146 (N_19146,N_12373,N_12679);
or U19147 (N_19147,N_12798,N_13430);
or U19148 (N_19148,N_12412,N_11464);
or U19149 (N_19149,N_14513,N_11377);
or U19150 (N_19150,N_12763,N_14524);
xor U19151 (N_19151,N_12068,N_11567);
xnor U19152 (N_19152,N_12276,N_12622);
or U19153 (N_19153,N_10002,N_11380);
nand U19154 (N_19154,N_14041,N_12540);
xor U19155 (N_19155,N_14326,N_11301);
xnor U19156 (N_19156,N_10258,N_11876);
xor U19157 (N_19157,N_14066,N_13380);
nor U19158 (N_19158,N_11320,N_12319);
nor U19159 (N_19159,N_12712,N_10817);
nand U19160 (N_19160,N_10601,N_13306);
and U19161 (N_19161,N_12040,N_13083);
and U19162 (N_19162,N_12937,N_13075);
nor U19163 (N_19163,N_13406,N_10504);
xor U19164 (N_19164,N_13939,N_12845);
and U19165 (N_19165,N_12207,N_11587);
nand U19166 (N_19166,N_11399,N_12478);
or U19167 (N_19167,N_10862,N_12846);
and U19168 (N_19168,N_10656,N_13948);
xor U19169 (N_19169,N_13642,N_10118);
nor U19170 (N_19170,N_11826,N_13222);
and U19171 (N_19171,N_14376,N_11362);
or U19172 (N_19172,N_14373,N_14691);
or U19173 (N_19173,N_13465,N_13039);
and U19174 (N_19174,N_12520,N_13694);
nand U19175 (N_19175,N_13132,N_10691);
and U19176 (N_19176,N_12732,N_11367);
xor U19177 (N_19177,N_11577,N_14832);
or U19178 (N_19178,N_13203,N_14559);
or U19179 (N_19179,N_13628,N_12396);
nand U19180 (N_19180,N_11458,N_10573);
and U19181 (N_19181,N_13273,N_10605);
or U19182 (N_19182,N_11863,N_10175);
nor U19183 (N_19183,N_11162,N_14611);
or U19184 (N_19184,N_11096,N_11795);
and U19185 (N_19185,N_12413,N_14276);
nand U19186 (N_19186,N_11943,N_14192);
and U19187 (N_19187,N_11298,N_13218);
nand U19188 (N_19188,N_14866,N_11722);
and U19189 (N_19189,N_14940,N_12179);
nand U19190 (N_19190,N_14878,N_12289);
or U19191 (N_19191,N_11475,N_13636);
nand U19192 (N_19192,N_13426,N_10916);
or U19193 (N_19193,N_10477,N_12130);
xnor U19194 (N_19194,N_13614,N_14651);
nand U19195 (N_19195,N_14619,N_14935);
and U19196 (N_19196,N_13852,N_13331);
nor U19197 (N_19197,N_14474,N_10016);
or U19198 (N_19198,N_13264,N_10290);
nor U19199 (N_19199,N_13099,N_13859);
xnor U19200 (N_19200,N_11130,N_13517);
and U19201 (N_19201,N_10821,N_13033);
or U19202 (N_19202,N_10815,N_12347);
nor U19203 (N_19203,N_14989,N_13000);
xor U19204 (N_19204,N_11985,N_14069);
or U19205 (N_19205,N_13097,N_12855);
and U19206 (N_19206,N_12712,N_10246);
nand U19207 (N_19207,N_14906,N_11000);
and U19208 (N_19208,N_14189,N_10796);
and U19209 (N_19209,N_10228,N_11721);
nor U19210 (N_19210,N_11990,N_11932);
nand U19211 (N_19211,N_10071,N_11403);
or U19212 (N_19212,N_10880,N_12541);
or U19213 (N_19213,N_10746,N_14186);
or U19214 (N_19214,N_10535,N_11651);
nor U19215 (N_19215,N_13349,N_13646);
xnor U19216 (N_19216,N_10121,N_13952);
nor U19217 (N_19217,N_10738,N_13739);
and U19218 (N_19218,N_12716,N_10270);
and U19219 (N_19219,N_12464,N_13895);
or U19220 (N_19220,N_14785,N_14622);
nand U19221 (N_19221,N_10503,N_12400);
and U19222 (N_19222,N_11211,N_11250);
nand U19223 (N_19223,N_14025,N_14830);
and U19224 (N_19224,N_10875,N_12190);
and U19225 (N_19225,N_12215,N_12452);
and U19226 (N_19226,N_12154,N_13005);
and U19227 (N_19227,N_14576,N_13160);
nand U19228 (N_19228,N_13471,N_13696);
nand U19229 (N_19229,N_14405,N_12588);
nor U19230 (N_19230,N_11290,N_10418);
or U19231 (N_19231,N_11056,N_11506);
nand U19232 (N_19232,N_13404,N_12292);
and U19233 (N_19233,N_13050,N_10465);
nor U19234 (N_19234,N_11578,N_12133);
xor U19235 (N_19235,N_10203,N_12808);
nand U19236 (N_19236,N_10268,N_10224);
nand U19237 (N_19237,N_13342,N_13737);
and U19238 (N_19238,N_10610,N_12816);
or U19239 (N_19239,N_13182,N_10656);
nand U19240 (N_19240,N_12763,N_14360);
xor U19241 (N_19241,N_10543,N_12002);
nor U19242 (N_19242,N_12543,N_11882);
or U19243 (N_19243,N_11481,N_12427);
nor U19244 (N_19244,N_10075,N_13773);
nor U19245 (N_19245,N_11213,N_11172);
or U19246 (N_19246,N_13921,N_12660);
xnor U19247 (N_19247,N_12608,N_12762);
and U19248 (N_19248,N_14140,N_12560);
nand U19249 (N_19249,N_12979,N_12405);
nor U19250 (N_19250,N_14001,N_12559);
or U19251 (N_19251,N_12190,N_10236);
nand U19252 (N_19252,N_12602,N_10434);
and U19253 (N_19253,N_11147,N_11638);
nand U19254 (N_19254,N_14526,N_13381);
nor U19255 (N_19255,N_10822,N_14470);
nand U19256 (N_19256,N_12395,N_13044);
or U19257 (N_19257,N_14873,N_10386);
nand U19258 (N_19258,N_12441,N_11029);
nand U19259 (N_19259,N_13551,N_10676);
nor U19260 (N_19260,N_14521,N_12452);
and U19261 (N_19261,N_12045,N_13694);
or U19262 (N_19262,N_10931,N_13474);
nand U19263 (N_19263,N_12468,N_10013);
nor U19264 (N_19264,N_12607,N_13487);
or U19265 (N_19265,N_14642,N_12804);
nor U19266 (N_19266,N_10041,N_11963);
nor U19267 (N_19267,N_13594,N_13859);
xor U19268 (N_19268,N_11937,N_14957);
and U19269 (N_19269,N_14892,N_10628);
nor U19270 (N_19270,N_13226,N_11855);
and U19271 (N_19271,N_10134,N_10588);
nor U19272 (N_19272,N_10911,N_11516);
xnor U19273 (N_19273,N_10059,N_10235);
nor U19274 (N_19274,N_10329,N_10185);
and U19275 (N_19275,N_10140,N_12685);
nand U19276 (N_19276,N_13052,N_12458);
or U19277 (N_19277,N_10338,N_14094);
xor U19278 (N_19278,N_13970,N_12911);
or U19279 (N_19279,N_10100,N_14122);
nor U19280 (N_19280,N_10302,N_13709);
or U19281 (N_19281,N_12491,N_12765);
nand U19282 (N_19282,N_11770,N_13897);
and U19283 (N_19283,N_10025,N_14227);
and U19284 (N_19284,N_11282,N_13270);
nor U19285 (N_19285,N_10501,N_10717);
nand U19286 (N_19286,N_12328,N_13457);
nor U19287 (N_19287,N_13642,N_10365);
xor U19288 (N_19288,N_13370,N_11803);
nor U19289 (N_19289,N_12176,N_12209);
xnor U19290 (N_19290,N_12222,N_13450);
nand U19291 (N_19291,N_12381,N_13085);
and U19292 (N_19292,N_10627,N_13188);
xor U19293 (N_19293,N_10533,N_10718);
nand U19294 (N_19294,N_13135,N_13102);
or U19295 (N_19295,N_13138,N_14509);
and U19296 (N_19296,N_12606,N_12795);
and U19297 (N_19297,N_11798,N_13548);
or U19298 (N_19298,N_12241,N_12920);
nand U19299 (N_19299,N_11834,N_12900);
nand U19300 (N_19300,N_13535,N_11474);
xor U19301 (N_19301,N_14239,N_11174);
or U19302 (N_19302,N_11427,N_12025);
nand U19303 (N_19303,N_12577,N_11172);
xnor U19304 (N_19304,N_12335,N_10836);
nand U19305 (N_19305,N_11417,N_14049);
nor U19306 (N_19306,N_11856,N_11350);
xnor U19307 (N_19307,N_11948,N_10326);
nand U19308 (N_19308,N_12227,N_12076);
xnor U19309 (N_19309,N_11888,N_10093);
nand U19310 (N_19310,N_11116,N_14679);
or U19311 (N_19311,N_10161,N_11370);
nor U19312 (N_19312,N_10385,N_10889);
xnor U19313 (N_19313,N_13495,N_13273);
nand U19314 (N_19314,N_11998,N_10871);
or U19315 (N_19315,N_14453,N_14972);
nand U19316 (N_19316,N_10693,N_10942);
nand U19317 (N_19317,N_14765,N_11863);
xnor U19318 (N_19318,N_11895,N_10972);
nor U19319 (N_19319,N_11252,N_11267);
or U19320 (N_19320,N_14018,N_10666);
xnor U19321 (N_19321,N_11079,N_12880);
nand U19322 (N_19322,N_14386,N_13575);
or U19323 (N_19323,N_12165,N_11944);
or U19324 (N_19324,N_14265,N_14970);
nor U19325 (N_19325,N_14060,N_14590);
and U19326 (N_19326,N_11185,N_11709);
xnor U19327 (N_19327,N_12708,N_14559);
xor U19328 (N_19328,N_14258,N_11110);
nor U19329 (N_19329,N_14337,N_13844);
and U19330 (N_19330,N_14865,N_12087);
nor U19331 (N_19331,N_11528,N_11433);
or U19332 (N_19332,N_13604,N_13579);
nor U19333 (N_19333,N_13662,N_12181);
and U19334 (N_19334,N_12547,N_13710);
nor U19335 (N_19335,N_13012,N_12971);
and U19336 (N_19336,N_12143,N_10818);
nor U19337 (N_19337,N_11818,N_12144);
nand U19338 (N_19338,N_11121,N_10902);
nand U19339 (N_19339,N_14964,N_13359);
nor U19340 (N_19340,N_12579,N_12777);
xor U19341 (N_19341,N_13649,N_14420);
nor U19342 (N_19342,N_12612,N_14592);
nor U19343 (N_19343,N_11065,N_13605);
and U19344 (N_19344,N_11923,N_13377);
xor U19345 (N_19345,N_11384,N_12551);
nor U19346 (N_19346,N_13522,N_12534);
nand U19347 (N_19347,N_13319,N_11012);
nand U19348 (N_19348,N_14079,N_14927);
and U19349 (N_19349,N_12797,N_11947);
and U19350 (N_19350,N_13265,N_10654);
xnor U19351 (N_19351,N_11157,N_10559);
and U19352 (N_19352,N_11023,N_10713);
nor U19353 (N_19353,N_13113,N_13173);
xor U19354 (N_19354,N_11837,N_10709);
xor U19355 (N_19355,N_14253,N_11461);
xnor U19356 (N_19356,N_11222,N_10503);
or U19357 (N_19357,N_10701,N_13977);
nor U19358 (N_19358,N_11623,N_10620);
nand U19359 (N_19359,N_10884,N_11085);
or U19360 (N_19360,N_12443,N_10030);
and U19361 (N_19361,N_13644,N_13241);
and U19362 (N_19362,N_13843,N_12425);
or U19363 (N_19363,N_14320,N_11680);
nand U19364 (N_19364,N_12372,N_13662);
or U19365 (N_19365,N_12834,N_11266);
and U19366 (N_19366,N_10350,N_11802);
nor U19367 (N_19367,N_11585,N_11842);
nand U19368 (N_19368,N_14704,N_13031);
xor U19369 (N_19369,N_11485,N_10749);
xor U19370 (N_19370,N_14293,N_11160);
or U19371 (N_19371,N_13809,N_12097);
xnor U19372 (N_19372,N_13152,N_11306);
or U19373 (N_19373,N_10935,N_12818);
or U19374 (N_19374,N_13280,N_13001);
and U19375 (N_19375,N_11573,N_14511);
or U19376 (N_19376,N_10448,N_10141);
xor U19377 (N_19377,N_10942,N_11778);
or U19378 (N_19378,N_12297,N_10807);
and U19379 (N_19379,N_10338,N_13526);
or U19380 (N_19380,N_13942,N_13077);
or U19381 (N_19381,N_13813,N_11025);
or U19382 (N_19382,N_10436,N_12532);
nor U19383 (N_19383,N_11482,N_14846);
and U19384 (N_19384,N_11029,N_11591);
nand U19385 (N_19385,N_11200,N_12248);
nand U19386 (N_19386,N_12273,N_11969);
nand U19387 (N_19387,N_11824,N_13480);
nor U19388 (N_19388,N_12853,N_10102);
and U19389 (N_19389,N_10561,N_11849);
or U19390 (N_19390,N_14748,N_14853);
nor U19391 (N_19391,N_11136,N_11303);
nor U19392 (N_19392,N_11724,N_12858);
and U19393 (N_19393,N_13773,N_14621);
xor U19394 (N_19394,N_11805,N_10680);
nor U19395 (N_19395,N_10201,N_12566);
nor U19396 (N_19396,N_12867,N_10326);
or U19397 (N_19397,N_10790,N_10875);
and U19398 (N_19398,N_11825,N_12283);
or U19399 (N_19399,N_12928,N_11971);
nor U19400 (N_19400,N_10237,N_13742);
nand U19401 (N_19401,N_10434,N_11473);
and U19402 (N_19402,N_10919,N_14319);
nand U19403 (N_19403,N_11706,N_14197);
and U19404 (N_19404,N_13848,N_10670);
xor U19405 (N_19405,N_10321,N_13395);
and U19406 (N_19406,N_11441,N_13857);
nor U19407 (N_19407,N_13024,N_12182);
and U19408 (N_19408,N_12452,N_11868);
nor U19409 (N_19409,N_10897,N_14377);
xnor U19410 (N_19410,N_14155,N_10492);
or U19411 (N_19411,N_13642,N_10314);
or U19412 (N_19412,N_12456,N_11589);
nand U19413 (N_19413,N_12211,N_10259);
xor U19414 (N_19414,N_11584,N_11033);
nand U19415 (N_19415,N_10465,N_10229);
and U19416 (N_19416,N_12766,N_10678);
nor U19417 (N_19417,N_14659,N_10640);
or U19418 (N_19418,N_13144,N_11353);
or U19419 (N_19419,N_13600,N_11380);
nor U19420 (N_19420,N_12697,N_14218);
or U19421 (N_19421,N_10676,N_10073);
nor U19422 (N_19422,N_14851,N_12485);
xnor U19423 (N_19423,N_10159,N_13305);
and U19424 (N_19424,N_10283,N_14589);
or U19425 (N_19425,N_12253,N_13322);
or U19426 (N_19426,N_12392,N_12930);
or U19427 (N_19427,N_12046,N_13550);
or U19428 (N_19428,N_10267,N_13817);
xnor U19429 (N_19429,N_13744,N_14104);
xor U19430 (N_19430,N_13796,N_14105);
nor U19431 (N_19431,N_11754,N_11064);
or U19432 (N_19432,N_13873,N_14784);
nand U19433 (N_19433,N_14703,N_12588);
nand U19434 (N_19434,N_13433,N_10645);
nor U19435 (N_19435,N_13192,N_13428);
and U19436 (N_19436,N_10649,N_14804);
or U19437 (N_19437,N_14403,N_10115);
nand U19438 (N_19438,N_13487,N_14902);
nand U19439 (N_19439,N_14287,N_12802);
nor U19440 (N_19440,N_11279,N_11921);
nand U19441 (N_19441,N_12631,N_13628);
xnor U19442 (N_19442,N_14911,N_10125);
or U19443 (N_19443,N_12011,N_14198);
xor U19444 (N_19444,N_11356,N_14490);
nand U19445 (N_19445,N_11871,N_13825);
xor U19446 (N_19446,N_14803,N_10619);
or U19447 (N_19447,N_10907,N_14878);
or U19448 (N_19448,N_12767,N_13181);
nor U19449 (N_19449,N_11970,N_14958);
nor U19450 (N_19450,N_10754,N_11306);
and U19451 (N_19451,N_10839,N_12862);
nand U19452 (N_19452,N_12565,N_14418);
or U19453 (N_19453,N_14004,N_13871);
nand U19454 (N_19454,N_14039,N_11490);
nand U19455 (N_19455,N_13822,N_13504);
and U19456 (N_19456,N_14218,N_13450);
nand U19457 (N_19457,N_10751,N_12181);
or U19458 (N_19458,N_12567,N_10981);
xnor U19459 (N_19459,N_11521,N_12695);
nand U19460 (N_19460,N_13404,N_11126);
or U19461 (N_19461,N_11467,N_10930);
nand U19462 (N_19462,N_14334,N_11645);
nand U19463 (N_19463,N_10910,N_12348);
xnor U19464 (N_19464,N_11796,N_14931);
and U19465 (N_19465,N_14393,N_13661);
xor U19466 (N_19466,N_12817,N_14040);
or U19467 (N_19467,N_13149,N_12290);
nor U19468 (N_19468,N_14690,N_12753);
nor U19469 (N_19469,N_14538,N_14455);
and U19470 (N_19470,N_12489,N_12076);
and U19471 (N_19471,N_12150,N_11580);
nor U19472 (N_19472,N_14020,N_12913);
or U19473 (N_19473,N_14716,N_11093);
nor U19474 (N_19474,N_11707,N_11380);
and U19475 (N_19475,N_14748,N_14001);
and U19476 (N_19476,N_10497,N_11952);
or U19477 (N_19477,N_13608,N_14975);
and U19478 (N_19478,N_10863,N_11193);
nand U19479 (N_19479,N_11187,N_13279);
nand U19480 (N_19480,N_11190,N_12405);
or U19481 (N_19481,N_14571,N_13806);
nand U19482 (N_19482,N_13313,N_12051);
nor U19483 (N_19483,N_11125,N_12622);
nand U19484 (N_19484,N_12612,N_12363);
nor U19485 (N_19485,N_11873,N_13833);
xnor U19486 (N_19486,N_10559,N_14664);
nand U19487 (N_19487,N_12566,N_10606);
nand U19488 (N_19488,N_11438,N_14313);
nand U19489 (N_19489,N_11553,N_14604);
nand U19490 (N_19490,N_10232,N_11925);
or U19491 (N_19491,N_14891,N_12380);
nor U19492 (N_19492,N_10950,N_12857);
nor U19493 (N_19493,N_12600,N_14337);
nor U19494 (N_19494,N_11360,N_13573);
nor U19495 (N_19495,N_11245,N_13312);
xnor U19496 (N_19496,N_12630,N_13799);
and U19497 (N_19497,N_10198,N_14812);
nand U19498 (N_19498,N_12271,N_12895);
nand U19499 (N_19499,N_11228,N_12033);
and U19500 (N_19500,N_12850,N_14996);
and U19501 (N_19501,N_13671,N_11849);
nor U19502 (N_19502,N_14587,N_11650);
xor U19503 (N_19503,N_13660,N_13425);
or U19504 (N_19504,N_14393,N_14091);
or U19505 (N_19505,N_14281,N_14986);
nand U19506 (N_19506,N_11387,N_14914);
nor U19507 (N_19507,N_12051,N_10469);
nand U19508 (N_19508,N_14002,N_13236);
nand U19509 (N_19509,N_13213,N_12760);
or U19510 (N_19510,N_14597,N_14431);
and U19511 (N_19511,N_13467,N_14634);
or U19512 (N_19512,N_11896,N_13927);
nor U19513 (N_19513,N_12856,N_14737);
nor U19514 (N_19514,N_13348,N_11778);
xnor U19515 (N_19515,N_10468,N_10173);
and U19516 (N_19516,N_14799,N_10603);
or U19517 (N_19517,N_14204,N_13353);
and U19518 (N_19518,N_10003,N_14596);
and U19519 (N_19519,N_13546,N_11734);
nor U19520 (N_19520,N_14614,N_10829);
nand U19521 (N_19521,N_14087,N_12692);
nor U19522 (N_19522,N_12504,N_12795);
nor U19523 (N_19523,N_10071,N_14428);
nand U19524 (N_19524,N_12573,N_11646);
and U19525 (N_19525,N_14453,N_13630);
or U19526 (N_19526,N_10158,N_11254);
nand U19527 (N_19527,N_11720,N_14365);
or U19528 (N_19528,N_14985,N_14291);
or U19529 (N_19529,N_12725,N_11398);
nor U19530 (N_19530,N_12020,N_10524);
or U19531 (N_19531,N_12130,N_12381);
nand U19532 (N_19532,N_10128,N_11260);
nand U19533 (N_19533,N_11989,N_14741);
nor U19534 (N_19534,N_10589,N_11325);
nor U19535 (N_19535,N_10891,N_11379);
and U19536 (N_19536,N_13074,N_13562);
nor U19537 (N_19537,N_10729,N_14950);
nor U19538 (N_19538,N_14817,N_12368);
xor U19539 (N_19539,N_14944,N_11151);
or U19540 (N_19540,N_10981,N_12765);
or U19541 (N_19541,N_13767,N_12945);
nor U19542 (N_19542,N_13707,N_12463);
nand U19543 (N_19543,N_13985,N_14114);
or U19544 (N_19544,N_11490,N_11867);
nor U19545 (N_19545,N_14157,N_11091);
and U19546 (N_19546,N_10947,N_13663);
nand U19547 (N_19547,N_13307,N_13181);
nand U19548 (N_19548,N_14753,N_10683);
and U19549 (N_19549,N_13207,N_14132);
xnor U19550 (N_19550,N_14090,N_12560);
and U19551 (N_19551,N_10505,N_14234);
nand U19552 (N_19552,N_11777,N_12960);
or U19553 (N_19553,N_10469,N_13157);
xnor U19554 (N_19554,N_12143,N_10150);
nor U19555 (N_19555,N_10042,N_11849);
and U19556 (N_19556,N_14567,N_13892);
nor U19557 (N_19557,N_12704,N_11858);
or U19558 (N_19558,N_11781,N_14498);
nor U19559 (N_19559,N_14324,N_12024);
or U19560 (N_19560,N_11874,N_10262);
xor U19561 (N_19561,N_13595,N_10846);
xnor U19562 (N_19562,N_13356,N_11334);
nand U19563 (N_19563,N_11521,N_14990);
or U19564 (N_19564,N_11852,N_11109);
and U19565 (N_19565,N_11926,N_10747);
and U19566 (N_19566,N_14293,N_10750);
xor U19567 (N_19567,N_10295,N_13224);
or U19568 (N_19568,N_11361,N_10464);
and U19569 (N_19569,N_10519,N_13319);
xnor U19570 (N_19570,N_12976,N_11419);
nor U19571 (N_19571,N_14934,N_11040);
xnor U19572 (N_19572,N_10710,N_10614);
nand U19573 (N_19573,N_11322,N_11136);
nor U19574 (N_19574,N_14254,N_14359);
nand U19575 (N_19575,N_10113,N_10527);
or U19576 (N_19576,N_11813,N_13877);
nand U19577 (N_19577,N_12804,N_12303);
xnor U19578 (N_19578,N_10752,N_11488);
nand U19579 (N_19579,N_10313,N_11881);
or U19580 (N_19580,N_12682,N_10674);
nor U19581 (N_19581,N_11445,N_11433);
or U19582 (N_19582,N_13571,N_14985);
or U19583 (N_19583,N_13327,N_13258);
xor U19584 (N_19584,N_11655,N_14399);
and U19585 (N_19585,N_14264,N_13334);
and U19586 (N_19586,N_12162,N_12589);
xor U19587 (N_19587,N_13957,N_12563);
nand U19588 (N_19588,N_13315,N_14833);
or U19589 (N_19589,N_10001,N_11606);
and U19590 (N_19590,N_13815,N_10696);
and U19591 (N_19591,N_13213,N_11301);
nor U19592 (N_19592,N_12305,N_13740);
nor U19593 (N_19593,N_13133,N_10852);
or U19594 (N_19594,N_13611,N_10942);
xor U19595 (N_19595,N_14719,N_12826);
nand U19596 (N_19596,N_10435,N_13562);
xor U19597 (N_19597,N_13741,N_13699);
nand U19598 (N_19598,N_10000,N_10504);
nand U19599 (N_19599,N_11532,N_14903);
xnor U19600 (N_19600,N_14488,N_10517);
nand U19601 (N_19601,N_11597,N_14562);
or U19602 (N_19602,N_13854,N_14394);
xnor U19603 (N_19603,N_12455,N_14308);
nand U19604 (N_19604,N_14010,N_10015);
nor U19605 (N_19605,N_14125,N_13583);
nor U19606 (N_19606,N_14512,N_14523);
and U19607 (N_19607,N_14007,N_14182);
nand U19608 (N_19608,N_14876,N_11332);
and U19609 (N_19609,N_14103,N_13987);
or U19610 (N_19610,N_13314,N_10494);
or U19611 (N_19611,N_10986,N_10405);
nand U19612 (N_19612,N_10027,N_13770);
nor U19613 (N_19613,N_13248,N_13126);
nand U19614 (N_19614,N_12760,N_12783);
nand U19615 (N_19615,N_14339,N_11873);
and U19616 (N_19616,N_11719,N_12137);
and U19617 (N_19617,N_14062,N_10741);
or U19618 (N_19618,N_14708,N_10344);
or U19619 (N_19619,N_11871,N_11406);
nor U19620 (N_19620,N_10273,N_11522);
xor U19621 (N_19621,N_11535,N_13486);
xor U19622 (N_19622,N_12160,N_14760);
nand U19623 (N_19623,N_12547,N_10651);
nand U19624 (N_19624,N_14263,N_11966);
xor U19625 (N_19625,N_10934,N_12699);
nand U19626 (N_19626,N_14851,N_11271);
or U19627 (N_19627,N_11502,N_11692);
xnor U19628 (N_19628,N_13957,N_10737);
nand U19629 (N_19629,N_12036,N_14770);
nor U19630 (N_19630,N_13222,N_12214);
nor U19631 (N_19631,N_14082,N_13637);
or U19632 (N_19632,N_12073,N_14068);
and U19633 (N_19633,N_13532,N_14734);
nand U19634 (N_19634,N_13050,N_11528);
xnor U19635 (N_19635,N_12729,N_12442);
and U19636 (N_19636,N_11373,N_14773);
nor U19637 (N_19637,N_13295,N_13643);
nor U19638 (N_19638,N_13600,N_14377);
xnor U19639 (N_19639,N_12357,N_10677);
nor U19640 (N_19640,N_11436,N_11513);
xnor U19641 (N_19641,N_13972,N_12318);
nor U19642 (N_19642,N_12732,N_14414);
nor U19643 (N_19643,N_11691,N_11501);
or U19644 (N_19644,N_12816,N_14636);
and U19645 (N_19645,N_14519,N_12041);
nand U19646 (N_19646,N_14072,N_12907);
nor U19647 (N_19647,N_12597,N_13039);
nor U19648 (N_19648,N_13991,N_10990);
nand U19649 (N_19649,N_10930,N_14544);
nand U19650 (N_19650,N_13537,N_14438);
nand U19651 (N_19651,N_11206,N_12697);
xnor U19652 (N_19652,N_13687,N_11687);
nand U19653 (N_19653,N_10573,N_13383);
and U19654 (N_19654,N_12034,N_10567);
and U19655 (N_19655,N_11276,N_12116);
xor U19656 (N_19656,N_12181,N_10150);
or U19657 (N_19657,N_14865,N_12074);
nor U19658 (N_19658,N_14727,N_11070);
or U19659 (N_19659,N_12920,N_12949);
nor U19660 (N_19660,N_10030,N_14852);
and U19661 (N_19661,N_12781,N_11265);
nand U19662 (N_19662,N_13337,N_10529);
nor U19663 (N_19663,N_14492,N_11362);
and U19664 (N_19664,N_13675,N_11465);
nand U19665 (N_19665,N_12443,N_10034);
and U19666 (N_19666,N_10878,N_14585);
or U19667 (N_19667,N_13233,N_10462);
and U19668 (N_19668,N_14026,N_10944);
and U19669 (N_19669,N_14168,N_12997);
nand U19670 (N_19670,N_13777,N_11332);
nor U19671 (N_19671,N_14256,N_12789);
nor U19672 (N_19672,N_13037,N_12635);
or U19673 (N_19673,N_12158,N_14475);
xnor U19674 (N_19674,N_11445,N_11893);
nand U19675 (N_19675,N_14892,N_13251);
and U19676 (N_19676,N_14645,N_11026);
or U19677 (N_19677,N_12819,N_13755);
nor U19678 (N_19678,N_13965,N_10747);
xor U19679 (N_19679,N_14972,N_11831);
and U19680 (N_19680,N_14192,N_11818);
xnor U19681 (N_19681,N_12278,N_11242);
nor U19682 (N_19682,N_11579,N_14670);
nor U19683 (N_19683,N_10777,N_13029);
or U19684 (N_19684,N_13288,N_13885);
xor U19685 (N_19685,N_10548,N_13652);
nand U19686 (N_19686,N_14311,N_10213);
nand U19687 (N_19687,N_13075,N_11105);
xor U19688 (N_19688,N_13277,N_11092);
and U19689 (N_19689,N_10042,N_14366);
nor U19690 (N_19690,N_13131,N_13182);
xor U19691 (N_19691,N_14675,N_10062);
xnor U19692 (N_19692,N_10207,N_13252);
and U19693 (N_19693,N_10002,N_12358);
xnor U19694 (N_19694,N_13213,N_10065);
nand U19695 (N_19695,N_13739,N_12331);
nor U19696 (N_19696,N_14676,N_13500);
xnor U19697 (N_19697,N_10179,N_12896);
and U19698 (N_19698,N_11949,N_10651);
xnor U19699 (N_19699,N_11607,N_11316);
nand U19700 (N_19700,N_12383,N_13289);
nor U19701 (N_19701,N_11704,N_13219);
nor U19702 (N_19702,N_13565,N_10150);
xnor U19703 (N_19703,N_12253,N_10963);
nor U19704 (N_19704,N_14814,N_11960);
xnor U19705 (N_19705,N_14430,N_14707);
nor U19706 (N_19706,N_10985,N_12764);
xnor U19707 (N_19707,N_14331,N_10116);
and U19708 (N_19708,N_13220,N_13563);
nand U19709 (N_19709,N_10878,N_11906);
nor U19710 (N_19710,N_11841,N_10092);
and U19711 (N_19711,N_10160,N_14281);
or U19712 (N_19712,N_11325,N_10398);
or U19713 (N_19713,N_12664,N_10125);
xor U19714 (N_19714,N_12720,N_11159);
xor U19715 (N_19715,N_13693,N_14656);
nor U19716 (N_19716,N_13166,N_12520);
and U19717 (N_19717,N_10148,N_11808);
nand U19718 (N_19718,N_14298,N_14856);
xor U19719 (N_19719,N_14529,N_12010);
nand U19720 (N_19720,N_10191,N_11364);
nand U19721 (N_19721,N_14316,N_12744);
and U19722 (N_19722,N_10603,N_13019);
and U19723 (N_19723,N_14240,N_12470);
nand U19724 (N_19724,N_10925,N_14346);
nand U19725 (N_19725,N_12612,N_11429);
or U19726 (N_19726,N_12453,N_10919);
xnor U19727 (N_19727,N_13399,N_14057);
and U19728 (N_19728,N_14287,N_11309);
nor U19729 (N_19729,N_10049,N_11857);
nor U19730 (N_19730,N_12011,N_11763);
xnor U19731 (N_19731,N_14575,N_13873);
xor U19732 (N_19732,N_10150,N_12659);
xor U19733 (N_19733,N_12392,N_12318);
or U19734 (N_19734,N_13884,N_10954);
nand U19735 (N_19735,N_13973,N_11396);
nand U19736 (N_19736,N_10825,N_12656);
nor U19737 (N_19737,N_10979,N_11212);
nor U19738 (N_19738,N_12664,N_14145);
xor U19739 (N_19739,N_14257,N_10893);
or U19740 (N_19740,N_13834,N_13356);
nand U19741 (N_19741,N_14815,N_10024);
and U19742 (N_19742,N_14075,N_14339);
or U19743 (N_19743,N_12516,N_13025);
xnor U19744 (N_19744,N_14317,N_12032);
or U19745 (N_19745,N_12579,N_11539);
xor U19746 (N_19746,N_12373,N_11875);
nor U19747 (N_19747,N_11760,N_10804);
and U19748 (N_19748,N_14374,N_12280);
xnor U19749 (N_19749,N_11215,N_12326);
nand U19750 (N_19750,N_10794,N_12881);
and U19751 (N_19751,N_10298,N_12687);
nor U19752 (N_19752,N_11247,N_12835);
nand U19753 (N_19753,N_12523,N_14872);
and U19754 (N_19754,N_14510,N_12476);
or U19755 (N_19755,N_10448,N_10544);
or U19756 (N_19756,N_14336,N_13078);
nand U19757 (N_19757,N_12547,N_14269);
and U19758 (N_19758,N_11651,N_10876);
nand U19759 (N_19759,N_11573,N_10416);
or U19760 (N_19760,N_13319,N_11268);
and U19761 (N_19761,N_11603,N_14833);
nor U19762 (N_19762,N_14261,N_11361);
and U19763 (N_19763,N_14153,N_14934);
and U19764 (N_19764,N_14602,N_13454);
or U19765 (N_19765,N_10154,N_11026);
nand U19766 (N_19766,N_14795,N_14175);
xor U19767 (N_19767,N_13452,N_10795);
xor U19768 (N_19768,N_14822,N_11471);
nor U19769 (N_19769,N_13276,N_13014);
nand U19770 (N_19770,N_12739,N_11072);
nand U19771 (N_19771,N_13729,N_12793);
nor U19772 (N_19772,N_12323,N_12071);
nor U19773 (N_19773,N_12023,N_13252);
nand U19774 (N_19774,N_10560,N_13775);
or U19775 (N_19775,N_14588,N_12490);
nand U19776 (N_19776,N_14673,N_11381);
xnor U19777 (N_19777,N_11314,N_13791);
nor U19778 (N_19778,N_12476,N_12183);
nand U19779 (N_19779,N_12580,N_10862);
nand U19780 (N_19780,N_11741,N_14413);
nand U19781 (N_19781,N_10414,N_12060);
nor U19782 (N_19782,N_14614,N_10169);
xor U19783 (N_19783,N_11365,N_11677);
or U19784 (N_19784,N_12112,N_14113);
nor U19785 (N_19785,N_11139,N_14946);
or U19786 (N_19786,N_11793,N_14778);
and U19787 (N_19787,N_10861,N_11846);
nor U19788 (N_19788,N_14642,N_10190);
and U19789 (N_19789,N_11033,N_14689);
and U19790 (N_19790,N_10333,N_13486);
xor U19791 (N_19791,N_12671,N_10032);
xnor U19792 (N_19792,N_11681,N_12867);
and U19793 (N_19793,N_13832,N_11078);
xnor U19794 (N_19794,N_14787,N_13061);
and U19795 (N_19795,N_14194,N_11539);
xor U19796 (N_19796,N_14683,N_12533);
nand U19797 (N_19797,N_11091,N_12014);
or U19798 (N_19798,N_11889,N_11626);
xor U19799 (N_19799,N_13596,N_10012);
or U19800 (N_19800,N_10583,N_14958);
nand U19801 (N_19801,N_10650,N_11916);
nor U19802 (N_19802,N_11952,N_14043);
or U19803 (N_19803,N_13238,N_14502);
and U19804 (N_19804,N_12888,N_12437);
nor U19805 (N_19805,N_14877,N_14487);
nor U19806 (N_19806,N_13694,N_13731);
or U19807 (N_19807,N_10075,N_11653);
xor U19808 (N_19808,N_10876,N_10260);
nand U19809 (N_19809,N_11942,N_12591);
nand U19810 (N_19810,N_14031,N_14231);
and U19811 (N_19811,N_14920,N_14760);
nor U19812 (N_19812,N_11319,N_13627);
nor U19813 (N_19813,N_13846,N_11869);
or U19814 (N_19814,N_10043,N_14051);
xor U19815 (N_19815,N_12403,N_12114);
xor U19816 (N_19816,N_13354,N_12684);
nor U19817 (N_19817,N_10289,N_13596);
nor U19818 (N_19818,N_14305,N_13600);
and U19819 (N_19819,N_13525,N_14713);
and U19820 (N_19820,N_11033,N_12811);
nand U19821 (N_19821,N_13226,N_11096);
xor U19822 (N_19822,N_13686,N_13217);
nand U19823 (N_19823,N_12269,N_14229);
or U19824 (N_19824,N_13684,N_11153);
nand U19825 (N_19825,N_13559,N_10190);
or U19826 (N_19826,N_10177,N_11289);
nand U19827 (N_19827,N_11014,N_10154);
xnor U19828 (N_19828,N_13853,N_11081);
nand U19829 (N_19829,N_14722,N_12478);
nor U19830 (N_19830,N_12228,N_13285);
or U19831 (N_19831,N_10754,N_14169);
and U19832 (N_19832,N_10647,N_10086);
or U19833 (N_19833,N_11472,N_13907);
xor U19834 (N_19834,N_11497,N_13007);
nor U19835 (N_19835,N_14936,N_12194);
xor U19836 (N_19836,N_11837,N_12065);
and U19837 (N_19837,N_11258,N_11659);
nand U19838 (N_19838,N_11535,N_14100);
nand U19839 (N_19839,N_13071,N_13534);
xor U19840 (N_19840,N_11372,N_11938);
nor U19841 (N_19841,N_10259,N_14335);
nand U19842 (N_19842,N_14943,N_14231);
and U19843 (N_19843,N_12548,N_10815);
xnor U19844 (N_19844,N_13476,N_11762);
nand U19845 (N_19845,N_11820,N_14769);
nand U19846 (N_19846,N_12675,N_14887);
xor U19847 (N_19847,N_10800,N_13487);
nor U19848 (N_19848,N_12408,N_12636);
or U19849 (N_19849,N_14393,N_11535);
nand U19850 (N_19850,N_14084,N_14520);
nand U19851 (N_19851,N_10131,N_13489);
or U19852 (N_19852,N_11075,N_10910);
or U19853 (N_19853,N_11775,N_12879);
nor U19854 (N_19854,N_11194,N_13488);
xnor U19855 (N_19855,N_14970,N_14342);
xor U19856 (N_19856,N_13900,N_14838);
nand U19857 (N_19857,N_13307,N_11585);
or U19858 (N_19858,N_14372,N_11258);
or U19859 (N_19859,N_14423,N_10253);
xor U19860 (N_19860,N_12373,N_10386);
or U19861 (N_19861,N_10238,N_12113);
nand U19862 (N_19862,N_14121,N_11217);
nand U19863 (N_19863,N_11220,N_11300);
xnor U19864 (N_19864,N_11978,N_13920);
xnor U19865 (N_19865,N_10104,N_10557);
nand U19866 (N_19866,N_14259,N_12999);
xor U19867 (N_19867,N_12721,N_12638);
xor U19868 (N_19868,N_10691,N_11335);
or U19869 (N_19869,N_12178,N_12490);
and U19870 (N_19870,N_14212,N_11812);
and U19871 (N_19871,N_11426,N_11150);
or U19872 (N_19872,N_13358,N_10770);
xor U19873 (N_19873,N_12960,N_10555);
nand U19874 (N_19874,N_14409,N_10638);
nand U19875 (N_19875,N_11232,N_13002);
and U19876 (N_19876,N_12333,N_14553);
nor U19877 (N_19877,N_13910,N_13232);
nor U19878 (N_19878,N_13394,N_12658);
or U19879 (N_19879,N_11811,N_11892);
xnor U19880 (N_19880,N_11717,N_14663);
nor U19881 (N_19881,N_13019,N_12812);
or U19882 (N_19882,N_14092,N_14961);
and U19883 (N_19883,N_12902,N_13172);
or U19884 (N_19884,N_11052,N_11304);
nand U19885 (N_19885,N_11980,N_10254);
nand U19886 (N_19886,N_13292,N_12811);
nor U19887 (N_19887,N_14768,N_14770);
nor U19888 (N_19888,N_13752,N_13017);
xnor U19889 (N_19889,N_12184,N_14992);
or U19890 (N_19890,N_13398,N_14497);
or U19891 (N_19891,N_14939,N_11269);
xor U19892 (N_19892,N_10069,N_12105);
and U19893 (N_19893,N_10431,N_11178);
nor U19894 (N_19894,N_13375,N_12186);
or U19895 (N_19895,N_14866,N_13885);
xnor U19896 (N_19896,N_10548,N_10359);
xnor U19897 (N_19897,N_12810,N_11359);
nand U19898 (N_19898,N_11349,N_13196);
and U19899 (N_19899,N_11671,N_13187);
and U19900 (N_19900,N_12806,N_12492);
nand U19901 (N_19901,N_12158,N_11598);
xor U19902 (N_19902,N_12877,N_12543);
nand U19903 (N_19903,N_11868,N_12531);
xor U19904 (N_19904,N_14878,N_11129);
nand U19905 (N_19905,N_10538,N_11269);
xnor U19906 (N_19906,N_13334,N_14576);
or U19907 (N_19907,N_13849,N_10294);
xnor U19908 (N_19908,N_10510,N_10093);
or U19909 (N_19909,N_11343,N_10581);
nand U19910 (N_19910,N_13023,N_13182);
or U19911 (N_19911,N_14752,N_14638);
and U19912 (N_19912,N_11694,N_14036);
xor U19913 (N_19913,N_10970,N_14105);
and U19914 (N_19914,N_11678,N_13240);
nand U19915 (N_19915,N_10577,N_14671);
or U19916 (N_19916,N_14098,N_11962);
or U19917 (N_19917,N_10150,N_13144);
xnor U19918 (N_19918,N_13847,N_10054);
nor U19919 (N_19919,N_12752,N_11764);
and U19920 (N_19920,N_14501,N_13270);
nor U19921 (N_19921,N_13452,N_12448);
nor U19922 (N_19922,N_11166,N_11675);
xor U19923 (N_19923,N_11704,N_10697);
and U19924 (N_19924,N_10609,N_11581);
xnor U19925 (N_19925,N_11582,N_13375);
and U19926 (N_19926,N_13518,N_12503);
and U19927 (N_19927,N_13692,N_10768);
xnor U19928 (N_19928,N_10679,N_13179);
or U19929 (N_19929,N_10902,N_11958);
or U19930 (N_19930,N_14815,N_12283);
nor U19931 (N_19931,N_13789,N_11039);
or U19932 (N_19932,N_11038,N_14067);
xnor U19933 (N_19933,N_13939,N_11290);
xor U19934 (N_19934,N_12657,N_11731);
or U19935 (N_19935,N_10217,N_12290);
nand U19936 (N_19936,N_12786,N_11818);
or U19937 (N_19937,N_11929,N_14652);
nor U19938 (N_19938,N_10487,N_10143);
nand U19939 (N_19939,N_12280,N_10795);
or U19940 (N_19940,N_14678,N_10154);
and U19941 (N_19941,N_11047,N_11189);
and U19942 (N_19942,N_14159,N_12779);
nand U19943 (N_19943,N_13315,N_13489);
xor U19944 (N_19944,N_12525,N_10821);
and U19945 (N_19945,N_12258,N_11677);
and U19946 (N_19946,N_14492,N_12722);
nor U19947 (N_19947,N_12237,N_11920);
xor U19948 (N_19948,N_12165,N_13045);
or U19949 (N_19949,N_10851,N_12353);
xnor U19950 (N_19950,N_14398,N_12073);
and U19951 (N_19951,N_13085,N_12366);
xnor U19952 (N_19952,N_14938,N_13885);
and U19953 (N_19953,N_12450,N_12152);
xnor U19954 (N_19954,N_11696,N_10055);
or U19955 (N_19955,N_11377,N_11579);
nor U19956 (N_19956,N_10061,N_12864);
nor U19957 (N_19957,N_12234,N_14292);
nand U19958 (N_19958,N_11695,N_12794);
nand U19959 (N_19959,N_14863,N_13325);
xor U19960 (N_19960,N_12600,N_10491);
nand U19961 (N_19961,N_10103,N_10796);
xnor U19962 (N_19962,N_13644,N_14233);
and U19963 (N_19963,N_11538,N_10720);
nor U19964 (N_19964,N_12574,N_11479);
and U19965 (N_19965,N_12051,N_11503);
nand U19966 (N_19966,N_12969,N_13449);
xnor U19967 (N_19967,N_11031,N_10934);
nor U19968 (N_19968,N_11471,N_10182);
nand U19969 (N_19969,N_14878,N_12115);
xor U19970 (N_19970,N_14713,N_14862);
xor U19971 (N_19971,N_10027,N_10551);
and U19972 (N_19972,N_11578,N_12616);
and U19973 (N_19973,N_11635,N_13774);
nand U19974 (N_19974,N_14128,N_10604);
and U19975 (N_19975,N_14524,N_13766);
nor U19976 (N_19976,N_11414,N_12759);
nor U19977 (N_19977,N_12026,N_14324);
xor U19978 (N_19978,N_14749,N_11587);
nor U19979 (N_19979,N_11794,N_14136);
and U19980 (N_19980,N_13410,N_12780);
nor U19981 (N_19981,N_14016,N_10842);
nand U19982 (N_19982,N_13156,N_14095);
or U19983 (N_19983,N_14186,N_13929);
nor U19984 (N_19984,N_11304,N_14818);
and U19985 (N_19985,N_13462,N_14219);
nor U19986 (N_19986,N_14743,N_14370);
xnor U19987 (N_19987,N_11454,N_11018);
or U19988 (N_19988,N_11694,N_10937);
nor U19989 (N_19989,N_14947,N_14534);
and U19990 (N_19990,N_11651,N_10285);
nand U19991 (N_19991,N_12819,N_14293);
xor U19992 (N_19992,N_13348,N_13094);
and U19993 (N_19993,N_14183,N_14252);
nand U19994 (N_19994,N_12420,N_14208);
nand U19995 (N_19995,N_11634,N_11448);
nand U19996 (N_19996,N_10567,N_12343);
and U19997 (N_19997,N_12306,N_13465);
and U19998 (N_19998,N_12615,N_13831);
nor U19999 (N_19999,N_13092,N_12717);
nor U20000 (N_20000,N_18345,N_18416);
xnor U20001 (N_20001,N_19848,N_16662);
xnor U20002 (N_20002,N_19031,N_16121);
or U20003 (N_20003,N_15910,N_18055);
xor U20004 (N_20004,N_17263,N_16174);
or U20005 (N_20005,N_18157,N_15419);
nand U20006 (N_20006,N_16430,N_17866);
and U20007 (N_20007,N_18901,N_16023);
nor U20008 (N_20008,N_19711,N_19621);
xor U20009 (N_20009,N_18703,N_15523);
nand U20010 (N_20010,N_19782,N_19952);
nor U20011 (N_20011,N_15513,N_18717);
xor U20012 (N_20012,N_15722,N_16675);
nor U20013 (N_20013,N_15948,N_17771);
and U20014 (N_20014,N_17510,N_17923);
xor U20015 (N_20015,N_16288,N_17737);
nor U20016 (N_20016,N_16775,N_19875);
xnor U20017 (N_20017,N_15347,N_16927);
nand U20018 (N_20018,N_16556,N_16116);
nand U20019 (N_20019,N_15842,N_17566);
nor U20020 (N_20020,N_19077,N_16876);
xor U20021 (N_20021,N_17709,N_19399);
and U20022 (N_20022,N_19421,N_17700);
and U20023 (N_20023,N_15575,N_18760);
xor U20024 (N_20024,N_15705,N_19974);
nand U20025 (N_20025,N_16328,N_16141);
or U20026 (N_20026,N_15240,N_17909);
nand U20027 (N_20027,N_19430,N_19284);
nand U20028 (N_20028,N_19573,N_16567);
nand U20029 (N_20029,N_16364,N_19454);
or U20030 (N_20030,N_18212,N_15412);
and U20031 (N_20031,N_19027,N_17849);
nand U20032 (N_20032,N_16578,N_19617);
and U20033 (N_20033,N_16041,N_16710);
or U20034 (N_20034,N_15537,N_17169);
nand U20035 (N_20035,N_18814,N_16083);
xor U20036 (N_20036,N_19498,N_18040);
and U20037 (N_20037,N_15595,N_19096);
nor U20038 (N_20038,N_17026,N_19536);
xnor U20039 (N_20039,N_19802,N_18639);
and U20040 (N_20040,N_15304,N_16696);
nand U20041 (N_20041,N_19619,N_19339);
nand U20042 (N_20042,N_19938,N_18253);
nand U20043 (N_20043,N_17409,N_16924);
and U20044 (N_20044,N_15009,N_19458);
and U20045 (N_20045,N_16185,N_19721);
and U20046 (N_20046,N_18326,N_16469);
or U20047 (N_20047,N_18608,N_17388);
or U20048 (N_20048,N_18296,N_17405);
xnor U20049 (N_20049,N_18482,N_18089);
nor U20050 (N_20050,N_15225,N_15796);
and U20051 (N_20051,N_18561,N_16977);
xnor U20052 (N_20052,N_19372,N_18336);
or U20053 (N_20053,N_19423,N_18099);
and U20054 (N_20054,N_19086,N_19712);
xor U20055 (N_20055,N_17525,N_18074);
nand U20056 (N_20056,N_19507,N_16045);
nand U20057 (N_20057,N_17425,N_15132);
xor U20058 (N_20058,N_15971,N_17784);
or U20059 (N_20059,N_17432,N_17747);
and U20060 (N_20060,N_16758,N_15089);
and U20061 (N_20061,N_19715,N_16750);
nor U20062 (N_20062,N_17427,N_16978);
nor U20063 (N_20063,N_19590,N_19456);
xnor U20064 (N_20064,N_15039,N_16705);
and U20065 (N_20065,N_19940,N_16094);
xor U20066 (N_20066,N_15086,N_16511);
or U20067 (N_20067,N_16741,N_19744);
or U20068 (N_20068,N_15250,N_17777);
and U20069 (N_20069,N_15564,N_19116);
xnor U20070 (N_20070,N_19867,N_18420);
nor U20071 (N_20071,N_19969,N_19470);
and U20072 (N_20072,N_19831,N_17887);
nor U20073 (N_20073,N_17442,N_15552);
or U20074 (N_20074,N_15876,N_19413);
nor U20075 (N_20075,N_17318,N_16381);
or U20076 (N_20076,N_18949,N_18769);
nor U20077 (N_20077,N_16080,N_16579);
xor U20078 (N_20078,N_17103,N_19980);
or U20079 (N_20079,N_18110,N_16812);
or U20080 (N_20080,N_16767,N_19455);
xnor U20081 (N_20081,N_15596,N_19177);
nor U20082 (N_20082,N_18294,N_18105);
nand U20083 (N_20083,N_16995,N_15848);
nand U20084 (N_20084,N_15553,N_19883);
nor U20085 (N_20085,N_19179,N_17512);
nor U20086 (N_20086,N_16936,N_15047);
nor U20087 (N_20087,N_16058,N_15667);
nor U20088 (N_20088,N_15287,N_19231);
nand U20089 (N_20089,N_17038,N_17650);
xnor U20090 (N_20090,N_16335,N_16310);
xnor U20091 (N_20091,N_18875,N_17195);
or U20092 (N_20092,N_19864,N_17822);
xor U20093 (N_20093,N_18831,N_15181);
nand U20094 (N_20094,N_16265,N_19428);
nor U20095 (N_20095,N_19663,N_19502);
nor U20096 (N_20096,N_15407,N_16904);
xnor U20097 (N_20097,N_17679,N_18515);
or U20098 (N_20098,N_17443,N_17988);
xnor U20099 (N_20099,N_19305,N_18953);
and U20100 (N_20100,N_19923,N_15744);
and U20101 (N_20101,N_19679,N_19680);
nand U20102 (N_20102,N_19494,N_18232);
and U20103 (N_20103,N_16580,N_16882);
nand U20104 (N_20104,N_16745,N_15815);
and U20105 (N_20105,N_16458,N_18377);
nor U20106 (N_20106,N_16838,N_16703);
nand U20107 (N_20107,N_18268,N_16278);
or U20108 (N_20108,N_19288,N_19855);
or U20109 (N_20109,N_17548,N_17553);
xor U20110 (N_20110,N_18629,N_17785);
nor U20111 (N_20111,N_16197,N_17722);
nand U20112 (N_20112,N_16907,N_19095);
nand U20113 (N_20113,N_15014,N_19208);
and U20114 (N_20114,N_15103,N_15411);
nor U20115 (N_20115,N_19579,N_17502);
nand U20116 (N_20116,N_19996,N_19154);
or U20117 (N_20117,N_19566,N_19303);
xnor U20118 (N_20118,N_18596,N_16102);
xnor U20119 (N_20119,N_17825,N_18847);
or U20120 (N_20120,N_18026,N_15137);
and U20121 (N_20121,N_17326,N_18557);
and U20122 (N_20122,N_16901,N_15912);
nand U20123 (N_20123,N_17915,N_19337);
or U20124 (N_20124,N_16455,N_19894);
xnor U20125 (N_20125,N_19829,N_18250);
xor U20126 (N_20126,N_17963,N_18928);
or U20127 (N_20127,N_17082,N_17561);
xor U20128 (N_20128,N_18293,N_15024);
xnor U20129 (N_20129,N_15550,N_18886);
and U20130 (N_20130,N_16176,N_18239);
xnor U20131 (N_20131,N_19283,N_15594);
nand U20132 (N_20132,N_19635,N_17092);
xnor U20133 (N_20133,N_15882,N_18960);
or U20134 (N_20134,N_17515,N_18659);
and U20135 (N_20135,N_17691,N_15058);
and U20136 (N_20136,N_15237,N_19104);
xor U20137 (N_20137,N_18371,N_19534);
xnor U20138 (N_20138,N_17532,N_16358);
xor U20139 (N_20139,N_16735,N_17122);
and U20140 (N_20140,N_18910,N_18190);
and U20141 (N_20141,N_15380,N_16314);
xor U20142 (N_20142,N_16725,N_15975);
and U20143 (N_20143,N_17436,N_17213);
xor U20144 (N_20144,N_15269,N_17274);
or U20145 (N_20145,N_18564,N_16206);
xnor U20146 (N_20146,N_19261,N_18828);
and U20147 (N_20147,N_17652,N_19447);
and U20148 (N_20148,N_17005,N_15774);
xor U20149 (N_20149,N_19808,N_16896);
nor U20150 (N_20150,N_18255,N_17363);
or U20151 (N_20151,N_16478,N_16914);
and U20152 (N_20152,N_17007,N_15475);
nand U20153 (N_20153,N_15004,N_15308);
nor U20154 (N_20154,N_16600,N_17071);
xnor U20155 (N_20155,N_18327,N_16397);
xor U20156 (N_20156,N_19709,N_16963);
xor U20157 (N_20157,N_17661,N_19967);
and U20158 (N_20158,N_16437,N_18305);
and U20159 (N_20159,N_19134,N_18687);
and U20160 (N_20160,N_18600,N_17475);
nor U20161 (N_20161,N_18003,N_19748);
and U20162 (N_20162,N_19859,N_16866);
nand U20163 (N_20163,N_16602,N_15660);
and U20164 (N_20164,N_19331,N_19604);
or U20165 (N_20165,N_15914,N_15296);
or U20166 (N_20166,N_18675,N_18784);
or U20167 (N_20167,N_16378,N_15029);
nor U20168 (N_20168,N_18500,N_15453);
nor U20169 (N_20169,N_16454,N_15258);
or U20170 (N_20170,N_17114,N_17403);
xnor U20171 (N_20171,N_15630,N_19863);
nor U20172 (N_20172,N_19384,N_16755);
xnor U20173 (N_20173,N_19195,N_17659);
or U20174 (N_20174,N_17707,N_17831);
nand U20175 (N_20175,N_15054,N_16671);
and U20176 (N_20176,N_15434,N_18702);
xor U20177 (N_20177,N_15900,N_16188);
nand U20178 (N_20178,N_15316,N_17738);
or U20179 (N_20179,N_16574,N_18489);
nand U20180 (N_20180,N_15557,N_19238);
nand U20181 (N_20181,N_15471,N_18914);
or U20182 (N_20182,N_18501,N_19818);
and U20183 (N_20183,N_15694,N_16819);
nand U20184 (N_20184,N_18131,N_19559);
xor U20185 (N_20185,N_15042,N_19248);
and U20186 (N_20186,N_18033,N_19388);
nor U20187 (N_20187,N_15606,N_17145);
xnor U20188 (N_20188,N_18867,N_19176);
xnor U20189 (N_20189,N_17226,N_19106);
nand U20190 (N_20190,N_16944,N_18604);
and U20191 (N_20191,N_15941,N_17489);
xnor U20192 (N_20192,N_15916,N_18794);
nand U20193 (N_20193,N_18854,N_16740);
nor U20194 (N_20194,N_16443,N_17015);
and U20195 (N_20195,N_16404,N_16809);
and U20196 (N_20196,N_18559,N_16193);
nor U20197 (N_20197,N_19210,N_17762);
xnor U20198 (N_20198,N_17615,N_16958);
xor U20199 (N_20199,N_18699,N_18865);
nand U20200 (N_20200,N_19737,N_16425);
or U20201 (N_20201,N_15260,N_16692);
nand U20202 (N_20202,N_19196,N_19939);
nor U20203 (N_20203,N_16731,N_17695);
nand U20204 (N_20204,N_17225,N_19278);
or U20205 (N_20205,N_18850,N_18350);
or U20206 (N_20206,N_17046,N_18050);
nor U20207 (N_20207,N_19508,N_17074);
nor U20208 (N_20208,N_18355,N_15979);
nand U20209 (N_20209,N_16349,N_18285);
xor U20210 (N_20210,N_17928,N_17060);
or U20211 (N_20211,N_19243,N_19274);
nand U20212 (N_20212,N_17578,N_15442);
and U20213 (N_20213,N_16969,N_17338);
nor U20214 (N_20214,N_19697,N_17540);
nand U20215 (N_20215,N_16402,N_18488);
or U20216 (N_20216,N_19794,N_18085);
nand U20217 (N_20217,N_17730,N_19783);
or U20218 (N_20218,N_18307,N_17829);
and U20219 (N_20219,N_18973,N_18452);
or U20220 (N_20220,N_18548,N_15091);
or U20221 (N_20221,N_18918,N_15644);
nand U20222 (N_20222,N_16150,N_16405);
xor U20223 (N_20223,N_16672,N_19011);
nor U20224 (N_20224,N_15708,N_17669);
nor U20225 (N_20225,N_18696,N_19004);
and U20226 (N_20226,N_17876,N_19126);
xor U20227 (N_20227,N_19541,N_18676);
nand U20228 (N_20228,N_19913,N_18047);
and U20229 (N_20229,N_19580,N_15886);
nand U20230 (N_20230,N_17451,N_17976);
xor U20231 (N_20231,N_15546,N_18933);
nor U20232 (N_20232,N_17830,N_19739);
nand U20233 (N_20233,N_19899,N_15239);
xnor U20234 (N_20234,N_16148,N_15362);
or U20235 (N_20235,N_16067,N_16024);
nor U20236 (N_20236,N_15271,N_18861);
nor U20237 (N_20237,N_19771,N_15893);
nor U20238 (N_20238,N_15952,N_19067);
nor U20239 (N_20239,N_18383,N_17729);
xor U20240 (N_20240,N_19268,N_15885);
or U20241 (N_20241,N_15970,N_19395);
and U20242 (N_20242,N_15289,N_16620);
xnor U20243 (N_20243,N_17025,N_17841);
nand U20244 (N_20244,N_16363,N_16413);
nand U20245 (N_20245,N_16689,N_19091);
and U20246 (N_20246,N_19553,N_16903);
xnor U20247 (N_20247,N_15802,N_18185);
and U20248 (N_20248,N_15603,N_19595);
xor U20249 (N_20249,N_16064,N_19693);
and U20250 (N_20250,N_15996,N_16260);
nor U20251 (N_20251,N_17073,N_19120);
nor U20252 (N_20252,N_18147,N_17401);
nor U20253 (N_20253,N_19902,N_18691);
xor U20254 (N_20254,N_17477,N_19074);
xnor U20255 (N_20255,N_19018,N_19620);
nor U20256 (N_20256,N_15932,N_18922);
xnor U20257 (N_20257,N_15593,N_17522);
nand U20258 (N_20258,N_18481,N_15637);
and U20259 (N_20259,N_19526,N_16270);
or U20260 (N_20260,N_15457,N_16048);
xnor U20261 (N_20261,N_16302,N_15843);
nand U20262 (N_20262,N_15211,N_17224);
nor U20263 (N_20263,N_17488,N_15006);
or U20264 (N_20264,N_16274,N_17415);
or U20265 (N_20265,N_17386,N_17437);
nor U20266 (N_20266,N_18808,N_16322);
xor U20267 (N_20267,N_18491,N_16918);
nand U20268 (N_20268,N_17311,N_17462);
xor U20269 (N_20269,N_16249,N_19719);
or U20270 (N_20270,N_17797,N_16716);
xnor U20271 (N_20271,N_16514,N_18889);
or U20272 (N_20272,N_17343,N_16658);
xnor U20273 (N_20273,N_15819,N_15653);
nand U20274 (N_20274,N_17420,N_16594);
and U20275 (N_20275,N_16124,N_18267);
or U20276 (N_20276,N_16611,N_16037);
xnor U20277 (N_20277,N_17296,N_16075);
xnor U20278 (N_20278,N_16138,N_16486);
and U20279 (N_20279,N_16199,N_17003);
nand U20280 (N_20280,N_15389,N_19189);
nand U20281 (N_20281,N_18112,N_15410);
and U20282 (N_20282,N_17971,N_16244);
and U20283 (N_20283,N_16329,N_19797);
nand U20284 (N_20284,N_16475,N_19618);
nor U20285 (N_20285,N_19518,N_15465);
xnor U20286 (N_20286,N_19460,N_19493);
nand U20287 (N_20287,N_18537,N_19503);
or U20288 (N_20288,N_15018,N_15884);
or U20289 (N_20289,N_19695,N_18401);
xnor U20290 (N_20290,N_15915,N_15549);
and U20291 (N_20291,N_19049,N_18408);
or U20292 (N_20292,N_15727,N_18181);
nor U20293 (N_20293,N_18031,N_18762);
and U20294 (N_20294,N_16590,N_19515);
and U20295 (N_20295,N_17643,N_17336);
xor U20296 (N_20296,N_16247,N_19954);
nor U20297 (N_20297,N_18980,N_19167);
nand U20298 (N_20298,N_17516,N_18014);
nand U20299 (N_20299,N_18011,N_18028);
and U20300 (N_20300,N_16756,N_15711);
nand U20301 (N_20301,N_17799,N_16836);
nand U20302 (N_20302,N_16572,N_17470);
and U20303 (N_20303,N_19474,N_19240);
nand U20304 (N_20304,N_15157,N_17396);
nand U20305 (N_20305,N_18096,N_15439);
nand U20306 (N_20306,N_16240,N_19482);
xor U20307 (N_20307,N_19191,N_16316);
or U20308 (N_20308,N_19706,N_17593);
nand U20309 (N_20309,N_19173,N_16615);
and U20310 (N_20310,N_18988,N_15934);
nor U20311 (N_20311,N_15195,N_19997);
nor U20312 (N_20312,N_16742,N_18091);
or U20313 (N_20313,N_16976,N_15298);
xor U20314 (N_20314,N_17259,N_19778);
xnor U20315 (N_20315,N_19634,N_16828);
nor U20316 (N_20316,N_16863,N_18137);
or U20317 (N_20317,N_15045,N_15219);
or U20318 (N_20318,N_18480,N_19277);
and U20319 (N_20319,N_19381,N_17180);
xor U20320 (N_20320,N_17057,N_16427);
or U20321 (N_20321,N_17332,N_18194);
xnor U20322 (N_20322,N_19731,N_19033);
or U20323 (N_20323,N_15251,N_16899);
xor U20324 (N_20324,N_17345,N_18220);
and U20325 (N_20325,N_19492,N_17791);
nor U20326 (N_20326,N_19057,N_18492);
or U20327 (N_20327,N_18843,N_16779);
nand U20328 (N_20328,N_15128,N_17204);
or U20329 (N_20329,N_16444,N_17733);
nand U20330 (N_20330,N_18499,N_17239);
xor U20331 (N_20331,N_18923,N_16849);
and U20332 (N_20332,N_19266,N_16186);
xnor U20333 (N_20333,N_16479,N_17146);
or U20334 (N_20334,N_16218,N_15203);
nand U20335 (N_20335,N_18810,N_19042);
and U20336 (N_20336,N_19574,N_18739);
or U20337 (N_20337,N_16312,N_17858);
nor U20338 (N_20338,N_18102,N_19486);
and U20339 (N_20339,N_19982,N_17769);
nor U20340 (N_20340,N_16563,N_16338);
nand U20341 (N_20341,N_16081,N_17466);
nand U20342 (N_20342,N_15095,N_16362);
and U20343 (N_20343,N_18568,N_19107);
xnor U20344 (N_20344,N_17133,N_17222);
or U20345 (N_20345,N_19187,N_17148);
nand U20346 (N_20346,N_17938,N_15627);
or U20347 (N_20347,N_17585,N_17511);
or U20348 (N_20348,N_18913,N_15720);
xor U20349 (N_20349,N_17247,N_19038);
nand U20350 (N_20350,N_16902,N_16575);
and U20351 (N_20351,N_16179,N_17151);
or U20352 (N_20352,N_16588,N_17616);
xnor U20353 (N_20353,N_18799,N_16182);
xor U20354 (N_20354,N_18970,N_16348);
and U20355 (N_20355,N_18330,N_15182);
xnor U20356 (N_20356,N_15671,N_16679);
xnor U20357 (N_20357,N_15762,N_17803);
and U20358 (N_20358,N_19965,N_17605);
xor U20359 (N_20359,N_18978,N_16399);
nor U20360 (N_20360,N_17818,N_18990);
xor U20361 (N_20361,N_16554,N_16929);
or U20362 (N_20362,N_15124,N_19162);
nor U20363 (N_20363,N_18882,N_19365);
nand U20364 (N_20364,N_17235,N_19254);
xnor U20365 (N_20365,N_15282,N_18007);
xor U20366 (N_20366,N_17586,N_19908);
nor U20367 (N_20367,N_17921,N_15960);
nor U20368 (N_20368,N_18378,N_15535);
nand U20369 (N_20369,N_16212,N_18313);
xor U20370 (N_20370,N_19583,N_16057);
and U20371 (N_20371,N_17991,N_17061);
nor U20372 (N_20372,N_17482,N_18016);
xor U20373 (N_20373,N_18898,N_15052);
or U20374 (N_20374,N_16090,N_18376);
nor U20375 (N_20375,N_18167,N_19698);
xnor U20376 (N_20376,N_16625,N_16543);
nor U20377 (N_20377,N_18362,N_17016);
and U20378 (N_20378,N_18486,N_19289);
nand U20379 (N_20379,N_19669,N_18211);
and U20380 (N_20380,N_19202,N_15277);
nand U20381 (N_20381,N_18547,N_17383);
xnor U20382 (N_20382,N_16885,N_18792);
nand U20383 (N_20383,N_15267,N_17757);
nand U20384 (N_20384,N_19605,N_17251);
nand U20385 (N_20385,N_16926,N_16595);
or U20386 (N_20386,N_17968,N_18752);
nand U20387 (N_20387,N_15143,N_18614);
or U20388 (N_20388,N_17983,N_16386);
and U20389 (N_20389,N_18858,N_15992);
and U20390 (N_20390,N_17790,N_16493);
or U20391 (N_20391,N_18974,N_15082);
and U20392 (N_20392,N_16304,N_18780);
or U20393 (N_20393,N_16237,N_15878);
nor U20394 (N_20394,N_16773,N_16714);
xor U20395 (N_20395,N_15490,N_17198);
or U20396 (N_20396,N_15395,N_16101);
nor U20397 (N_20397,N_16521,N_18409);
nand U20398 (N_20398,N_15171,N_17844);
nor U20399 (N_20399,N_16718,N_16177);
xor U20400 (N_20400,N_18292,N_15418);
and U20401 (N_20401,N_18763,N_18952);
or U20402 (N_20402,N_17644,N_18588);
xor U20403 (N_20403,N_15591,N_17211);
and U20404 (N_20404,N_19054,N_17568);
or U20405 (N_20405,N_15937,N_16825);
or U20406 (N_20406,N_16181,N_17233);
nand U20407 (N_20407,N_17013,N_16568);
nor U20408 (N_20408,N_19757,N_17666);
xnor U20409 (N_20409,N_17055,N_19119);
nand U20410 (N_20410,N_15619,N_17348);
nand U20411 (N_20411,N_15373,N_17164);
or U20412 (N_20412,N_16988,N_18123);
or U20413 (N_20413,N_19045,N_17816);
or U20414 (N_20414,N_16009,N_15738);
or U20415 (N_20415,N_17600,N_16311);
xor U20416 (N_20416,N_19557,N_17970);
xnor U20417 (N_20417,N_16467,N_16173);
xor U20418 (N_20418,N_18654,N_19844);
and U20419 (N_20419,N_18463,N_18361);
nand U20420 (N_20420,N_17189,N_17723);
or U20421 (N_20421,N_18522,N_17717);
or U20422 (N_20422,N_15943,N_16034);
nor U20423 (N_20423,N_15767,N_15567);
and U20424 (N_20424,N_17767,N_16752);
xnor U20425 (N_20425,N_17842,N_18874);
xor U20426 (N_20426,N_18335,N_15002);
nand U20427 (N_20427,N_16688,N_17072);
nor U20428 (N_20428,N_15639,N_15822);
nor U20429 (N_20429,N_17414,N_15431);
nand U20430 (N_20430,N_18902,N_18385);
or U20431 (N_20431,N_17152,N_18410);
xnor U20432 (N_20432,N_19761,N_15577);
and U20433 (N_20433,N_18215,N_18636);
nor U20434 (N_20434,N_17130,N_18349);
and U20435 (N_20435,N_16373,N_19714);
nand U20436 (N_20436,N_15944,N_19007);
nand U20437 (N_20437,N_17335,N_15334);
xor U20438 (N_20438,N_15984,N_16571);
nand U20439 (N_20439,N_15894,N_17187);
xor U20440 (N_20440,N_16233,N_15413);
xnor U20441 (N_20441,N_15655,N_16269);
nand U20442 (N_20442,N_17051,N_15645);
nor U20443 (N_20443,N_18041,N_19009);
xnor U20444 (N_20444,N_15750,N_19514);
xnor U20445 (N_20445,N_16431,N_19571);
and U20446 (N_20446,N_17531,N_18516);
nand U20447 (N_20447,N_16162,N_15860);
xor U20448 (N_20448,N_15766,N_15468);
nor U20449 (N_20449,N_18878,N_18958);
or U20450 (N_20450,N_17182,N_16711);
and U20451 (N_20451,N_16137,N_18994);
or U20452 (N_20452,N_16895,N_15071);
nor U20453 (N_20453,N_19576,N_17624);
xnor U20454 (N_20454,N_18414,N_16930);
xnor U20455 (N_20455,N_18530,N_18407);
and U20456 (N_20456,N_16236,N_16076);
xnor U20457 (N_20457,N_16423,N_18161);
nor U20458 (N_20458,N_15336,N_18075);
or U20459 (N_20459,N_17932,N_17395);
or U20460 (N_20460,N_19710,N_19296);
and U20461 (N_20461,N_18969,N_15174);
nand U20462 (N_20462,N_15017,N_19759);
or U20463 (N_20463,N_18068,N_15193);
xor U20464 (N_20464,N_16131,N_15066);
or U20465 (N_20465,N_17351,N_19551);
or U20466 (N_20466,N_19876,N_16051);
xnor U20467 (N_20467,N_17091,N_19249);
nand U20468 (N_20468,N_18817,N_17285);
and U20469 (N_20469,N_19889,N_19358);
and U20470 (N_20470,N_19570,N_16981);
xnor U20471 (N_20471,N_19080,N_19427);
xor U20472 (N_20472,N_18299,N_18004);
and U20473 (N_20473,N_18248,N_16585);
and U20474 (N_20474,N_16518,N_18712);
nand U20475 (N_20475,N_19310,N_15922);
nor U20476 (N_20476,N_17583,N_19951);
or U20477 (N_20477,N_16693,N_19419);
and U20478 (N_20478,N_17557,N_18263);
or U20479 (N_20479,N_19985,N_15392);
or U20480 (N_20480,N_18719,N_17885);
xor U20481 (N_20481,N_19849,N_17746);
or U20482 (N_20482,N_16350,N_15828);
xor U20483 (N_20483,N_15909,N_18101);
xnor U20484 (N_20484,N_18938,N_17127);
nor U20485 (N_20485,N_17813,N_18511);
or U20486 (N_20486,N_18742,N_19724);
and U20487 (N_20487,N_18174,N_16935);
xor U20488 (N_20488,N_17307,N_15617);
or U20489 (N_20489,N_16219,N_16547);
nor U20490 (N_20490,N_18896,N_17337);
nand U20491 (N_20491,N_17109,N_15273);
nand U20492 (N_20492,N_16320,N_19836);
and U20493 (N_20493,N_15949,N_15479);
xnor U20494 (N_20494,N_18987,N_16529);
and U20495 (N_20495,N_16898,N_15683);
nor U20496 (N_20496,N_17174,N_18643);
nor U20497 (N_20497,N_18162,N_17562);
nor U20498 (N_20498,N_17939,N_19260);
or U20499 (N_20499,N_15859,N_18158);
xnor U20500 (N_20500,N_16354,N_18054);
and U20501 (N_20501,N_17163,N_16577);
or U20502 (N_20502,N_18713,N_18044);
or U20503 (N_20503,N_17249,N_19993);
and U20504 (N_20504,N_16496,N_16852);
xor U20505 (N_20505,N_17366,N_19665);
nor U20506 (N_20506,N_19313,N_16721);
nor U20507 (N_20507,N_19804,N_16729);
nand U20508 (N_20508,N_17119,N_15343);
xor U20509 (N_20509,N_18171,N_19528);
nand U20510 (N_20510,N_19340,N_18768);
nand U20511 (N_20511,N_19144,N_15135);
nand U20512 (N_20512,N_19642,N_16229);
or U20513 (N_20513,N_19151,N_19070);
nand U20514 (N_20514,N_16071,N_15437);
nor U20515 (N_20515,N_17854,N_15167);
xnor U20516 (N_20516,N_15090,N_18015);
and U20517 (N_20517,N_18417,N_15424);
and U20518 (N_20518,N_15699,N_15152);
nor U20519 (N_20519,N_15543,N_18322);
and U20520 (N_20520,N_16743,N_15070);
nand U20521 (N_20521,N_16307,N_15825);
xor U20522 (N_20522,N_15514,N_16843);
xor U20523 (N_20523,N_18478,N_15209);
nand U20524 (N_20524,N_15742,N_15175);
or U20525 (N_20525,N_16604,N_17868);
and U20526 (N_20526,N_17209,N_18388);
nor U20527 (N_20527,N_15365,N_16343);
nand U20528 (N_20528,N_15458,N_18440);
xnor U20529 (N_20529,N_15811,N_16516);
nand U20530 (N_20530,N_18072,N_18531);
xor U20531 (N_20531,N_17856,N_16428);
nand U20532 (N_20532,N_16847,N_19856);
nor U20533 (N_20533,N_17535,N_18804);
or U20534 (N_20534,N_15093,N_17676);
or U20535 (N_20535,N_19275,N_17865);
nor U20536 (N_20536,N_19821,N_17892);
or U20537 (N_20537,N_16488,N_17647);
nor U20538 (N_20538,N_15281,N_16078);
or U20539 (N_20539,N_16873,N_19575);
xnor U20540 (N_20540,N_15721,N_19935);
or U20541 (N_20541,N_19262,N_17863);
nand U20542 (N_20542,N_18733,N_16539);
and U20543 (N_20543,N_17284,N_18093);
xor U20544 (N_20544,N_17875,N_18855);
nand U20545 (N_20545,N_15651,N_15544);
nand U20546 (N_20546,N_19853,N_18453);
or U20547 (N_20547,N_17083,N_19568);
xor U20548 (N_20548,N_18372,N_15133);
xor U20549 (N_20549,N_17677,N_18037);
nand U20550 (N_20550,N_15746,N_18609);
nand U20551 (N_20551,N_18256,N_16874);
and U20552 (N_20552,N_15151,N_19718);
xor U20553 (N_20553,N_16991,N_16570);
nor U20554 (N_20554,N_17178,N_19907);
nor U20555 (N_20555,N_18776,N_16528);
and U20556 (N_20556,N_19694,N_19563);
or U20557 (N_20557,N_17408,N_18183);
nor U20558 (N_20558,N_19677,N_17683);
or U20559 (N_20559,N_16168,N_18485);
and U20560 (N_20560,N_18318,N_16490);
and U20561 (N_20561,N_17308,N_15771);
and U20562 (N_20562,N_19449,N_17397);
and U20563 (N_20563,N_15806,N_15657);
or U20564 (N_20564,N_15116,N_18700);
nand U20565 (N_20565,N_16189,N_18427);
xor U20566 (N_20566,N_17852,N_19688);
or U20567 (N_20567,N_15989,N_15556);
or U20568 (N_20568,N_17845,N_16336);
xor U20569 (N_20569,N_17468,N_18118);
and U20570 (N_20570,N_15980,N_17521);
xor U20571 (N_20571,N_19942,N_15920);
nor U20572 (N_20572,N_18580,N_16256);
and U20573 (N_20573,N_17523,N_17798);
and U20574 (N_20574,N_18711,N_19885);
or U20575 (N_20575,N_19496,N_15154);
nand U20576 (N_20576,N_18748,N_16861);
xnor U20577 (N_20577,N_19682,N_18800);
or U20578 (N_20578,N_16359,N_15685);
nor U20579 (N_20579,N_17040,N_19966);
or U20580 (N_20580,N_18127,N_19309);
and U20581 (N_20581,N_16530,N_15677);
or U20582 (N_20582,N_18661,N_19717);
and U20583 (N_20583,N_16195,N_18231);
and U20584 (N_20584,N_17269,N_15732);
nand U20585 (N_20585,N_18467,N_19445);
nand U20586 (N_20586,N_18944,N_16115);
and U20587 (N_20587,N_16650,N_16424);
nor U20588 (N_20588,N_19847,N_18346);
or U20589 (N_20589,N_19976,N_16897);
or U20590 (N_20590,N_15686,N_19562);
xor U20591 (N_20591,N_15108,N_16802);
and U20592 (N_20592,N_18397,N_18701);
nor U20593 (N_20593,N_15724,N_18806);
xor U20594 (N_20594,N_17480,N_18698);
nor U20595 (N_20595,N_15508,N_15274);
xor U20596 (N_20596,N_17256,N_18877);
and U20597 (N_20597,N_18668,N_17411);
and U20598 (N_20598,N_16789,N_15228);
nand U20599 (N_20599,N_19652,N_16638);
or U20600 (N_20600,N_18718,N_15986);
nor U20601 (N_20601,N_15033,N_15578);
nand U20602 (N_20602,N_19886,N_15364);
nor U20603 (N_20603,N_17879,N_15307);
and U20604 (N_20604,N_16133,N_18280);
and U20605 (N_20605,N_18906,N_18544);
nand U20606 (N_20606,N_19433,N_19334);
or U20607 (N_20607,N_16548,N_19659);
nor U20608 (N_20608,N_15499,N_17279);
nor U20609 (N_20609,N_16313,N_16028);
or U20610 (N_20610,N_15626,N_18603);
nor U20611 (N_20611,N_18226,N_17126);
and U20612 (N_20612,N_19699,N_16442);
nor U20613 (N_20613,N_15879,N_17157);
nor U20614 (N_20614,N_17066,N_18502);
xor U20615 (N_20615,N_17254,N_15393);
nor U20616 (N_20616,N_16107,N_15755);
or U20617 (N_20617,N_16817,N_16837);
nor U20618 (N_20618,N_16295,N_16410);
or U20619 (N_20619,N_18724,N_17393);
nand U20620 (N_20620,N_16132,N_18690);
or U20621 (N_20621,N_19352,N_15020);
or U20622 (N_20622,N_16792,N_19992);
nand U20623 (N_20623,N_18429,N_19397);
or U20624 (N_20624,N_15104,N_17619);
xor U20625 (N_20625,N_15291,N_18389);
and U20626 (N_20626,N_15445,N_15302);
nor U20627 (N_20627,N_15566,N_16125);
xnor U20628 (N_20628,N_16283,N_16139);
or U20629 (N_20629,N_19168,N_15861);
xnor U20630 (N_20630,N_18080,N_19950);
nor U20631 (N_20631,N_18968,N_18442);
nor U20632 (N_20632,N_19668,N_17592);
xnor U20633 (N_20633,N_16535,N_15688);
and U20634 (N_20634,N_18298,N_17449);
xnor U20635 (N_20635,N_16786,N_16119);
and U20636 (N_20636,N_19893,N_16617);
and U20637 (N_20637,N_16673,N_15185);
and U20638 (N_20638,N_16726,N_15658);
or U20639 (N_20639,N_17020,N_17917);
xor U20640 (N_20640,N_18144,N_17686);
nor U20641 (N_20641,N_15177,N_15656);
or U20642 (N_20642,N_18084,N_16993);
nand U20643 (N_20643,N_15235,N_18967);
nor U20644 (N_20644,N_18605,N_17612);
xor U20645 (N_20645,N_17725,N_18747);
xor U20646 (N_20646,N_17238,N_19307);
or U20647 (N_20647,N_15643,N_18034);
and U20648 (N_20648,N_18295,N_16109);
xnor U20649 (N_20649,N_18672,N_16190);
or U20650 (N_20650,N_18807,N_15923);
or U20651 (N_20651,N_18943,N_19174);
xnor U20652 (N_20652,N_19606,N_16723);
nand U20653 (N_20653,N_15398,N_18270);
nor U20654 (N_20654,N_19860,N_18618);
or U20655 (N_20655,N_18862,N_16416);
or U20656 (N_20656,N_17713,N_18077);
nand U20657 (N_20657,N_17448,N_19929);
and U20658 (N_20658,N_19084,N_18575);
xnor U20659 (N_20659,N_17004,N_19314);
xnor U20660 (N_20660,N_18168,N_19285);
nor U20661 (N_20661,N_15161,N_17372);
and U20662 (N_20662,N_18424,N_16583);
nor U20663 (N_20663,N_19653,N_17620);
xnor U20664 (N_20664,N_17871,N_17193);
or U20665 (N_20665,N_19491,N_19851);
nand U20666 (N_20666,N_15217,N_19128);
xor U20667 (N_20667,N_18199,N_16647);
xor U20668 (N_20668,N_15214,N_16146);
and U20669 (N_20669,N_16216,N_17710);
and U20670 (N_20670,N_15509,N_16739);
xor U20671 (N_20671,N_19556,N_15201);
nand U20672 (N_20672,N_16674,N_15852);
and U20673 (N_20673,N_18686,N_19905);
xnor U20674 (N_20674,N_18798,N_17430);
and U20675 (N_20675,N_16450,N_16909);
or U20676 (N_20676,N_15725,N_16781);
xnor U20677 (N_20677,N_16161,N_16072);
nor U20678 (N_20678,N_15252,N_18272);
nor U20679 (N_20679,N_15080,N_17670);
and U20680 (N_20680,N_17667,N_17356);
or U20681 (N_20681,N_16446,N_15197);
or U20682 (N_20682,N_18281,N_15710);
xor U20683 (N_20683,N_19141,N_16565);
nand U20684 (N_20684,N_15075,N_16821);
xnor U20685 (N_20685,N_15779,N_17590);
xnor U20686 (N_20686,N_17471,N_15600);
and U20687 (N_20687,N_17253,N_18036);
and U20688 (N_20688,N_15121,N_15496);
or U20689 (N_20689,N_19100,N_18543);
and U20690 (N_20690,N_16347,N_16073);
or U20691 (N_20691,N_15814,N_15801);
nand U20692 (N_20692,N_16297,N_15841);
nand U20693 (N_20693,N_19158,N_18087);
nand U20694 (N_20694,N_15753,N_15472);
nand U20695 (N_20695,N_18140,N_15872);
xnor U20696 (N_20696,N_19544,N_17293);
and U20697 (N_20697,N_16344,N_15056);
nor U20698 (N_20698,N_15976,N_18598);
nand U20699 (N_20699,N_15034,N_19672);
xor U20700 (N_20700,N_18051,N_15330);
or U20701 (N_20701,N_17904,N_15297);
nand U20702 (N_20702,N_18904,N_19034);
and U20703 (N_20703,N_16652,N_18848);
nor U20704 (N_20704,N_19040,N_18984);
and U20705 (N_20705,N_18254,N_15520);
or U20706 (N_20706,N_15938,N_15117);
and U20707 (N_20707,N_16601,N_18986);
or U20708 (N_20708,N_17215,N_15001);
nand U20709 (N_20709,N_16134,N_19921);
nand U20710 (N_20710,N_19259,N_18321);
nand U20711 (N_20711,N_18823,N_16560);
xor U20712 (N_20712,N_19527,N_17602);
nor U20713 (N_20713,N_15763,N_19988);
nor U20714 (N_20714,N_18146,N_18338);
nor U20715 (N_20715,N_15510,N_16167);
nand U20716 (N_20716,N_19843,N_18444);
nor U20717 (N_20717,N_19046,N_16239);
xor U20718 (N_20718,N_15638,N_19366);
xor U20719 (N_20719,N_15569,N_19704);
or U20720 (N_20720,N_15172,N_17435);
or U20721 (N_20721,N_17481,N_18785);
xnor U20722 (N_20722,N_19393,N_16463);
and U20723 (N_20723,N_18065,N_19175);
nor U20724 (N_20724,N_19110,N_16844);
nand U20725 (N_20725,N_17258,N_18628);
and U20726 (N_20726,N_15110,N_18852);
xor U20727 (N_20727,N_15669,N_15040);
and U20728 (N_20728,N_18956,N_17870);
nand U20729 (N_20729,N_15858,N_18461);
or U20730 (N_20730,N_17966,N_15790);
xnor U20731 (N_20731,N_16122,N_16200);
or U20732 (N_20732,N_15945,N_15690);
nor U20733 (N_20733,N_15118,N_16749);
xnor U20734 (N_20734,N_17701,N_17538);
or U20735 (N_20735,N_19845,N_15311);
and U20736 (N_20736,N_15332,N_18098);
nor U20737 (N_20737,N_18340,N_16114);
and U20738 (N_20738,N_17069,N_17271);
nand U20739 (N_20739,N_15497,N_15028);
and U20740 (N_20740,N_17095,N_19150);
and U20741 (N_20741,N_17859,N_19183);
and U20742 (N_20742,N_17431,N_16418);
xor U20743 (N_20743,N_16782,N_17552);
or U20744 (N_20744,N_19287,N_19394);
xor U20745 (N_20745,N_16306,N_15032);
nor U20746 (N_20746,N_19359,N_17776);
nand U20747 (N_20747,N_17520,N_19180);
nand U20748 (N_20748,N_19983,N_18526);
xor U20749 (N_20749,N_16184,N_16271);
or U20750 (N_20750,N_18069,N_18435);
xor U20751 (N_20751,N_16355,N_18957);
xor U20752 (N_20752,N_15588,N_18134);
and U20753 (N_20753,N_15506,N_16962);
xor U20754 (N_20754,N_17257,N_19097);
nor U20755 (N_20755,N_19764,N_16651);
xnor U20756 (N_20756,N_18940,N_18457);
and U20757 (N_20757,N_17246,N_19006);
nand U20758 (N_20758,N_18527,N_15830);
nand U20759 (N_20759,N_16085,N_15820);
and U20760 (N_20760,N_19071,N_17281);
nand U20761 (N_20761,N_16648,N_18258);
or U20762 (N_20762,N_16420,N_19140);
or U20763 (N_20763,N_15730,N_16736);
nand U20764 (N_20764,N_16762,N_15839);
or U20765 (N_20765,N_16803,N_17277);
nor U20766 (N_20766,N_15850,N_19169);
xor U20767 (N_20767,N_16145,N_16815);
nor U20768 (N_20768,N_18704,N_16561);
or U20769 (N_20769,N_16810,N_15318);
nor U20770 (N_20770,N_16751,N_19660);
or U20771 (N_20771,N_15101,N_17651);
nor U20772 (N_20772,N_18018,N_19751);
and U20773 (N_20773,N_19509,N_17260);
and U20774 (N_20774,N_16489,N_15610);
nand U20775 (N_20775,N_18216,N_17526);
and U20776 (N_20776,N_17890,N_15581);
nand U20777 (N_20777,N_16923,N_16152);
or U20778 (N_20778,N_16717,N_19295);
xnor U20779 (N_20779,N_16629,N_15069);
nand U20780 (N_20780,N_18403,N_19832);
or U20781 (N_20781,N_17899,N_15043);
or U20782 (N_20782,N_18121,N_15012);
and U20783 (N_20783,N_17565,N_19505);
or U20784 (N_20784,N_16939,N_15565);
and U20785 (N_20785,N_17749,N_16656);
xor U20786 (N_20786,N_15718,N_19755);
nand U20787 (N_20787,N_17081,N_16111);
nand U20788 (N_20788,N_17929,N_16613);
nand U20789 (N_20789,N_18916,N_19589);
nand U20790 (N_20790,N_15887,N_15706);
nand U20791 (N_20791,N_18597,N_16769);
xor U20792 (N_20792,N_16032,N_17627);
xor U20793 (N_20793,N_16610,N_17668);
nor U20794 (N_20794,N_16784,N_18507);
xnor U20795 (N_20795,N_16321,N_16558);
nor U20796 (N_20796,N_17457,N_19255);
xor U20797 (N_20797,N_19085,N_15461);
nor U20798 (N_20798,N_17792,N_15249);
nor U20799 (N_20799,N_15085,N_16070);
xor U20800 (N_20800,N_15625,N_18135);
nand U20801 (N_20801,N_16449,N_15844);
or U20802 (N_20802,N_19880,N_18271);
nor U20803 (N_20803,N_15968,N_18781);
xnor U20804 (N_20804,N_18663,N_18632);
xor U20805 (N_20805,N_18851,N_16056);
xor U20806 (N_20806,N_16841,N_16532);
nand U20807 (N_20807,N_18309,N_17375);
nand U20808 (N_20808,N_16263,N_19994);
nand U20809 (N_20809,N_15464,N_17077);
nor U20810 (N_20810,N_17160,N_16222);
nand U20811 (N_20811,N_16733,N_18459);
xor U20812 (N_20812,N_16842,N_18819);
xor U20813 (N_20813,N_15366,N_17349);
nand U20814 (N_20814,N_18242,N_17546);
xor U20815 (N_20815,N_18539,N_19000);
xnor U20816 (N_20816,N_18822,N_19131);
nand U20817 (N_20817,N_19917,N_17847);
and U20818 (N_20818,N_19615,N_19858);
nor U20819 (N_20819,N_19933,N_18616);
nand U20820 (N_20820,N_18057,N_19800);
nor U20821 (N_20821,N_15786,N_15036);
or U20822 (N_20822,N_19519,N_19549);
or U20823 (N_20823,N_18224,N_17551);
xnor U20824 (N_20824,N_16018,N_19752);
nor U20825 (N_20825,N_18128,N_19117);
xor U20826 (N_20826,N_17969,N_16156);
nand U20827 (N_20827,N_18514,N_17878);
and U20828 (N_20828,N_15597,N_15913);
and U20829 (N_20829,N_19250,N_17387);
or U20830 (N_20830,N_15372,N_16388);
nor U20831 (N_20831,N_17702,N_19172);
or U20832 (N_20832,N_17604,N_15760);
xnor U20833 (N_20833,N_16129,N_15122);
nor U20834 (N_20834,N_17705,N_18642);
nor U20835 (N_20835,N_15173,N_16401);
xor U20836 (N_20836,N_17699,N_18497);
nor U20837 (N_20837,N_17171,N_18965);
nor U20838 (N_20838,N_19934,N_16171);
and U20839 (N_20839,N_17452,N_18450);
xnor U20840 (N_20840,N_15276,N_16598);
nor U20841 (N_20841,N_16906,N_16207);
nand U20842 (N_20842,N_19654,N_15019);
xnor U20843 (N_20843,N_19914,N_18551);
nor U20844 (N_20844,N_17838,N_19953);
and U20845 (N_20845,N_19485,N_16957);
nand U20846 (N_20846,N_17315,N_16196);
and U20847 (N_20847,N_19702,N_19488);
nor U20848 (N_20848,N_15474,N_17138);
xor U20849 (N_20849,N_17309,N_19376);
nor U20850 (N_20850,N_15572,N_18151);
xor U20851 (N_20851,N_19405,N_17295);
and U20852 (N_20852,N_15571,N_16997);
or U20853 (N_20853,N_16464,N_19233);
or U20854 (N_20854,N_16941,N_16827);
or U20855 (N_20855,N_16722,N_15939);
or U20856 (N_20856,N_19181,N_15102);
or U20857 (N_20857,N_17381,N_16164);
nand U20858 (N_20858,N_16025,N_18541);
xor U20859 (N_20859,N_16870,N_15256);
nand U20860 (N_20860,N_16985,N_17316);
xnor U20861 (N_20861,N_15067,N_19558);
nand U20862 (N_20862,N_16395,N_15908);
or U20863 (N_20863,N_18549,N_15929);
and U20864 (N_20864,N_15959,N_17693);
or U20865 (N_20865,N_17994,N_18838);
nand U20866 (N_20866,N_17385,N_15268);
xnor U20867 (N_20867,N_19594,N_17544);
xor U20868 (N_20868,N_18059,N_19326);
nand U20869 (N_20869,N_19351,N_15190);
nand U20870 (N_20870,N_16959,N_15477);
xnor U20871 (N_20871,N_19685,N_16495);
or U20872 (N_20872,N_15060,N_19723);
or U20873 (N_20873,N_19461,N_15300);
xor U20874 (N_20874,N_17268,N_16940);
nor U20875 (N_20875,N_16992,N_17242);
and U20876 (N_20876,N_19707,N_19462);
nand U20877 (N_20877,N_17884,N_17150);
nor U20878 (N_20878,N_16606,N_15542);
or U20879 (N_20879,N_16960,N_17499);
or U20880 (N_20880,N_16118,N_17500);
nand U20881 (N_20881,N_18907,N_17370);
nor U20882 (N_20882,N_19321,N_15483);
or U20883 (N_20883,N_15866,N_18813);
nand U20884 (N_20884,N_15376,N_18660);
xor U20885 (N_20885,N_19200,N_17974);
xor U20886 (N_20886,N_18116,N_16088);
nor U20887 (N_20887,N_16805,N_18149);
or U20888 (N_20888,N_15119,N_18774);
nor U20889 (N_20889,N_19674,N_18201);
nor U20890 (N_20890,N_18535,N_19079);
nand U20891 (N_20891,N_19868,N_16050);
or U20892 (N_20892,N_17485,N_16231);
nor U20893 (N_20893,N_18816,N_17220);
and U20894 (N_20894,N_19497,N_16862);
nor U20895 (N_20895,N_16452,N_19991);
xnor U20896 (N_20896,N_17794,N_18964);
nor U20897 (N_20897,N_17880,N_18627);
or U20898 (N_20898,N_16994,N_16546);
or U20899 (N_20899,N_16948,N_18773);
or U20900 (N_20900,N_19087,N_19839);
xnor U20901 (N_20901,N_18684,N_19315);
xnor U20902 (N_20902,N_15428,N_16707);
and U20903 (N_20903,N_15664,N_15072);
and U20904 (N_20904,N_19713,N_18257);
or U20905 (N_20905,N_15025,N_17995);
or U20906 (N_20906,N_17267,N_15568);
nor U20907 (N_20907,N_16720,N_17298);
and U20908 (N_20908,N_16884,N_18963);
and U20909 (N_20909,N_19385,N_18221);
and U20910 (N_20910,N_17759,N_18885);
xor U20911 (N_20911,N_19638,N_17965);
nor U20912 (N_20912,N_16245,N_15263);
nand U20913 (N_20913,N_16676,N_19632);
nand U20914 (N_20914,N_17836,N_18857);
nor U20915 (N_20915,N_15353,N_18382);
nand U20916 (N_20916,N_19193,N_15397);
or U20917 (N_20917,N_19958,N_15700);
nand U20918 (N_20918,N_19483,N_18837);
xor U20919 (N_20919,N_16666,N_16391);
nand U20920 (N_20920,N_17108,N_17487);
nand U20921 (N_20921,N_19543,N_16255);
or U20922 (N_20922,N_17840,N_18750);
nor U20923 (N_20923,N_16645,N_15607);
xor U20924 (N_20924,N_17417,N_18662);
nor U20925 (N_20925,N_19197,N_16377);
nor U20926 (N_20926,N_15752,N_19675);
and U20927 (N_20927,N_19513,N_19228);
xor U20928 (N_20928,N_15507,N_19247);
or U20929 (N_20929,N_17428,N_18787);
xor U20930 (N_20930,N_15935,N_19328);
or U20931 (N_20931,N_17554,N_17632);
or U20932 (N_20932,N_16796,N_16062);
nor U20933 (N_20933,N_15816,N_18607);
and U20934 (N_20934,N_15585,N_19869);
and U20935 (N_20935,N_19588,N_16217);
xnor U20936 (N_20936,N_19264,N_18302);
nor U20937 (N_20937,N_17231,N_17179);
nor U20938 (N_20938,N_18468,N_17099);
nand U20939 (N_20939,N_17513,N_19063);
and U20940 (N_20940,N_16612,N_17294);
nand U20941 (N_20941,N_19147,N_16509);
nor U20942 (N_20942,N_15470,N_19598);
or U20943 (N_20943,N_15130,N_19391);
xor U20944 (N_20944,N_19477,N_15484);
nand U20945 (N_20945,N_18593,N_18010);
nor U20946 (N_20946,N_16603,N_15061);
or U20947 (N_20947,N_19532,N_19548);
xnor U20948 (N_20948,N_15374,N_18494);
xnor U20949 (N_20949,N_15974,N_15622);
and U20950 (N_20950,N_15773,N_15361);
and U20951 (N_20951,N_17735,N_19170);
and U20952 (N_20952,N_19014,N_19451);
xnor U20953 (N_20953,N_18081,N_19919);
xor U20954 (N_20954,N_17273,N_18058);
and U20955 (N_20955,N_16266,N_15519);
nor U20956 (N_20956,N_18786,N_17465);
nor U20957 (N_20957,N_15207,N_16761);
nand U20958 (N_20958,N_19222,N_18312);
nor U20959 (N_20959,N_16757,N_17914);
and U20960 (N_20960,N_19795,N_19290);
or U20961 (N_20961,N_16091,N_15073);
nand U20962 (N_20962,N_19148,N_15204);
xnor U20963 (N_20963,N_16406,N_17469);
nand U20964 (N_20964,N_15670,N_18709);
nand U20965 (N_20965,N_17637,N_18590);
or U20966 (N_20966,N_18899,N_18954);
or U20967 (N_20967,N_18612,N_19051);
nor U20968 (N_20968,N_15809,N_19466);
nor U20969 (N_20969,N_17474,N_19016);
nand U20970 (N_20970,N_18680,N_19017);
nand U20971 (N_20971,N_19186,N_18177);
nand U20972 (N_20972,N_15966,N_15077);
or U20973 (N_20973,N_17216,N_16390);
and U20974 (N_20974,N_18103,N_19572);
nand U20975 (N_20975,N_19542,N_19846);
xor U20976 (N_20976,N_15713,N_18789);
nand U20977 (N_20977,N_18360,N_16533);
or U20978 (N_20978,N_17115,N_16589);
or U20979 (N_20979,N_16910,N_16592);
nor U20980 (N_20980,N_15538,N_17931);
and U20981 (N_20981,N_17903,N_19152);
or U20982 (N_20982,N_15231,N_16531);
nand U20983 (N_20983,N_16943,N_17205);
xnor U20984 (N_20984,N_16007,N_17458);
or U20985 (N_20985,N_16501,N_18623);
nand U20986 (N_20986,N_16066,N_16630);
and U20987 (N_20987,N_18311,N_15855);
xnor U20988 (N_20988,N_16795,N_16952);
or U20989 (N_20989,N_16996,N_16917);
and U20990 (N_20990,N_18589,N_15096);
and U20991 (N_20991,N_16931,N_17860);
and U20992 (N_20992,N_19920,N_16013);
nor U20993 (N_20993,N_16858,N_17400);
or U20994 (N_20994,N_15749,N_17951);
or U20995 (N_20995,N_18667,N_16211);
and U20996 (N_20996,N_15761,N_18035);
nor U20997 (N_20997,N_18165,N_18438);
xnor U20998 (N_20998,N_18503,N_18610);
xor U20999 (N_20999,N_17287,N_19226);
nor U21000 (N_21000,N_18772,N_16582);
and U21001 (N_21001,N_16919,N_15294);
xnor U21002 (N_21002,N_16655,N_15881);
nor U21003 (N_21003,N_19758,N_17110);
xnor U21004 (N_21004,N_19772,N_15805);
nand U21005 (N_21005,N_18620,N_18656);
xnor U21006 (N_21006,N_18714,N_15379);
nor U21007 (N_21007,N_16154,N_19145);
or U21008 (N_21008,N_19489,N_15794);
nand U21009 (N_21009,N_16559,N_16380);
nor U21010 (N_21010,N_15498,N_19380);
or U21011 (N_21011,N_19838,N_18880);
nor U21012 (N_21012,N_17804,N_19516);
nor U21013 (N_21013,N_16642,N_17517);
and U21014 (N_21014,N_16848,N_17881);
xnor U21015 (N_21015,N_17325,N_19891);
and U21016 (N_21016,N_16684,N_18150);
or U21017 (N_21017,N_15672,N_16175);
or U21018 (N_21018,N_17084,N_15401);
and U21019 (N_21019,N_19112,N_18423);
and U21020 (N_21020,N_15309,N_18584);
or U21021 (N_21021,N_16492,N_15099);
nor U21022 (N_21022,N_19325,N_19414);
or U21023 (N_21023,N_15114,N_15162);
and U21024 (N_21024,N_19925,N_18477);
nor U21025 (N_21025,N_17662,N_16878);
and U21026 (N_21026,N_17987,N_19970);
nand U21027 (N_21027,N_16473,N_15942);
nand U21028 (N_21028,N_16883,N_19865);
xnor U21029 (N_21029,N_16780,N_19409);
or U21030 (N_21030,N_18446,N_19901);
or U21031 (N_21031,N_17223,N_16794);
or U21032 (N_21032,N_18225,N_19336);
nand U21033 (N_21033,N_15450,N_17823);
nor U21034 (N_21034,N_19368,N_15386);
nand U21035 (N_21035,N_15704,N_18173);
or U21036 (N_21036,N_18977,N_16643);
or U21037 (N_21037,N_19930,N_15532);
xor U21038 (N_21038,N_15854,N_16932);
and U21039 (N_21039,N_16526,N_15776);
nor U21040 (N_21040,N_15286,N_16130);
xor U21041 (N_21041,N_17775,N_18245);
and U21042 (N_21042,N_15719,N_16550);
nand U21043 (N_21043,N_15517,N_18303);
nand U21044 (N_21044,N_17068,N_19484);
nor U21045 (N_21045,N_19780,N_16510);
xnor U21046 (N_21046,N_18834,N_15707);
nand U21047 (N_21047,N_15521,N_17537);
or U21048 (N_21048,N_15196,N_16953);
or U21049 (N_21049,N_19236,N_15329);
and U21050 (N_21050,N_18411,N_17895);
nor U21051 (N_21051,N_17460,N_17703);
xor U21052 (N_21052,N_16774,N_17750);
nor U21053 (N_21053,N_15088,N_17461);
and U21054 (N_21054,N_15238,N_19874);
and U21055 (N_21055,N_16084,N_17851);
and U21056 (N_21056,N_19253,N_19171);
or U21057 (N_21057,N_16986,N_19044);
or U21058 (N_21058,N_15387,N_19184);
and U21059 (N_21059,N_16331,N_16632);
or U21060 (N_21060,N_15241,N_17404);
and U21061 (N_21061,N_16581,N_15982);
or U21062 (N_21062,N_15422,N_19356);
or U21063 (N_21063,N_16503,N_16942);
and U21064 (N_21064,N_19153,N_19465);
xor U21065 (N_21065,N_19282,N_17869);
xnor U21066 (N_21066,N_18622,N_19630);
xor U21067 (N_21067,N_16279,N_19749);
or U21068 (N_21068,N_17125,N_18455);
and U21069 (N_21069,N_18370,N_19830);
xor U21070 (N_21070,N_18124,N_17802);
nor U21071 (N_21071,N_16727,N_19178);
or U21072 (N_21072,N_19163,N_17367);
nor U21073 (N_21073,N_17493,N_15325);
and U21074 (N_21074,N_19005,N_17288);
and U21075 (N_21075,N_19481,N_15777);
or U21076 (N_21076,N_18895,N_18646);
nand U21077 (N_21077,N_15446,N_19870);
nand U21078 (N_21078,N_16243,N_15737);
xor U21079 (N_21079,N_16937,N_18317);
nand U21080 (N_21080,N_18993,N_15772);
or U21081 (N_21081,N_17812,N_17959);
and U21082 (N_21082,N_16887,N_19407);
nor U21083 (N_21083,N_19624,N_15541);
or U21084 (N_21084,N_19776,N_19342);
nor U21085 (N_21085,N_17990,N_18005);
nor U21086 (N_21086,N_17188,N_16797);
nor U21087 (N_21087,N_17030,N_17560);
nor U21088 (N_21088,N_18520,N_15262);
nor U21089 (N_21089,N_18139,N_18979);
nor U21090 (N_21090,N_17322,N_18046);
xnor U21091 (N_21091,N_16626,N_19578);
nand U21092 (N_21092,N_16527,N_17800);
nand U21093 (N_21093,N_16202,N_18523);
nor U21094 (N_21094,N_17947,N_18519);
and U21095 (N_21095,N_19892,N_16854);
and U21096 (N_21096,N_18966,N_19602);
or U21097 (N_21097,N_15899,N_18197);
or U21098 (N_21098,N_19367,N_16252);
or U21099 (N_21099,N_18578,N_19977);
or U21100 (N_21100,N_15955,N_16361);
and U21101 (N_21101,N_15621,N_19024);
and U21102 (N_21102,N_19400,N_17558);
nor U21103 (N_21103,N_16515,N_19671);
xor U21104 (N_21104,N_19457,N_16470);
and U21105 (N_21105,N_19135,N_18844);
nor U21106 (N_21106,N_16205,N_18941);
and U21107 (N_21107,N_18159,N_18120);
or U21108 (N_21108,N_19347,N_17292);
nor U21109 (N_21109,N_18189,N_16210);
nand U21110 (N_21110,N_17894,N_17626);
nor U21111 (N_21111,N_18237,N_15927);
nand U21112 (N_21112,N_18697,N_17997);
xor U21113 (N_21113,N_15115,N_18573);
or U21114 (N_21114,N_18261,N_17159);
nand U21115 (N_21115,N_19647,N_19912);
nor U21116 (N_21116,N_16337,N_15662);
nand U21117 (N_21117,N_16147,N_17498);
nand U21118 (N_21118,N_18669,N_16664);
nor U21119 (N_21119,N_19809,N_16022);
nand U21120 (N_21120,N_16191,N_17217);
xnor U21121 (N_21121,N_19218,N_17450);
xor U21122 (N_21122,N_17497,N_17166);
nor U21123 (N_21123,N_19655,N_16089);
and U21124 (N_21124,N_18019,N_16826);
nand U21125 (N_21125,N_15192,N_16077);
and U21126 (N_21126,N_17534,N_19293);
nand U21127 (N_21127,N_15339,N_15612);
or U21128 (N_21128,N_18991,N_18872);
or U21129 (N_21129,N_16947,N_18809);
nand U21130 (N_21130,N_19069,N_19678);
nand U21131 (N_21131,N_19308,N_18534);
nor U21132 (N_21132,N_17341,N_15487);
nor U21133 (N_21133,N_19631,N_18290);
xnor U21134 (N_21134,N_17781,N_15107);
or U21135 (N_21135,N_19857,N_15632);
xnor U21136 (N_21136,N_19387,N_17808);
xnor U21137 (N_21137,N_16542,N_18744);
nor U21138 (N_21138,N_15026,N_18802);
or U21139 (N_21139,N_19790,N_19657);
nor U21140 (N_21140,N_16801,N_19036);
and U21141 (N_21141,N_18341,N_19622);
nand U21142 (N_21142,N_19650,N_17673);
nor U21143 (N_21143,N_16069,N_18846);
nor U21144 (N_21144,N_16494,N_16429);
and U21145 (N_21145,N_15838,N_18947);
xor U21146 (N_21146,N_19130,N_17312);
nor U21147 (N_21147,N_19986,N_19937);
xor U21148 (N_21148,N_18869,N_18793);
nor U21149 (N_21149,N_19770,N_15160);
or U21150 (N_21150,N_18020,N_19754);
nand U21151 (N_21151,N_18621,N_15661);
or U21152 (N_21152,N_19810,N_16719);
xor U21153 (N_21153,N_16277,N_16308);
nand U21154 (N_21154,N_19981,N_15159);
nand U21155 (N_21155,N_18790,N_19476);
nand U21156 (N_21156,N_16591,N_17696);
or U21157 (N_21157,N_18771,N_16635);
or U21158 (N_21158,N_15106,N_17418);
nand U21159 (N_21159,N_18125,N_15757);
or U21160 (N_21160,N_19026,N_18631);
or U21161 (N_21161,N_16846,N_17144);
xor U21162 (N_21162,N_16232,N_15205);
or U21163 (N_21163,N_19032,N_16833);
xor U21164 (N_21164,N_18836,N_19025);
and U21165 (N_21165,N_17631,N_19146);
nor U21166 (N_21166,N_18483,N_17248);
nand U21167 (N_21167,N_19345,N_15533);
nand U21168 (N_21168,N_19312,N_19560);
nor U21169 (N_21169,N_15531,N_19099);
or U21170 (N_21170,N_17519,N_17674);
nand U21171 (N_21171,N_18767,N_19792);
nand U21172 (N_21172,N_15403,N_17270);
xnor U21173 (N_21173,N_18630,N_17574);
or U21174 (N_21174,N_15835,N_15186);
xor U21175 (N_21175,N_18903,N_19842);
xnor U21176 (N_21176,N_18884,N_17070);
and U21177 (N_21177,N_15441,N_18465);
or U21178 (N_21178,N_18756,N_15074);
nor U21179 (N_21179,N_16325,N_17429);
and U21180 (N_21180,N_17098,N_17053);
nand U21181 (N_21181,N_16324,N_18332);
xor U21182 (N_21182,N_19684,N_17719);
or U21183 (N_21183,N_15997,N_18487);
or U21184 (N_21184,N_15076,N_16586);
nand U21185 (N_21185,N_15180,N_16657);
xnor U21186 (N_21186,N_18655,N_16220);
xnor U21187 (N_21187,N_19510,N_15836);
nor U21188 (N_21188,N_16772,N_18778);
nand U21189 (N_21189,N_17940,N_16834);
or U21190 (N_21190,N_19823,N_19341);
or U21191 (N_21191,N_15798,N_19374);
nand U21192 (N_21192,N_15455,N_19160);
nor U21193 (N_21193,N_15972,N_15863);
nand U21194 (N_21194,N_18945,N_19065);
xor U21195 (N_21195,N_19127,N_19332);
and U21196 (N_21196,N_15780,N_17768);
or U21197 (N_21197,N_16128,N_15016);
nand U21198 (N_21198,N_15602,N_18745);
or U21199 (N_21199,N_17136,N_19762);
and U21200 (N_21200,N_19437,N_19279);
nand U21201 (N_21201,N_18741,N_17376);
nor U21202 (N_21202,N_15808,N_18830);
nor U21203 (N_21203,N_15037,N_17219);
or U21204 (N_21204,N_18306,N_19055);
nor U21205 (N_21205,N_15511,N_19911);
nor U21206 (N_21206,N_17230,N_17949);
and U21207 (N_21207,N_17394,N_15904);
xnor U21208 (N_21208,N_17773,N_18008);
and U21209 (N_21209,N_17595,N_15356);
nand U21210 (N_21210,N_18090,N_19645);
nor U21211 (N_21211,N_17031,N_16989);
xnor U21212 (N_21212,N_19691,N_19251);
or U21213 (N_21213,N_16971,N_16280);
nand U21214 (N_21214,N_16113,N_18308);
nor U21215 (N_21215,N_18606,N_17629);
and U21216 (N_21216,N_16016,N_19265);
nand U21217 (N_21217,N_17406,N_15246);
and U21218 (N_21218,N_18876,N_17826);
nor U21219 (N_21219,N_19319,N_17922);
nand U21220 (N_21220,N_19725,N_15452);
nor U21221 (N_21221,N_16621,N_19703);
and U21222 (N_21222,N_15868,N_19524);
and U21223 (N_21223,N_19411,N_16871);
and U21224 (N_21224,N_15522,N_18365);
xor U21225 (N_21225,N_18038,N_18832);
or U21226 (N_21226,N_19246,N_17536);
and U21227 (N_21227,N_15245,N_15284);
and U21228 (N_21228,N_15723,N_15405);
and U21229 (N_21229,N_18924,N_18191);
or U21230 (N_21230,N_15156,N_17636);
and U21231 (N_21231,N_19765,N_17962);
nand U21232 (N_21232,N_16448,N_17036);
and U21233 (N_21233,N_16214,N_17439);
or U21234 (N_21234,N_18013,N_18094);
nand U21235 (N_21235,N_15703,N_15640);
xor U21236 (N_21236,N_15964,N_15494);
nor U21237 (N_21237,N_15283,N_16549);
xor U21238 (N_21238,N_16286,N_18000);
or U21239 (N_21239,N_16865,N_19593);
nand U21240 (N_21240,N_17505,N_18681);
nand U21241 (N_21241,N_16576,N_17342);
nor U21242 (N_21242,N_17228,N_17104);
nand U21243 (N_21243,N_19648,N_17105);
nor U21244 (N_21244,N_17272,N_16020);
nor U21245 (N_21245,N_18842,N_18379);
xnor U21246 (N_21246,N_15608,N_15140);
nor U21247 (N_21247,N_18553,N_17956);
nor U21248 (N_21248,N_15791,N_17793);
nand U21249 (N_21249,N_16668,N_18368);
or U21250 (N_21250,N_15335,N_16172);
nor U21251 (N_21251,N_17898,N_18252);
nand U21252 (N_21252,N_17085,N_19552);
or U21253 (N_21253,N_17011,N_17809);
nand U21254 (N_21254,N_16019,N_16938);
nand U21255 (N_21255,N_15234,N_17464);
nand U21256 (N_21256,N_17846,N_16701);
nand U21257 (N_21257,N_15279,N_15293);
or U21258 (N_21258,N_18563,N_19298);
and U21259 (N_21259,N_19083,N_19142);
xnor U21260 (N_21260,N_19803,N_18448);
nor U21261 (N_21261,N_18645,N_17579);
and U21262 (N_21262,N_19729,N_15864);
nand U21263 (N_21263,N_15576,N_19201);
nor U21264 (N_21264,N_18473,N_17441);
nand U21265 (N_21265,N_19444,N_18710);
xor U21266 (N_21266,N_17883,N_16890);
and U21267 (N_21267,N_15983,N_17623);
and U21268 (N_21268,N_15141,N_18394);
nand U21269 (N_21269,N_16641,N_17576);
or U21270 (N_21270,N_19811,N_19008);
nor U21271 (N_21271,N_15420,N_16552);
nand U21272 (N_21272,N_16117,N_17199);
nand U21273 (N_21273,N_18251,N_18163);
nor U21274 (N_21274,N_15756,N_15561);
nand U21275 (N_21275,N_16691,N_15883);
nand U21276 (N_21276,N_18024,N_15988);
and U21277 (N_21277,N_18812,N_15275);
and U21278 (N_21278,N_15953,N_17671);
xor U21279 (N_21279,N_15385,N_17058);
nand U21280 (N_21280,N_18999,N_19775);
and U21281 (N_21281,N_17280,N_17421);
or U21282 (N_21282,N_17158,N_18650);
nor U21283 (N_21283,N_17657,N_18062);
xnor U21284 (N_21284,N_16379,N_17655);
and U21285 (N_21285,N_17744,N_17194);
xor U21286 (N_21286,N_16194,N_16860);
nor U21287 (N_21287,N_17556,N_19473);
or U21288 (N_21288,N_15280,N_15473);
nand U21289 (N_21289,N_15648,N_17346);
xnor U21290 (N_21290,N_16573,N_15829);
xnor U21291 (N_21291,N_15327,N_19132);
nand U21292 (N_21292,N_16975,N_18209);
and U21293 (N_21293,N_17716,N_19434);
or U21294 (N_21294,N_15481,N_18304);
nor U21295 (N_21295,N_18683,N_19957);
nand U21296 (N_21296,N_19735,N_15918);
xor U21297 (N_21297,N_17240,N_19750);
nand U21298 (N_21298,N_18141,N_15163);
nand U21299 (N_21299,N_15875,N_15501);
and U21300 (N_21300,N_16006,N_15230);
and U21301 (N_21301,N_19060,N_17559);
nand U21302 (N_21302,N_17208,N_15692);
and U21303 (N_21303,N_17741,N_17328);
or U21304 (N_21304,N_15399,N_19114);
nand U21305 (N_21305,N_16912,N_15615);
or U21306 (N_21306,N_15200,N_16990);
and U21307 (N_21307,N_17543,N_18536);
or U21308 (N_21308,N_15592,N_19623);
xnor U21309 (N_21309,N_17190,N_16697);
xor U21310 (N_21310,N_16545,N_18348);
or U21311 (N_21311,N_17726,N_18236);
and U21312 (N_21312,N_16460,N_16699);
nand U21313 (N_21313,N_17527,N_19435);
nor U21314 (N_21314,N_19760,N_19232);
or U21315 (N_21315,N_16680,N_18339);
xor U21316 (N_21316,N_16284,N_16808);
nor U21317 (N_21317,N_15255,N_18839);
nor U21318 (N_21318,N_16440,N_16998);
or U21319 (N_21319,N_18415,N_17850);
xnor U21320 (N_21320,N_16737,N_16082);
nand U21321 (N_21321,N_18156,N_17438);
xnor U21322 (N_21322,N_18073,N_16793);
xnor U21323 (N_21323,N_18288,N_16264);
nor U21324 (N_21324,N_15212,N_17304);
or U21325 (N_21325,N_15800,N_19501);
or U21326 (N_21326,N_15676,N_19777);
or U21327 (N_21327,N_16517,N_17227);
or U21328 (N_21328,N_17192,N_18178);
xnor U21329 (N_21329,N_19814,N_16033);
xor U21330 (N_21330,N_16272,N_18217);
xor U21331 (N_21331,N_18219,N_19089);
nor U21332 (N_21332,N_16259,N_16042);
nor U21333 (N_21333,N_16685,N_16644);
and U21334 (N_21334,N_16002,N_17639);
nand U21335 (N_21335,N_18095,N_15183);
or U21336 (N_21336,N_16956,N_16704);
nand U21337 (N_21337,N_19281,N_17483);
and U21338 (N_21338,N_17390,N_18920);
or U21339 (N_21339,N_18860,N_18180);
xnor U21340 (N_21340,N_17196,N_19964);
nand U21341 (N_21341,N_18275,N_18347);
and U21342 (N_21342,N_18053,N_17817);
nor U21343 (N_21343,N_19806,N_16879);
xnor U21344 (N_21344,N_16049,N_17740);
nor U21345 (N_21345,N_16318,N_17314);
and U21346 (N_21346,N_17434,N_17135);
and U21347 (N_21347,N_18025,N_16453);
xor U21348 (N_21348,N_16623,N_17916);
nand U21349 (N_21349,N_16300,N_17097);
and U21350 (N_21350,N_19237,N_18897);
or U21351 (N_21351,N_16776,N_16524);
nor U21352 (N_21352,N_18753,N_15153);
xor U21353 (N_21353,N_19469,N_19003);
or U21354 (N_21354,N_15459,N_18204);
xor U21355 (N_21355,N_16339,N_19204);
and U21356 (N_21356,N_16624,N_17323);
nor U21357 (N_21357,N_16970,N_18097);
and U21358 (N_21358,N_19357,N_15221);
nor U21359 (N_21359,N_16183,N_17472);
nand U21360 (N_21360,N_18061,N_19586);
nor U21361 (N_21361,N_18472,N_17289);
nor U21362 (N_21362,N_15547,N_15179);
or U21363 (N_21363,N_18529,N_19971);
or U21364 (N_21364,N_17622,N_19019);
and U21365 (N_21365,N_15611,N_16353);
xnor U21366 (N_21366,N_15598,N_17889);
xnor U21367 (N_21367,N_16471,N_17913);
xor U21368 (N_21368,N_17286,N_17609);
or U21369 (N_21369,N_19789,N_19242);
nand U21370 (N_21370,N_19495,N_18119);
nand U21371 (N_21371,N_15113,N_19798);
nor U21372 (N_21372,N_17299,N_18998);
xnor U21373 (N_21373,N_15150,N_19108);
nand U21374 (N_21374,N_19540,N_18777);
xnor U21375 (N_21375,N_19463,N_18571);
xnor U21376 (N_21376,N_16287,N_17855);
xnor U21377 (N_21377,N_18202,N_16426);
and U21378 (N_21378,N_18722,N_17751);
xor U21379 (N_21379,N_18985,N_16596);
and U21380 (N_21380,N_17392,N_16747);
and U21381 (N_21381,N_16872,N_19943);
nor U21382 (N_21382,N_16880,N_18863);
nor U21383 (N_21383,N_19835,N_19216);
and U21384 (N_21384,N_19490,N_16634);
or U21385 (N_21385,N_15583,N_17827);
or U21386 (N_21386,N_15454,N_17736);
or U21387 (N_21387,N_17243,N_18975);
xor U21388 (N_21388,N_19774,N_16715);
nor U21389 (N_21389,N_15358,N_18976);
nor U21390 (N_21390,N_15402,N_17143);
or U21391 (N_21391,N_15869,N_19375);
or U21392 (N_21392,N_16345,N_15078);
or U21393 (N_21393,N_15349,N_16628);
or U21394 (N_21394,N_19182,N_18002);
or U21395 (N_21395,N_15803,N_19545);
or U21396 (N_21396,N_18367,N_19263);
xnor U21397 (N_21397,N_19267,N_18935);
and U21398 (N_21398,N_15891,N_16063);
or U21399 (N_21399,N_17232,N_17589);
nor U21400 (N_21400,N_19353,N_18283);
nor U21401 (N_21401,N_16771,N_19646);
xor U21402 (N_21402,N_17206,N_18815);
xnor U21403 (N_21403,N_16500,N_15890);
or U21404 (N_21404,N_16417,N_15338);
nor U21405 (N_21405,N_17419,N_16972);
nand U21406 (N_21406,N_19102,N_16061);
or U21407 (N_21407,N_18866,N_19257);
nor U21408 (N_21408,N_15363,N_15394);
nand U21409 (N_21409,N_17774,N_16922);
nor U21410 (N_21410,N_16451,N_17814);
nand U21411 (N_21411,N_18431,N_19224);
and U21412 (N_21412,N_19354,N_17241);
nand U21413 (N_21413,N_19878,N_18971);
xnor U21414 (N_21414,N_15877,N_15466);
and U21415 (N_21415,N_16112,N_15924);
or U21416 (N_21416,N_15649,N_19948);
and U21417 (N_21417,N_15493,N_19972);
and U21418 (N_21418,N_16010,N_19995);
and U21419 (N_21419,N_15673,N_17896);
nor U21420 (N_21420,N_18129,N_16822);
or U21421 (N_21421,N_17948,N_15111);
and U21422 (N_21422,N_15337,N_18108);
nand U21423 (N_21423,N_16894,N_19924);
xor U21424 (N_21424,N_19234,N_19683);
xor U21425 (N_21425,N_18783,N_16385);
nand U21426 (N_21426,N_17034,N_19022);
nor U21427 (N_21427,N_18196,N_15663);
and U21428 (N_21428,N_19440,N_16055);
xnor U21429 (N_21429,N_19511,N_15369);
or U21430 (N_21430,N_15485,N_16868);
or U21431 (N_21431,N_17014,N_19377);
nand U21432 (N_21432,N_17945,N_17943);
and U21433 (N_21433,N_15259,N_18208);
nand U21434 (N_21434,N_19664,N_16908);
nand U21435 (N_21435,N_19841,N_16877);
xnor U21436 (N_21436,N_19787,N_15144);
nor U21437 (N_21437,N_19012,N_16093);
or U21438 (N_21438,N_15931,N_19121);
or U21439 (N_21439,N_15906,N_18392);
nand U21440 (N_21440,N_15299,N_17486);
nand U21441 (N_21441,N_18166,N_18754);
or U21442 (N_21442,N_15977,N_19467);
and U21443 (N_21443,N_17926,N_15166);
nand U21444 (N_21444,N_16813,N_19998);
nand U21445 (N_21445,N_18437,N_18464);
and U21446 (N_21446,N_18841,N_15551);
nand U21447 (N_21447,N_17021,N_18634);
nor U21448 (N_21448,N_17265,N_17646);
nor U21449 (N_21449,N_15807,N_15226);
nand U21450 (N_21450,N_18113,N_18132);
and U21451 (N_21451,N_19412,N_18495);
xor U21452 (N_21452,N_18413,N_15092);
nand U21453 (N_21453,N_18594,N_15264);
nand U21454 (N_21454,N_15003,N_18708);
or U21455 (N_21455,N_17379,N_18533);
nand U21456 (N_21456,N_17580,N_16945);
nor U21457 (N_21457,N_19188,N_17918);
nand U21458 (N_21458,N_17175,N_19612);
nor U21459 (N_21459,N_18155,N_16001);
xor U21460 (N_21460,N_17978,N_15384);
nor U21461 (N_21461,N_17440,N_17183);
nand U21462 (N_21462,N_19390,N_19922);
or U21463 (N_21463,N_16618,N_17371);
and U21464 (N_21464,N_19753,N_18587);
or U21465 (N_21465,N_17805,N_18470);
nand U21466 (N_21466,N_16888,N_18927);
nand U21467 (N_21467,N_19701,N_15495);
nor U21468 (N_21468,N_15741,N_18565);
or U21469 (N_21469,N_16768,N_18264);
nand U21470 (N_21470,N_16609,N_15254);
and U21471 (N_21471,N_19766,N_17330);
xnor U21472 (N_21472,N_17711,N_18821);
xnor U21473 (N_21473,N_19139,N_16698);
xnor U21474 (N_21474,N_16098,N_16238);
or U21475 (N_21475,N_17571,N_16968);
and U21476 (N_21476,N_17587,N_18826);
xnor U21477 (N_21477,N_17925,N_15155);
or U21478 (N_21478,N_15759,N_19230);
nor U21479 (N_21479,N_19928,N_15272);
xor U21480 (N_21480,N_17229,N_19155);
nand U21481 (N_21481,N_16487,N_16964);
or U21482 (N_21482,N_15098,N_18356);
and U21483 (N_21483,N_15208,N_17087);
and U21484 (N_21484,N_19613,N_17358);
nor U21485 (N_21485,N_17090,N_18136);
and U21486 (N_21486,N_19537,N_15007);
and U21487 (N_21487,N_17630,N_18779);
nor U21488 (N_21488,N_15315,N_19781);
xor U21489 (N_21489,N_15770,N_16965);
or U21490 (N_21490,N_16973,N_16096);
nand U21491 (N_21491,N_17972,N_15840);
or U21492 (N_21492,N_16654,N_17564);
and U21493 (N_21493,N_18344,N_18357);
nand U21494 (N_21494,N_18791,N_18517);
xor U21495 (N_21495,N_18182,N_16474);
and U21496 (N_21496,N_19480,N_17141);
and U21497 (N_21497,N_17577,N_18301);
xnor U21498 (N_21498,N_18870,N_16439);
nor U21499 (N_21499,N_17780,N_18788);
or U21500 (N_21500,N_16759,N_19123);
nor U21501 (N_21501,N_19335,N_19945);
nand U21502 (N_21502,N_19452,N_18820);
nand U21503 (N_21503,N_17495,N_16472);
xnor U21504 (N_21504,N_19286,N_17955);
nand U21505 (N_21505,N_15684,N_15083);
nand U21506 (N_21506,N_18504,N_18458);
and U21507 (N_21507,N_16254,N_16333);
xnor U21508 (N_21508,N_16407,N_18490);
and U21509 (N_21509,N_15396,N_15540);
xor U21510 (N_21510,N_15728,N_19877);
nor U21511 (N_21511,N_18805,N_17964);
and U21512 (N_21512,N_19164,N_18310);
nor U21513 (N_21513,N_19448,N_19906);
nor U21514 (N_21514,N_15370,N_17494);
xor U21515 (N_21515,N_16765,N_18154);
xor U21516 (N_21516,N_17327,N_16289);
or U21517 (N_21517,N_19105,N_16047);
or U21518 (N_21518,N_15440,N_19221);
nand U21519 (N_21519,N_15381,N_17897);
or U21520 (N_21520,N_15382,N_17333);
or U21521 (N_21521,N_19166,N_18759);
nand U21522 (N_21522,N_17357,N_16551);
xnor U21523 (N_21523,N_19927,N_15064);
nand U21524 (N_21524,N_15862,N_17207);
xor U21525 (N_21525,N_19030,N_18909);
or U21526 (N_21526,N_18613,N_17054);
or U21527 (N_21527,N_19273,N_19871);
or U21528 (N_21528,N_19317,N_16438);
xnor U21529 (N_21529,N_18374,N_19968);
or U21530 (N_21530,N_16537,N_19522);
nor U21531 (N_21531,N_18419,N_15799);
nor U21532 (N_21532,N_19956,N_18126);
nand U21533 (N_21533,N_16788,N_18291);
nor U21534 (N_21534,N_16144,N_16900);
or U21535 (N_21535,N_17518,N_15650);
or U21536 (N_21536,N_19746,N_16298);
nor U21537 (N_21537,N_16393,N_17479);
nand U21538 (N_21538,N_16223,N_17734);
nand U21539 (N_21539,N_19446,N_16135);
and U21540 (N_21540,N_17433,N_16305);
nor U21541 (N_21541,N_17009,N_15063);
or U21542 (N_21542,N_19670,N_18373);
nor U21543 (N_21543,N_18017,N_15326);
nor U21544 (N_21544,N_19020,N_15202);
nor U21545 (N_21545,N_16766,N_16151);
nand U21546 (N_21546,N_16555,N_15967);
nor U21547 (N_21547,N_17355,N_18570);
xor U21548 (N_21548,N_19211,N_17715);
or U21549 (N_21549,N_16607,N_15528);
nand U21550 (N_21550,N_17369,N_19897);
or U21551 (N_21551,N_16054,N_17530);
nand U21552 (N_21552,N_17910,N_15486);
nor U21553 (N_21553,N_15871,N_16065);
xor U21554 (N_21554,N_15870,N_17039);
nor U21555 (N_21555,N_19733,N_16506);
or U21556 (N_21556,N_15947,N_16411);
nor U21557 (N_21557,N_19944,N_16857);
and U21558 (N_21558,N_17202,N_19828);
nor U21559 (N_21559,N_19094,N_18579);
or U21560 (N_21560,N_18512,N_19333);
nand U21561 (N_21561,N_16770,N_18331);
and U21562 (N_21562,N_19763,N_17698);
and U21563 (N_21563,N_19379,N_17610);
and U21564 (N_21564,N_19979,N_19827);
and U21565 (N_21565,N_16859,N_15698);
xnor U21566 (N_21566,N_17377,N_16215);
and U21567 (N_21567,N_15328,N_18961);
or U21568 (N_21568,N_19072,N_18323);
nand U21569 (N_21569,N_18707,N_15367);
and U21570 (N_21570,N_15408,N_18576);
xor U21571 (N_21571,N_17492,N_19209);
nor U21572 (N_21572,N_15950,N_16523);
nand U21573 (N_21573,N_17642,N_15492);
or U21574 (N_21574,N_19276,N_16724);
or U21575 (N_21575,N_16387,N_15084);
xnor U21576 (N_21576,N_17786,N_17019);
or U21577 (N_21577,N_16738,N_17591);
nand U21578 (N_21578,N_17902,N_17048);
or U21579 (N_21579,N_16225,N_19001);
xor U21580 (N_21580,N_18951,N_19840);
xor U21581 (N_21581,N_19539,N_19705);
and U21582 (N_21582,N_17380,N_15270);
xor U21583 (N_21583,N_18905,N_18353);
nor U21584 (N_21584,N_17010,N_19667);
or U21585 (N_21585,N_17362,N_19887);
nand U21586 (N_21586,N_16686,N_15793);
and U21587 (N_21587,N_19609,N_17982);
xor U21588 (N_21588,N_17165,N_15675);
nor U21589 (N_21589,N_16106,N_17137);
nand U21590 (N_21590,N_18766,N_17893);
nor U21591 (N_21591,N_19156,N_16734);
nand U21592 (N_21592,N_19915,N_17770);
nor U21593 (N_21593,N_16383,N_17788);
nand U21594 (N_21594,N_17754,N_19738);
nand U21595 (N_21595,N_15747,N_17942);
nor U21596 (N_21596,N_19378,N_18387);
nor U21597 (N_21597,N_18449,N_15295);
or U21598 (N_21598,N_19092,N_18325);
xnor U21599 (N_21599,N_18693,N_19822);
nand U21600 (N_21600,N_15993,N_15831);
or U21601 (N_21601,N_19910,N_16017);
xnor U21602 (N_21602,N_16614,N_16433);
or U21603 (N_21603,N_18948,N_15489);
and U21604 (N_21604,N_17107,N_16178);
and U21605 (N_21605,N_16208,N_19062);
xor U21606 (N_21606,N_16100,N_18983);
xnor U21607 (N_21607,N_15623,N_15319);
or U21608 (N_21608,N_19637,N_17321);
nor U21609 (N_21609,N_16309,N_17742);
nand U21610 (N_21610,N_16835,N_15257);
xnor U21611 (N_21611,N_16659,N_18066);
xor U21612 (N_21612,N_15584,N_17708);
or U21613 (N_21613,N_18282,N_18160);
or U21614 (N_21614,N_17359,N_16798);
and U21615 (N_21615,N_19716,N_17862);
or U21616 (N_21616,N_18917,N_18740);
and U21617 (N_21617,N_17398,N_16484);
xnor U21618 (N_21618,N_18234,N_17638);
or U21619 (N_21619,N_19649,N_19547);
nand U21620 (N_21620,N_19607,N_15897);
xor U21621 (N_21621,N_17996,N_17944);
and U21622 (N_21622,N_15775,N_17688);
and U21623 (N_21623,N_17824,N_19346);
and U21624 (N_21624,N_16830,N_17811);
nand U21625 (N_21625,N_18934,N_18546);
nor U21626 (N_21626,N_17012,N_18045);
nand U21627 (N_21627,N_15901,N_15817);
nor U21628 (N_21628,N_17953,N_15178);
nand U21629 (N_21629,N_16627,N_16228);
nand U21630 (N_21630,N_16445,N_19824);
or U21631 (N_21631,N_15035,N_16060);
and U21632 (N_21632,N_15194,N_15999);
or U21633 (N_21633,N_17177,N_17906);
or U21634 (N_21634,N_16319,N_17484);
and U21635 (N_21635,N_15589,N_18679);
or U21636 (N_21636,N_17665,N_15266);
xnor U21637 (N_21637,N_17176,N_18887);
nand U21638 (N_21638,N_15120,N_16384);
nor U21639 (N_21639,N_15031,N_18893);
xor U21640 (N_21640,N_16414,N_19807);
nor U21641 (N_21641,N_19529,N_18506);
and U21642 (N_21642,N_18314,N_15687);
and U21643 (N_21643,N_17912,N_18241);
xor U21644 (N_21644,N_19687,N_19442);
or U21645 (N_21645,N_19402,N_15444);
or U21646 (N_21646,N_15605,N_15691);
nand U21647 (N_21647,N_15731,N_15907);
or U21648 (N_21648,N_17447,N_17641);
xor U21649 (N_21649,N_19561,N_15136);
xor U21650 (N_21650,N_19424,N_18475);
and U21651 (N_21651,N_16021,N_18337);
xor U21652 (N_21652,N_19225,N_17384);
nand U21653 (N_21653,N_16683,N_15758);
nor U21654 (N_21654,N_18591,N_15702);
or U21655 (N_21655,N_19043,N_15451);
nor U21656 (N_21656,N_17310,N_17184);
and U21657 (N_21657,N_17712,N_18092);
or U21658 (N_21658,N_16584,N_15229);
and U21659 (N_21659,N_18329,N_18391);
nor U21660 (N_21660,N_16730,N_18319);
nor U21661 (N_21661,N_18509,N_18380);
or U21662 (N_21662,N_15081,N_18277);
and U21663 (N_21663,N_16257,N_16954);
nor U21664 (N_21664,N_18919,N_16811);
nor U21665 (N_21665,N_18582,N_18063);
or U21666 (N_21666,N_15682,N_15624);
xnor U21667 (N_21667,N_15818,N_18334);
and U21668 (N_21668,N_16403,N_17088);
nand U21669 (N_21669,N_18122,N_19898);
nor U21670 (N_21670,N_16136,N_19300);
xor U21671 (N_21671,N_17391,N_19438);
and U21672 (N_21672,N_19002,N_15210);
and U21673 (N_21673,N_16892,N_19306);
xor U21674 (N_21674,N_16346,N_16512);
nand U21675 (N_21675,N_17714,N_17503);
and U21676 (N_21676,N_17721,N_15044);
or U21677 (N_21677,N_16480,N_15680);
nand U21678 (N_21678,N_17867,N_17067);
nand U21679 (N_21679,N_17981,N_17635);
and U21680 (N_21680,N_15961,N_17350);
and U21681 (N_21681,N_17617,N_18021);
and U21682 (N_21682,N_15526,N_16661);
xnor U21683 (N_21683,N_18908,N_15129);
and U21684 (N_21684,N_16392,N_19990);
or U21685 (N_21685,N_15355,N_15354);
nor U21686 (N_21686,N_17018,N_16681);
or U21687 (N_21687,N_15512,N_18164);
or U21688 (N_21688,N_18552,N_16818);
xor U21689 (N_21689,N_18939,N_19819);
or U21690 (N_21690,N_16036,N_19538);
xor U21691 (N_21691,N_15856,N_17000);
and U21692 (N_21692,N_17056,N_16441);
nor U21693 (N_21693,N_18210,N_15261);
and U21694 (N_21694,N_16005,N_18276);
nand U21695 (N_21695,N_15628,N_15554);
xnor U21696 (N_21696,N_15109,N_17106);
nor U21697 (N_21697,N_18583,N_15783);
nand U21698 (N_21698,N_16640,N_19048);
or U21699 (N_21699,N_15740,N_19686);
and U21700 (N_21700,N_18638,N_15919);
nand U21701 (N_21701,N_17704,N_15351);
or U21702 (N_21702,N_19389,N_18214);
or U21703 (N_21703,N_19799,N_17900);
xor U21704 (N_21704,N_18421,N_16201);
nor U21705 (N_21705,N_15824,N_18279);
or U21706 (N_21706,N_19658,N_16881);
or U21707 (N_21707,N_15784,N_15951);
xnor U21708 (N_21708,N_18274,N_18524);
nand U21709 (N_21709,N_15787,N_19690);
or U21710 (N_21710,N_18569,N_19330);
nor U21711 (N_21711,N_18521,N_17121);
nand U21712 (N_21712,N_17967,N_16507);
and U21713 (N_21713,N_19327,N_15206);
and U21714 (N_21714,N_16732,N_15320);
xnor U21715 (N_21715,N_19504,N_19416);
and U21716 (N_21716,N_16855,N_18652);
or U21717 (N_21717,N_15011,N_18496);
nand U21718 (N_21718,N_15665,N_16268);
xor U21719 (N_21719,N_18868,N_18188);
nor U21720 (N_21720,N_17843,N_19740);
or U21721 (N_21721,N_15278,N_15812);
or U21722 (N_21722,N_17724,N_19386);
and U21723 (N_21723,N_19165,N_16544);
nor U21724 (N_21724,N_17045,N_16605);
and U21725 (N_21725,N_16893,N_16660);
xnor U21726 (N_21726,N_15236,N_18758);
or U21727 (N_21727,N_18032,N_19199);
xnor U21728 (N_21728,N_16708,N_18727);
nand U21729 (N_21729,N_18729,N_19628);
or U21730 (N_21730,N_18824,N_15215);
nor U21731 (N_21731,N_16250,N_16777);
and U21732 (N_21732,N_17907,N_18343);
and U21733 (N_21733,N_15616,N_16508);
nand U21734 (N_21734,N_16293,N_18811);
xor U21735 (N_21735,N_16099,N_18400);
or U21736 (N_21736,N_15027,N_17347);
xnor U21737 (N_21737,N_16966,N_17815);
xnor U21738 (N_21738,N_17234,N_15022);
nand U21739 (N_21739,N_16949,N_17334);
nor U21740 (N_21740,N_16505,N_17111);
xnor U21741 (N_21741,N_17682,N_15896);
and U21742 (N_21742,N_15529,N_15005);
or U21743 (N_21743,N_16352,N_19520);
xor U21744 (N_21744,N_15733,N_17728);
nand U21745 (N_21745,N_19311,N_15391);
xnor U21746 (N_21746,N_17035,N_15743);
nor U21747 (N_21747,N_17628,N_15227);
and U21748 (N_21748,N_15438,N_19373);
or U21749 (N_21749,N_17660,N_18079);
and U21750 (N_21750,N_19633,N_18352);
and U21751 (N_21751,N_15641,N_16712);
xor U21752 (N_21752,N_18682,N_19569);
and U21753 (N_21753,N_19035,N_17806);
xnor U21754 (N_21754,N_17692,N_17382);
and U21755 (N_21755,N_16665,N_18601);
nor U21756 (N_21756,N_17663,N_17250);
or U21757 (N_21757,N_16764,N_19587);
or U21758 (N_21758,N_17423,N_17614);
xor U21759 (N_21759,N_19872,N_15994);
xor U21760 (N_21760,N_18765,N_18925);
or U21761 (N_21761,N_19383,N_18273);
or U21762 (N_21762,N_15768,N_18647);
xnor U21763 (N_21763,N_18932,N_15936);
xnor U21764 (N_21764,N_18730,N_16465);
nand U21765 (N_21765,N_16637,N_18022);
nand U21766 (N_21766,N_19873,N_19768);
xnor U21767 (N_21767,N_16622,N_17984);
nor U21768 (N_21768,N_19118,N_19747);
xor U21769 (N_21769,N_19304,N_15134);
xor U21770 (N_21770,N_18138,N_18725);
or U21771 (N_21771,N_19722,N_16459);
and U21772 (N_21772,N_16291,N_19861);
nand U21773 (N_21773,N_16690,N_17324);
nand U21774 (N_21774,N_16961,N_18441);
nand U21775 (N_21775,N_18206,N_19203);
nor U21776 (N_21776,N_17731,N_16702);
nand U21777 (N_21777,N_15832,N_18775);
nand U21778 (N_21778,N_18300,N_19616);
nand U21779 (N_21779,N_18364,N_18479);
xnor U21780 (N_21780,N_17134,N_19487);
nand U21781 (N_21781,N_17919,N_16869);
or U21782 (N_21782,N_19439,N_18109);
nor U21783 (N_21783,N_17023,N_19103);
nand U21784 (N_21784,N_18230,N_16253);
nand U21785 (N_21785,N_17986,N_15105);
nor U21786 (N_21786,N_17149,N_17032);
or U21787 (N_21787,N_18229,N_17504);
and U21788 (N_21788,N_15963,N_18218);
nand U21789 (N_21789,N_18049,N_18060);
xor U21790 (N_21790,N_16967,N_17857);
and U21791 (N_21791,N_15068,N_18395);
or U21792 (N_21792,N_16408,N_15804);
or U21793 (N_21793,N_18023,N_18657);
and U21794 (N_21794,N_15788,N_19363);
nand U21795 (N_21795,N_19426,N_16587);
xor U21796 (N_21796,N_19143,N_18422);
xnor U21797 (N_21797,N_17828,N_16275);
and U21798 (N_21798,N_16251,N_18207);
and U21799 (N_21799,N_15168,N_19252);
or U21800 (N_21800,N_19136,N_15668);
nand U21801 (N_21801,N_16120,N_15301);
and U21802 (N_21802,N_16044,N_18205);
xor U21803 (N_21803,N_15536,N_17930);
nand U21804 (N_21804,N_18677,N_19343);
xnor U21805 (N_21805,N_18619,N_15789);
xor U21806 (N_21806,N_15169,N_16886);
or U21807 (N_21807,N_16087,N_15674);
or U21808 (N_21808,N_19410,N_18363);
xor U21809 (N_21809,N_16636,N_16248);
xnor U21810 (N_21810,N_19791,N_17042);
xor U21811 (N_21811,N_19788,N_16143);
xor U21812 (N_21812,N_18599,N_19833);
or U21813 (N_21813,N_19961,N_19113);
or U21814 (N_21814,N_19190,N_17024);
and U21815 (N_21815,N_17924,N_18833);
or U21816 (N_21816,N_17101,N_15614);
nor U21817 (N_21817,N_17093,N_19441);
xor U21818 (N_21818,N_16669,N_15973);
or U21819 (N_21819,N_19198,N_18375);
or U21820 (N_21820,N_17236,N_19280);
nor U21821 (N_21821,N_19736,N_19371);
or U21822 (N_21822,N_15515,N_15810);
nor U21823 (N_21823,N_18082,N_16435);
nor U21824 (N_21824,N_19909,N_15456);
xnor U21825 (N_21825,N_17687,N_17936);
nand U21826 (N_21826,N_16706,N_15898);
nor U21827 (N_21827,N_16086,N_18432);
and U21828 (N_21828,N_16950,N_18172);
or U21829 (N_21829,N_18556,N_17410);
and U21830 (N_21830,N_18959,N_18456);
xor U21831 (N_21831,N_18540,N_19815);
xor U21832 (N_21832,N_18142,N_15404);
nand U21833 (N_21833,N_19676,N_18946);
xor U21834 (N_21834,N_19614,N_15940);
and U21835 (N_21835,N_18962,N_16763);
and U21836 (N_21836,N_18981,N_16370);
xor U21837 (N_21837,N_17001,N_17533);
or U21838 (N_21838,N_17313,N_19550);
nor U21839 (N_21839,N_15851,N_18333);
or U21840 (N_21840,N_18474,N_17153);
nand U21841 (N_21841,N_16108,N_17049);
xnor U21842 (N_21842,N_17653,N_16369);
or U21843 (N_21843,N_18320,N_18651);
or U21844 (N_21844,N_15423,N_18558);
or U21845 (N_21845,N_15248,N_18130);
and U21846 (N_21846,N_19053,N_17961);
and U21847 (N_21847,N_18369,N_18770);
xor U21848 (N_21848,N_16525,N_15448);
nor U21849 (N_21849,N_19406,N_15406);
or U21850 (N_21850,N_17634,N_18581);
nand U21851 (N_21851,N_15146,N_18009);
xor U21852 (N_21852,N_15290,N_19926);
and U21853 (N_21853,N_15421,N_16303);
xor U21854 (N_21854,N_18287,N_16376);
nor U21855 (N_21855,N_18070,N_15925);
or U21856 (N_21856,N_18176,N_17476);
and U21857 (N_21857,N_19611,N_19932);
and U21858 (N_21858,N_16799,N_17541);
and U21859 (N_21859,N_18674,N_18731);
xor U21860 (N_21860,N_17509,N_17848);
nand U21861 (N_21861,N_17078,N_17426);
nand U21862 (N_21862,N_15764,N_15191);
xor U21863 (N_21863,N_19229,N_18562);
xnor U21864 (N_21864,N_15371,N_18560);
and U21865 (N_21865,N_19812,N_16012);
and U21866 (N_21866,N_17985,N_17597);
nand U21867 (N_21867,N_15642,N_15021);
nor U21868 (N_21868,N_19436,N_16713);
nor U21869 (N_21869,N_15926,N_17361);
or U21870 (N_21870,N_18996,N_17473);
or U21871 (N_21871,N_17569,N_17064);
nor U21872 (N_21872,N_16851,N_19058);
nand U21873 (N_21873,N_17172,N_17290);
nor U21874 (N_21874,N_19641,N_17853);
nand U21875 (N_21875,N_16856,N_15985);
xor U21876 (N_21876,N_17264,N_18755);
xnor U21877 (N_21877,N_19115,N_17739);
or U21878 (N_21878,N_18803,N_19061);
nand U21879 (N_21879,N_16422,N_15652);
xor U21880 (N_21880,N_17043,N_16983);
nand U21881 (N_21881,N_17245,N_17080);
xor U21882 (N_21882,N_16933,N_16340);
xor U21883 (N_21883,N_17041,N_15911);
nor U21884 (N_21884,N_16746,N_16915);
nand U21885 (N_21885,N_17300,N_19882);
and U21886 (N_21886,N_17821,N_15647);
nor U21887 (N_21887,N_17340,N_18635);
nor U21888 (N_21888,N_19850,N_17297);
nor U21889 (N_21889,N_18351,N_19499);
xor U21890 (N_21890,N_18735,N_19554);
nand U21891 (N_21891,N_15534,N_18937);
nor U21892 (N_21892,N_16029,N_18266);
or U21893 (N_21893,N_16227,N_17941);
or U21894 (N_21894,N_15853,N_15199);
or U21895 (N_21895,N_15736,N_19370);
and U21896 (N_21896,N_18067,N_15712);
nand U21897 (N_21897,N_15065,N_18749);
nor U21898 (N_21898,N_18493,N_15312);
xnor U21899 (N_21899,N_18386,N_19302);
and U21900 (N_21900,N_15678,N_15322);
xnor U21901 (N_21901,N_18484,N_17237);
or U21902 (N_21902,N_18982,N_17575);
xnor U21903 (N_21903,N_16296,N_15654);
nor U21904 (N_21904,N_17839,N_19052);
nor U21905 (N_21905,N_17888,N_17874);
xor U21906 (N_21906,N_15930,N_19235);
nor U21907 (N_21907,N_17911,N_19577);
xnor U21908 (N_21908,N_18595,N_17344);
or U21909 (N_21909,N_19834,N_18640);
nor U21910 (N_21910,N_19963,N_16299);
nand U21911 (N_21911,N_15849,N_15969);
or U21912 (N_21912,N_15559,N_17901);
xnor U21913 (N_21913,N_17506,N_15378);
and U21914 (N_21914,N_17573,N_19047);
nor U21915 (N_21915,N_16804,N_16351);
or U21916 (N_21916,N_18354,N_15430);
xor U21917 (N_21917,N_16791,N_16553);
and U21918 (N_21918,N_15435,N_19403);
or U21919 (N_21919,N_18043,N_16853);
or U21920 (N_21920,N_15505,N_16011);
or U21921 (N_21921,N_17685,N_18152);
nand U21922 (N_21922,N_16317,N_15928);
xor U21923 (N_21923,N_16079,N_15956);
or U21924 (N_21924,N_15220,N_17765);
nor U21925 (N_21925,N_17864,N_15243);
xnor U21926 (N_21926,N_19517,N_17453);
nor U21927 (N_21927,N_16785,N_18265);
xor U21928 (N_21928,N_15443,N_19297);
nor U21929 (N_21929,N_19784,N_16149);
and U21930 (N_21930,N_17261,N_16974);
xor U21931 (N_21931,N_19656,N_18454);
nor U21932 (N_21932,N_19090,N_15138);
nand U21933 (N_21933,N_17958,N_18827);
xnor U21934 (N_21934,N_15558,N_19610);
or U21935 (N_21935,N_15059,N_18665);
or U21936 (N_21936,N_19088,N_15244);
and U21937 (N_21937,N_15895,N_16140);
nor U21938 (N_21938,N_15488,N_16000);
nand U21939 (N_21939,N_17117,N_17720);
or U21940 (N_21940,N_19392,N_15390);
and U21941 (N_21941,N_15560,N_16365);
and U21942 (N_21942,N_15232,N_17718);
nor U21943 (N_21943,N_17603,N_19398);
nand U21944 (N_21944,N_17507,N_18797);
nor U21945 (N_21945,N_15933,N_17276);
xor U21946 (N_21946,N_18849,N_19068);
or U21947 (N_21947,N_19093,N_18891);
or U21948 (N_21948,N_16160,N_18451);
or U21949 (N_21949,N_16221,N_17877);
nand U21950 (N_21950,N_15265,N_15754);
nand U21951 (N_21951,N_19450,N_18195);
xnor U21952 (N_21952,N_19629,N_15903);
xnor U21953 (N_21953,N_16224,N_18436);
and U21954 (N_21954,N_17789,N_19382);
nor U21955 (N_21955,N_18864,N_19269);
nor U21956 (N_21956,N_16330,N_19959);
and U21957 (N_21957,N_15340,N_16462);
nand U21958 (N_21958,N_17588,N_19881);
xnor U21959 (N_21959,N_16504,N_16027);
and U21960 (N_21960,N_15636,N_19936);
and U21961 (N_21961,N_17008,N_18653);
and U21962 (N_21962,N_15176,N_16934);
and U21963 (N_21963,N_19817,N_18881);
and U21964 (N_21964,N_18505,N_16382);
and U21965 (N_21965,N_18088,N_15131);
nor U21966 (N_21966,N_17835,N_19533);
xnor U21967 (N_21967,N_19918,N_17933);
or U21968 (N_21968,N_15613,N_18955);
xnor U21969 (N_21969,N_16357,N_17156);
and U21970 (N_21970,N_19272,N_19837);
and U21971 (N_21971,N_18825,N_19608);
and U21972 (N_21972,N_19129,N_17212);
nand U21973 (N_21973,N_16389,N_17278);
xor U21974 (N_21974,N_19769,N_19021);
and U21975 (N_21975,N_15503,N_19348);
and U21976 (N_21976,N_16694,N_15375);
and U21977 (N_21977,N_19708,N_15482);
nand U21978 (N_21978,N_17123,N_18289);
or U21979 (N_21979,N_19661,N_15429);
xnor U21980 (N_21980,N_16557,N_16700);
or U21981 (N_21981,N_19506,N_18260);
or U21982 (N_21982,N_19987,N_16476);
nand U21983 (N_21983,N_19316,N_18186);
and U21984 (N_21984,N_17764,N_19291);
nand U21985 (N_21985,N_18641,N_15646);
and U21986 (N_21986,N_19890,N_17167);
or U21987 (N_21987,N_17672,N_15580);
and U21988 (N_21988,N_17354,N_16334);
nor U21989 (N_21989,N_19418,N_15548);
nand U21990 (N_21990,N_16649,N_16169);
or U21991 (N_21991,N_18764,N_17570);
and U21992 (N_21992,N_19584,N_17191);
and U21993 (N_21993,N_18732,N_18577);
nor U21994 (N_21994,N_17037,N_15527);
nor U21995 (N_21995,N_15765,N_16951);
nor U21996 (N_21996,N_19256,N_16323);
and U21997 (N_21997,N_18052,N_15462);
nand U21998 (N_21998,N_15545,N_15958);
and U21999 (N_21999,N_17675,N_16541);
nand U22000 (N_22000,N_18930,N_16946);
nand U22001 (N_22001,N_17203,N_15242);
xnor U22002 (N_22002,N_19468,N_17689);
or U22003 (N_22003,N_18078,N_19734);
xor U22004 (N_22004,N_19582,N_18695);
and U22005 (N_22005,N_18198,N_18249);
nor U22006 (N_22006,N_16891,N_15701);
nor U22007 (N_22007,N_17490,N_18936);
nor U22008 (N_22008,N_17282,N_17096);
nor U22009 (N_22009,N_18286,N_15224);
or U22010 (N_22010,N_17373,N_19431);
and U22011 (N_22011,N_15792,N_16371);
xor U22012 (N_22012,N_16074,N_18315);
nand U22013 (N_22013,N_17542,N_15946);
nor U22014 (N_22014,N_17170,N_16203);
or U22015 (N_22015,N_19564,N_15164);
nor U22016 (N_22016,N_19408,N_17102);
nor U22017 (N_22017,N_16744,N_18143);
or U22018 (N_22018,N_18039,N_19344);
nand U22019 (N_22019,N_17753,N_16246);
or U22020 (N_22020,N_19603,N_18284);
or U22021 (N_22021,N_15570,N_18117);
nand U22022 (N_22022,N_15586,N_19220);
or U22023 (N_22023,N_16783,N_19420);
and U22024 (N_22024,N_18883,N_18728);
or U22025 (N_22025,N_18406,N_18737);
or U22026 (N_22026,N_16999,N_18566);
xnor U22027 (N_22027,N_15874,N_17317);
nand U22028 (N_22028,N_17120,N_15659);
xor U22029 (N_22029,N_15013,N_19689);
xor U22030 (N_22030,N_18324,N_18716);
xnor U22031 (N_22031,N_16670,N_19793);
nor U22032 (N_22032,N_19639,N_16599);
nand U22033 (N_22033,N_16326,N_19862);
nand U22034 (N_22034,N_16290,N_17467);
xor U22035 (N_22035,N_15735,N_19662);
nand U22036 (N_22036,N_15223,N_16258);
nor U22037 (N_22037,N_17407,N_17162);
nor U22038 (N_22038,N_16889,N_18890);
nand U22039 (N_22039,N_15417,N_16540);
nand U22040 (N_22040,N_16984,N_15751);
nor U22041 (N_22041,N_18648,N_19720);
xor U22042 (N_22042,N_19362,N_16204);
and U22043 (N_22043,N_16864,N_19523);
and U22044 (N_22044,N_17819,N_17155);
and U22045 (N_22045,N_16126,N_15769);
nor U22046 (N_22046,N_17006,N_19059);
and U22047 (N_22047,N_19640,N_16366);
and U22048 (N_22048,N_19989,N_18723);
and U22049 (N_22049,N_16092,N_18498);
nor U22050 (N_22050,N_16979,N_16616);
or U22051 (N_22051,N_17154,N_15990);
or U22052 (N_22052,N_17422,N_16053);
xnor U22053 (N_22053,N_15530,N_18200);
and U22054 (N_22054,N_19879,N_19627);
xnor U22055 (N_22055,N_15400,N_19585);
xnor U22056 (N_22056,N_15305,N_15409);
and U22057 (N_22057,N_18203,N_17886);
and U22058 (N_22058,N_16639,N_16421);
nor U22059 (N_22059,N_16748,N_19323);
xor U22060 (N_22060,N_18114,N_18615);
nand U22061 (N_22061,N_16180,N_16165);
or U22062 (N_22062,N_15590,N_16273);
nand U22063 (N_22063,N_17613,N_16097);
or U22064 (N_22064,N_17732,N_19270);
nand U22065 (N_22065,N_16814,N_15695);
xor U22066 (N_22066,N_19010,N_15480);
nor U22067 (N_22067,N_16867,N_16157);
nand U22068 (N_22068,N_17545,N_17957);
nand U22069 (N_22069,N_18942,N_19565);
nand U22070 (N_22070,N_17861,N_18513);
nand U22071 (N_22071,N_17186,N_18412);
xor U22072 (N_22072,N_16030,N_18921);
xor U22073 (N_22073,N_16127,N_17168);
and U22074 (N_22074,N_15187,N_17596);
and U22075 (N_22075,N_18100,N_19745);
xnor U22076 (N_22076,N_19600,N_16059);
and U22077 (N_22077,N_19422,N_18555);
nand U22078 (N_22078,N_17412,N_19360);
nor U22079 (N_22079,N_15049,N_15716);
nand U22080 (N_22080,N_15125,N_15478);
xnor U22081 (N_22081,N_15288,N_18586);
xor U22082 (N_22082,N_18617,N_17937);
or U22083 (N_22083,N_17291,N_17218);
nand U22084 (N_22084,N_17779,N_19396);
or U22085 (N_22085,N_17374,N_15635);
xnor U22086 (N_22086,N_18694,N_16367);
nand U22087 (N_22087,N_15449,N_15213);
xnor U22088 (N_22088,N_17139,N_19056);
xor U22089 (N_22089,N_16593,N_19530);
xor U22090 (N_22090,N_15127,N_15123);
xor U22091 (N_22091,N_16192,N_18342);
nand U22092 (N_22092,N_15303,N_18518);
or U22093 (N_22093,N_17305,N_16235);
nor U22094 (N_22094,N_19013,N_16840);
and U22095 (N_22095,N_15587,N_16663);
or U22096 (N_22096,N_17606,N_15426);
or U22097 (N_22097,N_18029,N_18550);
or U22098 (N_22098,N_18153,N_17834);
xnor U22099 (N_22099,N_17654,N_17766);
or U22100 (N_22100,N_15846,N_16790);
nor U22101 (N_22101,N_16905,N_19597);
nor U22102 (N_22102,N_19214,N_16166);
nor U22103 (N_22103,N_15821,N_16372);
nor U22104 (N_22104,N_18083,N_17266);
and U22105 (N_22105,N_17221,N_15055);
nand U22106 (N_22106,N_15573,N_16534);
nand U22107 (N_22107,N_17599,N_17873);
nand U22108 (N_22108,N_17989,N_17549);
xnor U22109 (N_22109,N_17491,N_19028);
xnor U22110 (N_22110,N_17301,N_19756);
nand U22111 (N_22111,N_17658,N_15629);
and U22112 (N_22112,N_18278,N_15147);
and U22113 (N_22113,N_18056,N_18757);
xor U22114 (N_22114,N_17872,N_18673);
or U22115 (N_22115,N_15962,N_18892);
or U22116 (N_22116,N_16522,N_16262);
and U22117 (N_22117,N_18915,N_18358);
or U22118 (N_22118,N_16158,N_18434);
nand U22119 (N_22119,N_15813,N_18931);
nor U22120 (N_22120,N_17052,N_17528);
nor U22121 (N_22121,N_18366,N_16261);
and U22122 (N_22122,N_17076,N_17697);
and U22123 (N_22123,N_15218,N_17302);
nor U22124 (N_22124,N_16110,N_19478);
and U22125 (N_22125,N_17244,N_18433);
xor U22126 (N_22126,N_16267,N_17681);
nand U22127 (N_22127,N_15198,N_18170);
or U22128 (N_22128,N_17680,N_15516);
nor U22129 (N_22129,N_16631,N_17181);
nand U22130 (N_22130,N_15253,N_16980);
nor U22131 (N_22131,N_16562,N_19369);
nor U22132 (N_22132,N_18443,N_16394);
nor U22133 (N_22133,N_19029,N_18328);
nor U22134 (N_22134,N_18006,N_15469);
and U22135 (N_22135,N_18398,N_16282);
nor U22136 (N_22136,N_17275,N_18228);
and U22137 (N_22137,N_17954,N_16281);
xor U22138 (N_22138,N_15905,N_15460);
nand U22139 (N_22139,N_16230,N_17147);
and U22140 (N_22140,N_16198,N_17684);
or U22141 (N_22141,N_18071,N_17640);
nor U22142 (N_22142,N_19111,N_16597);
nor U22143 (N_22143,N_19700,N_18384);
nand U22144 (N_22144,N_15604,N_17706);
xor U22145 (N_22145,N_17648,N_15000);
nor U22146 (N_22146,N_18950,N_15023);
nor U22147 (N_22147,N_16824,N_17214);
nand U22148 (N_22148,N_18048,N_15415);
and U22149 (N_22149,N_17075,N_15170);
or U22150 (N_22150,N_19161,N_19075);
nor U22151 (N_22151,N_18929,N_18175);
nand U22152 (N_22152,N_15008,N_18169);
or U22153 (N_22153,N_19884,N_17508);
or U22154 (N_22154,N_18637,N_15563);
nand U22155 (N_22155,N_18462,N_15352);
xor U22156 (N_22156,N_17402,N_16800);
nor U22157 (N_22157,N_15324,N_19258);
xor U22158 (N_22158,N_19292,N_15184);
xor U22159 (N_22159,N_17028,N_18030);
and U22160 (N_22160,N_17882,N_16159);
or U22161 (N_22161,N_19681,N_18585);
nand U22162 (N_22162,N_18592,N_18997);
nand U22163 (N_22163,N_18835,N_19984);
xnor U22164 (N_22164,N_18736,N_16187);
and U22165 (N_22165,N_15360,N_15609);
and U22166 (N_22166,N_16035,N_19073);
and U22167 (N_22167,N_15889,N_18469);
xor U22168 (N_22168,N_17201,N_16003);
nor U22169 (N_22169,N_18845,N_17795);
and U22170 (N_22170,N_16806,N_15149);
and U22171 (N_22171,N_17761,N_19643);
nor U22172 (N_22172,N_17303,N_18086);
xnor U22173 (N_22173,N_16502,N_19599);
and U22174 (N_22174,N_15433,N_15778);
xnor U22175 (N_22175,N_19404,N_18995);
nor U22176 (N_22176,N_17745,N_18567);
and U22177 (N_22177,N_17975,N_19205);
and U22178 (N_22178,N_18972,N_16104);
xnor U22179 (N_22179,N_15965,N_17378);
and U22180 (N_22180,N_15917,N_15348);
xnor U22181 (N_22181,N_16068,N_17783);
xnor U22182 (N_22182,N_17645,N_16341);
and U22183 (N_22183,N_16142,N_17514);
nor U22184 (N_22184,N_17934,N_15321);
nor U22185 (N_22185,N_17772,N_19472);
and U22186 (N_22186,N_17820,N_19078);
or U22187 (N_22187,N_16456,N_18192);
and U22188 (N_22188,N_15978,N_19895);
xnor U22189 (N_22189,N_15709,N_16536);
or U22190 (N_22190,N_19728,N_16285);
xor U22191 (N_22191,N_19779,N_18685);
and U22192 (N_22192,N_18532,N_19318);
nor U22193 (N_22193,N_15051,N_17283);
and U22194 (N_22194,N_18572,N_16447);
or U22195 (N_22195,N_16038,N_15050);
nand U22196 (N_22196,N_16436,N_17352);
nor U22197 (N_22197,N_15795,N_19064);
nand U22198 (N_22198,N_16434,N_18179);
xnor U22199 (N_22199,N_19941,N_17992);
nor U22200 (N_22200,N_17129,N_15350);
nand U22201 (N_22201,N_16052,N_15345);
and U22202 (N_22202,N_17142,N_19946);
and U22203 (N_22203,N_15087,N_17262);
xor U22204 (N_22204,N_18390,N_17100);
xnor U22205 (N_22205,N_19109,N_15579);
nand U22206 (N_22206,N_15599,N_18233);
or U22207 (N_22207,N_17094,N_15357);
and U22208 (N_22208,N_16241,N_17210);
and U22209 (N_22209,N_15714,N_17979);
and U22210 (N_22210,N_19429,N_18430);
and U22211 (N_22211,N_17044,N_18751);
nor U22212 (N_22212,N_16477,N_15987);
or U22213 (N_22213,N_17413,N_15314);
nand U22214 (N_22214,N_15504,N_18545);
nor U22215 (N_22215,N_16982,N_15377);
nand U22216 (N_22216,N_15633,N_17601);
or U22217 (N_22217,N_16415,N_17062);
nor U22218 (N_22218,N_16315,N_19213);
or U22219 (N_22219,N_18542,N_15524);
xor U22220 (N_22220,N_15491,N_15726);
nor U22221 (N_22221,N_15041,N_15292);
xnor U22222 (N_22222,N_16921,N_19098);
nor U22223 (N_22223,N_16807,N_15957);
and U22224 (N_22224,N_18602,N_19039);
and U22225 (N_22225,N_15748,N_18688);
or U22226 (N_22226,N_17539,N_15631);
or U22227 (N_22227,N_18705,N_17927);
and U22228 (N_22228,N_15425,N_15826);
nand U22229 (N_22229,N_15432,N_17353);
xnor U22230 (N_22230,N_17047,N_19320);
nor U22231 (N_22231,N_16816,N_19826);
xor U22232 (N_22232,N_16728,N_19157);
and U22233 (N_22233,N_19546,N_19219);
and U22234 (N_22234,N_15048,N_18738);
nand U22235 (N_22235,N_17787,N_15689);
nor U22236 (N_22236,N_19159,N_16466);
and U22237 (N_22237,N_18396,N_15847);
or U22238 (N_22238,N_19361,N_15837);
and U22239 (N_22239,N_17582,N_19727);
nor U22240 (N_22240,N_15715,N_16356);
xnor U22241 (N_22241,N_16103,N_18644);
xor U22242 (N_22242,N_19567,N_17445);
nor U22243 (N_22243,N_18460,N_18782);
or U22244 (N_22244,N_16155,N_16276);
nand U22245 (N_22245,N_15696,N_15383);
and U22246 (N_22246,N_19916,N_17694);
and U22247 (N_22247,N_17002,N_17796);
nand U22248 (N_22248,N_16342,N_15693);
or U22249 (N_22249,N_15921,N_18989);
xor U22250 (N_22250,N_17758,N_18670);
xor U22251 (N_22251,N_18689,N_17118);
xnor U22252 (N_22252,N_19931,N_18829);
xor U22253 (N_22253,N_19037,N_19050);
xnor U22254 (N_22254,N_17905,N_18193);
nor U22255 (N_22255,N_15734,N_16646);
or U22256 (N_22256,N_19531,N_19244);
nand U22257 (N_22257,N_18626,N_19122);
and U22258 (N_22258,N_18222,N_19801);
nor U22259 (N_22259,N_19082,N_17017);
nand U22260 (N_22260,N_16760,N_19555);
nand U22261 (N_22261,N_15562,N_17416);
nor U22262 (N_22262,N_15888,N_15046);
or U22263 (N_22263,N_19417,N_16153);
or U22264 (N_22264,N_17760,N_19227);
nand U22265 (N_22265,N_17572,N_17331);
xnor U22266 (N_22266,N_17778,N_18213);
nand U22267 (N_22267,N_17748,N_19816);
xnor U22268 (N_22268,N_19786,N_18184);
xnor U22269 (N_22269,N_19015,N_17618);
xor U22270 (N_22270,N_19813,N_19743);
nand U22271 (N_22271,N_16046,N_15100);
and U22272 (N_22272,N_18246,N_17059);
xor U22273 (N_22273,N_17547,N_16687);
xor U22274 (N_22274,N_16396,N_15463);
or U22275 (N_22275,N_17810,N_19512);
or U22276 (N_22276,N_16499,N_19904);
nor U22277 (N_22277,N_17128,N_16820);
xor U22278 (N_22278,N_19975,N_18418);
nand U22279 (N_22279,N_17124,N_19625);
xnor U22280 (N_22280,N_17952,N_18678);
and U22281 (N_22281,N_17339,N_18746);
or U22282 (N_22282,N_16213,N_16482);
nand U22283 (N_22283,N_17161,N_19732);
nor U22284 (N_22284,N_16778,N_19101);
nand U22285 (N_22285,N_18721,N_18715);
nor U22286 (N_22286,N_18262,N_18525);
nand U22287 (N_22287,N_16497,N_15015);
nand U22288 (N_22288,N_17950,N_19773);
nor U22289 (N_22289,N_15717,N_19767);
nor U22290 (N_22290,N_18873,N_17664);
or U22291 (N_22291,N_15062,N_17920);
nor U22292 (N_22292,N_17079,N_15998);
nor U22293 (N_22293,N_19601,N_17478);
and U22294 (N_22294,N_18734,N_19673);
nor U22295 (N_22295,N_19207,N_19223);
or U22296 (N_22296,N_19066,N_17584);
nor U22297 (N_22297,N_15539,N_19459);
nor U22298 (N_22298,N_15342,N_16695);
nor U22299 (N_22299,N_19726,N_17255);
nor U22300 (N_22300,N_16461,N_17364);
nor U22301 (N_22301,N_18692,N_17463);
nor U22302 (N_22302,N_17529,N_15995);
or U22303 (N_22303,N_15785,N_18104);
and U22304 (N_22304,N_17611,N_19041);
nor U22305 (N_22305,N_15057,N_18223);
xnor U22306 (N_22306,N_19521,N_19217);
or U22307 (N_22307,N_19525,N_16375);
or U22308 (N_22308,N_15892,N_19696);
nor U22309 (N_22309,N_15618,N_15666);
nand U22310 (N_22310,N_16409,N_18911);
or U22311 (N_22311,N_18912,N_19947);
or U22312 (N_22312,N_17608,N_19692);
and U22313 (N_22313,N_17607,N_16916);
nand U22314 (N_22314,N_18554,N_16026);
nand U22315 (N_22315,N_15414,N_15781);
nor U22316 (N_22316,N_17727,N_17444);
nand U22317 (N_22317,N_17807,N_16368);
xor U22318 (N_22318,N_19432,N_19350);
nor U22319 (N_22319,N_18243,N_19206);
nor U22320 (N_22320,N_15555,N_19453);
and U22321 (N_22321,N_17973,N_16913);
nor U22322 (N_22322,N_19338,N_19866);
nor U22323 (N_22323,N_18428,N_17649);
and U22324 (N_22324,N_18853,N_19581);
and U22325 (N_22325,N_16653,N_19854);
and U22326 (N_22326,N_16398,N_17306);
or U22327 (N_22327,N_17625,N_15620);
and U22328 (N_22328,N_17999,N_17022);
xor U22329 (N_22329,N_16105,N_16234);
or U22330 (N_22330,N_15079,N_18859);
xnor U22331 (N_22331,N_17656,N_19215);
and U22332 (N_22332,N_18471,N_18900);
xor U22333 (N_22333,N_17782,N_19271);
xor U22334 (N_22334,N_18439,N_15317);
nand U22335 (N_22335,N_15097,N_16787);
xor U22336 (N_22336,N_17832,N_19955);
xor U22337 (N_22337,N_16678,N_15865);
nor U22338 (N_22338,N_19888,N_15833);
and U22339 (N_22339,N_17360,N_18894);
and U22340 (N_22340,N_17368,N_18316);
xor U22341 (N_22341,N_19443,N_19896);
xor U22342 (N_22342,N_19591,N_18145);
and U22343 (N_22343,N_18064,N_19301);
and U22344 (N_22344,N_17459,N_16513);
and U22345 (N_22345,N_18871,N_16014);
nor U22346 (N_22346,N_15436,N_17946);
nand U22347 (N_22347,N_19364,N_17455);
nor U22348 (N_22348,N_16677,N_18240);
xor U22349 (N_22349,N_15188,N_17837);
xnor U22350 (N_22350,N_18247,N_16004);
and U22351 (N_22351,N_18664,N_19820);
nor U22352 (N_22352,N_19666,N_17960);
or U22353 (N_22353,N_15359,N_18148);
nor U22354 (N_22354,N_15148,N_15857);
and U22355 (N_22355,N_16850,N_18111);
xor U22356 (N_22356,N_16170,N_19212);
nor U22357 (N_22357,N_15697,N_15158);
nand U22358 (N_22358,N_19192,N_17567);
nand U22359 (N_22359,N_19355,N_17319);
or U22360 (N_22360,N_18761,N_16360);
or U22361 (N_22361,N_17581,N_16123);
and U22362 (N_22362,N_18426,N_19592);
and U22363 (N_22363,N_16412,N_19425);
and U22364 (N_22364,N_15447,N_15679);
or U22365 (N_22365,N_17454,N_17550);
xnor U22366 (N_22366,N_16569,N_16043);
xnor U22367 (N_22367,N_15247,N_16432);
and U22368 (N_22368,N_17033,N_18856);
and U22369 (N_22369,N_18528,N_17140);
nor U22370 (N_22370,N_19825,N_17173);
xor U22371 (N_22371,N_18706,N_19962);
and U22372 (N_22372,N_16491,N_15954);
and U22373 (N_22373,N_16294,N_18001);
or U22374 (N_22374,N_15500,N_17456);
or U22375 (N_22375,N_17185,N_16468);
xor U22376 (N_22376,N_19241,N_18649);
xor U22377 (N_22377,N_15525,N_15601);
nand U22378 (N_22378,N_16831,N_19138);
nor U22379 (N_22379,N_19133,N_15306);
or U22380 (N_22380,N_18671,N_19349);
and U22381 (N_22381,N_16709,N_16566);
nand U22382 (N_22382,N_17743,N_16928);
nor U22383 (N_22383,N_18115,N_16754);
nand U22384 (N_22384,N_16301,N_17029);
xor U22385 (N_22385,N_16485,N_19322);
nor U22386 (N_22386,N_19294,N_15873);
and U22387 (N_22387,N_17399,N_15189);
nor U22388 (N_22388,N_19299,N_16374);
or U22389 (N_22389,N_19960,N_17977);
nor U22390 (N_22390,N_16987,N_16400);
or U22391 (N_22391,N_19805,N_19785);
xor U22392 (N_22392,N_18405,N_16520);
or U22393 (N_22393,N_16564,N_18259);
nand U22394 (N_22394,N_16829,N_19125);
nor U22395 (N_22395,N_16332,N_19651);
or U22396 (N_22396,N_19324,N_15823);
xor U22397 (N_22397,N_17801,N_17891);
and U22398 (N_22398,N_15313,N_15745);
or U22399 (N_22399,N_16327,N_17752);
and U22400 (N_22400,N_15126,N_18133);
and U22401 (N_22401,N_15038,N_19415);
nand U22402 (N_22402,N_16209,N_18726);
xnor U22403 (N_22403,N_15222,N_15053);
and U22404 (N_22404,N_15467,N_17678);
nor U22405 (N_22405,N_17089,N_16481);
nand U22406 (N_22406,N_15681,N_15880);
xnor U22407 (N_22407,N_16920,N_18402);
xor U22408 (N_22408,N_19796,N_17690);
or U22409 (N_22409,N_18801,N_15112);
or U22410 (N_22410,N_15368,N_18888);
xor U22411 (N_22411,N_16419,N_15388);
or U22412 (N_22412,N_17594,N_15142);
and U22413 (N_22413,N_17112,N_18447);
or U22414 (N_22414,N_16163,N_17446);
nor U22415 (N_22415,N_16955,N_17116);
xor U22416 (N_22416,N_17633,N_15216);
or U22417 (N_22417,N_19149,N_16483);
or U22418 (N_22418,N_19500,N_19479);
nor U22419 (N_22419,N_16292,N_19245);
nor U22420 (N_22420,N_16682,N_16875);
xnor U22421 (N_22421,N_18244,N_19194);
xnor U22422 (N_22422,N_17763,N_18012);
and U22423 (N_22423,N_19999,N_18476);
and U22424 (N_22424,N_17993,N_19185);
and U22425 (N_22425,N_19081,N_16498);
nand U22426 (N_22426,N_19596,N_17501);
and U22427 (N_22427,N_16538,N_15834);
xor U22428 (N_22428,N_18107,N_17027);
nor U22429 (N_22429,N_15729,N_16832);
and U22430 (N_22430,N_18720,N_18633);
nand U22431 (N_22431,N_19124,N_15518);
or U22432 (N_22432,N_19852,N_15323);
nor U22433 (N_22433,N_16608,N_18027);
xnor U22434 (N_22434,N_18658,N_15416);
nor U22435 (N_22435,N_19973,N_16015);
nand U22436 (N_22436,N_15797,N_18042);
nor U22437 (N_22437,N_18187,N_16457);
xnor U22438 (N_22438,N_17320,N_17424);
nor U22439 (N_22439,N_19742,N_15427);
or U22440 (N_22440,N_18538,N_18992);
or U22441 (N_22441,N_15145,N_17197);
or U22442 (N_22442,N_17200,N_17598);
and U22443 (N_22443,N_17063,N_17563);
xnor U22444 (N_22444,N_16040,N_17980);
xnor U22445 (N_22445,N_16845,N_15634);
nor U22446 (N_22446,N_15845,N_16519);
or U22447 (N_22447,N_15867,N_19076);
and U22448 (N_22448,N_19239,N_18106);
or U22449 (N_22449,N_18425,N_16039);
and U22450 (N_22450,N_18404,N_19900);
xnor U22451 (N_22451,N_17555,N_15341);
xor U22452 (N_22452,N_18666,N_15827);
nand U22453 (N_22453,N_19741,N_19137);
xnor U22454 (N_22454,N_17524,N_16633);
and U22455 (N_22455,N_16242,N_16095);
nor U22456 (N_22456,N_15331,N_15574);
nand U22457 (N_22457,N_15233,N_16753);
nor U22458 (N_22458,N_15991,N_16667);
nor U22459 (N_22459,N_17389,N_17998);
nor U22460 (N_22460,N_15310,N_17833);
or U22461 (N_22461,N_18510,N_16226);
xnor U22462 (N_22462,N_19636,N_19464);
nand U22463 (N_22463,N_18466,N_18611);
xnor U22464 (N_22464,N_19903,N_17086);
xnor U22465 (N_22465,N_17908,N_15502);
and U22466 (N_22466,N_18238,N_19626);
nor U22467 (N_22467,N_18879,N_19644);
nor U22468 (N_22468,N_15346,N_18269);
xor U22469 (N_22469,N_16925,N_15030);
and U22470 (N_22470,N_17755,N_17132);
or U22471 (N_22471,N_15902,N_18796);
and U22472 (N_22472,N_15333,N_18625);
nor U22473 (N_22473,N_15094,N_19475);
nor U22474 (N_22474,N_18743,N_18445);
and U22475 (N_22475,N_15344,N_19401);
nand U22476 (N_22476,N_19535,N_15782);
xnor U22477 (N_22477,N_15285,N_15139);
nor U22478 (N_22478,N_18235,N_18926);
and U22479 (N_22479,N_17621,N_17365);
and U22480 (N_22480,N_17935,N_18393);
nand U22481 (N_22481,N_16031,N_15010);
nor U22482 (N_22482,N_19978,N_18840);
nor U22483 (N_22483,N_18399,N_17756);
nand U22484 (N_22484,N_18076,N_17113);
and U22485 (N_22485,N_15739,N_16823);
xor U22486 (N_22486,N_15476,N_18381);
nand U22487 (N_22487,N_15165,N_17050);
or U22488 (N_22488,N_18297,N_19730);
xor U22489 (N_22489,N_17131,N_18818);
and U22490 (N_22490,N_16008,N_17329);
xnor U22491 (N_22491,N_15582,N_16839);
and U22492 (N_22492,N_19023,N_19949);
nor U22493 (N_22493,N_18227,N_15981);
xor U22494 (N_22494,N_16911,N_18795);
or U22495 (N_22495,N_19329,N_18508);
and U22496 (N_22496,N_17065,N_17252);
nand U22497 (N_22497,N_19471,N_16619);
nand U22498 (N_22498,N_18624,N_18359);
nor U22499 (N_22499,N_17496,N_18574);
and U22500 (N_22500,N_18674,N_15108);
and U22501 (N_22501,N_16191,N_18425);
nor U22502 (N_22502,N_16369,N_19736);
or U22503 (N_22503,N_16033,N_15188);
or U22504 (N_22504,N_17894,N_15060);
nor U22505 (N_22505,N_19662,N_18311);
or U22506 (N_22506,N_17884,N_17615);
and U22507 (N_22507,N_15716,N_17867);
or U22508 (N_22508,N_16347,N_19775);
or U22509 (N_22509,N_15919,N_16028);
and U22510 (N_22510,N_18546,N_15952);
or U22511 (N_22511,N_19908,N_19842);
or U22512 (N_22512,N_19634,N_19976);
nor U22513 (N_22513,N_17746,N_17692);
or U22514 (N_22514,N_16273,N_16018);
nor U22515 (N_22515,N_19215,N_16850);
or U22516 (N_22516,N_17516,N_15150);
and U22517 (N_22517,N_19925,N_19045);
nor U22518 (N_22518,N_15347,N_18063);
nand U22519 (N_22519,N_19638,N_17163);
xor U22520 (N_22520,N_18065,N_17605);
or U22521 (N_22521,N_19317,N_17930);
nand U22522 (N_22522,N_17305,N_17037);
nand U22523 (N_22523,N_15188,N_17602);
nand U22524 (N_22524,N_19764,N_16600);
xor U22525 (N_22525,N_16161,N_19906);
nor U22526 (N_22526,N_15987,N_17627);
nand U22527 (N_22527,N_18238,N_15519);
xnor U22528 (N_22528,N_19965,N_19153);
nand U22529 (N_22529,N_15892,N_19718);
or U22530 (N_22530,N_18377,N_18390);
or U22531 (N_22531,N_19824,N_19797);
xor U22532 (N_22532,N_19710,N_15282);
xor U22533 (N_22533,N_15716,N_16344);
and U22534 (N_22534,N_16133,N_17385);
and U22535 (N_22535,N_18611,N_19907);
xnor U22536 (N_22536,N_17898,N_18864);
nand U22537 (N_22537,N_16304,N_16147);
xnor U22538 (N_22538,N_18272,N_17757);
xnor U22539 (N_22539,N_16501,N_16706);
xor U22540 (N_22540,N_16842,N_19238);
nand U22541 (N_22541,N_15927,N_18998);
or U22542 (N_22542,N_19808,N_15050);
and U22543 (N_22543,N_18311,N_15719);
or U22544 (N_22544,N_16101,N_18316);
or U22545 (N_22545,N_15275,N_15347);
nand U22546 (N_22546,N_16981,N_19256);
or U22547 (N_22547,N_18875,N_17219);
nor U22548 (N_22548,N_18619,N_19787);
nand U22549 (N_22549,N_19365,N_18814);
or U22550 (N_22550,N_19616,N_19005);
or U22551 (N_22551,N_18576,N_16541);
nand U22552 (N_22552,N_18906,N_17919);
and U22553 (N_22553,N_19336,N_19843);
xor U22554 (N_22554,N_19146,N_18923);
and U22555 (N_22555,N_15066,N_16491);
nand U22556 (N_22556,N_15277,N_17638);
and U22557 (N_22557,N_18528,N_18777);
or U22558 (N_22558,N_19815,N_17548);
or U22559 (N_22559,N_16547,N_19076);
and U22560 (N_22560,N_16337,N_16989);
nand U22561 (N_22561,N_17737,N_19781);
nor U22562 (N_22562,N_19080,N_17633);
nand U22563 (N_22563,N_15794,N_16690);
nand U22564 (N_22564,N_18364,N_18856);
and U22565 (N_22565,N_19853,N_19723);
and U22566 (N_22566,N_17438,N_18997);
nand U22567 (N_22567,N_19948,N_19541);
nor U22568 (N_22568,N_18257,N_15307);
nor U22569 (N_22569,N_17555,N_19383);
or U22570 (N_22570,N_18318,N_18145);
nand U22571 (N_22571,N_18598,N_18601);
xnor U22572 (N_22572,N_17059,N_19996);
or U22573 (N_22573,N_19014,N_19886);
or U22574 (N_22574,N_16649,N_17317);
or U22575 (N_22575,N_18762,N_18912);
nor U22576 (N_22576,N_15995,N_16841);
xor U22577 (N_22577,N_18795,N_18093);
nand U22578 (N_22578,N_15211,N_16567);
nor U22579 (N_22579,N_17292,N_15030);
or U22580 (N_22580,N_19818,N_16580);
or U22581 (N_22581,N_17308,N_17553);
xor U22582 (N_22582,N_17337,N_16217);
and U22583 (N_22583,N_18386,N_19218);
nand U22584 (N_22584,N_19634,N_19000);
nor U22585 (N_22585,N_17159,N_17792);
and U22586 (N_22586,N_19021,N_15780);
nor U22587 (N_22587,N_15904,N_17648);
nor U22588 (N_22588,N_18177,N_17723);
or U22589 (N_22589,N_16806,N_17722);
or U22590 (N_22590,N_18474,N_18034);
and U22591 (N_22591,N_17230,N_17800);
and U22592 (N_22592,N_16297,N_19387);
nand U22593 (N_22593,N_15651,N_16517);
nand U22594 (N_22594,N_17111,N_18988);
xor U22595 (N_22595,N_19352,N_16934);
xnor U22596 (N_22596,N_19003,N_19567);
nand U22597 (N_22597,N_17206,N_19839);
xnor U22598 (N_22598,N_18225,N_18829);
or U22599 (N_22599,N_18719,N_17323);
and U22600 (N_22600,N_15475,N_15357);
and U22601 (N_22601,N_17296,N_15518);
and U22602 (N_22602,N_17892,N_19164);
nand U22603 (N_22603,N_17647,N_18779);
nand U22604 (N_22604,N_15946,N_15599);
nand U22605 (N_22605,N_19725,N_15955);
and U22606 (N_22606,N_16546,N_17829);
xor U22607 (N_22607,N_16532,N_19914);
xor U22608 (N_22608,N_18552,N_16771);
nand U22609 (N_22609,N_15944,N_19675);
nor U22610 (N_22610,N_18196,N_17599);
nor U22611 (N_22611,N_15106,N_15919);
nor U22612 (N_22612,N_17599,N_16315);
and U22613 (N_22613,N_19409,N_17940);
xor U22614 (N_22614,N_17328,N_18482);
nand U22615 (N_22615,N_15642,N_15910);
xor U22616 (N_22616,N_16699,N_17037);
nand U22617 (N_22617,N_17412,N_16563);
nor U22618 (N_22618,N_17992,N_16493);
nand U22619 (N_22619,N_19673,N_17223);
xor U22620 (N_22620,N_17837,N_17421);
nand U22621 (N_22621,N_18138,N_15642);
or U22622 (N_22622,N_15900,N_15420);
nand U22623 (N_22623,N_18703,N_18990);
or U22624 (N_22624,N_17033,N_19409);
or U22625 (N_22625,N_15880,N_18096);
and U22626 (N_22626,N_15251,N_17940);
and U22627 (N_22627,N_15398,N_16113);
nand U22628 (N_22628,N_18111,N_17789);
nor U22629 (N_22629,N_17948,N_19257);
and U22630 (N_22630,N_15797,N_18094);
and U22631 (N_22631,N_16905,N_19639);
and U22632 (N_22632,N_15853,N_16013);
nor U22633 (N_22633,N_16022,N_19805);
nand U22634 (N_22634,N_17519,N_17303);
and U22635 (N_22635,N_15111,N_16534);
and U22636 (N_22636,N_15839,N_19351);
nand U22637 (N_22637,N_17714,N_17935);
nor U22638 (N_22638,N_19822,N_15463);
and U22639 (N_22639,N_18159,N_19579);
nand U22640 (N_22640,N_17073,N_16046);
xor U22641 (N_22641,N_17508,N_15825);
and U22642 (N_22642,N_19600,N_17815);
xor U22643 (N_22643,N_16969,N_17249);
or U22644 (N_22644,N_15943,N_16077);
nand U22645 (N_22645,N_18811,N_17764);
and U22646 (N_22646,N_19497,N_17488);
nor U22647 (N_22647,N_17182,N_19169);
or U22648 (N_22648,N_16099,N_17722);
nor U22649 (N_22649,N_15558,N_15988);
or U22650 (N_22650,N_15311,N_19571);
nand U22651 (N_22651,N_16562,N_17793);
or U22652 (N_22652,N_19976,N_18585);
and U22653 (N_22653,N_18522,N_18616);
nand U22654 (N_22654,N_17851,N_17375);
nor U22655 (N_22655,N_19939,N_17207);
xor U22656 (N_22656,N_17888,N_16118);
and U22657 (N_22657,N_17507,N_17387);
nor U22658 (N_22658,N_19578,N_16971);
and U22659 (N_22659,N_18799,N_15829);
nor U22660 (N_22660,N_19806,N_17968);
xnor U22661 (N_22661,N_18266,N_15446);
nand U22662 (N_22662,N_16887,N_15644);
xor U22663 (N_22663,N_16113,N_16992);
xnor U22664 (N_22664,N_15858,N_18348);
or U22665 (N_22665,N_17426,N_18111);
nand U22666 (N_22666,N_18299,N_17463);
xnor U22667 (N_22667,N_16449,N_19498);
xor U22668 (N_22668,N_16520,N_19720);
or U22669 (N_22669,N_16983,N_16310);
nor U22670 (N_22670,N_19989,N_15141);
and U22671 (N_22671,N_15654,N_16137);
or U22672 (N_22672,N_15044,N_18972);
nor U22673 (N_22673,N_18641,N_18062);
and U22674 (N_22674,N_18918,N_19900);
or U22675 (N_22675,N_17162,N_16980);
nand U22676 (N_22676,N_15466,N_18351);
nand U22677 (N_22677,N_17761,N_17127);
nand U22678 (N_22678,N_16130,N_19315);
nand U22679 (N_22679,N_18208,N_19206);
or U22680 (N_22680,N_16814,N_16043);
or U22681 (N_22681,N_18053,N_15379);
nand U22682 (N_22682,N_17982,N_16416);
nor U22683 (N_22683,N_19968,N_18861);
nand U22684 (N_22684,N_17744,N_17862);
xnor U22685 (N_22685,N_16596,N_18791);
or U22686 (N_22686,N_19735,N_17244);
xnor U22687 (N_22687,N_17786,N_15744);
or U22688 (N_22688,N_18481,N_18888);
or U22689 (N_22689,N_18660,N_16777);
nor U22690 (N_22690,N_16156,N_19521);
nor U22691 (N_22691,N_18274,N_15110);
or U22692 (N_22692,N_16171,N_17025);
nand U22693 (N_22693,N_19730,N_16185);
and U22694 (N_22694,N_17970,N_19395);
or U22695 (N_22695,N_16745,N_15089);
and U22696 (N_22696,N_16489,N_15095);
nor U22697 (N_22697,N_16572,N_17451);
nand U22698 (N_22698,N_18695,N_17717);
nand U22699 (N_22699,N_18937,N_19720);
nor U22700 (N_22700,N_16108,N_18794);
nor U22701 (N_22701,N_18718,N_19867);
xor U22702 (N_22702,N_18289,N_16884);
xnor U22703 (N_22703,N_17816,N_18851);
nor U22704 (N_22704,N_17797,N_15598);
xnor U22705 (N_22705,N_19184,N_18509);
or U22706 (N_22706,N_16363,N_18220);
or U22707 (N_22707,N_19522,N_15055);
and U22708 (N_22708,N_15145,N_18410);
and U22709 (N_22709,N_16483,N_16201);
nand U22710 (N_22710,N_19241,N_17959);
nor U22711 (N_22711,N_17000,N_16501);
nor U22712 (N_22712,N_17987,N_19424);
xnor U22713 (N_22713,N_16989,N_17744);
and U22714 (N_22714,N_19550,N_17547);
nand U22715 (N_22715,N_19953,N_19400);
and U22716 (N_22716,N_16739,N_17707);
nand U22717 (N_22717,N_15606,N_19196);
nor U22718 (N_22718,N_19776,N_19693);
xor U22719 (N_22719,N_18442,N_16482);
nor U22720 (N_22720,N_17481,N_17823);
nand U22721 (N_22721,N_19557,N_16780);
and U22722 (N_22722,N_18534,N_18820);
nor U22723 (N_22723,N_18619,N_17290);
nand U22724 (N_22724,N_18375,N_15898);
xor U22725 (N_22725,N_16080,N_15405);
and U22726 (N_22726,N_17333,N_17634);
and U22727 (N_22727,N_18134,N_16805);
and U22728 (N_22728,N_15465,N_17209);
nand U22729 (N_22729,N_19461,N_16833);
nand U22730 (N_22730,N_18776,N_19493);
and U22731 (N_22731,N_18590,N_17621);
nor U22732 (N_22732,N_15608,N_17199);
nor U22733 (N_22733,N_17717,N_16033);
xor U22734 (N_22734,N_19612,N_16897);
nand U22735 (N_22735,N_16583,N_17368);
and U22736 (N_22736,N_15438,N_19419);
and U22737 (N_22737,N_19534,N_19510);
or U22738 (N_22738,N_17116,N_15611);
xnor U22739 (N_22739,N_18672,N_19166);
or U22740 (N_22740,N_19544,N_19526);
xnor U22741 (N_22741,N_17552,N_17568);
or U22742 (N_22742,N_19736,N_19447);
nand U22743 (N_22743,N_15152,N_16767);
nor U22744 (N_22744,N_16882,N_16696);
and U22745 (N_22745,N_18011,N_16667);
xor U22746 (N_22746,N_15696,N_18030);
or U22747 (N_22747,N_16297,N_17420);
or U22748 (N_22748,N_15441,N_16987);
or U22749 (N_22749,N_15184,N_18364);
nor U22750 (N_22750,N_19033,N_15030);
or U22751 (N_22751,N_19697,N_19830);
xor U22752 (N_22752,N_18557,N_17940);
nand U22753 (N_22753,N_19369,N_15520);
nand U22754 (N_22754,N_19837,N_15307);
nor U22755 (N_22755,N_17653,N_19570);
xnor U22756 (N_22756,N_16614,N_15981);
nand U22757 (N_22757,N_17438,N_19718);
xnor U22758 (N_22758,N_16689,N_15505);
xnor U22759 (N_22759,N_16347,N_18612);
nor U22760 (N_22760,N_15033,N_15162);
or U22761 (N_22761,N_19193,N_19815);
nand U22762 (N_22762,N_17236,N_18217);
nor U22763 (N_22763,N_16184,N_18490);
nor U22764 (N_22764,N_16075,N_16544);
nand U22765 (N_22765,N_18719,N_19646);
nor U22766 (N_22766,N_17971,N_15881);
nor U22767 (N_22767,N_18245,N_19810);
xnor U22768 (N_22768,N_17254,N_19330);
xnor U22769 (N_22769,N_15126,N_18191);
or U22770 (N_22770,N_15714,N_18554);
xnor U22771 (N_22771,N_16701,N_16320);
nor U22772 (N_22772,N_15108,N_19855);
nand U22773 (N_22773,N_19252,N_15552);
nand U22774 (N_22774,N_19607,N_17122);
nor U22775 (N_22775,N_18501,N_16117);
or U22776 (N_22776,N_15620,N_17631);
nor U22777 (N_22777,N_16337,N_17290);
xnor U22778 (N_22778,N_15346,N_17689);
nor U22779 (N_22779,N_18606,N_19897);
xor U22780 (N_22780,N_19737,N_19252);
or U22781 (N_22781,N_17997,N_15728);
nor U22782 (N_22782,N_16145,N_18551);
xnor U22783 (N_22783,N_15199,N_16597);
xnor U22784 (N_22784,N_16042,N_15902);
xor U22785 (N_22785,N_19649,N_16401);
and U22786 (N_22786,N_19576,N_15805);
or U22787 (N_22787,N_15525,N_16464);
nor U22788 (N_22788,N_16479,N_15149);
and U22789 (N_22789,N_15389,N_15469);
nand U22790 (N_22790,N_16547,N_15745);
xor U22791 (N_22791,N_17425,N_16278);
or U22792 (N_22792,N_19504,N_17996);
nand U22793 (N_22793,N_16838,N_19369);
or U22794 (N_22794,N_16712,N_15277);
and U22795 (N_22795,N_16885,N_18022);
nor U22796 (N_22796,N_15291,N_16115);
nor U22797 (N_22797,N_18171,N_15504);
and U22798 (N_22798,N_19698,N_15609);
xnor U22799 (N_22799,N_18878,N_16532);
and U22800 (N_22800,N_19390,N_15970);
nand U22801 (N_22801,N_16944,N_18148);
or U22802 (N_22802,N_17692,N_18462);
and U22803 (N_22803,N_19342,N_16374);
xnor U22804 (N_22804,N_19105,N_19809);
nand U22805 (N_22805,N_17644,N_19967);
or U22806 (N_22806,N_19800,N_18193);
nor U22807 (N_22807,N_16865,N_19964);
xnor U22808 (N_22808,N_16320,N_18154);
nor U22809 (N_22809,N_15208,N_17927);
nor U22810 (N_22810,N_17396,N_15659);
nor U22811 (N_22811,N_15880,N_18418);
nand U22812 (N_22812,N_17301,N_15220);
xor U22813 (N_22813,N_16632,N_17874);
nand U22814 (N_22814,N_17480,N_19807);
and U22815 (N_22815,N_19049,N_19493);
nor U22816 (N_22816,N_17439,N_16570);
nand U22817 (N_22817,N_18055,N_19265);
nand U22818 (N_22818,N_15181,N_16542);
xnor U22819 (N_22819,N_17125,N_15616);
and U22820 (N_22820,N_18806,N_15682);
nor U22821 (N_22821,N_15575,N_18862);
nand U22822 (N_22822,N_15360,N_17771);
nor U22823 (N_22823,N_17132,N_18862);
and U22824 (N_22824,N_19166,N_18198);
xnor U22825 (N_22825,N_17862,N_16724);
nor U22826 (N_22826,N_17235,N_19504);
or U22827 (N_22827,N_19224,N_19533);
xor U22828 (N_22828,N_19787,N_18909);
or U22829 (N_22829,N_15671,N_19167);
nor U22830 (N_22830,N_16211,N_18217);
or U22831 (N_22831,N_19015,N_19010);
nand U22832 (N_22832,N_17609,N_16970);
nand U22833 (N_22833,N_16989,N_19698);
xor U22834 (N_22834,N_15055,N_15694);
or U22835 (N_22835,N_18754,N_16789);
and U22836 (N_22836,N_18275,N_16597);
xor U22837 (N_22837,N_16817,N_18928);
or U22838 (N_22838,N_16149,N_19587);
and U22839 (N_22839,N_18277,N_16256);
or U22840 (N_22840,N_15102,N_17505);
and U22841 (N_22841,N_15766,N_19933);
nor U22842 (N_22842,N_19522,N_19250);
xnor U22843 (N_22843,N_17898,N_17360);
and U22844 (N_22844,N_15621,N_16484);
xor U22845 (N_22845,N_17206,N_17357);
nand U22846 (N_22846,N_17864,N_19882);
nor U22847 (N_22847,N_19145,N_19975);
xor U22848 (N_22848,N_16796,N_18507);
nor U22849 (N_22849,N_19158,N_16985);
or U22850 (N_22850,N_15194,N_17715);
or U22851 (N_22851,N_19323,N_19887);
or U22852 (N_22852,N_15203,N_19859);
nor U22853 (N_22853,N_19088,N_19891);
nand U22854 (N_22854,N_19726,N_18501);
nand U22855 (N_22855,N_17979,N_15416);
xnor U22856 (N_22856,N_15689,N_18233);
nor U22857 (N_22857,N_19978,N_18313);
nor U22858 (N_22858,N_16385,N_18700);
nand U22859 (N_22859,N_19048,N_19844);
and U22860 (N_22860,N_15435,N_18304);
or U22861 (N_22861,N_18547,N_18242);
and U22862 (N_22862,N_17852,N_17792);
nor U22863 (N_22863,N_15762,N_18869);
nand U22864 (N_22864,N_15826,N_19018);
nand U22865 (N_22865,N_18396,N_18630);
nor U22866 (N_22866,N_18272,N_17319);
and U22867 (N_22867,N_15956,N_19510);
or U22868 (N_22868,N_16658,N_15684);
xor U22869 (N_22869,N_18672,N_15077);
or U22870 (N_22870,N_15559,N_18482);
xnor U22871 (N_22871,N_18686,N_15329);
or U22872 (N_22872,N_18683,N_19681);
nand U22873 (N_22873,N_17520,N_19268);
nand U22874 (N_22874,N_17916,N_18627);
and U22875 (N_22875,N_15960,N_17558);
or U22876 (N_22876,N_16593,N_17309);
nand U22877 (N_22877,N_18242,N_16992);
or U22878 (N_22878,N_19066,N_18401);
and U22879 (N_22879,N_15945,N_18539);
and U22880 (N_22880,N_17790,N_16636);
and U22881 (N_22881,N_16321,N_15105);
nand U22882 (N_22882,N_15584,N_18167);
nand U22883 (N_22883,N_15997,N_15826);
nor U22884 (N_22884,N_18178,N_16251);
or U22885 (N_22885,N_15196,N_19958);
xor U22886 (N_22886,N_15644,N_15289);
or U22887 (N_22887,N_18409,N_15815);
xnor U22888 (N_22888,N_18771,N_16104);
nand U22889 (N_22889,N_19300,N_17375);
or U22890 (N_22890,N_15470,N_18484);
xor U22891 (N_22891,N_19058,N_17716);
xor U22892 (N_22892,N_16225,N_17630);
or U22893 (N_22893,N_19513,N_18187);
and U22894 (N_22894,N_16283,N_19280);
xnor U22895 (N_22895,N_18815,N_15142);
nand U22896 (N_22896,N_17887,N_15368);
xnor U22897 (N_22897,N_15333,N_18017);
nor U22898 (N_22898,N_18766,N_18320);
and U22899 (N_22899,N_15203,N_17351);
or U22900 (N_22900,N_19973,N_16945);
or U22901 (N_22901,N_18112,N_17965);
or U22902 (N_22902,N_18712,N_16050);
nor U22903 (N_22903,N_16741,N_16277);
and U22904 (N_22904,N_17798,N_17525);
xnor U22905 (N_22905,N_19526,N_19440);
nand U22906 (N_22906,N_18221,N_15954);
or U22907 (N_22907,N_16879,N_17659);
or U22908 (N_22908,N_17129,N_17625);
or U22909 (N_22909,N_19749,N_18490);
xor U22910 (N_22910,N_19956,N_16834);
xnor U22911 (N_22911,N_18786,N_15298);
nand U22912 (N_22912,N_17379,N_19192);
and U22913 (N_22913,N_18630,N_16380);
nor U22914 (N_22914,N_19208,N_19667);
and U22915 (N_22915,N_15772,N_16574);
nor U22916 (N_22916,N_19121,N_17388);
nor U22917 (N_22917,N_18378,N_15794);
or U22918 (N_22918,N_18465,N_18700);
and U22919 (N_22919,N_18556,N_19523);
nand U22920 (N_22920,N_16587,N_19741);
and U22921 (N_22921,N_18422,N_15403);
nand U22922 (N_22922,N_15855,N_17592);
xnor U22923 (N_22923,N_18212,N_15420);
xor U22924 (N_22924,N_17833,N_17553);
and U22925 (N_22925,N_15898,N_17726);
or U22926 (N_22926,N_17728,N_19642);
xnor U22927 (N_22927,N_16836,N_18069);
nor U22928 (N_22928,N_16643,N_16507);
and U22929 (N_22929,N_19043,N_15453);
xor U22930 (N_22930,N_17535,N_15743);
nor U22931 (N_22931,N_17738,N_19416);
and U22932 (N_22932,N_16284,N_16632);
xnor U22933 (N_22933,N_16099,N_15833);
xnor U22934 (N_22934,N_17165,N_17931);
xnor U22935 (N_22935,N_19511,N_16370);
nor U22936 (N_22936,N_19067,N_17230);
nor U22937 (N_22937,N_15686,N_17481);
nand U22938 (N_22938,N_19277,N_17078);
or U22939 (N_22939,N_17348,N_16971);
nor U22940 (N_22940,N_16604,N_18805);
nor U22941 (N_22941,N_16960,N_17846);
and U22942 (N_22942,N_16440,N_17456);
nand U22943 (N_22943,N_15426,N_15945);
nor U22944 (N_22944,N_16302,N_18438);
and U22945 (N_22945,N_16213,N_15913);
or U22946 (N_22946,N_18318,N_15383);
or U22947 (N_22947,N_16938,N_16854);
nand U22948 (N_22948,N_16110,N_18583);
nand U22949 (N_22949,N_18646,N_16862);
nand U22950 (N_22950,N_15012,N_18191);
nor U22951 (N_22951,N_19449,N_16683);
and U22952 (N_22952,N_16300,N_18826);
or U22953 (N_22953,N_17545,N_18643);
xor U22954 (N_22954,N_17103,N_16407);
and U22955 (N_22955,N_19837,N_15059);
nor U22956 (N_22956,N_18665,N_15105);
xnor U22957 (N_22957,N_19247,N_18567);
nor U22958 (N_22958,N_19596,N_17434);
or U22959 (N_22959,N_17069,N_16945);
nor U22960 (N_22960,N_16909,N_18266);
and U22961 (N_22961,N_16534,N_15390);
and U22962 (N_22962,N_18549,N_17016);
nand U22963 (N_22963,N_18697,N_18365);
or U22964 (N_22964,N_17190,N_19580);
nor U22965 (N_22965,N_15714,N_17149);
and U22966 (N_22966,N_19927,N_17702);
nand U22967 (N_22967,N_18266,N_18285);
nand U22968 (N_22968,N_16836,N_19559);
nor U22969 (N_22969,N_19293,N_18008);
xor U22970 (N_22970,N_19959,N_17624);
nor U22971 (N_22971,N_17212,N_17071);
and U22972 (N_22972,N_15246,N_16892);
and U22973 (N_22973,N_15380,N_15333);
nand U22974 (N_22974,N_18016,N_16508);
or U22975 (N_22975,N_18989,N_18759);
nand U22976 (N_22976,N_16593,N_15840);
xor U22977 (N_22977,N_16452,N_15142);
or U22978 (N_22978,N_15276,N_18280);
nand U22979 (N_22979,N_17880,N_16895);
nor U22980 (N_22980,N_16204,N_15573);
and U22981 (N_22981,N_18066,N_15976);
nor U22982 (N_22982,N_18494,N_17088);
nor U22983 (N_22983,N_15922,N_18827);
and U22984 (N_22984,N_17940,N_18835);
and U22985 (N_22985,N_16863,N_16454);
and U22986 (N_22986,N_18104,N_16218);
nor U22987 (N_22987,N_19989,N_16282);
or U22988 (N_22988,N_15511,N_18522);
and U22989 (N_22989,N_16176,N_16291);
xor U22990 (N_22990,N_19658,N_15380);
and U22991 (N_22991,N_15863,N_19816);
and U22992 (N_22992,N_15187,N_17603);
nand U22993 (N_22993,N_17403,N_15217);
nand U22994 (N_22994,N_15558,N_15901);
or U22995 (N_22995,N_15234,N_16724);
nor U22996 (N_22996,N_18882,N_17599);
or U22997 (N_22997,N_17239,N_17730);
xnor U22998 (N_22998,N_19185,N_16439);
or U22999 (N_22999,N_17523,N_18325);
or U23000 (N_23000,N_17125,N_17713);
xor U23001 (N_23001,N_17617,N_19255);
nor U23002 (N_23002,N_16519,N_16354);
nand U23003 (N_23003,N_17330,N_17020);
xor U23004 (N_23004,N_19703,N_19520);
and U23005 (N_23005,N_16943,N_17622);
or U23006 (N_23006,N_16423,N_18784);
nand U23007 (N_23007,N_18415,N_15429);
xnor U23008 (N_23008,N_17579,N_17848);
and U23009 (N_23009,N_15963,N_15309);
or U23010 (N_23010,N_16283,N_17464);
nand U23011 (N_23011,N_16127,N_15511);
xor U23012 (N_23012,N_19268,N_16971);
or U23013 (N_23013,N_17590,N_17232);
or U23014 (N_23014,N_16142,N_19864);
xor U23015 (N_23015,N_19818,N_16606);
or U23016 (N_23016,N_18557,N_15050);
xor U23017 (N_23017,N_15159,N_19331);
nand U23018 (N_23018,N_18698,N_19387);
and U23019 (N_23019,N_18861,N_19179);
and U23020 (N_23020,N_16731,N_16925);
and U23021 (N_23021,N_16384,N_17781);
xor U23022 (N_23022,N_16428,N_19471);
or U23023 (N_23023,N_16996,N_18611);
or U23024 (N_23024,N_15094,N_17186);
or U23025 (N_23025,N_19430,N_16349);
and U23026 (N_23026,N_17074,N_19988);
and U23027 (N_23027,N_15020,N_15240);
nand U23028 (N_23028,N_19555,N_19175);
nand U23029 (N_23029,N_18471,N_16003);
and U23030 (N_23030,N_17701,N_17912);
and U23031 (N_23031,N_17677,N_19034);
xor U23032 (N_23032,N_15761,N_15834);
and U23033 (N_23033,N_19108,N_15426);
or U23034 (N_23034,N_17331,N_19290);
or U23035 (N_23035,N_18809,N_17940);
and U23036 (N_23036,N_19102,N_19266);
xnor U23037 (N_23037,N_18635,N_19808);
or U23038 (N_23038,N_17965,N_16628);
nand U23039 (N_23039,N_15044,N_16890);
xor U23040 (N_23040,N_17866,N_18107);
nand U23041 (N_23041,N_17516,N_17368);
or U23042 (N_23042,N_19210,N_15361);
nand U23043 (N_23043,N_16991,N_18591);
xor U23044 (N_23044,N_16673,N_17552);
or U23045 (N_23045,N_19524,N_15155);
nor U23046 (N_23046,N_17472,N_17708);
or U23047 (N_23047,N_16963,N_16619);
and U23048 (N_23048,N_15820,N_19977);
nand U23049 (N_23049,N_19887,N_16429);
nand U23050 (N_23050,N_18296,N_19282);
nor U23051 (N_23051,N_16617,N_17112);
nand U23052 (N_23052,N_15506,N_19019);
xnor U23053 (N_23053,N_16812,N_19161);
and U23054 (N_23054,N_17009,N_19522);
nor U23055 (N_23055,N_19980,N_18710);
nor U23056 (N_23056,N_17262,N_19968);
xor U23057 (N_23057,N_15165,N_15424);
nand U23058 (N_23058,N_18706,N_18989);
or U23059 (N_23059,N_17128,N_18330);
and U23060 (N_23060,N_18140,N_18190);
nor U23061 (N_23061,N_15688,N_17205);
or U23062 (N_23062,N_16666,N_18399);
nand U23063 (N_23063,N_17983,N_18275);
nor U23064 (N_23064,N_16810,N_15380);
xor U23065 (N_23065,N_17911,N_16908);
or U23066 (N_23066,N_19128,N_18709);
nor U23067 (N_23067,N_17893,N_19803);
xnor U23068 (N_23068,N_19959,N_18746);
or U23069 (N_23069,N_17241,N_16429);
or U23070 (N_23070,N_18897,N_16066);
and U23071 (N_23071,N_17459,N_18427);
and U23072 (N_23072,N_17022,N_18717);
nor U23073 (N_23073,N_19138,N_19525);
nand U23074 (N_23074,N_19144,N_17065);
xor U23075 (N_23075,N_18907,N_16721);
nor U23076 (N_23076,N_16754,N_19031);
and U23077 (N_23077,N_16619,N_16364);
nand U23078 (N_23078,N_19615,N_15912);
or U23079 (N_23079,N_16297,N_15993);
nand U23080 (N_23080,N_15592,N_16008);
xnor U23081 (N_23081,N_16801,N_19313);
xnor U23082 (N_23082,N_15806,N_16619);
xor U23083 (N_23083,N_18028,N_16947);
nand U23084 (N_23084,N_15628,N_15580);
nor U23085 (N_23085,N_16336,N_17581);
nand U23086 (N_23086,N_15876,N_16227);
nand U23087 (N_23087,N_16740,N_19896);
or U23088 (N_23088,N_19332,N_18481);
or U23089 (N_23089,N_16582,N_16991);
nor U23090 (N_23090,N_17402,N_15144);
xor U23091 (N_23091,N_15809,N_16060);
and U23092 (N_23092,N_15689,N_15715);
and U23093 (N_23093,N_18801,N_17718);
nand U23094 (N_23094,N_19599,N_17845);
nand U23095 (N_23095,N_15143,N_16070);
nor U23096 (N_23096,N_17591,N_18246);
nor U23097 (N_23097,N_18626,N_16537);
nor U23098 (N_23098,N_17530,N_15176);
nand U23099 (N_23099,N_17266,N_18853);
nand U23100 (N_23100,N_17154,N_16963);
and U23101 (N_23101,N_16870,N_15670);
or U23102 (N_23102,N_17915,N_18773);
nand U23103 (N_23103,N_15531,N_18549);
xor U23104 (N_23104,N_19621,N_15490);
and U23105 (N_23105,N_17654,N_17147);
and U23106 (N_23106,N_16817,N_19803);
or U23107 (N_23107,N_17869,N_19204);
nor U23108 (N_23108,N_15455,N_16743);
xnor U23109 (N_23109,N_18261,N_18711);
xor U23110 (N_23110,N_15073,N_18799);
nand U23111 (N_23111,N_15477,N_18660);
and U23112 (N_23112,N_19685,N_18359);
xor U23113 (N_23113,N_16990,N_15317);
or U23114 (N_23114,N_16713,N_15013);
or U23115 (N_23115,N_17079,N_16719);
nand U23116 (N_23116,N_17347,N_15109);
and U23117 (N_23117,N_15676,N_15652);
or U23118 (N_23118,N_15977,N_19304);
and U23119 (N_23119,N_16749,N_16999);
nand U23120 (N_23120,N_15480,N_16332);
or U23121 (N_23121,N_19983,N_17937);
nor U23122 (N_23122,N_15955,N_19224);
or U23123 (N_23123,N_19713,N_18436);
nand U23124 (N_23124,N_18376,N_19390);
xor U23125 (N_23125,N_18767,N_16030);
and U23126 (N_23126,N_17257,N_15984);
nand U23127 (N_23127,N_19108,N_15038);
and U23128 (N_23128,N_19301,N_15491);
nor U23129 (N_23129,N_19544,N_15999);
xnor U23130 (N_23130,N_16812,N_18019);
nor U23131 (N_23131,N_17254,N_17602);
nand U23132 (N_23132,N_18266,N_19081);
or U23133 (N_23133,N_17476,N_15693);
nor U23134 (N_23134,N_19619,N_15291);
nor U23135 (N_23135,N_16325,N_18599);
and U23136 (N_23136,N_17954,N_19140);
xor U23137 (N_23137,N_17590,N_19657);
nand U23138 (N_23138,N_16731,N_17191);
or U23139 (N_23139,N_15223,N_19683);
and U23140 (N_23140,N_19941,N_18462);
nor U23141 (N_23141,N_19159,N_16579);
xnor U23142 (N_23142,N_18807,N_18842);
or U23143 (N_23143,N_18207,N_15983);
xor U23144 (N_23144,N_17519,N_18698);
nand U23145 (N_23145,N_15071,N_19957);
xnor U23146 (N_23146,N_19228,N_18820);
nand U23147 (N_23147,N_15353,N_19273);
or U23148 (N_23148,N_17252,N_17800);
nand U23149 (N_23149,N_16054,N_15223);
and U23150 (N_23150,N_18878,N_16918);
xnor U23151 (N_23151,N_15212,N_17284);
and U23152 (N_23152,N_16084,N_15916);
or U23153 (N_23153,N_15463,N_18112);
or U23154 (N_23154,N_19744,N_17446);
xnor U23155 (N_23155,N_16490,N_17649);
nor U23156 (N_23156,N_16862,N_15563);
and U23157 (N_23157,N_17277,N_16032);
and U23158 (N_23158,N_17142,N_19601);
or U23159 (N_23159,N_17677,N_18257);
or U23160 (N_23160,N_16008,N_16038);
or U23161 (N_23161,N_19546,N_18742);
xor U23162 (N_23162,N_16980,N_15316);
or U23163 (N_23163,N_15192,N_16133);
nor U23164 (N_23164,N_18220,N_17306);
nand U23165 (N_23165,N_18431,N_15245);
or U23166 (N_23166,N_18511,N_16258);
and U23167 (N_23167,N_17838,N_19341);
or U23168 (N_23168,N_16634,N_15286);
nand U23169 (N_23169,N_19709,N_15052);
nor U23170 (N_23170,N_19715,N_17832);
nand U23171 (N_23171,N_19871,N_19767);
xor U23172 (N_23172,N_16866,N_17948);
xor U23173 (N_23173,N_18019,N_16483);
nand U23174 (N_23174,N_15904,N_15701);
xnor U23175 (N_23175,N_18371,N_17675);
nor U23176 (N_23176,N_19205,N_18753);
and U23177 (N_23177,N_19613,N_15133);
xnor U23178 (N_23178,N_19032,N_16355);
or U23179 (N_23179,N_19972,N_15167);
nor U23180 (N_23180,N_19163,N_18630);
nand U23181 (N_23181,N_19875,N_15402);
or U23182 (N_23182,N_17764,N_16464);
xor U23183 (N_23183,N_18666,N_15043);
or U23184 (N_23184,N_16738,N_15511);
nand U23185 (N_23185,N_19359,N_17193);
and U23186 (N_23186,N_16534,N_19934);
xnor U23187 (N_23187,N_15324,N_16747);
nor U23188 (N_23188,N_15349,N_19601);
nand U23189 (N_23189,N_19367,N_17009);
xor U23190 (N_23190,N_16898,N_15288);
and U23191 (N_23191,N_15503,N_18462);
and U23192 (N_23192,N_16638,N_18704);
xor U23193 (N_23193,N_16629,N_16341);
xor U23194 (N_23194,N_15698,N_15213);
xor U23195 (N_23195,N_15501,N_17946);
nand U23196 (N_23196,N_15352,N_17068);
nor U23197 (N_23197,N_16193,N_15244);
or U23198 (N_23198,N_16750,N_17388);
or U23199 (N_23199,N_19994,N_16603);
nand U23200 (N_23200,N_19768,N_15023);
nand U23201 (N_23201,N_18208,N_15969);
xnor U23202 (N_23202,N_16214,N_17183);
or U23203 (N_23203,N_19810,N_17047);
and U23204 (N_23204,N_17399,N_17999);
nand U23205 (N_23205,N_17902,N_16053);
or U23206 (N_23206,N_19355,N_19184);
or U23207 (N_23207,N_15590,N_15148);
and U23208 (N_23208,N_17411,N_17900);
xor U23209 (N_23209,N_15021,N_15968);
nand U23210 (N_23210,N_16429,N_18261);
xnor U23211 (N_23211,N_19428,N_16412);
nand U23212 (N_23212,N_19938,N_16200);
xor U23213 (N_23213,N_15514,N_17906);
nor U23214 (N_23214,N_16538,N_16053);
and U23215 (N_23215,N_19885,N_16742);
xor U23216 (N_23216,N_16172,N_19920);
nor U23217 (N_23217,N_19554,N_17372);
xnor U23218 (N_23218,N_16955,N_17806);
nand U23219 (N_23219,N_15318,N_19517);
nor U23220 (N_23220,N_19070,N_19199);
xnor U23221 (N_23221,N_19854,N_15131);
nand U23222 (N_23222,N_15852,N_16470);
xnor U23223 (N_23223,N_18505,N_17634);
xor U23224 (N_23224,N_17179,N_17107);
and U23225 (N_23225,N_15702,N_19776);
xnor U23226 (N_23226,N_16683,N_18885);
nand U23227 (N_23227,N_16534,N_18802);
nand U23228 (N_23228,N_17597,N_18241);
and U23229 (N_23229,N_17287,N_15455);
and U23230 (N_23230,N_19499,N_18492);
nor U23231 (N_23231,N_16361,N_15269);
or U23232 (N_23232,N_18773,N_19665);
or U23233 (N_23233,N_16856,N_17388);
or U23234 (N_23234,N_16281,N_16590);
nor U23235 (N_23235,N_15728,N_18191);
nand U23236 (N_23236,N_19429,N_19431);
or U23237 (N_23237,N_16808,N_19647);
and U23238 (N_23238,N_16138,N_15735);
and U23239 (N_23239,N_18585,N_16824);
xnor U23240 (N_23240,N_17184,N_17197);
and U23241 (N_23241,N_15041,N_19390);
or U23242 (N_23242,N_18879,N_15647);
and U23243 (N_23243,N_18197,N_15434);
xor U23244 (N_23244,N_15129,N_15182);
nor U23245 (N_23245,N_17464,N_17825);
nor U23246 (N_23246,N_17604,N_16498);
xnor U23247 (N_23247,N_16600,N_17531);
or U23248 (N_23248,N_16281,N_18160);
nor U23249 (N_23249,N_19437,N_18255);
and U23250 (N_23250,N_16163,N_15165);
xnor U23251 (N_23251,N_18640,N_17646);
nor U23252 (N_23252,N_15760,N_19774);
or U23253 (N_23253,N_19641,N_16632);
xnor U23254 (N_23254,N_16295,N_16059);
or U23255 (N_23255,N_16897,N_19210);
and U23256 (N_23256,N_15290,N_16579);
nand U23257 (N_23257,N_18820,N_16543);
nand U23258 (N_23258,N_17216,N_17282);
nand U23259 (N_23259,N_17327,N_16224);
nand U23260 (N_23260,N_17389,N_19507);
or U23261 (N_23261,N_17843,N_17819);
xor U23262 (N_23262,N_15797,N_18499);
xnor U23263 (N_23263,N_15946,N_15458);
nor U23264 (N_23264,N_19466,N_17294);
nand U23265 (N_23265,N_18762,N_18813);
xnor U23266 (N_23266,N_19063,N_17872);
nor U23267 (N_23267,N_16129,N_17227);
nor U23268 (N_23268,N_16313,N_15886);
or U23269 (N_23269,N_17385,N_19964);
or U23270 (N_23270,N_19990,N_16704);
nand U23271 (N_23271,N_15559,N_19965);
and U23272 (N_23272,N_15671,N_15767);
or U23273 (N_23273,N_17314,N_17267);
xor U23274 (N_23274,N_15365,N_15095);
and U23275 (N_23275,N_15798,N_18925);
nand U23276 (N_23276,N_15269,N_15498);
xor U23277 (N_23277,N_15339,N_17041);
xor U23278 (N_23278,N_16324,N_16450);
or U23279 (N_23279,N_15743,N_17745);
xnor U23280 (N_23280,N_16030,N_15476);
nand U23281 (N_23281,N_16290,N_16105);
or U23282 (N_23282,N_17705,N_17259);
and U23283 (N_23283,N_18411,N_17406);
and U23284 (N_23284,N_19919,N_16658);
or U23285 (N_23285,N_19326,N_18510);
or U23286 (N_23286,N_15412,N_16578);
and U23287 (N_23287,N_18295,N_17030);
xor U23288 (N_23288,N_15223,N_16183);
xor U23289 (N_23289,N_15330,N_18815);
xnor U23290 (N_23290,N_15102,N_18090);
and U23291 (N_23291,N_18897,N_16160);
and U23292 (N_23292,N_19374,N_17687);
nand U23293 (N_23293,N_16787,N_15085);
nand U23294 (N_23294,N_17997,N_19430);
and U23295 (N_23295,N_19386,N_16757);
nor U23296 (N_23296,N_15255,N_17425);
and U23297 (N_23297,N_19585,N_18245);
nor U23298 (N_23298,N_18002,N_16867);
and U23299 (N_23299,N_16267,N_16502);
xor U23300 (N_23300,N_17288,N_19797);
nor U23301 (N_23301,N_15122,N_16726);
nor U23302 (N_23302,N_17539,N_18504);
or U23303 (N_23303,N_19548,N_16439);
nor U23304 (N_23304,N_18177,N_19074);
and U23305 (N_23305,N_18939,N_18493);
xnor U23306 (N_23306,N_16315,N_17606);
nand U23307 (N_23307,N_18505,N_18777);
and U23308 (N_23308,N_16455,N_18107);
nor U23309 (N_23309,N_17877,N_17472);
nor U23310 (N_23310,N_17005,N_15785);
and U23311 (N_23311,N_15716,N_16900);
nor U23312 (N_23312,N_19270,N_17087);
and U23313 (N_23313,N_16669,N_17788);
and U23314 (N_23314,N_17045,N_17991);
or U23315 (N_23315,N_17328,N_16698);
and U23316 (N_23316,N_17136,N_18826);
or U23317 (N_23317,N_18847,N_16626);
nand U23318 (N_23318,N_18122,N_15750);
nand U23319 (N_23319,N_19978,N_18608);
or U23320 (N_23320,N_16888,N_18139);
or U23321 (N_23321,N_19040,N_18739);
nor U23322 (N_23322,N_19417,N_16912);
or U23323 (N_23323,N_16300,N_17066);
nand U23324 (N_23324,N_17177,N_18049);
nor U23325 (N_23325,N_17740,N_15754);
nor U23326 (N_23326,N_19467,N_16593);
or U23327 (N_23327,N_17075,N_16550);
nand U23328 (N_23328,N_16116,N_19183);
or U23329 (N_23329,N_15223,N_19982);
nor U23330 (N_23330,N_17007,N_15388);
nor U23331 (N_23331,N_16065,N_18403);
or U23332 (N_23332,N_15635,N_15376);
nand U23333 (N_23333,N_15382,N_19002);
or U23334 (N_23334,N_19239,N_18486);
and U23335 (N_23335,N_19387,N_16901);
or U23336 (N_23336,N_18858,N_15798);
nor U23337 (N_23337,N_15191,N_16722);
and U23338 (N_23338,N_16539,N_17776);
nor U23339 (N_23339,N_15918,N_17239);
nor U23340 (N_23340,N_16413,N_19309);
and U23341 (N_23341,N_15374,N_16187);
nor U23342 (N_23342,N_15237,N_16725);
nor U23343 (N_23343,N_19558,N_15421);
nand U23344 (N_23344,N_17608,N_17800);
and U23345 (N_23345,N_15950,N_17398);
xor U23346 (N_23346,N_19057,N_15348);
nand U23347 (N_23347,N_17228,N_17875);
nand U23348 (N_23348,N_19599,N_17516);
or U23349 (N_23349,N_15098,N_15169);
nand U23350 (N_23350,N_16539,N_16971);
xor U23351 (N_23351,N_19311,N_15084);
xor U23352 (N_23352,N_17089,N_15883);
xnor U23353 (N_23353,N_17869,N_16532);
and U23354 (N_23354,N_19135,N_19666);
or U23355 (N_23355,N_17245,N_19160);
and U23356 (N_23356,N_18220,N_19783);
xnor U23357 (N_23357,N_18345,N_17178);
xor U23358 (N_23358,N_15275,N_17672);
or U23359 (N_23359,N_17593,N_15725);
and U23360 (N_23360,N_18297,N_17130);
and U23361 (N_23361,N_16943,N_19777);
nand U23362 (N_23362,N_18171,N_17750);
nor U23363 (N_23363,N_16254,N_16110);
nor U23364 (N_23364,N_17735,N_16494);
nand U23365 (N_23365,N_18495,N_15258);
nor U23366 (N_23366,N_16680,N_18014);
or U23367 (N_23367,N_15698,N_17917);
or U23368 (N_23368,N_19199,N_17450);
or U23369 (N_23369,N_15681,N_17320);
and U23370 (N_23370,N_15909,N_18308);
and U23371 (N_23371,N_19188,N_17172);
nor U23372 (N_23372,N_17696,N_19102);
nor U23373 (N_23373,N_17926,N_15945);
and U23374 (N_23374,N_17429,N_19343);
nand U23375 (N_23375,N_16328,N_19143);
xor U23376 (N_23376,N_19766,N_15261);
nor U23377 (N_23377,N_18432,N_15978);
nand U23378 (N_23378,N_18737,N_18065);
or U23379 (N_23379,N_17706,N_18334);
xor U23380 (N_23380,N_17468,N_19604);
or U23381 (N_23381,N_15850,N_18578);
nand U23382 (N_23382,N_19789,N_15260);
nand U23383 (N_23383,N_16503,N_16551);
or U23384 (N_23384,N_15414,N_19326);
nor U23385 (N_23385,N_17099,N_15651);
xnor U23386 (N_23386,N_16186,N_18387);
or U23387 (N_23387,N_19147,N_18221);
or U23388 (N_23388,N_19146,N_18432);
nor U23389 (N_23389,N_16133,N_17286);
and U23390 (N_23390,N_18697,N_15311);
nand U23391 (N_23391,N_19065,N_17124);
or U23392 (N_23392,N_19640,N_19452);
and U23393 (N_23393,N_19044,N_16225);
xnor U23394 (N_23394,N_15254,N_15850);
nor U23395 (N_23395,N_17589,N_16308);
nand U23396 (N_23396,N_19911,N_16699);
xnor U23397 (N_23397,N_15024,N_18663);
nand U23398 (N_23398,N_17922,N_17296);
xor U23399 (N_23399,N_18180,N_16664);
xor U23400 (N_23400,N_17724,N_19687);
and U23401 (N_23401,N_15412,N_17116);
nand U23402 (N_23402,N_17939,N_15404);
and U23403 (N_23403,N_19515,N_19444);
or U23404 (N_23404,N_17267,N_15217);
or U23405 (N_23405,N_15784,N_16863);
nand U23406 (N_23406,N_17498,N_15106);
or U23407 (N_23407,N_19212,N_19087);
nand U23408 (N_23408,N_15642,N_16258);
nand U23409 (N_23409,N_18635,N_19593);
nand U23410 (N_23410,N_16408,N_19635);
and U23411 (N_23411,N_15445,N_17957);
or U23412 (N_23412,N_19052,N_16003);
nand U23413 (N_23413,N_16217,N_16547);
and U23414 (N_23414,N_17049,N_15638);
or U23415 (N_23415,N_15647,N_15501);
and U23416 (N_23416,N_18098,N_18868);
xnor U23417 (N_23417,N_15291,N_17122);
xnor U23418 (N_23418,N_19135,N_16265);
nand U23419 (N_23419,N_18696,N_15358);
nand U23420 (N_23420,N_16444,N_16598);
nand U23421 (N_23421,N_19808,N_15098);
xnor U23422 (N_23422,N_15512,N_16651);
or U23423 (N_23423,N_18304,N_18356);
or U23424 (N_23424,N_19270,N_19553);
nor U23425 (N_23425,N_18759,N_15305);
or U23426 (N_23426,N_18409,N_15228);
nor U23427 (N_23427,N_15712,N_15850);
nand U23428 (N_23428,N_16368,N_15725);
or U23429 (N_23429,N_15533,N_16018);
nand U23430 (N_23430,N_17630,N_19874);
nor U23431 (N_23431,N_19772,N_16122);
nor U23432 (N_23432,N_18121,N_15170);
and U23433 (N_23433,N_16145,N_18290);
nand U23434 (N_23434,N_16298,N_19206);
nand U23435 (N_23435,N_18207,N_15201);
or U23436 (N_23436,N_18869,N_15021);
xnor U23437 (N_23437,N_15636,N_16199);
xnor U23438 (N_23438,N_16712,N_19769);
or U23439 (N_23439,N_15155,N_17688);
nor U23440 (N_23440,N_19605,N_17706);
and U23441 (N_23441,N_17671,N_17258);
and U23442 (N_23442,N_19770,N_19776);
xor U23443 (N_23443,N_19589,N_19701);
nor U23444 (N_23444,N_19537,N_17301);
nand U23445 (N_23445,N_17797,N_17402);
xor U23446 (N_23446,N_15880,N_16785);
nor U23447 (N_23447,N_18994,N_19398);
nor U23448 (N_23448,N_19879,N_17482);
or U23449 (N_23449,N_15391,N_16324);
or U23450 (N_23450,N_18707,N_18125);
and U23451 (N_23451,N_15265,N_16521);
nand U23452 (N_23452,N_18117,N_19895);
and U23453 (N_23453,N_15165,N_18967);
nor U23454 (N_23454,N_19885,N_19300);
or U23455 (N_23455,N_18053,N_16337);
and U23456 (N_23456,N_15914,N_19908);
xor U23457 (N_23457,N_17003,N_17004);
or U23458 (N_23458,N_19064,N_17631);
or U23459 (N_23459,N_15729,N_17624);
nand U23460 (N_23460,N_19493,N_15507);
nand U23461 (N_23461,N_19711,N_19412);
xor U23462 (N_23462,N_15674,N_19715);
nor U23463 (N_23463,N_15458,N_15512);
nor U23464 (N_23464,N_17584,N_18891);
or U23465 (N_23465,N_17277,N_18844);
nand U23466 (N_23466,N_17468,N_15294);
and U23467 (N_23467,N_17680,N_19301);
xnor U23468 (N_23468,N_19743,N_19079);
or U23469 (N_23469,N_19346,N_18381);
xor U23470 (N_23470,N_16615,N_17509);
and U23471 (N_23471,N_17309,N_16315);
nand U23472 (N_23472,N_17695,N_18195);
and U23473 (N_23473,N_17149,N_19773);
and U23474 (N_23474,N_17750,N_19224);
nor U23475 (N_23475,N_16887,N_17107);
and U23476 (N_23476,N_17260,N_19972);
xnor U23477 (N_23477,N_15597,N_19452);
nand U23478 (N_23478,N_18797,N_19983);
nand U23479 (N_23479,N_19063,N_18299);
nor U23480 (N_23480,N_15154,N_15758);
nor U23481 (N_23481,N_18206,N_17022);
or U23482 (N_23482,N_19739,N_16852);
and U23483 (N_23483,N_17918,N_18150);
and U23484 (N_23484,N_15163,N_18368);
xor U23485 (N_23485,N_17622,N_18762);
and U23486 (N_23486,N_19671,N_16670);
or U23487 (N_23487,N_18227,N_15675);
nand U23488 (N_23488,N_16775,N_18640);
nand U23489 (N_23489,N_19705,N_16352);
and U23490 (N_23490,N_16901,N_18588);
xor U23491 (N_23491,N_16450,N_16705);
nor U23492 (N_23492,N_16012,N_16463);
nor U23493 (N_23493,N_15805,N_17626);
or U23494 (N_23494,N_16962,N_18493);
xor U23495 (N_23495,N_18896,N_17657);
nor U23496 (N_23496,N_15704,N_19827);
or U23497 (N_23497,N_16257,N_15941);
xnor U23498 (N_23498,N_16330,N_18694);
and U23499 (N_23499,N_17810,N_15024);
nor U23500 (N_23500,N_18110,N_16625);
nand U23501 (N_23501,N_17687,N_17676);
or U23502 (N_23502,N_18115,N_18730);
or U23503 (N_23503,N_18632,N_15487);
and U23504 (N_23504,N_17936,N_18971);
or U23505 (N_23505,N_17744,N_19033);
and U23506 (N_23506,N_18994,N_16117);
or U23507 (N_23507,N_19510,N_17403);
xnor U23508 (N_23508,N_19029,N_17370);
or U23509 (N_23509,N_18102,N_15482);
nand U23510 (N_23510,N_15072,N_15755);
nand U23511 (N_23511,N_15940,N_19957);
and U23512 (N_23512,N_15434,N_18097);
or U23513 (N_23513,N_16869,N_16880);
or U23514 (N_23514,N_19106,N_19163);
nand U23515 (N_23515,N_15611,N_15913);
nor U23516 (N_23516,N_18471,N_16408);
and U23517 (N_23517,N_19174,N_15148);
and U23518 (N_23518,N_18981,N_17306);
and U23519 (N_23519,N_18648,N_17776);
xor U23520 (N_23520,N_15765,N_17726);
nor U23521 (N_23521,N_16766,N_17115);
and U23522 (N_23522,N_18889,N_16641);
nand U23523 (N_23523,N_17943,N_19258);
xnor U23524 (N_23524,N_15045,N_19400);
xor U23525 (N_23525,N_17733,N_19404);
nor U23526 (N_23526,N_18205,N_17180);
nor U23527 (N_23527,N_18666,N_17690);
xnor U23528 (N_23528,N_16416,N_16584);
xnor U23529 (N_23529,N_18107,N_17743);
or U23530 (N_23530,N_15993,N_16194);
and U23531 (N_23531,N_17677,N_19093);
or U23532 (N_23532,N_15044,N_19629);
and U23533 (N_23533,N_16603,N_17051);
and U23534 (N_23534,N_18088,N_18781);
nor U23535 (N_23535,N_19067,N_17922);
nor U23536 (N_23536,N_16855,N_15053);
or U23537 (N_23537,N_17567,N_18103);
xnor U23538 (N_23538,N_17754,N_19206);
or U23539 (N_23539,N_18526,N_16425);
nor U23540 (N_23540,N_17625,N_18277);
nand U23541 (N_23541,N_15872,N_19535);
nor U23542 (N_23542,N_18984,N_19904);
nand U23543 (N_23543,N_18663,N_16892);
or U23544 (N_23544,N_18150,N_19205);
or U23545 (N_23545,N_17784,N_15783);
nand U23546 (N_23546,N_17802,N_17581);
nor U23547 (N_23547,N_17006,N_17499);
xnor U23548 (N_23548,N_19711,N_18035);
and U23549 (N_23549,N_18910,N_15447);
nor U23550 (N_23550,N_19008,N_17595);
and U23551 (N_23551,N_17956,N_18539);
and U23552 (N_23552,N_19963,N_18871);
nor U23553 (N_23553,N_16859,N_15515);
and U23554 (N_23554,N_17471,N_19160);
or U23555 (N_23555,N_17620,N_15637);
nand U23556 (N_23556,N_15222,N_18822);
and U23557 (N_23557,N_19993,N_15002);
xor U23558 (N_23558,N_19610,N_18188);
and U23559 (N_23559,N_17715,N_16495);
and U23560 (N_23560,N_15297,N_15451);
xor U23561 (N_23561,N_16071,N_19110);
xnor U23562 (N_23562,N_16259,N_18586);
or U23563 (N_23563,N_19584,N_16786);
nor U23564 (N_23564,N_18227,N_15200);
xor U23565 (N_23565,N_16305,N_16968);
xor U23566 (N_23566,N_17457,N_19796);
nand U23567 (N_23567,N_18679,N_15803);
nor U23568 (N_23568,N_15176,N_19768);
or U23569 (N_23569,N_17921,N_17074);
nor U23570 (N_23570,N_16682,N_18483);
nor U23571 (N_23571,N_19981,N_16085);
nor U23572 (N_23572,N_15903,N_17521);
and U23573 (N_23573,N_15314,N_17204);
or U23574 (N_23574,N_18359,N_15500);
xor U23575 (N_23575,N_16188,N_16086);
nor U23576 (N_23576,N_19831,N_15291);
or U23577 (N_23577,N_15190,N_17688);
nand U23578 (N_23578,N_15021,N_18009);
and U23579 (N_23579,N_19941,N_16393);
nor U23580 (N_23580,N_18551,N_18376);
or U23581 (N_23581,N_19027,N_18398);
nand U23582 (N_23582,N_16716,N_17956);
and U23583 (N_23583,N_16938,N_17790);
nand U23584 (N_23584,N_16381,N_16967);
nor U23585 (N_23585,N_17155,N_18933);
xnor U23586 (N_23586,N_17761,N_18993);
nor U23587 (N_23587,N_17673,N_17229);
xor U23588 (N_23588,N_15990,N_15883);
xor U23589 (N_23589,N_16916,N_19024);
and U23590 (N_23590,N_19763,N_15665);
nor U23591 (N_23591,N_18898,N_15258);
nor U23592 (N_23592,N_16925,N_16161);
xor U23593 (N_23593,N_18839,N_15834);
nand U23594 (N_23594,N_16002,N_17495);
or U23595 (N_23595,N_16916,N_18685);
nand U23596 (N_23596,N_18757,N_16820);
xor U23597 (N_23597,N_18325,N_18356);
or U23598 (N_23598,N_18550,N_15598);
and U23599 (N_23599,N_19660,N_18762);
and U23600 (N_23600,N_18406,N_15913);
or U23601 (N_23601,N_16689,N_19954);
and U23602 (N_23602,N_17223,N_18097);
nand U23603 (N_23603,N_17840,N_17320);
and U23604 (N_23604,N_17185,N_16242);
or U23605 (N_23605,N_18356,N_16708);
or U23606 (N_23606,N_16902,N_19847);
or U23607 (N_23607,N_16048,N_19265);
or U23608 (N_23608,N_16113,N_17052);
xor U23609 (N_23609,N_16803,N_15398);
xor U23610 (N_23610,N_17613,N_18788);
nor U23611 (N_23611,N_17153,N_17262);
nor U23612 (N_23612,N_15925,N_19661);
nor U23613 (N_23613,N_19368,N_19018);
or U23614 (N_23614,N_15333,N_18433);
nand U23615 (N_23615,N_17112,N_16410);
nor U23616 (N_23616,N_19071,N_15238);
nor U23617 (N_23617,N_17819,N_18379);
nor U23618 (N_23618,N_18043,N_16793);
or U23619 (N_23619,N_18030,N_15438);
and U23620 (N_23620,N_18477,N_19649);
xnor U23621 (N_23621,N_19323,N_16216);
nor U23622 (N_23622,N_15568,N_18669);
nor U23623 (N_23623,N_18266,N_18111);
nand U23624 (N_23624,N_19138,N_19560);
xnor U23625 (N_23625,N_16795,N_15485);
and U23626 (N_23626,N_15394,N_17269);
and U23627 (N_23627,N_17828,N_16323);
and U23628 (N_23628,N_19483,N_18488);
xor U23629 (N_23629,N_17385,N_16531);
or U23630 (N_23630,N_17461,N_19256);
nand U23631 (N_23631,N_16787,N_16430);
nor U23632 (N_23632,N_17300,N_15171);
or U23633 (N_23633,N_16277,N_18782);
xor U23634 (N_23634,N_15281,N_16393);
or U23635 (N_23635,N_15453,N_19153);
nand U23636 (N_23636,N_16098,N_16153);
or U23637 (N_23637,N_18051,N_16663);
xnor U23638 (N_23638,N_15857,N_18378);
and U23639 (N_23639,N_16041,N_16805);
and U23640 (N_23640,N_15343,N_18528);
nor U23641 (N_23641,N_17450,N_17004);
or U23642 (N_23642,N_19871,N_19573);
and U23643 (N_23643,N_17710,N_19330);
and U23644 (N_23644,N_18356,N_15052);
xor U23645 (N_23645,N_18403,N_17258);
or U23646 (N_23646,N_18620,N_16556);
and U23647 (N_23647,N_19047,N_16792);
and U23648 (N_23648,N_15163,N_18942);
nand U23649 (N_23649,N_17843,N_19436);
xor U23650 (N_23650,N_17403,N_15083);
and U23651 (N_23651,N_19247,N_15321);
nand U23652 (N_23652,N_17969,N_19713);
nand U23653 (N_23653,N_18895,N_17107);
nor U23654 (N_23654,N_18135,N_18347);
nand U23655 (N_23655,N_17443,N_17221);
or U23656 (N_23656,N_18533,N_15474);
and U23657 (N_23657,N_15806,N_15755);
nor U23658 (N_23658,N_17791,N_19381);
or U23659 (N_23659,N_17059,N_15552);
nand U23660 (N_23660,N_16097,N_17953);
or U23661 (N_23661,N_17184,N_19415);
nand U23662 (N_23662,N_16396,N_15987);
and U23663 (N_23663,N_17987,N_15266);
or U23664 (N_23664,N_16718,N_19740);
nand U23665 (N_23665,N_19750,N_17130);
and U23666 (N_23666,N_15883,N_19205);
xor U23667 (N_23667,N_15925,N_19232);
or U23668 (N_23668,N_19986,N_18963);
nand U23669 (N_23669,N_17910,N_15770);
nor U23670 (N_23670,N_15451,N_16939);
and U23671 (N_23671,N_17028,N_17222);
nand U23672 (N_23672,N_16056,N_15129);
and U23673 (N_23673,N_19168,N_16601);
nand U23674 (N_23674,N_18476,N_15277);
and U23675 (N_23675,N_16176,N_17736);
nand U23676 (N_23676,N_17922,N_17727);
nand U23677 (N_23677,N_15705,N_17671);
and U23678 (N_23678,N_15213,N_15328);
xnor U23679 (N_23679,N_16302,N_15327);
nor U23680 (N_23680,N_15979,N_16479);
xnor U23681 (N_23681,N_18119,N_19863);
or U23682 (N_23682,N_18611,N_15530);
xnor U23683 (N_23683,N_18684,N_19908);
nor U23684 (N_23684,N_16080,N_15305);
xor U23685 (N_23685,N_16740,N_18509);
nor U23686 (N_23686,N_16269,N_19189);
or U23687 (N_23687,N_15570,N_19362);
or U23688 (N_23688,N_19904,N_17429);
xor U23689 (N_23689,N_19483,N_18514);
or U23690 (N_23690,N_17551,N_16167);
and U23691 (N_23691,N_18772,N_18285);
and U23692 (N_23692,N_17462,N_18524);
and U23693 (N_23693,N_19986,N_17547);
nand U23694 (N_23694,N_15716,N_18933);
or U23695 (N_23695,N_17727,N_18540);
and U23696 (N_23696,N_17840,N_17103);
and U23697 (N_23697,N_17351,N_17400);
nor U23698 (N_23698,N_17629,N_15179);
and U23699 (N_23699,N_18339,N_17262);
nor U23700 (N_23700,N_18054,N_18384);
xor U23701 (N_23701,N_17788,N_15802);
xor U23702 (N_23702,N_18479,N_18467);
nand U23703 (N_23703,N_16740,N_18570);
and U23704 (N_23704,N_16723,N_15616);
and U23705 (N_23705,N_19806,N_15743);
nand U23706 (N_23706,N_18288,N_18950);
nor U23707 (N_23707,N_15385,N_18139);
or U23708 (N_23708,N_18338,N_19007);
or U23709 (N_23709,N_18104,N_16183);
and U23710 (N_23710,N_17257,N_17979);
nor U23711 (N_23711,N_17601,N_15997);
xor U23712 (N_23712,N_18363,N_18838);
nor U23713 (N_23713,N_19890,N_15435);
nor U23714 (N_23714,N_15090,N_15792);
or U23715 (N_23715,N_17932,N_19269);
and U23716 (N_23716,N_16204,N_18579);
or U23717 (N_23717,N_19433,N_19001);
or U23718 (N_23718,N_16795,N_15180);
nor U23719 (N_23719,N_19004,N_16691);
and U23720 (N_23720,N_18642,N_15456);
nor U23721 (N_23721,N_19862,N_18127);
and U23722 (N_23722,N_16487,N_17234);
xor U23723 (N_23723,N_17270,N_18666);
and U23724 (N_23724,N_15828,N_15754);
nand U23725 (N_23725,N_19137,N_18454);
and U23726 (N_23726,N_17007,N_19542);
and U23727 (N_23727,N_18594,N_19857);
nor U23728 (N_23728,N_15281,N_15930);
or U23729 (N_23729,N_17221,N_18362);
or U23730 (N_23730,N_15344,N_18434);
or U23731 (N_23731,N_18411,N_19220);
nor U23732 (N_23732,N_19273,N_17472);
and U23733 (N_23733,N_16718,N_19441);
or U23734 (N_23734,N_18333,N_17860);
nand U23735 (N_23735,N_19030,N_15593);
nand U23736 (N_23736,N_19371,N_18074);
and U23737 (N_23737,N_15323,N_17010);
or U23738 (N_23738,N_16993,N_18606);
nand U23739 (N_23739,N_17993,N_18167);
or U23740 (N_23740,N_18135,N_16864);
xnor U23741 (N_23741,N_17981,N_17674);
nor U23742 (N_23742,N_18720,N_16739);
or U23743 (N_23743,N_16933,N_18974);
nand U23744 (N_23744,N_15112,N_16308);
and U23745 (N_23745,N_15562,N_17104);
nor U23746 (N_23746,N_18076,N_17741);
and U23747 (N_23747,N_15649,N_17193);
nor U23748 (N_23748,N_18143,N_19209);
nand U23749 (N_23749,N_19098,N_18639);
and U23750 (N_23750,N_15604,N_18937);
xor U23751 (N_23751,N_15669,N_19712);
xnor U23752 (N_23752,N_19158,N_17408);
or U23753 (N_23753,N_16467,N_18600);
and U23754 (N_23754,N_15518,N_16192);
or U23755 (N_23755,N_15692,N_18784);
nor U23756 (N_23756,N_15127,N_16245);
xor U23757 (N_23757,N_16111,N_16624);
xor U23758 (N_23758,N_15155,N_15123);
nand U23759 (N_23759,N_17275,N_15113);
xor U23760 (N_23760,N_15806,N_19931);
and U23761 (N_23761,N_17773,N_19394);
nand U23762 (N_23762,N_18296,N_16431);
nand U23763 (N_23763,N_16407,N_18998);
nand U23764 (N_23764,N_17018,N_15158);
or U23765 (N_23765,N_15748,N_17155);
nor U23766 (N_23766,N_18283,N_17449);
nor U23767 (N_23767,N_18199,N_16356);
or U23768 (N_23768,N_19811,N_19859);
xnor U23769 (N_23769,N_15954,N_17265);
and U23770 (N_23770,N_17471,N_16840);
xnor U23771 (N_23771,N_18042,N_16815);
nand U23772 (N_23772,N_15850,N_19513);
nor U23773 (N_23773,N_16302,N_17867);
and U23774 (N_23774,N_19662,N_16274);
and U23775 (N_23775,N_19179,N_19178);
and U23776 (N_23776,N_17927,N_18273);
and U23777 (N_23777,N_19794,N_19025);
xnor U23778 (N_23778,N_16920,N_19971);
nand U23779 (N_23779,N_17050,N_19112);
xor U23780 (N_23780,N_15419,N_19600);
and U23781 (N_23781,N_16576,N_16046);
nor U23782 (N_23782,N_19588,N_16639);
nand U23783 (N_23783,N_15007,N_19895);
or U23784 (N_23784,N_17768,N_15527);
nor U23785 (N_23785,N_19689,N_17431);
and U23786 (N_23786,N_15046,N_19653);
nand U23787 (N_23787,N_16919,N_15889);
xor U23788 (N_23788,N_18350,N_18078);
nand U23789 (N_23789,N_15973,N_16027);
nor U23790 (N_23790,N_18048,N_16803);
nor U23791 (N_23791,N_17014,N_19002);
xnor U23792 (N_23792,N_19842,N_16491);
nand U23793 (N_23793,N_16593,N_15385);
nand U23794 (N_23794,N_17347,N_19896);
xor U23795 (N_23795,N_17754,N_19122);
and U23796 (N_23796,N_19062,N_16111);
or U23797 (N_23797,N_15543,N_17992);
nor U23798 (N_23798,N_17490,N_19971);
and U23799 (N_23799,N_16663,N_17378);
or U23800 (N_23800,N_15588,N_17363);
and U23801 (N_23801,N_16275,N_17597);
xor U23802 (N_23802,N_17642,N_16085);
nor U23803 (N_23803,N_18888,N_18719);
nand U23804 (N_23804,N_19261,N_19064);
and U23805 (N_23805,N_19810,N_16993);
nand U23806 (N_23806,N_18368,N_15034);
nand U23807 (N_23807,N_17832,N_17689);
or U23808 (N_23808,N_19890,N_16635);
xor U23809 (N_23809,N_17836,N_19245);
nor U23810 (N_23810,N_18917,N_15231);
nand U23811 (N_23811,N_16579,N_19550);
and U23812 (N_23812,N_15432,N_15592);
and U23813 (N_23813,N_16444,N_18298);
xnor U23814 (N_23814,N_18659,N_15681);
nor U23815 (N_23815,N_19894,N_15355);
or U23816 (N_23816,N_17627,N_15497);
or U23817 (N_23817,N_16898,N_19756);
or U23818 (N_23818,N_18240,N_15996);
and U23819 (N_23819,N_19773,N_18272);
nand U23820 (N_23820,N_19608,N_17787);
nor U23821 (N_23821,N_15168,N_18112);
or U23822 (N_23822,N_19086,N_19002);
xor U23823 (N_23823,N_15276,N_15951);
or U23824 (N_23824,N_17525,N_17297);
or U23825 (N_23825,N_19673,N_15292);
nand U23826 (N_23826,N_15253,N_16504);
or U23827 (N_23827,N_15452,N_18766);
xor U23828 (N_23828,N_18385,N_17647);
nand U23829 (N_23829,N_17588,N_17391);
and U23830 (N_23830,N_15958,N_18730);
nor U23831 (N_23831,N_18007,N_17541);
and U23832 (N_23832,N_16880,N_19101);
nand U23833 (N_23833,N_18385,N_18003);
or U23834 (N_23834,N_16369,N_18518);
or U23835 (N_23835,N_19171,N_15466);
nor U23836 (N_23836,N_16603,N_18157);
and U23837 (N_23837,N_16113,N_18480);
nor U23838 (N_23838,N_17034,N_18307);
nand U23839 (N_23839,N_15009,N_16097);
nor U23840 (N_23840,N_15300,N_18883);
xnor U23841 (N_23841,N_15466,N_15929);
or U23842 (N_23842,N_19362,N_18590);
and U23843 (N_23843,N_16882,N_16657);
xnor U23844 (N_23844,N_16804,N_19530);
nand U23845 (N_23845,N_17557,N_18450);
or U23846 (N_23846,N_15742,N_17168);
and U23847 (N_23847,N_19263,N_16784);
nand U23848 (N_23848,N_19980,N_17712);
and U23849 (N_23849,N_19676,N_17477);
nor U23850 (N_23850,N_15670,N_16374);
xor U23851 (N_23851,N_18827,N_19647);
xor U23852 (N_23852,N_17606,N_19908);
xor U23853 (N_23853,N_18057,N_18450);
xor U23854 (N_23854,N_18284,N_16141);
or U23855 (N_23855,N_18802,N_17333);
xor U23856 (N_23856,N_15359,N_15580);
and U23857 (N_23857,N_19323,N_19013);
nand U23858 (N_23858,N_18950,N_18423);
or U23859 (N_23859,N_17514,N_16855);
nand U23860 (N_23860,N_15748,N_17632);
and U23861 (N_23861,N_17235,N_16519);
xnor U23862 (N_23862,N_19529,N_16207);
nand U23863 (N_23863,N_19935,N_16014);
and U23864 (N_23864,N_19239,N_18230);
or U23865 (N_23865,N_15157,N_17030);
and U23866 (N_23866,N_19111,N_15133);
xnor U23867 (N_23867,N_16546,N_19975);
nand U23868 (N_23868,N_15589,N_18772);
nand U23869 (N_23869,N_17111,N_15111);
xnor U23870 (N_23870,N_18143,N_16560);
xor U23871 (N_23871,N_16495,N_17839);
and U23872 (N_23872,N_19730,N_19062);
xnor U23873 (N_23873,N_16482,N_15179);
and U23874 (N_23874,N_18573,N_16427);
xnor U23875 (N_23875,N_16052,N_18134);
and U23876 (N_23876,N_18215,N_19037);
and U23877 (N_23877,N_16822,N_17961);
or U23878 (N_23878,N_15760,N_18480);
nand U23879 (N_23879,N_17630,N_18544);
nor U23880 (N_23880,N_18560,N_15626);
nand U23881 (N_23881,N_16618,N_19821);
nand U23882 (N_23882,N_16589,N_16816);
or U23883 (N_23883,N_16354,N_18772);
nor U23884 (N_23884,N_18417,N_17846);
and U23885 (N_23885,N_17528,N_17036);
nand U23886 (N_23886,N_16517,N_16816);
and U23887 (N_23887,N_15878,N_15613);
and U23888 (N_23888,N_19899,N_15736);
nor U23889 (N_23889,N_19040,N_19344);
nand U23890 (N_23890,N_16533,N_16055);
nor U23891 (N_23891,N_18720,N_19404);
nand U23892 (N_23892,N_19192,N_17131);
xnor U23893 (N_23893,N_15364,N_19528);
and U23894 (N_23894,N_17093,N_17104);
nor U23895 (N_23895,N_18251,N_16227);
and U23896 (N_23896,N_17283,N_19577);
xor U23897 (N_23897,N_16051,N_15880);
and U23898 (N_23898,N_19274,N_17553);
xor U23899 (N_23899,N_18739,N_16482);
nor U23900 (N_23900,N_18817,N_17175);
nor U23901 (N_23901,N_18866,N_18196);
nor U23902 (N_23902,N_16400,N_16310);
or U23903 (N_23903,N_17056,N_19578);
nor U23904 (N_23904,N_17192,N_15730);
and U23905 (N_23905,N_19436,N_17477);
xor U23906 (N_23906,N_17573,N_17785);
xor U23907 (N_23907,N_15745,N_17644);
or U23908 (N_23908,N_16687,N_17581);
xor U23909 (N_23909,N_18516,N_17359);
nor U23910 (N_23910,N_17308,N_17722);
nand U23911 (N_23911,N_15777,N_15602);
and U23912 (N_23912,N_16591,N_15889);
or U23913 (N_23913,N_19989,N_17579);
nor U23914 (N_23914,N_17587,N_19896);
xnor U23915 (N_23915,N_16751,N_19487);
or U23916 (N_23916,N_19284,N_18757);
or U23917 (N_23917,N_19654,N_16565);
nor U23918 (N_23918,N_18564,N_17909);
nor U23919 (N_23919,N_19507,N_15546);
and U23920 (N_23920,N_17166,N_16791);
or U23921 (N_23921,N_18267,N_17897);
nor U23922 (N_23922,N_19597,N_18260);
or U23923 (N_23923,N_15878,N_15629);
nor U23924 (N_23924,N_19855,N_17531);
xor U23925 (N_23925,N_15599,N_15563);
nand U23926 (N_23926,N_17237,N_16144);
nand U23927 (N_23927,N_15181,N_15952);
nor U23928 (N_23928,N_15146,N_18376);
xnor U23929 (N_23929,N_18011,N_17394);
xnor U23930 (N_23930,N_15434,N_18189);
xor U23931 (N_23931,N_17435,N_18580);
nor U23932 (N_23932,N_19750,N_18433);
xor U23933 (N_23933,N_19254,N_19056);
nor U23934 (N_23934,N_19420,N_19914);
nor U23935 (N_23935,N_17364,N_16000);
or U23936 (N_23936,N_15602,N_19349);
xor U23937 (N_23937,N_19381,N_16399);
and U23938 (N_23938,N_18900,N_18306);
or U23939 (N_23939,N_15129,N_19718);
or U23940 (N_23940,N_19708,N_16744);
xnor U23941 (N_23941,N_19895,N_18869);
or U23942 (N_23942,N_17562,N_18663);
or U23943 (N_23943,N_15403,N_16275);
nand U23944 (N_23944,N_18782,N_18985);
or U23945 (N_23945,N_16132,N_18772);
and U23946 (N_23946,N_17330,N_16525);
xor U23947 (N_23947,N_15544,N_18987);
and U23948 (N_23948,N_15648,N_16780);
xnor U23949 (N_23949,N_17949,N_19239);
xor U23950 (N_23950,N_19780,N_16459);
nor U23951 (N_23951,N_16411,N_15184);
nor U23952 (N_23952,N_18430,N_16786);
and U23953 (N_23953,N_15190,N_17643);
nand U23954 (N_23954,N_17641,N_18339);
and U23955 (N_23955,N_15963,N_15133);
or U23956 (N_23956,N_19575,N_17922);
or U23957 (N_23957,N_17604,N_18295);
and U23958 (N_23958,N_18286,N_17926);
or U23959 (N_23959,N_17901,N_15361);
xor U23960 (N_23960,N_16133,N_15615);
and U23961 (N_23961,N_16340,N_16636);
nand U23962 (N_23962,N_18233,N_18197);
xnor U23963 (N_23963,N_16064,N_15416);
nand U23964 (N_23964,N_15346,N_16145);
and U23965 (N_23965,N_18943,N_18987);
and U23966 (N_23966,N_16795,N_16299);
xor U23967 (N_23967,N_18348,N_15795);
nand U23968 (N_23968,N_19547,N_16901);
or U23969 (N_23969,N_16547,N_19245);
nand U23970 (N_23970,N_15080,N_15407);
and U23971 (N_23971,N_16100,N_18786);
nor U23972 (N_23972,N_19311,N_15330);
nor U23973 (N_23973,N_16371,N_17968);
nor U23974 (N_23974,N_17153,N_19718);
xor U23975 (N_23975,N_15998,N_18457);
nor U23976 (N_23976,N_16643,N_19359);
nor U23977 (N_23977,N_16917,N_18037);
or U23978 (N_23978,N_17108,N_15858);
nand U23979 (N_23979,N_18340,N_16797);
xor U23980 (N_23980,N_16261,N_19014);
xnor U23981 (N_23981,N_15597,N_18347);
nand U23982 (N_23982,N_19527,N_15643);
nand U23983 (N_23983,N_16156,N_18984);
and U23984 (N_23984,N_16600,N_17150);
xnor U23985 (N_23985,N_17667,N_17952);
nor U23986 (N_23986,N_17421,N_15997);
xor U23987 (N_23987,N_18406,N_15183);
nand U23988 (N_23988,N_16153,N_18458);
xor U23989 (N_23989,N_16323,N_18591);
or U23990 (N_23990,N_18569,N_17469);
nor U23991 (N_23991,N_18991,N_16783);
nor U23992 (N_23992,N_19173,N_15547);
nand U23993 (N_23993,N_19214,N_18561);
and U23994 (N_23994,N_18483,N_19139);
nand U23995 (N_23995,N_16142,N_17919);
and U23996 (N_23996,N_18116,N_18205);
nor U23997 (N_23997,N_17918,N_16142);
or U23998 (N_23998,N_15428,N_15247);
and U23999 (N_23999,N_19159,N_19522);
or U24000 (N_24000,N_17079,N_16324);
or U24001 (N_24001,N_19409,N_16163);
xnor U24002 (N_24002,N_17145,N_16727);
nor U24003 (N_24003,N_19276,N_16694);
xor U24004 (N_24004,N_19885,N_15414);
and U24005 (N_24005,N_15677,N_15052);
or U24006 (N_24006,N_16968,N_15947);
xnor U24007 (N_24007,N_15391,N_15813);
xnor U24008 (N_24008,N_17951,N_16968);
nor U24009 (N_24009,N_18921,N_17372);
and U24010 (N_24010,N_19677,N_18947);
or U24011 (N_24011,N_18136,N_15933);
xor U24012 (N_24012,N_19214,N_17668);
xor U24013 (N_24013,N_17200,N_18770);
or U24014 (N_24014,N_18279,N_16844);
or U24015 (N_24015,N_16788,N_15070);
xor U24016 (N_24016,N_16477,N_16038);
or U24017 (N_24017,N_17359,N_18954);
or U24018 (N_24018,N_17480,N_18147);
or U24019 (N_24019,N_17932,N_15079);
and U24020 (N_24020,N_17143,N_17486);
nand U24021 (N_24021,N_15038,N_19668);
xor U24022 (N_24022,N_19717,N_19532);
nor U24023 (N_24023,N_19659,N_15420);
xnor U24024 (N_24024,N_17131,N_16455);
and U24025 (N_24025,N_19524,N_17247);
nand U24026 (N_24026,N_17635,N_18634);
or U24027 (N_24027,N_16489,N_17729);
or U24028 (N_24028,N_17824,N_15387);
nand U24029 (N_24029,N_18384,N_19864);
xnor U24030 (N_24030,N_17300,N_16372);
xnor U24031 (N_24031,N_15937,N_15135);
nor U24032 (N_24032,N_15358,N_15162);
and U24033 (N_24033,N_15457,N_16540);
nor U24034 (N_24034,N_15683,N_15014);
nand U24035 (N_24035,N_18048,N_17624);
nand U24036 (N_24036,N_18327,N_19082);
and U24037 (N_24037,N_15444,N_15198);
and U24038 (N_24038,N_15782,N_19122);
and U24039 (N_24039,N_16828,N_19327);
or U24040 (N_24040,N_15899,N_18755);
nand U24041 (N_24041,N_17046,N_17708);
nor U24042 (N_24042,N_19597,N_19681);
and U24043 (N_24043,N_19025,N_17634);
xnor U24044 (N_24044,N_18589,N_18249);
or U24045 (N_24045,N_19569,N_16203);
nor U24046 (N_24046,N_16607,N_19332);
and U24047 (N_24047,N_15297,N_17863);
or U24048 (N_24048,N_15464,N_19537);
or U24049 (N_24049,N_17605,N_18756);
nor U24050 (N_24050,N_17748,N_17889);
and U24051 (N_24051,N_18822,N_18942);
or U24052 (N_24052,N_16302,N_15787);
xnor U24053 (N_24053,N_18609,N_15281);
and U24054 (N_24054,N_16101,N_18249);
xnor U24055 (N_24055,N_17724,N_15536);
and U24056 (N_24056,N_15705,N_15606);
nand U24057 (N_24057,N_18960,N_16412);
or U24058 (N_24058,N_18380,N_19190);
nor U24059 (N_24059,N_16448,N_19197);
xnor U24060 (N_24060,N_19291,N_19898);
or U24061 (N_24061,N_19417,N_16770);
xor U24062 (N_24062,N_15448,N_16931);
xnor U24063 (N_24063,N_18989,N_15804);
nand U24064 (N_24064,N_15072,N_19716);
nor U24065 (N_24065,N_15779,N_16223);
nand U24066 (N_24066,N_16194,N_15285);
and U24067 (N_24067,N_16673,N_16889);
nand U24068 (N_24068,N_19903,N_17130);
nor U24069 (N_24069,N_16366,N_19754);
nor U24070 (N_24070,N_17278,N_18358);
nor U24071 (N_24071,N_18927,N_19913);
nor U24072 (N_24072,N_19773,N_15318);
or U24073 (N_24073,N_18468,N_17212);
xnor U24074 (N_24074,N_18724,N_15345);
nand U24075 (N_24075,N_16414,N_15126);
or U24076 (N_24076,N_16831,N_18399);
and U24077 (N_24077,N_15543,N_18838);
nand U24078 (N_24078,N_17723,N_15541);
nand U24079 (N_24079,N_16085,N_17492);
xor U24080 (N_24080,N_19757,N_17047);
nand U24081 (N_24081,N_19004,N_18388);
or U24082 (N_24082,N_17343,N_15231);
or U24083 (N_24083,N_16318,N_19454);
nand U24084 (N_24084,N_19037,N_18714);
or U24085 (N_24085,N_15283,N_15859);
nor U24086 (N_24086,N_18796,N_19772);
or U24087 (N_24087,N_19929,N_16266);
xnor U24088 (N_24088,N_15046,N_16893);
or U24089 (N_24089,N_18300,N_15295);
or U24090 (N_24090,N_15414,N_16514);
or U24091 (N_24091,N_17136,N_15681);
xnor U24092 (N_24092,N_16156,N_17519);
or U24093 (N_24093,N_16471,N_18302);
nand U24094 (N_24094,N_17779,N_15337);
xor U24095 (N_24095,N_15151,N_16945);
or U24096 (N_24096,N_15961,N_16285);
xnor U24097 (N_24097,N_16512,N_19913);
or U24098 (N_24098,N_15926,N_19703);
nor U24099 (N_24099,N_18636,N_18635);
xnor U24100 (N_24100,N_17649,N_15145);
and U24101 (N_24101,N_15289,N_19952);
and U24102 (N_24102,N_17291,N_18358);
nand U24103 (N_24103,N_15397,N_19479);
nand U24104 (N_24104,N_15508,N_17123);
xnor U24105 (N_24105,N_17125,N_16928);
xnor U24106 (N_24106,N_18060,N_18961);
xor U24107 (N_24107,N_16130,N_18871);
and U24108 (N_24108,N_18765,N_16963);
and U24109 (N_24109,N_19346,N_15903);
or U24110 (N_24110,N_16877,N_15367);
nor U24111 (N_24111,N_17844,N_18601);
or U24112 (N_24112,N_19741,N_17691);
nand U24113 (N_24113,N_15982,N_17457);
xnor U24114 (N_24114,N_18154,N_15354);
nand U24115 (N_24115,N_18718,N_17302);
nand U24116 (N_24116,N_16786,N_19387);
xnor U24117 (N_24117,N_17097,N_18082);
xor U24118 (N_24118,N_18895,N_16806);
nor U24119 (N_24119,N_15378,N_18834);
nand U24120 (N_24120,N_19126,N_16001);
nor U24121 (N_24121,N_17041,N_16400);
and U24122 (N_24122,N_15236,N_15331);
or U24123 (N_24123,N_15908,N_19038);
nor U24124 (N_24124,N_16874,N_17178);
xnor U24125 (N_24125,N_19521,N_19704);
and U24126 (N_24126,N_18234,N_19217);
and U24127 (N_24127,N_15240,N_16454);
and U24128 (N_24128,N_16600,N_16164);
xor U24129 (N_24129,N_17229,N_16166);
nand U24130 (N_24130,N_19668,N_16802);
xor U24131 (N_24131,N_19598,N_16504);
nor U24132 (N_24132,N_15480,N_18491);
nand U24133 (N_24133,N_19081,N_16290);
xnor U24134 (N_24134,N_19397,N_15262);
nor U24135 (N_24135,N_17888,N_16602);
nor U24136 (N_24136,N_15023,N_15297);
nor U24137 (N_24137,N_18842,N_18134);
nand U24138 (N_24138,N_15424,N_18683);
nand U24139 (N_24139,N_16259,N_19021);
and U24140 (N_24140,N_17292,N_17523);
xor U24141 (N_24141,N_19370,N_19901);
nor U24142 (N_24142,N_18032,N_17829);
xnor U24143 (N_24143,N_15631,N_17015);
or U24144 (N_24144,N_19063,N_19956);
nor U24145 (N_24145,N_16785,N_15087);
nor U24146 (N_24146,N_15260,N_15812);
xnor U24147 (N_24147,N_16124,N_18207);
and U24148 (N_24148,N_17341,N_17712);
xnor U24149 (N_24149,N_19564,N_18090);
nand U24150 (N_24150,N_18658,N_15297);
nand U24151 (N_24151,N_18399,N_18470);
nand U24152 (N_24152,N_19949,N_15311);
xor U24153 (N_24153,N_19054,N_18577);
and U24154 (N_24154,N_19779,N_17946);
nand U24155 (N_24155,N_19800,N_19098);
xnor U24156 (N_24156,N_19053,N_18741);
and U24157 (N_24157,N_18635,N_17892);
and U24158 (N_24158,N_17088,N_19621);
and U24159 (N_24159,N_15322,N_16111);
or U24160 (N_24160,N_18572,N_18604);
or U24161 (N_24161,N_19343,N_18115);
nor U24162 (N_24162,N_18947,N_19719);
and U24163 (N_24163,N_17742,N_18254);
xor U24164 (N_24164,N_15139,N_19147);
and U24165 (N_24165,N_18866,N_19616);
nor U24166 (N_24166,N_16136,N_15241);
xnor U24167 (N_24167,N_17534,N_16647);
xnor U24168 (N_24168,N_15086,N_16264);
or U24169 (N_24169,N_15323,N_19212);
xor U24170 (N_24170,N_19362,N_16949);
xor U24171 (N_24171,N_17494,N_19389);
xor U24172 (N_24172,N_15099,N_16864);
nand U24173 (N_24173,N_16549,N_18394);
or U24174 (N_24174,N_15492,N_17890);
nor U24175 (N_24175,N_17204,N_19649);
or U24176 (N_24176,N_19236,N_17560);
xor U24177 (N_24177,N_19429,N_19343);
xnor U24178 (N_24178,N_17655,N_19214);
and U24179 (N_24179,N_19786,N_17070);
and U24180 (N_24180,N_19429,N_15129);
or U24181 (N_24181,N_16549,N_16740);
and U24182 (N_24182,N_17439,N_18655);
nor U24183 (N_24183,N_19621,N_17039);
or U24184 (N_24184,N_17499,N_19020);
xor U24185 (N_24185,N_18887,N_15771);
or U24186 (N_24186,N_16042,N_18760);
and U24187 (N_24187,N_16674,N_17892);
nor U24188 (N_24188,N_19099,N_19207);
xor U24189 (N_24189,N_19685,N_19244);
nor U24190 (N_24190,N_18485,N_18589);
xnor U24191 (N_24191,N_17941,N_16810);
xor U24192 (N_24192,N_19508,N_19702);
and U24193 (N_24193,N_15488,N_19208);
xor U24194 (N_24194,N_17394,N_19125);
nor U24195 (N_24195,N_16092,N_16525);
nor U24196 (N_24196,N_19065,N_19471);
nor U24197 (N_24197,N_17269,N_17472);
and U24198 (N_24198,N_18479,N_18615);
and U24199 (N_24199,N_16687,N_19600);
xor U24200 (N_24200,N_16535,N_19767);
nand U24201 (N_24201,N_16175,N_15320);
nand U24202 (N_24202,N_17178,N_19498);
nor U24203 (N_24203,N_18981,N_19496);
nand U24204 (N_24204,N_19802,N_17545);
and U24205 (N_24205,N_17490,N_19599);
and U24206 (N_24206,N_16922,N_15286);
nand U24207 (N_24207,N_17863,N_17566);
nor U24208 (N_24208,N_15283,N_16038);
nand U24209 (N_24209,N_18264,N_17885);
nand U24210 (N_24210,N_17466,N_17023);
xnor U24211 (N_24211,N_17211,N_18923);
xnor U24212 (N_24212,N_16941,N_18490);
xnor U24213 (N_24213,N_16950,N_19752);
nor U24214 (N_24214,N_18486,N_18596);
nor U24215 (N_24215,N_18928,N_19230);
xor U24216 (N_24216,N_18169,N_19715);
and U24217 (N_24217,N_18605,N_19541);
nor U24218 (N_24218,N_15622,N_15879);
nand U24219 (N_24219,N_19069,N_15236);
and U24220 (N_24220,N_16304,N_19712);
or U24221 (N_24221,N_19732,N_15283);
and U24222 (N_24222,N_18450,N_19235);
xor U24223 (N_24223,N_19209,N_15285);
nand U24224 (N_24224,N_17699,N_18201);
or U24225 (N_24225,N_15557,N_16173);
or U24226 (N_24226,N_17672,N_15771);
nor U24227 (N_24227,N_15690,N_19183);
nand U24228 (N_24228,N_16174,N_15063);
xnor U24229 (N_24229,N_19070,N_18726);
nor U24230 (N_24230,N_15335,N_17440);
or U24231 (N_24231,N_16617,N_15549);
nor U24232 (N_24232,N_19266,N_18354);
nand U24233 (N_24233,N_16753,N_16674);
nor U24234 (N_24234,N_17181,N_15403);
and U24235 (N_24235,N_15696,N_18845);
nand U24236 (N_24236,N_15544,N_15206);
or U24237 (N_24237,N_15383,N_16598);
nor U24238 (N_24238,N_19928,N_18650);
xor U24239 (N_24239,N_17786,N_16259);
or U24240 (N_24240,N_17985,N_15248);
nor U24241 (N_24241,N_19823,N_19004);
or U24242 (N_24242,N_18281,N_19370);
xor U24243 (N_24243,N_15958,N_18481);
nand U24244 (N_24244,N_18184,N_16994);
xor U24245 (N_24245,N_19241,N_17017);
nand U24246 (N_24246,N_16551,N_16249);
nand U24247 (N_24247,N_15970,N_19255);
nor U24248 (N_24248,N_17507,N_19024);
xor U24249 (N_24249,N_18707,N_18066);
xor U24250 (N_24250,N_16953,N_19490);
xnor U24251 (N_24251,N_15580,N_16562);
xnor U24252 (N_24252,N_16820,N_15549);
xnor U24253 (N_24253,N_16650,N_16257);
nor U24254 (N_24254,N_17227,N_15085);
and U24255 (N_24255,N_19675,N_16895);
nor U24256 (N_24256,N_16245,N_18027);
and U24257 (N_24257,N_15348,N_16751);
xnor U24258 (N_24258,N_18996,N_15446);
nor U24259 (N_24259,N_17666,N_17446);
nor U24260 (N_24260,N_18133,N_18061);
and U24261 (N_24261,N_18015,N_15660);
nor U24262 (N_24262,N_17596,N_19466);
nor U24263 (N_24263,N_18309,N_17527);
nor U24264 (N_24264,N_15715,N_16557);
nand U24265 (N_24265,N_17249,N_17737);
or U24266 (N_24266,N_16437,N_15766);
or U24267 (N_24267,N_19033,N_16983);
xnor U24268 (N_24268,N_19758,N_18635);
and U24269 (N_24269,N_16744,N_19936);
nor U24270 (N_24270,N_18448,N_16930);
xor U24271 (N_24271,N_15360,N_17593);
nor U24272 (N_24272,N_18841,N_15258);
nand U24273 (N_24273,N_17371,N_19625);
xnor U24274 (N_24274,N_17352,N_16143);
xnor U24275 (N_24275,N_19883,N_17031);
xor U24276 (N_24276,N_17656,N_15362);
nor U24277 (N_24277,N_16501,N_15279);
and U24278 (N_24278,N_17981,N_16561);
nor U24279 (N_24279,N_19331,N_17029);
xnor U24280 (N_24280,N_19238,N_16872);
and U24281 (N_24281,N_17388,N_19564);
xnor U24282 (N_24282,N_16503,N_17703);
nand U24283 (N_24283,N_19584,N_16131);
nand U24284 (N_24284,N_18560,N_19743);
and U24285 (N_24285,N_16240,N_16523);
and U24286 (N_24286,N_19016,N_16403);
nand U24287 (N_24287,N_15669,N_16457);
xor U24288 (N_24288,N_18461,N_19988);
or U24289 (N_24289,N_15422,N_18705);
or U24290 (N_24290,N_15001,N_15286);
and U24291 (N_24291,N_17199,N_19611);
nor U24292 (N_24292,N_19153,N_15207);
and U24293 (N_24293,N_19480,N_17146);
or U24294 (N_24294,N_15293,N_19968);
or U24295 (N_24295,N_17608,N_19711);
or U24296 (N_24296,N_18139,N_16438);
and U24297 (N_24297,N_19002,N_18134);
nand U24298 (N_24298,N_18517,N_19750);
xnor U24299 (N_24299,N_17849,N_18578);
and U24300 (N_24300,N_17754,N_17573);
or U24301 (N_24301,N_15044,N_15753);
xor U24302 (N_24302,N_19351,N_15893);
nor U24303 (N_24303,N_17932,N_16400);
nand U24304 (N_24304,N_15115,N_19506);
nand U24305 (N_24305,N_16060,N_18664);
nor U24306 (N_24306,N_17343,N_16769);
nor U24307 (N_24307,N_18226,N_17406);
or U24308 (N_24308,N_18547,N_18027);
xor U24309 (N_24309,N_17831,N_19669);
or U24310 (N_24310,N_19248,N_16175);
nand U24311 (N_24311,N_15641,N_18337);
xnor U24312 (N_24312,N_19293,N_15293);
xor U24313 (N_24313,N_17719,N_16214);
xnor U24314 (N_24314,N_16359,N_17444);
and U24315 (N_24315,N_16374,N_17431);
and U24316 (N_24316,N_17337,N_19859);
xor U24317 (N_24317,N_16106,N_15728);
nor U24318 (N_24318,N_19773,N_18936);
nor U24319 (N_24319,N_16833,N_19133);
nand U24320 (N_24320,N_17307,N_17686);
or U24321 (N_24321,N_17996,N_18445);
nand U24322 (N_24322,N_16169,N_16375);
nor U24323 (N_24323,N_19168,N_15892);
nor U24324 (N_24324,N_15964,N_15632);
xor U24325 (N_24325,N_19198,N_19577);
nor U24326 (N_24326,N_15975,N_17152);
or U24327 (N_24327,N_18215,N_15614);
xnor U24328 (N_24328,N_17059,N_16739);
nor U24329 (N_24329,N_18496,N_16109);
nor U24330 (N_24330,N_17592,N_18791);
xor U24331 (N_24331,N_16150,N_16238);
xnor U24332 (N_24332,N_17987,N_18594);
xnor U24333 (N_24333,N_19100,N_19968);
nor U24334 (N_24334,N_17577,N_16453);
or U24335 (N_24335,N_18343,N_19753);
and U24336 (N_24336,N_18831,N_19561);
or U24337 (N_24337,N_16116,N_15427);
and U24338 (N_24338,N_18338,N_19006);
xor U24339 (N_24339,N_16833,N_17042);
and U24340 (N_24340,N_18312,N_15979);
or U24341 (N_24341,N_17437,N_15057);
and U24342 (N_24342,N_18845,N_17807);
nand U24343 (N_24343,N_16219,N_15989);
and U24344 (N_24344,N_18131,N_19121);
nand U24345 (N_24345,N_15047,N_17134);
nor U24346 (N_24346,N_19099,N_15707);
or U24347 (N_24347,N_16071,N_16048);
or U24348 (N_24348,N_16510,N_15295);
nor U24349 (N_24349,N_16898,N_19664);
nand U24350 (N_24350,N_16177,N_19832);
or U24351 (N_24351,N_15932,N_15555);
xnor U24352 (N_24352,N_15661,N_19518);
nand U24353 (N_24353,N_16046,N_17857);
and U24354 (N_24354,N_18449,N_16817);
or U24355 (N_24355,N_18355,N_17617);
or U24356 (N_24356,N_16175,N_19991);
or U24357 (N_24357,N_15930,N_19107);
nor U24358 (N_24358,N_15227,N_17774);
xor U24359 (N_24359,N_17473,N_17694);
or U24360 (N_24360,N_15111,N_19868);
or U24361 (N_24361,N_19527,N_19560);
and U24362 (N_24362,N_15520,N_19015);
xor U24363 (N_24363,N_16724,N_17103);
xnor U24364 (N_24364,N_15090,N_19538);
nor U24365 (N_24365,N_18376,N_19384);
nor U24366 (N_24366,N_15250,N_18893);
nand U24367 (N_24367,N_18579,N_17486);
or U24368 (N_24368,N_18393,N_17318);
nand U24369 (N_24369,N_19967,N_15277);
xor U24370 (N_24370,N_15989,N_19789);
or U24371 (N_24371,N_18202,N_16972);
nand U24372 (N_24372,N_18447,N_18816);
and U24373 (N_24373,N_16082,N_15950);
nor U24374 (N_24374,N_18946,N_17744);
nand U24375 (N_24375,N_17494,N_18638);
or U24376 (N_24376,N_18469,N_15146);
nand U24377 (N_24377,N_16489,N_15707);
and U24378 (N_24378,N_17076,N_17278);
and U24379 (N_24379,N_16394,N_15500);
and U24380 (N_24380,N_18701,N_17933);
nor U24381 (N_24381,N_19533,N_19968);
and U24382 (N_24382,N_17166,N_15883);
and U24383 (N_24383,N_16034,N_16690);
and U24384 (N_24384,N_15004,N_15993);
and U24385 (N_24385,N_16873,N_18677);
nand U24386 (N_24386,N_16971,N_18502);
nand U24387 (N_24387,N_18869,N_17165);
xor U24388 (N_24388,N_18337,N_15293);
nand U24389 (N_24389,N_18281,N_19513);
xor U24390 (N_24390,N_19034,N_18982);
nor U24391 (N_24391,N_16199,N_15500);
or U24392 (N_24392,N_16866,N_15811);
nand U24393 (N_24393,N_16940,N_15219);
and U24394 (N_24394,N_15773,N_16297);
nand U24395 (N_24395,N_18635,N_19946);
xor U24396 (N_24396,N_19335,N_17842);
nor U24397 (N_24397,N_17027,N_15605);
nor U24398 (N_24398,N_15276,N_16520);
nand U24399 (N_24399,N_19296,N_19484);
or U24400 (N_24400,N_18114,N_17841);
nand U24401 (N_24401,N_16663,N_16608);
nand U24402 (N_24402,N_16888,N_18087);
and U24403 (N_24403,N_15200,N_19287);
and U24404 (N_24404,N_18580,N_16405);
xor U24405 (N_24405,N_17709,N_15794);
or U24406 (N_24406,N_17029,N_18447);
or U24407 (N_24407,N_19356,N_18474);
xnor U24408 (N_24408,N_17567,N_17281);
and U24409 (N_24409,N_18077,N_16353);
or U24410 (N_24410,N_15991,N_16156);
nand U24411 (N_24411,N_15393,N_15503);
nor U24412 (N_24412,N_19634,N_19172);
nor U24413 (N_24413,N_19087,N_15640);
xor U24414 (N_24414,N_16605,N_19901);
and U24415 (N_24415,N_17992,N_15128);
xnor U24416 (N_24416,N_19643,N_17676);
or U24417 (N_24417,N_16785,N_18036);
nand U24418 (N_24418,N_15058,N_15156);
xnor U24419 (N_24419,N_15949,N_16182);
nand U24420 (N_24420,N_16721,N_15493);
nor U24421 (N_24421,N_18408,N_15414);
nand U24422 (N_24422,N_15174,N_19844);
xor U24423 (N_24423,N_18753,N_16218);
or U24424 (N_24424,N_16651,N_18133);
and U24425 (N_24425,N_17903,N_18044);
nor U24426 (N_24426,N_16620,N_18942);
nand U24427 (N_24427,N_16446,N_19658);
nand U24428 (N_24428,N_15400,N_17860);
xnor U24429 (N_24429,N_17159,N_15412);
nand U24430 (N_24430,N_18081,N_19006);
xnor U24431 (N_24431,N_19546,N_18930);
xor U24432 (N_24432,N_17367,N_18945);
nand U24433 (N_24433,N_16345,N_16737);
nor U24434 (N_24434,N_18694,N_16174);
xnor U24435 (N_24435,N_19129,N_19580);
and U24436 (N_24436,N_17660,N_17176);
nand U24437 (N_24437,N_18075,N_18797);
nand U24438 (N_24438,N_15962,N_16916);
nor U24439 (N_24439,N_16722,N_16940);
nor U24440 (N_24440,N_15239,N_18404);
nand U24441 (N_24441,N_16268,N_15789);
nand U24442 (N_24442,N_17787,N_19440);
nand U24443 (N_24443,N_15156,N_15446);
and U24444 (N_24444,N_17955,N_15168);
or U24445 (N_24445,N_17723,N_15444);
xnor U24446 (N_24446,N_18906,N_16935);
and U24447 (N_24447,N_16512,N_19689);
nor U24448 (N_24448,N_18568,N_19481);
and U24449 (N_24449,N_19659,N_17598);
xnor U24450 (N_24450,N_19751,N_17870);
nor U24451 (N_24451,N_19070,N_16399);
xnor U24452 (N_24452,N_18606,N_19800);
and U24453 (N_24453,N_16494,N_19841);
or U24454 (N_24454,N_15204,N_18269);
nand U24455 (N_24455,N_19436,N_17355);
nor U24456 (N_24456,N_16432,N_16586);
xnor U24457 (N_24457,N_15047,N_17576);
xnor U24458 (N_24458,N_16724,N_18037);
or U24459 (N_24459,N_16769,N_18588);
and U24460 (N_24460,N_15690,N_16954);
xor U24461 (N_24461,N_17037,N_16557);
or U24462 (N_24462,N_17551,N_19904);
nand U24463 (N_24463,N_17452,N_15701);
or U24464 (N_24464,N_16684,N_18685);
xnor U24465 (N_24465,N_18846,N_18121);
nand U24466 (N_24466,N_17803,N_17334);
or U24467 (N_24467,N_15582,N_16576);
xor U24468 (N_24468,N_15313,N_19650);
xor U24469 (N_24469,N_17634,N_15009);
xor U24470 (N_24470,N_16942,N_15136);
nand U24471 (N_24471,N_16388,N_18412);
nor U24472 (N_24472,N_19507,N_15636);
nor U24473 (N_24473,N_18178,N_18881);
and U24474 (N_24474,N_19315,N_19350);
nand U24475 (N_24475,N_15945,N_18735);
xnor U24476 (N_24476,N_17472,N_19942);
xnor U24477 (N_24477,N_18691,N_16212);
nor U24478 (N_24478,N_17442,N_16394);
and U24479 (N_24479,N_18963,N_17991);
xor U24480 (N_24480,N_15818,N_16124);
nand U24481 (N_24481,N_15698,N_15646);
xnor U24482 (N_24482,N_18502,N_17932);
nand U24483 (N_24483,N_16760,N_17254);
nand U24484 (N_24484,N_16447,N_18106);
or U24485 (N_24485,N_16166,N_19567);
xor U24486 (N_24486,N_17854,N_18383);
nor U24487 (N_24487,N_18037,N_19571);
or U24488 (N_24488,N_15990,N_18884);
and U24489 (N_24489,N_17517,N_17295);
and U24490 (N_24490,N_18911,N_18947);
and U24491 (N_24491,N_18571,N_19466);
and U24492 (N_24492,N_17765,N_16937);
nand U24493 (N_24493,N_18086,N_19058);
nor U24494 (N_24494,N_18659,N_16077);
xor U24495 (N_24495,N_15125,N_15384);
nand U24496 (N_24496,N_18056,N_19275);
xor U24497 (N_24497,N_15929,N_18777);
nand U24498 (N_24498,N_18467,N_15463);
and U24499 (N_24499,N_18207,N_19228);
or U24500 (N_24500,N_15414,N_15762);
xnor U24501 (N_24501,N_17025,N_17503);
xor U24502 (N_24502,N_16486,N_18689);
nand U24503 (N_24503,N_17882,N_16550);
nor U24504 (N_24504,N_15309,N_16960);
and U24505 (N_24505,N_17584,N_17190);
or U24506 (N_24506,N_19026,N_15044);
xnor U24507 (N_24507,N_17579,N_15301);
nand U24508 (N_24508,N_16171,N_17581);
and U24509 (N_24509,N_18831,N_18935);
nor U24510 (N_24510,N_19665,N_19906);
xnor U24511 (N_24511,N_15544,N_16433);
nand U24512 (N_24512,N_18444,N_19164);
and U24513 (N_24513,N_18459,N_18886);
nand U24514 (N_24514,N_16299,N_15256);
and U24515 (N_24515,N_19201,N_18907);
nand U24516 (N_24516,N_15066,N_17157);
nand U24517 (N_24517,N_15067,N_15464);
nand U24518 (N_24518,N_19255,N_15881);
nand U24519 (N_24519,N_19364,N_15790);
nor U24520 (N_24520,N_15254,N_15200);
and U24521 (N_24521,N_15524,N_18117);
nor U24522 (N_24522,N_15959,N_16297);
nor U24523 (N_24523,N_19319,N_19125);
xnor U24524 (N_24524,N_17707,N_17538);
nor U24525 (N_24525,N_19913,N_16594);
or U24526 (N_24526,N_16811,N_17703);
or U24527 (N_24527,N_19871,N_16123);
or U24528 (N_24528,N_19230,N_16710);
xor U24529 (N_24529,N_19029,N_15269);
or U24530 (N_24530,N_18688,N_16548);
or U24531 (N_24531,N_18026,N_16698);
nand U24532 (N_24532,N_18544,N_15160);
nor U24533 (N_24533,N_17095,N_16283);
xnor U24534 (N_24534,N_16573,N_15794);
nor U24535 (N_24535,N_18131,N_18551);
nand U24536 (N_24536,N_18939,N_16135);
nor U24537 (N_24537,N_17378,N_19000);
or U24538 (N_24538,N_19189,N_18956);
and U24539 (N_24539,N_18280,N_19608);
or U24540 (N_24540,N_17391,N_17811);
nor U24541 (N_24541,N_16319,N_15888);
and U24542 (N_24542,N_19157,N_18459);
xor U24543 (N_24543,N_15630,N_18781);
nor U24544 (N_24544,N_18290,N_18421);
or U24545 (N_24545,N_19698,N_19934);
and U24546 (N_24546,N_17123,N_15013);
or U24547 (N_24547,N_15497,N_15457);
nor U24548 (N_24548,N_18270,N_17717);
or U24549 (N_24549,N_16178,N_17253);
nand U24550 (N_24550,N_17285,N_16134);
nand U24551 (N_24551,N_18512,N_15470);
nand U24552 (N_24552,N_15816,N_17048);
nor U24553 (N_24553,N_17824,N_15634);
or U24554 (N_24554,N_17115,N_18141);
nand U24555 (N_24555,N_19705,N_17855);
or U24556 (N_24556,N_15103,N_16523);
and U24557 (N_24557,N_19254,N_19711);
xnor U24558 (N_24558,N_17860,N_15809);
or U24559 (N_24559,N_17444,N_18376);
nor U24560 (N_24560,N_19608,N_18041);
xor U24561 (N_24561,N_19188,N_16534);
and U24562 (N_24562,N_17166,N_18234);
nor U24563 (N_24563,N_18508,N_17244);
nor U24564 (N_24564,N_16441,N_18589);
and U24565 (N_24565,N_18351,N_19099);
xor U24566 (N_24566,N_19172,N_15973);
xor U24567 (N_24567,N_17339,N_18600);
nor U24568 (N_24568,N_17455,N_18223);
xor U24569 (N_24569,N_17333,N_17187);
xnor U24570 (N_24570,N_18088,N_19776);
nor U24571 (N_24571,N_16463,N_16544);
nand U24572 (N_24572,N_16324,N_18041);
and U24573 (N_24573,N_17587,N_17582);
nand U24574 (N_24574,N_18851,N_18469);
nor U24575 (N_24575,N_16132,N_17179);
nand U24576 (N_24576,N_19817,N_15750);
nor U24577 (N_24577,N_17747,N_18112);
nand U24578 (N_24578,N_19238,N_19771);
or U24579 (N_24579,N_17612,N_15331);
nor U24580 (N_24580,N_16809,N_19328);
nand U24581 (N_24581,N_19646,N_18501);
or U24582 (N_24582,N_16662,N_15796);
or U24583 (N_24583,N_15143,N_15139);
nand U24584 (N_24584,N_16458,N_17199);
and U24585 (N_24585,N_17534,N_16497);
and U24586 (N_24586,N_16722,N_16782);
or U24587 (N_24587,N_17532,N_19256);
nor U24588 (N_24588,N_17402,N_19652);
nand U24589 (N_24589,N_19998,N_15998);
xnor U24590 (N_24590,N_19213,N_15109);
nor U24591 (N_24591,N_17799,N_19606);
or U24592 (N_24592,N_15664,N_16681);
or U24593 (N_24593,N_18382,N_16321);
and U24594 (N_24594,N_18223,N_16633);
nor U24595 (N_24595,N_18505,N_17503);
and U24596 (N_24596,N_15400,N_19846);
or U24597 (N_24597,N_17941,N_17904);
or U24598 (N_24598,N_19667,N_18611);
and U24599 (N_24599,N_16586,N_15629);
and U24600 (N_24600,N_15746,N_16288);
and U24601 (N_24601,N_15498,N_18959);
nand U24602 (N_24602,N_19394,N_15483);
xnor U24603 (N_24603,N_15162,N_19307);
and U24604 (N_24604,N_16035,N_18055);
nand U24605 (N_24605,N_15409,N_15586);
or U24606 (N_24606,N_15686,N_15697);
nor U24607 (N_24607,N_18617,N_19082);
and U24608 (N_24608,N_16305,N_17006);
and U24609 (N_24609,N_18387,N_15652);
nor U24610 (N_24610,N_17708,N_19724);
and U24611 (N_24611,N_15155,N_16214);
nand U24612 (N_24612,N_19373,N_18094);
and U24613 (N_24613,N_18172,N_15270);
nor U24614 (N_24614,N_16681,N_15174);
or U24615 (N_24615,N_18850,N_16282);
xor U24616 (N_24616,N_16318,N_19096);
nand U24617 (N_24617,N_15745,N_17508);
nand U24618 (N_24618,N_16603,N_15127);
or U24619 (N_24619,N_17092,N_18532);
xor U24620 (N_24620,N_19897,N_18147);
nor U24621 (N_24621,N_18332,N_15943);
nand U24622 (N_24622,N_19507,N_19098);
nand U24623 (N_24623,N_15865,N_16038);
and U24624 (N_24624,N_18259,N_15183);
nand U24625 (N_24625,N_16634,N_18943);
nor U24626 (N_24626,N_17645,N_19203);
nor U24627 (N_24627,N_18473,N_19120);
or U24628 (N_24628,N_17831,N_18432);
nor U24629 (N_24629,N_18966,N_16439);
xnor U24630 (N_24630,N_17016,N_19899);
nor U24631 (N_24631,N_15377,N_15858);
or U24632 (N_24632,N_19044,N_17893);
and U24633 (N_24633,N_17272,N_18283);
or U24634 (N_24634,N_18626,N_16505);
xor U24635 (N_24635,N_19498,N_18570);
xnor U24636 (N_24636,N_18213,N_15029);
nor U24637 (N_24637,N_19616,N_19786);
xnor U24638 (N_24638,N_17898,N_19018);
and U24639 (N_24639,N_19298,N_19378);
xnor U24640 (N_24640,N_19764,N_19871);
and U24641 (N_24641,N_18284,N_17958);
nand U24642 (N_24642,N_19767,N_16081);
nor U24643 (N_24643,N_15290,N_15650);
nand U24644 (N_24644,N_15764,N_15765);
nand U24645 (N_24645,N_15655,N_17305);
xor U24646 (N_24646,N_19440,N_15296);
nor U24647 (N_24647,N_16059,N_17273);
and U24648 (N_24648,N_16388,N_19152);
and U24649 (N_24649,N_15675,N_17226);
or U24650 (N_24650,N_16912,N_15943);
or U24651 (N_24651,N_16353,N_16175);
or U24652 (N_24652,N_19521,N_17638);
nand U24653 (N_24653,N_19047,N_17735);
xnor U24654 (N_24654,N_16199,N_16303);
nand U24655 (N_24655,N_18598,N_16145);
and U24656 (N_24656,N_15771,N_15809);
xnor U24657 (N_24657,N_15088,N_17482);
nand U24658 (N_24658,N_18622,N_19147);
nand U24659 (N_24659,N_15995,N_17243);
nand U24660 (N_24660,N_18094,N_18770);
nor U24661 (N_24661,N_17936,N_16592);
nand U24662 (N_24662,N_18549,N_18377);
or U24663 (N_24663,N_17751,N_19196);
or U24664 (N_24664,N_19468,N_17440);
and U24665 (N_24665,N_17375,N_19487);
and U24666 (N_24666,N_18196,N_17507);
nand U24667 (N_24667,N_17562,N_16314);
or U24668 (N_24668,N_15271,N_16757);
xnor U24669 (N_24669,N_19747,N_18057);
nor U24670 (N_24670,N_17161,N_16122);
xor U24671 (N_24671,N_16306,N_19492);
nand U24672 (N_24672,N_15199,N_15183);
and U24673 (N_24673,N_18777,N_16051);
xor U24674 (N_24674,N_19767,N_17293);
xnor U24675 (N_24675,N_15104,N_15731);
and U24676 (N_24676,N_17015,N_18946);
xnor U24677 (N_24677,N_15949,N_16761);
and U24678 (N_24678,N_17877,N_16042);
xnor U24679 (N_24679,N_18873,N_16075);
nand U24680 (N_24680,N_15224,N_17836);
nand U24681 (N_24681,N_18849,N_18466);
nor U24682 (N_24682,N_15780,N_16449);
nand U24683 (N_24683,N_17214,N_15080);
and U24684 (N_24684,N_19106,N_18256);
and U24685 (N_24685,N_16818,N_15101);
nand U24686 (N_24686,N_17903,N_16743);
or U24687 (N_24687,N_15092,N_19701);
nand U24688 (N_24688,N_17726,N_16101);
nand U24689 (N_24689,N_16202,N_18422);
or U24690 (N_24690,N_19318,N_17412);
nor U24691 (N_24691,N_17327,N_19493);
nand U24692 (N_24692,N_15031,N_15371);
nand U24693 (N_24693,N_18743,N_17736);
nand U24694 (N_24694,N_19518,N_15434);
or U24695 (N_24695,N_16571,N_16140);
or U24696 (N_24696,N_18178,N_17392);
nand U24697 (N_24697,N_17754,N_15946);
nand U24698 (N_24698,N_16496,N_19615);
nor U24699 (N_24699,N_15999,N_19598);
nand U24700 (N_24700,N_19713,N_19717);
nand U24701 (N_24701,N_17212,N_18000);
and U24702 (N_24702,N_16380,N_17144);
xor U24703 (N_24703,N_15892,N_16972);
nand U24704 (N_24704,N_19169,N_16691);
nor U24705 (N_24705,N_17499,N_18029);
nand U24706 (N_24706,N_15584,N_19974);
nor U24707 (N_24707,N_17814,N_18153);
or U24708 (N_24708,N_17930,N_19942);
nor U24709 (N_24709,N_19111,N_18765);
xnor U24710 (N_24710,N_18528,N_19023);
nand U24711 (N_24711,N_16627,N_19960);
nand U24712 (N_24712,N_16903,N_15832);
or U24713 (N_24713,N_16661,N_16601);
xnor U24714 (N_24714,N_18207,N_19827);
nand U24715 (N_24715,N_18742,N_15266);
or U24716 (N_24716,N_18455,N_17274);
nor U24717 (N_24717,N_17258,N_18939);
or U24718 (N_24718,N_15893,N_15869);
xor U24719 (N_24719,N_15514,N_16709);
nand U24720 (N_24720,N_15023,N_16266);
nor U24721 (N_24721,N_17949,N_15276);
xor U24722 (N_24722,N_18115,N_15169);
and U24723 (N_24723,N_17564,N_19775);
nand U24724 (N_24724,N_19525,N_15169);
nor U24725 (N_24725,N_15170,N_17156);
nand U24726 (N_24726,N_16080,N_16624);
or U24727 (N_24727,N_18894,N_15872);
nor U24728 (N_24728,N_18625,N_16790);
or U24729 (N_24729,N_17876,N_16834);
nor U24730 (N_24730,N_17116,N_16797);
or U24731 (N_24731,N_15215,N_15543);
and U24732 (N_24732,N_17329,N_17646);
xnor U24733 (N_24733,N_17441,N_18241);
nand U24734 (N_24734,N_19908,N_19118);
xor U24735 (N_24735,N_19635,N_18317);
nand U24736 (N_24736,N_16378,N_16544);
and U24737 (N_24737,N_18459,N_19567);
nand U24738 (N_24738,N_16360,N_17860);
or U24739 (N_24739,N_16411,N_17309);
and U24740 (N_24740,N_17516,N_15004);
nor U24741 (N_24741,N_17304,N_17906);
nor U24742 (N_24742,N_16221,N_16393);
nand U24743 (N_24743,N_15553,N_15560);
xor U24744 (N_24744,N_16457,N_19799);
xor U24745 (N_24745,N_17299,N_15350);
or U24746 (N_24746,N_16364,N_19971);
and U24747 (N_24747,N_17553,N_17568);
xor U24748 (N_24748,N_15966,N_17318);
or U24749 (N_24749,N_19613,N_16110);
nand U24750 (N_24750,N_17778,N_15999);
and U24751 (N_24751,N_17273,N_15521);
or U24752 (N_24752,N_17713,N_18257);
xnor U24753 (N_24753,N_16451,N_18504);
xor U24754 (N_24754,N_16088,N_16487);
nand U24755 (N_24755,N_17851,N_15159);
xor U24756 (N_24756,N_15199,N_18666);
or U24757 (N_24757,N_17126,N_18135);
and U24758 (N_24758,N_15372,N_17615);
or U24759 (N_24759,N_19986,N_17942);
and U24760 (N_24760,N_19665,N_15906);
nor U24761 (N_24761,N_16583,N_15030);
nor U24762 (N_24762,N_19664,N_18739);
or U24763 (N_24763,N_16617,N_16307);
and U24764 (N_24764,N_15748,N_15413);
nand U24765 (N_24765,N_18474,N_17284);
nand U24766 (N_24766,N_17365,N_18908);
nand U24767 (N_24767,N_19934,N_18953);
and U24768 (N_24768,N_15140,N_18974);
or U24769 (N_24769,N_17001,N_18954);
and U24770 (N_24770,N_18570,N_19371);
or U24771 (N_24771,N_17830,N_18241);
xnor U24772 (N_24772,N_15133,N_17231);
or U24773 (N_24773,N_16108,N_16411);
xor U24774 (N_24774,N_15057,N_16370);
and U24775 (N_24775,N_15954,N_16363);
xor U24776 (N_24776,N_15055,N_19047);
nand U24777 (N_24777,N_18058,N_16697);
xnor U24778 (N_24778,N_18540,N_18515);
nor U24779 (N_24779,N_18728,N_16626);
xor U24780 (N_24780,N_19123,N_19721);
xor U24781 (N_24781,N_15486,N_17950);
nor U24782 (N_24782,N_16468,N_19454);
or U24783 (N_24783,N_15403,N_16468);
xor U24784 (N_24784,N_15506,N_17294);
xnor U24785 (N_24785,N_19911,N_15350);
nor U24786 (N_24786,N_16379,N_17592);
nor U24787 (N_24787,N_16771,N_19761);
and U24788 (N_24788,N_19388,N_15614);
xor U24789 (N_24789,N_17683,N_16999);
nor U24790 (N_24790,N_18612,N_17936);
nand U24791 (N_24791,N_15718,N_16906);
nor U24792 (N_24792,N_15173,N_17312);
and U24793 (N_24793,N_18065,N_16954);
nand U24794 (N_24794,N_18016,N_19367);
nor U24795 (N_24795,N_17158,N_18823);
nand U24796 (N_24796,N_16509,N_16074);
or U24797 (N_24797,N_16276,N_17173);
and U24798 (N_24798,N_16166,N_18049);
or U24799 (N_24799,N_19720,N_19549);
nand U24800 (N_24800,N_17248,N_15161);
and U24801 (N_24801,N_15139,N_15596);
nand U24802 (N_24802,N_19380,N_16262);
or U24803 (N_24803,N_18054,N_19751);
xor U24804 (N_24804,N_15695,N_15330);
nand U24805 (N_24805,N_15525,N_15988);
or U24806 (N_24806,N_19082,N_19422);
nor U24807 (N_24807,N_16662,N_15893);
nand U24808 (N_24808,N_17178,N_17730);
nand U24809 (N_24809,N_16863,N_19945);
nor U24810 (N_24810,N_16565,N_16971);
or U24811 (N_24811,N_18430,N_15121);
or U24812 (N_24812,N_15259,N_17073);
xor U24813 (N_24813,N_16025,N_16228);
or U24814 (N_24814,N_19497,N_19177);
xor U24815 (N_24815,N_17354,N_17476);
nor U24816 (N_24816,N_17898,N_19591);
nor U24817 (N_24817,N_17736,N_16106);
nand U24818 (N_24818,N_18973,N_16901);
or U24819 (N_24819,N_18120,N_15814);
or U24820 (N_24820,N_17852,N_18812);
nand U24821 (N_24821,N_17133,N_18252);
nor U24822 (N_24822,N_15855,N_18416);
nand U24823 (N_24823,N_16253,N_16450);
nor U24824 (N_24824,N_18389,N_17810);
and U24825 (N_24825,N_16162,N_16330);
nor U24826 (N_24826,N_18644,N_17989);
or U24827 (N_24827,N_18852,N_17685);
nor U24828 (N_24828,N_15376,N_19047);
xnor U24829 (N_24829,N_19216,N_15120);
or U24830 (N_24830,N_16573,N_17177);
and U24831 (N_24831,N_17844,N_17094);
and U24832 (N_24832,N_19833,N_15837);
nor U24833 (N_24833,N_17999,N_19506);
or U24834 (N_24834,N_15910,N_17220);
and U24835 (N_24835,N_17981,N_17248);
or U24836 (N_24836,N_16708,N_15009);
and U24837 (N_24837,N_18869,N_19026);
xor U24838 (N_24838,N_17722,N_15074);
xnor U24839 (N_24839,N_19603,N_15263);
nand U24840 (N_24840,N_17040,N_15725);
xnor U24841 (N_24841,N_15169,N_19637);
and U24842 (N_24842,N_15251,N_16546);
nor U24843 (N_24843,N_15665,N_19568);
or U24844 (N_24844,N_19208,N_19567);
or U24845 (N_24845,N_17370,N_17024);
xor U24846 (N_24846,N_16276,N_17999);
nand U24847 (N_24847,N_19487,N_18223);
xnor U24848 (N_24848,N_19281,N_19983);
and U24849 (N_24849,N_18644,N_15474);
nand U24850 (N_24850,N_15162,N_16216);
xnor U24851 (N_24851,N_18222,N_16736);
or U24852 (N_24852,N_19150,N_18950);
nand U24853 (N_24853,N_18307,N_17352);
xnor U24854 (N_24854,N_19687,N_16650);
and U24855 (N_24855,N_18400,N_16011);
xor U24856 (N_24856,N_16507,N_18495);
or U24857 (N_24857,N_18478,N_18516);
nand U24858 (N_24858,N_18468,N_16806);
nor U24859 (N_24859,N_19418,N_17864);
xor U24860 (N_24860,N_19074,N_15694);
nand U24861 (N_24861,N_19461,N_17534);
and U24862 (N_24862,N_17564,N_15772);
and U24863 (N_24863,N_18322,N_15674);
nand U24864 (N_24864,N_19902,N_16754);
nor U24865 (N_24865,N_17056,N_16046);
xor U24866 (N_24866,N_18664,N_16247);
xor U24867 (N_24867,N_15162,N_19241);
or U24868 (N_24868,N_15970,N_17328);
or U24869 (N_24869,N_17118,N_19566);
nand U24870 (N_24870,N_15180,N_17810);
xnor U24871 (N_24871,N_19327,N_17679);
nand U24872 (N_24872,N_17270,N_19060);
nand U24873 (N_24873,N_17842,N_18200);
xor U24874 (N_24874,N_18287,N_17777);
nor U24875 (N_24875,N_15292,N_18728);
nor U24876 (N_24876,N_18502,N_18954);
xor U24877 (N_24877,N_19802,N_19835);
and U24878 (N_24878,N_15808,N_19814);
and U24879 (N_24879,N_17372,N_17380);
or U24880 (N_24880,N_19265,N_15894);
nand U24881 (N_24881,N_17782,N_17378);
xnor U24882 (N_24882,N_16199,N_18435);
xnor U24883 (N_24883,N_18457,N_19219);
nor U24884 (N_24884,N_16247,N_18266);
or U24885 (N_24885,N_18461,N_17485);
nor U24886 (N_24886,N_16469,N_15257);
and U24887 (N_24887,N_15614,N_19774);
and U24888 (N_24888,N_18549,N_17636);
or U24889 (N_24889,N_19139,N_16888);
nand U24890 (N_24890,N_19979,N_17795);
nand U24891 (N_24891,N_17096,N_19982);
nor U24892 (N_24892,N_19657,N_18051);
nor U24893 (N_24893,N_19799,N_16717);
nand U24894 (N_24894,N_16402,N_19449);
or U24895 (N_24895,N_17880,N_19981);
xnor U24896 (N_24896,N_19883,N_19458);
nor U24897 (N_24897,N_15189,N_15536);
nor U24898 (N_24898,N_16164,N_18097);
and U24899 (N_24899,N_18111,N_17176);
xor U24900 (N_24900,N_19022,N_16403);
xnor U24901 (N_24901,N_19396,N_17432);
and U24902 (N_24902,N_17932,N_17601);
nor U24903 (N_24903,N_18026,N_16801);
xnor U24904 (N_24904,N_16384,N_15242);
nand U24905 (N_24905,N_18563,N_16991);
and U24906 (N_24906,N_15484,N_18662);
and U24907 (N_24907,N_15242,N_18877);
nor U24908 (N_24908,N_17314,N_19823);
xor U24909 (N_24909,N_16432,N_17619);
nand U24910 (N_24910,N_18202,N_17199);
xnor U24911 (N_24911,N_17399,N_18846);
nand U24912 (N_24912,N_16438,N_17565);
xnor U24913 (N_24913,N_17370,N_15184);
and U24914 (N_24914,N_17602,N_18214);
xor U24915 (N_24915,N_15159,N_19321);
nor U24916 (N_24916,N_16283,N_19769);
xnor U24917 (N_24917,N_17153,N_15374);
xnor U24918 (N_24918,N_18675,N_18505);
or U24919 (N_24919,N_17628,N_17884);
xnor U24920 (N_24920,N_15246,N_19744);
and U24921 (N_24921,N_16606,N_15091);
and U24922 (N_24922,N_17681,N_18575);
or U24923 (N_24923,N_19476,N_17249);
nand U24924 (N_24924,N_18657,N_18887);
and U24925 (N_24925,N_19546,N_19132);
nand U24926 (N_24926,N_18623,N_16113);
nand U24927 (N_24927,N_16443,N_19940);
nand U24928 (N_24928,N_17241,N_17365);
and U24929 (N_24929,N_18600,N_16843);
xor U24930 (N_24930,N_16945,N_16817);
nor U24931 (N_24931,N_18385,N_18991);
nor U24932 (N_24932,N_19938,N_17121);
and U24933 (N_24933,N_18384,N_18040);
and U24934 (N_24934,N_15417,N_16281);
and U24935 (N_24935,N_16736,N_19467);
xnor U24936 (N_24936,N_17008,N_16272);
and U24937 (N_24937,N_17436,N_18827);
nand U24938 (N_24938,N_18374,N_19961);
or U24939 (N_24939,N_19976,N_15898);
nand U24940 (N_24940,N_16493,N_18997);
or U24941 (N_24941,N_16810,N_16576);
nor U24942 (N_24942,N_17874,N_16341);
or U24943 (N_24943,N_18544,N_16164);
xnor U24944 (N_24944,N_16387,N_17640);
or U24945 (N_24945,N_16732,N_19422);
or U24946 (N_24946,N_16814,N_18466);
xor U24947 (N_24947,N_19287,N_18865);
and U24948 (N_24948,N_18364,N_17885);
nand U24949 (N_24949,N_16514,N_17148);
nand U24950 (N_24950,N_15658,N_19244);
nand U24951 (N_24951,N_16299,N_18203);
xnor U24952 (N_24952,N_17524,N_19363);
xnor U24953 (N_24953,N_19456,N_16309);
xnor U24954 (N_24954,N_17753,N_19307);
nor U24955 (N_24955,N_18063,N_19914);
or U24956 (N_24956,N_17643,N_16870);
or U24957 (N_24957,N_16542,N_18196);
xor U24958 (N_24958,N_19254,N_18527);
or U24959 (N_24959,N_18561,N_16707);
xor U24960 (N_24960,N_16376,N_19423);
xnor U24961 (N_24961,N_16205,N_19905);
xor U24962 (N_24962,N_16619,N_19334);
xnor U24963 (N_24963,N_19502,N_16921);
and U24964 (N_24964,N_18931,N_17095);
or U24965 (N_24965,N_16601,N_15901);
or U24966 (N_24966,N_15561,N_16051);
nor U24967 (N_24967,N_17627,N_18098);
xnor U24968 (N_24968,N_17349,N_16667);
or U24969 (N_24969,N_15067,N_17717);
or U24970 (N_24970,N_15692,N_15836);
or U24971 (N_24971,N_17716,N_16837);
or U24972 (N_24972,N_19086,N_18281);
nand U24973 (N_24973,N_18722,N_19364);
or U24974 (N_24974,N_17098,N_19045);
and U24975 (N_24975,N_17318,N_17356);
and U24976 (N_24976,N_18290,N_19956);
and U24977 (N_24977,N_15469,N_18288);
and U24978 (N_24978,N_17430,N_18244);
xnor U24979 (N_24979,N_16865,N_18785);
nand U24980 (N_24980,N_16861,N_18406);
xnor U24981 (N_24981,N_15823,N_19933);
or U24982 (N_24982,N_17317,N_15622);
nand U24983 (N_24983,N_17089,N_19523);
nor U24984 (N_24984,N_15747,N_19503);
and U24985 (N_24985,N_16483,N_16550);
nand U24986 (N_24986,N_15325,N_17399);
xnor U24987 (N_24987,N_18382,N_18030);
xnor U24988 (N_24988,N_17211,N_18762);
or U24989 (N_24989,N_18565,N_16066);
nand U24990 (N_24990,N_19668,N_19847);
nand U24991 (N_24991,N_18734,N_18786);
nand U24992 (N_24992,N_15687,N_17033);
or U24993 (N_24993,N_18959,N_19445);
nor U24994 (N_24994,N_19286,N_18500);
nand U24995 (N_24995,N_19976,N_19870);
and U24996 (N_24996,N_19352,N_17249);
nor U24997 (N_24997,N_16613,N_16158);
nand U24998 (N_24998,N_17198,N_16416);
nand U24999 (N_24999,N_16459,N_18572);
xor UO_0 (O_0,N_21087,N_23069);
and UO_1 (O_1,N_22154,N_22315);
nor UO_2 (O_2,N_20732,N_20830);
and UO_3 (O_3,N_24845,N_23198);
nor UO_4 (O_4,N_21939,N_24920);
nand UO_5 (O_5,N_23763,N_24215);
nand UO_6 (O_6,N_21821,N_24690);
and UO_7 (O_7,N_20667,N_21469);
nor UO_8 (O_8,N_20398,N_21603);
xnor UO_9 (O_9,N_24676,N_21443);
or UO_10 (O_10,N_23964,N_24990);
nand UO_11 (O_11,N_21880,N_24239);
nor UO_12 (O_12,N_23614,N_24014);
or UO_13 (O_13,N_23825,N_24592);
xor UO_14 (O_14,N_20976,N_24611);
xnor UO_15 (O_15,N_22935,N_23701);
nor UO_16 (O_16,N_22449,N_21446);
nand UO_17 (O_17,N_21452,N_21424);
xor UO_18 (O_18,N_21702,N_20767);
or UO_19 (O_19,N_20046,N_20781);
nand UO_20 (O_20,N_23549,N_20442);
xor UO_21 (O_21,N_24143,N_20605);
and UO_22 (O_22,N_23298,N_23903);
xnor UO_23 (O_23,N_20344,N_20162);
and UO_24 (O_24,N_24222,N_21607);
or UO_25 (O_25,N_22396,N_23735);
nand UO_26 (O_26,N_21455,N_23263);
nor UO_27 (O_27,N_24644,N_23906);
nor UO_28 (O_28,N_23514,N_22827);
and UO_29 (O_29,N_23843,N_22503);
or UO_30 (O_30,N_21260,N_24955);
or UO_31 (O_31,N_20588,N_22608);
or UO_32 (O_32,N_20299,N_21206);
nand UO_33 (O_33,N_24498,N_22453);
nor UO_34 (O_34,N_21368,N_23796);
xnor UO_35 (O_35,N_23869,N_24240);
xnor UO_36 (O_36,N_22340,N_20078);
xnor UO_37 (O_37,N_21136,N_24178);
nand UO_38 (O_38,N_20674,N_21833);
or UO_39 (O_39,N_20967,N_20713);
or UO_40 (O_40,N_20384,N_21273);
and UO_41 (O_41,N_23540,N_23545);
or UO_42 (O_42,N_23314,N_22530);
and UO_43 (O_43,N_22986,N_21406);
xnor UO_44 (O_44,N_23303,N_22591);
nor UO_45 (O_45,N_22290,N_23343);
xnor UO_46 (O_46,N_22870,N_22890);
xor UO_47 (O_47,N_21681,N_20677);
or UO_48 (O_48,N_20289,N_20184);
or UO_49 (O_49,N_24510,N_22136);
xor UO_50 (O_50,N_23768,N_20323);
nor UO_51 (O_51,N_22514,N_20353);
or UO_52 (O_52,N_22966,N_23911);
nor UO_53 (O_53,N_24581,N_20678);
nor UO_54 (O_54,N_20108,N_20064);
or UO_55 (O_55,N_24162,N_20471);
nor UO_56 (O_56,N_22920,N_23334);
nor UO_57 (O_57,N_22317,N_23460);
nand UO_58 (O_58,N_24088,N_22145);
nand UO_59 (O_59,N_23889,N_24457);
nand UO_60 (O_60,N_24115,N_22465);
nor UO_61 (O_61,N_21106,N_20861);
or UO_62 (O_62,N_21505,N_22872);
xor UO_63 (O_63,N_21881,N_24259);
or UO_64 (O_64,N_20187,N_23446);
nor UO_65 (O_65,N_24632,N_21388);
and UO_66 (O_66,N_24709,N_23943);
or UO_67 (O_67,N_21180,N_24749);
and UO_68 (O_68,N_21904,N_21060);
nand UO_69 (O_69,N_20082,N_24898);
nor UO_70 (O_70,N_20230,N_24811);
nand UO_71 (O_71,N_21430,N_21027);
and UO_72 (O_72,N_24782,N_21875);
nand UO_73 (O_73,N_23815,N_20419);
nor UO_74 (O_74,N_23861,N_24145);
nand UO_75 (O_75,N_23018,N_21310);
or UO_76 (O_76,N_24347,N_21265);
and UO_77 (O_77,N_21634,N_20107);
nor UO_78 (O_78,N_20610,N_23956);
and UO_79 (O_79,N_21924,N_20087);
xor UO_80 (O_80,N_22841,N_22450);
nand UO_81 (O_81,N_22907,N_23800);
and UO_82 (O_82,N_23270,N_20517);
nand UO_83 (O_83,N_24140,N_22210);
nand UO_84 (O_84,N_22753,N_23132);
nor UO_85 (O_85,N_20603,N_20691);
nor UO_86 (O_86,N_20349,N_24905);
xor UO_87 (O_87,N_23096,N_20488);
nor UO_88 (O_88,N_21520,N_21364);
nor UO_89 (O_89,N_21556,N_20232);
nand UO_90 (O_90,N_23135,N_23526);
nand UO_91 (O_91,N_23332,N_24667);
and UO_92 (O_92,N_22008,N_21357);
nand UO_93 (O_93,N_21767,N_21781);
or UO_94 (O_94,N_24480,N_24999);
xnor UO_95 (O_95,N_20446,N_23422);
xnor UO_96 (O_96,N_23575,N_21196);
nand UO_97 (O_97,N_23715,N_21033);
xor UO_98 (O_98,N_24303,N_20258);
nor UO_99 (O_99,N_22551,N_21183);
and UO_100 (O_100,N_21646,N_21705);
xor UO_101 (O_101,N_21089,N_21953);
nand UO_102 (O_102,N_20979,N_22233);
nand UO_103 (O_103,N_21928,N_24937);
and UO_104 (O_104,N_23083,N_21951);
nand UO_105 (O_105,N_21411,N_20559);
and UO_106 (O_106,N_20277,N_24291);
and UO_107 (O_107,N_21504,N_22940);
xnor UO_108 (O_108,N_21380,N_20506);
nand UO_109 (O_109,N_23729,N_24852);
xor UO_110 (O_110,N_22401,N_23027);
and UO_111 (O_111,N_23536,N_24979);
and UO_112 (O_112,N_23783,N_21529);
or UO_113 (O_113,N_24664,N_23791);
and UO_114 (O_114,N_23011,N_23838);
or UO_115 (O_115,N_20362,N_20854);
xor UO_116 (O_116,N_23180,N_21020);
and UO_117 (O_117,N_22652,N_24702);
xor UO_118 (O_118,N_20132,N_23014);
and UO_119 (O_119,N_22319,N_20098);
nand UO_120 (O_120,N_20381,N_21171);
and UO_121 (O_121,N_22772,N_23564);
or UO_122 (O_122,N_24833,N_21476);
and UO_123 (O_123,N_24666,N_21382);
xor UO_124 (O_124,N_22217,N_23146);
nor UO_125 (O_125,N_24573,N_23899);
and UO_126 (O_126,N_21137,N_23853);
nor UO_127 (O_127,N_20965,N_21842);
and UO_128 (O_128,N_23053,N_21207);
nand UO_129 (O_129,N_20804,N_24562);
and UO_130 (O_130,N_21495,N_20298);
and UO_131 (O_131,N_24152,N_22277);
or UO_132 (O_132,N_20879,N_23055);
nor UO_133 (O_133,N_24229,N_21947);
and UO_134 (O_134,N_23659,N_22385);
nor UO_135 (O_135,N_24725,N_24308);
xor UO_136 (O_136,N_24362,N_21844);
and UO_137 (O_137,N_23913,N_24385);
and UO_138 (O_138,N_22538,N_20399);
xor UO_139 (O_139,N_21254,N_22049);
or UO_140 (O_140,N_21537,N_23547);
nor UO_141 (O_141,N_23704,N_24449);
nand UO_142 (O_142,N_20460,N_24302);
or UO_143 (O_143,N_24181,N_20757);
nand UO_144 (O_144,N_21262,N_20573);
xor UO_145 (O_145,N_21800,N_20891);
nand UO_146 (O_146,N_22331,N_24430);
nand UO_147 (O_147,N_22961,N_22824);
xor UO_148 (O_148,N_22087,N_22207);
nor UO_149 (O_149,N_23076,N_24049);
nand UO_150 (O_150,N_23483,N_22932);
xor UO_151 (O_151,N_24057,N_20139);
and UO_152 (O_152,N_23808,N_23229);
or UO_153 (O_153,N_20120,N_21783);
xor UO_154 (O_154,N_20012,N_24093);
nor UO_155 (O_155,N_23551,N_23125);
nand UO_156 (O_156,N_23289,N_22904);
nand UO_157 (O_157,N_22433,N_21801);
nor UO_158 (O_158,N_20008,N_21226);
nor UO_159 (O_159,N_21331,N_22967);
nor UO_160 (O_160,N_21359,N_23066);
nand UO_161 (O_161,N_22659,N_21722);
nor UO_162 (O_162,N_23522,N_20953);
and UO_163 (O_163,N_23003,N_20073);
xor UO_164 (O_164,N_22146,N_20943);
nand UO_165 (O_165,N_21779,N_23831);
nor UO_166 (O_166,N_20500,N_24962);
xnor UO_167 (O_167,N_23578,N_23766);
xnor UO_168 (O_168,N_23231,N_21124);
or UO_169 (O_169,N_22731,N_23778);
xnor UO_170 (O_170,N_22378,N_24201);
and UO_171 (O_171,N_20646,N_21069);
nand UO_172 (O_172,N_22209,N_20328);
xor UO_173 (O_173,N_24647,N_24807);
xor UO_174 (O_174,N_20701,N_20870);
nor UO_175 (O_175,N_22786,N_22617);
nand UO_176 (O_176,N_21894,N_20027);
xnor UO_177 (O_177,N_24295,N_20496);
and UO_178 (O_178,N_20877,N_24860);
nor UO_179 (O_179,N_20351,N_24559);
xor UO_180 (O_180,N_22436,N_22257);
xor UO_181 (O_181,N_22911,N_22603);
or UO_182 (O_182,N_24328,N_22361);
nor UO_183 (O_183,N_23423,N_23161);
or UO_184 (O_184,N_21445,N_21140);
nor UO_185 (O_185,N_21503,N_20156);
or UO_186 (O_186,N_21019,N_21150);
and UO_187 (O_187,N_22583,N_24515);
xnor UO_188 (O_188,N_20819,N_23216);
nand UO_189 (O_189,N_22736,N_21478);
xnor UO_190 (O_190,N_23739,N_22339);
and UO_191 (O_191,N_23010,N_24585);
nor UO_192 (O_192,N_20695,N_24820);
or UO_193 (O_193,N_21237,N_20878);
and UO_194 (O_194,N_22393,N_22611);
and UO_195 (O_195,N_24940,N_24475);
nand UO_196 (O_196,N_21270,N_24848);
nor UO_197 (O_197,N_24520,N_22579);
nand UO_198 (O_198,N_21619,N_20458);
nor UO_199 (O_199,N_24441,N_24737);
nand UO_200 (O_200,N_23392,N_24629);
and UO_201 (O_201,N_20658,N_21696);
and UO_202 (O_202,N_21194,N_20746);
nor UO_203 (O_203,N_24624,N_20850);
nand UO_204 (O_204,N_22461,N_20478);
and UO_205 (O_205,N_22797,N_21458);
xor UO_206 (O_206,N_22712,N_24231);
nor UO_207 (O_207,N_24293,N_21795);
or UO_208 (O_208,N_24822,N_24204);
nand UO_209 (O_209,N_24696,N_23622);
xnor UO_210 (O_210,N_24772,N_24356);
xnor UO_211 (O_211,N_23108,N_23344);
nor UO_212 (O_212,N_23759,N_24733);
or UO_213 (O_213,N_23402,N_23686);
nor UO_214 (O_214,N_24275,N_20911);
and UO_215 (O_215,N_21958,N_20459);
or UO_216 (O_216,N_22180,N_24658);
nand UO_217 (O_217,N_24729,N_21519);
or UO_218 (O_218,N_22025,N_23394);
or UO_219 (O_219,N_24031,N_21094);
nor UO_220 (O_220,N_20743,N_22467);
xnor UO_221 (O_221,N_21363,N_21267);
nand UO_222 (O_222,N_24048,N_21949);
xor UO_223 (O_223,N_22586,N_21749);
nand UO_224 (O_224,N_22948,N_21885);
or UO_225 (O_225,N_22404,N_23100);
nor UO_226 (O_226,N_20973,N_24880);
and UO_227 (O_227,N_22009,N_20243);
and UO_228 (O_228,N_22446,N_21046);
and UO_229 (O_229,N_20469,N_23897);
nand UO_230 (O_230,N_22704,N_23994);
xor UO_231 (O_231,N_20699,N_23958);
nor UO_232 (O_232,N_23874,N_23833);
nor UO_233 (O_233,N_23465,N_23002);
or UO_234 (O_234,N_23090,N_22545);
nor UO_235 (O_235,N_22980,N_24333);
nor UO_236 (O_236,N_23682,N_21630);
nor UO_237 (O_237,N_24731,N_22163);
and UO_238 (O_238,N_23203,N_21921);
xor UO_239 (O_239,N_24587,N_24500);
nor UO_240 (O_240,N_24353,N_24675);
nand UO_241 (O_241,N_21620,N_22480);
nor UO_242 (O_242,N_22610,N_22318);
or UO_243 (O_243,N_23837,N_24322);
nand UO_244 (O_244,N_20515,N_23208);
nand UO_245 (O_245,N_22165,N_22645);
nand UO_246 (O_246,N_23746,N_23388);
nand UO_247 (O_247,N_24311,N_20915);
nand UO_248 (O_248,N_21311,N_24223);
and UO_249 (O_249,N_23859,N_22255);
nor UO_250 (O_250,N_24509,N_20609);
nor UO_251 (O_251,N_20267,N_23482);
nor UO_252 (O_252,N_21272,N_20571);
xor UO_253 (O_253,N_22684,N_23890);
and UO_254 (O_254,N_22701,N_24174);
nand UO_255 (O_255,N_21733,N_24608);
nand UO_256 (O_256,N_22239,N_22708);
or UO_257 (O_257,N_21605,N_23111);
nor UO_258 (O_258,N_23472,N_23745);
or UO_259 (O_259,N_20251,N_21253);
or UO_260 (O_260,N_23645,N_21465);
nor UO_261 (O_261,N_22240,N_23519);
or UO_262 (O_262,N_22153,N_22668);
and UO_263 (O_263,N_23448,N_23271);
and UO_264 (O_264,N_22418,N_24993);
nand UO_265 (O_265,N_24859,N_24580);
or UO_266 (O_266,N_21299,N_20708);
xnor UO_267 (O_267,N_21610,N_22375);
or UO_268 (O_268,N_21732,N_22624);
nand UO_269 (O_269,N_24444,N_23753);
and UO_270 (O_270,N_21297,N_23374);
nand UO_271 (O_271,N_21650,N_23356);
or UO_272 (O_272,N_22099,N_24506);
nor UO_273 (O_273,N_21355,N_23795);
or UO_274 (O_274,N_23417,N_21164);
and UO_275 (O_275,N_24554,N_22291);
xor UO_276 (O_276,N_21523,N_22666);
nor UO_277 (O_277,N_22280,N_21026);
or UO_278 (O_278,N_24829,N_23470);
and UO_279 (O_279,N_24134,N_21028);
or UO_280 (O_280,N_21551,N_24996);
nor UO_281 (O_281,N_20433,N_24892);
xor UO_282 (O_282,N_24938,N_21323);
xor UO_283 (O_283,N_20210,N_24242);
and UO_284 (O_284,N_21441,N_21405);
nand UO_285 (O_285,N_23754,N_22581);
nor UO_286 (O_286,N_21641,N_22327);
nand UO_287 (O_287,N_24361,N_20390);
xnor UO_288 (O_288,N_21582,N_20016);
xor UO_289 (O_289,N_20339,N_24751);
nand UO_290 (O_290,N_24808,N_23406);
nand UO_291 (O_291,N_24989,N_21809);
xnor UO_292 (O_292,N_23802,N_21437);
or UO_293 (O_293,N_24071,N_20633);
nand UO_294 (O_294,N_24233,N_21855);
or UO_295 (O_295,N_23077,N_20436);
nor UO_296 (O_296,N_23663,N_22761);
and UO_297 (O_297,N_22542,N_23342);
xor UO_298 (O_298,N_20581,N_23565);
nand UO_299 (O_299,N_20839,N_21662);
nor UO_300 (O_300,N_20017,N_23299);
and UO_301 (O_301,N_20921,N_21989);
or UO_302 (O_302,N_20712,N_21473);
and UO_303 (O_303,N_22588,N_20681);
and UO_304 (O_304,N_24793,N_21922);
nor UO_305 (O_305,N_20060,N_24327);
and UO_306 (O_306,N_22281,N_20733);
and UO_307 (O_307,N_24387,N_20179);
xnor UO_308 (O_308,N_23484,N_20616);
or UO_309 (O_309,N_24916,N_22929);
or UO_310 (O_310,N_21806,N_23331);
nand UO_311 (O_311,N_23431,N_20273);
and UO_312 (O_312,N_24238,N_23941);
xor UO_313 (O_313,N_23412,N_23553);
nand UO_314 (O_314,N_24493,N_24505);
nand UO_315 (O_315,N_23247,N_23137);
xnor UO_316 (O_316,N_21526,N_23477);
nor UO_317 (O_317,N_21825,N_22424);
xnor UO_318 (O_318,N_21577,N_20578);
nor UO_319 (O_319,N_20324,N_20791);
or UO_320 (O_320,N_22429,N_23278);
nor UO_321 (O_321,N_23613,N_21366);
nand UO_322 (O_322,N_24078,N_20473);
nand UO_323 (O_323,N_23914,N_22286);
nor UO_324 (O_324,N_23839,N_20426);
or UO_325 (O_325,N_20760,N_21711);
and UO_326 (O_326,N_20929,N_23325);
and UO_327 (O_327,N_21750,N_24159);
xor UO_328 (O_328,N_20524,N_20306);
xor UO_329 (O_329,N_20886,N_24487);
or UO_330 (O_330,N_21828,N_23366);
nand UO_331 (O_331,N_24199,N_20874);
nand UO_332 (O_332,N_21317,N_22633);
or UO_333 (O_333,N_24502,N_23269);
and UO_334 (O_334,N_20159,N_21788);
or UO_335 (O_335,N_21500,N_21914);
and UO_336 (O_336,N_22459,N_20872);
nand UO_337 (O_337,N_21704,N_24074);
or UO_338 (O_338,N_23318,N_23886);
nor UO_339 (O_339,N_22970,N_23139);
or UO_340 (O_340,N_22862,N_24906);
or UO_341 (O_341,N_24879,N_20574);
nand UO_342 (O_342,N_24010,N_22580);
nand UO_343 (O_343,N_21707,N_21148);
and UO_344 (O_344,N_24352,N_21775);
nor UO_345 (O_345,N_24455,N_23749);
nor UO_346 (O_346,N_24728,N_20183);
or UO_347 (O_347,N_21435,N_21906);
xor UO_348 (O_348,N_24830,N_20577);
nand UO_349 (O_349,N_20882,N_24260);
nor UO_350 (O_350,N_24389,N_21127);
or UO_351 (O_351,N_21490,N_23871);
nor UO_352 (O_352,N_24818,N_24411);
or UO_353 (O_353,N_23166,N_23326);
xor UO_354 (O_354,N_20317,N_24698);
xnor UO_355 (O_355,N_22560,N_22715);
xnor UO_356 (O_356,N_22440,N_23103);
and UO_357 (O_357,N_21964,N_20754);
nand UO_358 (O_358,N_20376,N_20498);
nand UO_359 (O_359,N_22190,N_23275);
xnor UO_360 (O_360,N_23721,N_24780);
and UO_361 (O_361,N_24123,N_20736);
nand UO_362 (O_362,N_24301,N_23567);
nand UO_363 (O_363,N_23133,N_24410);
and UO_364 (O_364,N_22636,N_23028);
xor UO_365 (O_365,N_22962,N_21428);
and UO_366 (O_366,N_20989,N_24715);
xnor UO_367 (O_367,N_23487,N_24972);
or UO_368 (O_368,N_23572,N_22294);
xor UO_369 (O_369,N_22139,N_22822);
nand UO_370 (O_370,N_23489,N_20123);
nand UO_371 (O_371,N_20218,N_23718);
or UO_372 (O_372,N_21623,N_22628);
and UO_373 (O_373,N_21167,N_22350);
nand UO_374 (O_374,N_20962,N_23820);
xor UO_375 (O_375,N_20029,N_20537);
nand UO_376 (O_376,N_21116,N_20494);
nor UO_377 (O_377,N_22695,N_20966);
nor UO_378 (O_378,N_24288,N_24236);
nand UO_379 (O_379,N_24439,N_20355);
nand UO_380 (O_380,N_21118,N_22839);
nand UO_381 (O_381,N_22992,N_24628);
nor UO_382 (O_382,N_20930,N_20836);
nor UO_383 (O_383,N_24104,N_20824);
or UO_384 (O_384,N_24743,N_23782);
nor UO_385 (O_385,N_23576,N_23873);
xor UO_386 (O_386,N_20007,N_23401);
nor UO_387 (O_387,N_20203,N_22760);
or UO_388 (O_388,N_21786,N_24366);
and UO_389 (O_389,N_24679,N_23142);
nand UO_390 (O_390,N_22046,N_23641);
nor UO_391 (O_391,N_21008,N_21957);
and UO_392 (O_392,N_20093,N_24452);
xor UO_393 (O_393,N_23979,N_21778);
and UO_394 (O_394,N_24792,N_22464);
nand UO_395 (O_395,N_22263,N_22482);
nor UO_396 (O_396,N_22414,N_22421);
xor UO_397 (O_397,N_20904,N_20271);
or UO_398 (O_398,N_21793,N_24893);
nand UO_399 (O_399,N_20845,N_24528);
nor UO_400 (O_400,N_24736,N_23305);
nor UO_401 (O_401,N_21349,N_23041);
and UO_402 (O_402,N_21021,N_20825);
nor UO_403 (O_403,N_23781,N_20794);
or UO_404 (O_404,N_23692,N_20618);
nor UO_405 (O_405,N_20084,N_21474);
and UO_406 (O_406,N_23091,N_20660);
or UO_407 (O_407,N_23651,N_20716);
xor UO_408 (O_408,N_22178,N_23123);
and UO_409 (O_409,N_21528,N_20717);
or UO_410 (O_410,N_21549,N_21065);
nor UO_411 (O_411,N_22887,N_23189);
nand UO_412 (O_412,N_20422,N_22654);
or UO_413 (O_413,N_23209,N_20253);
nand UO_414 (O_414,N_21747,N_21758);
nand UO_415 (O_415,N_20725,N_23084);
nor UO_416 (O_416,N_24851,N_24801);
nor UO_417 (O_417,N_21316,N_20615);
and UO_418 (O_418,N_22305,N_21499);
and UO_419 (O_419,N_21764,N_23416);
nor UO_420 (O_420,N_22381,N_24396);
nor UO_421 (O_421,N_24928,N_23670);
nand UO_422 (O_422,N_23360,N_23094);
nor UO_423 (O_423,N_20063,N_23454);
xnor UO_424 (O_424,N_22594,N_24519);
and UO_425 (O_425,N_24331,N_22050);
nand UO_426 (O_426,N_24276,N_22973);
xnor UO_427 (O_427,N_20849,N_23061);
nand UO_428 (O_428,N_24418,N_20127);
nor UO_429 (O_429,N_20800,N_24492);
or UO_430 (O_430,N_24100,N_20670);
xor UO_431 (O_431,N_20745,N_21755);
and UO_432 (O_432,N_22958,N_24533);
xor UO_433 (O_433,N_23677,N_24307);
xor UO_434 (O_434,N_21043,N_20690);
nand UO_435 (O_435,N_21687,N_20675);
xnor UO_436 (O_436,N_22079,N_22916);
nand UO_437 (O_437,N_20213,N_24176);
and UO_438 (O_438,N_21050,N_21063);
nor UO_439 (O_439,N_22223,N_21352);
or UO_440 (O_440,N_20613,N_22292);
or UO_441 (O_441,N_20897,N_24981);
or UO_442 (O_442,N_20417,N_20360);
nor UO_443 (O_443,N_21946,N_23953);
nor UO_444 (O_444,N_24129,N_23998);
nor UO_445 (O_445,N_23188,N_20224);
and UO_446 (O_446,N_24287,N_24324);
nand UO_447 (O_447,N_21120,N_23297);
nand UO_448 (O_448,N_22460,N_21291);
nand UO_449 (O_449,N_21330,N_21131);
xor UO_450 (O_450,N_22574,N_24403);
or UO_451 (O_451,N_20236,N_22891);
or UO_452 (O_452,N_24392,N_22819);
nand UO_453 (O_453,N_21768,N_23447);
nor UO_454 (O_454,N_20579,N_24000);
nor UO_455 (O_455,N_23373,N_23354);
nor UO_456 (O_456,N_23070,N_20553);
xnor UO_457 (O_457,N_24391,N_24024);
or UO_458 (O_458,N_21548,N_22639);
or UO_459 (O_459,N_24791,N_22109);
or UO_460 (O_460,N_22289,N_20510);
nor UO_461 (O_461,N_22805,N_24577);
nand UO_462 (O_462,N_20254,N_22895);
xor UO_463 (O_463,N_20055,N_24740);
nor UO_464 (O_464,N_21570,N_24251);
nor UO_465 (O_465,N_22908,N_24813);
or UO_466 (O_466,N_22376,N_20563);
and UO_467 (O_467,N_20304,N_22673);
nor UO_468 (O_468,N_22549,N_23451);
and UO_469 (O_469,N_21999,N_24045);
nor UO_470 (O_470,N_21918,N_21176);
xor UO_471 (O_471,N_22287,N_23805);
or UO_472 (O_472,N_21190,N_22380);
and UO_473 (O_473,N_20434,N_24289);
and UO_474 (O_474,N_21817,N_22898);
nand UO_475 (O_475,N_22495,N_21153);
and UO_476 (O_476,N_22926,N_22295);
xor UO_477 (O_477,N_20922,N_22686);
xor UO_478 (O_478,N_20913,N_21123);
nor UO_479 (O_479,N_21119,N_21048);
or UO_480 (O_480,N_22325,N_24337);
nand UO_481 (O_481,N_22110,N_22052);
or UO_482 (O_482,N_22373,N_20952);
nand UO_483 (O_483,N_22638,N_21727);
nand UO_484 (O_484,N_23852,N_23822);
nor UO_485 (O_485,N_21514,N_22937);
nor UO_486 (O_486,N_21340,N_23154);
nand UO_487 (O_487,N_23801,N_24163);
and UO_488 (O_488,N_20890,N_23282);
or UO_489 (O_489,N_22179,N_22936);
nand UO_490 (O_490,N_21007,N_21587);
nand UO_491 (O_491,N_23976,N_21155);
nor UO_492 (O_492,N_20439,N_22425);
or UO_493 (O_493,N_20161,N_20977);
and UO_494 (O_494,N_23246,N_23844);
and UO_495 (O_495,N_22757,N_21135);
and UO_496 (O_496,N_24727,N_21487);
nor UO_497 (O_497,N_21369,N_23065);
nor UO_498 (O_498,N_20373,N_20540);
nand UO_499 (O_499,N_21491,N_22730);
nand UO_500 (O_500,N_23301,N_21114);
and UO_501 (O_501,N_22111,N_22525);
or UO_502 (O_502,N_21203,N_20015);
nand UO_503 (O_503,N_20024,N_22707);
and UO_504 (O_504,N_24386,N_23977);
xor UO_505 (O_505,N_22405,N_23039);
xnor UO_506 (O_506,N_23136,N_24683);
xnor UO_507 (O_507,N_20643,N_24089);
nor UO_508 (O_508,N_22546,N_22752);
xor UO_509 (O_509,N_22273,N_22648);
xnor UO_510 (O_510,N_22500,N_22452);
xnor UO_511 (O_511,N_24384,N_21418);
xor UO_512 (O_512,N_20207,N_20405);
and UO_513 (O_513,N_20867,N_20786);
nor UO_514 (O_514,N_20441,N_20639);
nand UO_515 (O_515,N_20350,N_24266);
or UO_516 (O_516,N_21154,N_20764);
nand UO_517 (O_517,N_20755,N_22090);
nand UO_518 (O_518,N_20407,N_21796);
nand UO_519 (O_519,N_23695,N_22466);
nor UO_520 (O_520,N_24125,N_22172);
and UO_521 (O_521,N_20451,N_24931);
xor UO_522 (O_522,N_24547,N_21538);
nand UO_523 (O_523,N_21149,N_23279);
nand UO_524 (O_524,N_21085,N_23044);
nand UO_525 (O_525,N_21572,N_24207);
nor UO_526 (O_526,N_22488,N_21575);
xnor UO_527 (O_527,N_20461,N_24036);
xor UO_528 (O_528,N_22397,N_23458);
nor UO_529 (O_529,N_23038,N_24858);
or UO_530 (O_530,N_24825,N_22523);
nor UO_531 (O_531,N_22147,N_24061);
and UO_532 (O_532,N_23635,N_23957);
or UO_533 (O_533,N_20375,N_24286);
nand UO_534 (O_534,N_23328,N_20283);
and UO_535 (O_535,N_22829,N_23508);
xnor UO_536 (O_536,N_22148,N_20305);
nor UO_537 (O_537,N_23767,N_22828);
and UO_538 (O_538,N_23790,N_20204);
and UO_539 (O_539,N_20910,N_21709);
nand UO_540 (O_540,N_21017,N_20641);
nand UO_541 (O_541,N_23654,N_20898);
or UO_542 (O_542,N_23058,N_22541);
nor UO_543 (O_543,N_23684,N_23047);
nor UO_544 (O_544,N_23528,N_21756);
nand UO_545 (O_545,N_22785,N_22925);
or UO_546 (O_546,N_24596,N_24622);
or UO_547 (O_547,N_22511,N_22477);
nor UO_548 (O_548,N_23436,N_22213);
or UO_549 (O_549,N_24499,N_24323);
nor UO_550 (O_550,N_22930,N_21542);
or UO_551 (O_551,N_20068,N_23673);
and UO_552 (O_552,N_22494,N_21362);
and UO_553 (O_553,N_24535,N_21969);
and UO_554 (O_554,N_21434,N_24175);
nand UO_555 (O_555,N_20126,N_22748);
and UO_556 (O_556,N_22640,N_23232);
or UO_557 (O_557,N_22934,N_20424);
xor UO_558 (O_558,N_21975,N_23597);
nand UO_559 (O_559,N_24075,N_21680);
nor UO_560 (O_560,N_21615,N_22114);
or UO_561 (O_561,N_23437,N_21147);
xor UO_562 (O_562,N_20533,N_22484);
nor UO_563 (O_563,N_22363,N_22774);
and UO_564 (O_564,N_21227,N_23449);
nor UO_565 (O_565,N_22762,N_24939);
nor UO_566 (O_566,N_21617,N_22691);
nor UO_567 (O_567,N_23720,N_24081);
and UO_568 (O_568,N_24472,N_24778);
nand UO_569 (O_569,N_21501,N_21025);
or UO_570 (O_570,N_20659,N_20154);
and UO_571 (O_571,N_24722,N_22854);
and UO_572 (O_572,N_23598,N_24694);
nor UO_573 (O_573,N_21893,N_21054);
xor UO_574 (O_574,N_20916,N_22320);
nor UO_575 (O_575,N_20429,N_24247);
and UO_576 (O_576,N_24522,N_22100);
and UO_577 (O_577,N_24209,N_20173);
nand UO_578 (O_578,N_20340,N_21613);
xnor UO_579 (O_579,N_22042,N_20917);
nand UO_580 (O_580,N_20516,N_20428);
or UO_581 (O_581,N_22568,N_21279);
xnor UO_582 (O_582,N_21863,N_23586);
or UO_583 (O_583,N_21823,N_24855);
or UO_584 (O_584,N_23336,N_23410);
nand UO_585 (O_585,N_24202,N_21962);
or UO_586 (O_586,N_21822,N_21618);
nand UO_587 (O_587,N_22818,N_21410);
or UO_588 (O_588,N_20171,N_21235);
or UO_589 (O_589,N_22019,N_23592);
nor UO_590 (O_590,N_23201,N_21333);
nand UO_591 (O_591,N_22422,N_20318);
or UO_592 (O_592,N_20457,N_23945);
nand UO_593 (O_593,N_20813,N_22602);
nor UO_594 (O_594,N_21166,N_24165);
nor UO_595 (O_595,N_20352,N_22905);
xnor UO_596 (O_596,N_22412,N_21923);
and UO_597 (O_597,N_22983,N_24105);
xor UO_598 (O_598,N_22642,N_21168);
nand UO_599 (O_599,N_24437,N_22529);
nand UO_600 (O_600,N_23060,N_21769);
or UO_601 (O_601,N_20924,N_24077);
nor UO_602 (O_602,N_21280,N_24412);
or UO_603 (O_603,N_21315,N_23008);
nand UO_604 (O_604,N_24821,N_23934);
and UO_605 (O_605,N_21416,N_20889);
nand UO_606 (O_606,N_20086,N_23868);
or UO_607 (O_607,N_23707,N_23938);
and UO_608 (O_608,N_22518,N_23688);
and UO_609 (O_609,N_23177,N_24245);
nand UO_610 (O_610,N_22946,N_23608);
xor UO_611 (O_611,N_24052,N_24206);
xnor UO_612 (O_612,N_21771,N_24713);
xnor UO_613 (O_613,N_23794,N_21506);
and UO_614 (O_614,N_24866,N_22744);
or UO_615 (O_615,N_24482,N_24954);
or UO_616 (O_616,N_24831,N_22587);
nor UO_617 (O_617,N_22791,N_21011);
and UO_618 (O_618,N_24561,N_21950);
or UO_619 (O_619,N_23542,N_20102);
nand UO_620 (O_620,N_24874,N_20088);
or UO_621 (O_621,N_20208,N_20486);
xor UO_622 (O_622,N_20443,N_21471);
nor UO_623 (O_623,N_22208,N_24545);
nand UO_624 (O_624,N_22717,N_23590);
nor UO_625 (O_625,N_23340,N_20155);
nor UO_626 (O_626,N_24369,N_20704);
or UO_627 (O_627,N_22048,N_20808);
nand UO_628 (O_628,N_22871,N_22997);
nand UO_629 (O_629,N_22155,N_24150);
xor UO_630 (O_630,N_24431,N_24754);
or UO_631 (O_631,N_20403,N_24968);
xor UO_632 (O_632,N_23310,N_22951);
nand UO_633 (O_633,N_23380,N_23120);
and UO_634 (O_634,N_21353,N_21271);
and UO_635 (O_635,N_22582,N_24082);
or UO_636 (O_636,N_23591,N_21606);
nor UO_637 (O_637,N_22651,N_20054);
nor UO_638 (O_638,N_24220,N_23929);
xnor UO_639 (O_639,N_23712,N_22310);
nor UO_640 (O_640,N_23475,N_23602);
and UO_641 (O_641,N_20759,N_22265);
and UO_642 (O_642,N_21004,N_23516);
xor UO_643 (O_643,N_24985,N_22367);
nand UO_644 (O_644,N_22776,N_20655);
or UO_645 (O_645,N_22653,N_22313);
nand UO_646 (O_646,N_24558,N_24013);
nor UO_647 (O_647,N_20552,N_21649);
nor UO_648 (O_648,N_20038,N_22910);
xnor UO_649 (O_649,N_22420,N_24018);
xnor UO_650 (O_650,N_21459,N_20002);
nor UO_651 (O_651,N_20149,N_20025);
nor UO_652 (O_652,N_23969,N_23743);
xnor UO_653 (O_653,N_22437,N_23867);
and UO_654 (O_654,N_22275,N_24172);
or UO_655 (O_655,N_24648,N_22795);
and UO_656 (O_656,N_22272,N_22116);
or UO_657 (O_657,N_21701,N_21614);
and UO_658 (O_658,N_23679,N_23150);
or UO_659 (O_659,N_24670,N_23535);
nand UO_660 (O_660,N_20069,N_24399);
or UO_661 (O_661,N_23089,N_24154);
nand UO_662 (O_662,N_20884,N_24474);
nand UO_663 (O_663,N_20797,N_24321);
nand UO_664 (O_664,N_23359,N_22716);
nand UO_665 (O_665,N_23046,N_24524);
nor UO_666 (O_666,N_20167,N_23607);
nand UO_667 (O_667,N_20168,N_20385);
xnor UO_668 (O_668,N_23321,N_21961);
nand UO_669 (O_669,N_21772,N_22219);
and UO_670 (O_670,N_22977,N_24228);
nor UO_671 (O_671,N_22918,N_23569);
xnor UO_672 (O_672,N_23494,N_22244);
xnor UO_673 (O_673,N_22194,N_20893);
or UO_674 (O_674,N_24423,N_21450);
and UO_675 (O_675,N_21275,N_22445);
and UO_676 (O_676,N_20594,N_23587);
nand UO_677 (O_677,N_23115,N_21920);
or UO_678 (O_678,N_21288,N_22532);
xor UO_679 (O_679,N_22185,N_20389);
nand UO_680 (O_680,N_21757,N_22386);
xor UO_681 (O_681,N_21375,N_20316);
nor UO_682 (O_682,N_21157,N_20566);
xor UO_683 (O_683,N_22635,N_20118);
nand UO_684 (O_684,N_22041,N_20590);
and UO_685 (O_685,N_20131,N_20817);
nor UO_686 (O_686,N_20509,N_24020);
nand UO_687 (O_687,N_22075,N_23490);
nor UO_688 (O_688,N_21042,N_23894);
nor UO_689 (O_689,N_20607,N_20112);
and UO_690 (O_690,N_20300,N_23057);
nand UO_691 (O_691,N_24109,N_24190);
xor UO_692 (O_692,N_20829,N_21632);
nand UO_693 (O_693,N_21161,N_24806);
xor UO_694 (O_694,N_22592,N_23316);
nor UO_695 (O_695,N_23238,N_24213);
nor UO_696 (O_696,N_24297,N_23995);
or UO_697 (O_697,N_24258,N_23353);
and UO_698 (O_698,N_22823,N_23505);
xor UO_699 (O_699,N_22321,N_23296);
or UO_700 (O_700,N_20364,N_23311);
and UO_701 (O_701,N_21395,N_21694);
nand UO_702 (O_702,N_21959,N_24758);
and UO_703 (O_703,N_24185,N_20201);
or UO_704 (O_704,N_23330,N_21006);
xor UO_705 (O_705,N_22473,N_22764);
xnor UO_706 (O_706,N_24936,N_21414);
nand UO_707 (O_707,N_22094,N_23818);
xor UO_708 (O_708,N_22830,N_22669);
nor UO_709 (O_709,N_23042,N_20174);
nor UO_710 (O_710,N_20177,N_22347);
xor UO_711 (O_711,N_20083,N_24618);
nor UO_712 (O_712,N_23885,N_22108);
and UO_713 (O_713,N_21000,N_20440);
and UO_714 (O_714,N_20780,N_22913);
nand UO_715 (O_715,N_22416,N_22881);
xnor UO_716 (O_716,N_22729,N_22798);
or UO_717 (O_717,N_20175,N_20512);
or UO_718 (O_718,N_23249,N_22508);
and UO_719 (O_719,N_23481,N_22531);
or UO_720 (O_720,N_23875,N_20136);
nor UO_721 (O_721,N_22472,N_21558);
nand UO_722 (O_722,N_24844,N_24062);
nand UO_723 (O_723,N_23560,N_21905);
and UO_724 (O_724,N_20923,N_23828);
and UO_725 (O_725,N_22026,N_22982);
nor UO_726 (O_726,N_23181,N_20835);
or UO_727 (O_727,N_21631,N_23533);
and UO_728 (O_728,N_24417,N_24933);
nor UO_729 (O_729,N_23068,N_20888);
and UO_730 (O_730,N_24932,N_22067);
nand UO_731 (O_731,N_22251,N_23155);
or UO_732 (O_732,N_21312,N_24325);
nor UO_733 (O_733,N_24614,N_22737);
nor UO_734 (O_734,N_20447,N_22411);
or UO_735 (O_735,N_21228,N_22301);
nand UO_736 (O_736,N_22117,N_23532);
and UO_737 (O_737,N_22124,N_22693);
nor UO_738 (O_738,N_23086,N_22129);
or UO_739 (O_739,N_23922,N_21095);
and UO_740 (O_740,N_21963,N_20856);
and UO_741 (O_741,N_24882,N_23153);
or UO_742 (O_742,N_22242,N_24203);
nor UO_743 (O_743,N_23074,N_22343);
and UO_744 (O_744,N_20961,N_22096);
nor UO_745 (O_745,N_23615,N_22502);
xor UO_746 (O_746,N_21125,N_20286);
xnor UO_747 (O_747,N_20592,N_24443);
nand UO_748 (O_748,N_21718,N_23192);
xnor UO_749 (O_749,N_21189,N_22953);
or UO_750 (O_750,N_20152,N_23304);
or UO_751 (O_751,N_23004,N_24415);
and UO_752 (O_752,N_24574,N_23661);
nand UO_753 (O_753,N_24718,N_20348);
and UO_754 (O_754,N_23372,N_22721);
and UO_755 (O_755,N_22066,N_23062);
xnor UO_756 (O_756,N_20022,N_21177);
and UO_757 (O_757,N_21753,N_21591);
and UO_758 (O_758,N_20810,N_24659);
and UO_759 (O_759,N_23085,N_24182);
xor UO_760 (O_760,N_20206,N_21419);
and UO_761 (O_761,N_23877,N_24047);
and UO_762 (O_762,N_20188,N_23207);
or UO_763 (O_763,N_21878,N_21648);
and UO_764 (O_764,N_20621,N_24612);
nand UO_765 (O_765,N_20104,N_21872);
and UO_766 (O_766,N_21966,N_24687);
and UO_767 (O_767,N_22996,N_24642);
and UO_768 (O_768,N_22850,N_21225);
and UO_769 (O_769,N_21976,N_20396);
or UO_770 (O_770,N_20374,N_23963);
and UO_771 (O_771,N_23143,N_21100);
nor UO_772 (O_772,N_24451,N_20282);
and UO_773 (O_773,N_24101,N_20013);
and UO_774 (O_774,N_23375,N_22014);
nand UO_775 (O_775,N_21294,N_23409);
xor UO_776 (O_776,N_20071,N_21126);
and UO_777 (O_777,N_20843,N_21695);
or UO_778 (O_778,N_22335,N_22123);
and UO_779 (O_779,N_20193,N_21462);
or UO_780 (O_780,N_21892,N_24767);
nor UO_781 (O_781,N_20365,N_24414);
and UO_782 (O_782,N_20771,N_22566);
nor UO_783 (O_783,N_24619,N_20169);
nand UO_784 (O_784,N_22312,N_21320);
nand UO_785 (O_785,N_20070,N_22083);
xor UO_786 (O_786,N_24029,N_24429);
and UO_787 (O_787,N_23294,N_21543);
or UO_788 (O_788,N_21192,N_20925);
or UO_789 (O_789,N_23741,N_21798);
or UO_790 (O_790,N_22709,N_22329);
or UO_791 (O_791,N_21927,N_21789);
nand UO_792 (O_792,N_22988,N_20255);
nor UO_793 (O_793,N_23165,N_23452);
and UO_794 (O_794,N_22949,N_23352);
nand UO_795 (O_795,N_23078,N_24413);
xnor UO_796 (O_796,N_23093,N_23462);
nor UO_797 (O_797,N_20604,N_22553);
or UO_798 (O_798,N_23151,N_22504);
nand UO_799 (O_799,N_21744,N_20338);
nor UO_800 (O_800,N_24085,N_23443);
nand UO_801 (O_801,N_23625,N_23517);
and UO_802 (O_802,N_22689,N_23648);
or UO_803 (O_803,N_23724,N_23760);
xor UO_804 (O_804,N_24122,N_20532);
xnor UO_805 (O_805,N_21093,N_21891);
and UO_806 (O_806,N_23742,N_20080);
xor UO_807 (O_807,N_23104,N_23302);
nor UO_808 (O_808,N_22054,N_20652);
or UO_809 (O_809,N_24540,N_24269);
and UO_810 (O_810,N_21724,N_20887);
nor UO_811 (O_811,N_20729,N_24575);
nand UO_812 (O_812,N_20933,N_21993);
nand UO_813 (O_813,N_20682,N_22725);
nor UO_814 (O_814,N_22069,N_24598);
and UO_815 (O_815,N_22848,N_24007);
nand UO_816 (O_816,N_24686,N_24992);
nor UO_817 (O_817,N_21911,N_22998);
or UO_818 (O_818,N_21666,N_22188);
nand UO_819 (O_819,N_21595,N_22415);
or UO_820 (O_820,N_22241,N_23121);
and UO_821 (O_821,N_20959,N_22627);
nor UO_822 (O_822,N_20792,N_23847);
nor UO_823 (O_823,N_23986,N_24672);
nand UO_824 (O_824,N_24708,N_21210);
nor UO_825 (O_825,N_23389,N_23217);
or UO_826 (O_826,N_20238,N_22575);
or UO_827 (O_827,N_22789,N_21852);
xor UO_828 (O_828,N_23792,N_24513);
nand UO_829 (O_829,N_21274,N_23399);
nor UO_830 (O_830,N_20409,N_22990);
xnor UO_831 (O_831,N_24117,N_24781);
and UO_832 (O_832,N_23358,N_20192);
xor UO_833 (O_833,N_23933,N_20301);
xor UO_834 (O_834,N_24891,N_24986);
xor UO_835 (O_835,N_21651,N_23703);
and UO_836 (O_836,N_23113,N_21826);
nand UO_837 (O_837,N_24111,N_24401);
nand UO_838 (O_838,N_21854,N_20688);
and UO_839 (O_839,N_20750,N_24250);
nor UO_840 (O_840,N_20227,N_21689);
xor UO_841 (O_841,N_22360,N_24946);
nand UO_842 (O_842,N_24741,N_20528);
nor UO_843 (O_843,N_20261,N_21421);
and UO_844 (O_844,N_23685,N_23034);
and UO_845 (O_845,N_20319,N_21715);
xor UO_846 (O_846,N_24923,N_20821);
xor UO_847 (O_847,N_22471,N_22509);
nor UO_848 (O_848,N_24056,N_24342);
xnor UO_849 (O_849,N_21979,N_21673);
nor UO_850 (O_850,N_24871,N_24218);
nand UO_851 (O_851,N_23147,N_20421);
nand UO_852 (O_852,N_23491,N_20949);
xor UO_853 (O_853,N_24248,N_23864);
xnor UO_854 (O_854,N_21864,N_23571);
nand UO_855 (O_855,N_20209,N_20964);
xnor UO_856 (O_856,N_23900,N_23725);
and UO_857 (O_857,N_22556,N_21109);
nor UO_858 (O_858,N_20583,N_23705);
or UO_859 (O_859,N_22493,N_21456);
nand UO_860 (O_860,N_21945,N_21432);
nand UO_861 (O_861,N_20816,N_22351);
and UO_862 (O_862,N_22886,N_23210);
nor UO_863 (O_863,N_22267,N_24157);
xnor UO_864 (O_864,N_21211,N_20900);
nand UO_865 (O_865,N_24496,N_24271);
nand UO_866 (O_866,N_24097,N_22134);
nor UO_867 (O_867,N_24908,N_21973);
nand UO_868 (O_868,N_24009,N_21101);
nor UO_869 (O_869,N_22520,N_24854);
xnor UO_870 (O_870,N_21994,N_23435);
and UO_871 (O_871,N_22402,N_23736);
xor UO_872 (O_872,N_24599,N_22861);
xor UO_873 (O_873,N_23432,N_24774);
nor UO_874 (O_874,N_22012,N_21064);
nor UO_875 (O_875,N_23904,N_21047);
nor UO_876 (O_876,N_24495,N_21625);
nor UO_877 (O_877,N_20256,N_24953);
and UO_878 (O_878,N_21719,N_21931);
and UO_879 (O_879,N_23118,N_21594);
and UO_880 (O_880,N_20538,N_23019);
nand UO_881 (O_881,N_20585,N_20595);
and UO_882 (O_882,N_23365,N_23772);
and UO_883 (O_883,N_24043,N_20310);
and UO_884 (O_884,N_22022,N_21740);
and UO_885 (O_885,N_20565,N_24810);
and UO_886 (O_886,N_23176,N_20128);
or UO_887 (O_887,N_20815,N_23322);
or UO_888 (O_888,N_24652,N_20903);
and UO_889 (O_889,N_23520,N_23709);
xnor UO_890 (O_890,N_21839,N_21281);
and UO_891 (O_891,N_24494,N_22900);
nand UO_892 (O_892,N_21581,N_21342);
or UO_893 (O_893,N_21639,N_20665);
xnor UO_894 (O_894,N_23175,N_20722);
and UO_895 (O_895,N_23382,N_20564);
or UO_896 (O_896,N_24763,N_22011);
nand UO_897 (O_897,N_23942,N_20844);
and UO_898 (O_898,N_23748,N_20307);
nand UO_899 (O_899,N_20285,N_20030);
nor UO_900 (O_900,N_23738,N_23223);
nand UO_901 (O_901,N_20138,N_22612);
xnor UO_902 (O_902,N_20601,N_21883);
xnor UO_903 (O_903,N_21187,N_21846);
xor UO_904 (O_904,N_20453,N_23033);
or UO_905 (O_905,N_22282,N_22815);
and UO_906 (O_906,N_20620,N_23327);
and UO_907 (O_907,N_24961,N_23983);
or UO_908 (O_908,N_21516,N_21729);
nor UO_909 (O_909,N_23730,N_24184);
nand UO_910 (O_910,N_21377,N_20753);
and UO_911 (O_911,N_21877,N_20569);
nor UO_912 (O_912,N_23281,N_22021);
or UO_913 (O_913,N_22237,N_22832);
or UO_914 (O_914,N_22458,N_22755);
nor UO_915 (O_915,N_24514,N_22835);
nand UO_916 (O_916,N_20738,N_24995);
nand UO_917 (O_917,N_23195,N_20857);
and UO_918 (O_918,N_21561,N_21181);
or UO_919 (O_919,N_20697,N_20720);
nand UO_920 (O_920,N_21909,N_23395);
nand UO_921 (O_921,N_21269,N_22699);
nand UO_922 (O_922,N_22068,N_22454);
nand UO_923 (O_923,N_24677,N_20470);
and UO_924 (O_924,N_21103,N_22833);
xor UO_925 (O_925,N_20415,N_23858);
xor UO_926 (O_926,N_24394,N_24864);
and UO_927 (O_927,N_23681,N_22357);
xor UO_928 (O_928,N_24377,N_21851);
nor UO_929 (O_929,N_20806,N_22107);
and UO_930 (O_930,N_23205,N_21059);
nand UO_931 (O_931,N_20683,N_24354);
nor UO_932 (O_932,N_24357,N_23106);
and UO_933 (O_933,N_22002,N_21351);
nor UO_934 (O_934,N_24119,N_22876);
nor UO_935 (O_935,N_21365,N_22417);
or UO_936 (O_936,N_21710,N_22016);
and UO_937 (O_937,N_21409,N_23383);
nor UO_938 (O_938,N_23144,N_24744);
nor UO_939 (O_939,N_24967,N_21566);
nor UO_940 (O_940,N_23035,N_22234);
or UO_941 (O_941,N_21929,N_22181);
nand UO_942 (O_942,N_22298,N_20773);
nor UO_943 (O_943,N_21489,N_23734);
xnor UO_944 (O_944,N_24232,N_20983);
and UO_945 (O_945,N_22915,N_22727);
nor UO_946 (O_946,N_20495,N_20752);
and UO_947 (O_947,N_20784,N_21553);
and UO_948 (O_948,N_22846,N_20020);
nor UO_949 (O_949,N_24988,N_24699);
and UO_950 (O_950,N_24517,N_22858);
or UO_951 (O_951,N_22485,N_21056);
nand UO_952 (O_952,N_22960,N_24761);
and UO_953 (O_953,N_21699,N_21152);
and UO_954 (O_954,N_20371,N_22133);
nand UO_955 (O_955,N_24445,N_23468);
xor UO_956 (O_956,N_21010,N_23274);
or UO_957 (O_957,N_22200,N_23368);
or UO_958 (O_958,N_23676,N_22954);
and UO_959 (O_959,N_20625,N_24571);
nand UO_960 (O_960,N_24966,N_22191);
and UO_961 (O_961,N_20242,N_20160);
and UO_962 (O_962,N_23918,N_20679);
and UO_963 (O_963,N_24605,N_23756);
or UO_964 (O_964,N_23393,N_20556);
nor UO_965 (O_965,N_22554,N_22001);
and UO_966 (O_966,N_20265,N_22768);
xor UO_967 (O_967,N_21652,N_24634);
nand UO_968 (O_968,N_20342,N_22247);
or UO_969 (O_969,N_24507,N_20935);
or UO_970 (O_970,N_24877,N_24252);
xor UO_971 (O_971,N_20672,N_21403);
nor UO_972 (O_972,N_24929,N_22232);
and UO_973 (O_973,N_21292,N_21887);
and UO_974 (O_974,N_23114,N_23988);
nor UO_975 (O_975,N_20281,N_22374);
and UO_976 (O_976,N_21256,N_22314);
or UO_977 (O_977,N_21965,N_24530);
nor UO_978 (O_978,N_24978,N_20326);
nand UO_979 (O_979,N_23901,N_21521);
or UO_980 (O_980,N_21640,N_23227);
and UO_981 (O_981,N_21030,N_22674);
xnor UO_982 (O_982,N_22702,N_20309);
or UO_983 (O_983,N_20394,N_22976);
and UO_984 (O_984,N_23313,N_21385);
or UO_985 (O_985,N_22238,N_24351);
or UO_986 (O_986,N_21890,N_24483);
xnor UO_987 (O_987,N_24320,N_21308);
nand UO_988 (O_988,N_22922,N_22658);
and UO_989 (O_989,N_21977,N_24977);
xnor UO_990 (O_990,N_21138,N_20799);
xnor UO_991 (O_991,N_22964,N_20619);
nor UO_992 (O_992,N_23949,N_20341);
or UO_993 (O_993,N_22778,N_21948);
xnor UO_994 (O_994,N_21079,N_24584);
nand UO_995 (O_995,N_23655,N_23292);
nor UO_996 (O_996,N_23775,N_22324);
or UO_997 (O_997,N_24594,N_22337);
or UO_998 (O_998,N_20549,N_22028);
or UO_999 (O_999,N_23530,N_21586);
xor UO_1000 (O_1000,N_20687,N_24576);
xor UO_1001 (O_1001,N_23936,N_24775);
xnor UO_1002 (O_1002,N_23687,N_22005);
or UO_1003 (O_1003,N_20770,N_24838);
nand UO_1004 (O_1004,N_20802,N_20377);
nand UO_1005 (O_1005,N_23434,N_21860);
nand UO_1006 (O_1006,N_23202,N_22793);
nand UO_1007 (O_1007,N_21714,N_21402);
xnor UO_1008 (O_1008,N_20503,N_23731);
nand UO_1009 (O_1009,N_21213,N_23506);
nor UO_1010 (O_1010,N_23445,N_20748);
nor UO_1011 (O_1011,N_24755,N_24609);
and UO_1012 (O_1012,N_24032,N_24186);
nand UO_1013 (O_1013,N_24113,N_22671);
or UO_1014 (O_1014,N_21751,N_22955);
xnor UO_1015 (O_1015,N_24355,N_23814);
xor UO_1016 (O_1016,N_21442,N_24161);
and UO_1017 (O_1017,N_23832,N_24406);
xnor UO_1018 (O_1018,N_20696,N_20295);
or UO_1019 (O_1019,N_20508,N_21761);
nor UO_1020 (O_1020,N_23961,N_20111);
xor UO_1021 (O_1021,N_24131,N_24899);
xor UO_1022 (O_1022,N_23908,N_21743);
and UO_1023 (O_1023,N_21672,N_21900);
and UO_1024 (O_1024,N_21117,N_20103);
xor UO_1025 (O_1025,N_20057,N_20116);
and UO_1026 (O_1026,N_23719,N_24853);
xnor UO_1027 (O_1027,N_23059,N_21374);
and UO_1028 (O_1028,N_20011,N_20325);
nor UO_1029 (O_1029,N_21128,N_21243);
and UO_1030 (O_1030,N_24262,N_23618);
or UO_1031 (O_1031,N_21926,N_24765);
nand UO_1032 (O_1032,N_23081,N_23830);
and UO_1033 (O_1033,N_24281,N_22619);
xor UO_1034 (O_1034,N_22945,N_20811);
and UO_1035 (O_1035,N_23978,N_20456);
xnor UO_1036 (O_1036,N_24099,N_24927);
xor UO_1037 (O_1037,N_24552,N_24560);
or UO_1038 (O_1038,N_21230,N_21433);
nor UO_1039 (O_1039,N_24984,N_24895);
xnor UO_1040 (O_1040,N_21250,N_20768);
nand UO_1041 (O_1041,N_24193,N_20205);
or UO_1042 (O_1042,N_22126,N_22777);
nand UO_1043 (O_1043,N_24869,N_20499);
or UO_1044 (O_1044,N_23463,N_24668);
xnor UO_1045 (O_1045,N_24750,N_22073);
or UO_1046 (O_1046,N_21295,N_23643);
xnor UO_1047 (O_1047,N_24408,N_21562);
xor UO_1048 (O_1048,N_20366,N_20463);
and UO_1049 (O_1049,N_23164,N_20049);
or UO_1050 (O_1050,N_23762,N_21787);
and UO_1051 (O_1051,N_23907,N_20761);
and UO_1052 (O_1052,N_21242,N_21249);
nor UO_1053 (O_1053,N_23159,N_23242);
nor UO_1054 (O_1054,N_20663,N_23267);
xnor UO_1055 (O_1055,N_22297,N_22842);
xor UO_1056 (O_1056,N_23955,N_23130);
xor UO_1057 (O_1057,N_21588,N_21115);
nand UO_1058 (O_1058,N_22196,N_22615);
xnor UO_1059 (O_1059,N_24397,N_23459);
nor UO_1060 (O_1060,N_21726,N_23697);
nor UO_1061 (O_1061,N_22088,N_24873);
and UO_1062 (O_1062,N_23786,N_20431);
nand UO_1063 (O_1063,N_24022,N_23966);
and UO_1064 (O_1064,N_22264,N_24335);
and UO_1065 (O_1065,N_24582,N_22080);
nor UO_1066 (O_1066,N_21261,N_24625);
xnor UO_1067 (O_1067,N_23224,N_24794);
xor UO_1068 (O_1068,N_20130,N_21068);
xnor UO_1069 (O_1069,N_22195,N_20638);
nor UO_1070 (O_1070,N_20798,N_20153);
nor UO_1071 (O_1071,N_22634,N_23538);
or UO_1072 (O_1072,N_20513,N_21832);
xnor UO_1073 (O_1073,N_20805,N_21508);
nor UO_1074 (O_1074,N_24479,N_20311);
xor UO_1075 (O_1075,N_22696,N_24426);
and UO_1076 (O_1076,N_23821,N_23225);
nor UO_1077 (O_1077,N_21344,N_22821);
nor UO_1078 (O_1078,N_20637,N_22741);
xnor UO_1079 (O_1079,N_21022,N_23951);
and UO_1080 (O_1080,N_23097,N_22092);
nor UO_1081 (O_1081,N_23243,N_23623);
nand UO_1082 (O_1082,N_20274,N_24380);
nor UO_1083 (O_1083,N_24420,N_22826);
and UO_1084 (O_1084,N_23355,N_21799);
xor UO_1085 (O_1085,N_22081,N_20693);
or UO_1086 (O_1086,N_23450,N_20586);
and UO_1087 (O_1087,N_22573,N_22840);
nor UO_1088 (O_1088,N_22051,N_21944);
xor UO_1089 (O_1089,N_20105,N_24141);
or UO_1090 (O_1090,N_21098,N_23031);
nand UO_1091 (O_1091,N_21236,N_24620);
xor UO_1092 (O_1092,N_22852,N_24809);
or UO_1093 (O_1093,N_23699,N_22724);
nand UO_1094 (O_1094,N_24300,N_20157);
or UO_1095 (O_1095,N_21698,N_23425);
and UO_1096 (O_1096,N_22227,N_22177);
nand UO_1097 (O_1097,N_23427,N_20858);
xnor UO_1098 (O_1098,N_22284,N_21791);
nor UO_1099 (O_1099,N_24799,N_23082);
nor UO_1100 (O_1100,N_21510,N_23277);
or UO_1101 (O_1101,N_20796,N_24590);
xor UO_1102 (O_1102,N_21684,N_22388);
and UO_1103 (O_1103,N_22889,N_21092);
xor UO_1104 (O_1104,N_21647,N_24976);
xnor UO_1105 (O_1105,N_24678,N_23991);
or UO_1106 (O_1106,N_23433,N_20662);
xor UO_1107 (O_1107,N_20598,N_23129);
and UO_1108 (O_1108,N_23419,N_23893);
and UO_1109 (O_1109,N_20150,N_22995);
and UO_1110 (O_1110,N_24069,N_20535);
xor UO_1111 (O_1111,N_21071,N_23616);
xnor UO_1112 (O_1112,N_23092,N_20749);
xnor UO_1113 (O_1113,N_22370,N_22332);
and UO_1114 (O_1114,N_24712,N_24130);
nor UO_1115 (O_1115,N_21014,N_24549);
xnor UO_1116 (O_1116,N_23418,N_21327);
nor UO_1117 (O_1117,N_21132,N_20418);
and UO_1118 (O_1118,N_23158,N_20636);
and UO_1119 (O_1119,N_24363,N_21940);
or UO_1120 (O_1120,N_20220,N_20941);
xnor UO_1121 (O_1121,N_21319,N_22236);
nand UO_1122 (O_1122,N_22045,N_20346);
or UO_1123 (O_1123,N_23583,N_23905);
or UO_1124 (O_1124,N_24912,N_20730);
nand UO_1125 (O_1125,N_23087,N_21665);
and UO_1126 (O_1126,N_22391,N_21457);
nor UO_1127 (O_1127,N_20246,N_21759);
and UO_1128 (O_1128,N_22400,N_20984);
xnor UO_1129 (O_1129,N_20591,N_23600);
or UO_1130 (O_1130,N_22348,N_23333);
nand UO_1131 (O_1131,N_20189,N_20596);
xor UO_1132 (O_1132,N_24034,N_20998);
nand UO_1133 (O_1133,N_21412,N_21568);
nor UO_1134 (O_1134,N_24795,N_22901);
nand UO_1135 (O_1135,N_20548,N_22269);
and UO_1136 (O_1136,N_21195,N_20834);
or UO_1137 (O_1137,N_21745,N_20747);
xor UO_1138 (O_1138,N_21384,N_24003);
or UO_1139 (O_1139,N_23789,N_22175);
xnor UO_1140 (O_1140,N_22817,N_24035);
xor UO_1141 (O_1141,N_24835,N_24216);
or UO_1142 (O_1142,N_20124,N_24187);
or UO_1143 (O_1143,N_24447,N_21313);
xor UO_1144 (O_1144,N_22515,N_21360);
nor UO_1145 (O_1145,N_20629,N_23429);
nor UO_1146 (O_1146,N_21448,N_21264);
nand UO_1147 (O_1147,N_24002,N_21917);
and UO_1148 (O_1148,N_22033,N_20536);
or UO_1149 (O_1149,N_20741,N_24164);
and UO_1150 (O_1150,N_21995,N_23376);
and UO_1151 (O_1151,N_20191,N_24310);
and UO_1152 (O_1152,N_24945,N_20452);
xor UO_1153 (O_1153,N_24705,N_22132);
nor UO_1154 (O_1154,N_21055,N_23307);
nand UO_1155 (O_1155,N_21836,N_20401);
and UO_1156 (O_1156,N_21038,N_23633);
xor UO_1157 (O_1157,N_23122,N_24110);
or UO_1158 (O_1158,N_20228,N_23799);
and UO_1159 (O_1159,N_20000,N_22865);
nand UO_1160 (O_1160,N_21593,N_22250);
nor UO_1161 (O_1161,N_24726,N_20391);
nor UO_1162 (O_1162,N_20731,N_23025);
or UO_1163 (O_1163,N_23172,N_23456);
xor UO_1164 (O_1164,N_23752,N_20758);
and UO_1165 (O_1165,N_23478,N_24277);
or UO_1166 (O_1166,N_23032,N_23722);
nand UO_1167 (O_1167,N_22311,N_24438);
nor UO_1168 (O_1168,N_22974,N_20166);
xor UO_1169 (O_1169,N_22723,N_22705);
or UO_1170 (O_1170,N_24244,N_23385);
nor UO_1171 (O_1171,N_24464,N_24497);
xor UO_1172 (O_1172,N_22266,N_21970);
nand UO_1173 (O_1173,N_24704,N_22137);
xnor UO_1174 (O_1174,N_23498,N_23582);
or UO_1175 (O_1175,N_23254,N_20197);
and UO_1176 (O_1176,N_21609,N_20240);
or UO_1177 (O_1177,N_23234,N_23559);
and UO_1178 (O_1178,N_21337,N_22142);
and UO_1179 (O_1179,N_24292,N_23184);
nor UO_1180 (O_1180,N_20940,N_21635);
nor UO_1181 (O_1181,N_21464,N_23693);
nor UO_1182 (O_1182,N_20718,N_22439);
or UO_1183 (O_1183,N_24604,N_23993);
and UO_1184 (O_1184,N_21686,N_20257);
and UO_1185 (O_1185,N_21306,N_23902);
and UO_1186 (O_1186,N_21345,N_21616);
xor UO_1187 (O_1187,N_23898,N_23056);
or UO_1188 (O_1188,N_20165,N_21741);
nand UO_1189 (O_1189,N_23512,N_22883);
and UO_1190 (O_1190,N_22766,N_23013);
nand UO_1191 (O_1191,N_20042,N_24787);
nand UO_1192 (O_1192,N_21113,N_24613);
nand UO_1193 (O_1193,N_22252,N_24226);
nor UO_1194 (O_1194,N_21933,N_23630);
or UO_1195 (O_1195,N_21660,N_21468);
and UO_1196 (O_1196,N_23212,N_20065);
nand UO_1197 (O_1197,N_22747,N_21867);
or UO_1198 (O_1198,N_24080,N_22379);
nand UO_1199 (O_1199,N_20627,N_23573);
xnor UO_1200 (O_1200,N_24816,N_21324);
nor UO_1201 (O_1201,N_23840,N_22816);
and UO_1202 (O_1202,N_21358,N_21378);
nand UO_1203 (O_1203,N_21982,N_22563);
nor UO_1204 (O_1204,N_22448,N_20425);
or UO_1205 (O_1205,N_22205,N_22498);
or UO_1206 (O_1206,N_23599,N_22524);
xnor UO_1207 (O_1207,N_24234,N_21777);
nor UO_1208 (O_1208,N_22923,N_21144);
and UO_1209 (O_1209,N_23634,N_23323);
or UO_1210 (O_1210,N_21907,N_20489);
nand UO_1211 (O_1211,N_23824,N_24264);
nand UO_1212 (O_1212,N_20997,N_23924);
and UO_1213 (O_1213,N_22535,N_20245);
nand UO_1214 (O_1214,N_21440,N_20694);
or UO_1215 (O_1215,N_23319,N_21942);
xor UO_1216 (O_1216,N_23764,N_21309);
or UO_1217 (O_1217,N_23309,N_20711);
and UO_1218 (O_1218,N_23774,N_21658);
nor UO_1219 (O_1219,N_22253,N_23959);
nand UO_1220 (O_1220,N_24491,N_20950);
xnor UO_1221 (O_1221,N_20986,N_24856);
xnor UO_1222 (O_1222,N_21902,N_20624);
xor UO_1223 (O_1223,N_23226,N_21774);
or UO_1224 (O_1224,N_20912,N_23716);
nand UO_1225 (O_1225,N_22434,N_23531);
nor UO_1226 (O_1226,N_21204,N_23384);
xor UO_1227 (O_1227,N_22024,N_20404);
nor UO_1228 (O_1228,N_22125,N_21597);
nor UO_1229 (O_1229,N_20270,N_20058);
or UO_1230 (O_1230,N_22663,N_20567);
and UO_1231 (O_1231,N_24459,N_22299);
xnor UO_1232 (O_1232,N_23017,N_20842);
nor UO_1233 (O_1233,N_20777,N_23220);
and UO_1234 (O_1234,N_20520,N_21287);
nor UO_1235 (O_1235,N_22334,N_22944);
xnor UO_1236 (O_1236,N_24146,N_20059);
nor UO_1237 (O_1237,N_21830,N_20367);
and UO_1238 (O_1238,N_20076,N_22259);
and UO_1239 (O_1239,N_24752,N_24897);
xnor UO_1240 (O_1240,N_22576,N_24090);
nand UO_1241 (O_1241,N_23788,N_24753);
or UO_1242 (O_1242,N_23639,N_20560);
nand UO_1243 (O_1243,N_22303,N_22221);
nor UO_1244 (O_1244,N_22279,N_21585);
nor UO_1245 (O_1245,N_20357,N_21974);
nand UO_1246 (O_1246,N_22316,N_24481);
xor UO_1247 (O_1247,N_24888,N_23603);
or UO_1248 (O_1248,N_21599,N_23529);
nor UO_1249 (O_1249,N_20504,N_20380);
nand UO_1250 (O_1250,N_20827,N_21584);
or UO_1251 (O_1251,N_20034,N_24382);
and UO_1252 (O_1252,N_21392,N_24011);
and UO_1253 (O_1253,N_23064,N_24166);
nand UO_1254 (O_1254,N_24044,N_24739);
xor UO_1255 (O_1255,N_20252,N_24942);
nand UO_1256 (O_1256,N_20995,N_21367);
xor UO_1257 (O_1257,N_22989,N_21677);
nand UO_1258 (O_1258,N_24365,N_24635);
nor UO_1259 (O_1259,N_21990,N_23525);
or UO_1260 (O_1260,N_20873,N_23486);
xnor UO_1261 (O_1261,N_20483,N_24641);
nand UO_1262 (O_1262,N_23049,N_21058);
xnor UO_1263 (O_1263,N_24681,N_24896);
or UO_1264 (O_1264,N_21018,N_23127);
nor UO_1265 (O_1265,N_23152,N_22552);
and UO_1266 (O_1266,N_24211,N_21853);
nand UO_1267 (O_1267,N_21233,N_20505);
nor UO_1268 (O_1268,N_23048,N_23842);
and UO_1269 (O_1269,N_21223,N_22152);
or UO_1270 (O_1270,N_20809,N_20530);
nand UO_1271 (O_1271,N_22571,N_21559);
or UO_1272 (O_1272,N_21576,N_23678);
xor UO_1273 (O_1273,N_22893,N_24485);
or UO_1274 (O_1274,N_23769,N_24606);
xnor UO_1275 (O_1275,N_20212,N_21185);
nand UO_1276 (O_1276,N_23258,N_21257);
and UO_1277 (O_1277,N_21782,N_20721);
xnor UO_1278 (O_1278,N_23662,N_21484);
nand UO_1279 (O_1279,N_24012,N_23737);
nand UO_1280 (O_1280,N_22533,N_24654);
and UO_1281 (O_1281,N_23485,N_21277);
and UO_1282 (O_1282,N_23257,N_22596);
and UO_1283 (O_1283,N_20321,N_21869);
xnor UO_1284 (O_1284,N_20047,N_22030);
nor UO_1285 (O_1285,N_23493,N_23105);
nand UO_1286 (O_1286,N_24124,N_22897);
nand UO_1287 (O_1287,N_21831,N_24863);
nand UO_1288 (O_1288,N_20492,N_24706);
nand UO_1289 (O_1289,N_21086,N_24194);
nand UO_1290 (O_1290,N_24151,N_23408);
nor UO_1291 (O_1291,N_21598,N_20932);
and UO_1292 (O_1292,N_23541,N_20710);
xor UO_1293 (O_1293,N_22151,N_24108);
and UO_1294 (O_1294,N_23674,N_22463);
or UO_1295 (O_1295,N_22204,N_20315);
nand UO_1296 (O_1296,N_23222,N_24033);
and UO_1297 (O_1297,N_21554,N_24532);
nand UO_1298 (O_1298,N_21214,N_21564);
and UO_1299 (O_1299,N_21897,N_22230);
nor UO_1300 (O_1300,N_21502,N_24427);
nand UO_1301 (O_1301,N_20479,N_23241);
and UO_1302 (O_1302,N_24521,N_22243);
xnor UO_1303 (O_1303,N_21343,N_23967);
nand UO_1304 (O_1304,N_21073,N_20960);
or UO_1305 (O_1305,N_22063,N_22775);
or UO_1306 (O_1306,N_24197,N_21238);
xnor UO_1307 (O_1307,N_21602,N_22879);
and UO_1308 (O_1308,N_22387,N_24910);
nand UO_1309 (O_1309,N_21524,N_23636);
and UO_1310 (O_1310,N_24636,N_21222);
nor UO_1311 (O_1311,N_24435,N_21748);
or UO_1312 (O_1312,N_20502,N_21803);
nand UO_1313 (O_1313,N_24167,N_24370);
and UO_1314 (O_1314,N_22003,N_23985);
nor UO_1315 (O_1315,N_23317,N_23170);
nand UO_1316 (O_1316,N_22084,N_21997);
or UO_1317 (O_1317,N_23026,N_23870);
nor UO_1318 (O_1318,N_22368,N_22811);
or UO_1319 (O_1319,N_23464,N_21498);
nor UO_1320 (O_1320,N_23518,N_20599);
xnor UO_1321 (O_1321,N_23664,N_23848);
or UO_1322 (O_1322,N_21925,N_20523);
and UO_1323 (O_1323,N_23141,N_21988);
and UO_1324 (O_1324,N_24568,N_24265);
and UO_1325 (O_1325,N_20653,N_20198);
nor UO_1326 (O_1326,N_22655,N_21624);
nor UO_1327 (O_1327,N_20626,N_22746);
nor UO_1328 (O_1328,N_21547,N_23827);
nand UO_1329 (O_1329,N_24796,N_24156);
or UO_1330 (O_1330,N_24461,N_24028);
nand UO_1331 (O_1331,N_20823,N_23968);
and UO_1332 (O_1332,N_23523,N_24777);
nand UO_1333 (O_1333,N_21346,N_23109);
and UO_1334 (O_1334,N_22166,N_21091);
or UO_1335 (O_1335,N_24617,N_23751);
or UO_1336 (O_1336,N_21182,N_22224);
or UO_1337 (O_1337,N_21482,N_23865);
xnor UO_1338 (O_1338,N_21379,N_23854);
and UO_1339 (O_1339,N_23128,N_21332);
and UO_1340 (O_1340,N_21857,N_22868);
nand UO_1341 (O_1341,N_24504,N_22176);
nand UO_1342 (O_1342,N_24424,N_20501);
xor UO_1343 (O_1343,N_20954,N_21036);
xor UO_1344 (O_1344,N_22749,N_21099);
nor UO_1345 (O_1345,N_24091,N_20028);
nor UO_1346 (O_1346,N_24345,N_20993);
xnor UO_1347 (O_1347,N_23439,N_23747);
and UO_1348 (O_1348,N_23585,N_20669);
or UO_1349 (O_1349,N_24058,N_24764);
or UO_1350 (O_1350,N_20994,N_22838);
and UO_1351 (O_1351,N_22156,N_20728);
or UO_1352 (O_1352,N_20992,N_20018);
xor UO_1353 (O_1353,N_23823,N_24973);
nor UO_1354 (O_1354,N_22661,N_21080);
and UO_1355 (O_1355,N_20689,N_20045);
or UO_1356 (O_1356,N_22547,N_22589);
and UO_1357 (O_1357,N_22593,N_22825);
or UO_1358 (O_1358,N_20957,N_23364);
and UO_1359 (O_1359,N_24103,N_24407);
or UO_1360 (O_1360,N_21215,N_23324);
xnor UO_1361 (O_1361,N_22431,N_21339);
nor UO_1362 (O_1362,N_22199,N_24316);
nor UO_1363 (O_1363,N_23345,N_21205);
nand UO_1364 (O_1364,N_21143,N_21108);
and UO_1365 (O_1365,N_21159,N_20547);
and UO_1366 (O_1366,N_21682,N_23946);
nand UO_1367 (O_1367,N_22198,N_21284);
xor UO_1368 (O_1368,N_20010,N_24332);
nand UO_1369 (O_1369,N_21296,N_21837);
xor UO_1370 (O_1370,N_20782,N_24930);
nand UO_1371 (O_1371,N_24849,N_24314);
nand UO_1372 (O_1372,N_22047,N_21735);
and UO_1373 (O_1373,N_22044,N_24087);
nor UO_1374 (O_1374,N_24997,N_24516);
nand UO_1375 (O_1375,N_20801,N_22469);
or UO_1376 (O_1376,N_23251,N_21871);
or UO_1377 (O_1377,N_20337,N_22489);
xor UO_1378 (O_1378,N_20195,N_23916);
xnor UO_1379 (O_1379,N_21626,N_23256);
nor UO_1380 (O_1380,N_24465,N_23915);
nand UO_1381 (O_1381,N_23975,N_23629);
nand UO_1382 (O_1382,N_20400,N_22683);
xor UO_1383 (O_1383,N_21444,N_22186);
nor UO_1384 (O_1384,N_20467,N_22864);
and UO_1385 (O_1385,N_23390,N_21971);
nor UO_1386 (O_1386,N_24019,N_20332);
or UO_1387 (O_1387,N_23067,N_23400);
or UO_1388 (O_1388,N_22056,N_23917);
and UO_1389 (O_1389,N_20739,N_20724);
nor UO_1390 (O_1390,N_24135,N_24747);
nor UO_1391 (O_1391,N_24723,N_21876);
and UO_1392 (O_1392,N_20476,N_21956);
nand UO_1393 (O_1393,N_20544,N_21184);
or UO_1394 (O_1394,N_23239,N_21657);
nand UO_1395 (O_1395,N_24569,N_20420);
or UO_1396 (O_1396,N_23029,N_20649);
nor UO_1397 (O_1397,N_24987,N_24862);
or UO_1398 (O_1398,N_23273,N_20826);
and UO_1399 (O_1399,N_23420,N_22564);
or UO_1400 (O_1400,N_20895,N_21387);
or UO_1401 (O_1401,N_22522,N_23700);
or UO_1402 (O_1402,N_22943,N_23992);
xnor UO_1403 (O_1403,N_24691,N_22614);
xor UO_1404 (O_1404,N_20751,N_20477);
xnor UO_1405 (O_1405,N_23671,N_20474);
nor UO_1406 (O_1406,N_23080,N_22013);
and UO_1407 (O_1407,N_20386,N_23605);
and UO_1408 (O_1408,N_22698,N_21496);
and UO_1409 (O_1409,N_24336,N_21850);
and UO_1410 (O_1410,N_22034,N_21263);
or UO_1411 (O_1411,N_23581,N_20735);
nand UO_1412 (O_1412,N_21286,N_20493);
xnor UO_1413 (O_1413,N_20032,N_21169);
or UO_1414 (O_1414,N_20186,N_22739);
and UO_1415 (O_1415,N_20021,N_23421);
nand UO_1416 (O_1416,N_20775,N_21130);
xnor UO_1417 (O_1417,N_22130,N_24046);
and UO_1418 (O_1418,N_24823,N_20635);
nor UO_1419 (O_1419,N_20259,N_21611);
and UO_1420 (O_1420,N_24748,N_20529);
and UO_1421 (O_1421,N_21301,N_23812);
nand UO_1422 (O_1422,N_22623,N_20671);
and UO_1423 (O_1423,N_24279,N_24364);
and UO_1424 (O_1424,N_21057,N_20859);
or UO_1425 (O_1425,N_22276,N_21636);
and UO_1426 (O_1426,N_20686,N_24350);
xnor UO_1427 (O_1427,N_23023,N_24221);
or UO_1428 (O_1428,N_22103,N_22141);
xnor UO_1429 (O_1429,N_23228,N_24655);
or UO_1430 (O_1430,N_21304,N_22959);
nor UO_1431 (O_1431,N_20314,N_20393);
and UO_1432 (O_1432,N_24732,N_23131);
or UO_1433 (O_1433,N_20988,N_20412);
xor UO_1434 (O_1434,N_21952,N_21105);
and UO_1435 (O_1435,N_22371,N_21697);
xnor UO_1436 (O_1436,N_23981,N_21984);
and UO_1437 (O_1437,N_20557,N_24958);
nand UO_1438 (O_1438,N_24142,N_24039);
xor UO_1439 (O_1439,N_20145,N_23378);
nand UO_1440 (O_1440,N_22300,N_21633);
xnor UO_1441 (O_1441,N_20705,N_22182);
or UO_1442 (O_1442,N_20247,N_20094);
or UO_1443 (O_1443,N_24313,N_23510);
nand UO_1444 (O_1444,N_21865,N_20050);
nand UO_1445 (O_1445,N_23036,N_22738);
and UO_1446 (O_1446,N_23148,N_24645);
nor UO_1447 (O_1447,N_23811,N_23444);
or UO_1448 (O_1448,N_21555,N_21070);
nor UO_1449 (O_1449,N_21814,N_21515);
nand UO_1450 (O_1450,N_21404,N_24205);
nor UO_1451 (O_1451,N_20909,N_21511);
nand UO_1452 (O_1452,N_20871,N_23691);
and UO_1453 (O_1453,N_21628,N_22687);
nand UO_1454 (O_1454,N_21713,N_24537);
and UO_1455 (O_1455,N_24850,N_22787);
or UO_1456 (O_1456,N_23230,N_24489);
or UO_1457 (O_1457,N_22506,N_21044);
nor UO_1458 (O_1458,N_21298,N_21721);
nor UO_1459 (O_1459,N_20125,N_20684);
and UO_1460 (O_1460,N_22390,N_20763);
or UO_1461 (O_1461,N_21717,N_22106);
or UO_1462 (O_1462,N_20644,N_22754);
or UO_1463 (O_1463,N_22621,N_23338);
nand UO_1464 (O_1464,N_24883,N_22218);
or UO_1465 (O_1465,N_22344,N_24267);
or UO_1466 (O_1466,N_20468,N_21967);
nand UO_1467 (O_1467,N_20855,N_22248);
and UO_1468 (O_1468,N_23921,N_22769);
and UO_1469 (O_1469,N_23320,N_24602);
xor UO_1470 (O_1470,N_21968,N_21941);
nand UO_1471 (O_1471,N_24975,N_21165);
nor UO_1472 (O_1472,N_22342,N_22975);
nand UO_1473 (O_1473,N_21335,N_21838);
or UO_1474 (O_1474,N_24914,N_20602);
nor UO_1475 (O_1475,N_20490,N_20623);
and UO_1476 (O_1476,N_22444,N_21870);
nor UO_1477 (O_1477,N_24073,N_22740);
nor UO_1478 (O_1478,N_23561,N_23740);
nand UO_1479 (O_1479,N_20853,N_22039);
and UO_1480 (O_1480,N_21494,N_20151);
or UO_1481 (O_1481,N_20134,N_23926);
nor UO_1482 (O_1482,N_24319,N_22931);
nor UO_1483 (O_1483,N_23555,N_23606);
and UO_1484 (O_1484,N_23776,N_20896);
or UO_1485 (O_1485,N_24876,N_20378);
nand UO_1486 (O_1486,N_22468,N_24926);
and UO_1487 (O_1487,N_21915,N_22710);
xnor UO_1488 (O_1488,N_22670,N_21668);
nand UO_1489 (O_1489,N_23770,N_21912);
xnor UO_1490 (O_1490,N_21077,N_21475);
or UO_1491 (O_1491,N_20936,N_24980);
nand UO_1492 (O_1492,N_21991,N_24680);
xnor UO_1493 (O_1493,N_22796,N_20814);
xnor UO_1494 (O_1494,N_24246,N_24017);
nand UO_1495 (O_1495,N_24329,N_24383);
or UO_1496 (O_1496,N_24881,N_21938);
nor UO_1497 (O_1497,N_21654,N_23841);
xnor UO_1498 (O_1498,N_20846,N_23807);
and UO_1499 (O_1499,N_20302,N_21935);
xnor UO_1500 (O_1500,N_24230,N_23554);
and UO_1501 (O_1501,N_23965,N_22260);
and UO_1502 (O_1502,N_23079,N_20014);
nor UO_1503 (O_1503,N_24759,N_23407);
and UO_1504 (O_1504,N_24285,N_20987);
xnor UO_1505 (O_1505,N_24274,N_22928);
xnor UO_1506 (O_1506,N_23910,N_24841);
xnor UO_1507 (O_1507,N_23568,N_22369);
or UO_1508 (O_1508,N_22169,N_23213);
and UO_1509 (O_1509,N_24998,N_23250);
nand UO_1510 (O_1510,N_22880,N_24027);
nand UO_1511 (O_1511,N_24467,N_23293);
or UO_1512 (O_1512,N_20875,N_24261);
or UO_1513 (O_1513,N_23930,N_23300);
nor UO_1514 (O_1514,N_20410,N_24374);
or UO_1515 (O_1515,N_21102,N_21536);
nor UO_1516 (O_1516,N_23088,N_22394);
nor UO_1517 (O_1517,N_23116,N_20129);
nor UO_1518 (O_1518,N_20526,N_20727);
and UO_1519 (O_1519,N_20947,N_24757);
nor UO_1520 (O_1520,N_24440,N_23404);
nand UO_1521 (O_1521,N_20647,N_24189);
xnor UO_1522 (O_1522,N_24917,N_21051);
and UO_1523 (O_1523,N_24536,N_20133);
nand UO_1524 (O_1524,N_20225,N_21678);
nand UO_1525 (O_1525,N_21218,N_22867);
and UO_1526 (O_1526,N_24826,N_20106);
and UO_1527 (O_1527,N_21532,N_22162);
or UO_1528 (O_1528,N_23534,N_20634);
xor UO_1529 (O_1529,N_20894,N_21693);
nor UO_1530 (O_1530,N_23168,N_24798);
and UO_1531 (O_1531,N_24805,N_20719);
nor UO_1532 (O_1532,N_22613,N_20956);
xnor UO_1533 (O_1533,N_22616,N_20543);
and UO_1534 (O_1534,N_20445,N_23396);
nand UO_1535 (O_1535,N_21731,N_24511);
or UO_1536 (O_1536,N_23562,N_20052);
or UO_1537 (O_1537,N_22667,N_21201);
or UO_1538 (O_1538,N_22507,N_23862);
or UO_1539 (O_1539,N_21460,N_21336);
nor UO_1540 (O_1540,N_22010,N_22647);
and UO_1541 (O_1541,N_22836,N_23972);
xnor UO_1542 (O_1542,N_24525,N_20628);
xnor UO_1543 (O_1543,N_24868,N_24671);
nand UO_1544 (O_1544,N_24651,N_21341);
or UO_1545 (O_1545,N_20334,N_21076);
and UO_1546 (O_1546,N_20387,N_24219);
xnor UO_1547 (O_1547,N_22135,N_22053);
or UO_1548 (O_1548,N_24884,N_20918);
and UO_1549 (O_1549,N_24273,N_24478);
nand UO_1550 (O_1550,N_24432,N_20978);
and UO_1551 (O_1551,N_24253,N_20531);
nor UO_1552 (O_1552,N_20788,N_24419);
or UO_1553 (O_1553,N_21513,N_20043);
or UO_1554 (O_1554,N_24400,N_21736);
xor UO_1555 (O_1555,N_24890,N_21398);
or UO_1556 (O_1556,N_23357,N_21390);
or UO_1557 (O_1557,N_20919,N_23480);
nand UO_1558 (O_1558,N_23194,N_20522);
or UO_1559 (O_1559,N_21552,N_23502);
nand UO_1560 (O_1560,N_24557,N_20408);
or UO_1561 (O_1561,N_21252,N_20361);
xnor UO_1562 (O_1562,N_23816,N_24421);
nand UO_1563 (O_1563,N_20906,N_24913);
xor UO_1564 (O_1564,N_21066,N_20772);
nand UO_1565 (O_1565,N_24092,N_23714);
nand UO_1566 (O_1566,N_20176,N_24692);
and UO_1567 (O_1567,N_24788,N_20969);
xor UO_1568 (O_1568,N_22903,N_22578);
and UO_1569 (O_1569,N_22781,N_21784);
nor UO_1570 (O_1570,N_24623,N_21420);
nand UO_1571 (O_1571,N_23063,N_24886);
or UO_1572 (O_1572,N_24843,N_23683);
or UO_1573 (O_1573,N_20178,N_24473);
nor UO_1574 (O_1574,N_23024,N_23706);
nand UO_1575 (O_1575,N_20497,N_24969);
nand UO_1576 (O_1576,N_20881,N_23476);
or UO_1577 (O_1577,N_20580,N_24255);
nand UO_1578 (O_1578,N_23813,N_24834);
and UO_1579 (O_1579,N_23075,N_20945);
and UO_1580 (O_1580,N_22158,N_22383);
nand UO_1581 (O_1581,N_24241,N_24306);
or UO_1582 (O_1582,N_23186,N_24304);
xor UO_1583 (O_1583,N_23461,N_23276);
nand UO_1584 (O_1584,N_24526,N_23974);
nand UO_1585 (O_1585,N_22419,N_22790);
nor UO_1586 (O_1586,N_22268,N_22971);
nand UO_1587 (O_1587,N_23960,N_22697);
nor UO_1588 (O_1588,N_23253,N_24660);
and UO_1589 (O_1589,N_24711,N_20942);
nand UO_1590 (O_1590,N_21372,N_20803);
and UO_1591 (O_1591,N_24935,N_24527);
nand UO_1592 (O_1592,N_23612,N_21525);
nand UO_1593 (O_1593,N_23755,N_22491);
nand UO_1594 (O_1594,N_21134,N_22919);
nand UO_1595 (O_1595,N_20164,N_20056);
nand UO_1596 (O_1596,N_22157,N_23984);
xnor UO_1597 (O_1597,N_21629,N_21574);
nor UO_1598 (O_1598,N_20221,N_23680);
nor UO_1599 (O_1599,N_20432,N_23632);
nand UO_1600 (O_1600,N_22837,N_22834);
nand UO_1601 (O_1601,N_21879,N_24965);
xor UO_1602 (O_1602,N_23593,N_24963);
xor UO_1603 (O_1603,N_24878,N_21557);
nor UO_1604 (O_1604,N_20296,N_21107);
nand UO_1605 (O_1605,N_23500,N_23690);
and UO_1606 (O_1606,N_21507,N_24177);
or UO_1607 (O_1607,N_21874,N_22894);
nand UO_1608 (O_1608,N_22427,N_24867);
and UO_1609 (O_1609,N_23173,N_23932);
nor UO_1610 (O_1610,N_21539,N_20280);
nand UO_1611 (O_1611,N_24934,N_21245);
xnor UO_1612 (O_1612,N_22061,N_22599);
nand UO_1613 (O_1613,N_21198,N_22187);
or UO_1614 (O_1614,N_23628,N_23784);
and UO_1615 (O_1615,N_24746,N_22354);
xor UO_1616 (O_1616,N_24784,N_22082);
or UO_1617 (O_1617,N_23005,N_21259);
nand UO_1618 (O_1618,N_21888,N_22941);
xnor UO_1619 (O_1619,N_21807,N_20437);
xnor UO_1620 (O_1620,N_20135,N_22521);
or UO_1621 (O_1621,N_23206,N_22070);
nor UO_1622 (O_1622,N_21413,N_24477);
and UO_1623 (O_1623,N_20090,N_22389);
nor UO_1624 (O_1624,N_21146,N_24388);
and UO_1625 (O_1625,N_24284,N_22211);
nor UO_1626 (O_1626,N_21908,N_24824);
or UO_1627 (O_1627,N_24565,N_20214);
or UO_1628 (O_1628,N_20216,N_23574);
and UO_1629 (O_1629,N_24249,N_20141);
nor UO_1630 (O_1630,N_23954,N_23896);
and UO_1631 (O_1631,N_22121,N_22308);
and UO_1632 (O_1632,N_24716,N_21397);
xor UO_1633 (O_1633,N_23675,N_20215);
and UO_1634 (O_1634,N_20863,N_21859);
nor UO_1635 (O_1635,N_21700,N_23335);
nand UO_1636 (O_1636,N_24948,N_20276);
nand UO_1637 (O_1637,N_22921,N_20464);
xor UO_1638 (O_1638,N_23287,N_22972);
xnor UO_1639 (O_1639,N_24214,N_24827);
xor UO_1640 (O_1640,N_23037,N_23826);
or UO_1641 (O_1641,N_20958,N_20423);
nor UO_1642 (O_1642,N_22000,N_23793);
or UO_1643 (O_1643,N_20774,N_22501);
nor UO_1644 (O_1644,N_21112,N_21427);
or UO_1645 (O_1645,N_21096,N_23430);
nor UO_1646 (O_1646,N_21209,N_21992);
nor UO_1647 (O_1647,N_24428,N_20485);
or UO_1648 (O_1648,N_24828,N_21896);
nor UO_1649 (O_1649,N_23698,N_22572);
nand UO_1650 (O_1650,N_21716,N_21972);
and UO_1651 (O_1651,N_24298,N_23937);
xnor UO_1652 (O_1652,N_21268,N_24944);
or UO_1653 (O_1653,N_22601,N_23040);
and UO_1654 (O_1654,N_21354,N_21258);
xnor UO_1655 (O_1655,N_22168,N_20449);
and UO_1656 (O_1656,N_20551,N_23211);
and UO_1657 (O_1657,N_24603,N_22018);
and UO_1658 (O_1658,N_23240,N_21834);
xor UO_1659 (O_1659,N_20661,N_24343);
xor UO_1660 (O_1660,N_20182,N_23883);
nor UO_1661 (O_1661,N_20862,N_20035);
and UO_1662 (O_1662,N_23264,N_24633);
xor UO_1663 (O_1663,N_23771,N_22036);
nand UO_1664 (O_1664,N_20142,N_21399);
nor UO_1665 (O_1665,N_20902,N_24053);
nor UO_1666 (O_1666,N_20740,N_20920);
nand UO_1667 (O_1667,N_20472,N_22451);
and UO_1668 (O_1668,N_20331,N_22512);
nand UO_1669 (O_1669,N_21685,N_24409);
nor UO_1670 (O_1670,N_20036,N_21328);
nor UO_1671 (O_1671,N_21550,N_24037);
nand UO_1672 (O_1672,N_22478,N_23604);
and UO_1673 (O_1673,N_21645,N_23140);
or UO_1674 (O_1674,N_24050,N_21541);
or UO_1675 (O_1675,N_24922,N_21321);
nor UO_1676 (O_1676,N_23647,N_24040);
nand UO_1677 (O_1677,N_21361,N_21866);
or UO_1678 (O_1678,N_22662,N_22353);
and UO_1679 (O_1679,N_20640,N_23190);
xor UO_1680 (O_1680,N_24646,N_20600);
and UO_1681 (O_1681,N_23548,N_24042);
and UO_1682 (O_1682,N_24703,N_23214);
nor UO_1683 (O_1683,N_20521,N_22779);
and UO_1684 (O_1684,N_21347,N_20099);
xor UO_1685 (O_1685,N_20262,N_24315);
and UO_1686 (O_1686,N_24771,N_24662);
nor UO_1687 (O_1687,N_24179,N_23939);
or UO_1688 (O_1688,N_24529,N_24359);
nor UO_1689 (O_1689,N_22202,N_23488);
xnor UO_1690 (O_1690,N_22430,N_23346);
or UO_1691 (O_1691,N_24889,N_22222);
nand UO_1692 (O_1692,N_20550,N_21061);
xor UO_1693 (O_1693,N_24153,N_24171);
nand UO_1694 (O_1694,N_21383,N_22820);
or UO_1695 (O_1695,N_23474,N_20703);
xor UO_1696 (O_1696,N_22170,N_22706);
or UO_1697 (O_1697,N_24173,N_23179);
xnor UO_1698 (O_1698,N_24640,N_21590);
or UO_1699 (O_1699,N_24921,N_24785);
nand UO_1700 (O_1700,N_23912,N_22692);
xor UO_1701 (O_1701,N_22942,N_21708);
xor UO_1702 (O_1702,N_24023,N_21170);
xnor UO_1703 (O_1703,N_24237,N_21763);
nor UO_1704 (O_1704,N_24422,N_24970);
nor UO_1705 (O_1705,N_23672,N_21376);
or UO_1706 (O_1706,N_21282,N_23370);
or UO_1707 (O_1707,N_23920,N_21173);
and UO_1708 (O_1708,N_20611,N_24563);
nor UO_1709 (O_1709,N_22632,N_24317);
nand UO_1710 (O_1710,N_24693,N_24270);
xnor UO_1711 (O_1711,N_20004,N_24294);
or UO_1712 (O_1712,N_20723,N_21216);
nand UO_1713 (O_1713,N_24994,N_22751);
or UO_1714 (O_1714,N_20294,N_20545);
nor UO_1715 (O_1715,N_23987,N_22607);
nor UO_1716 (O_1716,N_21841,N_22212);
xnor UO_1717 (O_1717,N_23288,N_23546);
nand UO_1718 (O_1718,N_23285,N_23438);
or UO_1719 (O_1719,N_23527,N_23935);
nor UO_1720 (O_1720,N_20554,N_21041);
and UO_1721 (O_1721,N_22118,N_20617);
nand UO_1722 (O_1722,N_24597,N_24544);
xor UO_1723 (O_1723,N_21067,N_22600);
or UO_1724 (O_1724,N_20005,N_23544);
xnor UO_1725 (O_1725,N_24591,N_24402);
nand UO_1726 (O_1726,N_20100,N_24235);
and UO_1727 (O_1727,N_21835,N_21241);
and UO_1728 (O_1728,N_23909,N_22304);
nand UO_1729 (O_1729,N_23339,N_20181);
and UO_1730 (O_1730,N_21175,N_20170);
nor UO_1731 (O_1731,N_21470,N_21661);
xnor UO_1732 (O_1732,N_21692,N_20868);
nor UO_1733 (O_1733,N_21179,N_23733);
nor UO_1734 (O_1734,N_21737,N_20692);
and UO_1735 (O_1735,N_24553,N_22456);
nand UO_1736 (O_1736,N_21386,N_21493);
and UO_1737 (O_1737,N_23779,N_24490);
nand UO_1738 (O_1738,N_24674,N_22487);
or UO_1739 (O_1739,N_21596,N_24786);
and UO_1740 (O_1740,N_21488,N_21937);
xor UO_1741 (O_1741,N_20109,N_20491);
or UO_1742 (O_1742,N_24299,N_21943);
or UO_1743 (O_1743,N_20077,N_23007);
nor UO_1744 (O_1744,N_20336,N_20241);
or UO_1745 (O_1745,N_22428,N_20726);
and UO_1746 (O_1746,N_22510,N_21431);
and UO_1747 (O_1747,N_23157,N_22201);
or UO_1748 (O_1748,N_24344,N_24615);
nand UO_1749 (O_1749,N_20832,N_21178);
and UO_1750 (O_1750,N_21326,N_24373);
nor UO_1751 (O_1751,N_22665,N_21224);
or UO_1752 (O_1752,N_21097,N_21845);
or UO_1753 (O_1753,N_24538,N_24008);
or UO_1754 (O_1754,N_21005,N_20576);
xor UO_1755 (O_1755,N_23145,N_24257);
xnor UO_1756 (O_1756,N_20907,N_20122);
xnor UO_1757 (O_1757,N_23642,N_21802);
xor UO_1758 (O_1758,N_24393,N_20388);
and UO_1759 (O_1759,N_24523,N_22559);
nand UO_1760 (O_1760,N_22399,N_20444);
and UO_1761 (O_1761,N_22878,N_20864);
nand UO_1762 (O_1762,N_24390,N_24947);
and UO_1763 (O_1763,N_22694,N_23479);
xor UO_1764 (O_1764,N_20023,N_24817);
nor UO_1765 (O_1765,N_23758,N_24128);
nor UO_1766 (O_1766,N_23990,N_23245);
or UO_1767 (O_1767,N_23665,N_24503);
nand UO_1768 (O_1768,N_22093,N_22479);
nand UO_1769 (O_1769,N_21987,N_21533);
or UO_1770 (O_1770,N_22438,N_23259);
nor UO_1771 (O_1771,N_22801,N_22866);
xor UO_1772 (O_1772,N_23850,N_22086);
nand UO_1773 (O_1773,N_21370,N_24282);
nand UO_1774 (O_1774,N_24126,N_21884);
and UO_1775 (O_1775,N_22625,N_23457);
and UO_1776 (O_1776,N_22254,N_24595);
nand UO_1777 (O_1777,N_23689,N_22101);
or UO_1778 (O_1778,N_21160,N_20656);
or UO_1779 (O_1779,N_22492,N_24941);
and UO_1780 (O_1780,N_22537,N_20383);
xnor UO_1781 (O_1781,N_23215,N_20980);
nand UO_1782 (O_1782,N_21023,N_21391);
or UO_1783 (O_1783,N_21158,N_20430);
or UO_1784 (O_1784,N_21811,N_24376);
xnor UO_1785 (O_1785,N_21121,N_21483);
nand UO_1786 (O_1786,N_21232,N_20632);
and UO_1787 (O_1787,N_22609,N_21898);
xnor UO_1788 (O_1788,N_20288,N_21314);
nand UO_1789 (O_1789,N_23455,N_22765);
and UO_1790 (O_1790,N_24579,N_23845);
nand UO_1791 (O_1791,N_20673,N_21725);
nor UO_1792 (O_1792,N_22680,N_23377);
xor UO_1793 (O_1793,N_21151,N_22952);
xnor UO_1794 (O_1794,N_21454,N_20787);
xnor UO_1795 (O_1795,N_21612,N_20934);
or UO_1796 (O_1796,N_23398,N_22912);
nor UO_1797 (O_1797,N_22035,N_20113);
or UO_1798 (O_1798,N_23102,N_24065);
and UO_1799 (O_1799,N_20631,N_20290);
nand UO_1800 (O_1800,N_22899,N_23499);
and UO_1801 (O_1801,N_20223,N_23660);
and UO_1802 (O_1802,N_24280,N_22206);
and UO_1803 (O_1803,N_21840,N_23117);
and UO_1804 (O_1804,N_20680,N_24038);
nand UO_1805 (O_1805,N_22924,N_22763);
and UO_1806 (O_1806,N_23261,N_23197);
or UO_1807 (O_1807,N_20075,N_20330);
nor UO_1808 (O_1808,N_23773,N_24583);
nor UO_1809 (O_1809,N_23702,N_24001);
nor UO_1810 (O_1810,N_23515,N_21810);
nand UO_1811 (O_1811,N_23556,N_22882);
or UO_1812 (O_1812,N_21996,N_20742);
nor UO_1813 (O_1813,N_24653,N_21078);
and UO_1814 (O_1814,N_24556,N_21090);
xnor UO_1815 (O_1815,N_24486,N_23881);
nor UO_1816 (O_1816,N_22902,N_24566);
nor UO_1817 (O_1817,N_22293,N_24309);
xnor UO_1818 (O_1818,N_22831,N_24254);
xor UO_1819 (O_1819,N_21436,N_20148);
nand UO_1820 (O_1820,N_20092,N_23015);
nor UO_1821 (O_1821,N_24116,N_21217);
and UO_1822 (O_1822,N_23866,N_20235);
and UO_1823 (O_1823,N_22732,N_23563);
or UO_1824 (O_1824,N_20363,N_23982);
and UO_1825 (O_1825,N_21653,N_20196);
nand UO_1826 (O_1826,N_23940,N_23621);
xnor UO_1827 (O_1827,N_23524,N_24745);
nand UO_1828 (O_1828,N_21746,N_20462);
nand UO_1829 (O_1829,N_21567,N_21642);
nor UO_1830 (O_1830,N_20783,N_21053);
xor UO_1831 (O_1831,N_22330,N_22306);
and UO_1832 (O_1832,N_22214,N_21754);
and UO_1833 (O_1833,N_21229,N_21322);
xor UO_1834 (O_1834,N_21983,N_21002);
nand UO_1835 (O_1835,N_21579,N_22845);
and UO_1836 (O_1836,N_20199,N_21197);
and UO_1837 (O_1837,N_24138,N_20144);
xor UO_1838 (O_1838,N_21829,N_23996);
nor UO_1839 (O_1839,N_21522,N_22802);
nor UO_1840 (O_1840,N_24072,N_22875);
nor UO_1841 (O_1841,N_24721,N_24059);
and UO_1842 (O_1842,N_22808,N_23878);
nor UO_1843 (O_1843,N_20438,N_22225);
and UO_1844 (O_1844,N_21773,N_23000);
or UO_1845 (O_1845,N_23424,N_23272);
or UO_1846 (O_1846,N_20880,N_20584);
or UO_1847 (O_1847,N_21035,N_22577);
or UO_1848 (O_1848,N_24875,N_22877);
nor UO_1849 (O_1849,N_20200,N_22516);
xor UO_1850 (O_1850,N_24296,N_22392);
nor UO_1851 (O_1851,N_22409,N_22540);
xor UO_1852 (O_1852,N_24217,N_23283);
nor UO_1853 (O_1853,N_22927,N_20865);
or UO_1854 (O_1854,N_22528,N_20312);
xnor UO_1855 (O_1855,N_20219,N_21770);
nor UO_1856 (O_1856,N_24158,N_23440);
or UO_1857 (O_1857,N_23182,N_22788);
nor UO_1858 (O_1858,N_20044,N_21293);
and UO_1859 (O_1859,N_23806,N_22362);
or UO_1860 (O_1860,N_21251,N_21527);
nor UO_1861 (O_1861,N_22164,N_24210);
xnor UO_1862 (O_1862,N_20272,N_21032);
or UO_1863 (O_1863,N_24804,N_23804);
and UO_1864 (O_1864,N_20852,N_24268);
nand UO_1865 (O_1865,N_20333,N_22722);
xor UO_1866 (O_1866,N_24925,N_20519);
nand UO_1867 (O_1867,N_22604,N_23073);
xor UO_1868 (O_1868,N_24865,N_22307);
xor UO_1869 (O_1869,N_23539,N_21535);
and UO_1870 (O_1870,N_20287,N_21583);
nand UO_1871 (O_1871,N_24548,N_20233);
xor UO_1872 (O_1872,N_22004,N_22015);
nand UO_1873 (O_1873,N_21913,N_21266);
and UO_1874 (O_1874,N_20837,N_24076);
or UO_1875 (O_1875,N_23872,N_23846);
or UO_1876 (O_1876,N_24227,N_22055);
or UO_1877 (O_1877,N_23948,N_24484);
or UO_1878 (O_1878,N_21039,N_22969);
xor UO_1879 (O_1879,N_21804,N_24136);
and UO_1880 (O_1880,N_20041,N_24026);
and UO_1881 (O_1881,N_20359,N_20668);
nor UO_1882 (O_1882,N_22605,N_24196);
nor UO_1883 (O_1883,N_23156,N_23879);
and UO_1884 (O_1884,N_24800,N_21200);
nand UO_1885 (O_1885,N_21081,N_20908);
nor UO_1886 (O_1886,N_24564,N_23442);
nand UO_1887 (O_1887,N_20546,N_24803);
or UO_1888 (O_1888,N_20970,N_22384);
xor UO_1889 (O_1889,N_21589,N_22847);
xnor UO_1890 (O_1890,N_24372,N_23803);
nor UO_1891 (O_1891,N_23329,N_24832);
and UO_1892 (O_1892,N_22713,N_24626);
and UO_1893 (O_1893,N_22382,N_24779);
xnor UO_1894 (O_1894,N_21015,N_24339);
nand UO_1895 (O_1895,N_20572,N_24368);
nor UO_1896 (O_1896,N_24688,N_20074);
and UO_1897 (O_1897,N_22065,N_21285);
or UO_1898 (O_1898,N_20833,N_22703);
and UO_1899 (O_1899,N_23405,N_22585);
xnor UO_1900 (O_1900,N_21981,N_22728);
xor UO_1901 (O_1901,N_23471,N_20110);
or UO_1902 (O_1902,N_20244,N_24840);
xor UO_1903 (O_1903,N_22426,N_24661);
and UO_1904 (O_1904,N_20840,N_21082);
nand UO_1905 (O_1905,N_21472,N_21571);
or UO_1906 (O_1906,N_20948,N_21278);
and UO_1907 (O_1907,N_22112,N_24601);
or UO_1908 (O_1908,N_21813,N_20180);
or UO_1909 (O_1909,N_21667,N_23627);
xor UO_1910 (O_1910,N_23107,N_20926);
or UO_1911 (O_1911,N_22352,N_24607);
nand UO_1912 (O_1912,N_20266,N_22938);
nor UO_1913 (O_1913,N_23163,N_23658);
or UO_1914 (O_1914,N_24148,N_22078);
and UO_1915 (O_1915,N_22947,N_24107);
nor UO_1916 (O_1916,N_21734,N_23045);
nand UO_1917 (O_1917,N_23095,N_24717);
and UO_1918 (O_1918,N_22784,N_21381);
xor UO_1919 (O_1919,N_23566,N_21300);
nand UO_1920 (O_1920,N_20248,N_21862);
and UO_1921 (O_1921,N_20737,N_24067);
or UO_1922 (O_1922,N_20263,N_22249);
xnor UO_1923 (O_1923,N_22993,N_20795);
or UO_1924 (O_1924,N_20860,N_20507);
xnor UO_1925 (O_1925,N_23619,N_22517);
nor UO_1926 (O_1926,N_23503,N_23550);
and UO_1927 (O_1927,N_24839,N_20313);
or UO_1928 (O_1928,N_21683,N_24446);
or UO_1929 (O_1929,N_22443,N_20648);
xor UO_1930 (O_1930,N_24155,N_20379);
or UO_1931 (O_1931,N_23726,N_24453);
nor UO_1932 (O_1932,N_20614,N_24469);
and UO_1933 (O_1933,N_22646,N_20769);
or UO_1934 (O_1934,N_20487,N_22138);
xor UO_1935 (O_1935,N_24991,N_23403);
nand UO_1936 (O_1936,N_22183,N_22758);
and UO_1937 (O_1937,N_23244,N_21425);
or UO_1938 (O_1938,N_23149,N_23570);
nor UO_1939 (O_1939,N_20279,N_23337);
or UO_1940 (O_1940,N_24802,N_23617);
or UO_1941 (O_1941,N_23507,N_22309);
or UO_1942 (O_1942,N_22338,N_23521);
or UO_1943 (O_1943,N_24112,N_24719);
nand UO_1944 (O_1944,N_22105,N_22322);
or UO_1945 (O_1945,N_23694,N_20026);
and UO_1946 (O_1946,N_24682,N_23884);
xor UO_1947 (O_1947,N_23856,N_23944);
nor UO_1948 (O_1948,N_21219,N_20582);
and UO_1949 (O_1949,N_22358,N_24730);
or UO_1950 (O_1950,N_22672,N_21231);
or UO_1951 (O_1951,N_22742,N_22950);
xor UO_1952 (O_1952,N_21426,N_23637);
nand UO_1953 (O_1953,N_21886,N_22807);
nor UO_1954 (O_1954,N_20820,N_22660);
and UO_1955 (O_1955,N_24133,N_21706);
nand UO_1956 (O_1956,N_20115,N_24318);
xnor UO_1957 (O_1957,N_24243,N_22483);
nand UO_1958 (O_1958,N_22641,N_23927);
nor UO_1959 (O_1959,N_22102,N_20883);
or UO_1960 (O_1960,N_21193,N_22447);
and UO_1961 (O_1961,N_23174,N_23887);
nand UO_1962 (O_1962,N_21199,N_22569);
nor UO_1963 (O_1963,N_23295,N_21656);
or UO_1964 (O_1964,N_21608,N_21517);
xnor UO_1965 (O_1965,N_24139,N_21676);
nor UO_1966 (O_1966,N_22097,N_23308);
and UO_1967 (O_1967,N_21819,N_23379);
or UO_1968 (O_1968,N_22203,N_23006);
nor UO_1969 (O_1969,N_24137,N_21477);
or UO_1970 (O_1970,N_22649,N_23919);
or UO_1971 (O_1971,N_22981,N_24326);
xnor UO_1972 (O_1972,N_23237,N_22346);
xor UO_1973 (O_1973,N_21356,N_21573);
nand UO_1974 (O_1974,N_22892,N_21307);
nor UO_1975 (O_1975,N_21348,N_24720);
nand UO_1976 (O_1976,N_23112,N_22851);
and UO_1977 (O_1977,N_20480,N_22160);
or UO_1978 (O_1978,N_20789,N_23925);
nor UO_1979 (O_1979,N_23653,N_24915);
or UO_1980 (O_1980,N_23187,N_22519);
xor UO_1981 (O_1981,N_21492,N_20392);
nand UO_1982 (O_1982,N_23492,N_21467);
nor UO_1983 (O_1983,N_20511,N_20484);
nor UO_1984 (O_1984,N_22688,N_20053);
and UO_1985 (O_1985,N_24861,N_24621);
xor UO_1986 (O_1986,N_21029,N_22077);
xor UO_1987 (O_1987,N_23001,N_23016);
nor UO_1988 (O_1988,N_21302,N_21407);
or UO_1989 (O_1989,N_20031,N_23732);
or UO_1990 (O_1990,N_24450,N_24918);
nor UO_1991 (O_1991,N_21659,N_23501);
and UO_1992 (O_1992,N_20575,N_23252);
xnor UO_1993 (O_1993,N_24425,N_24638);
xnor UO_1994 (O_1994,N_21861,N_24436);
or UO_1995 (O_1995,N_21451,N_24956);
nand UO_1996 (O_1996,N_21671,N_22359);
and UO_1997 (O_1997,N_20202,N_21396);
nor UO_1998 (O_1998,N_22470,N_24900);
nor UO_1999 (O_1999,N_21486,N_20963);
or UO_2000 (O_2000,N_23248,N_22626);
nor UO_2001 (O_2001,N_23467,N_22413);
xnor UO_2002 (O_2002,N_23624,N_21738);
nor UO_2003 (O_2003,N_24086,N_22557);
and UO_2004 (O_2004,N_21003,N_24570);
xor UO_2005 (O_2005,N_22555,N_20411);
or UO_2006 (O_2006,N_21290,N_21998);
nand UO_2007 (O_2007,N_23950,N_24616);
xor UO_2008 (O_2008,N_22800,N_24015);
and UO_2009 (O_2009,N_22490,N_20001);
nand UO_2010 (O_2010,N_21129,N_22377);
nor UO_2011 (O_2011,N_20527,N_22991);
nor UO_2012 (O_2012,N_22590,N_20822);
xnor UO_2013 (O_2013,N_20542,N_20744);
nor UO_2014 (O_2014,N_24734,N_24121);
or UO_2015 (O_2015,N_21901,N_20250);
or UO_2016 (O_2016,N_24341,N_21325);
or UO_2017 (O_2017,N_21530,N_21644);
xor UO_2018 (O_2018,N_22984,N_20972);
xnor UO_2019 (O_2019,N_20101,N_22804);
nand UO_2020 (O_2020,N_23723,N_22682);
nor UO_2021 (O_2021,N_24263,N_21794);
nand UO_2022 (O_2022,N_21186,N_22406);
xnor UO_2023 (O_2023,N_21481,N_21847);
and UO_2024 (O_2024,N_21919,N_21512);
xnor UO_2025 (O_2025,N_22398,N_20091);
or UO_2026 (O_2026,N_22031,N_23160);
and UO_2027 (O_2027,N_20715,N_22366);
nor UO_2028 (O_2028,N_20914,N_22957);
nor UO_2029 (O_2029,N_20901,N_23191);
nand UO_2030 (O_2030,N_24534,N_24395);
nand UO_2031 (O_2031,N_22884,N_20327);
or UO_2032 (O_2032,N_21849,N_24192);
or UO_2033 (O_2033,N_22173,N_21449);
nor UO_2034 (O_2034,N_20217,N_24684);
xnor UO_2035 (O_2035,N_20892,N_22999);
or UO_2036 (O_2036,N_21329,N_23030);
and UO_2037 (O_2037,N_21930,N_23371);
and UO_2038 (O_2038,N_22917,N_23880);
xor UO_2039 (O_2039,N_20303,N_24695);
nand UO_2040 (O_2040,N_20698,N_21240);
xnor UO_2041 (O_2041,N_20095,N_22174);
or UO_2042 (O_2042,N_24783,N_20778);
or UO_2043 (O_2043,N_24685,N_22676);
nor UO_2044 (O_2044,N_22365,N_24959);
nand UO_2045 (O_2045,N_20372,N_21012);
xor UO_2046 (O_2046,N_21723,N_23441);
nand UO_2047 (O_2047,N_20606,N_22144);
and UO_2048 (O_2048,N_24904,N_23196);
and UO_2049 (O_2049,N_20291,N_20264);
or UO_2050 (O_2050,N_24127,N_22874);
nand UO_2051 (O_2051,N_22032,N_22159);
nand UO_2052 (O_2052,N_23099,N_23255);
and UO_2053 (O_2053,N_24819,N_23610);
nand UO_2054 (O_2054,N_22863,N_20143);
nand UO_2055 (O_2055,N_22994,N_24283);
nand UO_2056 (O_2056,N_23835,N_21423);
xnor UO_2057 (O_2057,N_22869,N_23361);
nor UO_2058 (O_2058,N_24030,N_22735);
xnor UO_2059 (O_2059,N_23928,N_24330);
nor UO_2060 (O_2060,N_21439,N_20848);
nor UO_2061 (O_2061,N_21305,N_24041);
nor UO_2062 (O_2062,N_24102,N_21805);
nor UO_2063 (O_2063,N_22029,N_23834);
nand UO_2064 (O_2064,N_22171,N_22007);
or UO_2065 (O_2065,N_24169,N_24416);
and UO_2066 (O_2066,N_24982,N_22285);
and UO_2067 (O_2067,N_20700,N_24096);
nor UO_2068 (O_2068,N_21247,N_21955);
xor UO_2069 (O_2069,N_20776,N_24543);
xor UO_2070 (O_2070,N_20089,N_23595);
and UO_2071 (O_2071,N_24471,N_23387);
and UO_2072 (O_2072,N_24200,N_20414);
nand UO_2073 (O_2073,N_20838,N_24842);
xor UO_2074 (O_2074,N_24334,N_23167);
nor UO_2075 (O_2075,N_21776,N_24278);
nor UO_2076 (O_2076,N_21895,N_24433);
and UO_2077 (O_2077,N_21049,N_24735);
nand UO_2078 (O_2078,N_21960,N_23280);
nor UO_2079 (O_2079,N_22229,N_20335);
or UO_2080 (O_2080,N_21824,N_24463);
nand UO_2081 (O_2081,N_21172,N_23351);
nor UO_2082 (O_2082,N_21248,N_20539);
xor UO_2083 (O_2083,N_23473,N_20081);
nor UO_2084 (O_2084,N_24951,N_23386);
nand UO_2085 (O_2085,N_20664,N_21373);
and UO_2086 (O_2086,N_23728,N_22475);
and UO_2087 (O_2087,N_22064,N_21565);
and UO_2088 (O_2088,N_24700,N_24770);
nand UO_2089 (O_2089,N_22794,N_23367);
or UO_2090 (O_2090,N_22956,N_20869);
or UO_2091 (O_2091,N_23290,N_21163);
xnor UO_2092 (O_2092,N_20812,N_23596);
nor UO_2093 (O_2093,N_22150,N_23962);
and UO_2094 (O_2094,N_22246,N_23557);
or UO_2095 (O_2095,N_22584,N_22037);
and UO_2096 (O_2096,N_20137,N_24971);
nor UO_2097 (O_2097,N_21221,N_24586);
nor UO_2098 (O_2098,N_21350,N_20654);
nand UO_2099 (O_2099,N_24776,N_21785);
or UO_2100 (O_2100,N_21246,N_22074);
and UO_2101 (O_2101,N_24195,N_20971);
nand UO_2102 (O_2102,N_20096,N_21873);
xnor UO_2103 (O_2103,N_24084,N_22403);
or UO_2104 (O_2104,N_24593,N_21703);
and UO_2105 (O_2105,N_23589,N_24132);
nor UO_2106 (O_2106,N_23895,N_22770);
xnor UO_2107 (O_2107,N_22597,N_21739);
and UO_2108 (O_2108,N_20981,N_20048);
xor UO_2109 (O_2109,N_20555,N_23054);
or UO_2110 (O_2110,N_24631,N_24021);
and UO_2111 (O_2111,N_20937,N_23601);
nor UO_2112 (O_2112,N_22979,N_24256);
and UO_2113 (O_2113,N_21985,N_22685);
and UO_2114 (O_2114,N_23626,N_21111);
nand UO_2115 (O_2115,N_20642,N_23552);
and UO_2116 (O_2116,N_23260,N_20951);
xnor UO_2117 (O_2117,N_20040,N_21674);
and UO_2118 (O_2118,N_22364,N_21212);
or UO_2119 (O_2119,N_22906,N_22283);
nor UO_2120 (O_2120,N_20779,N_22978);
xnor UO_2121 (O_2121,N_23265,N_22677);
nor UO_2122 (O_2122,N_24005,N_20612);
or UO_2123 (O_2123,N_23980,N_24657);
nand UO_2124 (O_2124,N_23744,N_22328);
nor UO_2125 (O_2125,N_24847,N_23284);
or UO_2126 (O_2126,N_20657,N_20079);
and UO_2127 (O_2127,N_22606,N_24773);
or UO_2128 (O_2128,N_24060,N_21899);
and UO_2129 (O_2129,N_22714,N_22410);
or UO_2130 (O_2130,N_24643,N_23646);
and UO_2131 (O_2131,N_23381,N_21663);
and UO_2132 (O_2132,N_22071,N_22143);
and UO_2133 (O_2133,N_23138,N_24106);
nand UO_2134 (O_2134,N_22679,N_20395);
or UO_2135 (O_2135,N_24909,N_23952);
nand UO_2136 (O_2136,N_22803,N_23291);
and UO_2137 (O_2137,N_21848,N_21986);
or UO_2138 (O_2138,N_23882,N_21534);
nor UO_2139 (O_2139,N_20876,N_20666);
or UO_2140 (O_2140,N_22128,N_24518);
or UO_2141 (O_2141,N_20114,N_24887);
and UO_2142 (O_2142,N_20345,N_24663);
nor UO_2143 (O_2143,N_21544,N_22496);
nand UO_2144 (O_2144,N_20185,N_20356);
xor UO_2145 (O_2145,N_20593,N_21234);
or UO_2146 (O_2146,N_21139,N_24114);
and UO_2147 (O_2147,N_21415,N_23640);
nor UO_2148 (O_2148,N_21461,N_20194);
xnor UO_2149 (O_2149,N_20019,N_20037);
nor UO_2150 (O_2150,N_22618,N_22771);
or UO_2151 (O_2151,N_22486,N_23708);
or UO_2152 (O_2152,N_22657,N_22149);
and UO_2153 (O_2153,N_20650,N_24358);
xor UO_2154 (O_2154,N_22193,N_22192);
and UO_2155 (O_2155,N_23266,N_21141);
nand UO_2156 (O_2156,N_22720,N_23810);
and UO_2157 (O_2157,N_24610,N_22558);
xor UO_2158 (O_2158,N_22565,N_20368);
or UO_2159 (O_2159,N_22120,N_24051);
nor UO_2160 (O_2160,N_20899,N_21688);
or UO_2161 (O_2161,N_22017,N_20211);
and UO_2162 (O_2162,N_22189,N_21936);
nor UO_2163 (O_2163,N_23020,N_22476);
xnor UO_2164 (O_2164,N_22043,N_22743);
nor UO_2165 (O_2165,N_23022,N_22888);
or UO_2166 (O_2166,N_21255,N_22548);
nor UO_2167 (O_2167,N_22726,N_23594);
and UO_2168 (O_2168,N_23757,N_24147);
and UO_2169 (O_2169,N_23199,N_20067);
and UO_2170 (O_2170,N_21600,N_23072);
nand UO_2171 (O_2171,N_21816,N_21083);
xnor UO_2172 (O_2172,N_23428,N_21303);
xor UO_2173 (O_2173,N_22228,N_22711);
and UO_2174 (O_2174,N_24550,N_20072);
xor UO_2175 (O_2175,N_23218,N_24797);
nor UO_2176 (O_2176,N_22356,N_23466);
nor UO_2177 (O_2177,N_22629,N_22656);
and UO_2178 (O_2178,N_23620,N_22062);
nand UO_2179 (O_2179,N_21580,N_23558);
or UO_2180 (O_2180,N_24769,N_20158);
or UO_2181 (O_2181,N_20645,N_21690);
nand UO_2182 (O_2182,N_24901,N_20562);
and UO_2183 (O_2183,N_21142,N_23426);
nor UO_2184 (O_2184,N_23348,N_21417);
and UO_2185 (O_2185,N_24697,N_20756);
and UO_2186 (O_2186,N_22756,N_24488);
xor UO_2187 (O_2187,N_21276,N_20009);
nor UO_2188 (O_2188,N_20709,N_23860);
or UO_2189 (O_2189,N_24815,N_22345);
and UO_2190 (O_2190,N_22262,N_24578);
nor UO_2191 (O_2191,N_24188,N_22278);
nor UO_2192 (O_2192,N_21978,N_24183);
nor UO_2193 (O_2193,N_24079,N_22076);
nand UO_2194 (O_2194,N_22985,N_20996);
xnor UO_2195 (O_2195,N_22783,N_20222);
xnor UO_2196 (O_2196,N_23836,N_22630);
nand UO_2197 (O_2197,N_23631,N_23219);
nor UO_2198 (O_2198,N_24144,N_20066);
nand UO_2199 (O_2199,N_23997,N_20589);
nand UO_2200 (O_2200,N_22288,N_21934);
and UO_2201 (O_2201,N_20702,N_22780);
or UO_2202 (O_2202,N_24468,N_22933);
nor UO_2203 (O_2203,N_21338,N_24381);
nor UO_2204 (O_2204,N_23931,N_24630);
xor UO_2205 (O_2205,N_23513,N_20269);
nand UO_2206 (O_2206,N_22231,N_23537);
nor UO_2207 (O_2207,N_23391,N_22631);
and UO_2208 (O_2208,N_20413,N_22113);
nand UO_2209 (O_2209,N_23970,N_20597);
xnor UO_2210 (O_2210,N_22539,N_21013);
xor UO_2211 (O_2211,N_21790,N_22091);
and UO_2212 (O_2212,N_22140,N_20293);
nor UO_2213 (O_2213,N_23652,N_22810);
xnor UO_2214 (O_2214,N_21289,N_24812);
nand UO_2215 (O_2215,N_21815,N_24627);
nor UO_2216 (O_2216,N_20481,N_22750);
and UO_2217 (O_2217,N_20534,N_20999);
xnor UO_2218 (O_2218,N_22215,N_22773);
and UO_2219 (O_2219,N_23369,N_23110);
xnor UO_2220 (O_2220,N_21408,N_21592);
nor UO_2221 (O_2221,N_22027,N_21569);
xnor UO_2222 (O_2222,N_24068,N_21531);
or UO_2223 (O_2223,N_21797,N_24338);
xor UO_2224 (O_2224,N_24789,N_23923);
and UO_2225 (O_2225,N_23817,N_24952);
or UO_2226 (O_2226,N_23819,N_22855);
xnor UO_2227 (O_2227,N_20525,N_21389);
nand UO_2228 (O_2228,N_22987,N_20622);
and UO_2229 (O_2229,N_22799,N_21518);
nand UO_2230 (O_2230,N_23577,N_20239);
nor UO_2231 (O_2231,N_21540,N_21318);
nor UO_2232 (O_2232,N_24025,N_22526);
or UO_2233 (O_2233,N_23580,N_20358);
nand UO_2234 (O_2234,N_22474,N_24790);
xor UO_2235 (O_2235,N_21084,N_24919);
or UO_2236 (O_2236,N_20062,N_24120);
xnor UO_2237 (O_2237,N_22072,N_20818);
or UO_2238 (O_2238,N_24846,N_20172);
and UO_2239 (O_2239,N_22271,N_20955);
nand UO_2240 (O_2240,N_24224,N_22395);
and UO_2241 (O_2241,N_23999,N_22372);
nor UO_2242 (O_2242,N_21882,N_21601);
and UO_2243 (O_2243,N_24656,N_24371);
nor UO_2244 (O_2244,N_21009,N_21239);
and UO_2245 (O_2245,N_23414,N_20033);
nor UO_2246 (O_2246,N_23497,N_24742);
or UO_2247 (O_2247,N_20982,N_21932);
or UO_2248 (O_2248,N_20406,N_24983);
and UO_2249 (O_2249,N_20475,N_21244);
nand UO_2250 (O_2250,N_21447,N_24551);
and UO_2251 (O_2251,N_20561,N_24639);
nand UO_2252 (O_2252,N_21220,N_22274);
nor UO_2253 (O_2253,N_21638,N_20793);
nor UO_2254 (O_2254,N_22965,N_21560);
or UO_2255 (O_2255,N_20275,N_22497);
nand UO_2256 (O_2256,N_20765,N_22006);
and UO_2257 (O_2257,N_22302,N_22527);
or UO_2258 (O_2258,N_20946,N_20292);
or UO_2259 (O_2259,N_22085,N_24456);
nand UO_2260 (O_2260,N_21438,N_23098);
or UO_2261 (O_2261,N_23051,N_22622);
nand UO_2262 (O_2262,N_21637,N_23415);
nor UO_2263 (O_2263,N_24272,N_24004);
nand UO_2264 (O_2264,N_21394,N_23644);
and UO_2265 (O_2265,N_21622,N_24501);
xor UO_2266 (O_2266,N_22161,N_24760);
nand UO_2267 (O_2267,N_20343,N_20146);
or UO_2268 (O_2268,N_20975,N_20397);
nor UO_2269 (O_2269,N_22323,N_21712);
nor UO_2270 (O_2270,N_20938,N_23347);
xor UO_2271 (O_2271,N_21497,N_21910);
and UO_2272 (O_2272,N_20237,N_23666);
xnor UO_2273 (O_2273,N_24476,N_24673);
and UO_2274 (O_2274,N_22258,N_21031);
nand UO_2275 (O_2275,N_24083,N_24814);
nor UO_2276 (O_2276,N_24149,N_22849);
xnor UO_2277 (O_2277,N_24589,N_20322);
nand UO_2278 (O_2278,N_24168,N_21578);
xor UO_2279 (O_2279,N_23971,N_24070);
and UO_2280 (O_2280,N_22432,N_21627);
xnor UO_2281 (O_2281,N_21480,N_23233);
xnor UO_2282 (O_2282,N_21208,N_22296);
or UO_2283 (O_2283,N_24349,N_23761);
nand UO_2284 (O_2284,N_24170,N_21675);
and UO_2285 (O_2285,N_22058,N_23312);
nor UO_2286 (O_2286,N_22885,N_22718);
and UO_2287 (O_2287,N_22650,N_20944);
nor UO_2288 (O_2288,N_20260,N_21104);
nor UO_2289 (O_2289,N_23315,N_22089);
or UO_2290 (O_2290,N_23235,N_23579);
and UO_2291 (O_2291,N_23713,N_24911);
nand UO_2292 (O_2292,N_24903,N_24470);
and UO_2293 (O_2293,N_22423,N_21792);
and UO_2294 (O_2294,N_23857,N_22435);
nor UO_2295 (O_2295,N_22536,N_21400);
or UO_2296 (O_2296,N_23511,N_23193);
or UO_2297 (O_2297,N_23469,N_23183);
nand UO_2298 (O_2298,N_22131,N_24756);
or UO_2299 (O_2299,N_21371,N_21655);
nor UO_2300 (O_2300,N_24312,N_20706);
nor UO_2301 (O_2301,N_23509,N_22859);
xor UO_2302 (O_2302,N_24531,N_24054);
or UO_2303 (O_2303,N_24949,N_24340);
and UO_2304 (O_2304,N_20147,N_21024);
nand UO_2305 (O_2305,N_22562,N_20630);
or UO_2306 (O_2306,N_24398,N_24442);
nor UO_2307 (O_2307,N_21664,N_20685);
nand UO_2308 (O_2308,N_21174,N_21429);
nand UO_2309 (O_2309,N_21334,N_23021);
or UO_2310 (O_2310,N_23777,N_20003);
nor UO_2311 (O_2311,N_22261,N_21563);
or UO_2312 (O_2312,N_24055,N_21401);
xor UO_2313 (O_2313,N_22664,N_23656);
xnor UO_2314 (O_2314,N_23134,N_20766);
xnor UO_2315 (O_2315,N_20939,N_23012);
xnor UO_2316 (O_2316,N_21463,N_22637);
nor UO_2317 (O_2317,N_20734,N_24458);
xnor UO_2318 (O_2318,N_24539,N_24707);
and UO_2319 (O_2319,N_24857,N_24466);
xor UO_2320 (O_2320,N_20308,N_23668);
nand UO_2321 (O_2321,N_23204,N_21765);
nand UO_2322 (O_2322,N_20514,N_20568);
nand UO_2323 (O_2323,N_23798,N_21045);
and UO_2324 (O_2324,N_20465,N_21679);
and UO_2325 (O_2325,N_23543,N_24669);
nor UO_2326 (O_2326,N_24924,N_21858);
nor UO_2327 (O_2327,N_22543,N_21110);
xnor UO_2328 (O_2328,N_24943,N_23504);
and UO_2329 (O_2329,N_22119,N_20435);
or UO_2330 (O_2330,N_22598,N_22220);
nor UO_2331 (O_2331,N_21856,N_22326);
and UO_2332 (O_2332,N_20455,N_22184);
nor UO_2333 (O_2333,N_24710,N_23849);
xnor UO_2334 (O_2334,N_23863,N_22806);
or UO_2335 (O_2335,N_21954,N_22857);
or UO_2336 (O_2336,N_21643,N_20354);
nor UO_2337 (O_2337,N_20985,N_23876);
nor UO_2338 (O_2338,N_21760,N_24006);
and UO_2339 (O_2339,N_24367,N_22792);
nor UO_2340 (O_2340,N_20866,N_22963);
nand UO_2341 (O_2341,N_20427,N_23119);
nor UO_2342 (O_2342,N_22057,N_24588);
nor UO_2343 (O_2343,N_22843,N_22127);
nand UO_2344 (O_2344,N_22235,N_23609);
xor UO_2345 (O_2345,N_23286,N_23397);
and UO_2346 (O_2346,N_20085,N_21162);
or UO_2347 (O_2347,N_22700,N_20790);
xnor UO_2348 (O_2348,N_24508,N_22462);
or UO_2349 (O_2349,N_24650,N_21889);
xnor UO_2350 (O_2350,N_22733,N_23711);
nand UO_2351 (O_2351,N_23236,N_23363);
and UO_2352 (O_2352,N_23043,N_24118);
nand UO_2353 (O_2353,N_22759,N_24974);
xnor UO_2354 (O_2354,N_21156,N_20329);
or UO_2355 (O_2355,N_22349,N_21691);
nand UO_2356 (O_2356,N_22038,N_20851);
nor UO_2357 (O_2357,N_24016,N_24689);
and UO_2358 (O_2358,N_22782,N_22060);
xnor UO_2359 (O_2359,N_22550,N_21742);
or UO_2360 (O_2360,N_21072,N_20061);
nor UO_2361 (O_2361,N_23162,N_24907);
or UO_2362 (O_2362,N_22873,N_23989);
nand UO_2363 (O_2363,N_22095,N_22896);
xor UO_2364 (O_2364,N_20466,N_20518);
nor UO_2365 (O_2365,N_24225,N_20676);
and UO_2366 (O_2366,N_20931,N_24378);
nor UO_2367 (O_2367,N_23262,N_24872);
nand UO_2368 (O_2368,N_23611,N_23071);
nor UO_2369 (O_2369,N_24348,N_23780);
xnor UO_2370 (O_2370,N_23101,N_21762);
xnor UO_2371 (O_2371,N_22455,N_22567);
or UO_2372 (O_2372,N_24208,N_22914);
xor UO_2373 (O_2373,N_24460,N_22812);
or UO_2374 (O_2374,N_24305,N_23667);
and UO_2375 (O_2375,N_23124,N_23787);
nor UO_2376 (O_2376,N_21145,N_21669);
or UO_2377 (O_2377,N_21812,N_22457);
nand UO_2378 (O_2378,N_21485,N_24902);
xnor UO_2379 (O_2379,N_22167,N_22681);
or UO_2380 (O_2380,N_21466,N_22909);
and UO_2381 (O_2381,N_24512,N_23350);
or UO_2382 (O_2382,N_22355,N_20482);
nor UO_2383 (O_2383,N_23411,N_23495);
or UO_2384 (O_2384,N_23185,N_21621);
xnor UO_2385 (O_2385,N_20369,N_21075);
nand UO_2386 (O_2386,N_20284,N_24546);
xnor UO_2387 (O_2387,N_21133,N_20163);
or UO_2388 (O_2388,N_22968,N_24836);
nand UO_2389 (O_2389,N_22675,N_24885);
nand UO_2390 (O_2390,N_24637,N_20991);
nand UO_2391 (O_2391,N_22643,N_22226);
and UO_2392 (O_2392,N_23765,N_22333);
nand UO_2393 (O_2393,N_20119,N_22336);
or UO_2394 (O_2394,N_23638,N_22734);
nor UO_2395 (O_2395,N_24404,N_24964);
or UO_2396 (O_2396,N_20450,N_24762);
nand UO_2397 (O_2397,N_22644,N_22020);
and UO_2398 (O_2398,N_24665,N_21122);
nor UO_2399 (O_2399,N_21728,N_24191);
nand UO_2400 (O_2400,N_21808,N_24957);
nor UO_2401 (O_2401,N_23785,N_24960);
nand UO_2402 (O_2402,N_20448,N_21730);
nor UO_2403 (O_2403,N_21820,N_20968);
or UO_2404 (O_2404,N_23710,N_21903);
nor UO_2405 (O_2405,N_23888,N_22104);
xnor UO_2406 (O_2406,N_22040,N_24701);
nor UO_2407 (O_2407,N_21818,N_23657);
nand UO_2408 (O_2408,N_22595,N_23052);
nand UO_2409 (O_2409,N_23727,N_20927);
or UO_2410 (O_2410,N_21766,N_20714);
and UO_2411 (O_2411,N_23050,N_24180);
and UO_2412 (O_2412,N_20608,N_20297);
or UO_2413 (O_2413,N_23829,N_22216);
or UO_2414 (O_2414,N_24064,N_20558);
nand UO_2415 (O_2415,N_20249,N_20370);
or UO_2416 (O_2416,N_21034,N_21720);
xor UO_2417 (O_2417,N_21843,N_22481);
nand UO_2418 (O_2418,N_22115,N_21037);
xnor UO_2419 (O_2419,N_20974,N_24724);
xnor UO_2420 (O_2420,N_22561,N_20347);
xor UO_2421 (O_2421,N_22197,N_20831);
or UO_2422 (O_2422,N_22341,N_24198);
and UO_2423 (O_2423,N_20117,N_20402);
xnor UO_2424 (O_2424,N_24375,N_23221);
nor UO_2425 (O_2425,N_21980,N_24714);
or UO_2426 (O_2426,N_22256,N_22678);
and UO_2427 (O_2427,N_23268,N_22767);
nand UO_2428 (O_2428,N_24950,N_23126);
xnor UO_2429 (O_2429,N_21752,N_23669);
and UO_2430 (O_2430,N_20140,N_24567);
xor UO_2431 (O_2431,N_21062,N_24649);
nor UO_2432 (O_2432,N_22544,N_22270);
and UO_2433 (O_2433,N_21001,N_21780);
nor UO_2434 (O_2434,N_24063,N_21509);
or UO_2435 (O_2435,N_22939,N_22441);
and UO_2436 (O_2436,N_21604,N_24555);
and UO_2437 (O_2437,N_21546,N_21393);
nand UO_2438 (O_2438,N_24346,N_23851);
and UO_2439 (O_2439,N_20454,N_23349);
nor UO_2440 (O_2440,N_24434,N_24379);
or UO_2441 (O_2441,N_20841,N_24160);
and UO_2442 (O_2442,N_20587,N_22534);
or UO_2443 (O_2443,N_24360,N_20121);
nor UO_2444 (O_2444,N_20807,N_24462);
nand UO_2445 (O_2445,N_20885,N_20229);
or UO_2446 (O_2446,N_24870,N_20320);
or UO_2447 (O_2447,N_23200,N_22059);
and UO_2448 (O_2448,N_20039,N_23306);
nor UO_2449 (O_2449,N_21868,N_21052);
nor UO_2450 (O_2450,N_23973,N_23891);
or UO_2451 (O_2451,N_22122,N_23750);
and UO_2452 (O_2452,N_23797,N_23947);
nor UO_2453 (O_2453,N_21016,N_24290);
nor UO_2454 (O_2454,N_24454,N_20707);
or UO_2455 (O_2455,N_22442,N_22745);
xor UO_2456 (O_2456,N_21283,N_21074);
nor UO_2457 (O_2457,N_22499,N_24094);
xor UO_2458 (O_2458,N_21088,N_22513);
nand UO_2459 (O_2459,N_23650,N_22620);
nand UO_2460 (O_2460,N_23892,N_23009);
xnor UO_2461 (O_2461,N_23649,N_20006);
and UO_2462 (O_2462,N_20541,N_23696);
or UO_2463 (O_2463,N_21188,N_20051);
or UO_2464 (O_2464,N_23809,N_22023);
nor UO_2465 (O_2465,N_20905,N_21545);
or UO_2466 (O_2466,N_24894,N_23178);
and UO_2467 (O_2467,N_21916,N_24738);
nor UO_2468 (O_2468,N_21040,N_22719);
nor UO_2469 (O_2469,N_20570,N_22245);
or UO_2470 (O_2470,N_24600,N_23341);
nor UO_2471 (O_2471,N_20234,N_20990);
xnor UO_2472 (O_2472,N_24212,N_20762);
nand UO_2473 (O_2473,N_22407,N_22853);
nand UO_2474 (O_2474,N_22814,N_21670);
nor UO_2475 (O_2475,N_21422,N_22813);
nand UO_2476 (O_2476,N_22856,N_23169);
nor UO_2477 (O_2477,N_23496,N_20226);
or UO_2478 (O_2478,N_22570,N_24098);
or UO_2479 (O_2479,N_23588,N_24066);
nand UO_2480 (O_2480,N_20785,N_23453);
nand UO_2481 (O_2481,N_20382,N_20847);
nor UO_2482 (O_2482,N_20231,N_22408);
nor UO_2483 (O_2483,N_20828,N_24572);
nand UO_2484 (O_2484,N_21191,N_23717);
or UO_2485 (O_2485,N_23855,N_22098);
xnor UO_2486 (O_2486,N_20928,N_22809);
nor UO_2487 (O_2487,N_24095,N_24768);
nor UO_2488 (O_2488,N_24541,N_22860);
xnor UO_2489 (O_2489,N_24405,N_20097);
nand UO_2490 (O_2490,N_20416,N_23362);
or UO_2491 (O_2491,N_20190,N_21827);
and UO_2492 (O_2492,N_23584,N_23171);
and UO_2493 (O_2493,N_20278,N_24766);
nor UO_2494 (O_2494,N_21453,N_21202);
nand UO_2495 (O_2495,N_22505,N_22844);
or UO_2496 (O_2496,N_21479,N_23413);
xnor UO_2497 (O_2497,N_24448,N_22690);
and UO_2498 (O_2498,N_20651,N_24542);
and UO_2499 (O_2499,N_20268,N_24837);
nand UO_2500 (O_2500,N_21956,N_21525);
xnor UO_2501 (O_2501,N_21988,N_23850);
nor UO_2502 (O_2502,N_23765,N_20870);
nand UO_2503 (O_2503,N_24818,N_23333);
or UO_2504 (O_2504,N_20515,N_22056);
xor UO_2505 (O_2505,N_23697,N_22491);
nand UO_2506 (O_2506,N_23813,N_23927);
or UO_2507 (O_2507,N_24942,N_21336);
nor UO_2508 (O_2508,N_24089,N_23550);
or UO_2509 (O_2509,N_23988,N_21538);
and UO_2510 (O_2510,N_21870,N_24131);
xor UO_2511 (O_2511,N_21674,N_21538);
xor UO_2512 (O_2512,N_24541,N_24732);
nor UO_2513 (O_2513,N_23419,N_21185);
and UO_2514 (O_2514,N_21177,N_22444);
nand UO_2515 (O_2515,N_21379,N_24446);
or UO_2516 (O_2516,N_24350,N_21150);
nor UO_2517 (O_2517,N_20792,N_23267);
and UO_2518 (O_2518,N_24306,N_22016);
or UO_2519 (O_2519,N_20219,N_21400);
xor UO_2520 (O_2520,N_22034,N_21599);
xnor UO_2521 (O_2521,N_22426,N_21092);
xnor UO_2522 (O_2522,N_24785,N_24560);
xnor UO_2523 (O_2523,N_23128,N_23866);
or UO_2524 (O_2524,N_24924,N_22368);
or UO_2525 (O_2525,N_20962,N_21542);
xnor UO_2526 (O_2526,N_21462,N_23181);
xnor UO_2527 (O_2527,N_24309,N_21178);
xnor UO_2528 (O_2528,N_24120,N_20899);
xor UO_2529 (O_2529,N_22622,N_22548);
xor UO_2530 (O_2530,N_21900,N_24995);
nor UO_2531 (O_2531,N_21550,N_20636);
nand UO_2532 (O_2532,N_23272,N_20032);
or UO_2533 (O_2533,N_24581,N_24319);
or UO_2534 (O_2534,N_23293,N_20271);
nand UO_2535 (O_2535,N_22257,N_23402);
nor UO_2536 (O_2536,N_21890,N_21429);
or UO_2537 (O_2537,N_21723,N_24414);
nand UO_2538 (O_2538,N_20945,N_23740);
or UO_2539 (O_2539,N_22976,N_23262);
xnor UO_2540 (O_2540,N_22573,N_22728);
xnor UO_2541 (O_2541,N_23635,N_22914);
xnor UO_2542 (O_2542,N_20662,N_24974);
nand UO_2543 (O_2543,N_23027,N_21130);
nand UO_2544 (O_2544,N_22944,N_23331);
nand UO_2545 (O_2545,N_24526,N_23015);
and UO_2546 (O_2546,N_23638,N_20618);
or UO_2547 (O_2547,N_21243,N_23175);
nand UO_2548 (O_2548,N_24114,N_23413);
and UO_2549 (O_2549,N_23725,N_21471);
xor UO_2550 (O_2550,N_21485,N_20406);
nor UO_2551 (O_2551,N_21977,N_23658);
nor UO_2552 (O_2552,N_20720,N_24223);
nand UO_2553 (O_2553,N_22336,N_23180);
and UO_2554 (O_2554,N_24605,N_24250);
nor UO_2555 (O_2555,N_22806,N_22381);
and UO_2556 (O_2556,N_24278,N_23157);
nor UO_2557 (O_2557,N_21848,N_20583);
or UO_2558 (O_2558,N_22698,N_21176);
nand UO_2559 (O_2559,N_23181,N_21499);
xnor UO_2560 (O_2560,N_22887,N_20393);
xor UO_2561 (O_2561,N_24333,N_21411);
nor UO_2562 (O_2562,N_23536,N_21793);
nand UO_2563 (O_2563,N_20418,N_23237);
and UO_2564 (O_2564,N_23722,N_24882);
nand UO_2565 (O_2565,N_23681,N_21534);
or UO_2566 (O_2566,N_22173,N_24116);
or UO_2567 (O_2567,N_20541,N_22242);
xor UO_2568 (O_2568,N_20640,N_20088);
nor UO_2569 (O_2569,N_21079,N_22026);
xnor UO_2570 (O_2570,N_21116,N_24072);
or UO_2571 (O_2571,N_21124,N_21031);
nor UO_2572 (O_2572,N_22405,N_21756);
or UO_2573 (O_2573,N_23339,N_24640);
nor UO_2574 (O_2574,N_22102,N_21806);
and UO_2575 (O_2575,N_23385,N_24977);
and UO_2576 (O_2576,N_23183,N_21472);
or UO_2577 (O_2577,N_21643,N_24928);
and UO_2578 (O_2578,N_23928,N_24017);
xor UO_2579 (O_2579,N_21795,N_22766);
and UO_2580 (O_2580,N_22222,N_22792);
or UO_2581 (O_2581,N_22171,N_20459);
nor UO_2582 (O_2582,N_20030,N_20908);
or UO_2583 (O_2583,N_23726,N_23716);
or UO_2584 (O_2584,N_23722,N_22012);
and UO_2585 (O_2585,N_24600,N_23637);
nor UO_2586 (O_2586,N_20124,N_24009);
nand UO_2587 (O_2587,N_21511,N_23728);
nor UO_2588 (O_2588,N_21051,N_21384);
nor UO_2589 (O_2589,N_24276,N_20215);
xnor UO_2590 (O_2590,N_21614,N_23423);
and UO_2591 (O_2591,N_21587,N_22930);
nor UO_2592 (O_2592,N_22106,N_21606);
and UO_2593 (O_2593,N_21240,N_21065);
or UO_2594 (O_2594,N_21437,N_20720);
nor UO_2595 (O_2595,N_21905,N_21088);
xnor UO_2596 (O_2596,N_23340,N_20683);
and UO_2597 (O_2597,N_22658,N_24370);
or UO_2598 (O_2598,N_23065,N_20630);
or UO_2599 (O_2599,N_21167,N_22332);
and UO_2600 (O_2600,N_22829,N_24012);
xnor UO_2601 (O_2601,N_23834,N_20842);
nand UO_2602 (O_2602,N_20735,N_20095);
or UO_2603 (O_2603,N_23947,N_24302);
or UO_2604 (O_2604,N_20508,N_24021);
xor UO_2605 (O_2605,N_22269,N_24368);
xnor UO_2606 (O_2606,N_20909,N_22103);
and UO_2607 (O_2607,N_24416,N_20486);
or UO_2608 (O_2608,N_21323,N_23587);
nand UO_2609 (O_2609,N_20055,N_21453);
or UO_2610 (O_2610,N_22330,N_20101);
nor UO_2611 (O_2611,N_23114,N_21153);
nand UO_2612 (O_2612,N_21982,N_23853);
nand UO_2613 (O_2613,N_22602,N_23646);
nor UO_2614 (O_2614,N_23666,N_22302);
or UO_2615 (O_2615,N_24803,N_24199);
and UO_2616 (O_2616,N_21495,N_23849);
and UO_2617 (O_2617,N_21095,N_21778);
xor UO_2618 (O_2618,N_23722,N_20641);
nand UO_2619 (O_2619,N_23170,N_20898);
and UO_2620 (O_2620,N_24853,N_20911);
or UO_2621 (O_2621,N_22274,N_24123);
xor UO_2622 (O_2622,N_24705,N_21825);
and UO_2623 (O_2623,N_20694,N_24289);
and UO_2624 (O_2624,N_22469,N_23220);
nor UO_2625 (O_2625,N_20166,N_20604);
nor UO_2626 (O_2626,N_20712,N_23299);
nand UO_2627 (O_2627,N_24350,N_22511);
or UO_2628 (O_2628,N_21666,N_24410);
or UO_2629 (O_2629,N_23842,N_20538);
xnor UO_2630 (O_2630,N_21746,N_22435);
nand UO_2631 (O_2631,N_24453,N_20700);
nor UO_2632 (O_2632,N_22763,N_24456);
nand UO_2633 (O_2633,N_20801,N_24268);
and UO_2634 (O_2634,N_24590,N_22204);
and UO_2635 (O_2635,N_21873,N_24542);
nor UO_2636 (O_2636,N_22583,N_21196);
nand UO_2637 (O_2637,N_22737,N_22368);
or UO_2638 (O_2638,N_23766,N_22307);
and UO_2639 (O_2639,N_22673,N_21278);
xnor UO_2640 (O_2640,N_24577,N_20883);
xnor UO_2641 (O_2641,N_21516,N_21751);
nor UO_2642 (O_2642,N_21299,N_21832);
and UO_2643 (O_2643,N_23245,N_21049);
nand UO_2644 (O_2644,N_20806,N_22575);
nor UO_2645 (O_2645,N_24578,N_24821);
or UO_2646 (O_2646,N_24839,N_20267);
or UO_2647 (O_2647,N_24067,N_20136);
and UO_2648 (O_2648,N_23366,N_21189);
nand UO_2649 (O_2649,N_22588,N_23249);
xor UO_2650 (O_2650,N_21155,N_24597);
or UO_2651 (O_2651,N_20547,N_22708);
nand UO_2652 (O_2652,N_20848,N_24889);
nand UO_2653 (O_2653,N_23292,N_22975);
and UO_2654 (O_2654,N_21196,N_20860);
and UO_2655 (O_2655,N_24065,N_23381);
nor UO_2656 (O_2656,N_22646,N_24631);
xnor UO_2657 (O_2657,N_24715,N_20624);
nor UO_2658 (O_2658,N_24467,N_23961);
nand UO_2659 (O_2659,N_24156,N_23686);
nor UO_2660 (O_2660,N_21616,N_21575);
or UO_2661 (O_2661,N_24442,N_22629);
nand UO_2662 (O_2662,N_20931,N_22760);
or UO_2663 (O_2663,N_20219,N_24836);
xor UO_2664 (O_2664,N_22046,N_22037);
or UO_2665 (O_2665,N_24724,N_21608);
or UO_2666 (O_2666,N_21034,N_21025);
or UO_2667 (O_2667,N_21592,N_23576);
and UO_2668 (O_2668,N_20119,N_23870);
xnor UO_2669 (O_2669,N_20247,N_22887);
nand UO_2670 (O_2670,N_22790,N_23304);
xor UO_2671 (O_2671,N_22282,N_24428);
and UO_2672 (O_2672,N_22736,N_24920);
or UO_2673 (O_2673,N_20008,N_20474);
xnor UO_2674 (O_2674,N_23959,N_21153);
xnor UO_2675 (O_2675,N_22204,N_20256);
or UO_2676 (O_2676,N_22897,N_23382);
or UO_2677 (O_2677,N_23266,N_22536);
nor UO_2678 (O_2678,N_24911,N_22591);
or UO_2679 (O_2679,N_23131,N_24012);
and UO_2680 (O_2680,N_24924,N_22497);
nand UO_2681 (O_2681,N_24167,N_22659);
xor UO_2682 (O_2682,N_21746,N_21909);
xnor UO_2683 (O_2683,N_24649,N_22262);
nand UO_2684 (O_2684,N_20437,N_23150);
nand UO_2685 (O_2685,N_20762,N_24995);
and UO_2686 (O_2686,N_23114,N_24857);
and UO_2687 (O_2687,N_21192,N_23022);
nand UO_2688 (O_2688,N_20293,N_23774);
and UO_2689 (O_2689,N_23682,N_20998);
nor UO_2690 (O_2690,N_21359,N_22320);
and UO_2691 (O_2691,N_20412,N_23861);
or UO_2692 (O_2692,N_22086,N_21919);
nand UO_2693 (O_2693,N_23749,N_24333);
and UO_2694 (O_2694,N_22137,N_21869);
xor UO_2695 (O_2695,N_24137,N_20428);
nand UO_2696 (O_2696,N_20513,N_21560);
xor UO_2697 (O_2697,N_24405,N_21924);
or UO_2698 (O_2698,N_21851,N_22554);
and UO_2699 (O_2699,N_24179,N_23922);
nor UO_2700 (O_2700,N_21371,N_20447);
or UO_2701 (O_2701,N_20151,N_20441);
xnor UO_2702 (O_2702,N_20898,N_21237);
xor UO_2703 (O_2703,N_21244,N_20445);
xor UO_2704 (O_2704,N_22367,N_24845);
nand UO_2705 (O_2705,N_22743,N_23129);
or UO_2706 (O_2706,N_23789,N_24428);
nand UO_2707 (O_2707,N_23350,N_21143);
nand UO_2708 (O_2708,N_20479,N_21958);
nand UO_2709 (O_2709,N_21789,N_23538);
and UO_2710 (O_2710,N_20930,N_21589);
xnor UO_2711 (O_2711,N_23742,N_20948);
nor UO_2712 (O_2712,N_20451,N_20416);
nand UO_2713 (O_2713,N_23700,N_24566);
and UO_2714 (O_2714,N_23283,N_22101);
nor UO_2715 (O_2715,N_20908,N_21936);
nor UO_2716 (O_2716,N_20480,N_24951);
xnor UO_2717 (O_2717,N_21948,N_21286);
or UO_2718 (O_2718,N_24387,N_24969);
and UO_2719 (O_2719,N_20633,N_21810);
xor UO_2720 (O_2720,N_24488,N_22294);
nand UO_2721 (O_2721,N_23687,N_22463);
or UO_2722 (O_2722,N_23146,N_20873);
nor UO_2723 (O_2723,N_21464,N_24658);
nand UO_2724 (O_2724,N_22628,N_23985);
and UO_2725 (O_2725,N_22934,N_23393);
and UO_2726 (O_2726,N_23963,N_22090);
nor UO_2727 (O_2727,N_23234,N_21536);
nand UO_2728 (O_2728,N_22353,N_20026);
and UO_2729 (O_2729,N_22424,N_23993);
or UO_2730 (O_2730,N_22771,N_24740);
nand UO_2731 (O_2731,N_20695,N_20292);
xor UO_2732 (O_2732,N_22847,N_23381);
or UO_2733 (O_2733,N_20660,N_21135);
and UO_2734 (O_2734,N_20317,N_24920);
or UO_2735 (O_2735,N_22506,N_20571);
or UO_2736 (O_2736,N_21092,N_24229);
nor UO_2737 (O_2737,N_22927,N_24724);
nand UO_2738 (O_2738,N_21727,N_24672);
and UO_2739 (O_2739,N_23635,N_21964);
nor UO_2740 (O_2740,N_20370,N_22798);
or UO_2741 (O_2741,N_24079,N_20903);
nor UO_2742 (O_2742,N_23083,N_23105);
or UO_2743 (O_2743,N_23267,N_21258);
or UO_2744 (O_2744,N_20231,N_23836);
or UO_2745 (O_2745,N_23191,N_24930);
nand UO_2746 (O_2746,N_24611,N_24164);
nand UO_2747 (O_2747,N_22896,N_20994);
or UO_2748 (O_2748,N_23103,N_22592);
xor UO_2749 (O_2749,N_24488,N_20406);
nor UO_2750 (O_2750,N_24207,N_24834);
xnor UO_2751 (O_2751,N_23948,N_22418);
and UO_2752 (O_2752,N_21275,N_24121);
xor UO_2753 (O_2753,N_21371,N_23424);
nor UO_2754 (O_2754,N_21140,N_21662);
or UO_2755 (O_2755,N_20925,N_21784);
or UO_2756 (O_2756,N_22931,N_24232);
nor UO_2757 (O_2757,N_20639,N_22127);
nand UO_2758 (O_2758,N_20874,N_22035);
nor UO_2759 (O_2759,N_20469,N_22522);
and UO_2760 (O_2760,N_22052,N_22988);
xnor UO_2761 (O_2761,N_21441,N_20579);
xor UO_2762 (O_2762,N_21103,N_23752);
xor UO_2763 (O_2763,N_21387,N_21099);
nor UO_2764 (O_2764,N_23679,N_21616);
xor UO_2765 (O_2765,N_23372,N_23528);
or UO_2766 (O_2766,N_20455,N_24655);
nor UO_2767 (O_2767,N_24525,N_21108);
xor UO_2768 (O_2768,N_23715,N_21305);
or UO_2769 (O_2769,N_21106,N_20436);
nand UO_2770 (O_2770,N_20147,N_20897);
xnor UO_2771 (O_2771,N_24736,N_20684);
nor UO_2772 (O_2772,N_22626,N_24396);
nand UO_2773 (O_2773,N_22004,N_24684);
xor UO_2774 (O_2774,N_24850,N_20119);
nor UO_2775 (O_2775,N_23488,N_24206);
xor UO_2776 (O_2776,N_24708,N_20466);
or UO_2777 (O_2777,N_23901,N_24595);
nand UO_2778 (O_2778,N_21726,N_22792);
xor UO_2779 (O_2779,N_22634,N_20170);
nand UO_2780 (O_2780,N_24922,N_22819);
nand UO_2781 (O_2781,N_21141,N_22706);
or UO_2782 (O_2782,N_22118,N_22690);
nor UO_2783 (O_2783,N_23585,N_23268);
xor UO_2784 (O_2784,N_24234,N_21727);
nor UO_2785 (O_2785,N_21211,N_24366);
nor UO_2786 (O_2786,N_21160,N_24427);
nand UO_2787 (O_2787,N_20292,N_21174);
or UO_2788 (O_2788,N_24961,N_23714);
and UO_2789 (O_2789,N_22781,N_20520);
or UO_2790 (O_2790,N_20682,N_23680);
xnor UO_2791 (O_2791,N_23775,N_22718);
and UO_2792 (O_2792,N_20995,N_20702);
or UO_2793 (O_2793,N_20982,N_22046);
or UO_2794 (O_2794,N_20093,N_22639);
and UO_2795 (O_2795,N_20850,N_22988);
nand UO_2796 (O_2796,N_23041,N_20254);
or UO_2797 (O_2797,N_23716,N_24652);
xor UO_2798 (O_2798,N_24733,N_21193);
nand UO_2799 (O_2799,N_20204,N_20792);
nor UO_2800 (O_2800,N_20246,N_24063);
nor UO_2801 (O_2801,N_21250,N_22809);
or UO_2802 (O_2802,N_24787,N_24989);
or UO_2803 (O_2803,N_21039,N_22860);
nor UO_2804 (O_2804,N_22193,N_20428);
nand UO_2805 (O_2805,N_23707,N_23741);
or UO_2806 (O_2806,N_23849,N_24234);
nand UO_2807 (O_2807,N_24644,N_20463);
xnor UO_2808 (O_2808,N_21146,N_22818);
nor UO_2809 (O_2809,N_23135,N_20421);
or UO_2810 (O_2810,N_23712,N_24974);
and UO_2811 (O_2811,N_24802,N_22042);
and UO_2812 (O_2812,N_23398,N_24772);
and UO_2813 (O_2813,N_20670,N_22372);
and UO_2814 (O_2814,N_21029,N_22555);
and UO_2815 (O_2815,N_20096,N_21403);
xnor UO_2816 (O_2816,N_21382,N_20108);
or UO_2817 (O_2817,N_21621,N_24951);
xnor UO_2818 (O_2818,N_21857,N_20927);
nand UO_2819 (O_2819,N_22096,N_20878);
xor UO_2820 (O_2820,N_22410,N_21593);
nand UO_2821 (O_2821,N_20956,N_21830);
nand UO_2822 (O_2822,N_21268,N_23940);
xor UO_2823 (O_2823,N_24476,N_20069);
or UO_2824 (O_2824,N_22841,N_22274);
or UO_2825 (O_2825,N_21387,N_21018);
nor UO_2826 (O_2826,N_22026,N_24984);
xor UO_2827 (O_2827,N_22138,N_21132);
xor UO_2828 (O_2828,N_21754,N_22425);
and UO_2829 (O_2829,N_24924,N_22786);
or UO_2830 (O_2830,N_24243,N_24728);
nor UO_2831 (O_2831,N_20096,N_20775);
nor UO_2832 (O_2832,N_23403,N_21605);
and UO_2833 (O_2833,N_21824,N_22492);
or UO_2834 (O_2834,N_24709,N_21021);
nand UO_2835 (O_2835,N_24990,N_20689);
xnor UO_2836 (O_2836,N_21367,N_21365);
nand UO_2837 (O_2837,N_21280,N_24846);
or UO_2838 (O_2838,N_22294,N_20519);
xnor UO_2839 (O_2839,N_23459,N_24168);
or UO_2840 (O_2840,N_20170,N_22799);
and UO_2841 (O_2841,N_23962,N_23974);
nand UO_2842 (O_2842,N_21231,N_21227);
nor UO_2843 (O_2843,N_20582,N_20442);
or UO_2844 (O_2844,N_22703,N_24540);
or UO_2845 (O_2845,N_20788,N_20067);
nand UO_2846 (O_2846,N_24097,N_24483);
xnor UO_2847 (O_2847,N_23103,N_24946);
or UO_2848 (O_2848,N_21254,N_23324);
or UO_2849 (O_2849,N_22115,N_23356);
nor UO_2850 (O_2850,N_21885,N_24943);
or UO_2851 (O_2851,N_24391,N_22576);
and UO_2852 (O_2852,N_22000,N_21730);
xor UO_2853 (O_2853,N_21693,N_20227);
xor UO_2854 (O_2854,N_22745,N_21750);
nor UO_2855 (O_2855,N_21180,N_22086);
nor UO_2856 (O_2856,N_22417,N_24481);
nor UO_2857 (O_2857,N_20563,N_22415);
nor UO_2858 (O_2858,N_23341,N_23797);
or UO_2859 (O_2859,N_23332,N_24472);
nor UO_2860 (O_2860,N_20426,N_23392);
or UO_2861 (O_2861,N_20129,N_21064);
and UO_2862 (O_2862,N_20745,N_21864);
and UO_2863 (O_2863,N_20599,N_23630);
and UO_2864 (O_2864,N_20316,N_24185);
nor UO_2865 (O_2865,N_21566,N_24358);
or UO_2866 (O_2866,N_23810,N_21254);
nand UO_2867 (O_2867,N_24219,N_22176);
or UO_2868 (O_2868,N_22109,N_20809);
nand UO_2869 (O_2869,N_20782,N_21624);
xor UO_2870 (O_2870,N_24486,N_22774);
or UO_2871 (O_2871,N_21773,N_23844);
nand UO_2872 (O_2872,N_24802,N_23484);
or UO_2873 (O_2873,N_22932,N_20189);
xnor UO_2874 (O_2874,N_21492,N_20964);
or UO_2875 (O_2875,N_21447,N_20706);
xor UO_2876 (O_2876,N_21867,N_21355);
xnor UO_2877 (O_2877,N_20877,N_24426);
nand UO_2878 (O_2878,N_21689,N_22925);
and UO_2879 (O_2879,N_20074,N_24864);
or UO_2880 (O_2880,N_20355,N_23003);
or UO_2881 (O_2881,N_24489,N_24258);
or UO_2882 (O_2882,N_21641,N_22817);
nand UO_2883 (O_2883,N_23839,N_24142);
nor UO_2884 (O_2884,N_21514,N_21630);
nor UO_2885 (O_2885,N_20616,N_23518);
nor UO_2886 (O_2886,N_21462,N_22249);
xor UO_2887 (O_2887,N_21559,N_24950);
and UO_2888 (O_2888,N_20157,N_20680);
nor UO_2889 (O_2889,N_23003,N_20225);
xnor UO_2890 (O_2890,N_24650,N_23303);
nor UO_2891 (O_2891,N_24064,N_24470);
nand UO_2892 (O_2892,N_20752,N_21823);
nand UO_2893 (O_2893,N_23737,N_20514);
nand UO_2894 (O_2894,N_20405,N_22097);
and UO_2895 (O_2895,N_23769,N_24849);
nor UO_2896 (O_2896,N_20798,N_20294);
and UO_2897 (O_2897,N_20090,N_20756);
or UO_2898 (O_2898,N_20854,N_20102);
or UO_2899 (O_2899,N_22843,N_20646);
nand UO_2900 (O_2900,N_22614,N_23041);
and UO_2901 (O_2901,N_20736,N_21414);
nand UO_2902 (O_2902,N_24515,N_20713);
xor UO_2903 (O_2903,N_20263,N_21801);
and UO_2904 (O_2904,N_21460,N_22876);
nand UO_2905 (O_2905,N_24928,N_20506);
xor UO_2906 (O_2906,N_23637,N_22550);
xor UO_2907 (O_2907,N_22069,N_23211);
xnor UO_2908 (O_2908,N_23845,N_22824);
xor UO_2909 (O_2909,N_21442,N_24815);
xor UO_2910 (O_2910,N_23567,N_21703);
and UO_2911 (O_2911,N_20921,N_22710);
nand UO_2912 (O_2912,N_24757,N_23281);
and UO_2913 (O_2913,N_23514,N_24463);
and UO_2914 (O_2914,N_23239,N_20096);
or UO_2915 (O_2915,N_21988,N_20464);
or UO_2916 (O_2916,N_21209,N_21035);
xor UO_2917 (O_2917,N_22297,N_24888);
and UO_2918 (O_2918,N_22437,N_22261);
and UO_2919 (O_2919,N_20496,N_22168);
and UO_2920 (O_2920,N_21747,N_23279);
or UO_2921 (O_2921,N_20545,N_23085);
nor UO_2922 (O_2922,N_23148,N_24164);
nor UO_2923 (O_2923,N_20529,N_22161);
nand UO_2924 (O_2924,N_21754,N_20556);
and UO_2925 (O_2925,N_23011,N_24093);
and UO_2926 (O_2926,N_22607,N_23771);
or UO_2927 (O_2927,N_22452,N_20526);
xor UO_2928 (O_2928,N_21654,N_21044);
nand UO_2929 (O_2929,N_22013,N_22559);
nor UO_2930 (O_2930,N_22176,N_21506);
and UO_2931 (O_2931,N_20864,N_22565);
xnor UO_2932 (O_2932,N_24841,N_23585);
or UO_2933 (O_2933,N_23850,N_21463);
or UO_2934 (O_2934,N_23640,N_23727);
or UO_2935 (O_2935,N_22885,N_22059);
xor UO_2936 (O_2936,N_24000,N_20767);
or UO_2937 (O_2937,N_20321,N_20190);
nor UO_2938 (O_2938,N_24678,N_24544);
and UO_2939 (O_2939,N_21819,N_20280);
and UO_2940 (O_2940,N_20980,N_22707);
and UO_2941 (O_2941,N_20889,N_21931);
or UO_2942 (O_2942,N_22282,N_23088);
xnor UO_2943 (O_2943,N_22560,N_23764);
or UO_2944 (O_2944,N_20067,N_22709);
nor UO_2945 (O_2945,N_22379,N_21276);
and UO_2946 (O_2946,N_22848,N_20402);
or UO_2947 (O_2947,N_22707,N_23345);
nand UO_2948 (O_2948,N_21899,N_21325);
nor UO_2949 (O_2949,N_24816,N_20686);
and UO_2950 (O_2950,N_24296,N_22176);
nor UO_2951 (O_2951,N_22237,N_22813);
xnor UO_2952 (O_2952,N_22312,N_22460);
and UO_2953 (O_2953,N_24141,N_22800);
or UO_2954 (O_2954,N_22939,N_24681);
or UO_2955 (O_2955,N_21256,N_21398);
nand UO_2956 (O_2956,N_23710,N_20975);
or UO_2957 (O_2957,N_24231,N_21742);
nor UO_2958 (O_2958,N_22730,N_22679);
nor UO_2959 (O_2959,N_24207,N_24179);
and UO_2960 (O_2960,N_23805,N_20620);
and UO_2961 (O_2961,N_24028,N_23979);
nor UO_2962 (O_2962,N_20828,N_20776);
xnor UO_2963 (O_2963,N_24960,N_20114);
and UO_2964 (O_2964,N_21965,N_24070);
or UO_2965 (O_2965,N_20379,N_23492);
or UO_2966 (O_2966,N_21739,N_21911);
xor UO_2967 (O_2967,N_24131,N_20970);
and UO_2968 (O_2968,N_22390,N_24590);
nor UO_2969 (O_2969,N_20297,N_23242);
and UO_2970 (O_2970,N_24324,N_20361);
and UO_2971 (O_2971,N_24366,N_22674);
nor UO_2972 (O_2972,N_21052,N_23211);
nand UO_2973 (O_2973,N_22065,N_24406);
xnor UO_2974 (O_2974,N_21584,N_21961);
nand UO_2975 (O_2975,N_23891,N_20371);
nand UO_2976 (O_2976,N_20387,N_20855);
nand UO_2977 (O_2977,N_21440,N_24938);
xor UO_2978 (O_2978,N_22984,N_21930);
nor UO_2979 (O_2979,N_20716,N_24668);
xnor UO_2980 (O_2980,N_24658,N_24071);
or UO_2981 (O_2981,N_21863,N_21286);
nand UO_2982 (O_2982,N_21128,N_22878);
nor UO_2983 (O_2983,N_24293,N_23251);
nand UO_2984 (O_2984,N_24428,N_21499);
and UO_2985 (O_2985,N_24117,N_20495);
and UO_2986 (O_2986,N_22690,N_21140);
nand UO_2987 (O_2987,N_20335,N_24876);
xor UO_2988 (O_2988,N_21210,N_21899);
and UO_2989 (O_2989,N_23775,N_23386);
xnor UO_2990 (O_2990,N_21992,N_21325);
nand UO_2991 (O_2991,N_21680,N_24785);
nand UO_2992 (O_2992,N_22841,N_23334);
and UO_2993 (O_2993,N_22094,N_21961);
nor UO_2994 (O_2994,N_21597,N_24199);
xnor UO_2995 (O_2995,N_22217,N_21357);
nand UO_2996 (O_2996,N_23740,N_22327);
nor UO_2997 (O_2997,N_24943,N_20455);
nand UO_2998 (O_2998,N_22923,N_23311);
xor UO_2999 (O_2999,N_20812,N_21651);
endmodule