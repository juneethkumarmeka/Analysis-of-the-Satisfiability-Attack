module basic_500_3000_500_50_levels_1xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_205,In_387);
or U1 (N_1,In_150,In_72);
nor U2 (N_2,In_273,In_130);
or U3 (N_3,In_44,In_473);
nand U4 (N_4,In_93,In_415);
nor U5 (N_5,In_78,In_177);
and U6 (N_6,In_460,In_185);
or U7 (N_7,In_295,In_179);
or U8 (N_8,In_359,In_99);
and U9 (N_9,In_430,In_138);
or U10 (N_10,In_164,In_155);
or U11 (N_11,In_300,In_367);
and U12 (N_12,In_21,In_431);
nand U13 (N_13,In_362,In_38);
nor U14 (N_14,In_453,In_70);
nor U15 (N_15,In_19,In_71);
and U16 (N_16,In_158,In_234);
nor U17 (N_17,In_161,In_497);
nand U18 (N_18,In_486,In_293);
nor U19 (N_19,In_88,In_271);
and U20 (N_20,In_7,In_207);
and U21 (N_21,In_268,In_356);
nand U22 (N_22,In_477,In_220);
nand U23 (N_23,In_303,In_421);
and U24 (N_24,In_14,In_364);
nand U25 (N_25,In_382,In_353);
nor U26 (N_26,In_376,In_11);
nand U27 (N_27,In_348,In_90);
and U28 (N_28,In_17,In_258);
and U29 (N_29,In_326,In_474);
or U30 (N_30,In_288,In_169);
nor U31 (N_31,In_314,In_468);
nor U32 (N_32,In_231,In_29);
or U33 (N_33,In_193,In_143);
nand U34 (N_34,In_168,In_266);
nor U35 (N_35,In_407,In_107);
nor U36 (N_36,In_2,In_311);
nand U37 (N_37,In_406,In_383);
or U38 (N_38,In_124,In_328);
and U39 (N_39,In_20,In_187);
nor U40 (N_40,In_375,In_381);
nor U41 (N_41,In_27,In_190);
nand U42 (N_42,In_191,In_126);
and U43 (N_43,In_246,In_308);
xor U44 (N_44,In_22,In_218);
nor U45 (N_45,In_250,In_197);
or U46 (N_46,In_346,In_410);
nand U47 (N_47,In_60,In_103);
nand U48 (N_48,In_104,In_449);
or U49 (N_49,In_46,In_74);
or U50 (N_50,In_132,In_263);
nor U51 (N_51,In_446,In_35);
nor U52 (N_52,In_42,In_23);
nor U53 (N_53,In_251,In_96);
and U54 (N_54,In_31,In_345);
and U55 (N_55,In_144,In_120);
xor U56 (N_56,In_463,In_276);
nor U57 (N_57,In_129,In_133);
and U58 (N_58,In_136,In_214);
or U59 (N_59,In_76,In_84);
or U60 (N_60,In_489,In_272);
nor U61 (N_61,In_58,In_432);
nand U62 (N_62,In_163,N_26);
nand U63 (N_63,In_373,In_285);
and U64 (N_64,In_264,In_330);
or U65 (N_65,In_494,In_149);
nor U66 (N_66,In_294,In_389);
and U67 (N_67,In_223,In_395);
and U68 (N_68,In_82,In_472);
nand U69 (N_69,In_301,In_122);
nor U70 (N_70,In_9,In_53);
or U71 (N_71,In_255,In_426);
or U72 (N_72,In_230,In_341);
nor U73 (N_73,In_202,In_384);
and U74 (N_74,In_480,N_49);
or U75 (N_75,N_10,In_420);
nor U76 (N_76,In_261,In_335);
nand U77 (N_77,In_405,In_3);
and U78 (N_78,In_305,In_418);
or U79 (N_79,In_113,In_352);
nand U80 (N_80,In_391,In_427);
nand U81 (N_81,In_342,In_317);
or U82 (N_82,In_236,In_227);
and U83 (N_83,In_248,N_42);
and U84 (N_84,In_444,In_438);
and U85 (N_85,In_313,In_215);
or U86 (N_86,In_487,In_488);
or U87 (N_87,In_119,In_262);
and U88 (N_88,In_94,N_9);
nor U89 (N_89,In_456,In_323);
and U90 (N_90,In_403,In_192);
and U91 (N_91,In_67,In_12);
nand U92 (N_92,In_279,In_278);
or U93 (N_93,In_404,In_157);
and U94 (N_94,In_361,In_217);
or U95 (N_95,In_57,In_265);
and U96 (N_96,In_457,N_16);
and U97 (N_97,In_422,N_2);
or U98 (N_98,N_23,In_189);
and U99 (N_99,N_20,In_254);
or U100 (N_100,In_43,In_399);
and U101 (N_101,In_483,In_36);
and U102 (N_102,In_225,In_165);
and U103 (N_103,N_57,In_203);
or U104 (N_104,In_269,In_388);
nand U105 (N_105,In_50,In_114);
and U106 (N_106,In_45,In_471);
nand U107 (N_107,N_31,In_172);
nand U108 (N_108,N_17,In_370);
nor U109 (N_109,In_439,In_13);
nand U110 (N_110,N_56,In_413);
or U111 (N_111,In_222,N_53);
and U112 (N_112,In_75,In_372);
nand U113 (N_113,In_343,In_182);
or U114 (N_114,In_175,In_379);
nand U115 (N_115,In_32,In_33);
and U116 (N_116,In_26,In_66);
nand U117 (N_117,In_434,In_321);
and U118 (N_118,In_18,In_15);
xnor U119 (N_119,In_425,In_493);
or U120 (N_120,In_451,In_226);
or U121 (N_121,In_318,In_257);
or U122 (N_122,In_319,In_54);
nor U123 (N_123,N_30,In_62);
or U124 (N_124,N_73,In_307);
nor U125 (N_125,In_243,In_210);
nor U126 (N_126,N_45,N_100);
nand U127 (N_127,In_491,In_117);
nor U128 (N_128,In_476,N_69);
nor U129 (N_129,In_495,In_141);
nor U130 (N_130,N_15,N_105);
nand U131 (N_131,In_454,N_114);
or U132 (N_132,In_30,In_28);
nand U133 (N_133,In_37,In_47);
or U134 (N_134,In_101,In_337);
or U135 (N_135,In_91,N_8);
and U136 (N_136,N_85,In_366);
and U137 (N_137,In_180,In_386);
or U138 (N_138,In_59,In_284);
nor U139 (N_139,In_152,In_398);
and U140 (N_140,In_332,In_436);
or U141 (N_141,N_93,In_83);
and U142 (N_142,N_34,In_482);
nor U143 (N_143,In_292,In_241);
or U144 (N_144,N_27,In_89);
nor U145 (N_145,In_208,In_419);
nand U146 (N_146,In_10,In_160);
or U147 (N_147,In_52,In_4);
and U148 (N_148,N_119,In_423);
nor U149 (N_149,In_167,N_11);
and U150 (N_150,N_51,N_102);
and U151 (N_151,In_100,N_71);
nor U152 (N_152,In_412,In_360);
and U153 (N_153,In_134,In_338);
nand U154 (N_154,In_238,In_183);
and U155 (N_155,In_242,In_390);
and U156 (N_156,In_414,In_291);
nor U157 (N_157,In_441,In_51);
or U158 (N_158,N_43,In_209);
nand U159 (N_159,In_170,In_385);
nand U160 (N_160,In_498,In_302);
nand U161 (N_161,In_123,In_184);
and U162 (N_162,N_13,In_137);
or U163 (N_163,In_277,N_7);
or U164 (N_164,In_485,In_440);
nand U165 (N_165,In_198,N_36);
or U166 (N_166,N_94,In_206);
and U167 (N_167,In_5,N_90);
nand U168 (N_168,N_83,N_54);
and U169 (N_169,In_105,In_232);
nand U170 (N_170,In_173,In_461);
or U171 (N_171,In_287,In_296);
and U172 (N_172,N_115,In_111);
nand U173 (N_173,In_380,N_21);
nand U174 (N_174,In_87,In_25);
nand U175 (N_175,N_81,N_68);
nor U176 (N_176,N_74,N_64);
and U177 (N_177,N_55,In_252);
and U178 (N_178,In_151,N_33);
nor U179 (N_179,In_65,In_139);
and U180 (N_180,N_88,In_479);
or U181 (N_181,N_108,In_229);
nor U182 (N_182,In_240,In_166);
nor U183 (N_183,In_153,In_200);
or U184 (N_184,In_79,N_132);
nor U185 (N_185,N_164,N_48);
nand U186 (N_186,In_216,In_336);
nand U187 (N_187,In_194,N_121);
or U188 (N_188,In_339,In_334);
and U189 (N_189,N_167,In_369);
and U190 (N_190,In_245,N_1);
or U191 (N_191,N_175,In_397);
and U192 (N_192,N_58,N_131);
or U193 (N_193,In_85,In_127);
nor U194 (N_194,In_73,N_47);
or U195 (N_195,N_5,N_32);
nor U196 (N_196,In_219,N_38);
nor U197 (N_197,In_462,In_40);
nand U198 (N_198,In_465,N_75);
nand U199 (N_199,N_169,In_316);
and U200 (N_200,In_401,In_249);
or U201 (N_201,In_56,N_126);
nor U202 (N_202,N_97,In_142);
nor U203 (N_203,In_327,N_25);
xnor U204 (N_204,In_95,In_154);
nand U205 (N_205,N_144,In_408);
nor U206 (N_206,In_81,In_253);
nand U207 (N_207,N_28,In_186);
and U208 (N_208,In_354,In_140);
nor U209 (N_209,N_176,N_162);
nor U210 (N_210,In_213,In_69);
or U211 (N_211,In_499,In_470);
nor U212 (N_212,In_61,In_299);
or U213 (N_213,In_309,N_62);
and U214 (N_214,In_351,N_128);
or U215 (N_215,N_77,In_8);
and U216 (N_216,N_37,N_124);
nand U217 (N_217,In_212,In_459);
nand U218 (N_218,N_18,In_298);
nand U219 (N_219,In_39,In_458);
and U220 (N_220,N_139,N_82);
nand U221 (N_221,N_12,In_237);
nand U222 (N_222,N_178,In_228);
and U223 (N_223,In_363,In_289);
and U224 (N_224,In_320,In_280);
or U225 (N_225,N_168,N_3);
nand U226 (N_226,In_371,N_35);
or U227 (N_227,N_52,In_159);
and U228 (N_228,N_155,In_125);
or U229 (N_229,N_120,N_103);
nand U230 (N_230,In_204,In_428);
and U231 (N_231,In_475,N_148);
and U232 (N_232,In_374,In_355);
nor U233 (N_233,In_411,N_99);
nor U234 (N_234,In_409,In_481);
or U235 (N_235,N_137,In_392);
and U236 (N_236,In_34,N_130);
nand U237 (N_237,In_68,In_448);
or U238 (N_238,In_171,N_106);
and U239 (N_239,N_14,In_115);
nor U240 (N_240,In_466,N_222);
nor U241 (N_241,N_95,In_282);
and U242 (N_242,N_174,In_195);
nand U243 (N_243,In_162,N_79);
and U244 (N_244,In_331,In_80);
nand U245 (N_245,N_238,In_41);
nand U246 (N_246,In_135,N_190);
or U247 (N_247,N_84,N_206);
nor U248 (N_248,N_4,N_142);
nor U249 (N_249,N_104,N_180);
nand U250 (N_250,N_232,N_110);
nand U251 (N_251,N_50,N_44);
nor U252 (N_252,N_29,In_98);
nand U253 (N_253,In_128,N_217);
or U254 (N_254,In_199,In_188);
and U255 (N_255,N_234,In_260);
nand U256 (N_256,N_40,In_147);
or U257 (N_257,N_239,In_347);
or U258 (N_258,N_150,N_233);
xor U259 (N_259,In_102,N_225);
or U260 (N_260,N_199,N_61);
and U261 (N_261,In_275,In_467);
and U262 (N_262,In_442,N_177);
nand U263 (N_263,In_148,N_186);
nor U264 (N_264,In_156,In_329);
nand U265 (N_265,N_163,N_191);
and U266 (N_266,N_149,N_91);
and U267 (N_267,N_189,N_229);
nand U268 (N_268,In_110,N_96);
nor U269 (N_269,In_286,N_202);
and U270 (N_270,N_160,In_55);
and U271 (N_271,N_182,In_417);
nand U272 (N_272,In_235,N_147);
nand U273 (N_273,In_1,N_165);
nand U274 (N_274,N_136,In_77);
or U275 (N_275,In_368,In_297);
and U276 (N_276,N_107,N_166);
nor U277 (N_277,N_123,N_111);
and U278 (N_278,N_22,N_0);
and U279 (N_279,In_118,In_344);
xnor U280 (N_280,N_195,N_109);
or U281 (N_281,In_315,In_131);
and U282 (N_282,In_433,N_101);
or U283 (N_283,N_70,N_135);
or U284 (N_284,In_450,N_172);
nor U285 (N_285,N_141,In_452);
or U286 (N_286,N_231,N_6);
and U287 (N_287,N_112,In_402);
or U288 (N_288,N_122,In_464);
nor U289 (N_289,In_396,N_86);
nand U290 (N_290,In_490,In_310);
nand U291 (N_291,In_306,In_247);
and U292 (N_292,N_67,N_138);
or U293 (N_293,N_146,N_192);
nand U294 (N_294,N_187,N_205);
and U295 (N_295,N_201,N_159);
nand U296 (N_296,N_204,In_16);
nand U297 (N_297,N_24,In_283);
nand U298 (N_298,N_78,In_357);
nand U299 (N_299,In_435,In_290);
or U300 (N_300,N_227,N_212);
nand U301 (N_301,N_197,In_181);
nand U302 (N_302,In_447,N_241);
nor U303 (N_303,N_243,N_157);
nor U304 (N_304,In_281,In_400);
nand U305 (N_305,N_170,In_201);
nor U306 (N_306,N_299,N_127);
or U307 (N_307,N_237,N_210);
or U308 (N_308,N_198,N_208);
and U309 (N_309,N_216,N_242);
nand U310 (N_310,N_60,N_219);
nand U311 (N_311,In_304,N_252);
nor U312 (N_312,N_98,N_113);
nand U313 (N_313,N_255,N_280);
or U314 (N_314,N_184,N_213);
nor U315 (N_315,N_275,N_161);
nand U316 (N_316,N_117,N_179);
nor U317 (N_317,N_193,In_244);
xor U318 (N_318,N_269,N_271);
and U319 (N_319,In_0,N_272);
nand U320 (N_320,N_277,In_86);
or U321 (N_321,N_220,N_223);
or U322 (N_322,In_322,In_211);
and U323 (N_323,N_188,N_218);
or U324 (N_324,N_289,In_377);
and U325 (N_325,In_393,N_285);
or U326 (N_326,N_288,N_283);
or U327 (N_327,N_134,N_265);
or U328 (N_328,N_295,N_129);
or U329 (N_329,In_358,N_273);
nor U330 (N_330,N_260,N_262);
and U331 (N_331,In_221,N_125);
nor U332 (N_332,N_63,N_72);
and U333 (N_333,N_39,N_118);
nor U334 (N_334,In_437,In_350);
nor U335 (N_335,In_108,In_270);
xor U336 (N_336,N_226,N_173);
or U337 (N_337,N_153,N_292);
nand U338 (N_338,N_264,In_496);
or U339 (N_339,In_224,N_256);
nand U340 (N_340,In_365,In_429);
and U341 (N_341,In_484,In_196);
and U342 (N_342,N_297,In_333);
nand U343 (N_343,N_247,N_298);
and U344 (N_344,N_282,N_251);
or U345 (N_345,N_263,In_259);
or U346 (N_346,N_66,N_181);
nor U347 (N_347,In_24,N_171);
nor U348 (N_348,N_215,In_340);
and U349 (N_349,N_293,In_378);
and U350 (N_350,In_445,N_143);
nor U351 (N_351,N_258,N_257);
nand U352 (N_352,In_176,N_151);
or U353 (N_353,In_174,N_291);
nor U354 (N_354,N_87,In_64);
nor U355 (N_355,N_250,N_224);
and U356 (N_356,N_281,N_268);
nand U357 (N_357,N_253,In_145);
or U358 (N_358,N_259,In_349);
or U359 (N_359,In_92,N_19);
and U360 (N_360,In_106,N_41);
nor U361 (N_361,N_357,N_306);
or U362 (N_362,N_65,In_455);
nor U363 (N_363,N_351,N_240);
or U364 (N_364,N_326,N_305);
nor U365 (N_365,N_350,N_156);
nor U366 (N_366,N_203,N_278);
and U367 (N_367,N_302,N_244);
nor U368 (N_368,In_146,N_185);
nand U369 (N_369,In_478,N_279);
or U370 (N_370,N_183,N_266);
or U371 (N_371,N_80,N_59);
nand U372 (N_372,N_246,N_319);
nand U373 (N_373,In_312,N_294);
nor U374 (N_374,In_121,In_49);
nor U375 (N_375,N_154,N_328);
nand U376 (N_376,N_194,N_316);
or U377 (N_377,In_112,In_492);
and U378 (N_378,N_356,In_233);
nor U379 (N_379,N_355,N_152);
nand U380 (N_380,N_330,N_300);
or U381 (N_381,N_347,N_140);
and U382 (N_382,N_286,N_344);
or U383 (N_383,N_230,N_335);
or U384 (N_384,N_318,N_274);
or U385 (N_385,N_320,N_327);
or U386 (N_386,N_248,N_329);
and U387 (N_387,N_236,N_304);
or U388 (N_388,N_287,N_290);
or U389 (N_389,N_196,N_235);
nand U390 (N_390,In_267,N_309);
or U391 (N_391,N_270,N_359);
and U392 (N_392,N_337,N_339);
nand U393 (N_393,In_6,N_349);
nor U394 (N_394,N_308,N_346);
nand U395 (N_395,N_46,N_145);
and U396 (N_396,In_178,In_469);
or U397 (N_397,N_343,N_207);
nand U398 (N_398,N_322,N_313);
and U399 (N_399,N_211,In_443);
nand U400 (N_400,N_334,N_303);
and U401 (N_401,In_97,N_341);
nor U402 (N_402,N_333,N_317);
nand U403 (N_403,N_296,In_239);
or U404 (N_404,N_332,N_301);
or U405 (N_405,N_276,In_416);
nand U406 (N_406,N_358,In_48);
nor U407 (N_407,In_324,N_133);
nand U408 (N_408,N_342,N_323);
or U409 (N_409,N_89,N_340);
or U410 (N_410,N_324,N_315);
and U411 (N_411,In_274,N_209);
nand U412 (N_412,In_325,N_116);
and U413 (N_413,N_311,N_352);
or U414 (N_414,N_321,N_249);
nor U415 (N_415,N_307,N_228);
and U416 (N_416,N_348,In_109);
or U417 (N_417,N_325,N_284);
or U418 (N_418,In_424,N_267);
nand U419 (N_419,N_214,N_221);
nor U420 (N_420,N_380,N_409);
nor U421 (N_421,In_116,N_398);
nand U422 (N_422,N_92,N_365);
nor U423 (N_423,N_362,N_368);
or U424 (N_424,N_367,N_415);
nor U425 (N_425,N_401,N_381);
or U426 (N_426,N_418,N_200);
nand U427 (N_427,N_387,In_256);
nand U428 (N_428,N_372,N_384);
or U429 (N_429,N_371,N_394);
nor U430 (N_430,N_416,In_394);
nor U431 (N_431,N_314,N_312);
nand U432 (N_432,N_361,N_386);
xnor U433 (N_433,N_392,N_374);
and U434 (N_434,N_245,N_366);
or U435 (N_435,N_389,N_405);
nor U436 (N_436,N_331,N_345);
and U437 (N_437,N_399,N_375);
and U438 (N_438,N_310,N_364);
nand U439 (N_439,N_377,In_63);
and U440 (N_440,N_390,N_376);
nand U441 (N_441,N_417,N_419);
nand U442 (N_442,N_158,N_402);
and U443 (N_443,N_412,N_370);
or U444 (N_444,N_378,N_369);
and U445 (N_445,N_353,N_414);
nand U446 (N_446,N_385,N_254);
nand U447 (N_447,N_338,N_261);
or U448 (N_448,N_76,N_393);
nor U449 (N_449,N_406,N_397);
nor U450 (N_450,N_410,N_403);
and U451 (N_451,N_411,N_407);
nor U452 (N_452,N_336,N_383);
or U453 (N_453,N_396,N_379);
and U454 (N_454,N_382,N_373);
or U455 (N_455,N_413,N_388);
nand U456 (N_456,N_395,N_363);
nor U457 (N_457,N_408,N_391);
and U458 (N_458,N_404,N_354);
and U459 (N_459,N_400,N_360);
or U460 (N_460,N_369,N_261);
nor U461 (N_461,N_388,N_407);
and U462 (N_462,N_261,N_372);
nand U463 (N_463,N_360,N_200);
and U464 (N_464,N_398,N_411);
or U465 (N_465,N_375,N_405);
nor U466 (N_466,N_407,N_380);
or U467 (N_467,N_410,N_331);
nand U468 (N_468,N_377,N_331);
or U469 (N_469,N_394,N_379);
and U470 (N_470,In_256,N_354);
or U471 (N_471,N_408,N_409);
and U472 (N_472,N_411,N_374);
nand U473 (N_473,N_380,N_375);
or U474 (N_474,N_418,N_408);
or U475 (N_475,N_76,N_314);
or U476 (N_476,N_374,In_116);
or U477 (N_477,N_374,N_400);
nor U478 (N_478,N_416,N_368);
nor U479 (N_479,N_389,N_200);
nand U480 (N_480,N_428,N_478);
and U481 (N_481,N_476,N_452);
and U482 (N_482,N_443,N_425);
or U483 (N_483,N_468,N_433);
nor U484 (N_484,N_451,N_436);
nor U485 (N_485,N_470,N_474);
and U486 (N_486,N_465,N_455);
nand U487 (N_487,N_466,N_467);
and U488 (N_488,N_460,N_462);
nand U489 (N_489,N_472,N_438);
or U490 (N_490,N_449,N_434);
or U491 (N_491,N_458,N_437);
nor U492 (N_492,N_473,N_477);
nor U493 (N_493,N_439,N_464);
and U494 (N_494,N_450,N_456);
or U495 (N_495,N_479,N_475);
and U496 (N_496,N_431,N_432);
and U497 (N_497,N_471,N_454);
nand U498 (N_498,N_444,N_429);
or U499 (N_499,N_426,N_435);
and U500 (N_500,N_463,N_422);
or U501 (N_501,N_457,N_427);
nor U502 (N_502,N_459,N_442);
or U503 (N_503,N_420,N_424);
nor U504 (N_504,N_430,N_448);
and U505 (N_505,N_440,N_441);
and U506 (N_506,N_469,N_446);
or U507 (N_507,N_423,N_421);
and U508 (N_508,N_447,N_445);
nand U509 (N_509,N_461,N_453);
nor U510 (N_510,N_424,N_475);
nand U511 (N_511,N_440,N_472);
nor U512 (N_512,N_446,N_455);
and U513 (N_513,N_475,N_449);
or U514 (N_514,N_422,N_433);
and U515 (N_515,N_447,N_469);
nand U516 (N_516,N_449,N_421);
or U517 (N_517,N_424,N_437);
and U518 (N_518,N_430,N_477);
nor U519 (N_519,N_463,N_444);
and U520 (N_520,N_476,N_464);
nor U521 (N_521,N_452,N_471);
nor U522 (N_522,N_469,N_439);
nor U523 (N_523,N_424,N_460);
nand U524 (N_524,N_447,N_436);
and U525 (N_525,N_430,N_466);
nand U526 (N_526,N_455,N_430);
nand U527 (N_527,N_433,N_432);
nor U528 (N_528,N_431,N_474);
nor U529 (N_529,N_479,N_422);
or U530 (N_530,N_441,N_422);
and U531 (N_531,N_469,N_453);
or U532 (N_532,N_461,N_431);
nand U533 (N_533,N_437,N_457);
nand U534 (N_534,N_434,N_473);
nand U535 (N_535,N_436,N_478);
or U536 (N_536,N_443,N_469);
and U537 (N_537,N_428,N_438);
nand U538 (N_538,N_468,N_459);
and U539 (N_539,N_443,N_431);
or U540 (N_540,N_510,N_499);
nand U541 (N_541,N_500,N_537);
or U542 (N_542,N_483,N_492);
nand U543 (N_543,N_505,N_528);
nand U544 (N_544,N_530,N_496);
and U545 (N_545,N_535,N_497);
nand U546 (N_546,N_490,N_498);
or U547 (N_547,N_495,N_489);
nor U548 (N_548,N_484,N_506);
nand U549 (N_549,N_526,N_508);
nand U550 (N_550,N_501,N_518);
xnor U551 (N_551,N_488,N_524);
nand U552 (N_552,N_482,N_487);
and U553 (N_553,N_480,N_533);
nand U554 (N_554,N_502,N_491);
or U555 (N_555,N_515,N_523);
nand U556 (N_556,N_521,N_522);
and U557 (N_557,N_517,N_514);
or U558 (N_558,N_531,N_529);
and U559 (N_559,N_532,N_481);
and U560 (N_560,N_516,N_511);
nand U561 (N_561,N_493,N_507);
nand U562 (N_562,N_485,N_486);
nand U563 (N_563,N_538,N_539);
and U564 (N_564,N_513,N_494);
and U565 (N_565,N_503,N_519);
nor U566 (N_566,N_525,N_504);
and U567 (N_567,N_512,N_527);
and U568 (N_568,N_534,N_520);
nand U569 (N_569,N_536,N_509);
nand U570 (N_570,N_511,N_523);
or U571 (N_571,N_533,N_535);
nand U572 (N_572,N_536,N_507);
nor U573 (N_573,N_495,N_490);
and U574 (N_574,N_514,N_507);
or U575 (N_575,N_525,N_505);
nand U576 (N_576,N_518,N_529);
nor U577 (N_577,N_493,N_516);
nor U578 (N_578,N_482,N_491);
nand U579 (N_579,N_508,N_503);
and U580 (N_580,N_534,N_526);
or U581 (N_581,N_485,N_519);
or U582 (N_582,N_526,N_512);
or U583 (N_583,N_490,N_527);
or U584 (N_584,N_488,N_482);
or U585 (N_585,N_534,N_480);
and U586 (N_586,N_526,N_495);
xnor U587 (N_587,N_528,N_500);
nor U588 (N_588,N_496,N_529);
nor U589 (N_589,N_495,N_504);
xnor U590 (N_590,N_524,N_487);
nand U591 (N_591,N_494,N_514);
nor U592 (N_592,N_490,N_522);
or U593 (N_593,N_507,N_535);
nand U594 (N_594,N_538,N_529);
or U595 (N_595,N_495,N_492);
and U596 (N_596,N_538,N_482);
nor U597 (N_597,N_523,N_500);
nand U598 (N_598,N_538,N_533);
nand U599 (N_599,N_496,N_536);
or U600 (N_600,N_575,N_554);
nand U601 (N_601,N_572,N_598);
or U602 (N_602,N_543,N_552);
nand U603 (N_603,N_591,N_541);
and U604 (N_604,N_563,N_585);
nor U605 (N_605,N_567,N_558);
or U606 (N_606,N_553,N_556);
nand U607 (N_607,N_562,N_548);
nand U608 (N_608,N_540,N_577);
nand U609 (N_609,N_549,N_544);
and U610 (N_610,N_586,N_593);
nand U611 (N_611,N_599,N_597);
or U612 (N_612,N_596,N_566);
nor U613 (N_613,N_564,N_588);
and U614 (N_614,N_550,N_560);
nor U615 (N_615,N_569,N_580);
and U616 (N_616,N_555,N_584);
nand U617 (N_617,N_568,N_590);
nor U618 (N_618,N_565,N_557);
nand U619 (N_619,N_579,N_578);
nand U620 (N_620,N_576,N_581);
and U621 (N_621,N_571,N_582);
nor U622 (N_622,N_559,N_587);
and U623 (N_623,N_570,N_573);
or U624 (N_624,N_595,N_592);
or U625 (N_625,N_547,N_594);
and U626 (N_626,N_546,N_583);
nand U627 (N_627,N_574,N_589);
nand U628 (N_628,N_551,N_545);
nand U629 (N_629,N_561,N_542);
nor U630 (N_630,N_546,N_584);
and U631 (N_631,N_569,N_585);
nand U632 (N_632,N_548,N_564);
nor U633 (N_633,N_559,N_597);
or U634 (N_634,N_543,N_576);
nor U635 (N_635,N_569,N_584);
and U636 (N_636,N_544,N_568);
nand U637 (N_637,N_590,N_588);
nand U638 (N_638,N_546,N_586);
or U639 (N_639,N_586,N_543);
nand U640 (N_640,N_566,N_554);
nand U641 (N_641,N_583,N_586);
and U642 (N_642,N_543,N_591);
nand U643 (N_643,N_550,N_586);
nand U644 (N_644,N_563,N_587);
and U645 (N_645,N_598,N_590);
nor U646 (N_646,N_559,N_599);
or U647 (N_647,N_579,N_581);
and U648 (N_648,N_575,N_577);
and U649 (N_649,N_549,N_589);
and U650 (N_650,N_554,N_570);
and U651 (N_651,N_563,N_558);
nand U652 (N_652,N_562,N_541);
and U653 (N_653,N_557,N_587);
or U654 (N_654,N_570,N_594);
or U655 (N_655,N_589,N_559);
nand U656 (N_656,N_564,N_589);
or U657 (N_657,N_549,N_550);
or U658 (N_658,N_599,N_546);
or U659 (N_659,N_589,N_569);
nor U660 (N_660,N_650,N_602);
or U661 (N_661,N_651,N_652);
or U662 (N_662,N_644,N_611);
and U663 (N_663,N_659,N_636);
or U664 (N_664,N_653,N_614);
or U665 (N_665,N_638,N_620);
nor U666 (N_666,N_641,N_631);
nor U667 (N_667,N_654,N_643);
nand U668 (N_668,N_633,N_626);
nor U669 (N_669,N_601,N_657);
nand U670 (N_670,N_608,N_649);
nand U671 (N_671,N_618,N_612);
nor U672 (N_672,N_645,N_634);
nor U673 (N_673,N_622,N_632);
nand U674 (N_674,N_621,N_640);
nand U675 (N_675,N_642,N_604);
nand U676 (N_676,N_616,N_628);
and U677 (N_677,N_623,N_610);
and U678 (N_678,N_639,N_615);
and U679 (N_679,N_624,N_629);
and U680 (N_680,N_646,N_635);
and U681 (N_681,N_605,N_613);
and U682 (N_682,N_617,N_619);
or U683 (N_683,N_606,N_609);
and U684 (N_684,N_647,N_627);
or U685 (N_685,N_656,N_658);
nor U686 (N_686,N_630,N_648);
nand U687 (N_687,N_607,N_600);
and U688 (N_688,N_603,N_637);
nor U689 (N_689,N_655,N_625);
and U690 (N_690,N_658,N_600);
nor U691 (N_691,N_635,N_615);
nor U692 (N_692,N_643,N_627);
and U693 (N_693,N_650,N_605);
or U694 (N_694,N_626,N_601);
nor U695 (N_695,N_618,N_659);
nor U696 (N_696,N_658,N_618);
or U697 (N_697,N_602,N_620);
and U698 (N_698,N_619,N_610);
and U699 (N_699,N_647,N_640);
nand U700 (N_700,N_658,N_643);
nor U701 (N_701,N_655,N_606);
nand U702 (N_702,N_641,N_614);
nand U703 (N_703,N_651,N_621);
nand U704 (N_704,N_621,N_647);
nor U705 (N_705,N_638,N_642);
nor U706 (N_706,N_658,N_657);
and U707 (N_707,N_637,N_656);
nor U708 (N_708,N_607,N_603);
nor U709 (N_709,N_633,N_637);
nor U710 (N_710,N_626,N_639);
nand U711 (N_711,N_644,N_634);
nor U712 (N_712,N_658,N_632);
and U713 (N_713,N_604,N_600);
and U714 (N_714,N_632,N_659);
or U715 (N_715,N_649,N_634);
and U716 (N_716,N_602,N_659);
or U717 (N_717,N_600,N_650);
or U718 (N_718,N_624,N_620);
and U719 (N_719,N_626,N_605);
nand U720 (N_720,N_710,N_680);
nor U721 (N_721,N_668,N_691);
nand U722 (N_722,N_719,N_706);
and U723 (N_723,N_699,N_684);
nor U724 (N_724,N_667,N_663);
nand U725 (N_725,N_716,N_709);
nor U726 (N_726,N_687,N_703);
and U727 (N_727,N_712,N_660);
and U728 (N_728,N_670,N_665);
nand U729 (N_729,N_672,N_713);
or U730 (N_730,N_696,N_689);
or U731 (N_731,N_682,N_679);
nand U732 (N_732,N_661,N_681);
and U733 (N_733,N_698,N_714);
nor U734 (N_734,N_675,N_666);
nand U735 (N_735,N_707,N_705);
nor U736 (N_736,N_683,N_694);
nand U737 (N_737,N_690,N_717);
nand U738 (N_738,N_711,N_685);
or U739 (N_739,N_686,N_697);
nand U740 (N_740,N_673,N_702);
nand U741 (N_741,N_693,N_715);
and U742 (N_742,N_704,N_674);
and U743 (N_743,N_701,N_669);
or U744 (N_744,N_708,N_677);
nand U745 (N_745,N_700,N_692);
nand U746 (N_746,N_662,N_676);
nor U747 (N_747,N_664,N_688);
nand U748 (N_748,N_695,N_678);
and U749 (N_749,N_671,N_718);
nand U750 (N_750,N_714,N_671);
nand U751 (N_751,N_670,N_709);
nand U752 (N_752,N_696,N_687);
nor U753 (N_753,N_673,N_710);
and U754 (N_754,N_716,N_686);
or U755 (N_755,N_672,N_719);
xnor U756 (N_756,N_667,N_688);
and U757 (N_757,N_713,N_691);
nand U758 (N_758,N_697,N_701);
nor U759 (N_759,N_715,N_714);
and U760 (N_760,N_710,N_678);
nor U761 (N_761,N_695,N_693);
nand U762 (N_762,N_693,N_689);
nor U763 (N_763,N_705,N_688);
or U764 (N_764,N_707,N_703);
or U765 (N_765,N_664,N_706);
nand U766 (N_766,N_690,N_704);
or U767 (N_767,N_688,N_715);
nand U768 (N_768,N_690,N_673);
or U769 (N_769,N_708,N_701);
or U770 (N_770,N_712,N_669);
nand U771 (N_771,N_716,N_668);
and U772 (N_772,N_715,N_689);
xor U773 (N_773,N_697,N_660);
or U774 (N_774,N_669,N_715);
nor U775 (N_775,N_703,N_666);
or U776 (N_776,N_716,N_670);
and U777 (N_777,N_699,N_716);
and U778 (N_778,N_670,N_686);
nand U779 (N_779,N_683,N_664);
nor U780 (N_780,N_760,N_739);
nand U781 (N_781,N_769,N_773);
nor U782 (N_782,N_774,N_765);
or U783 (N_783,N_761,N_766);
and U784 (N_784,N_771,N_749);
and U785 (N_785,N_736,N_724);
nor U786 (N_786,N_758,N_740);
and U787 (N_787,N_726,N_756);
or U788 (N_788,N_779,N_751);
and U789 (N_789,N_764,N_738);
nor U790 (N_790,N_746,N_770);
nor U791 (N_791,N_750,N_763);
nand U792 (N_792,N_747,N_730);
and U793 (N_793,N_733,N_755);
xor U794 (N_794,N_775,N_748);
or U795 (N_795,N_737,N_725);
nor U796 (N_796,N_752,N_745);
nand U797 (N_797,N_757,N_721);
nand U798 (N_798,N_731,N_744);
nand U799 (N_799,N_778,N_777);
nand U800 (N_800,N_772,N_729);
or U801 (N_801,N_728,N_768);
nor U802 (N_802,N_767,N_776);
or U803 (N_803,N_732,N_762);
xor U804 (N_804,N_759,N_720);
and U805 (N_805,N_753,N_742);
nor U806 (N_806,N_743,N_754);
and U807 (N_807,N_741,N_735);
nand U808 (N_808,N_722,N_727);
nand U809 (N_809,N_734,N_723);
or U810 (N_810,N_732,N_735);
nor U811 (N_811,N_751,N_743);
nor U812 (N_812,N_736,N_735);
nand U813 (N_813,N_730,N_779);
and U814 (N_814,N_734,N_721);
nand U815 (N_815,N_738,N_775);
nor U816 (N_816,N_730,N_773);
and U817 (N_817,N_760,N_746);
xnor U818 (N_818,N_732,N_720);
and U819 (N_819,N_758,N_744);
or U820 (N_820,N_747,N_733);
nand U821 (N_821,N_720,N_731);
nor U822 (N_822,N_769,N_734);
nand U823 (N_823,N_728,N_772);
and U824 (N_824,N_723,N_738);
nor U825 (N_825,N_732,N_775);
nand U826 (N_826,N_740,N_731);
nor U827 (N_827,N_741,N_730);
and U828 (N_828,N_744,N_739);
and U829 (N_829,N_766,N_737);
and U830 (N_830,N_767,N_769);
nand U831 (N_831,N_725,N_761);
and U832 (N_832,N_753,N_750);
and U833 (N_833,N_736,N_745);
and U834 (N_834,N_741,N_748);
or U835 (N_835,N_730,N_752);
nand U836 (N_836,N_748,N_750);
nor U837 (N_837,N_764,N_747);
or U838 (N_838,N_762,N_724);
nor U839 (N_839,N_735,N_769);
and U840 (N_840,N_801,N_825);
and U841 (N_841,N_816,N_826);
and U842 (N_842,N_824,N_790);
nor U843 (N_843,N_791,N_832);
and U844 (N_844,N_784,N_812);
or U845 (N_845,N_782,N_807);
and U846 (N_846,N_786,N_815);
nor U847 (N_847,N_796,N_811);
and U848 (N_848,N_835,N_785);
and U849 (N_849,N_802,N_799);
nor U850 (N_850,N_836,N_819);
or U851 (N_851,N_820,N_795);
and U852 (N_852,N_838,N_794);
and U853 (N_853,N_780,N_837);
nor U854 (N_854,N_797,N_827);
or U855 (N_855,N_813,N_798);
nor U856 (N_856,N_809,N_829);
and U857 (N_857,N_822,N_823);
nand U858 (N_858,N_818,N_803);
and U859 (N_859,N_788,N_800);
nand U860 (N_860,N_828,N_839);
or U861 (N_861,N_830,N_833);
or U862 (N_862,N_792,N_804);
xor U863 (N_863,N_806,N_834);
or U864 (N_864,N_789,N_781);
or U865 (N_865,N_821,N_831);
and U866 (N_866,N_808,N_817);
or U867 (N_867,N_793,N_783);
or U868 (N_868,N_810,N_805);
and U869 (N_869,N_787,N_814);
nand U870 (N_870,N_813,N_784);
or U871 (N_871,N_820,N_829);
and U872 (N_872,N_836,N_811);
nor U873 (N_873,N_791,N_787);
nand U874 (N_874,N_803,N_791);
nor U875 (N_875,N_786,N_839);
or U876 (N_876,N_808,N_807);
and U877 (N_877,N_796,N_828);
nor U878 (N_878,N_824,N_808);
nor U879 (N_879,N_830,N_794);
and U880 (N_880,N_795,N_816);
nor U881 (N_881,N_809,N_821);
or U882 (N_882,N_813,N_791);
nor U883 (N_883,N_830,N_807);
nor U884 (N_884,N_793,N_803);
and U885 (N_885,N_835,N_810);
and U886 (N_886,N_825,N_798);
nand U887 (N_887,N_825,N_805);
nor U888 (N_888,N_827,N_830);
nand U889 (N_889,N_833,N_801);
nor U890 (N_890,N_797,N_789);
nand U891 (N_891,N_812,N_826);
and U892 (N_892,N_801,N_783);
nand U893 (N_893,N_807,N_816);
nor U894 (N_894,N_791,N_819);
nor U895 (N_895,N_830,N_825);
nand U896 (N_896,N_824,N_811);
nor U897 (N_897,N_836,N_788);
and U898 (N_898,N_828,N_826);
nor U899 (N_899,N_792,N_836);
and U900 (N_900,N_875,N_873);
and U901 (N_901,N_872,N_888);
nor U902 (N_902,N_870,N_877);
and U903 (N_903,N_843,N_876);
nor U904 (N_904,N_846,N_887);
nor U905 (N_905,N_866,N_862);
nand U906 (N_906,N_856,N_880);
nand U907 (N_907,N_897,N_871);
nand U908 (N_908,N_869,N_864);
nand U909 (N_909,N_857,N_899);
nor U910 (N_910,N_844,N_885);
nand U911 (N_911,N_859,N_886);
nand U912 (N_912,N_847,N_881);
or U913 (N_913,N_867,N_842);
or U914 (N_914,N_860,N_863);
and U915 (N_915,N_865,N_849);
nor U916 (N_916,N_893,N_895);
and U917 (N_917,N_889,N_884);
or U918 (N_918,N_883,N_879);
nor U919 (N_919,N_850,N_891);
nor U920 (N_920,N_848,N_890);
and U921 (N_921,N_840,N_868);
nand U922 (N_922,N_894,N_898);
or U923 (N_923,N_861,N_855);
or U924 (N_924,N_858,N_854);
nor U925 (N_925,N_845,N_852);
nor U926 (N_926,N_851,N_892);
nand U927 (N_927,N_882,N_853);
nand U928 (N_928,N_841,N_874);
and U929 (N_929,N_896,N_878);
or U930 (N_930,N_899,N_877);
and U931 (N_931,N_843,N_877);
and U932 (N_932,N_877,N_872);
or U933 (N_933,N_894,N_855);
and U934 (N_934,N_896,N_852);
or U935 (N_935,N_861,N_883);
nand U936 (N_936,N_847,N_863);
nand U937 (N_937,N_858,N_842);
or U938 (N_938,N_893,N_871);
nand U939 (N_939,N_856,N_874);
or U940 (N_940,N_868,N_846);
nand U941 (N_941,N_896,N_847);
nand U942 (N_942,N_890,N_889);
nor U943 (N_943,N_860,N_868);
nor U944 (N_944,N_858,N_877);
nor U945 (N_945,N_858,N_859);
nor U946 (N_946,N_848,N_883);
or U947 (N_947,N_899,N_850);
or U948 (N_948,N_847,N_889);
nor U949 (N_949,N_864,N_861);
nand U950 (N_950,N_882,N_886);
nand U951 (N_951,N_857,N_853);
and U952 (N_952,N_845,N_863);
nand U953 (N_953,N_863,N_850);
nand U954 (N_954,N_897,N_841);
and U955 (N_955,N_881,N_891);
nor U956 (N_956,N_860,N_843);
or U957 (N_957,N_846,N_877);
or U958 (N_958,N_857,N_890);
nor U959 (N_959,N_897,N_881);
nor U960 (N_960,N_939,N_919);
or U961 (N_961,N_949,N_915);
nand U962 (N_962,N_913,N_920);
and U963 (N_963,N_931,N_954);
or U964 (N_964,N_922,N_951);
or U965 (N_965,N_943,N_900);
and U966 (N_966,N_953,N_932);
nor U967 (N_967,N_952,N_906);
and U968 (N_968,N_940,N_933);
and U969 (N_969,N_908,N_959);
and U970 (N_970,N_912,N_937);
nor U971 (N_971,N_910,N_930);
nor U972 (N_972,N_934,N_958);
or U973 (N_973,N_942,N_923);
nand U974 (N_974,N_909,N_901);
or U975 (N_975,N_944,N_957);
and U976 (N_976,N_914,N_929);
nor U977 (N_977,N_955,N_947);
nand U978 (N_978,N_924,N_950);
and U979 (N_979,N_911,N_945);
nor U980 (N_980,N_941,N_903);
or U981 (N_981,N_904,N_926);
and U982 (N_982,N_917,N_902);
and U983 (N_983,N_916,N_938);
nor U984 (N_984,N_921,N_907);
nand U985 (N_985,N_928,N_936);
nand U986 (N_986,N_918,N_925);
nand U987 (N_987,N_956,N_927);
or U988 (N_988,N_935,N_905);
and U989 (N_989,N_946,N_948);
nand U990 (N_990,N_948,N_936);
nor U991 (N_991,N_938,N_943);
or U992 (N_992,N_932,N_946);
nand U993 (N_993,N_946,N_938);
or U994 (N_994,N_914,N_923);
and U995 (N_995,N_947,N_952);
nand U996 (N_996,N_941,N_949);
xor U997 (N_997,N_908,N_940);
nand U998 (N_998,N_904,N_916);
nand U999 (N_999,N_950,N_946);
and U1000 (N_1000,N_935,N_953);
and U1001 (N_1001,N_947,N_922);
or U1002 (N_1002,N_924,N_945);
or U1003 (N_1003,N_922,N_953);
nor U1004 (N_1004,N_906,N_931);
or U1005 (N_1005,N_903,N_950);
and U1006 (N_1006,N_903,N_946);
xnor U1007 (N_1007,N_902,N_914);
and U1008 (N_1008,N_927,N_922);
nand U1009 (N_1009,N_917,N_931);
nor U1010 (N_1010,N_933,N_952);
or U1011 (N_1011,N_901,N_933);
nor U1012 (N_1012,N_924,N_930);
or U1013 (N_1013,N_910,N_937);
or U1014 (N_1014,N_931,N_942);
nand U1015 (N_1015,N_941,N_929);
or U1016 (N_1016,N_916,N_949);
nor U1017 (N_1017,N_907,N_925);
nor U1018 (N_1018,N_928,N_911);
or U1019 (N_1019,N_944,N_959);
or U1020 (N_1020,N_963,N_961);
or U1021 (N_1021,N_1013,N_978);
nand U1022 (N_1022,N_1003,N_997);
nand U1023 (N_1023,N_1004,N_994);
nor U1024 (N_1024,N_989,N_990);
nor U1025 (N_1025,N_995,N_972);
nand U1026 (N_1026,N_1010,N_980);
and U1027 (N_1027,N_960,N_971);
and U1028 (N_1028,N_965,N_962);
or U1029 (N_1029,N_964,N_984);
nor U1030 (N_1030,N_981,N_973);
nand U1031 (N_1031,N_1007,N_999);
or U1032 (N_1032,N_1019,N_966);
nand U1033 (N_1033,N_992,N_968);
nand U1034 (N_1034,N_982,N_1014);
nor U1035 (N_1035,N_987,N_1016);
or U1036 (N_1036,N_998,N_977);
and U1037 (N_1037,N_1006,N_1001);
nor U1038 (N_1038,N_988,N_993);
and U1039 (N_1039,N_1012,N_979);
or U1040 (N_1040,N_1002,N_1017);
and U1041 (N_1041,N_986,N_976);
or U1042 (N_1042,N_974,N_1015);
nand U1043 (N_1043,N_969,N_1011);
nor U1044 (N_1044,N_1008,N_1005);
nor U1045 (N_1045,N_1018,N_975);
or U1046 (N_1046,N_983,N_1009);
nand U1047 (N_1047,N_991,N_967);
and U1048 (N_1048,N_1000,N_985);
nor U1049 (N_1049,N_996,N_970);
or U1050 (N_1050,N_967,N_961);
or U1051 (N_1051,N_1002,N_1019);
and U1052 (N_1052,N_1003,N_975);
or U1053 (N_1053,N_1014,N_1001);
nand U1054 (N_1054,N_972,N_993);
nand U1055 (N_1055,N_1010,N_989);
and U1056 (N_1056,N_1014,N_999);
nand U1057 (N_1057,N_983,N_982);
and U1058 (N_1058,N_967,N_1014);
or U1059 (N_1059,N_1004,N_985);
or U1060 (N_1060,N_964,N_962);
nand U1061 (N_1061,N_961,N_993);
nand U1062 (N_1062,N_999,N_977);
nand U1063 (N_1063,N_1008,N_1011);
nand U1064 (N_1064,N_968,N_982);
and U1065 (N_1065,N_1016,N_997);
nand U1066 (N_1066,N_989,N_992);
or U1067 (N_1067,N_1008,N_983);
nand U1068 (N_1068,N_980,N_973);
nand U1069 (N_1069,N_989,N_994);
and U1070 (N_1070,N_1005,N_967);
or U1071 (N_1071,N_1015,N_996);
and U1072 (N_1072,N_1007,N_978);
nor U1073 (N_1073,N_966,N_962);
nor U1074 (N_1074,N_1011,N_988);
nor U1075 (N_1075,N_974,N_967);
nor U1076 (N_1076,N_973,N_972);
nand U1077 (N_1077,N_991,N_973);
and U1078 (N_1078,N_964,N_1004);
nor U1079 (N_1079,N_999,N_1005);
and U1080 (N_1080,N_1033,N_1021);
nand U1081 (N_1081,N_1068,N_1022);
nor U1082 (N_1082,N_1048,N_1026);
or U1083 (N_1083,N_1037,N_1027);
nor U1084 (N_1084,N_1047,N_1076);
nor U1085 (N_1085,N_1071,N_1023);
or U1086 (N_1086,N_1024,N_1043);
and U1087 (N_1087,N_1040,N_1060);
nor U1088 (N_1088,N_1035,N_1046);
nand U1089 (N_1089,N_1053,N_1074);
and U1090 (N_1090,N_1034,N_1059);
nor U1091 (N_1091,N_1025,N_1029);
nor U1092 (N_1092,N_1028,N_1078);
nand U1093 (N_1093,N_1045,N_1063);
or U1094 (N_1094,N_1077,N_1067);
nand U1095 (N_1095,N_1057,N_1061);
and U1096 (N_1096,N_1072,N_1041);
nand U1097 (N_1097,N_1049,N_1070);
and U1098 (N_1098,N_1052,N_1062);
and U1099 (N_1099,N_1036,N_1054);
nand U1100 (N_1100,N_1075,N_1055);
or U1101 (N_1101,N_1044,N_1032);
and U1102 (N_1102,N_1020,N_1079);
nor U1103 (N_1103,N_1065,N_1058);
and U1104 (N_1104,N_1038,N_1073);
nor U1105 (N_1105,N_1051,N_1050);
nor U1106 (N_1106,N_1031,N_1069);
and U1107 (N_1107,N_1042,N_1056);
nand U1108 (N_1108,N_1064,N_1030);
nand U1109 (N_1109,N_1066,N_1039);
nand U1110 (N_1110,N_1061,N_1055);
nand U1111 (N_1111,N_1042,N_1054);
or U1112 (N_1112,N_1035,N_1051);
nand U1113 (N_1113,N_1043,N_1077);
nand U1114 (N_1114,N_1033,N_1042);
and U1115 (N_1115,N_1036,N_1072);
nand U1116 (N_1116,N_1041,N_1065);
nor U1117 (N_1117,N_1026,N_1028);
nor U1118 (N_1118,N_1062,N_1045);
or U1119 (N_1119,N_1061,N_1027);
and U1120 (N_1120,N_1066,N_1048);
or U1121 (N_1121,N_1037,N_1024);
nor U1122 (N_1122,N_1028,N_1037);
and U1123 (N_1123,N_1075,N_1034);
nor U1124 (N_1124,N_1027,N_1035);
nand U1125 (N_1125,N_1069,N_1030);
nand U1126 (N_1126,N_1062,N_1056);
nor U1127 (N_1127,N_1021,N_1038);
and U1128 (N_1128,N_1079,N_1037);
nor U1129 (N_1129,N_1044,N_1064);
and U1130 (N_1130,N_1054,N_1026);
nor U1131 (N_1131,N_1034,N_1033);
or U1132 (N_1132,N_1058,N_1046);
nand U1133 (N_1133,N_1062,N_1033);
nand U1134 (N_1134,N_1073,N_1071);
and U1135 (N_1135,N_1045,N_1064);
nand U1136 (N_1136,N_1025,N_1030);
nand U1137 (N_1137,N_1022,N_1036);
and U1138 (N_1138,N_1052,N_1037);
and U1139 (N_1139,N_1053,N_1023);
nor U1140 (N_1140,N_1131,N_1123);
nor U1141 (N_1141,N_1097,N_1095);
nor U1142 (N_1142,N_1133,N_1135);
or U1143 (N_1143,N_1117,N_1108);
or U1144 (N_1144,N_1084,N_1089);
or U1145 (N_1145,N_1115,N_1101);
nor U1146 (N_1146,N_1091,N_1127);
nor U1147 (N_1147,N_1114,N_1126);
nand U1148 (N_1148,N_1119,N_1116);
or U1149 (N_1149,N_1093,N_1083);
nor U1150 (N_1150,N_1087,N_1138);
nor U1151 (N_1151,N_1085,N_1086);
or U1152 (N_1152,N_1102,N_1082);
or U1153 (N_1153,N_1081,N_1105);
or U1154 (N_1154,N_1100,N_1132);
and U1155 (N_1155,N_1106,N_1094);
nor U1156 (N_1156,N_1096,N_1125);
nor U1157 (N_1157,N_1137,N_1128);
or U1158 (N_1158,N_1099,N_1090);
and U1159 (N_1159,N_1112,N_1111);
and U1160 (N_1160,N_1110,N_1104);
nand U1161 (N_1161,N_1129,N_1113);
nand U1162 (N_1162,N_1109,N_1092);
or U1163 (N_1163,N_1124,N_1120);
nand U1164 (N_1164,N_1098,N_1139);
and U1165 (N_1165,N_1107,N_1121);
and U1166 (N_1166,N_1122,N_1134);
nand U1167 (N_1167,N_1130,N_1118);
and U1168 (N_1168,N_1103,N_1088);
nor U1169 (N_1169,N_1136,N_1080);
nor U1170 (N_1170,N_1107,N_1135);
and U1171 (N_1171,N_1086,N_1116);
and U1172 (N_1172,N_1127,N_1106);
and U1173 (N_1173,N_1085,N_1101);
and U1174 (N_1174,N_1111,N_1099);
and U1175 (N_1175,N_1099,N_1087);
nor U1176 (N_1176,N_1112,N_1100);
nor U1177 (N_1177,N_1090,N_1104);
and U1178 (N_1178,N_1114,N_1133);
or U1179 (N_1179,N_1090,N_1129);
nor U1180 (N_1180,N_1087,N_1081);
nand U1181 (N_1181,N_1087,N_1132);
xnor U1182 (N_1182,N_1137,N_1089);
or U1183 (N_1183,N_1089,N_1096);
nor U1184 (N_1184,N_1097,N_1091);
and U1185 (N_1185,N_1114,N_1112);
nand U1186 (N_1186,N_1137,N_1085);
nand U1187 (N_1187,N_1087,N_1093);
and U1188 (N_1188,N_1108,N_1106);
or U1189 (N_1189,N_1135,N_1104);
nand U1190 (N_1190,N_1091,N_1115);
or U1191 (N_1191,N_1083,N_1117);
nand U1192 (N_1192,N_1088,N_1100);
nand U1193 (N_1193,N_1102,N_1114);
nor U1194 (N_1194,N_1101,N_1118);
nand U1195 (N_1195,N_1083,N_1087);
or U1196 (N_1196,N_1085,N_1113);
and U1197 (N_1197,N_1091,N_1114);
nor U1198 (N_1198,N_1083,N_1134);
and U1199 (N_1199,N_1084,N_1130);
nor U1200 (N_1200,N_1177,N_1142);
nand U1201 (N_1201,N_1180,N_1140);
or U1202 (N_1202,N_1167,N_1199);
and U1203 (N_1203,N_1171,N_1196);
nand U1204 (N_1204,N_1194,N_1190);
or U1205 (N_1205,N_1143,N_1150);
nor U1206 (N_1206,N_1163,N_1181);
and U1207 (N_1207,N_1195,N_1191);
and U1208 (N_1208,N_1182,N_1186);
nand U1209 (N_1209,N_1164,N_1170);
nand U1210 (N_1210,N_1155,N_1189);
and U1211 (N_1211,N_1175,N_1146);
nand U1212 (N_1212,N_1185,N_1162);
nor U1213 (N_1213,N_1148,N_1149);
nor U1214 (N_1214,N_1197,N_1187);
and U1215 (N_1215,N_1188,N_1157);
and U1216 (N_1216,N_1161,N_1184);
and U1217 (N_1217,N_1160,N_1154);
nand U1218 (N_1218,N_1192,N_1173);
nand U1219 (N_1219,N_1141,N_1172);
nor U1220 (N_1220,N_1151,N_1174);
or U1221 (N_1221,N_1147,N_1153);
nand U1222 (N_1222,N_1176,N_1169);
xor U1223 (N_1223,N_1152,N_1156);
nor U1224 (N_1224,N_1178,N_1144);
or U1225 (N_1225,N_1159,N_1168);
nand U1226 (N_1226,N_1166,N_1158);
nand U1227 (N_1227,N_1193,N_1198);
and U1228 (N_1228,N_1165,N_1179);
nor U1229 (N_1229,N_1145,N_1183);
nor U1230 (N_1230,N_1140,N_1199);
nand U1231 (N_1231,N_1154,N_1146);
nor U1232 (N_1232,N_1158,N_1145);
nor U1233 (N_1233,N_1161,N_1179);
and U1234 (N_1234,N_1149,N_1164);
nand U1235 (N_1235,N_1198,N_1189);
nand U1236 (N_1236,N_1156,N_1151);
or U1237 (N_1237,N_1159,N_1167);
nand U1238 (N_1238,N_1170,N_1148);
nor U1239 (N_1239,N_1142,N_1194);
nor U1240 (N_1240,N_1145,N_1160);
nand U1241 (N_1241,N_1185,N_1179);
and U1242 (N_1242,N_1157,N_1143);
nand U1243 (N_1243,N_1192,N_1140);
nand U1244 (N_1244,N_1154,N_1156);
nor U1245 (N_1245,N_1166,N_1184);
and U1246 (N_1246,N_1140,N_1175);
and U1247 (N_1247,N_1144,N_1189);
nor U1248 (N_1248,N_1151,N_1143);
and U1249 (N_1249,N_1165,N_1161);
or U1250 (N_1250,N_1183,N_1169);
or U1251 (N_1251,N_1159,N_1199);
or U1252 (N_1252,N_1147,N_1196);
nor U1253 (N_1253,N_1167,N_1172);
nor U1254 (N_1254,N_1159,N_1145);
and U1255 (N_1255,N_1167,N_1175);
and U1256 (N_1256,N_1188,N_1150);
nand U1257 (N_1257,N_1184,N_1152);
nor U1258 (N_1258,N_1198,N_1188);
nand U1259 (N_1259,N_1178,N_1153);
and U1260 (N_1260,N_1202,N_1242);
and U1261 (N_1261,N_1229,N_1236);
nor U1262 (N_1262,N_1253,N_1252);
nor U1263 (N_1263,N_1208,N_1256);
nand U1264 (N_1264,N_1227,N_1245);
or U1265 (N_1265,N_1218,N_1221);
nand U1266 (N_1266,N_1235,N_1213);
and U1267 (N_1267,N_1222,N_1226);
nor U1268 (N_1268,N_1211,N_1248);
or U1269 (N_1269,N_1205,N_1203);
or U1270 (N_1270,N_1216,N_1206);
nor U1271 (N_1271,N_1234,N_1204);
and U1272 (N_1272,N_1228,N_1217);
or U1273 (N_1273,N_1241,N_1246);
nor U1274 (N_1274,N_1209,N_1220);
and U1275 (N_1275,N_1215,N_1231);
or U1276 (N_1276,N_1230,N_1225);
nand U1277 (N_1277,N_1237,N_1240);
and U1278 (N_1278,N_1249,N_1223);
nand U1279 (N_1279,N_1257,N_1200);
nor U1280 (N_1280,N_1255,N_1224);
nor U1281 (N_1281,N_1214,N_1250);
nor U1282 (N_1282,N_1254,N_1201);
and U1283 (N_1283,N_1259,N_1244);
nor U1284 (N_1284,N_1258,N_1232);
or U1285 (N_1285,N_1251,N_1219);
nor U1286 (N_1286,N_1243,N_1233);
nor U1287 (N_1287,N_1247,N_1239);
nor U1288 (N_1288,N_1212,N_1238);
nand U1289 (N_1289,N_1207,N_1210);
or U1290 (N_1290,N_1240,N_1229);
nor U1291 (N_1291,N_1235,N_1202);
and U1292 (N_1292,N_1219,N_1252);
nor U1293 (N_1293,N_1229,N_1218);
nor U1294 (N_1294,N_1238,N_1249);
or U1295 (N_1295,N_1257,N_1227);
nand U1296 (N_1296,N_1218,N_1236);
nor U1297 (N_1297,N_1200,N_1211);
or U1298 (N_1298,N_1203,N_1218);
and U1299 (N_1299,N_1223,N_1206);
or U1300 (N_1300,N_1215,N_1248);
nand U1301 (N_1301,N_1222,N_1236);
nor U1302 (N_1302,N_1259,N_1210);
or U1303 (N_1303,N_1209,N_1241);
nand U1304 (N_1304,N_1232,N_1202);
nor U1305 (N_1305,N_1219,N_1239);
nand U1306 (N_1306,N_1252,N_1229);
and U1307 (N_1307,N_1247,N_1252);
nor U1308 (N_1308,N_1206,N_1231);
nor U1309 (N_1309,N_1220,N_1225);
or U1310 (N_1310,N_1235,N_1220);
or U1311 (N_1311,N_1209,N_1226);
nand U1312 (N_1312,N_1232,N_1210);
nor U1313 (N_1313,N_1219,N_1215);
or U1314 (N_1314,N_1233,N_1220);
xnor U1315 (N_1315,N_1209,N_1206);
and U1316 (N_1316,N_1229,N_1204);
or U1317 (N_1317,N_1241,N_1206);
nand U1318 (N_1318,N_1258,N_1242);
or U1319 (N_1319,N_1229,N_1241);
nand U1320 (N_1320,N_1266,N_1278);
or U1321 (N_1321,N_1288,N_1303);
or U1322 (N_1322,N_1265,N_1306);
or U1323 (N_1323,N_1284,N_1262);
nor U1324 (N_1324,N_1290,N_1309);
nand U1325 (N_1325,N_1276,N_1314);
nor U1326 (N_1326,N_1298,N_1319);
nor U1327 (N_1327,N_1264,N_1275);
nand U1328 (N_1328,N_1286,N_1279);
nor U1329 (N_1329,N_1277,N_1318);
nor U1330 (N_1330,N_1263,N_1307);
nor U1331 (N_1331,N_1260,N_1268);
nor U1332 (N_1332,N_1289,N_1305);
or U1333 (N_1333,N_1274,N_1302);
and U1334 (N_1334,N_1273,N_1297);
nand U1335 (N_1335,N_1316,N_1300);
and U1336 (N_1336,N_1317,N_1301);
nor U1337 (N_1337,N_1315,N_1311);
nor U1338 (N_1338,N_1313,N_1312);
nand U1339 (N_1339,N_1283,N_1296);
and U1340 (N_1340,N_1271,N_1294);
nand U1341 (N_1341,N_1295,N_1293);
nand U1342 (N_1342,N_1292,N_1291);
and U1343 (N_1343,N_1287,N_1281);
and U1344 (N_1344,N_1267,N_1299);
or U1345 (N_1345,N_1304,N_1270);
nor U1346 (N_1346,N_1272,N_1261);
or U1347 (N_1347,N_1282,N_1269);
nand U1348 (N_1348,N_1285,N_1310);
or U1349 (N_1349,N_1308,N_1280);
or U1350 (N_1350,N_1278,N_1284);
nor U1351 (N_1351,N_1309,N_1262);
xor U1352 (N_1352,N_1319,N_1291);
nor U1353 (N_1353,N_1305,N_1267);
nand U1354 (N_1354,N_1273,N_1287);
or U1355 (N_1355,N_1288,N_1305);
nand U1356 (N_1356,N_1308,N_1288);
nor U1357 (N_1357,N_1297,N_1283);
nand U1358 (N_1358,N_1296,N_1266);
and U1359 (N_1359,N_1310,N_1297);
and U1360 (N_1360,N_1270,N_1276);
nor U1361 (N_1361,N_1271,N_1286);
or U1362 (N_1362,N_1317,N_1277);
nand U1363 (N_1363,N_1296,N_1265);
or U1364 (N_1364,N_1265,N_1312);
or U1365 (N_1365,N_1276,N_1262);
nor U1366 (N_1366,N_1260,N_1316);
and U1367 (N_1367,N_1312,N_1261);
or U1368 (N_1368,N_1267,N_1319);
or U1369 (N_1369,N_1267,N_1304);
or U1370 (N_1370,N_1282,N_1296);
nand U1371 (N_1371,N_1261,N_1318);
and U1372 (N_1372,N_1306,N_1290);
nor U1373 (N_1373,N_1269,N_1315);
or U1374 (N_1374,N_1266,N_1310);
nand U1375 (N_1375,N_1317,N_1285);
and U1376 (N_1376,N_1298,N_1301);
nand U1377 (N_1377,N_1270,N_1295);
or U1378 (N_1378,N_1300,N_1275);
nor U1379 (N_1379,N_1281,N_1269);
or U1380 (N_1380,N_1324,N_1323);
nor U1381 (N_1381,N_1334,N_1348);
nor U1382 (N_1382,N_1343,N_1350);
and U1383 (N_1383,N_1370,N_1353);
nor U1384 (N_1384,N_1341,N_1358);
and U1385 (N_1385,N_1378,N_1347);
and U1386 (N_1386,N_1373,N_1364);
nor U1387 (N_1387,N_1376,N_1321);
nor U1388 (N_1388,N_1344,N_1331);
and U1389 (N_1389,N_1379,N_1366);
nor U1390 (N_1390,N_1375,N_1371);
and U1391 (N_1391,N_1342,N_1363);
nor U1392 (N_1392,N_1356,N_1336);
or U1393 (N_1393,N_1368,N_1352);
nor U1394 (N_1394,N_1328,N_1322);
nor U1395 (N_1395,N_1330,N_1345);
and U1396 (N_1396,N_1335,N_1377);
or U1397 (N_1397,N_1354,N_1325);
and U1398 (N_1398,N_1337,N_1357);
nand U1399 (N_1399,N_1326,N_1332);
and U1400 (N_1400,N_1327,N_1365);
or U1401 (N_1401,N_1349,N_1372);
nand U1402 (N_1402,N_1333,N_1369);
nor U1403 (N_1403,N_1359,N_1340);
nand U1404 (N_1404,N_1320,N_1361);
and U1405 (N_1405,N_1346,N_1338);
nor U1406 (N_1406,N_1329,N_1360);
and U1407 (N_1407,N_1362,N_1351);
and U1408 (N_1408,N_1355,N_1367);
nand U1409 (N_1409,N_1339,N_1374);
or U1410 (N_1410,N_1343,N_1373);
nor U1411 (N_1411,N_1367,N_1335);
or U1412 (N_1412,N_1366,N_1329);
nor U1413 (N_1413,N_1358,N_1322);
nor U1414 (N_1414,N_1342,N_1335);
or U1415 (N_1415,N_1345,N_1375);
nand U1416 (N_1416,N_1350,N_1334);
or U1417 (N_1417,N_1332,N_1355);
and U1418 (N_1418,N_1340,N_1342);
nor U1419 (N_1419,N_1378,N_1345);
nor U1420 (N_1420,N_1325,N_1321);
and U1421 (N_1421,N_1366,N_1330);
nor U1422 (N_1422,N_1343,N_1323);
and U1423 (N_1423,N_1361,N_1339);
nand U1424 (N_1424,N_1337,N_1321);
and U1425 (N_1425,N_1364,N_1367);
nor U1426 (N_1426,N_1370,N_1362);
nand U1427 (N_1427,N_1364,N_1333);
nand U1428 (N_1428,N_1339,N_1337);
nand U1429 (N_1429,N_1350,N_1356);
and U1430 (N_1430,N_1357,N_1320);
nor U1431 (N_1431,N_1366,N_1361);
or U1432 (N_1432,N_1373,N_1355);
nand U1433 (N_1433,N_1328,N_1354);
nor U1434 (N_1434,N_1327,N_1378);
and U1435 (N_1435,N_1320,N_1341);
or U1436 (N_1436,N_1358,N_1329);
and U1437 (N_1437,N_1349,N_1325);
nand U1438 (N_1438,N_1339,N_1330);
nand U1439 (N_1439,N_1343,N_1349);
or U1440 (N_1440,N_1389,N_1412);
nor U1441 (N_1441,N_1413,N_1431);
xnor U1442 (N_1442,N_1395,N_1439);
nand U1443 (N_1443,N_1388,N_1390);
nand U1444 (N_1444,N_1429,N_1380);
nor U1445 (N_1445,N_1408,N_1419);
nand U1446 (N_1446,N_1384,N_1414);
nand U1447 (N_1447,N_1386,N_1434);
and U1448 (N_1448,N_1396,N_1432);
and U1449 (N_1449,N_1437,N_1430);
or U1450 (N_1450,N_1421,N_1410);
or U1451 (N_1451,N_1406,N_1405);
nor U1452 (N_1452,N_1397,N_1423);
nand U1453 (N_1453,N_1403,N_1426);
or U1454 (N_1454,N_1425,N_1407);
and U1455 (N_1455,N_1382,N_1438);
nand U1456 (N_1456,N_1433,N_1424);
and U1457 (N_1457,N_1381,N_1387);
nand U1458 (N_1458,N_1400,N_1420);
nor U1459 (N_1459,N_1402,N_1411);
or U1460 (N_1460,N_1428,N_1401);
nand U1461 (N_1461,N_1385,N_1418);
nand U1462 (N_1462,N_1436,N_1383);
or U1463 (N_1463,N_1422,N_1398);
and U1464 (N_1464,N_1394,N_1393);
or U1465 (N_1465,N_1435,N_1417);
nor U1466 (N_1466,N_1427,N_1416);
nor U1467 (N_1467,N_1404,N_1415);
and U1468 (N_1468,N_1391,N_1399);
nor U1469 (N_1469,N_1409,N_1392);
nor U1470 (N_1470,N_1435,N_1400);
nand U1471 (N_1471,N_1428,N_1396);
or U1472 (N_1472,N_1407,N_1423);
xnor U1473 (N_1473,N_1407,N_1411);
or U1474 (N_1474,N_1422,N_1433);
and U1475 (N_1475,N_1408,N_1404);
or U1476 (N_1476,N_1408,N_1391);
and U1477 (N_1477,N_1407,N_1394);
or U1478 (N_1478,N_1383,N_1432);
nand U1479 (N_1479,N_1392,N_1439);
and U1480 (N_1480,N_1402,N_1415);
nand U1481 (N_1481,N_1382,N_1415);
and U1482 (N_1482,N_1435,N_1431);
nand U1483 (N_1483,N_1395,N_1431);
nand U1484 (N_1484,N_1426,N_1424);
nand U1485 (N_1485,N_1434,N_1392);
nor U1486 (N_1486,N_1439,N_1428);
and U1487 (N_1487,N_1391,N_1385);
and U1488 (N_1488,N_1387,N_1434);
and U1489 (N_1489,N_1429,N_1423);
nand U1490 (N_1490,N_1433,N_1436);
and U1491 (N_1491,N_1422,N_1416);
nand U1492 (N_1492,N_1429,N_1424);
nor U1493 (N_1493,N_1437,N_1389);
and U1494 (N_1494,N_1389,N_1438);
and U1495 (N_1495,N_1420,N_1396);
and U1496 (N_1496,N_1397,N_1426);
and U1497 (N_1497,N_1428,N_1423);
nand U1498 (N_1498,N_1434,N_1423);
or U1499 (N_1499,N_1414,N_1395);
nand U1500 (N_1500,N_1478,N_1480);
and U1501 (N_1501,N_1448,N_1472);
nor U1502 (N_1502,N_1447,N_1444);
nand U1503 (N_1503,N_1471,N_1460);
or U1504 (N_1504,N_1459,N_1479);
nor U1505 (N_1505,N_1463,N_1491);
and U1506 (N_1506,N_1495,N_1464);
nor U1507 (N_1507,N_1476,N_1469);
nor U1508 (N_1508,N_1477,N_1490);
or U1509 (N_1509,N_1473,N_1466);
nand U1510 (N_1510,N_1456,N_1494);
and U1511 (N_1511,N_1441,N_1470);
or U1512 (N_1512,N_1485,N_1443);
nand U1513 (N_1513,N_1481,N_1453);
or U1514 (N_1514,N_1482,N_1461);
or U1515 (N_1515,N_1486,N_1468);
nand U1516 (N_1516,N_1488,N_1467);
or U1517 (N_1517,N_1458,N_1493);
and U1518 (N_1518,N_1487,N_1462);
nand U1519 (N_1519,N_1449,N_1483);
nor U1520 (N_1520,N_1452,N_1489);
and U1521 (N_1521,N_1455,N_1497);
nand U1522 (N_1522,N_1442,N_1499);
xnor U1523 (N_1523,N_1465,N_1445);
nor U1524 (N_1524,N_1474,N_1484);
and U1525 (N_1525,N_1440,N_1450);
nand U1526 (N_1526,N_1454,N_1457);
and U1527 (N_1527,N_1498,N_1475);
nand U1528 (N_1528,N_1492,N_1451);
or U1529 (N_1529,N_1446,N_1496);
nand U1530 (N_1530,N_1473,N_1456);
and U1531 (N_1531,N_1492,N_1486);
nand U1532 (N_1532,N_1475,N_1449);
or U1533 (N_1533,N_1480,N_1461);
nor U1534 (N_1534,N_1463,N_1499);
or U1535 (N_1535,N_1445,N_1466);
nand U1536 (N_1536,N_1455,N_1451);
and U1537 (N_1537,N_1474,N_1454);
nand U1538 (N_1538,N_1485,N_1481);
nor U1539 (N_1539,N_1471,N_1473);
nor U1540 (N_1540,N_1461,N_1465);
nor U1541 (N_1541,N_1466,N_1486);
nand U1542 (N_1542,N_1477,N_1487);
xnor U1543 (N_1543,N_1466,N_1487);
nand U1544 (N_1544,N_1440,N_1484);
nor U1545 (N_1545,N_1452,N_1459);
nor U1546 (N_1546,N_1471,N_1457);
nand U1547 (N_1547,N_1453,N_1466);
nand U1548 (N_1548,N_1442,N_1488);
and U1549 (N_1549,N_1472,N_1468);
and U1550 (N_1550,N_1491,N_1475);
nand U1551 (N_1551,N_1468,N_1491);
nand U1552 (N_1552,N_1440,N_1492);
nor U1553 (N_1553,N_1445,N_1485);
or U1554 (N_1554,N_1470,N_1462);
or U1555 (N_1555,N_1477,N_1454);
and U1556 (N_1556,N_1478,N_1454);
nand U1557 (N_1557,N_1462,N_1472);
and U1558 (N_1558,N_1465,N_1482);
and U1559 (N_1559,N_1474,N_1496);
nand U1560 (N_1560,N_1521,N_1551);
or U1561 (N_1561,N_1548,N_1528);
and U1562 (N_1562,N_1542,N_1547);
nor U1563 (N_1563,N_1518,N_1524);
nand U1564 (N_1564,N_1539,N_1534);
nor U1565 (N_1565,N_1501,N_1505);
nor U1566 (N_1566,N_1527,N_1517);
nand U1567 (N_1567,N_1559,N_1531);
or U1568 (N_1568,N_1510,N_1500);
nor U1569 (N_1569,N_1537,N_1503);
nor U1570 (N_1570,N_1502,N_1516);
nor U1571 (N_1571,N_1544,N_1532);
nor U1572 (N_1572,N_1536,N_1541);
or U1573 (N_1573,N_1526,N_1535);
nor U1574 (N_1574,N_1520,N_1558);
and U1575 (N_1575,N_1513,N_1543);
and U1576 (N_1576,N_1507,N_1538);
and U1577 (N_1577,N_1512,N_1508);
or U1578 (N_1578,N_1522,N_1550);
and U1579 (N_1579,N_1523,N_1552);
and U1580 (N_1580,N_1530,N_1554);
and U1581 (N_1581,N_1511,N_1514);
or U1582 (N_1582,N_1546,N_1556);
nand U1583 (N_1583,N_1529,N_1553);
nor U1584 (N_1584,N_1540,N_1504);
or U1585 (N_1585,N_1557,N_1525);
nand U1586 (N_1586,N_1519,N_1533);
and U1587 (N_1587,N_1549,N_1506);
and U1588 (N_1588,N_1545,N_1555);
and U1589 (N_1589,N_1509,N_1515);
nand U1590 (N_1590,N_1512,N_1514);
nor U1591 (N_1591,N_1506,N_1543);
or U1592 (N_1592,N_1545,N_1523);
xor U1593 (N_1593,N_1502,N_1547);
or U1594 (N_1594,N_1544,N_1528);
nor U1595 (N_1595,N_1549,N_1528);
and U1596 (N_1596,N_1504,N_1527);
nor U1597 (N_1597,N_1512,N_1520);
nand U1598 (N_1598,N_1524,N_1540);
or U1599 (N_1599,N_1531,N_1517);
and U1600 (N_1600,N_1538,N_1510);
or U1601 (N_1601,N_1556,N_1528);
nor U1602 (N_1602,N_1500,N_1541);
and U1603 (N_1603,N_1521,N_1511);
or U1604 (N_1604,N_1526,N_1543);
nor U1605 (N_1605,N_1523,N_1536);
nand U1606 (N_1606,N_1507,N_1533);
nand U1607 (N_1607,N_1513,N_1541);
nor U1608 (N_1608,N_1538,N_1525);
nand U1609 (N_1609,N_1529,N_1508);
or U1610 (N_1610,N_1552,N_1509);
or U1611 (N_1611,N_1509,N_1510);
nor U1612 (N_1612,N_1530,N_1503);
and U1613 (N_1613,N_1508,N_1546);
and U1614 (N_1614,N_1504,N_1519);
and U1615 (N_1615,N_1518,N_1540);
nand U1616 (N_1616,N_1548,N_1542);
and U1617 (N_1617,N_1553,N_1542);
and U1618 (N_1618,N_1537,N_1502);
nand U1619 (N_1619,N_1543,N_1556);
and U1620 (N_1620,N_1569,N_1608);
nor U1621 (N_1621,N_1586,N_1606);
nor U1622 (N_1622,N_1612,N_1596);
and U1623 (N_1623,N_1564,N_1618);
nor U1624 (N_1624,N_1619,N_1603);
and U1625 (N_1625,N_1589,N_1607);
or U1626 (N_1626,N_1571,N_1566);
and U1627 (N_1627,N_1575,N_1592);
nor U1628 (N_1628,N_1615,N_1578);
nand U1629 (N_1629,N_1576,N_1594);
or U1630 (N_1630,N_1609,N_1565);
nand U1631 (N_1631,N_1616,N_1563);
and U1632 (N_1632,N_1567,N_1568);
nand U1633 (N_1633,N_1604,N_1597);
nor U1634 (N_1634,N_1562,N_1572);
or U1635 (N_1635,N_1570,N_1573);
or U1636 (N_1636,N_1584,N_1613);
nand U1637 (N_1637,N_1611,N_1602);
or U1638 (N_1638,N_1614,N_1583);
or U1639 (N_1639,N_1605,N_1581);
xnor U1640 (N_1640,N_1585,N_1598);
nand U1641 (N_1641,N_1587,N_1591);
nor U1642 (N_1642,N_1582,N_1561);
or U1643 (N_1643,N_1580,N_1577);
nor U1644 (N_1644,N_1588,N_1574);
and U1645 (N_1645,N_1601,N_1560);
nor U1646 (N_1646,N_1593,N_1599);
nand U1647 (N_1647,N_1595,N_1590);
or U1648 (N_1648,N_1600,N_1610);
nor U1649 (N_1649,N_1617,N_1579);
nand U1650 (N_1650,N_1605,N_1607);
and U1651 (N_1651,N_1579,N_1613);
or U1652 (N_1652,N_1574,N_1607);
nor U1653 (N_1653,N_1601,N_1592);
or U1654 (N_1654,N_1604,N_1605);
nand U1655 (N_1655,N_1583,N_1564);
nor U1656 (N_1656,N_1617,N_1587);
nand U1657 (N_1657,N_1584,N_1561);
or U1658 (N_1658,N_1594,N_1589);
and U1659 (N_1659,N_1569,N_1572);
and U1660 (N_1660,N_1564,N_1589);
and U1661 (N_1661,N_1597,N_1590);
and U1662 (N_1662,N_1582,N_1594);
nor U1663 (N_1663,N_1563,N_1577);
and U1664 (N_1664,N_1578,N_1592);
and U1665 (N_1665,N_1593,N_1572);
nand U1666 (N_1666,N_1606,N_1585);
or U1667 (N_1667,N_1600,N_1581);
nor U1668 (N_1668,N_1580,N_1599);
or U1669 (N_1669,N_1608,N_1577);
nand U1670 (N_1670,N_1619,N_1583);
nor U1671 (N_1671,N_1575,N_1609);
or U1672 (N_1672,N_1573,N_1596);
nand U1673 (N_1673,N_1593,N_1586);
nor U1674 (N_1674,N_1573,N_1587);
and U1675 (N_1675,N_1574,N_1572);
or U1676 (N_1676,N_1571,N_1611);
and U1677 (N_1677,N_1578,N_1583);
nand U1678 (N_1678,N_1583,N_1601);
nand U1679 (N_1679,N_1577,N_1587);
nand U1680 (N_1680,N_1649,N_1656);
nor U1681 (N_1681,N_1675,N_1630);
nand U1682 (N_1682,N_1673,N_1662);
and U1683 (N_1683,N_1641,N_1626);
nand U1684 (N_1684,N_1647,N_1627);
nor U1685 (N_1685,N_1624,N_1661);
or U1686 (N_1686,N_1640,N_1650);
and U1687 (N_1687,N_1653,N_1671);
nand U1688 (N_1688,N_1637,N_1646);
or U1689 (N_1689,N_1625,N_1632);
or U1690 (N_1690,N_1629,N_1645);
nand U1691 (N_1691,N_1652,N_1677);
nor U1692 (N_1692,N_1678,N_1628);
or U1693 (N_1693,N_1672,N_1643);
nor U1694 (N_1694,N_1620,N_1679);
nand U1695 (N_1695,N_1667,N_1660);
or U1696 (N_1696,N_1659,N_1631);
nand U1697 (N_1697,N_1666,N_1638);
and U1698 (N_1698,N_1654,N_1648);
or U1699 (N_1699,N_1633,N_1664);
or U1700 (N_1700,N_1668,N_1621);
and U1701 (N_1701,N_1635,N_1663);
nand U1702 (N_1702,N_1676,N_1639);
nand U1703 (N_1703,N_1651,N_1642);
or U1704 (N_1704,N_1636,N_1669);
nor U1705 (N_1705,N_1634,N_1657);
nor U1706 (N_1706,N_1658,N_1665);
nand U1707 (N_1707,N_1622,N_1674);
and U1708 (N_1708,N_1670,N_1623);
nor U1709 (N_1709,N_1644,N_1655);
nor U1710 (N_1710,N_1638,N_1643);
or U1711 (N_1711,N_1629,N_1677);
nand U1712 (N_1712,N_1660,N_1638);
or U1713 (N_1713,N_1650,N_1674);
or U1714 (N_1714,N_1657,N_1633);
nor U1715 (N_1715,N_1624,N_1620);
nand U1716 (N_1716,N_1651,N_1647);
nand U1717 (N_1717,N_1656,N_1661);
nor U1718 (N_1718,N_1668,N_1673);
and U1719 (N_1719,N_1665,N_1652);
or U1720 (N_1720,N_1651,N_1672);
nor U1721 (N_1721,N_1660,N_1641);
or U1722 (N_1722,N_1679,N_1672);
nand U1723 (N_1723,N_1636,N_1647);
nand U1724 (N_1724,N_1667,N_1641);
nand U1725 (N_1725,N_1669,N_1646);
nor U1726 (N_1726,N_1637,N_1640);
nor U1727 (N_1727,N_1643,N_1665);
or U1728 (N_1728,N_1620,N_1641);
nor U1729 (N_1729,N_1655,N_1678);
nor U1730 (N_1730,N_1627,N_1650);
nor U1731 (N_1731,N_1642,N_1667);
nand U1732 (N_1732,N_1663,N_1660);
or U1733 (N_1733,N_1625,N_1638);
or U1734 (N_1734,N_1635,N_1665);
nor U1735 (N_1735,N_1653,N_1624);
or U1736 (N_1736,N_1659,N_1651);
and U1737 (N_1737,N_1629,N_1644);
nor U1738 (N_1738,N_1637,N_1662);
or U1739 (N_1739,N_1621,N_1677);
or U1740 (N_1740,N_1701,N_1706);
or U1741 (N_1741,N_1723,N_1682);
nand U1742 (N_1742,N_1693,N_1713);
and U1743 (N_1743,N_1695,N_1728);
nor U1744 (N_1744,N_1700,N_1685);
or U1745 (N_1745,N_1739,N_1686);
nor U1746 (N_1746,N_1691,N_1725);
nor U1747 (N_1747,N_1730,N_1689);
nor U1748 (N_1748,N_1736,N_1708);
or U1749 (N_1749,N_1735,N_1705);
nor U1750 (N_1750,N_1696,N_1698);
or U1751 (N_1751,N_1731,N_1710);
nor U1752 (N_1752,N_1738,N_1680);
nor U1753 (N_1753,N_1715,N_1720);
and U1754 (N_1754,N_1733,N_1714);
or U1755 (N_1755,N_1692,N_1694);
nor U1756 (N_1756,N_1712,N_1716);
and U1757 (N_1757,N_1702,N_1688);
nand U1758 (N_1758,N_1718,N_1721);
xnor U1759 (N_1759,N_1726,N_1699);
and U1760 (N_1760,N_1684,N_1681);
nor U1761 (N_1761,N_1737,N_1727);
nor U1762 (N_1762,N_1697,N_1687);
and U1763 (N_1763,N_1707,N_1734);
nor U1764 (N_1764,N_1709,N_1703);
nand U1765 (N_1765,N_1732,N_1717);
nor U1766 (N_1766,N_1711,N_1690);
or U1767 (N_1767,N_1704,N_1719);
nor U1768 (N_1768,N_1683,N_1729);
nand U1769 (N_1769,N_1724,N_1722);
nor U1770 (N_1770,N_1690,N_1724);
nand U1771 (N_1771,N_1702,N_1698);
and U1772 (N_1772,N_1718,N_1700);
and U1773 (N_1773,N_1722,N_1685);
nor U1774 (N_1774,N_1695,N_1722);
xor U1775 (N_1775,N_1711,N_1707);
nor U1776 (N_1776,N_1692,N_1729);
nand U1777 (N_1777,N_1718,N_1730);
nor U1778 (N_1778,N_1699,N_1690);
nand U1779 (N_1779,N_1709,N_1694);
or U1780 (N_1780,N_1699,N_1688);
and U1781 (N_1781,N_1729,N_1737);
or U1782 (N_1782,N_1694,N_1735);
nand U1783 (N_1783,N_1692,N_1739);
and U1784 (N_1784,N_1700,N_1727);
and U1785 (N_1785,N_1714,N_1694);
nor U1786 (N_1786,N_1697,N_1680);
nand U1787 (N_1787,N_1680,N_1715);
nand U1788 (N_1788,N_1707,N_1721);
or U1789 (N_1789,N_1683,N_1730);
nand U1790 (N_1790,N_1716,N_1727);
and U1791 (N_1791,N_1710,N_1686);
or U1792 (N_1792,N_1715,N_1698);
nor U1793 (N_1793,N_1706,N_1715);
nand U1794 (N_1794,N_1684,N_1701);
and U1795 (N_1795,N_1686,N_1713);
nor U1796 (N_1796,N_1686,N_1680);
and U1797 (N_1797,N_1698,N_1734);
and U1798 (N_1798,N_1704,N_1681);
nand U1799 (N_1799,N_1735,N_1689);
nor U1800 (N_1800,N_1776,N_1765);
or U1801 (N_1801,N_1774,N_1796);
nand U1802 (N_1802,N_1762,N_1793);
nor U1803 (N_1803,N_1757,N_1747);
nor U1804 (N_1804,N_1746,N_1761);
nor U1805 (N_1805,N_1783,N_1791);
or U1806 (N_1806,N_1792,N_1789);
nor U1807 (N_1807,N_1778,N_1798);
and U1808 (N_1808,N_1790,N_1740);
nor U1809 (N_1809,N_1743,N_1744);
and U1810 (N_1810,N_1781,N_1756);
and U1811 (N_1811,N_1753,N_1752);
and U1812 (N_1812,N_1794,N_1749);
or U1813 (N_1813,N_1773,N_1750);
nand U1814 (N_1814,N_1754,N_1787);
nor U1815 (N_1815,N_1766,N_1797);
nand U1816 (N_1816,N_1779,N_1777);
or U1817 (N_1817,N_1772,N_1784);
nor U1818 (N_1818,N_1755,N_1742);
nand U1819 (N_1819,N_1768,N_1760);
nor U1820 (N_1820,N_1786,N_1795);
and U1821 (N_1821,N_1758,N_1782);
and U1822 (N_1822,N_1788,N_1763);
and U1823 (N_1823,N_1751,N_1748);
nand U1824 (N_1824,N_1769,N_1745);
nor U1825 (N_1825,N_1775,N_1767);
nor U1826 (N_1826,N_1785,N_1771);
nand U1827 (N_1827,N_1741,N_1764);
nand U1828 (N_1828,N_1770,N_1780);
or U1829 (N_1829,N_1759,N_1799);
and U1830 (N_1830,N_1747,N_1753);
or U1831 (N_1831,N_1751,N_1799);
and U1832 (N_1832,N_1771,N_1794);
or U1833 (N_1833,N_1796,N_1743);
or U1834 (N_1834,N_1771,N_1758);
nand U1835 (N_1835,N_1746,N_1763);
nor U1836 (N_1836,N_1754,N_1781);
nand U1837 (N_1837,N_1793,N_1754);
or U1838 (N_1838,N_1772,N_1797);
nand U1839 (N_1839,N_1784,N_1747);
or U1840 (N_1840,N_1772,N_1769);
or U1841 (N_1841,N_1761,N_1779);
and U1842 (N_1842,N_1767,N_1742);
or U1843 (N_1843,N_1788,N_1789);
or U1844 (N_1844,N_1796,N_1741);
nor U1845 (N_1845,N_1745,N_1756);
nand U1846 (N_1846,N_1758,N_1773);
nor U1847 (N_1847,N_1761,N_1787);
and U1848 (N_1848,N_1748,N_1785);
nand U1849 (N_1849,N_1783,N_1751);
and U1850 (N_1850,N_1772,N_1777);
or U1851 (N_1851,N_1782,N_1788);
nor U1852 (N_1852,N_1758,N_1781);
nand U1853 (N_1853,N_1798,N_1797);
nor U1854 (N_1854,N_1756,N_1761);
and U1855 (N_1855,N_1799,N_1789);
and U1856 (N_1856,N_1781,N_1795);
or U1857 (N_1857,N_1778,N_1766);
and U1858 (N_1858,N_1747,N_1780);
nor U1859 (N_1859,N_1769,N_1777);
and U1860 (N_1860,N_1851,N_1805);
or U1861 (N_1861,N_1858,N_1840);
nor U1862 (N_1862,N_1857,N_1853);
or U1863 (N_1863,N_1847,N_1836);
and U1864 (N_1864,N_1821,N_1828);
nor U1865 (N_1865,N_1801,N_1823);
and U1866 (N_1866,N_1841,N_1845);
or U1867 (N_1867,N_1811,N_1849);
and U1868 (N_1868,N_1856,N_1803);
nor U1869 (N_1869,N_1855,N_1835);
and U1870 (N_1870,N_1819,N_1850);
and U1871 (N_1871,N_1815,N_1826);
or U1872 (N_1872,N_1800,N_1854);
nand U1873 (N_1873,N_1831,N_1852);
or U1874 (N_1874,N_1833,N_1813);
and U1875 (N_1875,N_1859,N_1844);
nor U1876 (N_1876,N_1808,N_1812);
nor U1877 (N_1877,N_1820,N_1829);
nand U1878 (N_1878,N_1816,N_1807);
nand U1879 (N_1879,N_1814,N_1842);
nor U1880 (N_1880,N_1846,N_1834);
or U1881 (N_1881,N_1822,N_1837);
or U1882 (N_1882,N_1832,N_1818);
nor U1883 (N_1883,N_1804,N_1809);
nor U1884 (N_1884,N_1802,N_1839);
nand U1885 (N_1885,N_1848,N_1810);
and U1886 (N_1886,N_1825,N_1817);
nor U1887 (N_1887,N_1843,N_1830);
nand U1888 (N_1888,N_1824,N_1827);
nor U1889 (N_1889,N_1838,N_1806);
or U1890 (N_1890,N_1840,N_1846);
or U1891 (N_1891,N_1813,N_1820);
nor U1892 (N_1892,N_1850,N_1847);
nand U1893 (N_1893,N_1837,N_1806);
or U1894 (N_1894,N_1806,N_1805);
nand U1895 (N_1895,N_1808,N_1817);
nand U1896 (N_1896,N_1815,N_1816);
and U1897 (N_1897,N_1828,N_1845);
nand U1898 (N_1898,N_1856,N_1830);
nand U1899 (N_1899,N_1837,N_1824);
or U1900 (N_1900,N_1845,N_1832);
nand U1901 (N_1901,N_1817,N_1815);
or U1902 (N_1902,N_1844,N_1846);
and U1903 (N_1903,N_1818,N_1842);
nand U1904 (N_1904,N_1835,N_1817);
and U1905 (N_1905,N_1800,N_1821);
nor U1906 (N_1906,N_1808,N_1825);
nor U1907 (N_1907,N_1828,N_1857);
nand U1908 (N_1908,N_1814,N_1800);
and U1909 (N_1909,N_1833,N_1828);
nand U1910 (N_1910,N_1801,N_1840);
or U1911 (N_1911,N_1836,N_1841);
or U1912 (N_1912,N_1803,N_1852);
nand U1913 (N_1913,N_1846,N_1808);
and U1914 (N_1914,N_1855,N_1821);
nand U1915 (N_1915,N_1847,N_1831);
or U1916 (N_1916,N_1826,N_1813);
and U1917 (N_1917,N_1832,N_1817);
or U1918 (N_1918,N_1810,N_1833);
nand U1919 (N_1919,N_1822,N_1838);
or U1920 (N_1920,N_1869,N_1894);
nand U1921 (N_1921,N_1883,N_1905);
or U1922 (N_1922,N_1862,N_1898);
or U1923 (N_1923,N_1876,N_1885);
nand U1924 (N_1924,N_1875,N_1896);
and U1925 (N_1925,N_1899,N_1863);
or U1926 (N_1926,N_1892,N_1881);
and U1927 (N_1927,N_1916,N_1888);
nor U1928 (N_1928,N_1884,N_1914);
or U1929 (N_1929,N_1890,N_1893);
nor U1930 (N_1930,N_1860,N_1874);
nor U1931 (N_1931,N_1872,N_1906);
and U1932 (N_1932,N_1919,N_1868);
or U1933 (N_1933,N_1913,N_1917);
and U1934 (N_1934,N_1880,N_1871);
and U1935 (N_1935,N_1904,N_1861);
or U1936 (N_1936,N_1915,N_1897);
or U1937 (N_1937,N_1873,N_1908);
nor U1938 (N_1938,N_1887,N_1886);
nand U1939 (N_1939,N_1910,N_1864);
and U1940 (N_1940,N_1882,N_1903);
nand U1941 (N_1941,N_1918,N_1870);
nand U1942 (N_1942,N_1878,N_1909);
and U1943 (N_1943,N_1867,N_1889);
or U1944 (N_1944,N_1911,N_1900);
nand U1945 (N_1945,N_1879,N_1907);
and U1946 (N_1946,N_1901,N_1877);
nand U1947 (N_1947,N_1902,N_1891);
nand U1948 (N_1948,N_1895,N_1912);
nor U1949 (N_1949,N_1865,N_1866);
and U1950 (N_1950,N_1898,N_1876);
or U1951 (N_1951,N_1877,N_1887);
and U1952 (N_1952,N_1885,N_1901);
nand U1953 (N_1953,N_1862,N_1918);
nor U1954 (N_1954,N_1882,N_1918);
and U1955 (N_1955,N_1888,N_1860);
nor U1956 (N_1956,N_1916,N_1873);
or U1957 (N_1957,N_1862,N_1866);
nand U1958 (N_1958,N_1898,N_1890);
or U1959 (N_1959,N_1873,N_1876);
or U1960 (N_1960,N_1907,N_1866);
nor U1961 (N_1961,N_1868,N_1900);
nand U1962 (N_1962,N_1898,N_1893);
nand U1963 (N_1963,N_1878,N_1896);
nand U1964 (N_1964,N_1900,N_1912);
or U1965 (N_1965,N_1870,N_1903);
or U1966 (N_1966,N_1908,N_1888);
nor U1967 (N_1967,N_1917,N_1877);
nand U1968 (N_1968,N_1916,N_1871);
or U1969 (N_1969,N_1898,N_1878);
nand U1970 (N_1970,N_1896,N_1886);
nor U1971 (N_1971,N_1891,N_1910);
nand U1972 (N_1972,N_1880,N_1883);
nor U1973 (N_1973,N_1871,N_1868);
and U1974 (N_1974,N_1874,N_1911);
or U1975 (N_1975,N_1887,N_1882);
or U1976 (N_1976,N_1866,N_1885);
or U1977 (N_1977,N_1909,N_1915);
nand U1978 (N_1978,N_1917,N_1874);
or U1979 (N_1979,N_1884,N_1874);
nand U1980 (N_1980,N_1956,N_1958);
nand U1981 (N_1981,N_1979,N_1961);
and U1982 (N_1982,N_1945,N_1921);
and U1983 (N_1983,N_1927,N_1960);
nor U1984 (N_1984,N_1976,N_1963);
or U1985 (N_1985,N_1970,N_1930);
or U1986 (N_1986,N_1966,N_1929);
nand U1987 (N_1987,N_1933,N_1935);
or U1988 (N_1988,N_1949,N_1941);
and U1989 (N_1989,N_1951,N_1962);
nor U1990 (N_1990,N_1923,N_1965);
and U1991 (N_1991,N_1971,N_1967);
and U1992 (N_1992,N_1924,N_1977);
and U1993 (N_1993,N_1946,N_1925);
and U1994 (N_1994,N_1937,N_1953);
nand U1995 (N_1995,N_1934,N_1959);
or U1996 (N_1996,N_1938,N_1974);
nand U1997 (N_1997,N_1931,N_1932);
and U1998 (N_1998,N_1939,N_1942);
nor U1999 (N_1999,N_1947,N_1964);
or U2000 (N_2000,N_1955,N_1928);
or U2001 (N_2001,N_1922,N_1950);
and U2002 (N_2002,N_1973,N_1944);
or U2003 (N_2003,N_1957,N_1968);
nand U2004 (N_2004,N_1936,N_1948);
and U2005 (N_2005,N_1972,N_1943);
or U2006 (N_2006,N_1940,N_1952);
and U2007 (N_2007,N_1978,N_1969);
nor U2008 (N_2008,N_1920,N_1975);
nand U2009 (N_2009,N_1954,N_1926);
and U2010 (N_2010,N_1934,N_1938);
and U2011 (N_2011,N_1924,N_1931);
nor U2012 (N_2012,N_1957,N_1935);
nand U2013 (N_2013,N_1934,N_1966);
nor U2014 (N_2014,N_1949,N_1956);
and U2015 (N_2015,N_1925,N_1962);
and U2016 (N_2016,N_1952,N_1957);
xnor U2017 (N_2017,N_1953,N_1956);
nand U2018 (N_2018,N_1937,N_1928);
nor U2019 (N_2019,N_1958,N_1924);
or U2020 (N_2020,N_1922,N_1947);
and U2021 (N_2021,N_1975,N_1966);
or U2022 (N_2022,N_1973,N_1947);
and U2023 (N_2023,N_1943,N_1939);
and U2024 (N_2024,N_1945,N_1979);
nand U2025 (N_2025,N_1964,N_1936);
or U2026 (N_2026,N_1979,N_1952);
nand U2027 (N_2027,N_1936,N_1933);
or U2028 (N_2028,N_1939,N_1944);
or U2029 (N_2029,N_1971,N_1922);
and U2030 (N_2030,N_1941,N_1961);
nand U2031 (N_2031,N_1970,N_1931);
nand U2032 (N_2032,N_1966,N_1923);
nor U2033 (N_2033,N_1966,N_1933);
nor U2034 (N_2034,N_1979,N_1927);
or U2035 (N_2035,N_1950,N_1936);
nand U2036 (N_2036,N_1961,N_1932);
or U2037 (N_2037,N_1923,N_1979);
and U2038 (N_2038,N_1970,N_1945);
nor U2039 (N_2039,N_1972,N_1948);
and U2040 (N_2040,N_2008,N_2002);
nand U2041 (N_2041,N_2018,N_2009);
nor U2042 (N_2042,N_1983,N_2003);
and U2043 (N_2043,N_2039,N_2034);
and U2044 (N_2044,N_2010,N_1990);
nor U2045 (N_2045,N_2016,N_2012);
nor U2046 (N_2046,N_1997,N_1982);
nand U2047 (N_2047,N_2029,N_2017);
and U2048 (N_2048,N_2014,N_2001);
and U2049 (N_2049,N_1996,N_1989);
nor U2050 (N_2050,N_2022,N_2013);
or U2051 (N_2051,N_2020,N_2025);
or U2052 (N_2052,N_2023,N_2011);
or U2053 (N_2053,N_2032,N_2035);
or U2054 (N_2054,N_2005,N_1984);
xor U2055 (N_2055,N_2026,N_1987);
nand U2056 (N_2056,N_2021,N_2024);
nor U2057 (N_2057,N_1995,N_1988);
or U2058 (N_2058,N_2036,N_1998);
or U2059 (N_2059,N_2007,N_2027);
and U2060 (N_2060,N_2019,N_2015);
nor U2061 (N_2061,N_2038,N_2000);
and U2062 (N_2062,N_1985,N_2037);
or U2063 (N_2063,N_1986,N_2028);
nand U2064 (N_2064,N_1993,N_2031);
or U2065 (N_2065,N_1991,N_1981);
and U2066 (N_2066,N_1994,N_2030);
or U2067 (N_2067,N_2004,N_1980);
or U2068 (N_2068,N_1992,N_2033);
nor U2069 (N_2069,N_1999,N_2006);
nor U2070 (N_2070,N_2001,N_2006);
and U2071 (N_2071,N_1988,N_2030);
nand U2072 (N_2072,N_1995,N_2011);
nor U2073 (N_2073,N_2039,N_1988);
or U2074 (N_2074,N_2014,N_1984);
xnor U2075 (N_2075,N_1999,N_2037);
or U2076 (N_2076,N_2014,N_2007);
or U2077 (N_2077,N_2023,N_2001);
or U2078 (N_2078,N_1988,N_2019);
and U2079 (N_2079,N_2003,N_2000);
nor U2080 (N_2080,N_2036,N_1991);
nor U2081 (N_2081,N_2035,N_2029);
nand U2082 (N_2082,N_1981,N_2014);
and U2083 (N_2083,N_2033,N_2026);
and U2084 (N_2084,N_1980,N_2036);
nand U2085 (N_2085,N_2014,N_2027);
nand U2086 (N_2086,N_2025,N_2032);
nor U2087 (N_2087,N_2005,N_2022);
or U2088 (N_2088,N_2030,N_2016);
or U2089 (N_2089,N_2029,N_1997);
nor U2090 (N_2090,N_2022,N_2012);
nand U2091 (N_2091,N_2030,N_2026);
or U2092 (N_2092,N_2022,N_2011);
or U2093 (N_2093,N_2024,N_1993);
nand U2094 (N_2094,N_1980,N_2007);
or U2095 (N_2095,N_2003,N_1996);
nor U2096 (N_2096,N_1992,N_1987);
or U2097 (N_2097,N_1984,N_2023);
and U2098 (N_2098,N_1981,N_2033);
nor U2099 (N_2099,N_1996,N_1982);
or U2100 (N_2100,N_2095,N_2061);
nor U2101 (N_2101,N_2096,N_2097);
nand U2102 (N_2102,N_2072,N_2083);
nor U2103 (N_2103,N_2075,N_2040);
or U2104 (N_2104,N_2064,N_2065);
or U2105 (N_2105,N_2047,N_2069);
or U2106 (N_2106,N_2068,N_2048);
or U2107 (N_2107,N_2078,N_2081);
and U2108 (N_2108,N_2062,N_2077);
nand U2109 (N_2109,N_2080,N_2067);
and U2110 (N_2110,N_2043,N_2098);
or U2111 (N_2111,N_2073,N_2054);
nand U2112 (N_2112,N_2051,N_2050);
nor U2113 (N_2113,N_2042,N_2085);
nand U2114 (N_2114,N_2059,N_2049);
nand U2115 (N_2115,N_2082,N_2086);
nor U2116 (N_2116,N_2056,N_2041);
nor U2117 (N_2117,N_2052,N_2045);
or U2118 (N_2118,N_2063,N_2084);
or U2119 (N_2119,N_2044,N_2091);
nor U2120 (N_2120,N_2099,N_2079);
nor U2121 (N_2121,N_2053,N_2058);
and U2122 (N_2122,N_2066,N_2071);
and U2123 (N_2123,N_2076,N_2090);
nor U2124 (N_2124,N_2055,N_2092);
and U2125 (N_2125,N_2060,N_2088);
or U2126 (N_2126,N_2093,N_2087);
or U2127 (N_2127,N_2057,N_2046);
and U2128 (N_2128,N_2089,N_2074);
nand U2129 (N_2129,N_2070,N_2094);
or U2130 (N_2130,N_2080,N_2066);
nor U2131 (N_2131,N_2056,N_2071);
nand U2132 (N_2132,N_2089,N_2079);
and U2133 (N_2133,N_2081,N_2064);
nand U2134 (N_2134,N_2086,N_2073);
nand U2135 (N_2135,N_2044,N_2055);
nor U2136 (N_2136,N_2046,N_2092);
nand U2137 (N_2137,N_2081,N_2072);
or U2138 (N_2138,N_2060,N_2048);
and U2139 (N_2139,N_2041,N_2053);
or U2140 (N_2140,N_2047,N_2061);
nor U2141 (N_2141,N_2096,N_2047);
nand U2142 (N_2142,N_2078,N_2090);
and U2143 (N_2143,N_2089,N_2096);
or U2144 (N_2144,N_2081,N_2098);
and U2145 (N_2145,N_2041,N_2071);
or U2146 (N_2146,N_2042,N_2095);
nor U2147 (N_2147,N_2073,N_2088);
nand U2148 (N_2148,N_2058,N_2096);
nor U2149 (N_2149,N_2093,N_2081);
and U2150 (N_2150,N_2082,N_2091);
and U2151 (N_2151,N_2068,N_2097);
nand U2152 (N_2152,N_2092,N_2071);
nor U2153 (N_2153,N_2084,N_2062);
and U2154 (N_2154,N_2072,N_2069);
nor U2155 (N_2155,N_2097,N_2076);
nor U2156 (N_2156,N_2061,N_2040);
nor U2157 (N_2157,N_2070,N_2068);
or U2158 (N_2158,N_2046,N_2088);
or U2159 (N_2159,N_2043,N_2065);
nand U2160 (N_2160,N_2103,N_2143);
and U2161 (N_2161,N_2154,N_2131);
or U2162 (N_2162,N_2151,N_2117);
or U2163 (N_2163,N_2104,N_2156);
or U2164 (N_2164,N_2109,N_2128);
nor U2165 (N_2165,N_2150,N_2135);
and U2166 (N_2166,N_2148,N_2124);
or U2167 (N_2167,N_2113,N_2138);
nand U2168 (N_2168,N_2100,N_2111);
nand U2169 (N_2169,N_2105,N_2102);
nor U2170 (N_2170,N_2125,N_2116);
or U2171 (N_2171,N_2122,N_2140);
or U2172 (N_2172,N_2141,N_2123);
or U2173 (N_2173,N_2108,N_2121);
nand U2174 (N_2174,N_2142,N_2139);
or U2175 (N_2175,N_2133,N_2158);
and U2176 (N_2176,N_2107,N_2101);
nor U2177 (N_2177,N_2119,N_2136);
nor U2178 (N_2178,N_2144,N_2153);
nor U2179 (N_2179,N_2132,N_2157);
nand U2180 (N_2180,N_2149,N_2145);
nand U2181 (N_2181,N_2152,N_2110);
nand U2182 (N_2182,N_2115,N_2112);
or U2183 (N_2183,N_2129,N_2126);
and U2184 (N_2184,N_2106,N_2130);
nand U2185 (N_2185,N_2134,N_2120);
or U2186 (N_2186,N_2127,N_2118);
and U2187 (N_2187,N_2146,N_2114);
nand U2188 (N_2188,N_2137,N_2147);
nand U2189 (N_2189,N_2155,N_2159);
nand U2190 (N_2190,N_2120,N_2149);
nand U2191 (N_2191,N_2127,N_2110);
nor U2192 (N_2192,N_2113,N_2155);
and U2193 (N_2193,N_2149,N_2143);
and U2194 (N_2194,N_2136,N_2117);
or U2195 (N_2195,N_2108,N_2114);
and U2196 (N_2196,N_2144,N_2101);
nand U2197 (N_2197,N_2159,N_2138);
nand U2198 (N_2198,N_2157,N_2113);
or U2199 (N_2199,N_2136,N_2113);
xnor U2200 (N_2200,N_2143,N_2113);
nand U2201 (N_2201,N_2134,N_2121);
nand U2202 (N_2202,N_2113,N_2154);
nand U2203 (N_2203,N_2116,N_2142);
nor U2204 (N_2204,N_2136,N_2134);
and U2205 (N_2205,N_2126,N_2125);
nand U2206 (N_2206,N_2123,N_2109);
nand U2207 (N_2207,N_2152,N_2147);
and U2208 (N_2208,N_2115,N_2144);
and U2209 (N_2209,N_2156,N_2105);
nand U2210 (N_2210,N_2120,N_2141);
and U2211 (N_2211,N_2117,N_2142);
or U2212 (N_2212,N_2129,N_2108);
or U2213 (N_2213,N_2134,N_2128);
nor U2214 (N_2214,N_2159,N_2110);
or U2215 (N_2215,N_2153,N_2111);
xor U2216 (N_2216,N_2115,N_2125);
nand U2217 (N_2217,N_2139,N_2117);
nor U2218 (N_2218,N_2128,N_2152);
or U2219 (N_2219,N_2110,N_2108);
nor U2220 (N_2220,N_2183,N_2177);
nand U2221 (N_2221,N_2180,N_2192);
nand U2222 (N_2222,N_2169,N_2200);
nand U2223 (N_2223,N_2202,N_2187);
and U2224 (N_2224,N_2206,N_2210);
nand U2225 (N_2225,N_2191,N_2170);
and U2226 (N_2226,N_2209,N_2184);
nand U2227 (N_2227,N_2161,N_2219);
and U2228 (N_2228,N_2162,N_2207);
nand U2229 (N_2229,N_2176,N_2185);
nand U2230 (N_2230,N_2201,N_2168);
nor U2231 (N_2231,N_2205,N_2163);
nand U2232 (N_2232,N_2165,N_2218);
nand U2233 (N_2233,N_2193,N_2199);
or U2234 (N_2234,N_2160,N_2212);
and U2235 (N_2235,N_2211,N_2213);
and U2236 (N_2236,N_2178,N_2167);
nand U2237 (N_2237,N_2203,N_2194);
or U2238 (N_2238,N_2172,N_2208);
and U2239 (N_2239,N_2216,N_2195);
or U2240 (N_2240,N_2166,N_2217);
nor U2241 (N_2241,N_2214,N_2179);
or U2242 (N_2242,N_2215,N_2196);
and U2243 (N_2243,N_2173,N_2186);
xor U2244 (N_2244,N_2181,N_2197);
and U2245 (N_2245,N_2182,N_2190);
nor U2246 (N_2246,N_2174,N_2164);
and U2247 (N_2247,N_2175,N_2188);
nand U2248 (N_2248,N_2198,N_2204);
nand U2249 (N_2249,N_2171,N_2189);
or U2250 (N_2250,N_2209,N_2176);
and U2251 (N_2251,N_2189,N_2199);
and U2252 (N_2252,N_2201,N_2167);
nand U2253 (N_2253,N_2167,N_2183);
or U2254 (N_2254,N_2180,N_2196);
nor U2255 (N_2255,N_2196,N_2162);
and U2256 (N_2256,N_2194,N_2189);
or U2257 (N_2257,N_2161,N_2190);
or U2258 (N_2258,N_2167,N_2169);
nand U2259 (N_2259,N_2186,N_2219);
and U2260 (N_2260,N_2216,N_2197);
or U2261 (N_2261,N_2171,N_2188);
and U2262 (N_2262,N_2201,N_2216);
nand U2263 (N_2263,N_2198,N_2206);
or U2264 (N_2264,N_2208,N_2185);
nor U2265 (N_2265,N_2177,N_2201);
nand U2266 (N_2266,N_2183,N_2212);
or U2267 (N_2267,N_2196,N_2168);
nor U2268 (N_2268,N_2200,N_2175);
nand U2269 (N_2269,N_2189,N_2168);
or U2270 (N_2270,N_2202,N_2198);
nand U2271 (N_2271,N_2216,N_2217);
nor U2272 (N_2272,N_2188,N_2167);
and U2273 (N_2273,N_2168,N_2166);
nor U2274 (N_2274,N_2210,N_2219);
nand U2275 (N_2275,N_2192,N_2179);
or U2276 (N_2276,N_2179,N_2211);
and U2277 (N_2277,N_2188,N_2207);
and U2278 (N_2278,N_2206,N_2185);
nor U2279 (N_2279,N_2209,N_2198);
nor U2280 (N_2280,N_2234,N_2233);
nand U2281 (N_2281,N_2275,N_2277);
nand U2282 (N_2282,N_2231,N_2269);
or U2283 (N_2283,N_2245,N_2248);
and U2284 (N_2284,N_2278,N_2273);
and U2285 (N_2285,N_2247,N_2223);
and U2286 (N_2286,N_2226,N_2240);
or U2287 (N_2287,N_2242,N_2246);
nand U2288 (N_2288,N_2261,N_2237);
nand U2289 (N_2289,N_2252,N_2249);
nand U2290 (N_2290,N_2239,N_2224);
and U2291 (N_2291,N_2236,N_2257);
and U2292 (N_2292,N_2279,N_2265);
nand U2293 (N_2293,N_2229,N_2258);
nor U2294 (N_2294,N_2274,N_2222);
and U2295 (N_2295,N_2271,N_2263);
nand U2296 (N_2296,N_2250,N_2228);
nor U2297 (N_2297,N_2244,N_2238);
xor U2298 (N_2298,N_2260,N_2251);
and U2299 (N_2299,N_2235,N_2262);
nand U2300 (N_2300,N_2221,N_2227);
nand U2301 (N_2301,N_2259,N_2270);
and U2302 (N_2302,N_2256,N_2268);
or U2303 (N_2303,N_2230,N_2225);
nor U2304 (N_2304,N_2276,N_2243);
nand U2305 (N_2305,N_2220,N_2255);
nor U2306 (N_2306,N_2272,N_2266);
or U2307 (N_2307,N_2267,N_2264);
nor U2308 (N_2308,N_2232,N_2253);
and U2309 (N_2309,N_2241,N_2254);
nor U2310 (N_2310,N_2255,N_2259);
and U2311 (N_2311,N_2276,N_2260);
xor U2312 (N_2312,N_2236,N_2234);
or U2313 (N_2313,N_2245,N_2258);
nor U2314 (N_2314,N_2232,N_2279);
and U2315 (N_2315,N_2223,N_2241);
or U2316 (N_2316,N_2241,N_2263);
xor U2317 (N_2317,N_2234,N_2267);
or U2318 (N_2318,N_2256,N_2278);
and U2319 (N_2319,N_2273,N_2267);
xor U2320 (N_2320,N_2272,N_2231);
nor U2321 (N_2321,N_2252,N_2266);
nor U2322 (N_2322,N_2267,N_2236);
and U2323 (N_2323,N_2244,N_2227);
nor U2324 (N_2324,N_2231,N_2260);
nand U2325 (N_2325,N_2256,N_2232);
nor U2326 (N_2326,N_2231,N_2271);
and U2327 (N_2327,N_2274,N_2272);
and U2328 (N_2328,N_2226,N_2277);
and U2329 (N_2329,N_2222,N_2252);
and U2330 (N_2330,N_2231,N_2257);
and U2331 (N_2331,N_2222,N_2271);
nor U2332 (N_2332,N_2273,N_2249);
and U2333 (N_2333,N_2264,N_2254);
and U2334 (N_2334,N_2245,N_2227);
or U2335 (N_2335,N_2264,N_2237);
nand U2336 (N_2336,N_2224,N_2227);
nor U2337 (N_2337,N_2242,N_2261);
and U2338 (N_2338,N_2225,N_2259);
nor U2339 (N_2339,N_2263,N_2273);
or U2340 (N_2340,N_2281,N_2311);
or U2341 (N_2341,N_2339,N_2316);
nor U2342 (N_2342,N_2329,N_2317);
nand U2343 (N_2343,N_2287,N_2321);
xor U2344 (N_2344,N_2332,N_2323);
or U2345 (N_2345,N_2327,N_2325);
nand U2346 (N_2346,N_2290,N_2333);
nand U2347 (N_2347,N_2320,N_2283);
or U2348 (N_2348,N_2330,N_2319);
nand U2349 (N_2349,N_2338,N_2324);
or U2350 (N_2350,N_2310,N_2299);
nor U2351 (N_2351,N_2280,N_2282);
or U2352 (N_2352,N_2308,N_2336);
nor U2353 (N_2353,N_2289,N_2295);
and U2354 (N_2354,N_2296,N_2326);
and U2355 (N_2355,N_2288,N_2335);
and U2356 (N_2356,N_2293,N_2309);
or U2357 (N_2357,N_2306,N_2337);
nor U2358 (N_2358,N_2304,N_2300);
nand U2359 (N_2359,N_2322,N_2331);
nor U2360 (N_2360,N_2303,N_2302);
nor U2361 (N_2361,N_2328,N_2298);
nor U2362 (N_2362,N_2297,N_2285);
or U2363 (N_2363,N_2334,N_2286);
nand U2364 (N_2364,N_2312,N_2314);
nand U2365 (N_2365,N_2301,N_2315);
nand U2366 (N_2366,N_2294,N_2318);
or U2367 (N_2367,N_2307,N_2291);
and U2368 (N_2368,N_2305,N_2284);
and U2369 (N_2369,N_2313,N_2292);
or U2370 (N_2370,N_2325,N_2306);
nand U2371 (N_2371,N_2319,N_2300);
and U2372 (N_2372,N_2302,N_2312);
and U2373 (N_2373,N_2317,N_2321);
nand U2374 (N_2374,N_2292,N_2309);
nand U2375 (N_2375,N_2300,N_2285);
and U2376 (N_2376,N_2284,N_2337);
or U2377 (N_2377,N_2308,N_2295);
xnor U2378 (N_2378,N_2324,N_2284);
nand U2379 (N_2379,N_2281,N_2308);
nand U2380 (N_2380,N_2306,N_2295);
nor U2381 (N_2381,N_2282,N_2306);
and U2382 (N_2382,N_2328,N_2322);
or U2383 (N_2383,N_2333,N_2338);
and U2384 (N_2384,N_2315,N_2330);
nor U2385 (N_2385,N_2308,N_2328);
or U2386 (N_2386,N_2305,N_2335);
nor U2387 (N_2387,N_2335,N_2326);
or U2388 (N_2388,N_2339,N_2294);
xnor U2389 (N_2389,N_2293,N_2332);
and U2390 (N_2390,N_2308,N_2303);
nor U2391 (N_2391,N_2330,N_2295);
nand U2392 (N_2392,N_2311,N_2338);
and U2393 (N_2393,N_2288,N_2332);
nor U2394 (N_2394,N_2307,N_2293);
nand U2395 (N_2395,N_2311,N_2303);
and U2396 (N_2396,N_2295,N_2291);
nor U2397 (N_2397,N_2289,N_2322);
nor U2398 (N_2398,N_2319,N_2329);
and U2399 (N_2399,N_2336,N_2298);
nand U2400 (N_2400,N_2383,N_2342);
and U2401 (N_2401,N_2393,N_2348);
and U2402 (N_2402,N_2340,N_2385);
and U2403 (N_2403,N_2362,N_2379);
and U2404 (N_2404,N_2352,N_2344);
nand U2405 (N_2405,N_2349,N_2341);
or U2406 (N_2406,N_2359,N_2372);
and U2407 (N_2407,N_2397,N_2384);
and U2408 (N_2408,N_2343,N_2370);
or U2409 (N_2409,N_2368,N_2363);
and U2410 (N_2410,N_2371,N_2369);
or U2411 (N_2411,N_2396,N_2376);
and U2412 (N_2412,N_2354,N_2391);
and U2413 (N_2413,N_2357,N_2386);
nor U2414 (N_2414,N_2398,N_2378);
and U2415 (N_2415,N_2367,N_2350);
nor U2416 (N_2416,N_2346,N_2380);
and U2417 (N_2417,N_2345,N_2377);
nor U2418 (N_2418,N_2353,N_2382);
or U2419 (N_2419,N_2360,N_2389);
and U2420 (N_2420,N_2373,N_2355);
and U2421 (N_2421,N_2390,N_2388);
nor U2422 (N_2422,N_2381,N_2394);
nand U2423 (N_2423,N_2347,N_2358);
nor U2424 (N_2424,N_2364,N_2351);
or U2425 (N_2425,N_2392,N_2395);
or U2426 (N_2426,N_2356,N_2366);
nor U2427 (N_2427,N_2387,N_2374);
or U2428 (N_2428,N_2399,N_2375);
nor U2429 (N_2429,N_2361,N_2365);
or U2430 (N_2430,N_2391,N_2382);
nor U2431 (N_2431,N_2393,N_2389);
and U2432 (N_2432,N_2370,N_2367);
nor U2433 (N_2433,N_2350,N_2353);
nand U2434 (N_2434,N_2349,N_2378);
and U2435 (N_2435,N_2360,N_2354);
nor U2436 (N_2436,N_2366,N_2354);
nand U2437 (N_2437,N_2390,N_2364);
nor U2438 (N_2438,N_2389,N_2354);
and U2439 (N_2439,N_2341,N_2345);
or U2440 (N_2440,N_2376,N_2362);
or U2441 (N_2441,N_2367,N_2354);
nor U2442 (N_2442,N_2383,N_2366);
or U2443 (N_2443,N_2346,N_2370);
nor U2444 (N_2444,N_2380,N_2364);
and U2445 (N_2445,N_2383,N_2345);
nor U2446 (N_2446,N_2389,N_2366);
nand U2447 (N_2447,N_2385,N_2387);
nand U2448 (N_2448,N_2383,N_2373);
and U2449 (N_2449,N_2363,N_2351);
and U2450 (N_2450,N_2378,N_2355);
nor U2451 (N_2451,N_2363,N_2354);
nor U2452 (N_2452,N_2357,N_2381);
nor U2453 (N_2453,N_2364,N_2385);
and U2454 (N_2454,N_2385,N_2362);
nand U2455 (N_2455,N_2384,N_2385);
nor U2456 (N_2456,N_2368,N_2349);
and U2457 (N_2457,N_2366,N_2380);
nor U2458 (N_2458,N_2367,N_2347);
nand U2459 (N_2459,N_2384,N_2383);
and U2460 (N_2460,N_2440,N_2424);
and U2461 (N_2461,N_2409,N_2439);
or U2462 (N_2462,N_2449,N_2432);
nand U2463 (N_2463,N_2457,N_2408);
and U2464 (N_2464,N_2407,N_2401);
or U2465 (N_2465,N_2448,N_2442);
xnor U2466 (N_2466,N_2412,N_2435);
and U2467 (N_2467,N_2433,N_2400);
or U2468 (N_2468,N_2431,N_2418);
and U2469 (N_2469,N_2417,N_2429);
nand U2470 (N_2470,N_2450,N_2416);
and U2471 (N_2471,N_2427,N_2410);
and U2472 (N_2472,N_2406,N_2455);
and U2473 (N_2473,N_2452,N_2423);
nor U2474 (N_2474,N_2414,N_2420);
nor U2475 (N_2475,N_2443,N_2438);
nor U2476 (N_2476,N_2458,N_2451);
nor U2477 (N_2477,N_2403,N_2436);
and U2478 (N_2478,N_2428,N_2402);
or U2479 (N_2479,N_2447,N_2453);
nand U2480 (N_2480,N_2434,N_2413);
nand U2481 (N_2481,N_2419,N_2415);
and U2482 (N_2482,N_2441,N_2445);
nand U2483 (N_2483,N_2454,N_2444);
nor U2484 (N_2484,N_2411,N_2437);
or U2485 (N_2485,N_2404,N_2456);
or U2486 (N_2486,N_2426,N_2446);
nor U2487 (N_2487,N_2422,N_2421);
or U2488 (N_2488,N_2459,N_2430);
and U2489 (N_2489,N_2425,N_2405);
and U2490 (N_2490,N_2401,N_2449);
nand U2491 (N_2491,N_2410,N_2455);
or U2492 (N_2492,N_2425,N_2424);
nor U2493 (N_2493,N_2450,N_2404);
and U2494 (N_2494,N_2401,N_2404);
nand U2495 (N_2495,N_2442,N_2429);
nand U2496 (N_2496,N_2425,N_2437);
or U2497 (N_2497,N_2441,N_2417);
nand U2498 (N_2498,N_2452,N_2407);
or U2499 (N_2499,N_2431,N_2438);
and U2500 (N_2500,N_2414,N_2402);
or U2501 (N_2501,N_2452,N_2455);
or U2502 (N_2502,N_2425,N_2433);
or U2503 (N_2503,N_2439,N_2457);
or U2504 (N_2504,N_2438,N_2400);
and U2505 (N_2505,N_2428,N_2447);
and U2506 (N_2506,N_2414,N_2412);
and U2507 (N_2507,N_2444,N_2421);
or U2508 (N_2508,N_2456,N_2444);
nand U2509 (N_2509,N_2443,N_2410);
or U2510 (N_2510,N_2425,N_2430);
nand U2511 (N_2511,N_2445,N_2452);
nor U2512 (N_2512,N_2432,N_2405);
and U2513 (N_2513,N_2413,N_2442);
xor U2514 (N_2514,N_2438,N_2425);
nor U2515 (N_2515,N_2415,N_2412);
or U2516 (N_2516,N_2449,N_2411);
and U2517 (N_2517,N_2446,N_2442);
nor U2518 (N_2518,N_2441,N_2402);
or U2519 (N_2519,N_2406,N_2435);
nor U2520 (N_2520,N_2462,N_2470);
nand U2521 (N_2521,N_2516,N_2496);
and U2522 (N_2522,N_2463,N_2482);
nor U2523 (N_2523,N_2494,N_2477);
nand U2524 (N_2524,N_2502,N_2484);
nand U2525 (N_2525,N_2472,N_2478);
nand U2526 (N_2526,N_2513,N_2508);
nor U2527 (N_2527,N_2510,N_2518);
and U2528 (N_2528,N_2467,N_2498);
or U2529 (N_2529,N_2506,N_2479);
nor U2530 (N_2530,N_2490,N_2514);
or U2531 (N_2531,N_2509,N_2493);
nor U2532 (N_2532,N_2476,N_2512);
nand U2533 (N_2533,N_2480,N_2471);
nor U2534 (N_2534,N_2517,N_2503);
nand U2535 (N_2535,N_2507,N_2489);
and U2536 (N_2536,N_2492,N_2515);
nor U2537 (N_2537,N_2466,N_2488);
nand U2538 (N_2538,N_2461,N_2469);
or U2539 (N_2539,N_2491,N_2505);
nor U2540 (N_2540,N_2468,N_2486);
and U2541 (N_2541,N_2465,N_2499);
or U2542 (N_2542,N_2500,N_2483);
or U2543 (N_2543,N_2495,N_2474);
nand U2544 (N_2544,N_2487,N_2501);
nand U2545 (N_2545,N_2519,N_2475);
nand U2546 (N_2546,N_2504,N_2511);
nor U2547 (N_2547,N_2473,N_2481);
xnor U2548 (N_2548,N_2464,N_2497);
nor U2549 (N_2549,N_2485,N_2460);
nor U2550 (N_2550,N_2481,N_2488);
and U2551 (N_2551,N_2497,N_2474);
and U2552 (N_2552,N_2467,N_2513);
nor U2553 (N_2553,N_2483,N_2511);
nand U2554 (N_2554,N_2469,N_2472);
nor U2555 (N_2555,N_2519,N_2476);
nand U2556 (N_2556,N_2468,N_2516);
and U2557 (N_2557,N_2465,N_2497);
nor U2558 (N_2558,N_2475,N_2481);
and U2559 (N_2559,N_2467,N_2469);
or U2560 (N_2560,N_2511,N_2486);
nor U2561 (N_2561,N_2506,N_2499);
or U2562 (N_2562,N_2479,N_2490);
and U2563 (N_2563,N_2474,N_2466);
and U2564 (N_2564,N_2476,N_2514);
and U2565 (N_2565,N_2479,N_2470);
nand U2566 (N_2566,N_2511,N_2509);
nor U2567 (N_2567,N_2510,N_2514);
nand U2568 (N_2568,N_2491,N_2495);
or U2569 (N_2569,N_2487,N_2469);
nor U2570 (N_2570,N_2507,N_2509);
nand U2571 (N_2571,N_2487,N_2515);
nor U2572 (N_2572,N_2506,N_2518);
and U2573 (N_2573,N_2471,N_2499);
or U2574 (N_2574,N_2488,N_2515);
nor U2575 (N_2575,N_2499,N_2492);
and U2576 (N_2576,N_2468,N_2461);
nor U2577 (N_2577,N_2501,N_2509);
nand U2578 (N_2578,N_2494,N_2509);
and U2579 (N_2579,N_2495,N_2509);
and U2580 (N_2580,N_2545,N_2567);
nand U2581 (N_2581,N_2522,N_2579);
and U2582 (N_2582,N_2530,N_2546);
or U2583 (N_2583,N_2529,N_2544);
and U2584 (N_2584,N_2563,N_2578);
nand U2585 (N_2585,N_2568,N_2561);
or U2586 (N_2586,N_2538,N_2573);
or U2587 (N_2587,N_2575,N_2521);
nand U2588 (N_2588,N_2559,N_2553);
or U2589 (N_2589,N_2569,N_2534);
and U2590 (N_2590,N_2539,N_2532);
nor U2591 (N_2591,N_2535,N_2551);
nand U2592 (N_2592,N_2574,N_2571);
nor U2593 (N_2593,N_2555,N_2531);
nor U2594 (N_2594,N_2577,N_2524);
nand U2595 (N_2595,N_2564,N_2552);
xnor U2596 (N_2596,N_2533,N_2547);
or U2597 (N_2597,N_2527,N_2557);
and U2598 (N_2598,N_2548,N_2562);
and U2599 (N_2599,N_2520,N_2558);
and U2600 (N_2600,N_2549,N_2526);
and U2601 (N_2601,N_2528,N_2572);
and U2602 (N_2602,N_2556,N_2537);
and U2603 (N_2603,N_2566,N_2576);
nor U2604 (N_2604,N_2523,N_2565);
or U2605 (N_2605,N_2540,N_2541);
nor U2606 (N_2606,N_2542,N_2536);
or U2607 (N_2607,N_2525,N_2554);
or U2608 (N_2608,N_2550,N_2543);
or U2609 (N_2609,N_2560,N_2570);
nand U2610 (N_2610,N_2537,N_2524);
nand U2611 (N_2611,N_2531,N_2562);
or U2612 (N_2612,N_2558,N_2577);
nor U2613 (N_2613,N_2565,N_2558);
and U2614 (N_2614,N_2521,N_2527);
nor U2615 (N_2615,N_2552,N_2540);
and U2616 (N_2616,N_2579,N_2558);
and U2617 (N_2617,N_2520,N_2577);
or U2618 (N_2618,N_2540,N_2565);
xor U2619 (N_2619,N_2561,N_2555);
and U2620 (N_2620,N_2551,N_2538);
nand U2621 (N_2621,N_2540,N_2564);
and U2622 (N_2622,N_2526,N_2540);
and U2623 (N_2623,N_2533,N_2568);
or U2624 (N_2624,N_2554,N_2574);
and U2625 (N_2625,N_2570,N_2544);
and U2626 (N_2626,N_2552,N_2551);
nand U2627 (N_2627,N_2525,N_2537);
and U2628 (N_2628,N_2522,N_2563);
nor U2629 (N_2629,N_2550,N_2563);
or U2630 (N_2630,N_2561,N_2527);
nor U2631 (N_2631,N_2570,N_2520);
nor U2632 (N_2632,N_2550,N_2570);
and U2633 (N_2633,N_2576,N_2521);
nand U2634 (N_2634,N_2530,N_2578);
nand U2635 (N_2635,N_2526,N_2544);
nand U2636 (N_2636,N_2524,N_2571);
nand U2637 (N_2637,N_2533,N_2539);
or U2638 (N_2638,N_2542,N_2568);
nand U2639 (N_2639,N_2541,N_2547);
nor U2640 (N_2640,N_2622,N_2612);
nor U2641 (N_2641,N_2611,N_2625);
nand U2642 (N_2642,N_2633,N_2620);
nor U2643 (N_2643,N_2606,N_2592);
and U2644 (N_2644,N_2610,N_2638);
or U2645 (N_2645,N_2607,N_2580);
or U2646 (N_2646,N_2632,N_2636);
nand U2647 (N_2647,N_2583,N_2624);
or U2648 (N_2648,N_2615,N_2596);
nand U2649 (N_2649,N_2605,N_2608);
nand U2650 (N_2650,N_2629,N_2600);
nand U2651 (N_2651,N_2617,N_2614);
nand U2652 (N_2652,N_2590,N_2637);
nor U2653 (N_2653,N_2623,N_2616);
nor U2654 (N_2654,N_2603,N_2588);
and U2655 (N_2655,N_2582,N_2593);
and U2656 (N_2656,N_2609,N_2621);
nand U2657 (N_2657,N_2628,N_2604);
nand U2658 (N_2658,N_2619,N_2601);
nand U2659 (N_2659,N_2626,N_2587);
nand U2660 (N_2660,N_2635,N_2630);
and U2661 (N_2661,N_2584,N_2585);
nor U2662 (N_2662,N_2597,N_2589);
nor U2663 (N_2663,N_2599,N_2595);
nor U2664 (N_2664,N_2602,N_2594);
nor U2665 (N_2665,N_2618,N_2639);
and U2666 (N_2666,N_2634,N_2613);
nor U2667 (N_2667,N_2591,N_2586);
or U2668 (N_2668,N_2631,N_2598);
nor U2669 (N_2669,N_2627,N_2581);
and U2670 (N_2670,N_2597,N_2583);
or U2671 (N_2671,N_2638,N_2618);
or U2672 (N_2672,N_2593,N_2621);
nand U2673 (N_2673,N_2604,N_2601);
and U2674 (N_2674,N_2610,N_2639);
nor U2675 (N_2675,N_2606,N_2595);
nor U2676 (N_2676,N_2582,N_2639);
and U2677 (N_2677,N_2605,N_2634);
nor U2678 (N_2678,N_2598,N_2626);
nor U2679 (N_2679,N_2624,N_2611);
xor U2680 (N_2680,N_2624,N_2587);
nor U2681 (N_2681,N_2613,N_2615);
or U2682 (N_2682,N_2593,N_2591);
and U2683 (N_2683,N_2580,N_2625);
nor U2684 (N_2684,N_2622,N_2602);
and U2685 (N_2685,N_2624,N_2598);
or U2686 (N_2686,N_2623,N_2639);
nor U2687 (N_2687,N_2613,N_2581);
nor U2688 (N_2688,N_2597,N_2603);
nand U2689 (N_2689,N_2589,N_2594);
nor U2690 (N_2690,N_2599,N_2592);
or U2691 (N_2691,N_2596,N_2621);
nor U2692 (N_2692,N_2617,N_2599);
or U2693 (N_2693,N_2593,N_2631);
nand U2694 (N_2694,N_2621,N_2601);
or U2695 (N_2695,N_2638,N_2580);
nand U2696 (N_2696,N_2602,N_2600);
nand U2697 (N_2697,N_2592,N_2614);
nor U2698 (N_2698,N_2633,N_2612);
nor U2699 (N_2699,N_2584,N_2616);
nor U2700 (N_2700,N_2673,N_2664);
nand U2701 (N_2701,N_2678,N_2680);
nor U2702 (N_2702,N_2655,N_2658);
and U2703 (N_2703,N_2679,N_2657);
nor U2704 (N_2704,N_2696,N_2651);
and U2705 (N_2705,N_2654,N_2669);
nand U2706 (N_2706,N_2670,N_2662);
and U2707 (N_2707,N_2697,N_2684);
or U2708 (N_2708,N_2681,N_2649);
and U2709 (N_2709,N_2686,N_2667);
and U2710 (N_2710,N_2693,N_2661);
and U2711 (N_2711,N_2688,N_2675);
and U2712 (N_2712,N_2640,N_2671);
nand U2713 (N_2713,N_2695,N_2653);
and U2714 (N_2714,N_2644,N_2652);
nand U2715 (N_2715,N_2646,N_2682);
nand U2716 (N_2716,N_2694,N_2699);
nor U2717 (N_2717,N_2647,N_2642);
and U2718 (N_2718,N_2687,N_2663);
nor U2719 (N_2719,N_2643,N_2668);
or U2720 (N_2720,N_2641,N_2659);
or U2721 (N_2721,N_2698,N_2692);
nor U2722 (N_2722,N_2689,N_2665);
and U2723 (N_2723,N_2677,N_2685);
nand U2724 (N_2724,N_2666,N_2656);
or U2725 (N_2725,N_2674,N_2672);
nand U2726 (N_2726,N_2648,N_2676);
xor U2727 (N_2727,N_2645,N_2650);
and U2728 (N_2728,N_2690,N_2683);
nor U2729 (N_2729,N_2691,N_2660);
nor U2730 (N_2730,N_2654,N_2698);
or U2731 (N_2731,N_2689,N_2640);
nor U2732 (N_2732,N_2672,N_2661);
or U2733 (N_2733,N_2647,N_2650);
or U2734 (N_2734,N_2652,N_2678);
or U2735 (N_2735,N_2667,N_2680);
and U2736 (N_2736,N_2684,N_2672);
and U2737 (N_2737,N_2653,N_2640);
nor U2738 (N_2738,N_2693,N_2665);
or U2739 (N_2739,N_2686,N_2688);
nand U2740 (N_2740,N_2691,N_2647);
and U2741 (N_2741,N_2677,N_2684);
nand U2742 (N_2742,N_2676,N_2677);
and U2743 (N_2743,N_2680,N_2692);
nor U2744 (N_2744,N_2677,N_2657);
nand U2745 (N_2745,N_2672,N_2657);
nand U2746 (N_2746,N_2674,N_2687);
nand U2747 (N_2747,N_2699,N_2684);
nand U2748 (N_2748,N_2655,N_2698);
nand U2749 (N_2749,N_2665,N_2688);
and U2750 (N_2750,N_2642,N_2669);
nor U2751 (N_2751,N_2655,N_2682);
nor U2752 (N_2752,N_2656,N_2685);
and U2753 (N_2753,N_2675,N_2655);
nor U2754 (N_2754,N_2686,N_2640);
nor U2755 (N_2755,N_2665,N_2676);
nand U2756 (N_2756,N_2648,N_2653);
or U2757 (N_2757,N_2659,N_2694);
and U2758 (N_2758,N_2674,N_2651);
and U2759 (N_2759,N_2691,N_2651);
nor U2760 (N_2760,N_2758,N_2713);
or U2761 (N_2761,N_2700,N_2740);
or U2762 (N_2762,N_2722,N_2732);
nand U2763 (N_2763,N_2731,N_2752);
or U2764 (N_2764,N_2719,N_2702);
and U2765 (N_2765,N_2756,N_2705);
and U2766 (N_2766,N_2707,N_2746);
and U2767 (N_2767,N_2735,N_2708);
nor U2768 (N_2768,N_2714,N_2716);
nand U2769 (N_2769,N_2753,N_2717);
and U2770 (N_2770,N_2754,N_2750);
or U2771 (N_2771,N_2739,N_2741);
nand U2772 (N_2772,N_2725,N_2744);
nand U2773 (N_2773,N_2738,N_2743);
nor U2774 (N_2774,N_2701,N_2742);
or U2775 (N_2775,N_2726,N_2755);
nand U2776 (N_2776,N_2721,N_2723);
nor U2777 (N_2777,N_2747,N_2737);
or U2778 (N_2778,N_2720,N_2711);
nor U2779 (N_2779,N_2724,N_2712);
or U2780 (N_2780,N_2745,N_2757);
or U2781 (N_2781,N_2751,N_2748);
xnor U2782 (N_2782,N_2733,N_2718);
nand U2783 (N_2783,N_2709,N_2728);
and U2784 (N_2784,N_2727,N_2730);
nand U2785 (N_2785,N_2759,N_2736);
nor U2786 (N_2786,N_2706,N_2710);
nand U2787 (N_2787,N_2749,N_2734);
or U2788 (N_2788,N_2729,N_2703);
and U2789 (N_2789,N_2704,N_2715);
and U2790 (N_2790,N_2714,N_2740);
nand U2791 (N_2791,N_2755,N_2753);
or U2792 (N_2792,N_2732,N_2703);
nand U2793 (N_2793,N_2704,N_2753);
nor U2794 (N_2794,N_2751,N_2708);
and U2795 (N_2795,N_2703,N_2742);
or U2796 (N_2796,N_2707,N_2724);
or U2797 (N_2797,N_2705,N_2747);
or U2798 (N_2798,N_2735,N_2730);
and U2799 (N_2799,N_2729,N_2706);
nor U2800 (N_2800,N_2755,N_2725);
or U2801 (N_2801,N_2759,N_2702);
nor U2802 (N_2802,N_2733,N_2703);
and U2803 (N_2803,N_2721,N_2754);
nand U2804 (N_2804,N_2734,N_2756);
and U2805 (N_2805,N_2702,N_2736);
and U2806 (N_2806,N_2726,N_2721);
nor U2807 (N_2807,N_2719,N_2729);
and U2808 (N_2808,N_2739,N_2718);
and U2809 (N_2809,N_2745,N_2714);
and U2810 (N_2810,N_2724,N_2736);
nand U2811 (N_2811,N_2716,N_2713);
and U2812 (N_2812,N_2742,N_2757);
nand U2813 (N_2813,N_2723,N_2704);
or U2814 (N_2814,N_2737,N_2723);
nand U2815 (N_2815,N_2725,N_2736);
and U2816 (N_2816,N_2736,N_2728);
or U2817 (N_2817,N_2712,N_2743);
nand U2818 (N_2818,N_2726,N_2750);
nand U2819 (N_2819,N_2721,N_2702);
nand U2820 (N_2820,N_2799,N_2793);
nor U2821 (N_2821,N_2779,N_2800);
or U2822 (N_2822,N_2814,N_2819);
nor U2823 (N_2823,N_2803,N_2797);
nor U2824 (N_2824,N_2762,N_2807);
nor U2825 (N_2825,N_2796,N_2783);
nor U2826 (N_2826,N_2795,N_2777);
and U2827 (N_2827,N_2761,N_2808);
nor U2828 (N_2828,N_2815,N_2792);
and U2829 (N_2829,N_2786,N_2813);
nor U2830 (N_2830,N_2809,N_2771);
or U2831 (N_2831,N_2767,N_2787);
nor U2832 (N_2832,N_2788,N_2818);
nand U2833 (N_2833,N_2765,N_2775);
nand U2834 (N_2834,N_2806,N_2778);
or U2835 (N_2835,N_2801,N_2781);
nand U2836 (N_2836,N_2805,N_2794);
nand U2837 (N_2837,N_2804,N_2773);
nor U2838 (N_2838,N_2816,N_2790);
or U2839 (N_2839,N_2812,N_2784);
or U2840 (N_2840,N_2764,N_2782);
nand U2841 (N_2841,N_2789,N_2802);
nor U2842 (N_2842,N_2769,N_2817);
or U2843 (N_2843,N_2811,N_2763);
nand U2844 (N_2844,N_2770,N_2780);
nand U2845 (N_2845,N_2774,N_2785);
nand U2846 (N_2846,N_2798,N_2760);
and U2847 (N_2847,N_2768,N_2776);
nor U2848 (N_2848,N_2810,N_2766);
and U2849 (N_2849,N_2772,N_2791);
and U2850 (N_2850,N_2815,N_2761);
or U2851 (N_2851,N_2769,N_2762);
and U2852 (N_2852,N_2771,N_2799);
nor U2853 (N_2853,N_2769,N_2819);
and U2854 (N_2854,N_2799,N_2814);
and U2855 (N_2855,N_2818,N_2761);
nor U2856 (N_2856,N_2818,N_2810);
nand U2857 (N_2857,N_2787,N_2788);
nand U2858 (N_2858,N_2815,N_2782);
nor U2859 (N_2859,N_2776,N_2810);
nor U2860 (N_2860,N_2791,N_2799);
and U2861 (N_2861,N_2778,N_2814);
or U2862 (N_2862,N_2818,N_2813);
or U2863 (N_2863,N_2769,N_2799);
nor U2864 (N_2864,N_2788,N_2797);
and U2865 (N_2865,N_2793,N_2818);
and U2866 (N_2866,N_2786,N_2788);
and U2867 (N_2867,N_2819,N_2796);
nand U2868 (N_2868,N_2784,N_2819);
nand U2869 (N_2869,N_2790,N_2812);
nand U2870 (N_2870,N_2810,N_2797);
and U2871 (N_2871,N_2790,N_2789);
or U2872 (N_2872,N_2815,N_2767);
or U2873 (N_2873,N_2781,N_2777);
nor U2874 (N_2874,N_2819,N_2790);
nor U2875 (N_2875,N_2800,N_2805);
or U2876 (N_2876,N_2768,N_2792);
nor U2877 (N_2877,N_2771,N_2803);
or U2878 (N_2878,N_2797,N_2765);
or U2879 (N_2879,N_2776,N_2795);
and U2880 (N_2880,N_2824,N_2872);
or U2881 (N_2881,N_2844,N_2842);
or U2882 (N_2882,N_2868,N_2826);
nand U2883 (N_2883,N_2867,N_2878);
and U2884 (N_2884,N_2827,N_2851);
or U2885 (N_2885,N_2846,N_2854);
nand U2886 (N_2886,N_2870,N_2835);
nand U2887 (N_2887,N_2833,N_2848);
nand U2888 (N_2888,N_2847,N_2820);
or U2889 (N_2889,N_2864,N_2861);
nand U2890 (N_2890,N_2830,N_2849);
or U2891 (N_2891,N_2850,N_2831);
nand U2892 (N_2892,N_2865,N_2856);
nand U2893 (N_2893,N_2859,N_2841);
and U2894 (N_2894,N_2838,N_2852);
and U2895 (N_2895,N_2839,N_2879);
or U2896 (N_2896,N_2825,N_2874);
xor U2897 (N_2897,N_2845,N_2860);
and U2898 (N_2898,N_2837,N_2828);
nand U2899 (N_2899,N_2858,N_2829);
and U2900 (N_2900,N_2832,N_2863);
or U2901 (N_2901,N_2866,N_2855);
or U2902 (N_2902,N_2840,N_2869);
and U2903 (N_2903,N_2836,N_2821);
or U2904 (N_2904,N_2871,N_2822);
nand U2905 (N_2905,N_2876,N_2877);
nor U2906 (N_2906,N_2857,N_2873);
or U2907 (N_2907,N_2843,N_2823);
or U2908 (N_2908,N_2834,N_2875);
nand U2909 (N_2909,N_2862,N_2853);
nand U2910 (N_2910,N_2855,N_2838);
nor U2911 (N_2911,N_2868,N_2836);
or U2912 (N_2912,N_2858,N_2845);
nor U2913 (N_2913,N_2826,N_2845);
nand U2914 (N_2914,N_2850,N_2846);
nand U2915 (N_2915,N_2853,N_2820);
and U2916 (N_2916,N_2844,N_2827);
nor U2917 (N_2917,N_2871,N_2836);
or U2918 (N_2918,N_2820,N_2874);
or U2919 (N_2919,N_2854,N_2847);
or U2920 (N_2920,N_2847,N_2834);
or U2921 (N_2921,N_2822,N_2845);
and U2922 (N_2922,N_2836,N_2840);
and U2923 (N_2923,N_2828,N_2861);
or U2924 (N_2924,N_2828,N_2847);
nor U2925 (N_2925,N_2834,N_2856);
and U2926 (N_2926,N_2847,N_2845);
nor U2927 (N_2927,N_2877,N_2824);
nand U2928 (N_2928,N_2879,N_2836);
nor U2929 (N_2929,N_2850,N_2837);
and U2930 (N_2930,N_2846,N_2860);
nor U2931 (N_2931,N_2857,N_2823);
nor U2932 (N_2932,N_2865,N_2852);
nor U2933 (N_2933,N_2846,N_2853);
nor U2934 (N_2934,N_2835,N_2869);
and U2935 (N_2935,N_2863,N_2853);
nor U2936 (N_2936,N_2833,N_2825);
nand U2937 (N_2937,N_2841,N_2867);
and U2938 (N_2938,N_2870,N_2837);
or U2939 (N_2939,N_2860,N_2825);
nand U2940 (N_2940,N_2906,N_2936);
or U2941 (N_2941,N_2929,N_2930);
and U2942 (N_2942,N_2883,N_2900);
and U2943 (N_2943,N_2914,N_2907);
nand U2944 (N_2944,N_2889,N_2933);
or U2945 (N_2945,N_2884,N_2928);
nand U2946 (N_2946,N_2922,N_2896);
nand U2947 (N_2947,N_2885,N_2912);
or U2948 (N_2948,N_2921,N_2939);
or U2949 (N_2949,N_2932,N_2938);
xor U2950 (N_2950,N_2908,N_2899);
nand U2951 (N_2951,N_2890,N_2935);
and U2952 (N_2952,N_2925,N_2927);
nor U2953 (N_2953,N_2919,N_2905);
nor U2954 (N_2954,N_2892,N_2913);
or U2955 (N_2955,N_2891,N_2909);
and U2956 (N_2956,N_2904,N_2934);
nand U2957 (N_2957,N_2893,N_2888);
and U2958 (N_2958,N_2916,N_2901);
nor U2959 (N_2959,N_2886,N_2882);
nor U2960 (N_2960,N_2895,N_2923);
nand U2961 (N_2961,N_2910,N_2915);
nand U2962 (N_2962,N_2917,N_2880);
nand U2963 (N_2963,N_2918,N_2926);
nor U2964 (N_2964,N_2924,N_2898);
nand U2965 (N_2965,N_2903,N_2902);
nand U2966 (N_2966,N_2911,N_2887);
nor U2967 (N_2967,N_2937,N_2897);
nand U2968 (N_2968,N_2920,N_2931);
and U2969 (N_2969,N_2881,N_2894);
and U2970 (N_2970,N_2886,N_2939);
nor U2971 (N_2971,N_2898,N_2932);
nand U2972 (N_2972,N_2916,N_2893);
nand U2973 (N_2973,N_2937,N_2911);
nor U2974 (N_2974,N_2923,N_2917);
nor U2975 (N_2975,N_2903,N_2880);
and U2976 (N_2976,N_2906,N_2886);
and U2977 (N_2977,N_2903,N_2932);
or U2978 (N_2978,N_2892,N_2905);
nor U2979 (N_2979,N_2906,N_2899);
nand U2980 (N_2980,N_2890,N_2914);
nor U2981 (N_2981,N_2920,N_2891);
or U2982 (N_2982,N_2927,N_2894);
nor U2983 (N_2983,N_2902,N_2926);
or U2984 (N_2984,N_2888,N_2887);
nand U2985 (N_2985,N_2883,N_2913);
and U2986 (N_2986,N_2909,N_2923);
or U2987 (N_2987,N_2891,N_2903);
or U2988 (N_2988,N_2909,N_2900);
and U2989 (N_2989,N_2921,N_2925);
nor U2990 (N_2990,N_2919,N_2937);
nand U2991 (N_2991,N_2905,N_2933);
nor U2992 (N_2992,N_2897,N_2922);
nor U2993 (N_2993,N_2928,N_2883);
or U2994 (N_2994,N_2884,N_2886);
nor U2995 (N_2995,N_2907,N_2881);
nand U2996 (N_2996,N_2916,N_2910);
nand U2997 (N_2997,N_2925,N_2926);
and U2998 (N_2998,N_2927,N_2881);
nand U2999 (N_2999,N_2939,N_2907);
or UO_0 (O_0,N_2960,N_2982);
or UO_1 (O_1,N_2957,N_2987);
and UO_2 (O_2,N_2964,N_2940);
or UO_3 (O_3,N_2945,N_2988);
nor UO_4 (O_4,N_2986,N_2998);
and UO_5 (O_5,N_2991,N_2954);
nor UO_6 (O_6,N_2949,N_2966);
nand UO_7 (O_7,N_2956,N_2971);
nand UO_8 (O_8,N_2952,N_2993);
or UO_9 (O_9,N_2996,N_2980);
nor UO_10 (O_10,N_2961,N_2942);
or UO_11 (O_11,N_2995,N_2990);
nand UO_12 (O_12,N_2997,N_2972);
nand UO_13 (O_13,N_2953,N_2999);
or UO_14 (O_14,N_2963,N_2970);
nand UO_15 (O_15,N_2974,N_2948);
or UO_16 (O_16,N_2944,N_2947);
nand UO_17 (O_17,N_2958,N_2946);
nor UO_18 (O_18,N_2994,N_2979);
nor UO_19 (O_19,N_2969,N_2981);
and UO_20 (O_20,N_2955,N_2975);
or UO_21 (O_21,N_2989,N_2950);
or UO_22 (O_22,N_2941,N_2973);
nor UO_23 (O_23,N_2983,N_2985);
nand UO_24 (O_24,N_2943,N_2976);
or UO_25 (O_25,N_2959,N_2951);
or UO_26 (O_26,N_2962,N_2977);
and UO_27 (O_27,N_2967,N_2965);
and UO_28 (O_28,N_2968,N_2992);
nor UO_29 (O_29,N_2978,N_2984);
nor UO_30 (O_30,N_2949,N_2977);
nand UO_31 (O_31,N_2961,N_2948);
nor UO_32 (O_32,N_2948,N_2986);
or UO_33 (O_33,N_2961,N_2969);
or UO_34 (O_34,N_2956,N_2978);
nor UO_35 (O_35,N_2983,N_2989);
or UO_36 (O_36,N_2998,N_2983);
or UO_37 (O_37,N_2998,N_2963);
and UO_38 (O_38,N_2982,N_2942);
nor UO_39 (O_39,N_2975,N_2967);
nand UO_40 (O_40,N_2978,N_2975);
nand UO_41 (O_41,N_2945,N_2977);
xnor UO_42 (O_42,N_2947,N_2982);
nor UO_43 (O_43,N_2942,N_2954);
and UO_44 (O_44,N_2988,N_2949);
nand UO_45 (O_45,N_2953,N_2950);
or UO_46 (O_46,N_2984,N_2948);
nand UO_47 (O_47,N_2962,N_2997);
or UO_48 (O_48,N_2965,N_2994);
and UO_49 (O_49,N_2959,N_2984);
nor UO_50 (O_50,N_2972,N_2971);
nor UO_51 (O_51,N_2949,N_2954);
nand UO_52 (O_52,N_2946,N_2966);
nand UO_53 (O_53,N_2948,N_2959);
and UO_54 (O_54,N_2975,N_2963);
nand UO_55 (O_55,N_2959,N_2998);
nand UO_56 (O_56,N_2946,N_2968);
nand UO_57 (O_57,N_2969,N_2953);
and UO_58 (O_58,N_2956,N_2972);
nand UO_59 (O_59,N_2958,N_2997);
and UO_60 (O_60,N_2963,N_2984);
nor UO_61 (O_61,N_2966,N_2955);
nor UO_62 (O_62,N_2965,N_2960);
or UO_63 (O_63,N_2986,N_2951);
and UO_64 (O_64,N_2965,N_2951);
or UO_65 (O_65,N_2953,N_2987);
nor UO_66 (O_66,N_2991,N_2955);
nand UO_67 (O_67,N_2987,N_2955);
nand UO_68 (O_68,N_2978,N_2971);
and UO_69 (O_69,N_2998,N_2956);
nand UO_70 (O_70,N_2940,N_2944);
and UO_71 (O_71,N_2992,N_2959);
nor UO_72 (O_72,N_2957,N_2942);
and UO_73 (O_73,N_2953,N_2983);
or UO_74 (O_74,N_2999,N_2951);
nor UO_75 (O_75,N_2967,N_2981);
and UO_76 (O_76,N_2957,N_2975);
or UO_77 (O_77,N_2998,N_2987);
and UO_78 (O_78,N_2940,N_2990);
nor UO_79 (O_79,N_2956,N_2986);
and UO_80 (O_80,N_2946,N_2988);
and UO_81 (O_81,N_2971,N_2998);
nor UO_82 (O_82,N_2953,N_2977);
nand UO_83 (O_83,N_2992,N_2961);
nor UO_84 (O_84,N_2974,N_2991);
nand UO_85 (O_85,N_2985,N_2940);
or UO_86 (O_86,N_2957,N_2959);
nor UO_87 (O_87,N_2979,N_2961);
and UO_88 (O_88,N_2968,N_2966);
nor UO_89 (O_89,N_2958,N_2973);
or UO_90 (O_90,N_2978,N_2992);
nor UO_91 (O_91,N_2946,N_2999);
nand UO_92 (O_92,N_2982,N_2979);
nor UO_93 (O_93,N_2943,N_2995);
nand UO_94 (O_94,N_2963,N_2961);
or UO_95 (O_95,N_2950,N_2969);
and UO_96 (O_96,N_2990,N_2963);
or UO_97 (O_97,N_2996,N_2983);
and UO_98 (O_98,N_2988,N_2954);
nand UO_99 (O_99,N_2982,N_2961);
xor UO_100 (O_100,N_2942,N_2964);
or UO_101 (O_101,N_2991,N_2978);
or UO_102 (O_102,N_2996,N_2997);
or UO_103 (O_103,N_2963,N_2958);
nand UO_104 (O_104,N_2967,N_2958);
nand UO_105 (O_105,N_2995,N_2962);
and UO_106 (O_106,N_2987,N_2994);
or UO_107 (O_107,N_2949,N_2943);
or UO_108 (O_108,N_2992,N_2947);
and UO_109 (O_109,N_2942,N_2987);
or UO_110 (O_110,N_2970,N_2955);
nor UO_111 (O_111,N_2952,N_2997);
or UO_112 (O_112,N_2941,N_2974);
nor UO_113 (O_113,N_2982,N_2949);
nor UO_114 (O_114,N_2956,N_2991);
or UO_115 (O_115,N_2944,N_2966);
or UO_116 (O_116,N_2991,N_2965);
nor UO_117 (O_117,N_2978,N_2979);
and UO_118 (O_118,N_2944,N_2973);
or UO_119 (O_119,N_2967,N_2995);
and UO_120 (O_120,N_2995,N_2988);
or UO_121 (O_121,N_2995,N_2985);
and UO_122 (O_122,N_2960,N_2942);
and UO_123 (O_123,N_2953,N_2965);
nand UO_124 (O_124,N_2942,N_2997);
and UO_125 (O_125,N_2977,N_2957);
or UO_126 (O_126,N_2945,N_2978);
and UO_127 (O_127,N_2948,N_2944);
and UO_128 (O_128,N_2954,N_2972);
and UO_129 (O_129,N_2992,N_2962);
nand UO_130 (O_130,N_2956,N_2969);
nor UO_131 (O_131,N_2963,N_2965);
nor UO_132 (O_132,N_2963,N_2979);
or UO_133 (O_133,N_2995,N_2966);
and UO_134 (O_134,N_2993,N_2979);
nor UO_135 (O_135,N_2951,N_2955);
and UO_136 (O_136,N_2969,N_2992);
and UO_137 (O_137,N_2950,N_2986);
and UO_138 (O_138,N_2995,N_2968);
or UO_139 (O_139,N_2961,N_2971);
nand UO_140 (O_140,N_2994,N_2960);
and UO_141 (O_141,N_2948,N_2985);
nand UO_142 (O_142,N_2982,N_2994);
nor UO_143 (O_143,N_2949,N_2942);
or UO_144 (O_144,N_2995,N_2972);
nor UO_145 (O_145,N_2967,N_2983);
nand UO_146 (O_146,N_2985,N_2979);
and UO_147 (O_147,N_2961,N_2943);
nand UO_148 (O_148,N_2960,N_2964);
and UO_149 (O_149,N_2991,N_2962);
and UO_150 (O_150,N_2963,N_2955);
nand UO_151 (O_151,N_2993,N_2989);
or UO_152 (O_152,N_2991,N_2992);
nor UO_153 (O_153,N_2990,N_2966);
nand UO_154 (O_154,N_2961,N_2967);
and UO_155 (O_155,N_2983,N_2961);
nor UO_156 (O_156,N_2970,N_2960);
and UO_157 (O_157,N_2945,N_2958);
nor UO_158 (O_158,N_2982,N_2963);
and UO_159 (O_159,N_2950,N_2946);
xnor UO_160 (O_160,N_2999,N_2970);
nand UO_161 (O_161,N_2948,N_2979);
nand UO_162 (O_162,N_2979,N_2940);
nand UO_163 (O_163,N_2990,N_2945);
and UO_164 (O_164,N_2948,N_2956);
nor UO_165 (O_165,N_2984,N_2954);
and UO_166 (O_166,N_2960,N_2983);
nand UO_167 (O_167,N_2958,N_2985);
nor UO_168 (O_168,N_2979,N_2991);
or UO_169 (O_169,N_2990,N_2997);
and UO_170 (O_170,N_2948,N_2942);
nand UO_171 (O_171,N_2990,N_2944);
nor UO_172 (O_172,N_2994,N_2973);
nand UO_173 (O_173,N_2954,N_2977);
nand UO_174 (O_174,N_2960,N_2969);
or UO_175 (O_175,N_2963,N_2964);
and UO_176 (O_176,N_2946,N_2953);
nor UO_177 (O_177,N_2999,N_2980);
nor UO_178 (O_178,N_2956,N_2988);
nor UO_179 (O_179,N_2983,N_2965);
nor UO_180 (O_180,N_2971,N_2999);
xor UO_181 (O_181,N_2993,N_2999);
nand UO_182 (O_182,N_2943,N_2975);
nor UO_183 (O_183,N_2967,N_2990);
or UO_184 (O_184,N_2969,N_2955);
nand UO_185 (O_185,N_2951,N_2987);
nand UO_186 (O_186,N_2964,N_2979);
nand UO_187 (O_187,N_2973,N_2978);
nor UO_188 (O_188,N_2987,N_2985);
nor UO_189 (O_189,N_2969,N_2991);
and UO_190 (O_190,N_2986,N_2963);
and UO_191 (O_191,N_2948,N_2962);
and UO_192 (O_192,N_2972,N_2949);
nor UO_193 (O_193,N_2979,N_2969);
and UO_194 (O_194,N_2997,N_2950);
and UO_195 (O_195,N_2962,N_2953);
nand UO_196 (O_196,N_2951,N_2994);
and UO_197 (O_197,N_2995,N_2984);
and UO_198 (O_198,N_2967,N_2996);
or UO_199 (O_199,N_2957,N_2992);
nand UO_200 (O_200,N_2949,N_2953);
nand UO_201 (O_201,N_2972,N_2945);
and UO_202 (O_202,N_2985,N_2956);
nor UO_203 (O_203,N_2974,N_2995);
or UO_204 (O_204,N_2985,N_2992);
nand UO_205 (O_205,N_2981,N_2956);
nand UO_206 (O_206,N_2973,N_2965);
and UO_207 (O_207,N_2966,N_2979);
nand UO_208 (O_208,N_2966,N_2976);
and UO_209 (O_209,N_2973,N_2987);
nand UO_210 (O_210,N_2992,N_2981);
nor UO_211 (O_211,N_2989,N_2960);
nand UO_212 (O_212,N_2987,N_2960);
nand UO_213 (O_213,N_2961,N_2968);
and UO_214 (O_214,N_2977,N_2959);
or UO_215 (O_215,N_2973,N_2977);
or UO_216 (O_216,N_2963,N_2988);
nand UO_217 (O_217,N_2965,N_2959);
or UO_218 (O_218,N_2999,N_2965);
nand UO_219 (O_219,N_2974,N_2945);
and UO_220 (O_220,N_2952,N_2968);
or UO_221 (O_221,N_2994,N_2972);
nand UO_222 (O_222,N_2970,N_2979);
or UO_223 (O_223,N_2991,N_2975);
and UO_224 (O_224,N_2955,N_2956);
nand UO_225 (O_225,N_2973,N_2948);
nor UO_226 (O_226,N_2988,N_2992);
and UO_227 (O_227,N_2994,N_2941);
or UO_228 (O_228,N_2940,N_2986);
or UO_229 (O_229,N_2988,N_2953);
and UO_230 (O_230,N_2956,N_2970);
or UO_231 (O_231,N_2980,N_2987);
or UO_232 (O_232,N_2974,N_2990);
nor UO_233 (O_233,N_2964,N_2987);
or UO_234 (O_234,N_2948,N_2969);
and UO_235 (O_235,N_2985,N_2976);
and UO_236 (O_236,N_2978,N_2954);
nand UO_237 (O_237,N_2958,N_2956);
and UO_238 (O_238,N_2951,N_2960);
nor UO_239 (O_239,N_2984,N_2957);
and UO_240 (O_240,N_2990,N_2985);
nor UO_241 (O_241,N_2980,N_2942);
or UO_242 (O_242,N_2986,N_2981);
or UO_243 (O_243,N_2968,N_2956);
nand UO_244 (O_244,N_2961,N_2990);
nor UO_245 (O_245,N_2997,N_2946);
nor UO_246 (O_246,N_2962,N_2957);
and UO_247 (O_247,N_2990,N_2954);
nand UO_248 (O_248,N_2943,N_2946);
nor UO_249 (O_249,N_2994,N_2991);
nor UO_250 (O_250,N_2953,N_2947);
or UO_251 (O_251,N_2954,N_2951);
nand UO_252 (O_252,N_2960,N_2958);
or UO_253 (O_253,N_2974,N_2992);
or UO_254 (O_254,N_2951,N_2973);
or UO_255 (O_255,N_2983,N_2946);
nor UO_256 (O_256,N_2973,N_2995);
and UO_257 (O_257,N_2974,N_2970);
nand UO_258 (O_258,N_2959,N_2971);
or UO_259 (O_259,N_2985,N_2993);
nor UO_260 (O_260,N_2973,N_2983);
or UO_261 (O_261,N_2966,N_2954);
or UO_262 (O_262,N_2988,N_2950);
nand UO_263 (O_263,N_2992,N_2948);
nand UO_264 (O_264,N_2971,N_2970);
and UO_265 (O_265,N_2974,N_2977);
xor UO_266 (O_266,N_2993,N_2994);
nand UO_267 (O_267,N_2946,N_2976);
nor UO_268 (O_268,N_2998,N_2992);
nand UO_269 (O_269,N_2955,N_2982);
nor UO_270 (O_270,N_2997,N_2992);
and UO_271 (O_271,N_2976,N_2963);
nor UO_272 (O_272,N_2967,N_2978);
nand UO_273 (O_273,N_2956,N_2983);
nand UO_274 (O_274,N_2989,N_2980);
and UO_275 (O_275,N_2990,N_2942);
nor UO_276 (O_276,N_2986,N_2962);
nor UO_277 (O_277,N_2989,N_2948);
and UO_278 (O_278,N_2955,N_2980);
nand UO_279 (O_279,N_2956,N_2944);
and UO_280 (O_280,N_2996,N_2945);
and UO_281 (O_281,N_2986,N_2985);
nor UO_282 (O_282,N_2948,N_2988);
or UO_283 (O_283,N_2985,N_2994);
nand UO_284 (O_284,N_2971,N_2991);
nor UO_285 (O_285,N_2976,N_2993);
nor UO_286 (O_286,N_2974,N_2976);
nand UO_287 (O_287,N_2956,N_2962);
nor UO_288 (O_288,N_2956,N_2940);
nand UO_289 (O_289,N_2962,N_2971);
and UO_290 (O_290,N_2985,N_2954);
nand UO_291 (O_291,N_2949,N_2984);
nand UO_292 (O_292,N_2948,N_2967);
or UO_293 (O_293,N_2949,N_2992);
or UO_294 (O_294,N_2981,N_2973);
or UO_295 (O_295,N_2949,N_2985);
or UO_296 (O_296,N_2956,N_2946);
nand UO_297 (O_297,N_2955,N_2950);
and UO_298 (O_298,N_2994,N_2995);
nand UO_299 (O_299,N_2987,N_2946);
or UO_300 (O_300,N_2960,N_2940);
nand UO_301 (O_301,N_2965,N_2968);
and UO_302 (O_302,N_2947,N_2995);
or UO_303 (O_303,N_2953,N_2985);
nor UO_304 (O_304,N_2971,N_2975);
and UO_305 (O_305,N_2941,N_2984);
nand UO_306 (O_306,N_2978,N_2976);
nand UO_307 (O_307,N_2998,N_2964);
nand UO_308 (O_308,N_2949,N_2980);
and UO_309 (O_309,N_2964,N_2994);
nand UO_310 (O_310,N_2989,N_2942);
or UO_311 (O_311,N_2975,N_2952);
or UO_312 (O_312,N_2993,N_2983);
xnor UO_313 (O_313,N_2996,N_2949);
nand UO_314 (O_314,N_2940,N_2966);
nand UO_315 (O_315,N_2959,N_2978);
nor UO_316 (O_316,N_2975,N_2997);
and UO_317 (O_317,N_2951,N_2991);
nand UO_318 (O_318,N_2990,N_2971);
and UO_319 (O_319,N_2958,N_2989);
or UO_320 (O_320,N_2994,N_2955);
or UO_321 (O_321,N_2975,N_2940);
nand UO_322 (O_322,N_2986,N_2978);
or UO_323 (O_323,N_2940,N_2965);
nand UO_324 (O_324,N_2985,N_2942);
nand UO_325 (O_325,N_2991,N_2970);
or UO_326 (O_326,N_2957,N_2971);
and UO_327 (O_327,N_2950,N_2974);
nor UO_328 (O_328,N_2962,N_2967);
nor UO_329 (O_329,N_2967,N_2982);
and UO_330 (O_330,N_2946,N_2977);
nand UO_331 (O_331,N_2977,N_2966);
nor UO_332 (O_332,N_2986,N_2987);
and UO_333 (O_333,N_2989,N_2992);
nand UO_334 (O_334,N_2958,N_2991);
and UO_335 (O_335,N_2998,N_2970);
nand UO_336 (O_336,N_2957,N_2966);
nand UO_337 (O_337,N_2950,N_2951);
nor UO_338 (O_338,N_2981,N_2944);
or UO_339 (O_339,N_2996,N_2944);
and UO_340 (O_340,N_2947,N_2981);
and UO_341 (O_341,N_2989,N_2978);
nor UO_342 (O_342,N_2967,N_2993);
nand UO_343 (O_343,N_2998,N_2990);
and UO_344 (O_344,N_2941,N_2987);
nor UO_345 (O_345,N_2959,N_2962);
or UO_346 (O_346,N_2966,N_2998);
nand UO_347 (O_347,N_2979,N_2942);
nor UO_348 (O_348,N_2996,N_2948);
nand UO_349 (O_349,N_2969,N_2999);
and UO_350 (O_350,N_2984,N_2947);
or UO_351 (O_351,N_2956,N_2976);
or UO_352 (O_352,N_2980,N_2979);
nor UO_353 (O_353,N_2984,N_2996);
and UO_354 (O_354,N_2984,N_2953);
and UO_355 (O_355,N_2965,N_2989);
or UO_356 (O_356,N_2973,N_2996);
and UO_357 (O_357,N_2941,N_2952);
and UO_358 (O_358,N_2958,N_2990);
or UO_359 (O_359,N_2971,N_2949);
and UO_360 (O_360,N_2970,N_2995);
and UO_361 (O_361,N_2970,N_2958);
or UO_362 (O_362,N_2956,N_2997);
or UO_363 (O_363,N_2940,N_2984);
or UO_364 (O_364,N_2989,N_2994);
nor UO_365 (O_365,N_2965,N_2978);
or UO_366 (O_366,N_2987,N_2991);
nor UO_367 (O_367,N_2950,N_2979);
and UO_368 (O_368,N_2971,N_2980);
nor UO_369 (O_369,N_2946,N_2998);
nor UO_370 (O_370,N_2957,N_2968);
nor UO_371 (O_371,N_2996,N_2993);
nor UO_372 (O_372,N_2975,N_2961);
nor UO_373 (O_373,N_2999,N_2998);
and UO_374 (O_374,N_2967,N_2970);
nand UO_375 (O_375,N_2975,N_2990);
nor UO_376 (O_376,N_2957,N_2979);
xor UO_377 (O_377,N_2998,N_2984);
nand UO_378 (O_378,N_2961,N_2960);
and UO_379 (O_379,N_2952,N_2996);
nor UO_380 (O_380,N_2975,N_2960);
or UO_381 (O_381,N_2944,N_2997);
nand UO_382 (O_382,N_2983,N_2963);
or UO_383 (O_383,N_2983,N_2984);
nand UO_384 (O_384,N_2970,N_2984);
or UO_385 (O_385,N_2999,N_2959);
nand UO_386 (O_386,N_2962,N_2940);
nand UO_387 (O_387,N_2995,N_2976);
nor UO_388 (O_388,N_2942,N_2965);
nand UO_389 (O_389,N_2980,N_2964);
nor UO_390 (O_390,N_2952,N_2998);
nor UO_391 (O_391,N_2947,N_2973);
nor UO_392 (O_392,N_2983,N_2949);
nand UO_393 (O_393,N_2968,N_2958);
nor UO_394 (O_394,N_2984,N_2958);
nor UO_395 (O_395,N_2955,N_2945);
nand UO_396 (O_396,N_2946,N_2991);
nand UO_397 (O_397,N_2940,N_2948);
nand UO_398 (O_398,N_2962,N_2964);
nand UO_399 (O_399,N_2949,N_2955);
nor UO_400 (O_400,N_2942,N_2955);
or UO_401 (O_401,N_2993,N_2968);
nor UO_402 (O_402,N_2947,N_2974);
or UO_403 (O_403,N_2960,N_2984);
and UO_404 (O_404,N_2988,N_2980);
nor UO_405 (O_405,N_2974,N_2957);
and UO_406 (O_406,N_2956,N_2951);
and UO_407 (O_407,N_2986,N_2972);
nand UO_408 (O_408,N_2993,N_2984);
or UO_409 (O_409,N_2992,N_2940);
or UO_410 (O_410,N_2990,N_2972);
nand UO_411 (O_411,N_2998,N_2972);
or UO_412 (O_412,N_2967,N_2949);
nor UO_413 (O_413,N_2986,N_2969);
nor UO_414 (O_414,N_2964,N_2999);
and UO_415 (O_415,N_2986,N_2942);
nor UO_416 (O_416,N_2971,N_2940);
nand UO_417 (O_417,N_2984,N_2980);
xnor UO_418 (O_418,N_2952,N_2949);
nand UO_419 (O_419,N_2958,N_2940);
and UO_420 (O_420,N_2940,N_2972);
and UO_421 (O_421,N_2968,N_2940);
nand UO_422 (O_422,N_2960,N_2952);
nand UO_423 (O_423,N_2951,N_2962);
nand UO_424 (O_424,N_2977,N_2981);
or UO_425 (O_425,N_2974,N_2952);
nor UO_426 (O_426,N_2981,N_2958);
and UO_427 (O_427,N_2990,N_2982);
nand UO_428 (O_428,N_2992,N_2941);
nand UO_429 (O_429,N_2948,N_2994);
nand UO_430 (O_430,N_2947,N_2957);
or UO_431 (O_431,N_2967,N_2940);
or UO_432 (O_432,N_2971,N_2983);
or UO_433 (O_433,N_2952,N_2988);
or UO_434 (O_434,N_2994,N_2997);
nor UO_435 (O_435,N_2962,N_2942);
xor UO_436 (O_436,N_2969,N_2995);
nor UO_437 (O_437,N_2957,N_2986);
nand UO_438 (O_438,N_2986,N_2982);
and UO_439 (O_439,N_2995,N_2993);
nor UO_440 (O_440,N_2941,N_2999);
and UO_441 (O_441,N_2954,N_2957);
or UO_442 (O_442,N_2967,N_2972);
nand UO_443 (O_443,N_2991,N_2980);
and UO_444 (O_444,N_2943,N_2998);
nor UO_445 (O_445,N_2968,N_2975);
or UO_446 (O_446,N_2951,N_2980);
nand UO_447 (O_447,N_2964,N_2954);
nor UO_448 (O_448,N_2968,N_2953);
or UO_449 (O_449,N_2979,N_2995);
nor UO_450 (O_450,N_2945,N_2946);
nor UO_451 (O_451,N_2976,N_2973);
and UO_452 (O_452,N_2985,N_2973);
and UO_453 (O_453,N_2943,N_2982);
or UO_454 (O_454,N_2970,N_2982);
nor UO_455 (O_455,N_2995,N_2954);
and UO_456 (O_456,N_2961,N_2954);
nor UO_457 (O_457,N_2991,N_2950);
and UO_458 (O_458,N_2998,N_2982);
and UO_459 (O_459,N_2977,N_2970);
and UO_460 (O_460,N_2989,N_2976);
nand UO_461 (O_461,N_2987,N_2974);
and UO_462 (O_462,N_2999,N_2967);
or UO_463 (O_463,N_2945,N_2941);
nor UO_464 (O_464,N_2969,N_2954);
or UO_465 (O_465,N_2986,N_2979);
nor UO_466 (O_466,N_2984,N_2987);
or UO_467 (O_467,N_2961,N_2981);
and UO_468 (O_468,N_2985,N_2957);
xor UO_469 (O_469,N_2964,N_2993);
nand UO_470 (O_470,N_2940,N_2947);
nand UO_471 (O_471,N_2975,N_2966);
and UO_472 (O_472,N_2965,N_2984);
nand UO_473 (O_473,N_2998,N_2969);
nor UO_474 (O_474,N_2975,N_2977);
or UO_475 (O_475,N_2988,N_2994);
xor UO_476 (O_476,N_2980,N_2966);
nand UO_477 (O_477,N_2965,N_2964);
and UO_478 (O_478,N_2982,N_2975);
xor UO_479 (O_479,N_2953,N_2998);
nand UO_480 (O_480,N_2980,N_2970);
or UO_481 (O_481,N_2978,N_2970);
and UO_482 (O_482,N_2968,N_2943);
or UO_483 (O_483,N_2952,N_2986);
nor UO_484 (O_484,N_2944,N_2959);
or UO_485 (O_485,N_2995,N_2956);
and UO_486 (O_486,N_2942,N_2951);
or UO_487 (O_487,N_2996,N_2977);
or UO_488 (O_488,N_2969,N_2957);
xnor UO_489 (O_489,N_2940,N_2977);
nor UO_490 (O_490,N_2943,N_2981);
nand UO_491 (O_491,N_2970,N_2981);
and UO_492 (O_492,N_2994,N_2980);
and UO_493 (O_493,N_2980,N_2972);
nor UO_494 (O_494,N_2995,N_2949);
nand UO_495 (O_495,N_2965,N_2987);
nor UO_496 (O_496,N_2980,N_2954);
or UO_497 (O_497,N_2957,N_2960);
nand UO_498 (O_498,N_2964,N_2943);
nand UO_499 (O_499,N_2997,N_2998);
endmodule