module basic_3000_30000_3500_30_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
xor U0 (N_0,In_2317,In_2096);
and U1 (N_1,In_2416,In_1479);
nand U2 (N_2,In_1851,In_1247);
nor U3 (N_3,In_61,In_552);
or U4 (N_4,In_1536,In_610);
and U5 (N_5,In_1015,In_2201);
or U6 (N_6,In_2490,In_884);
nand U7 (N_7,In_2629,In_2194);
nand U8 (N_8,In_476,In_1245);
or U9 (N_9,In_1850,In_1055);
or U10 (N_10,In_2315,In_238);
nor U11 (N_11,In_670,In_2918);
xor U12 (N_12,In_941,In_675);
nor U13 (N_13,In_2180,In_2961);
and U14 (N_14,In_876,In_25);
or U15 (N_15,In_472,In_1759);
and U16 (N_16,In_1209,In_548);
xnor U17 (N_17,In_2134,In_204);
nand U18 (N_18,In_2847,In_1868);
or U19 (N_19,In_1541,In_2343);
and U20 (N_20,In_2381,In_145);
or U21 (N_21,In_2541,In_8);
nor U22 (N_22,In_1783,In_1307);
xor U23 (N_23,In_1149,In_423);
xnor U24 (N_24,In_1235,In_668);
or U25 (N_25,In_579,In_939);
and U26 (N_26,In_1478,In_1776);
nand U27 (N_27,In_1,In_478);
or U28 (N_28,In_1809,In_509);
nor U29 (N_29,In_2928,In_177);
and U30 (N_30,In_350,In_2861);
nand U31 (N_31,In_1107,In_2648);
nand U32 (N_32,In_1582,In_2375);
xnor U33 (N_33,In_2692,In_1763);
or U34 (N_34,In_1983,In_953);
or U35 (N_35,In_1781,In_1442);
and U36 (N_36,In_2395,In_2810);
nor U37 (N_37,In_2011,In_754);
or U38 (N_38,In_2385,In_137);
and U39 (N_39,In_440,In_2752);
or U40 (N_40,In_2219,In_966);
nand U41 (N_41,In_1207,In_1921);
and U42 (N_42,In_530,In_1760);
or U43 (N_43,In_1404,In_919);
xor U44 (N_44,In_187,In_375);
xor U45 (N_45,In_1376,In_2045);
xnor U46 (N_46,In_1593,In_1237);
or U47 (N_47,In_349,In_2791);
nor U48 (N_48,In_604,In_1777);
or U49 (N_49,In_1772,In_2111);
xnor U50 (N_50,In_969,In_255);
and U51 (N_51,In_2034,In_2334);
or U52 (N_52,In_1801,In_1915);
and U53 (N_53,In_1356,In_230);
and U54 (N_54,In_1383,In_1256);
nor U55 (N_55,In_2402,In_2638);
or U56 (N_56,In_2026,In_1903);
and U57 (N_57,In_122,In_2710);
and U58 (N_58,In_457,In_1135);
nor U59 (N_59,In_748,In_2519);
or U60 (N_60,In_2420,In_381);
or U61 (N_61,In_2878,In_1949);
nor U62 (N_62,In_449,In_641);
and U63 (N_63,In_1026,In_1443);
nor U64 (N_64,In_1375,In_2732);
and U65 (N_65,In_625,In_1933);
xor U66 (N_66,In_44,In_2141);
xor U67 (N_67,In_411,In_424);
and U68 (N_68,In_2760,In_461);
nand U69 (N_69,In_2184,In_2972);
nor U70 (N_70,In_2244,In_1609);
xnor U71 (N_71,In_2192,In_1317);
xnor U72 (N_72,In_1714,In_1787);
nand U73 (N_73,In_2454,In_816);
nor U74 (N_74,In_1663,In_1615);
nand U75 (N_75,In_1412,In_1600);
and U76 (N_76,In_2537,In_791);
and U77 (N_77,In_2153,In_2340);
nand U78 (N_78,In_2666,In_1693);
or U79 (N_79,In_2683,In_2319);
or U80 (N_80,In_2390,In_609);
or U81 (N_81,In_1203,In_2126);
xnor U82 (N_82,In_1715,In_2550);
nand U83 (N_83,In_128,In_1489);
and U84 (N_84,In_2988,In_2772);
xnor U85 (N_85,In_1040,In_2964);
xnor U86 (N_86,In_1571,In_873);
and U87 (N_87,In_521,In_881);
and U88 (N_88,In_1870,In_157);
xor U89 (N_89,In_1409,In_1852);
and U90 (N_90,In_464,In_1349);
nor U91 (N_91,In_947,In_1445);
or U92 (N_92,In_2065,In_802);
nand U93 (N_93,In_1332,In_753);
xnor U94 (N_94,In_439,In_909);
or U95 (N_95,In_1434,In_860);
and U96 (N_96,In_1862,In_37);
nand U97 (N_97,In_404,In_2121);
nand U98 (N_98,In_1056,In_142);
xnor U99 (N_99,In_275,In_708);
nand U100 (N_100,In_713,In_1829);
or U101 (N_101,In_2608,In_1044);
nor U102 (N_102,In_729,In_2177);
nand U103 (N_103,In_2971,In_2151);
or U104 (N_104,In_2508,In_1914);
xnor U105 (N_105,In_907,In_2013);
or U106 (N_106,In_1539,In_1405);
nand U107 (N_107,In_429,In_2957);
nor U108 (N_108,In_2503,In_638);
xor U109 (N_109,In_1788,In_2884);
nand U110 (N_110,In_719,In_805);
nand U111 (N_111,In_896,In_815);
and U112 (N_112,In_2855,In_2076);
nor U113 (N_113,In_267,In_2584);
or U114 (N_114,In_655,In_1198);
nor U115 (N_115,In_2651,In_1296);
and U116 (N_116,In_2080,In_691);
xor U117 (N_117,In_2284,In_2359);
or U118 (N_118,In_1884,In_1795);
nand U119 (N_119,In_2149,In_2310);
nor U120 (N_120,In_2676,In_1608);
and U121 (N_121,In_812,In_563);
or U122 (N_122,In_2744,In_1395);
xor U123 (N_123,In_1290,In_1281);
and U124 (N_124,In_2902,In_1030);
and U125 (N_125,In_2798,In_367);
and U126 (N_126,In_2631,In_2101);
nand U127 (N_127,In_1299,In_2885);
nor U128 (N_128,In_1400,In_2804);
nand U129 (N_129,In_2784,In_1060);
and U130 (N_130,In_2759,In_2733);
and U131 (N_131,In_616,In_1746);
nor U132 (N_132,In_2057,In_1682);
and U133 (N_133,In_322,In_2906);
xnor U134 (N_134,In_402,In_810);
nor U135 (N_135,In_895,In_1729);
nor U136 (N_136,In_764,In_2127);
nor U137 (N_137,In_1258,In_2718);
or U138 (N_138,In_2768,In_2487);
or U139 (N_139,In_1537,In_2349);
xnor U140 (N_140,In_1849,In_1716);
nor U141 (N_141,In_555,In_2516);
nand U142 (N_142,In_2227,In_1988);
xor U143 (N_143,In_1461,In_2698);
nor U144 (N_144,In_2523,In_2697);
and U145 (N_145,In_692,In_2895);
and U146 (N_146,In_2448,In_244);
nor U147 (N_147,In_1354,In_1192);
and U148 (N_148,In_2886,In_1972);
or U149 (N_149,In_1213,In_2518);
nand U150 (N_150,In_649,In_2921);
and U151 (N_151,In_1554,In_2821);
and U152 (N_152,In_874,In_2967);
xor U153 (N_153,In_2348,In_498);
nor U154 (N_154,In_751,In_2112);
xor U155 (N_155,In_2642,In_1959);
and U156 (N_156,In_2331,In_57);
nor U157 (N_157,In_192,In_1200);
nand U158 (N_158,In_1004,In_2135);
nand U159 (N_159,In_600,In_2748);
and U160 (N_160,In_357,In_92);
xnor U161 (N_161,In_2216,In_2603);
nand U162 (N_162,In_2428,In_1257);
and U163 (N_163,In_1225,In_2394);
nand U164 (N_164,In_918,In_2222);
and U165 (N_165,In_1579,In_47);
nand U166 (N_166,In_1553,In_797);
xnor U167 (N_167,In_501,In_2577);
nand U168 (N_168,In_219,In_2368);
xor U169 (N_169,In_2538,In_1498);
and U170 (N_170,In_2463,In_1866);
nor U171 (N_171,In_1468,In_2363);
and U172 (N_172,In_1509,In_2499);
xor U173 (N_173,In_1009,In_2029);
nor U174 (N_174,In_294,In_1005);
nand U175 (N_175,In_2453,In_2412);
nor U176 (N_176,In_2293,In_793);
and U177 (N_177,In_2785,In_314);
nand U178 (N_178,In_510,In_2802);
or U179 (N_179,In_1337,In_262);
nand U180 (N_180,In_1587,In_952);
or U181 (N_181,In_27,In_2746);
or U182 (N_182,In_828,In_1758);
or U183 (N_183,In_1649,In_989);
or U184 (N_184,In_221,In_1270);
xnor U185 (N_185,In_782,In_2148);
and U186 (N_186,In_631,In_2636);
or U187 (N_187,In_174,In_2387);
or U188 (N_188,In_2292,In_2838);
and U189 (N_189,In_81,In_2280);
nand U190 (N_190,In_1062,In_596);
nor U191 (N_191,In_2346,In_743);
or U192 (N_192,In_716,In_777);
or U193 (N_193,In_1540,In_944);
and U194 (N_194,In_97,In_1646);
nand U195 (N_195,In_803,In_487);
and U196 (N_196,In_662,In_2751);
xor U197 (N_197,In_408,In_1335);
nand U198 (N_198,In_2484,In_2341);
xor U199 (N_199,In_2758,In_2393);
nor U200 (N_200,In_2517,In_1707);
nor U201 (N_201,In_1749,In_2823);
and U202 (N_202,In_1326,In_2370);
xor U203 (N_203,In_2500,In_454);
or U204 (N_204,In_2836,In_1944);
xnor U205 (N_205,In_1341,In_2413);
nand U206 (N_206,In_225,In_2747);
nor U207 (N_207,In_849,In_2702);
or U208 (N_208,In_2110,In_704);
xnor U209 (N_209,In_76,In_1698);
or U210 (N_210,In_1076,In_554);
nand U211 (N_211,In_1179,In_2031);
nor U212 (N_212,In_1033,In_1961);
nor U213 (N_213,In_2896,In_2994);
nor U214 (N_214,In_2862,In_181);
or U215 (N_215,In_223,In_2900);
or U216 (N_216,In_506,In_2806);
nor U217 (N_217,In_2047,In_861);
or U218 (N_218,In_2437,In_2399);
and U219 (N_219,In_2681,In_2777);
or U220 (N_220,In_2042,In_284);
and U221 (N_221,In_117,In_125);
and U222 (N_222,In_1289,In_1657);
or U223 (N_223,In_2833,In_292);
or U224 (N_224,In_2700,In_1043);
nand U225 (N_225,In_549,In_2980);
xnor U226 (N_226,In_804,In_2060);
xnor U227 (N_227,In_1229,In_1750);
or U228 (N_228,In_1941,In_879);
nor U229 (N_229,In_2593,In_1518);
nor U230 (N_230,In_1578,In_212);
xnor U231 (N_231,In_232,In_7);
nand U232 (N_232,In_1275,In_1967);
nand U233 (N_233,In_1742,In_285);
or U234 (N_234,In_976,In_1822);
xor U235 (N_235,In_734,In_528);
nand U236 (N_236,In_2471,In_1182);
nor U237 (N_237,In_1555,In_2946);
nand U238 (N_238,In_2087,In_848);
or U239 (N_239,In_1011,In_1981);
nand U240 (N_240,In_2050,In_1420);
and U241 (N_241,In_445,In_2941);
nand U242 (N_242,In_450,In_2513);
nand U243 (N_243,In_698,In_663);
and U244 (N_244,In_1806,In_2232);
and U245 (N_245,In_1073,In_1117);
xor U246 (N_246,In_826,In_1472);
or U247 (N_247,In_91,In_967);
and U248 (N_248,In_747,In_2701);
or U249 (N_249,In_2669,In_2212);
and U250 (N_250,In_1481,In_1877);
and U251 (N_251,In_1293,In_1007);
xnor U252 (N_252,In_2435,In_93);
nor U253 (N_253,In_2256,In_380);
xnor U254 (N_254,In_766,In_369);
xnor U255 (N_255,In_372,In_36);
and U256 (N_256,In_1067,In_1020);
and U257 (N_257,In_749,In_463);
nand U258 (N_258,In_234,In_795);
xnor U259 (N_259,In_1476,In_295);
and U260 (N_260,In_1132,In_899);
and U261 (N_261,In_1285,In_1956);
nand U262 (N_262,In_1090,In_1180);
nand U263 (N_263,In_739,In_2267);
or U264 (N_264,In_1912,In_2679);
xor U265 (N_265,In_695,In_1544);
xor U266 (N_266,In_2071,In_33);
and U267 (N_267,In_1310,In_200);
or U268 (N_268,In_1659,In_1993);
or U269 (N_269,In_1490,In_252);
nor U270 (N_270,In_26,In_2623);
or U271 (N_271,In_1145,In_1086);
nand U272 (N_272,In_1658,In_431);
and U273 (N_273,In_2734,In_1301);
or U274 (N_274,In_2796,In_2145);
nand U275 (N_275,In_176,In_1099);
xnor U276 (N_276,In_2671,In_948);
nand U277 (N_277,In_1466,In_1899);
nor U278 (N_278,In_446,In_2574);
or U279 (N_279,In_2816,In_2270);
nand U280 (N_280,In_980,In_540);
nand U281 (N_281,In_283,In_388);
and U282 (N_282,In_2466,In_2940);
nor U283 (N_283,In_2044,In_762);
and U284 (N_284,In_792,In_512);
xor U285 (N_285,In_1928,In_1268);
xnor U286 (N_286,In_1423,In_256);
or U287 (N_287,In_260,In_1484);
or U288 (N_288,In_316,In_2417);
and U289 (N_289,In_1745,In_1391);
and U290 (N_290,In_687,In_877);
or U291 (N_291,In_2067,In_1083);
xor U292 (N_292,In_1584,In_193);
or U293 (N_293,In_1504,In_1599);
or U294 (N_294,In_1163,In_1230);
nand U295 (N_295,In_1415,In_2820);
nor U296 (N_296,In_48,In_1176);
xnor U297 (N_297,In_2093,In_2354);
xnor U298 (N_298,In_86,In_1032);
or U299 (N_299,In_1406,In_2458);
nand U300 (N_300,In_2289,In_1598);
nand U301 (N_301,In_1796,In_923);
or U302 (N_302,In_1871,In_2269);
nor U303 (N_303,In_2327,In_266);
or U304 (N_304,In_1762,In_426);
nor U305 (N_305,In_2652,In_208);
or U306 (N_306,In_2092,In_1888);
and U307 (N_307,In_271,In_2268);
and U308 (N_308,In_2161,In_1875);
xor U309 (N_309,In_1641,In_2589);
or U310 (N_310,In_1670,In_781);
nor U311 (N_311,In_203,In_1617);
xor U312 (N_312,In_2709,In_324);
or U313 (N_313,In_1186,In_1926);
xor U314 (N_314,In_2723,In_2782);
xnor U315 (N_315,In_2665,In_1427);
and U316 (N_316,In_2372,In_399);
xor U317 (N_317,In_1761,In_2421);
xnor U318 (N_318,In_216,In_131);
xor U319 (N_319,In_2056,In_499);
and U320 (N_320,In_2274,In_2509);
and U321 (N_321,In_1522,In_1153);
xnor U322 (N_322,In_2389,In_851);
or U323 (N_323,In_1848,In_2588);
and U324 (N_324,In_1217,In_147);
and U325 (N_325,In_2251,In_110);
or U326 (N_326,In_482,In_705);
and U327 (N_327,In_1546,In_613);
or U328 (N_328,In_2364,In_2800);
and U329 (N_329,In_1042,In_1568);
or U330 (N_330,In_2680,In_1137);
nand U331 (N_331,In_857,In_2442);
xor U332 (N_332,In_2236,In_1187);
xnor U333 (N_333,In_798,In_2146);
and U334 (N_334,In_272,In_2398);
and U335 (N_335,In_2622,In_154);
xor U336 (N_336,In_251,In_2081);
and U337 (N_337,In_1890,In_992);
or U338 (N_338,In_2020,In_79);
and U339 (N_339,In_997,In_758);
xnor U340 (N_340,In_13,In_2848);
nor U341 (N_341,In_35,In_2826);
and U342 (N_342,In_2887,In_2933);
or U343 (N_343,In_201,In_2750);
xnor U344 (N_344,In_1911,In_210);
and U345 (N_345,In_1947,In_1764);
or U346 (N_346,In_1321,In_626);
and U347 (N_347,In_2302,In_2987);
nor U348 (N_348,In_524,In_1867);
xor U349 (N_349,In_1728,In_149);
nor U350 (N_350,In_2528,In_871);
or U351 (N_351,In_930,In_2504);
nor U352 (N_352,In_999,In_1712);
nand U353 (N_353,In_759,In_1036);
nor U354 (N_354,In_359,In_2423);
or U355 (N_355,In_2273,In_845);
and U356 (N_356,In_593,In_1152);
or U357 (N_357,In_2480,In_2787);
nor U358 (N_358,In_2834,In_1557);
and U359 (N_359,In_1328,In_2316);
nor U360 (N_360,In_650,In_1948);
and U361 (N_361,In_2446,In_2627);
nor U362 (N_362,In_811,In_1505);
xnor U363 (N_363,In_834,In_1046);
nand U364 (N_364,In_363,In_1699);
or U365 (N_365,In_1672,In_58);
or U366 (N_366,In_1106,In_1990);
nor U367 (N_367,In_1974,In_1847);
xnor U368 (N_368,In_1676,In_1041);
xnor U369 (N_369,In_2271,In_406);
nor U370 (N_370,In_2525,In_1873);
xnor U371 (N_371,In_492,In_652);
or U372 (N_372,In_2953,In_2647);
nand U373 (N_373,In_2737,In_50);
and U374 (N_374,In_85,In_1403);
xor U375 (N_375,In_1669,In_2465);
nand U376 (N_376,In_2386,In_842);
or U377 (N_377,In_2122,In_598);
xnor U378 (N_378,In_1826,In_1214);
or U379 (N_379,In_2260,In_2357);
xor U380 (N_380,In_1562,In_436);
nand U381 (N_381,In_553,In_1206);
nor U382 (N_382,In_1366,In_1902);
and U383 (N_383,In_2263,In_1683);
nand U384 (N_384,In_866,In_911);
nor U385 (N_385,In_2875,In_2615);
or U386 (N_386,In_468,In_1680);
nor U387 (N_387,In_1091,In_622);
xor U388 (N_388,In_2654,In_2220);
and U389 (N_389,In_2033,In_2590);
nor U390 (N_390,In_566,In_2473);
nor U391 (N_391,In_1114,In_2339);
nand U392 (N_392,In_1243,In_2297);
nor U393 (N_393,In_1689,In_20);
xor U394 (N_394,In_2054,In_2438);
and U395 (N_395,In_1070,In_2934);
nor U396 (N_396,In_2094,In_312);
or U397 (N_397,In_916,In_2632);
xor U398 (N_398,In_39,In_914);
or U399 (N_399,In_1778,In_1968);
nand U400 (N_400,In_772,In_2978);
nor U401 (N_401,In_2852,In_1297);
nor U402 (N_402,In_608,In_1793);
nor U403 (N_403,In_1602,In_1448);
nand U404 (N_404,In_2673,In_1782);
xnor U405 (N_405,In_162,In_740);
nand U406 (N_406,In_2223,In_2214);
nor U407 (N_407,In_685,In_100);
or U408 (N_408,In_332,In_1819);
nand U409 (N_409,In_1549,In_104);
or U410 (N_410,In_557,In_296);
nand U411 (N_411,In_371,In_550);
and U412 (N_412,In_942,In_2948);
nand U413 (N_413,In_1516,In_780);
nand U414 (N_414,In_2935,In_458);
xor U415 (N_415,In_1318,In_1216);
nor U416 (N_416,In_2986,In_2091);
nor U417 (N_417,In_1204,In_1197);
nand U418 (N_418,In_2380,In_2449);
or U419 (N_419,In_1477,In_151);
and U420 (N_420,In_586,In_265);
nor U421 (N_421,In_489,In_1561);
or U422 (N_422,In_636,In_1432);
nor U423 (N_423,In_2299,In_108);
nor U424 (N_424,In_2295,In_2844);
xnor U425 (N_425,In_1309,In_1320);
nor U426 (N_426,In_2021,In_1444);
and U427 (N_427,In_469,In_1426);
or U428 (N_428,In_2451,In_1013);
and U429 (N_429,In_2264,In_656);
nor U430 (N_430,In_198,In_2238);
nand U431 (N_431,In_1542,In_1820);
nand U432 (N_432,In_612,In_2337);
and U433 (N_433,In_2052,In_1458);
xnor U434 (N_434,In_2858,In_1674);
or U435 (N_435,In_2725,In_1525);
nand U436 (N_436,In_2450,In_1688);
nand U437 (N_437,In_435,In_118);
xnor U438 (N_438,In_932,In_121);
xor U439 (N_439,In_1396,In_1580);
nand U440 (N_440,In_1791,In_2536);
nor U441 (N_441,In_697,In_1459);
or U442 (N_442,In_2688,In_2108);
nor U443 (N_443,In_134,In_1906);
nor U444 (N_444,In_1227,In_2624);
nand U445 (N_445,In_2506,In_1939);
and U446 (N_446,In_1054,In_1465);
or U447 (N_447,In_456,In_844);
and U448 (N_448,In_1855,In_1808);
or U449 (N_449,In_2625,In_2495);
xor U450 (N_450,In_111,In_1088);
or U451 (N_451,In_1183,In_2560);
or U452 (N_452,In_2352,In_785);
or U453 (N_453,In_168,In_960);
xor U454 (N_454,In_1655,In_1975);
and U455 (N_455,In_508,In_1260);
or U456 (N_456,In_2614,In_937);
or U457 (N_457,In_2773,In_2189);
or U458 (N_458,In_2591,In_575);
nand U459 (N_459,In_211,In_527);
nor U460 (N_460,In_2131,In_1719);
or U461 (N_461,In_1018,In_2287);
or U462 (N_462,In_934,In_415);
or U463 (N_463,In_1987,In_1910);
nand U464 (N_464,In_1239,In_2678);
xnor U465 (N_465,In_2835,In_345);
nand U466 (N_466,In_576,In_2025);
xor U467 (N_467,In_2909,In_1422);
or U468 (N_468,In_2781,In_239);
xnor U469 (N_469,In_1766,In_1919);
and U470 (N_470,In_882,In_1951);
nand U471 (N_471,In_1526,In_717);
nor U472 (N_472,In_144,In_106);
nand U473 (N_473,In_2109,In_2937);
and U474 (N_474,In_387,In_2483);
or U475 (N_475,In_962,In_184);
nand U476 (N_476,In_619,In_2195);
nor U477 (N_477,In_398,In_870);
xnor U478 (N_478,In_855,In_846);
xor U479 (N_479,In_1418,In_202);
or U480 (N_480,In_1113,In_1531);
or U481 (N_481,In_1480,In_565);
and U482 (N_482,In_1722,In_2405);
nand U483 (N_483,In_1653,In_940);
xor U484 (N_484,In_2672,In_2350);
and U485 (N_485,In_1980,In_2741);
or U486 (N_486,In_888,In_183);
nor U487 (N_487,In_2656,In_206);
and U488 (N_488,In_253,In_2008);
nand U489 (N_489,In_1901,In_526);
nand U490 (N_490,In_1547,In_1384);
and U491 (N_491,In_1414,In_2307);
or U492 (N_492,In_123,In_1298);
and U493 (N_493,In_2261,In_2873);
or U494 (N_494,In_875,In_1606);
nor U495 (N_495,In_2258,In_71);
nor U496 (N_496,In_2932,In_2891);
nand U497 (N_497,In_2927,In_1164);
nor U498 (N_498,In_1934,In_585);
nor U499 (N_499,In_728,In_46);
or U500 (N_500,In_1343,In_297);
xor U501 (N_501,In_2606,In_894);
or U502 (N_502,In_801,In_2655);
nand U503 (N_503,In_105,In_1700);
and U504 (N_504,In_385,In_2839);
xor U505 (N_505,In_5,In_2605);
xnor U506 (N_506,In_2172,In_1386);
nand U507 (N_507,In_136,In_2845);
or U508 (N_508,In_2675,In_433);
nor U509 (N_509,In_2587,In_2086);
and U510 (N_510,In_2312,In_2720);
or U511 (N_511,In_229,In_1635);
nand U512 (N_512,In_823,In_2626);
nand U513 (N_513,In_2424,In_525);
nand U514 (N_514,In_683,In_1854);
nor U515 (N_515,In_287,In_640);
nand U516 (N_516,In_1125,In_2028);
nand U517 (N_517,In_346,In_1369);
nand U518 (N_518,In_1794,In_393);
nand U519 (N_519,In_1962,In_2924);
xor U520 (N_520,In_310,In_1999);
xor U521 (N_521,In_642,In_126);
or U522 (N_522,In_633,In_2841);
and U523 (N_523,In_24,In_2899);
xnor U524 (N_524,In_462,In_189);
or U525 (N_525,In_742,In_778);
or U526 (N_526,In_822,In_2567);
nor U527 (N_527,In_102,In_1059);
and U528 (N_528,In_2950,In_2695);
or U529 (N_529,In_2892,In_60);
or U530 (N_530,In_1610,In_1038);
and U531 (N_531,In_2410,In_2790);
xor U532 (N_532,In_516,In_1563);
xor U533 (N_533,In_1368,In_2371);
and U534 (N_534,In_1828,In_2842);
or U535 (N_535,In_286,In_854);
xnor U536 (N_536,In_1534,In_2202);
or U537 (N_537,In_968,In_1389);
nand U538 (N_538,In_1520,In_1751);
and U539 (N_539,In_1401,In_961);
xor U540 (N_540,In_2005,In_1800);
nor U541 (N_541,In_248,In_2757);
and U542 (N_542,In_2707,In_2440);
nand U543 (N_543,In_1277,In_65);
and U544 (N_544,In_1502,In_475);
and U545 (N_545,In_2770,In_2819);
or U546 (N_546,In_2213,In_83);
nor U547 (N_547,In_2006,In_2740);
nor U548 (N_548,In_2461,In_752);
xor U549 (N_549,In_1491,In_1222);
nand U550 (N_550,In_2118,In_2190);
or U551 (N_551,In_2464,In_11);
xor U552 (N_552,In_965,In_2443);
nor U553 (N_553,In_1346,In_1096);
nand U554 (N_554,In_2944,In_438);
and U555 (N_555,In_437,In_2956);
xor U556 (N_556,In_194,In_377);
nand U557 (N_557,In_1628,In_2);
nand U558 (N_558,In_2619,In_2532);
and U559 (N_559,In_1457,In_1569);
nand U560 (N_560,In_1253,In_1276);
nor U561 (N_561,In_1893,In_1976);
or U562 (N_562,In_1189,In_351);
xor U563 (N_563,In_1978,In_535);
and U564 (N_564,In_2846,In_2481);
or U565 (N_565,In_637,In_1585);
and U566 (N_566,In_541,In_1618);
xor U567 (N_567,In_1231,In_2296);
or U568 (N_568,In_1639,In_293);
and U569 (N_569,In_504,In_2609);
nor U570 (N_570,In_2123,In_2497);
and U571 (N_571,In_1311,In_2601);
nor U572 (N_572,In_571,In_1402);
xnor U573 (N_573,In_936,In_1813);
nand U574 (N_574,In_1586,In_338);
nand U575 (N_575,In_852,In_1904);
or U576 (N_576,In_1524,In_2889);
nand U577 (N_577,In_64,In_1154);
or U578 (N_578,In_1891,In_143);
xnor U579 (N_579,In_2221,In_671);
nand U580 (N_580,In_2951,In_1008);
nor U581 (N_581,In_2729,In_926);
xnor U582 (N_582,In_2230,In_605);
or U583 (N_583,In_68,In_2939);
nor U584 (N_584,In_1035,In_2769);
xor U585 (N_585,In_87,In_714);
nor U586 (N_586,In_1755,In_2397);
nand U587 (N_587,In_2207,In_278);
xor U588 (N_588,In_1066,In_2104);
nand U589 (N_589,In_1284,In_1141);
and U590 (N_590,In_1932,In_2272);
nor U591 (N_591,In_2320,In_488);
xnor U592 (N_592,In_496,In_2799);
nand U593 (N_593,In_1814,In_1946);
xnor U594 (N_594,In_2507,In_1249);
nor U595 (N_595,In_2136,In_1779);
or U596 (N_596,In_1234,In_1339);
nand U597 (N_597,In_2708,In_1199);
xnor U598 (N_598,In_59,In_2275);
nor U599 (N_599,In_2066,In_931);
or U600 (N_600,In_630,In_817);
nand U601 (N_601,In_2404,In_1467);
and U602 (N_602,In_1528,In_280);
nor U603 (N_603,In_2667,In_1648);
nor U604 (N_604,In_1223,In_2597);
and U605 (N_605,In_2919,In_1241);
nand U606 (N_606,In_1874,In_2637);
nand U607 (N_607,In_254,In_2566);
and U608 (N_608,In_624,In_2105);
xnor U609 (N_609,In_2183,In_644);
or U610 (N_610,In_1462,In_319);
nor U611 (N_611,In_2015,In_1388);
or U612 (N_612,In_1010,In_167);
nand U613 (N_613,In_1604,In_1570);
or U614 (N_614,In_786,In_2281);
or U615 (N_615,In_186,In_1330);
xnor U616 (N_616,In_1151,In_1701);
nand U617 (N_617,In_1964,In_1673);
nor U618 (N_618,In_14,In_1455);
or U619 (N_619,In_2690,In_2246);
nor U620 (N_620,In_1882,In_1031);
xor U621 (N_621,In_2406,In_833);
nand U622 (N_622,In_299,In_370);
nor U623 (N_623,In_1028,In_2003);
nor U624 (N_624,In_1834,In_755);
and U625 (N_625,In_1603,In_2308);
nor U626 (N_626,In_2907,In_305);
nor U627 (N_627,In_794,In_1470);
xnor U628 (N_628,In_1272,In_139);
and U629 (N_629,In_891,In_1651);
nor U630 (N_630,In_1898,In_1450);
nor U631 (N_631,In_1841,In_1697);
xnor U632 (N_632,In_1846,In_2882);
or U633 (N_633,In_1892,In_1861);
nor U634 (N_634,In_2585,In_477);
or U635 (N_635,In_2616,In_2169);
nor U636 (N_636,In_1196,In_723);
nor U637 (N_637,In_985,In_712);
and U638 (N_638,In_2103,In_1860);
or U639 (N_639,In_2196,In_2367);
nand U640 (N_640,In_1045,In_1160);
xor U641 (N_641,In_2685,In_459);
or U642 (N_642,In_559,In_1588);
nor U643 (N_643,In_1282,In_2290);
nor U644 (N_644,In_1897,In_2477);
nand U645 (N_645,In_2178,In_783);
xor U646 (N_646,In_1734,In_1625);
nand U647 (N_647,In_1686,In_453);
nand U648 (N_648,In_2068,In_242);
and U649 (N_649,In_1917,In_2570);
xnor U650 (N_650,In_573,In_2662);
nand U651 (N_651,In_790,In_2329);
or U652 (N_652,In_2494,In_2285);
xor U653 (N_653,In_329,In_1002);
nand U654 (N_654,In_1864,In_1238);
and U655 (N_655,In_682,In_1363);
nand U656 (N_656,In_311,In_1738);
or U657 (N_657,In_326,In_2279);
nor U658 (N_658,In_384,In_1181);
nor U659 (N_659,In_1958,In_1918);
or U660 (N_660,In_1666,In_2156);
or U661 (N_661,In_2425,In_1109);
and U662 (N_662,In_1342,In_546);
and U663 (N_663,In_2783,In_1740);
nand U664 (N_664,In_2309,In_1314);
nor U665 (N_665,In_425,In_954);
nor U666 (N_666,In_140,In_9);
and U667 (N_667,In_2018,In_1202);
nor U668 (N_668,In_1702,In_2400);
or U669 (N_669,In_1743,In_32);
nor U670 (N_670,In_2955,In_620);
nor U671 (N_671,In_1730,In_1908);
xnor U672 (N_672,In_654,In_1937);
or U673 (N_673,In_2217,In_99);
nor U674 (N_674,In_1817,In_927);
and U675 (N_675,In_2441,In_1840);
or U676 (N_676,In_2650,In_1092);
xor U677 (N_677,In_455,In_42);
xnor U678 (N_678,In_2072,In_218);
xnor U679 (N_679,In_2245,In_432);
nand U680 (N_680,In_1374,In_1175);
nand U681 (N_681,In_978,In_1831);
nand U682 (N_682,In_1594,In_422);
and U683 (N_683,In_1072,In_2162);
and U684 (N_684,In_720,In_1952);
nor U685 (N_685,In_394,In_2485);
nor U686 (N_686,In_1748,In_2705);
xor U687 (N_687,In_1607,In_1267);
and U688 (N_688,In_2335,In_1087);
nand U689 (N_689,In_1896,In_673);
and U690 (N_690,In_1638,In_2181);
nand U691 (N_691,In_2871,In_1074);
xnor U692 (N_692,In_1021,In_241);
or U693 (N_693,In_1095,In_1127);
and U694 (N_694,In_300,In_1889);
nand U695 (N_695,In_2938,In_1279);
xor U696 (N_696,In_1662,In_2125);
and U697 (N_697,In_1977,In_938);
nand U698 (N_698,In_2422,In_2032);
and U699 (N_699,In_1647,In_2883);
nor U700 (N_700,In_611,In_2639);
nand U701 (N_701,In_1287,In_1460);
or U702 (N_702,In_862,In_2512);
xor U703 (N_703,In_2225,In_77);
xor U704 (N_704,In_2117,In_1105);
nor U705 (N_705,In_1737,In_994);
nand U706 (N_706,In_1134,In_1739);
or U707 (N_707,In_1622,In_45);
xor U708 (N_708,In_1720,In_288);
and U709 (N_709,In_1259,In_577);
nor U710 (N_710,In_2874,In_12);
nand U711 (N_711,In_2716,In_2130);
nand U712 (N_712,In_2265,In_430);
nor U713 (N_713,In_2474,In_330);
nor U714 (N_714,In_231,In_1629);
or U715 (N_715,In_1312,In_2890);
xor U716 (N_716,In_707,In_2711);
nor U717 (N_717,In_119,In_1377);
and U718 (N_718,In_869,In_2224);
xor U719 (N_719,In_2305,In_2132);
or U720 (N_720,In_1507,In_1244);
and U721 (N_721,In_2433,In_412);
nor U722 (N_722,In_2573,In_2657);
nor U723 (N_723,In_2459,In_444);
xor U724 (N_724,In_1880,In_1097);
or U725 (N_725,In_282,In_2492);
and U726 (N_726,In_2789,In_950);
xor U727 (N_727,In_448,In_1325);
or U728 (N_728,In_1626,In_1344);
or U729 (N_729,In_539,In_1138);
xor U730 (N_730,In_418,In_1513);
or U731 (N_731,In_1986,In_1825);
nor U732 (N_732,In_1818,In_935);
nand U733 (N_733,In_2689,In_1945);
and U734 (N_734,In_2539,In_1156);
xnor U735 (N_735,In_963,In_2137);
xnor U736 (N_736,In_2968,In_1464);
xor U737 (N_737,In_486,In_2179);
or U738 (N_738,In_30,In_2097);
or U739 (N_739,In_807,In_672);
and U740 (N_740,In_922,In_841);
nor U741 (N_741,In_1078,In_2954);
nand U742 (N_742,In_146,In_103);
or U743 (N_743,In_2501,In_2152);
and U744 (N_744,In_2611,In_1262);
and U745 (N_745,In_2431,In_1413);
and U746 (N_746,In_2291,In_133);
nand U747 (N_747,In_366,In_1789);
or U748 (N_748,In_1929,In_1573);
nor U749 (N_749,In_1212,In_107);
and U750 (N_750,In_2009,In_473);
nor U751 (N_751,In_513,In_1264);
nor U752 (N_752,In_155,In_2610);
or U753 (N_753,In_2976,In_1023);
xnor U754 (N_754,In_518,In_269);
nand U755 (N_755,In_1756,In_2294);
nand U756 (N_756,In_72,In_809);
xnor U757 (N_757,In_1173,In_956);
and U758 (N_758,In_1446,In_2078);
or U759 (N_759,In_629,In_1390);
or U760 (N_760,In_2001,In_599);
and U761 (N_761,In_1581,In_2660);
and U762 (N_762,In_2313,In_666);
xnor U763 (N_763,In_2840,In_160);
and U764 (N_764,In_1685,In_1620);
and U765 (N_765,In_2099,In_382);
and U766 (N_766,In_2144,In_2325);
and U767 (N_767,In_245,In_990);
and U768 (N_768,In_2771,In_1188);
nor U769 (N_769,In_711,In_178);
or U770 (N_770,In_517,In_1302);
nand U771 (N_771,In_2996,In_1548);
nor U772 (N_772,In_2143,In_49);
or U773 (N_773,In_1969,In_1691);
and U774 (N_774,In_2869,In_112);
and U775 (N_775,In_318,In_750);
and U776 (N_776,In_1575,In_56);
and U777 (N_777,In_1266,In_465);
nor U778 (N_778,In_15,In_2975);
or U779 (N_779,In_1081,In_1304);
or U780 (N_780,In_2383,In_2408);
and U781 (N_781,In_2599,In_872);
and U782 (N_782,In_2301,In_951);
nand U783 (N_783,In_2602,In_500);
and U784 (N_784,In_323,In_2158);
and U785 (N_785,In_1177,In_606);
nand U786 (N_786,In_819,In_2989);
nor U787 (N_787,In_1417,In_1839);
xnor U788 (N_788,In_1633,In_591);
nor U789 (N_789,In_1265,In_1089);
and U790 (N_790,In_1886,In_568);
nor U791 (N_791,In_1103,In_368);
xnor U792 (N_792,In_2693,In_2984);
and U793 (N_793,In_2326,In_722);
or U794 (N_794,In_1922,In_1345);
and U795 (N_795,In_1997,In_1965);
xor U796 (N_796,In_442,In_2556);
nor U797 (N_797,In_2628,In_1744);
and U798 (N_798,In_2374,In_2476);
xnor U799 (N_799,In_397,In_2533);
nor U800 (N_800,In_376,In_41);
nor U801 (N_801,In_1843,In_2925);
nor U802 (N_802,In_1323,In_391);
xor U803 (N_803,In_1380,In_2894);
or U804 (N_804,In_2379,In_986);
xor U805 (N_805,In_1790,In_799);
xnor U806 (N_806,In_1624,In_2242);
or U807 (N_807,In_320,In_2229);
and U808 (N_808,In_1080,In_2554);
xnor U809 (N_809,In_2527,In_180);
xor U810 (N_810,In_2469,In_94);
or U811 (N_811,In_1924,In_1250);
xnor U812 (N_812,In_1016,In_523);
nor U813 (N_813,In_1121,In_1185);
nor U814 (N_814,In_972,In_1705);
xor U815 (N_815,In_2731,In_2344);
and U816 (N_816,In_2027,In_1495);
nand U817 (N_817,In_1724,In_2176);
and U818 (N_818,In_2159,In_1577);
xnor U819 (N_819,In_2969,In_361);
xnor U820 (N_820,In_2075,In_648);
and U821 (N_821,In_2981,In_2535);
and U822 (N_822,In_977,In_336);
xnor U823 (N_823,In_1077,In_534);
nor U824 (N_824,In_639,In_303);
nor U825 (N_825,In_788,In_1463);
nor U826 (N_826,In_1195,In_1085);
nand U827 (N_827,In_1131,In_2926);
xor U828 (N_828,In_2233,In_858);
nand U829 (N_829,In_1916,In_2592);
or U830 (N_830,In_1283,In_765);
or U831 (N_831,In_925,In_1142);
xor U832 (N_832,In_2062,In_902);
xnor U833 (N_833,In_1681,In_1120);
and U834 (N_834,In_1885,In_1425);
or U835 (N_835,In_2990,In_2663);
and U836 (N_836,In_1930,In_2048);
and U837 (N_837,In_2300,In_52);
xor U838 (N_838,In_261,In_1001);
nand U839 (N_839,In_2912,In_308);
xnor U840 (N_840,In_709,In_2468);
or U841 (N_841,In_2510,In_2429);
or U842 (N_842,In_1146,In_1452);
or U843 (N_843,In_1128,In_1803);
and U844 (N_844,In_1291,In_1352);
and U845 (N_845,In_1410,In_2797);
or U846 (N_846,In_1775,In_2306);
and U847 (N_847,In_737,In_2445);
and U848 (N_848,In_1347,In_2411);
nor U849 (N_849,In_55,In_1872);
nand U850 (N_850,In_414,In_1644);
nand U851 (N_851,In_2163,In_1771);
and U852 (N_852,In_1614,In_2721);
nand U853 (N_853,In_1486,In_313);
nor U854 (N_854,In_1589,In_1441);
nand U855 (N_855,In_88,In_18);
nand U856 (N_856,In_1361,In_2171);
or U857 (N_857,In_1876,In_84);
xnor U858 (N_858,In_1079,In_1710);
and U859 (N_859,In_831,In_2843);
nor U860 (N_860,In_2962,In_2792);
or U861 (N_861,In_2607,In_171);
nand U862 (N_862,In_1271,In_2565);
nor U863 (N_863,In_148,In_1218);
or U864 (N_864,In_1785,In_1357);
nor U865 (N_865,In_1497,In_2037);
or U866 (N_866,In_2640,In_850);
xnor U867 (N_867,In_481,In_1193);
or U868 (N_868,In_130,In_1118);
and U869 (N_869,In_2282,In_1483);
xor U870 (N_870,In_1069,In_2083);
or U871 (N_871,In_1338,In_837);
and U872 (N_872,In_2278,In_1449);
or U873 (N_873,In_1382,In_1159);
nand U874 (N_874,In_987,In_1844);
nor U875 (N_875,In_2762,In_1161);
nor U876 (N_876,In_674,In_2677);
xor U877 (N_877,In_1942,In_240);
or U878 (N_878,In_207,In_684);
and U879 (N_879,In_2714,In_2382);
or U880 (N_880,In_2767,In_522);
xnor U881 (N_881,In_718,In_2633);
nor U882 (N_882,In_900,In_2903);
and U883 (N_883,In_298,In_1294);
or U884 (N_884,In_643,In_2157);
nor U885 (N_885,In_1512,In_247);
xnor U886 (N_886,In_2321,In_532);
xor U887 (N_887,In_1913,In_2904);
nor U888 (N_888,In_1240,In_2049);
nor U889 (N_889,In_627,In_2830);
and U890 (N_890,In_1112,In_2203);
nand U891 (N_891,In_2726,In_80);
and U892 (N_892,In_2576,In_2470);
and U893 (N_893,In_471,In_2457);
nand U894 (N_894,In_2801,In_2728);
nand U895 (N_895,In_1473,In_2897);
and U896 (N_896,In_1333,In_2571);
xor U897 (N_897,In_1215,In_1695);
nand U898 (N_898,In_1909,In_1895);
xor U899 (N_899,In_706,In_564);
xor U900 (N_900,In_829,In_66);
or U901 (N_901,In_621,In_1058);
and U902 (N_902,In_2039,In_2795);
nor U903 (N_903,In_124,In_2288);
nor U904 (N_904,In_1157,In_1592);
and U905 (N_905,In_2778,In_1431);
and U906 (N_906,In_1550,In_2872);
nand U907 (N_907,In_1661,In_182);
nor U908 (N_908,In_618,In_1305);
or U909 (N_909,In_601,In_958);
and U910 (N_910,In_1654,In_2215);
or U911 (N_911,In_410,In_2674);
nand U912 (N_912,In_2979,In_689);
and U913 (N_913,In_1370,In_413);
nand U914 (N_914,In_1365,In_2557);
or U915 (N_915,In_395,In_2983);
and U916 (N_916,In_1971,In_1148);
or U917 (N_917,In_2074,In_2965);
nand U918 (N_918,In_2336,In_327);
nand U919 (N_919,In_2712,In_821);
and U920 (N_920,In_1601,In_1576);
and U921 (N_921,In_383,In_943);
or U922 (N_922,In_1656,In_2167);
nand U923 (N_923,In_2491,In_2040);
or U924 (N_924,In_2545,In_2358);
nor U925 (N_925,In_1665,In_897);
nand U926 (N_926,In_2811,In_887);
or U927 (N_927,In_114,In_825);
and U928 (N_928,In_2147,In_1433);
nor U929 (N_929,In_1006,In_1233);
nor U930 (N_930,In_2407,In_582);
nand U931 (N_931,In_1879,In_1050);
or U932 (N_932,In_1274,In_321);
and U933 (N_933,In_2043,In_2166);
and U934 (N_934,In_2479,In_1071);
xor U935 (N_935,In_519,In_2908);
xnor U936 (N_936,In_1984,In_906);
nand U937 (N_937,In_2620,In_1051);
nor U938 (N_938,In_62,In_628);
nor U939 (N_939,In_889,In_2853);
and U940 (N_940,In_1690,In_2730);
or U941 (N_941,In_567,In_362);
xnor U942 (N_942,In_2943,In_774);
and U943 (N_943,In_570,In_588);
and U944 (N_944,In_1853,In_224);
and U945 (N_945,In_2881,In_1167);
nand U946 (N_946,In_355,In_2743);
nand U947 (N_947,In_982,In_2496);
nand U948 (N_948,In_863,In_1907);
nor U949 (N_949,In_2763,In_1687);
or U950 (N_950,In_21,In_2373);
xnor U951 (N_951,In_2923,In_1170);
nor U952 (N_952,In_773,In_2362);
nand U953 (N_953,In_2259,In_646);
nand U954 (N_954,In_2682,In_400);
or U955 (N_955,In_2812,In_2715);
nand U956 (N_956,In_421,In_90);
nor U957 (N_957,In_233,In_1348);
and U958 (N_958,In_1367,In_724);
or U959 (N_959,In_1989,In_2444);
or U960 (N_960,In_2898,In_1733);
or U961 (N_961,In_756,In_1725);
and U962 (N_962,In_2736,In_768);
nor U963 (N_963,In_2249,In_1052);
nor U964 (N_964,In_427,In_2704);
xor U965 (N_965,In_2564,In_1824);
xnor U966 (N_966,In_2333,In_1567);
or U967 (N_967,In_2594,In_1288);
or U968 (N_968,In_595,In_2430);
and U969 (N_969,In_2016,In_1428);
nand U970 (N_970,In_2568,In_838);
nand U971 (N_971,In_2314,In_306);
xor U972 (N_972,In_1319,In_1381);
and U973 (N_973,In_1232,In_2745);
xnor U974 (N_974,In_2073,In_917);
nor U975 (N_975,In_1858,In_1155);
and U976 (N_976,In_2856,In_1407);
nand U977 (N_977,In_769,In_2462);
or U978 (N_978,In_1998,In_2867);
nand U979 (N_979,In_1144,In_2107);
xnor U980 (N_980,In_1726,In_2188);
nor U981 (N_981,In_2888,In_1936);
or U982 (N_982,In_2100,In_721);
or U983 (N_983,In_2549,In_903);
nor U984 (N_984,In_1802,In_1438);
nand U985 (N_985,In_1508,In_2558);
nand U986 (N_986,In_2447,In_1752);
and U987 (N_987,In_2502,In_2717);
xnor U988 (N_988,In_1583,In_2960);
and U989 (N_989,In_1126,In_374);
xor U990 (N_990,In_236,In_973);
or U991 (N_991,In_2646,In_1061);
xor U992 (N_992,In_196,In_2051);
or U993 (N_993,In_1551,In_2684);
xor U994 (N_994,In_617,In_775);
xnor U995 (N_995,In_2859,In_2920);
nor U996 (N_996,In_702,In_1399);
and U997 (N_997,In_2719,In_738);
and U998 (N_998,In_1488,In_2905);
or U999 (N_999,In_277,In_1242);
or U1000 (N_1000,In_681,N_143);
and U1001 (N_1001,N_509,In_1424);
xor U1002 (N_1002,In_912,In_205);
xor U1003 (N_1003,N_19,In_2562);
xnor U1004 (N_1004,In_480,In_2432);
and U1005 (N_1005,N_208,N_102);
nor U1006 (N_1006,N_595,N_785);
xnor U1007 (N_1007,In_2142,N_868);
and U1008 (N_1008,N_243,In_1812);
and U1009 (N_1009,N_370,In_2415);
xnor U1010 (N_1010,In_1530,In_615);
nand U1011 (N_1011,N_606,N_359);
or U1012 (N_1012,In_1408,N_696);
nor U1013 (N_1013,N_550,In_2418);
nand U1014 (N_1014,In_1025,N_909);
xnor U1015 (N_1015,In_1935,In_1224);
nor U1016 (N_1016,N_714,N_819);
or U1017 (N_1017,In_159,N_400);
and U1018 (N_1018,In_75,In_2831);
and U1019 (N_1019,In_2403,N_609);
xor U1020 (N_1020,N_150,In_1804);
or U1021 (N_1021,In_1535,In_199);
or U1022 (N_1022,N_495,In_645);
nor U1023 (N_1023,N_892,N_48);
and U1024 (N_1024,In_974,N_818);
xor U1025 (N_1025,In_1351,In_1063);
xor U1026 (N_1026,N_731,N_300);
or U1027 (N_1027,In_1955,N_457);
and U1028 (N_1028,N_860,In_2240);
nand U1029 (N_1029,N_981,In_2600);
nand U1030 (N_1030,In_686,N_753);
xor U1031 (N_1031,N_418,In_343);
nand U1032 (N_1032,N_893,In_614);
and U1033 (N_1033,N_412,In_607);
nor U1034 (N_1034,N_752,N_487);
xor U1035 (N_1035,In_2617,In_2780);
and U1036 (N_1036,N_730,N_494);
nand U1037 (N_1037,N_917,N_596);
and U1038 (N_1038,N_183,N_220);
or U1039 (N_1039,N_223,N_637);
and U1040 (N_1040,N_541,N_666);
or U1041 (N_1041,In_2193,In_2345);
nor U1042 (N_1042,N_958,In_991);
xor U1043 (N_1043,In_2644,N_771);
nand U1044 (N_1044,In_2958,In_214);
or U1045 (N_1045,In_2254,In_2168);
and U1046 (N_1046,In_1049,In_116);
and U1047 (N_1047,In_690,N_355);
nor U1048 (N_1048,In_1437,In_222);
nor U1049 (N_1049,In_228,In_760);
nand U1050 (N_1050,In_95,In_2880);
and U1051 (N_1051,In_2649,In_1122);
or U1052 (N_1052,In_1634,In_1104);
nor U1053 (N_1053,N_693,N_559);
nor U1054 (N_1054,In_1340,N_361);
nor U1055 (N_1055,In_2079,In_1116);
xor U1056 (N_1056,N_504,N_743);
nand U1057 (N_1057,In_1995,N_482);
xor U1058 (N_1058,N_451,N_554);
and U1059 (N_1059,In_1784,N_997);
xnor U1060 (N_1060,In_2722,N_66);
nor U1061 (N_1061,In_1201,N_969);
nand U1062 (N_1062,In_2396,In_2929);
and U1063 (N_1063,In_1660,N_147);
xnor U1064 (N_1064,N_832,In_677);
nand U1065 (N_1065,In_736,N_111);
nand U1066 (N_1066,In_409,In_560);
and U1067 (N_1067,N_564,In_289);
nor U1068 (N_1068,N_939,In_2061);
nor U1069 (N_1069,In_1836,N_280);
xnor U1070 (N_1070,In_407,N_81);
nand U1071 (N_1071,N_773,In_2914);
nand U1072 (N_1072,N_191,N_496);
xor U1073 (N_1073,In_784,N_789);
or U1074 (N_1074,In_727,In_1527);
nor U1075 (N_1075,In_1364,In_2000);
and U1076 (N_1076,In_1842,In_1037);
xor U1077 (N_1077,N_503,N_688);
or U1078 (N_1078,In_1950,N_960);
or U1079 (N_1079,N_650,In_1514);
or U1080 (N_1080,N_22,In_2531);
or U1081 (N_1081,In_983,N_281);
xnor U1082 (N_1082,In_507,In_138);
and U1083 (N_1083,In_325,In_2949);
xnor U1084 (N_1084,In_1636,N_757);
xnor U1085 (N_1085,N_101,In_1211);
nor U1086 (N_1086,N_110,N_410);
xnor U1087 (N_1087,In_551,In_54);
and U1088 (N_1088,N_404,In_113);
or U1089 (N_1089,In_1692,In_2997);
or U1090 (N_1090,In_1807,N_464);
or U1091 (N_1091,In_2893,In_1827);
and U1092 (N_1092,N_431,In_893);
and U1093 (N_1093,N_58,In_497);
nand U1094 (N_1094,N_718,In_304);
nand U1095 (N_1095,In_2298,N_29);
or U1096 (N_1096,In_101,N_69);
or U1097 (N_1097,N_423,N_240);
or U1098 (N_1098,N_970,In_2931);
and U1099 (N_1099,In_2250,In_2930);
or U1100 (N_1100,N_672,N_310);
nor U1101 (N_1101,In_28,N_536);
and U1102 (N_1102,N_699,In_2084);
and U1103 (N_1103,In_250,In_479);
nor U1104 (N_1104,In_1469,In_257);
or U1105 (N_1105,In_2774,In_1931);
nor U1106 (N_1106,N_252,N_669);
and U1107 (N_1107,In_1292,N_235);
nor U1108 (N_1108,N_364,N_739);
and U1109 (N_1109,In_2419,N_397);
xor U1110 (N_1110,N_354,N_14);
nand U1111 (N_1111,N_36,In_348);
xnor U1112 (N_1112,N_471,In_237);
or U1113 (N_1113,In_2901,In_984);
or U1114 (N_1114,N_237,N_684);
nor U1115 (N_1115,N_373,N_568);
nor U1116 (N_1116,N_758,N_141);
xor U1117 (N_1117,N_857,N_995);
xor U1118 (N_1118,In_904,N_184);
or U1119 (N_1119,N_793,N_203);
xnor U1120 (N_1120,N_545,N_13);
nor U1121 (N_1121,In_2866,N_999);
or U1122 (N_1122,In_2376,In_2520);
and U1123 (N_1123,N_906,In_578);
xor U1124 (N_1124,N_867,N_107);
nor U1125 (N_1125,In_259,N_941);
or U1126 (N_1126,In_657,In_2488);
xor U1127 (N_1127,In_531,N_133);
xnor U1128 (N_1128,N_389,N_705);
nor U1129 (N_1129,N_196,N_529);
and U1130 (N_1130,N_266,In_770);
xnor U1131 (N_1131,N_472,N_303);
xnor U1132 (N_1132,N_570,N_646);
nand U1133 (N_1133,N_493,In_651);
nand U1134 (N_1134,In_1940,In_915);
nand U1135 (N_1135,N_591,N_530);
xor U1136 (N_1136,In_544,In_864);
nand U1137 (N_1137,N_916,N_826);
or U1138 (N_1138,In_584,N_745);
nor U1139 (N_1139,In_2553,In_63);
nor U1140 (N_1140,N_314,In_2959);
and U1141 (N_1141,N_667,In_2786);
xnor U1142 (N_1142,N_862,In_2643);
or U1143 (N_1143,N_119,N_94);
xnor U1144 (N_1144,In_53,N_352);
and U1145 (N_1145,In_2035,N_113);
nand U1146 (N_1146,In_1708,In_2582);
and U1147 (N_1147,In_1261,In_2581);
or U1148 (N_1148,In_676,In_880);
and U1149 (N_1149,N_258,In_971);
xnor U1150 (N_1150,N_70,In_2187);
nor U1151 (N_1151,N_118,N_505);
or U1152 (N_1152,In_1816,In_2998);
nand U1153 (N_1153,In_2860,In_16);
nand U1154 (N_1154,N_889,N_134);
xor U1155 (N_1155,N_181,N_169);
nand U1156 (N_1156,N_348,N_976);
nor U1157 (N_1157,In_1613,In_1487);
or U1158 (N_1158,N_786,In_390);
or U1159 (N_1159,N_930,N_288);
nor U1160 (N_1160,N_876,In_744);
or U1161 (N_1161,N_737,In_279);
or U1162 (N_1162,In_1767,In_246);
nor U1163 (N_1163,N_656,In_2164);
and U1164 (N_1164,N_695,In_2113);
nor U1165 (N_1165,N_883,N_34);
xor U1166 (N_1166,In_1815,In_2255);
nor U1167 (N_1167,In_268,N_201);
or U1168 (N_1168,In_290,In_1979);
nor U1169 (N_1169,N_766,In_188);
and U1170 (N_1170,In_2452,In_1773);
nor U1171 (N_1171,N_160,N_61);
and U1172 (N_1172,N_242,N_172);
and U1173 (N_1173,In_291,In_1612);
xor U1174 (N_1174,In_1246,In_2191);
or U1175 (N_1175,In_2209,In_1226);
nor U1176 (N_1176,N_275,In_1596);
and U1177 (N_1177,N_468,N_709);
nand U1178 (N_1178,In_1597,In_416);
xor U1179 (N_1179,In_2243,In_1252);
or U1180 (N_1180,N_847,In_2154);
xnor U1181 (N_1181,In_746,N_946);
xor U1182 (N_1182,In_594,In_1165);
nor U1183 (N_1183,N_152,In_354);
nor U1184 (N_1184,In_1039,In_1552);
nand U1185 (N_1185,In_1331,N_136);
nand U1186 (N_1186,N_896,N_304);
xnor U1187 (N_1187,In_998,N_108);
nor U1188 (N_1188,N_95,In_2753);
nor U1189 (N_1189,N_987,In_2276);
nor U1190 (N_1190,N_131,In_70);
nor U1191 (N_1191,N_782,N_28);
xor U1192 (N_1192,N_578,In_1510);
nand U1193 (N_1193,In_2824,N_236);
or U1194 (N_1194,N_866,N_526);
nor U1195 (N_1195,N_700,In_2526);
or U1196 (N_1196,N_837,N_719);
nor U1197 (N_1197,N_791,N_406);
nand U1198 (N_1198,N_188,In_957);
xnor U1199 (N_1199,N_659,N_973);
xor U1200 (N_1200,In_1394,N_214);
or U1201 (N_1201,In_495,In_401);
and U1202 (N_1202,In_1315,N_881);
or U1203 (N_1203,N_60,In_490);
and U1204 (N_1204,In_757,In_2529);
or U1205 (N_1205,In_10,N_90);
xor U1206 (N_1206,In_2472,N_315);
or U1207 (N_1207,In_1334,In_31);
nor U1208 (N_1208,N_897,N_453);
nor U1209 (N_1209,In_1019,In_152);
nand U1210 (N_1210,N_522,N_600);
nand U1211 (N_1211,N_543,In_2814);
and U1212 (N_1212,N_694,N_843);
xnor U1213 (N_1213,N_372,In_2311);
nand U1214 (N_1214,N_575,In_2455);
or U1215 (N_1215,In_1353,N_53);
xnor U1216 (N_1216,In_2837,N_422);
xor U1217 (N_1217,In_2173,In_2578);
nor U1218 (N_1218,N_27,N_661);
nand U1219 (N_1219,N_754,In_1075);
nand U1220 (N_1220,N_768,In_688);
nor U1221 (N_1221,In_1678,N_935);
nor U1222 (N_1222,N_247,In_771);
xnor U1223 (N_1223,In_2945,In_78);
xor U1224 (N_1224,In_1171,N_31);
and U1225 (N_1225,In_2936,N_989);
and U1226 (N_1226,In_665,N_72);
nor U1227 (N_1227,In_933,N_100);
and U1228 (N_1228,In_1694,N_467);
and U1229 (N_1229,In_1047,In_2486);
or U1230 (N_1230,In_1101,In_2540);
nand U1231 (N_1231,In_405,N_460);
nand U1232 (N_1232,In_1048,In_867);
nor U1233 (N_1233,In_1894,N_475);
nor U1234 (N_1234,N_800,In_452);
xnor U1235 (N_1235,In_419,In_946);
xnor U1236 (N_1236,N_980,In_1313);
nor U1237 (N_1237,N_286,In_2661);
nor U1238 (N_1238,In_2825,N_702);
or U1239 (N_1239,In_2355,In_856);
nor U1240 (N_1240,N_648,In_533);
nor U1241 (N_1241,N_951,N_120);
nor U1242 (N_1242,In_165,In_2521);
xnor U1243 (N_1243,N_949,N_259);
xnor U1244 (N_1244,In_2756,N_498);
xnor U1245 (N_1245,In_908,N_879);
nor U1246 (N_1246,N_994,In_2974);
and U1247 (N_1247,In_2234,N_124);
nand U1248 (N_1248,In_1456,N_921);
nor U1249 (N_1249,N_50,In_337);
or U1250 (N_1250,In_2827,In_2815);
nor U1251 (N_1251,In_1677,In_1970);
nor U1252 (N_1252,N_337,N_357);
or U1253 (N_1253,N_846,In_1411);
nor U1254 (N_1254,In_169,In_467);
nand U1255 (N_1255,In_373,N_605);
or U1256 (N_1256,N_388,In_2023);
and U1257 (N_1257,In_1501,N_747);
xor U1258 (N_1258,In_1475,In_2641);
nor U1259 (N_1259,N_407,N_769);
xnor U1260 (N_1260,In_2911,In_693);
xor U1261 (N_1261,In_341,N_56);
nand U1262 (N_1262,In_1630,N_115);
xor U1263 (N_1263,In_2366,In_1856);
nor U1264 (N_1264,N_116,N_187);
xor U1265 (N_1265,In_2694,In_166);
nor U1266 (N_1266,N_226,In_2069);
or U1267 (N_1267,In_806,In_2813);
xor U1268 (N_1268,In_2779,N_566);
or U1269 (N_1269,In_2973,N_362);
nor U1270 (N_1270,N_391,N_828);
xnor U1271 (N_1271,N_74,In_43);
and U1272 (N_1272,N_379,N_200);
nor U1273 (N_1273,In_1565,N_142);
nand U1274 (N_1274,In_2658,In_1887);
nand U1275 (N_1275,In_96,In_2544);
and U1276 (N_1276,N_409,In_1845);
or U1277 (N_1277,In_2089,In_1003);
and U1278 (N_1278,N_830,N_783);
nand U1279 (N_1279,N_855,In_2493);
and U1280 (N_1280,N_256,N_603);
and U1281 (N_1281,In_981,In_1482);
nand U1282 (N_1282,N_154,In_29);
nand U1283 (N_1283,N_998,In_2952);
xnor U1284 (N_1284,In_379,In_964);
xor U1285 (N_1285,In_2456,N_540);
and U1286 (N_1286,In_1996,In_2205);
and U1287 (N_1287,N_628,N_427);
nor U1288 (N_1288,In_2776,In_2247);
xor U1289 (N_1289,In_562,In_1022);
and U1290 (N_1290,In_1511,N_399);
or U1291 (N_1291,N_80,In_2200);
nand U1292 (N_1292,N_485,N_219);
nand U1293 (N_1293,In_1273,N_531);
xnor U1294 (N_1294,N_905,N_318);
and U1295 (N_1295,N_283,In_2706);
nor U1296 (N_1296,In_2010,N_416);
nor U1297 (N_1297,In_694,In_924);
and U1298 (N_1298,N_307,In_1943);
nor U1299 (N_1299,N_320,N_452);
and U1300 (N_1300,N_164,In_1642);
nor U1301 (N_1301,N_454,N_98);
and U1302 (N_1302,In_2252,In_1278);
and U1303 (N_1303,In_263,In_2522);
nor U1304 (N_1304,In_832,N_805);
or U1305 (N_1305,In_1057,N_10);
or U1306 (N_1306,N_913,In_1703);
and U1307 (N_1307,In_2963,N_262);
nor U1308 (N_1308,N_105,In_886);
or U1309 (N_1309,In_2696,In_1938);
nand U1310 (N_1310,In_1566,N_647);
xor U1311 (N_1311,N_325,N_16);
xor U1312 (N_1312,In_2877,N_439);
and U1313 (N_1313,In_333,N_992);
xnor U1314 (N_1314,In_975,In_955);
xnor U1315 (N_1315,N_815,N_232);
xor U1316 (N_1316,In_859,N_971);
nor U1317 (N_1317,N_222,In_1416);
xnor U1318 (N_1318,In_466,N_518);
and U1319 (N_1319,In_2788,N_770);
nand U1320 (N_1320,In_2505,In_1506);
xnor U1321 (N_1321,N_25,N_49);
and U1322 (N_1322,N_681,N_502);
and U1323 (N_1323,In_2038,In_1082);
nor U1324 (N_1324,In_2237,N_724);
nor U1325 (N_1325,In_1360,In_1300);
and U1326 (N_1326,N_593,N_652);
and U1327 (N_1327,In_2384,In_602);
and U1328 (N_1328,In_1721,N_651);
nand U1329 (N_1329,In_270,N_145);
nand U1330 (N_1330,N_254,N_175);
or U1331 (N_1331,In_679,N_140);
nor U1332 (N_1332,N_982,In_309);
nor U1333 (N_1333,In_302,In_1529);
and U1334 (N_1334,In_1786,N_390);
or U1335 (N_1335,In_1519,N_0);
and U1336 (N_1336,N_733,In_334);
nor U1337 (N_1337,N_965,In_1430);
nand U1338 (N_1338,In_1905,N_51);
and U1339 (N_1339,N_177,In_2182);
or U1340 (N_1340,N_382,In_344);
xnor U1341 (N_1341,In_2534,N_420);
nor U1342 (N_1342,N_734,N_890);
nand U1343 (N_1343,In_725,N_195);
nand U1344 (N_1344,N_450,N_888);
nor U1345 (N_1345,In_1640,In_2204);
xnor U1346 (N_1346,N_12,N_332);
nand U1347 (N_1347,In_1440,In_2766);
or U1348 (N_1348,N_583,N_825);
xor U1349 (N_1349,N_852,N_1);
xnor U1350 (N_1350,N_761,N_89);
nor U1351 (N_1351,N_865,In_2543);
and U1352 (N_1352,In_1718,N_424);
nand U1353 (N_1353,N_17,N_817);
xnor U1354 (N_1354,N_231,N_269);
xor U1355 (N_1355,N_931,N_71);
nor U1356 (N_1356,N_189,N_573);
nand U1357 (N_1357,N_84,N_977);
or U1358 (N_1358,N_585,N_746);
xor U1359 (N_1359,N_166,In_741);
nor U1360 (N_1360,N_914,N_797);
or U1361 (N_1361,In_865,In_170);
and U1362 (N_1362,In_547,In_1994);
and U1363 (N_1363,N_972,In_945);
and U1364 (N_1364,N_807,In_474);
nand U1365 (N_1365,In_745,N_959);
and U1366 (N_1366,In_1731,In_1336);
or U1367 (N_1367,N_581,In_443);
nand U1368 (N_1368,In_2630,N_55);
or U1369 (N_1369,N_265,In_226);
and U1370 (N_1370,N_945,N_78);
and U1371 (N_1371,N_478,N_675);
or U1372 (N_1372,In_583,In_1869);
xnor U1373 (N_1373,In_2206,N_185);
and U1374 (N_1374,In_484,In_2579);
nor U1375 (N_1375,N_635,N_508);
xnor U1376 (N_1376,In_1255,In_264);
and U1377 (N_1377,In_814,N_574);
or U1378 (N_1378,In_2542,N_158);
xnor U1379 (N_1379,N_717,In_389);
nor U1380 (N_1380,In_1590,In_1447);
nand U1381 (N_1381,In_2257,N_333);
xor U1382 (N_1382,In_2645,In_710);
or U1383 (N_1383,In_696,In_2703);
and U1384 (N_1384,In_1805,In_2604);
nor U1385 (N_1385,N_443,N_330);
nor U1386 (N_1386,N_777,N_767);
nor U1387 (N_1387,N_221,N_948);
nand U1388 (N_1388,In_2724,In_1012);
or U1389 (N_1389,N_18,N_294);
and U1390 (N_1390,In_818,N_708);
nor U1391 (N_1391,N_295,N_827);
nor U1392 (N_1392,N_253,N_622);
nor U1393 (N_1393,In_949,N_4);
and U1394 (N_1394,In_2012,In_1329);
or U1395 (N_1395,N_756,N_173);
nor U1396 (N_1396,In_905,N_728);
and U1397 (N_1397,N_877,N_109);
xor U1398 (N_1398,In_2338,N_251);
nor U1399 (N_1399,In_1158,N_723);
nand U1400 (N_1400,N_532,In_735);
nand U1401 (N_1401,In_235,N_584);
xor U1402 (N_1402,N_886,In_1923);
nor U1403 (N_1403,In_1668,In_1713);
nor U1404 (N_1404,N_692,N_922);
nor U1405 (N_1405,N_239,N_365);
or U1406 (N_1406,N_393,N_349);
or U1407 (N_1407,In_1754,In_556);
and U1408 (N_1408,In_2749,N_334);
or U1409 (N_1409,N_831,In_1110);
or U1410 (N_1410,In_2401,N_156);
nand U1411 (N_1411,N_32,In_1774);
xnor U1412 (N_1412,N_511,In_835);
or U1413 (N_1413,In_1706,In_494);
nand U1414 (N_1414,N_597,In_2580);
nand U1415 (N_1415,N_139,N_356);
nor U1416 (N_1416,N_572,In_2017);
nand U1417 (N_1417,N_614,In_17);
xor U1418 (N_1418,In_890,N_447);
or U1419 (N_1419,N_556,In_378);
or U1420 (N_1420,In_634,N_748);
nor U1421 (N_1421,In_1645,In_1736);
or U1422 (N_1422,N_658,In_120);
xnor U1423 (N_1423,N_975,In_2917);
and U1424 (N_1424,In_1883,In_2742);
nor U1425 (N_1425,In_365,In_2489);
xnor U1426 (N_1426,In_574,N_368);
and U1427 (N_1427,N_515,N_241);
nand U1428 (N_1428,In_1835,N_908);
nand U1429 (N_1429,In_2328,In_1667);
or U1430 (N_1430,N_703,In_1453);
and U1431 (N_1431,In_1421,N_30);
and U1432 (N_1432,In_2586,N_455);
nor U1433 (N_1433,In_1823,N_710);
and U1434 (N_1434,In_808,N_864);
xnor U1435 (N_1435,In_703,In_434);
nor U1436 (N_1436,In_2555,N_274);
and U1437 (N_1437,N_47,N_621);
or U1438 (N_1438,In_1765,In_1623);
xor U1439 (N_1439,In_38,In_2266);
nand U1440 (N_1440,N_182,In_2699);
and U1441 (N_1441,N_735,In_1017);
or U1442 (N_1442,N_598,N_97);
nand U1443 (N_1443,In_2139,In_1147);
nor U1444 (N_1444,In_715,In_73);
xor U1445 (N_1445,N_796,In_209);
nand U1446 (N_1446,N_683,In_2439);
nand U1447 (N_1447,N_2,In_2727);
nand U1448 (N_1448,N_507,In_2475);
nor U1449 (N_1449,In_158,N_26);
xnor U1450 (N_1450,In_2409,N_329);
nand U1451 (N_1451,In_647,In_40);
or U1452 (N_1452,N_895,N_632);
nand U1453 (N_1453,N_804,N_126);
nand U1454 (N_1454,In_2621,N_387);
nand U1455 (N_1455,In_1140,In_1385);
and U1456 (N_1456,In_776,N_204);
or U1457 (N_1457,N_376,In_2283);
or U1458 (N_1458,In_161,N_808);
and U1459 (N_1459,N_492,N_79);
or U1460 (N_1460,In_661,In_2253);
nor U1461 (N_1461,N_962,In_1210);
nand U1462 (N_1462,In_156,N_278);
nor U1463 (N_1463,N_629,N_483);
xnor U1464 (N_1464,N_726,N_328);
nor U1465 (N_1465,N_856,N_762);
nor U1466 (N_1466,N_551,N_580);
nand U1467 (N_1467,In_2828,N_544);
nand U1468 (N_1468,In_763,In_733);
nor U1469 (N_1469,In_2595,In_2865);
or U1470 (N_1470,In_2863,N_103);
nor U1471 (N_1471,In_2775,In_109);
nor U1472 (N_1472,In_827,N_130);
nand U1473 (N_1473,N_513,N_198);
nor U1474 (N_1474,N_952,N_170);
nand U1475 (N_1475,In_1379,In_1166);
nor U1476 (N_1476,N_211,N_411);
or U1477 (N_1477,N_21,In_2436);
and U1478 (N_1478,N_179,N_839);
and U1479 (N_1479,N_686,In_789);
xnor U1480 (N_1480,In_220,N_729);
and U1481 (N_1481,In_1172,In_2063);
and U1482 (N_1482,N_678,In_173);
nand U1483 (N_1483,In_1435,In_2019);
nand U1484 (N_1484,In_2460,In_1741);
and U1485 (N_1485,In_1859,N_516);
nand U1486 (N_1486,N_153,In_569);
nand U1487 (N_1487,N_682,N_167);
and U1488 (N_1488,N_542,In_1220);
nand U1489 (N_1489,N_440,N_276);
and U1490 (N_1490,N_721,In_2228);
or U1491 (N_1491,In_653,N_697);
xnor U1492 (N_1492,In_995,In_928);
or U1493 (N_1493,In_69,N_901);
or U1494 (N_1494,In_2552,N_616);
nand U1495 (N_1495,N_957,N_685);
nand U1496 (N_1496,In_127,N_161);
and U1497 (N_1497,N_615,In_2303);
xor U1498 (N_1498,N_859,In_2548);
and U1499 (N_1499,N_290,In_1533);
or U1500 (N_1500,In_2427,In_1532);
and U1501 (N_1501,N_442,N_561);
xnor U1502 (N_1502,N_932,N_546);
nand U1503 (N_1503,N_456,In_2613);
or U1504 (N_1504,N_385,In_2318);
nor U1505 (N_1505,N_822,In_1543);
nand U1506 (N_1506,In_1014,In_1102);
nor U1507 (N_1507,In_1992,In_1350);
nor U1508 (N_1508,N_812,N_197);
and U1509 (N_1509,N_984,N_907);
nor U1510 (N_1510,In_1324,In_2817);
and U1511 (N_1511,N_428,In_1178);
nand U1512 (N_1512,N_57,N_813);
nor U1513 (N_1513,N_62,N_594);
nand U1514 (N_1514,N_327,N_375);
nor U1515 (N_1515,In_1768,In_2982);
and U1516 (N_1516,In_2818,N_91);
nand U1517 (N_1517,In_2053,In_2598);
and U1518 (N_1518,In_2119,In_868);
xor U1519 (N_1519,N_434,In_358);
or U1520 (N_1520,In_1920,N_346);
xnor U1521 (N_1521,N_792,In_386);
nor U1522 (N_1522,In_1558,N_514);
nor U1523 (N_1523,N_824,In_2879);
or U1524 (N_1524,In_2414,In_2174);
xor U1525 (N_1525,In_1308,N_64);
nand U1526 (N_1526,N_121,In_921);
xor U1527 (N_1527,In_2055,N_176);
or U1528 (N_1528,In_543,N_39);
xnor U1529 (N_1529,In_1627,N_885);
xor U1530 (N_1530,In_2208,In_2197);
or U1531 (N_1531,In_878,N_37);
nor U1532 (N_1532,N_955,N_159);
xnor U1533 (N_1533,N_33,In_1830);
and U1534 (N_1534,In_1303,In_2116);
and U1535 (N_1535,N_433,N_445);
and U1536 (N_1536,N_180,In_1757);
and U1537 (N_1537,N_560,N_823);
xor U1538 (N_1538,N_964,N_367);
nand U1539 (N_1539,N_784,N_293);
and U1540 (N_1540,In_163,In_580);
and U1541 (N_1541,N_395,In_2351);
xor U1542 (N_1542,In_2434,In_1632);
xor U1543 (N_1543,N_755,N_85);
or U1544 (N_1544,N_592,In_217);
and U1545 (N_1545,In_2498,In_2002);
or U1546 (N_1546,N_436,N_548);
or U1547 (N_1547,In_502,In_1454);
or U1548 (N_1548,In_1679,N_588);
and U1549 (N_1549,N_918,N_587);
xnor U1550 (N_1550,N_788,N_903);
xnor U1551 (N_1551,N_872,In_1957);
nor U1552 (N_1552,N_88,N_506);
or U1553 (N_1553,In_1133,In_1637);
and U1554 (N_1554,In_2569,In_1650);
nor U1555 (N_1555,In_1797,N_233);
nor U1556 (N_1556,In_2353,N_704);
or U1557 (N_1557,N_461,N_302);
or U1558 (N_1558,N_759,In_840);
and U1559 (N_1559,N_68,In_1838);
nor U1560 (N_1560,N_192,In_1591);
nand U1561 (N_1561,In_227,N_764);
nor U1562 (N_1562,N_558,In_1286);
or U1563 (N_1563,In_970,N_469);
nor U1564 (N_1564,N_23,In_796);
or U1565 (N_1565,In_2561,In_2803);
or U1566 (N_1566,N_342,In_2970);
nand U1567 (N_1567,N_900,N_245);
or U1568 (N_1568,N_537,In_2262);
nand U1569 (N_1569,In_215,N_634);
or U1570 (N_1570,In_74,N_15);
and U1571 (N_1571,In_307,N_816);
and U1572 (N_1572,In_993,In_135);
nor U1573 (N_1573,In_2664,N_794);
and U1574 (N_1574,In_2199,In_1652);
xnor U1575 (N_1575,In_2635,In_2077);
and U1576 (N_1576,N_711,In_824);
xnor U1577 (N_1577,In_664,In_2985);
nand U1578 (N_1578,N_380,N_535);
nor U1579 (N_1579,N_384,In_2388);
and U1580 (N_1580,In_561,In_1966);
and U1581 (N_1581,N_383,In_2088);
and U1582 (N_1582,N_814,N_476);
nor U1583 (N_1583,In_2128,In_1150);
or U1584 (N_1584,N_426,N_190);
or U1585 (N_1585,In_353,In_700);
and U1586 (N_1586,N_104,In_1372);
or U1587 (N_1587,In_1316,In_2849);
nand U1588 (N_1588,N_925,N_858);
xnor U1589 (N_1589,In_2064,In_317);
nor U1590 (N_1590,In_699,N_260);
or U1591 (N_1591,In_6,In_115);
nand U1592 (N_1592,N_985,In_2170);
nor U1593 (N_1593,In_726,N_93);
or U1594 (N_1594,In_243,In_2241);
and U1595 (N_1595,In_1451,N_899);
or U1596 (N_1596,N_910,In_356);
nand U1597 (N_1597,N_557,N_186);
or U1598 (N_1598,N_626,In_2356);
nand U1599 (N_1599,N_524,In_813);
or U1600 (N_1600,N_527,N_547);
nand U1601 (N_1601,N_128,In_1034);
nand U1602 (N_1602,In_191,N_414);
and U1603 (N_1603,In_2754,In_2612);
xor U1604 (N_1604,N_484,N_663);
and U1605 (N_1605,N_774,In_892);
xor U1606 (N_1606,N_967,N_929);
and U1607 (N_1607,N_249,In_1704);
nand U1608 (N_1608,N_41,N_59);
nand U1609 (N_1609,In_2870,In_347);
and U1610 (N_1610,N_500,N_44);
nand U1611 (N_1611,In_2392,In_1236);
or U1612 (N_1612,In_1129,In_175);
xnor U1613 (N_1613,In_331,N_636);
nor U1614 (N_1614,In_2851,In_1219);
nor U1615 (N_1615,In_1643,N_87);
xnor U1616 (N_1616,N_402,In_1717);
nor U1617 (N_1617,In_281,N_466);
nor U1618 (N_1618,N_904,In_1184);
nand U1619 (N_1619,N_915,N_270);
nor U1620 (N_1620,In_1538,In_1263);
or U1621 (N_1621,N_920,In_1500);
nor U1622 (N_1622,N_246,In_2618);
nand U1623 (N_1623,N_234,N_316);
or U1624 (N_1624,In_2739,N_465);
nor U1625 (N_1625,N_437,N_86);
or U1626 (N_1626,N_617,N_673);
and U1627 (N_1627,In_1960,N_778);
nor U1628 (N_1628,In_2041,In_572);
or U1629 (N_1629,N_521,N_619);
nor U1630 (N_1630,N_875,In_67);
nand U1631 (N_1631,N_438,In_22);
or U1632 (N_1632,N_45,N_377);
nand U1633 (N_1633,N_923,In_447);
or U1634 (N_1634,In_913,In_2808);
xnor U1635 (N_1635,N_713,N_291);
xor U1636 (N_1636,In_1136,In_2999);
xor U1637 (N_1637,In_1053,In_1832);
or U1638 (N_1638,N_474,N_607);
or U1639 (N_1639,N_555,N_927);
or U1640 (N_1640,N_565,In_536);
and U1641 (N_1641,In_2058,N_462);
or U1642 (N_1642,N_680,In_273);
or U1643 (N_1643,In_2014,In_132);
nor U1644 (N_1644,In_1094,N_149);
or U1645 (N_1645,In_1559,N_40);
nand U1646 (N_1646,N_491,In_2765);
nand U1647 (N_1647,N_210,N_122);
or U1648 (N_1648,In_1174,N_727);
and U1649 (N_1649,In_153,N_339);
nand U1650 (N_1650,In_1521,N_255);
nor U1651 (N_1651,N_851,N_207);
or U1652 (N_1652,N_802,In_1711);
xnor U1653 (N_1653,N_148,In_1753);
nand U1654 (N_1654,N_654,N_674);
xor U1655 (N_1655,In_1169,N_671);
nand U1656 (N_1656,N_963,In_164);
or U1657 (N_1657,In_503,In_1119);
and U1658 (N_1658,In_1295,In_1139);
nand U1659 (N_1659,N_217,N_112);
nand U1660 (N_1660,In_1143,In_2755);
xor U1661 (N_1661,N_640,In_1000);
nor U1662 (N_1662,N_458,N_571);
nand U1663 (N_1663,In_2186,In_2198);
xnor U1664 (N_1664,N_473,N_127);
nand U1665 (N_1665,N_38,N_54);
nor U1666 (N_1666,In_1611,N_289);
or U1667 (N_1667,N_277,N_282);
nor U1668 (N_1668,N_528,N_712);
xnor U1669 (N_1669,N_947,N_363);
xnor U1670 (N_1670,In_732,N_394);
and U1671 (N_1671,In_2090,In_2324);
xor U1672 (N_1672,N_228,In_2913);
and U1673 (N_1673,N_795,In_1397);
or U1674 (N_1674,N_613,N_919);
nor U1675 (N_1675,In_2175,In_2634);
or U1676 (N_1676,N_82,In_660);
xor U1677 (N_1677,In_213,N_218);
nand U1678 (N_1678,In_2596,N_638);
xnor U1679 (N_1679,In_1881,In_1564);
nor U1680 (N_1680,N_144,In_1398);
nor U1681 (N_1681,In_1545,N_205);
nor U1682 (N_1682,N_7,N_991);
or U1683 (N_1683,N_891,N_604);
xnor U1684 (N_1684,N_309,N_386);
and U1685 (N_1685,In_1517,N_489);
nor U1686 (N_1686,In_929,N_765);
or U1687 (N_1687,N_790,N_835);
xnor U1688 (N_1688,In_1769,In_1130);
xor U1689 (N_1689,N_162,In_2095);
nor U1690 (N_1690,N_838,N_301);
and U1691 (N_1691,N_216,N_772);
and U1692 (N_1692,In_2807,N_96);
and U1693 (N_1693,N_961,In_678);
and U1694 (N_1694,N_820,In_2114);
and U1695 (N_1695,N_313,In_1865);
or U1696 (N_1696,N_263,In_172);
and U1697 (N_1697,In_2124,In_417);
nor U1698 (N_1698,In_920,N_480);
or U1699 (N_1699,N_209,N_429);
nand U1700 (N_1700,In_2478,N_844);
and U1701 (N_1701,In_537,N_43);
or U1702 (N_1702,N_168,N_151);
nand U1703 (N_1703,N_928,N_523);
or U1704 (N_1704,In_1925,N_608);
xnor U1705 (N_1705,N_396,N_732);
nand U1706 (N_1706,N_408,In_1355);
nand U1707 (N_1707,In_632,In_2546);
xor U1708 (N_1708,N_562,N_486);
or U1709 (N_1709,In_589,In_538);
nor U1710 (N_1710,N_854,In_342);
or U1711 (N_1711,N_776,N_224);
or U1712 (N_1712,N_940,N_934);
or U1713 (N_1713,N_936,N_444);
xor U1714 (N_1714,N_35,In_1115);
xor U1715 (N_1715,In_1024,In_1927);
or U1716 (N_1716,N_193,N_336);
and U1717 (N_1717,In_328,N_586);
or U1718 (N_1718,N_751,In_988);
xor U1719 (N_1719,In_558,In_511);
or U1720 (N_1720,In_1254,In_1605);
nor U1721 (N_1721,N_655,N_311);
nand U1722 (N_1722,In_2024,N_326);
and U1723 (N_1723,N_871,In_2378);
or U1724 (N_1724,In_853,N_811);
or U1725 (N_1725,In_2942,N_741);
xnor U1726 (N_1726,In_2046,In_898);
xor U1727 (N_1727,In_197,N_842);
xnor U1728 (N_1728,N_911,In_885);
and U1729 (N_1729,N_988,N_202);
and U1730 (N_1730,In_392,N_398);
and U1731 (N_1731,N_392,N_481);
and U1732 (N_1732,In_339,In_581);
nand U1733 (N_1733,In_2583,In_2822);
and U1734 (N_1734,In_587,In_1560);
and U1735 (N_1735,N_742,In_2876);
nand U1736 (N_1736,In_352,In_3);
nor U1737 (N_1737,In_1027,N_833);
nand U1738 (N_1738,N_347,In_51);
nand U1739 (N_1739,N_691,In_301);
nand U1740 (N_1740,N_845,N_750);
xnor U1741 (N_1741,N_569,N_449);
nand U1742 (N_1742,In_1696,In_420);
nand U1743 (N_1743,In_2286,In_1954);
and U1744 (N_1744,N_787,N_421);
and U1745 (N_1745,In_1811,In_820);
and U1746 (N_1746,N_374,In_150);
nand U1747 (N_1747,In_520,In_483);
and U1748 (N_1748,In_1619,In_2511);
or U1749 (N_1749,N_135,N_510);
nor U1750 (N_1750,N_539,N_986);
and U1751 (N_1751,In_505,N_194);
xnor U1752 (N_1752,N_441,N_425);
and U1753 (N_1753,N_869,In_1436);
or U1754 (N_1754,In_2670,In_2102);
nand U1755 (N_1755,N_944,N_631);
and U1756 (N_1756,In_1098,In_1821);
and U1757 (N_1757,N_264,In_1228);
nor U1758 (N_1758,In_635,N_341);
nor U1759 (N_1759,In_2854,N_878);
xnor U1760 (N_1760,In_1162,In_542);
or U1761 (N_1761,In_2106,In_2082);
nor U1762 (N_1762,In_1616,In_1327);
nand U1763 (N_1763,N_296,In_2085);
nor U1764 (N_1764,In_1857,N_740);
xor U1765 (N_1765,In_2966,N_623);
nor U1766 (N_1766,N_477,N_882);
nand U1767 (N_1767,In_1168,In_658);
and U1768 (N_1768,N_533,In_2332);
xnor U1769 (N_1769,N_894,In_360);
xor U1770 (N_1770,N_553,N_470);
nand U1771 (N_1771,In_1523,N_687);
or U1772 (N_1772,In_2991,In_2248);
nor U1773 (N_1773,In_364,N_132);
xor U1774 (N_1774,N_137,In_2514);
xor U1775 (N_1775,In_2868,In_1985);
or U1776 (N_1776,In_2713,In_731);
nand U1777 (N_1777,N_630,In_597);
and U1778 (N_1778,N_248,In_2992);
xnor U1779 (N_1779,N_887,N_171);
xnor U1780 (N_1780,N_238,N_257);
nor U1781 (N_1781,In_2915,In_2515);
xnor U1782 (N_1782,In_2922,In_959);
xnor U1783 (N_1783,N_749,In_839);
nor U1784 (N_1784,In_2155,In_2211);
xnor U1785 (N_1785,N_129,In_1496);
or U1786 (N_1786,In_761,N_841);
or U1787 (N_1787,N_165,N_413);
nor U1788 (N_1788,N_279,In_2323);
xnor U1789 (N_1789,N_268,N_968);
and U1790 (N_1790,In_1393,N_589);
nand U1791 (N_1791,N_63,N_114);
nand U1792 (N_1792,N_350,N_801);
nor U1793 (N_1793,In_2850,N_979);
nand U1794 (N_1794,N_324,N_497);
and U1795 (N_1795,In_1574,N_690);
and U1796 (N_1796,In_0,In_2160);
xor U1797 (N_1797,N_618,In_1499);
xnor U1798 (N_1798,N_641,In_1727);
nand U1799 (N_1799,In_667,N_863);
or U1800 (N_1800,In_2864,N_323);
xnor U1801 (N_1801,N_321,In_2691);
and U1802 (N_1802,N_244,N_943);
and U1803 (N_1803,N_206,N_715);
and U1804 (N_1804,N_633,In_1671);
xor U1805 (N_1805,In_1068,In_1190);
and U1806 (N_1806,In_2098,N_369);
or U1807 (N_1807,In_249,In_883);
or U1808 (N_1808,N_657,In_428);
and U1809 (N_1809,N_125,In_1863);
nor U1810 (N_1810,In_847,In_335);
or U1811 (N_1811,N_435,In_1621);
or U1812 (N_1812,N_983,In_2563);
nand U1813 (N_1813,In_2115,In_1205);
xor U1814 (N_1814,In_2377,In_2947);
or U1815 (N_1815,N_448,N_744);
or U1816 (N_1816,In_2022,In_2794);
nor U1817 (N_1817,N_736,N_284);
nor U1818 (N_1818,In_2322,In_2235);
nor U1819 (N_1819,In_669,In_2687);
or U1820 (N_1820,N_660,N_11);
nand U1821 (N_1821,N_563,In_2330);
or U1822 (N_1822,In_1191,N_938);
and U1823 (N_1823,N_722,N_298);
and U1824 (N_1824,N_974,N_620);
and U1825 (N_1825,N_67,N_873);
nor U1826 (N_1826,N_624,In_2231);
xor U1827 (N_1827,In_1485,N_840);
xnor U1828 (N_1828,In_1392,In_315);
nor U1829 (N_1829,N_933,N_488);
xor U1830 (N_1830,N_538,N_668);
or U1831 (N_1831,In_1732,In_276);
and U1832 (N_1832,N_174,N_775);
xor U1833 (N_1833,In_1429,N_670);
xor U1834 (N_1834,In_470,N_937);
and U1835 (N_1835,In_2551,N_106);
nor U1836 (N_1836,N_861,In_2226);
nor U1837 (N_1837,N_199,N_76);
xor U1838 (N_1838,N_810,N_225);
xnor U1839 (N_1839,N_610,In_1100);
or U1840 (N_1840,In_258,N_157);
and U1841 (N_1841,N_954,N_577);
and U1842 (N_1842,N_297,In_2793);
and U1843 (N_1843,N_643,N_317);
nor U1844 (N_1844,N_212,In_1208);
nor U1845 (N_1845,N_75,In_779);
or U1846 (N_1846,In_451,In_1471);
nand U1847 (N_1847,In_89,N_912);
nand U1848 (N_1848,N_649,In_1248);
and U1849 (N_1849,In_185,In_996);
nand U1850 (N_1850,In_2150,In_1221);
nand U1851 (N_1851,In_2239,N_446);
nand U1852 (N_1852,N_602,In_2218);
xor U1853 (N_1853,In_1093,In_1572);
nor U1854 (N_1854,N_8,In_800);
and U1855 (N_1855,N_806,N_645);
or U1856 (N_1856,In_2070,N_853);
xor U1857 (N_1857,In_129,In_836);
and U1858 (N_1858,In_2133,N_490);
xnor U1859 (N_1859,In_2916,N_870);
or U1860 (N_1860,In_493,In_623);
or U1861 (N_1861,N_611,N_780);
and U1862 (N_1862,N_271,In_2210);
nand U1863 (N_1863,In_1798,In_659);
and U1864 (N_1864,N_625,N_779);
or U1865 (N_1865,N_950,In_141);
xnor U1866 (N_1866,N_123,N_292);
nand U1867 (N_1867,In_1837,N_20);
nand U1868 (N_1868,In_1359,In_730);
nor U1869 (N_1869,N_676,N_662);
nand U1870 (N_1870,In_1108,In_82);
xnor U1871 (N_1871,In_910,N_627);
and U1872 (N_1872,N_73,In_2277);
xnor U1873 (N_1873,N_665,In_2030);
and U1874 (N_1874,In_1419,In_2832);
nand U1875 (N_1875,N_65,N_340);
or U1876 (N_1876,In_1735,N_305);
nand U1877 (N_1877,In_1503,N_836);
or U1878 (N_1878,In_1595,N_582);
or U1879 (N_1879,In_179,N_898);
xnor U1880 (N_1880,In_2530,N_763);
or U1881 (N_1881,N_953,In_2165);
nor U1882 (N_1882,In_403,N_272);
or U1883 (N_1883,In_2185,In_2764);
nand U1884 (N_1884,In_1358,In_515);
xnor U1885 (N_1885,In_590,In_2007);
and U1886 (N_1886,In_340,In_514);
or U1887 (N_1887,N_479,N_344);
nand U1888 (N_1888,In_1373,N_52);
and U1889 (N_1889,N_966,In_2347);
or U1890 (N_1890,N_378,N_809);
xor U1891 (N_1891,In_2004,N_230);
and U1892 (N_1892,N_343,In_1515);
xnor U1893 (N_1893,In_2426,In_2977);
nand U1894 (N_1894,In_1770,N_720);
nor U1895 (N_1895,N_261,N_287);
xor U1896 (N_1896,In_787,In_2910);
nand U1897 (N_1897,In_529,N_117);
xor U1898 (N_1898,In_1029,In_843);
nand U1899 (N_1899,N_707,In_1709);
or U1900 (N_1900,In_1280,In_901);
nand U1901 (N_1901,In_2036,N_590);
nor U1902 (N_1902,In_680,In_592);
and U1903 (N_1903,N_698,N_401);
xor U1904 (N_1904,In_1084,N_517);
or U1905 (N_1905,In_1251,N_360);
or U1906 (N_1906,In_1378,In_2342);
or U1907 (N_1907,N_250,N_138);
and U1908 (N_1908,N_501,In_19);
xnor U1909 (N_1909,N_273,N_956);
nor U1910 (N_1910,N_978,N_689);
and U1911 (N_1911,N_5,N_335);
or U1912 (N_1912,N_415,In_2482);
nor U1913 (N_1913,N_215,In_1664);
or U1914 (N_1914,In_1780,In_1494);
or U1915 (N_1915,In_441,In_1474);
nand U1916 (N_1916,In_1833,N_338);
and U1917 (N_1917,N_552,In_34);
and U1918 (N_1918,N_706,In_1065);
nand U1919 (N_1919,N_77,N_677);
nor U1920 (N_1920,In_603,N_612);
or U1921 (N_1921,N_738,In_1492);
nor U1922 (N_1922,In_2805,In_1306);
and U1923 (N_1923,N_299,In_1556);
and U1924 (N_1924,N_829,N_3);
xnor U1925 (N_1925,N_353,N_417);
nand U1926 (N_1926,N_331,In_545);
xor U1927 (N_1927,N_459,In_2304);
nor U1928 (N_1928,In_2857,In_1123);
nand U1929 (N_1929,In_2138,N_419);
nor U1930 (N_1930,N_381,In_1269);
nand U1931 (N_1931,In_2467,N_799);
nor U1932 (N_1932,In_1064,In_2361);
nor U1933 (N_1933,In_1675,N_99);
xor U1934 (N_1934,N_993,N_308);
nor U1935 (N_1935,N_644,In_1973);
nor U1936 (N_1936,N_463,N_880);
and U1937 (N_1937,In_195,N_306);
or U1938 (N_1938,In_2559,N_874);
and U1939 (N_1939,N_358,In_2993);
or U1940 (N_1940,N_430,N_701);
xor U1941 (N_1941,In_2738,N_990);
xor U1942 (N_1942,In_1878,In_830);
or U1943 (N_1943,In_396,In_1684);
or U1944 (N_1944,N_760,N_716);
nor U1945 (N_1945,In_4,In_460);
nor U1946 (N_1946,In_190,In_1194);
and U1947 (N_1947,N_725,N_884);
or U1948 (N_1948,In_2360,In_701);
nand U1949 (N_1949,In_1982,N_9);
or U1950 (N_1950,In_767,In_1792);
and U1951 (N_1951,In_2995,In_98);
nand U1952 (N_1952,In_1493,In_1439);
nand U1953 (N_1953,In_2365,N_848);
and U1954 (N_1954,N_798,N_653);
nand U1955 (N_1955,N_576,In_2391);
or U1956 (N_1956,N_432,In_1124);
xor U1957 (N_1957,N_579,N_146);
and U1958 (N_1958,In_274,N_849);
nor U1959 (N_1959,N_996,N_803);
nand U1960 (N_1960,In_1371,N_403);
nand U1961 (N_1961,N_926,In_2735);
nor U1962 (N_1962,N_601,N_267);
xnor U1963 (N_1963,N_163,In_1111);
nor U1964 (N_1964,In_2668,N_213);
or U1965 (N_1965,In_979,N_92);
or U1966 (N_1966,In_1953,N_227);
and U1967 (N_1967,N_229,In_2369);
nor U1968 (N_1968,In_2140,In_1362);
xnor U1969 (N_1969,N_942,N_639);
and U1970 (N_1970,In_23,N_834);
xor U1971 (N_1971,In_1631,N_664);
nor U1972 (N_1972,N_924,In_1387);
nand U1973 (N_1973,N_371,N_549);
xnor U1974 (N_1974,N_351,N_83);
and U1975 (N_1975,In_2547,N_405);
or U1976 (N_1976,In_485,In_2686);
xor U1977 (N_1977,N_178,N_567);
nand U1978 (N_1978,N_902,N_821);
xnor U1979 (N_1979,N_345,N_679);
or U1980 (N_1980,N_781,N_850);
nand U1981 (N_1981,In_2059,N_42);
xor U1982 (N_1982,In_1900,N_525);
or U1983 (N_1983,In_2572,In_1799);
nor U1984 (N_1984,In_2129,N_534);
nor U1985 (N_1985,In_1322,In_2120);
nor U1986 (N_1986,N_46,In_1991);
nor U1987 (N_1987,N_285,In_1963);
xor U1988 (N_1988,N_155,N_24);
xnor U1989 (N_1989,In_1810,In_1723);
and U1990 (N_1990,In_2761,In_1747);
or U1991 (N_1991,In_491,N_642);
nor U1992 (N_1992,N_6,N_499);
nand U1993 (N_1993,N_599,In_2659);
xor U1994 (N_1994,In_2575,N_520);
xnor U1995 (N_1995,In_2829,In_2809);
nand U1996 (N_1996,N_322,N_512);
nand U1997 (N_1997,In_2524,N_366);
or U1998 (N_1998,In_2653,N_312);
nand U1999 (N_1999,N_519,N_319);
and U2000 (N_2000,N_1688,N_1626);
and U2001 (N_2001,N_1085,N_1064);
and U2002 (N_2002,N_1969,N_1202);
or U2003 (N_2003,N_1765,N_1229);
or U2004 (N_2004,N_1813,N_1574);
and U2005 (N_2005,N_1863,N_1750);
and U2006 (N_2006,N_1705,N_1590);
nor U2007 (N_2007,N_1474,N_1310);
and U2008 (N_2008,N_1281,N_1510);
nor U2009 (N_2009,N_1149,N_1161);
or U2010 (N_2010,N_1137,N_1562);
nor U2011 (N_2011,N_1177,N_1207);
and U2012 (N_2012,N_1026,N_1854);
nor U2013 (N_2013,N_1067,N_1054);
xnor U2014 (N_2014,N_1571,N_1350);
xnor U2015 (N_2015,N_1829,N_1358);
or U2016 (N_2016,N_1919,N_1640);
nor U2017 (N_2017,N_1236,N_1980);
nor U2018 (N_2018,N_1498,N_1699);
nand U2019 (N_2019,N_1484,N_1698);
and U2020 (N_2020,N_1951,N_1463);
nand U2021 (N_2021,N_1872,N_1645);
or U2022 (N_2022,N_1860,N_1652);
nand U2023 (N_2023,N_1375,N_1097);
nor U2024 (N_2024,N_1136,N_1904);
xnor U2025 (N_2025,N_1703,N_1925);
nand U2026 (N_2026,N_1158,N_1719);
nor U2027 (N_2027,N_1630,N_1106);
nand U2028 (N_2028,N_1727,N_1240);
or U2029 (N_2029,N_1857,N_1805);
or U2030 (N_2030,N_1117,N_1101);
nand U2031 (N_2031,N_1366,N_1609);
or U2032 (N_2032,N_1217,N_1776);
nor U2033 (N_2033,N_1532,N_1173);
or U2034 (N_2034,N_1911,N_1183);
nand U2035 (N_2035,N_1514,N_1086);
nand U2036 (N_2036,N_1282,N_1460);
and U2037 (N_2037,N_1603,N_1915);
or U2038 (N_2038,N_1267,N_1455);
and U2039 (N_2039,N_1615,N_1050);
nor U2040 (N_2040,N_1743,N_1305);
and U2041 (N_2041,N_1480,N_1001);
or U2042 (N_2042,N_1777,N_1081);
nand U2043 (N_2043,N_1008,N_1492);
or U2044 (N_2044,N_1541,N_1686);
nor U2045 (N_2045,N_1682,N_1493);
and U2046 (N_2046,N_1581,N_1570);
nand U2047 (N_2047,N_1822,N_1428);
or U2048 (N_2048,N_1667,N_1669);
xnor U2049 (N_2049,N_1212,N_1658);
or U2050 (N_2050,N_1759,N_1839);
or U2051 (N_2051,N_1304,N_1948);
and U2052 (N_2052,N_1663,N_1327);
nand U2053 (N_2053,N_1808,N_1594);
xor U2054 (N_2054,N_1061,N_1836);
nor U2055 (N_2055,N_1687,N_1632);
or U2056 (N_2056,N_1924,N_1223);
or U2057 (N_2057,N_1019,N_1251);
and U2058 (N_2058,N_1280,N_1079);
nand U2059 (N_2059,N_1968,N_1410);
or U2060 (N_2060,N_1192,N_1336);
xnor U2061 (N_2061,N_1981,N_1057);
nand U2062 (N_2062,N_1732,N_1725);
nor U2063 (N_2063,N_1031,N_1185);
nor U2064 (N_2064,N_1602,N_1296);
or U2065 (N_2065,N_1317,N_1029);
or U2066 (N_2066,N_1695,N_1913);
nor U2067 (N_2067,N_1840,N_1881);
nand U2068 (N_2068,N_1436,N_1341);
nor U2069 (N_2069,N_1735,N_1868);
nor U2070 (N_2070,N_1819,N_1773);
nand U2071 (N_2071,N_1423,N_1340);
or U2072 (N_2072,N_1367,N_1575);
nand U2073 (N_2073,N_1254,N_1309);
and U2074 (N_2074,N_1523,N_1264);
or U2075 (N_2075,N_1262,N_1553);
or U2076 (N_2076,N_1165,N_1121);
and U2077 (N_2077,N_1994,N_1613);
xor U2078 (N_2078,N_1119,N_1102);
and U2079 (N_2079,N_1406,N_1563);
nor U2080 (N_2080,N_1397,N_1027);
nor U2081 (N_2081,N_1799,N_1148);
or U2082 (N_2082,N_1661,N_1517);
or U2083 (N_2083,N_1960,N_1634);
and U2084 (N_2084,N_1627,N_1814);
and U2085 (N_2085,N_1780,N_1036);
nor U2086 (N_2086,N_1434,N_1624);
xor U2087 (N_2087,N_1831,N_1935);
and U2088 (N_2088,N_1611,N_1761);
nor U2089 (N_2089,N_1507,N_1692);
or U2090 (N_2090,N_1095,N_1084);
or U2091 (N_2091,N_1501,N_1905);
nor U2092 (N_2092,N_1748,N_1017);
nand U2093 (N_2093,N_1832,N_1151);
nor U2094 (N_2094,N_1790,N_1343);
nand U2095 (N_2095,N_1300,N_1355);
xor U2096 (N_2096,N_1647,N_1762);
nor U2097 (N_2097,N_1852,N_1697);
xnor U2098 (N_2098,N_1944,N_1153);
or U2099 (N_2099,N_1565,N_1864);
xnor U2100 (N_2100,N_1513,N_1014);
nor U2101 (N_2101,N_1522,N_1099);
nor U2102 (N_2102,N_1299,N_1239);
nand U2103 (N_2103,N_1897,N_1564);
nor U2104 (N_2104,N_1978,N_1483);
and U2105 (N_2105,N_1542,N_1593);
nor U2106 (N_2106,N_1015,N_1134);
nor U2107 (N_2107,N_1672,N_1823);
and U2108 (N_2108,N_1867,N_1975);
or U2109 (N_2109,N_1400,N_1856);
or U2110 (N_2110,N_1616,N_1444);
nand U2111 (N_2111,N_1419,N_1895);
or U2112 (N_2112,N_1744,N_1368);
and U2113 (N_2113,N_1936,N_1511);
and U2114 (N_2114,N_1345,N_1416);
nor U2115 (N_2115,N_1037,N_1006);
xnor U2116 (N_2116,N_1549,N_1046);
xnor U2117 (N_2117,N_1092,N_1926);
or U2118 (N_2118,N_1076,N_1133);
or U2119 (N_2119,N_1087,N_1472);
and U2120 (N_2120,N_1821,N_1107);
or U2121 (N_2121,N_1784,N_1963);
nor U2122 (N_2122,N_1620,N_1409);
xor U2123 (N_2123,N_1909,N_1861);
nand U2124 (N_2124,N_1334,N_1930);
and U2125 (N_2125,N_1786,N_1302);
nand U2126 (N_2126,N_1668,N_1722);
or U2127 (N_2127,N_1204,N_1674);
nor U2128 (N_2128,N_1740,N_1866);
nand U2129 (N_2129,N_1934,N_1998);
xnor U2130 (N_2130,N_1422,N_1398);
nand U2131 (N_2131,N_1335,N_1118);
nand U2132 (N_2132,N_1458,N_1918);
nand U2133 (N_2133,N_1530,N_1521);
nand U2134 (N_2134,N_1074,N_1432);
nand U2135 (N_2135,N_1502,N_1643);
and U2136 (N_2136,N_1670,N_1657);
nand U2137 (N_2137,N_1536,N_1021);
xor U2138 (N_2138,N_1869,N_1371);
and U2139 (N_2139,N_1795,N_1883);
or U2140 (N_2140,N_1465,N_1892);
xnor U2141 (N_2141,N_1506,N_1965);
nor U2142 (N_2142,N_1195,N_1120);
and U2143 (N_2143,N_1733,N_1078);
nor U2144 (N_2144,N_1701,N_1199);
xnor U2145 (N_2145,N_1424,N_1045);
nor U2146 (N_2146,N_1516,N_1982);
nand U2147 (N_2147,N_1189,N_1273);
or U2148 (N_2148,N_1587,N_1617);
xor U2149 (N_2149,N_1798,N_1105);
nand U2150 (N_2150,N_1504,N_1171);
nor U2151 (N_2151,N_1443,N_1650);
or U2152 (N_2152,N_1253,N_1421);
xor U2153 (N_2153,N_1131,N_1162);
nand U2154 (N_2154,N_1788,N_1793);
nor U2155 (N_2155,N_1741,N_1351);
nor U2156 (N_2156,N_1680,N_1870);
nor U2157 (N_2157,N_1537,N_1604);
nor U2158 (N_2158,N_1629,N_1454);
nor U2159 (N_2159,N_1804,N_1755);
or U2160 (N_2160,N_1572,N_1241);
xnor U2161 (N_2161,N_1734,N_1349);
or U2162 (N_2162,N_1952,N_1714);
or U2163 (N_2163,N_1708,N_1942);
xor U2164 (N_2164,N_1266,N_1344);
xnor U2165 (N_2165,N_1842,N_1882);
nor U2166 (N_2166,N_1292,N_1724);
xnor U2167 (N_2167,N_1450,N_1124);
or U2168 (N_2168,N_1083,N_1539);
xnor U2169 (N_2169,N_1082,N_1383);
or U2170 (N_2170,N_1828,N_1515);
nand U2171 (N_2171,N_1216,N_1311);
nor U2172 (N_2172,N_1880,N_1704);
xor U2173 (N_2173,N_1338,N_1332);
nor U2174 (N_2174,N_1983,N_1122);
and U2175 (N_2175,N_1374,N_1172);
nand U2176 (N_2176,N_1638,N_1258);
nor U2177 (N_2177,N_1841,N_1113);
and U2178 (N_2178,N_1816,N_1751);
xor U2179 (N_2179,N_1903,N_1991);
and U2180 (N_2180,N_1677,N_1614);
and U2181 (N_2181,N_1032,N_1114);
nor U2182 (N_2182,N_1048,N_1625);
xnor U2183 (N_2183,N_1269,N_1276);
or U2184 (N_2184,N_1939,N_1633);
nand U2185 (N_2185,N_1025,N_1268);
nor U2186 (N_2186,N_1376,N_1294);
xnor U2187 (N_2187,N_1414,N_1660);
nand U2188 (N_2188,N_1945,N_1599);
and U2189 (N_2189,N_1946,N_1543);
and U2190 (N_2190,N_1691,N_1033);
or U2191 (N_2191,N_1024,N_1179);
nor U2192 (N_2192,N_1073,N_1957);
nand U2193 (N_2193,N_1291,N_1979);
nand U2194 (N_2194,N_1089,N_1578);
nand U2195 (N_2195,N_1226,N_1846);
and U2196 (N_2196,N_1737,N_1713);
nor U2197 (N_2197,N_1221,N_1785);
nand U2198 (N_2198,N_1360,N_1038);
nand U2199 (N_2199,N_1175,N_1288);
or U2200 (N_2200,N_1491,N_1495);
xor U2201 (N_2201,N_1348,N_1147);
or U2202 (N_2202,N_1301,N_1889);
nand U2203 (N_2203,N_1481,N_1684);
xor U2204 (N_2204,N_1250,N_1205);
nand U2205 (N_2205,N_1853,N_1290);
and U2206 (N_2206,N_1916,N_1265);
or U2207 (N_2207,N_1818,N_1597);
xnor U2208 (N_2208,N_1094,N_1555);
or U2209 (N_2209,N_1768,N_1219);
xnor U2210 (N_2210,N_1896,N_1005);
or U2211 (N_2211,N_1844,N_1128);
nand U2212 (N_2212,N_1203,N_1649);
xor U2213 (N_2213,N_1170,N_1448);
nor U2214 (N_2214,N_1156,N_1888);
xnor U2215 (N_2215,N_1929,N_1509);
nor U2216 (N_2216,N_1865,N_1452);
nand U2217 (N_2217,N_1987,N_1508);
nand U2218 (N_2218,N_1244,N_1091);
and U2219 (N_2219,N_1096,N_1791);
or U2220 (N_2220,N_1373,N_1583);
or U2221 (N_2221,N_1407,N_1585);
or U2222 (N_2222,N_1020,N_1835);
xnor U2223 (N_2223,N_1731,N_1286);
and U2224 (N_2224,N_1742,N_1874);
and U2225 (N_2225,N_1811,N_1088);
or U2226 (N_2226,N_1546,N_1186);
or U2227 (N_2227,N_1004,N_1993);
or U2228 (N_2228,N_1477,N_1456);
and U2229 (N_2229,N_1182,N_1641);
nand U2230 (N_2230,N_1190,N_1132);
or U2231 (N_2231,N_1586,N_1110);
xor U2232 (N_2232,N_1573,N_1441);
or U2233 (N_2233,N_1550,N_1312);
nor U2234 (N_2234,N_1275,N_1797);
xnor U2235 (N_2235,N_1591,N_1430);
nand U2236 (N_2236,N_1928,N_1330);
or U2237 (N_2237,N_1858,N_1601);
nand U2238 (N_2238,N_1496,N_1547);
and U2239 (N_2239,N_1779,N_1706);
or U2240 (N_2240,N_1451,N_1529);
nand U2241 (N_2241,N_1966,N_1063);
and U2242 (N_2242,N_1125,N_1577);
nor U2243 (N_2243,N_1721,N_1908);
nor U2244 (N_2244,N_1610,N_1464);
and U2245 (N_2245,N_1770,N_1446);
or U2246 (N_2246,N_1940,N_1753);
xnor U2247 (N_2247,N_1035,N_1736);
nand U2248 (N_2248,N_1461,N_1651);
xnor U2249 (N_2249,N_1363,N_1738);
xnor U2250 (N_2250,N_1769,N_1758);
nor U2251 (N_2251,N_1700,N_1243);
xnor U2252 (N_2252,N_1702,N_1922);
nand U2253 (N_2253,N_1920,N_1152);
and U2254 (N_2254,N_1249,N_1320);
xnor U2255 (N_2255,N_1628,N_1447);
and U2256 (N_2256,N_1220,N_1385);
xor U2257 (N_2257,N_1115,N_1833);
nand U2258 (N_2258,N_1069,N_1381);
or U2259 (N_2259,N_1062,N_1248);
and U2260 (N_2260,N_1028,N_1557);
xnor U2261 (N_2261,N_1453,N_1402);
xor U2262 (N_2262,N_1353,N_1990);
and U2263 (N_2263,N_1678,N_1943);
or U2264 (N_2264,N_1298,N_1815);
or U2265 (N_2265,N_1431,N_1181);
nand U2266 (N_2266,N_1228,N_1321);
nand U2267 (N_2267,N_1016,N_1756);
or U2268 (N_2268,N_1080,N_1246);
xnor U2269 (N_2269,N_1955,N_1060);
or U2270 (N_2270,N_1612,N_1512);
xnor U2271 (N_2271,N_1885,N_1075);
nor U2272 (N_2272,N_1065,N_1098);
nand U2273 (N_2273,N_1323,N_1261);
and U2274 (N_2274,N_1961,N_1285);
nand U2275 (N_2275,N_1138,N_1307);
nor U2276 (N_2276,N_1973,N_1850);
xor U2277 (N_2277,N_1986,N_1426);
or U2278 (N_2278,N_1425,N_1322);
or U2279 (N_2279,N_1792,N_1230);
xnor U2280 (N_2280,N_1690,N_1435);
nand U2281 (N_2281,N_1442,N_1372);
nand U2282 (N_2282,N_1995,N_1168);
nor U2283 (N_2283,N_1242,N_1820);
and U2284 (N_2284,N_1654,N_1503);
or U2285 (N_2285,N_1396,N_1342);
nand U2286 (N_2286,N_1287,N_1675);
nand U2287 (N_2287,N_1794,N_1346);
nand U2288 (N_2288,N_1324,N_1109);
nand U2289 (N_2289,N_1568,N_1490);
or U2290 (N_2290,N_1333,N_1252);
xor U2291 (N_2291,N_1775,N_1146);
nand U2292 (N_2292,N_1938,N_1497);
nor U2293 (N_2293,N_1639,N_1764);
nor U2294 (N_2294,N_1042,N_1723);
or U2295 (N_2295,N_1193,N_1475);
nor U2296 (N_2296,N_1696,N_1313);
or U2297 (N_2297,N_1685,N_1274);
nor U2298 (N_2298,N_1235,N_1715);
nor U2299 (N_2299,N_1720,N_1540);
nand U2300 (N_2300,N_1745,N_1757);
or U2301 (N_2301,N_1160,N_1142);
nand U2302 (N_2302,N_1917,N_1180);
and U2303 (N_2303,N_1412,N_1257);
xor U2304 (N_2304,N_1711,N_1213);
nand U2305 (N_2305,N_1052,N_1459);
or U2306 (N_2306,N_1824,N_1356);
nand U2307 (N_2307,N_1393,N_1135);
xnor U2308 (N_2308,N_1893,N_1462);
and U2309 (N_2309,N_1314,N_1891);
or U2310 (N_2310,N_1278,N_1429);
and U2311 (N_2311,N_1681,N_1002);
nand U2312 (N_2312,N_1145,N_1093);
xor U2313 (N_2313,N_1653,N_1914);
and U2314 (N_2314,N_1116,N_1972);
nand U2315 (N_2315,N_1174,N_1782);
or U2316 (N_2316,N_1947,N_1659);
or U2317 (N_2317,N_1066,N_1988);
and U2318 (N_2318,N_1316,N_1921);
and U2319 (N_2319,N_1655,N_1469);
and U2320 (N_2320,N_1848,N_1403);
and U2321 (N_2321,N_1884,N_1315);
and U2322 (N_2322,N_1379,N_1646);
nor U2323 (N_2323,N_1387,N_1352);
nor U2324 (N_2324,N_1068,N_1297);
xnor U2325 (N_2325,N_1992,N_1150);
nor U2326 (N_2326,N_1642,N_1862);
xnor U2327 (N_2327,N_1598,N_1439);
xnor U2328 (N_2328,N_1072,N_1637);
or U2329 (N_2329,N_1875,N_1392);
nand U2330 (N_2330,N_1225,N_1879);
or U2331 (N_2331,N_1796,N_1802);
xor U2332 (N_2332,N_1801,N_1807);
or U2333 (N_2333,N_1218,N_1906);
and U2334 (N_2334,N_1817,N_1962);
nor U2335 (N_2335,N_1887,N_1279);
xnor U2336 (N_2336,N_1932,N_1662);
nor U2337 (N_2337,N_1886,N_1717);
nor U2338 (N_2338,N_1364,N_1144);
and U2339 (N_2339,N_1010,N_1104);
nor U2340 (N_2340,N_1608,N_1956);
and U2341 (N_2341,N_1766,N_1718);
xnor U2342 (N_2342,N_1184,N_1295);
nor U2343 (N_2343,N_1210,N_1789);
and U2344 (N_2344,N_1056,N_1198);
nand U2345 (N_2345,N_1528,N_1030);
nor U2346 (N_2346,N_1760,N_1605);
and U2347 (N_2347,N_1912,N_1534);
nand U2348 (N_2348,N_1233,N_1487);
and U2349 (N_2349,N_1810,N_1747);
xnor U2350 (N_2350,N_1022,N_1194);
xor U2351 (N_2351,N_1482,N_1976);
xor U2352 (N_2352,N_1166,N_1231);
nand U2353 (N_2353,N_1763,N_1197);
nand U2354 (N_2354,N_1538,N_1644);
xnor U2355 (N_2355,N_1825,N_1548);
nand U2356 (N_2356,N_1806,N_1059);
or U2357 (N_2357,N_1673,N_1556);
xor U2358 (N_2358,N_1671,N_1389);
nand U2359 (N_2359,N_1479,N_1354);
nand U2360 (N_2360,N_1103,N_1716);
nor U2361 (N_2361,N_1582,N_1489);
xor U2362 (N_2362,N_1964,N_1533);
xnor U2363 (N_2363,N_1471,N_1413);
xor U2364 (N_2364,N_1712,N_1812);
nor U2365 (N_2365,N_1211,N_1576);
xor U2366 (N_2366,N_1800,N_1559);
nor U2367 (N_2367,N_1749,N_1247);
xor U2368 (N_2368,N_1362,N_1418);
and U2369 (N_2369,N_1803,N_1849);
nor U2370 (N_2370,N_1159,N_1989);
nand U2371 (N_2371,N_1224,N_1283);
or U2372 (N_2372,N_1200,N_1531);
nor U2373 (N_2373,N_1551,N_1129);
nor U2374 (N_2374,N_1877,N_1873);
xnor U2375 (N_2375,N_1683,N_1237);
nor U2376 (N_2376,N_1847,N_1664);
and U2377 (N_2377,N_1837,N_1208);
and U2378 (N_2378,N_1622,N_1545);
or U2379 (N_2379,N_1589,N_1592);
xor U2380 (N_2380,N_1380,N_1826);
and U2381 (N_2381,N_1141,N_1227);
and U2382 (N_2382,N_1126,N_1289);
xnor U2383 (N_2383,N_1827,N_1927);
and U2384 (N_2384,N_1438,N_1427);
nor U2385 (N_2385,N_1369,N_1359);
xnor U2386 (N_2386,N_1325,N_1729);
nand U2387 (N_2387,N_1433,N_1855);
and U2388 (N_2388,N_1178,N_1499);
or U2389 (N_2389,N_1730,N_1377);
xnor U2390 (N_2390,N_1752,N_1967);
nand U2391 (N_2391,N_1127,N_1579);
nor U2392 (N_2392,N_1898,N_1399);
and U2393 (N_2393,N_1209,N_1196);
nor U2394 (N_2394,N_1485,N_1476);
xnor U2395 (N_2395,N_1746,N_1143);
and U2396 (N_2396,N_1596,N_1588);
xor U2397 (N_2397,N_1486,N_1552);
nor U2398 (N_2398,N_1473,N_1958);
and U2399 (N_2399,N_1636,N_1970);
nor U2400 (N_2400,N_1417,N_1384);
nor U2401 (N_2401,N_1023,N_1329);
or U2402 (N_2402,N_1923,N_1910);
nand U2403 (N_2403,N_1974,N_1238);
nand U2404 (N_2404,N_1679,N_1271);
and U2405 (N_2405,N_1370,N_1191);
or U2406 (N_2406,N_1259,N_1007);
and U2407 (N_2407,N_1018,N_1255);
nor U2408 (N_2408,N_1566,N_1984);
or U2409 (N_2409,N_1053,N_1838);
or U2410 (N_2410,N_1306,N_1772);
and U2411 (N_2411,N_1404,N_1580);
or U2412 (N_2412,N_1871,N_1937);
and U2413 (N_2413,N_1043,N_1996);
nand U2414 (N_2414,N_1739,N_1710);
and U2415 (N_2415,N_1058,N_1234);
or U2416 (N_2416,N_1277,N_1676);
and U2417 (N_2417,N_1326,N_1470);
or U2418 (N_2418,N_1999,N_1318);
or U2419 (N_2419,N_1112,N_1843);
nand U2420 (N_2420,N_1055,N_1378);
nor U2421 (N_2421,N_1090,N_1584);
nand U2422 (N_2422,N_1188,N_1631);
or U2423 (N_2423,N_1395,N_1270);
nand U2424 (N_2424,N_1411,N_1011);
nor U2425 (N_2425,N_1420,N_1977);
nor U2426 (N_2426,N_1890,N_1394);
nor U2427 (N_2427,N_1365,N_1830);
nand U2428 (N_2428,N_1051,N_1505);
nand U2429 (N_2429,N_1985,N_1535);
nand U2430 (N_2430,N_1959,N_1445);
nor U2431 (N_2431,N_1440,N_1108);
nor U2432 (N_2432,N_1569,N_1771);
xnor U2433 (N_2433,N_1245,N_1954);
xnor U2434 (N_2434,N_1859,N_1163);
nand U2435 (N_2435,N_1130,N_1809);
and U2436 (N_2436,N_1728,N_1899);
nor U2437 (N_2437,N_1328,N_1049);
and U2438 (N_2438,N_1357,N_1034);
or U2439 (N_2439,N_1176,N_1561);
xor U2440 (N_2440,N_1707,N_1595);
nor U2441 (N_2441,N_1100,N_1621);
xor U2442 (N_2442,N_1774,N_1900);
nor U2443 (N_2443,N_1787,N_1558);
or U2444 (N_2444,N_1648,N_1554);
xnor U2445 (N_2445,N_1997,N_1401);
or U2446 (N_2446,N_1876,N_1187);
or U2447 (N_2447,N_1894,N_1140);
or U2448 (N_2448,N_1263,N_1012);
xnor U2449 (N_2449,N_1519,N_1600);
or U2450 (N_2450,N_1303,N_1157);
or U2451 (N_2451,N_1781,N_1169);
nand U2452 (N_2452,N_1408,N_1520);
xor U2453 (N_2453,N_1449,N_1933);
nand U2454 (N_2454,N_1467,N_1390);
xor U2455 (N_2455,N_1003,N_1293);
nand U2456 (N_2456,N_1726,N_1386);
nand U2457 (N_2457,N_1111,N_1405);
nor U2458 (N_2458,N_1500,N_1524);
or U2459 (N_2459,N_1754,N_1525);
or U2460 (N_2460,N_1950,N_1767);
or U2461 (N_2461,N_1201,N_1139);
nor U2462 (N_2462,N_1155,N_1272);
nand U2463 (N_2463,N_1526,N_1013);
and U2464 (N_2464,N_1000,N_1931);
nor U2465 (N_2465,N_1222,N_1971);
xnor U2466 (N_2466,N_1337,N_1618);
or U2467 (N_2467,N_1232,N_1039);
and U2468 (N_2468,N_1901,N_1047);
or U2469 (N_2469,N_1851,N_1308);
or U2470 (N_2470,N_1665,N_1953);
nor U2471 (N_2471,N_1693,N_1215);
or U2472 (N_2472,N_1544,N_1382);
or U2473 (N_2473,N_1361,N_1656);
or U2474 (N_2474,N_1070,N_1941);
or U2475 (N_2475,N_1466,N_1077);
xnor U2476 (N_2476,N_1607,N_1415);
and U2477 (N_2477,N_1834,N_1256);
or U2478 (N_2478,N_1949,N_1167);
xor U2479 (N_2479,N_1845,N_1044);
xnor U2480 (N_2480,N_1040,N_1567);
xnor U2481 (N_2481,N_1623,N_1260);
and U2482 (N_2482,N_1437,N_1527);
xor U2483 (N_2483,N_1619,N_1494);
nand U2484 (N_2484,N_1339,N_1783);
xor U2485 (N_2485,N_1488,N_1164);
nor U2486 (N_2486,N_1902,N_1284);
xnor U2487 (N_2487,N_1606,N_1694);
nand U2488 (N_2488,N_1154,N_1457);
and U2489 (N_2489,N_1206,N_1071);
or U2490 (N_2490,N_1907,N_1478);
or U2491 (N_2491,N_1635,N_1689);
and U2492 (N_2492,N_1347,N_1331);
nor U2493 (N_2493,N_1214,N_1709);
xnor U2494 (N_2494,N_1391,N_1468);
xnor U2495 (N_2495,N_1518,N_1388);
and U2496 (N_2496,N_1666,N_1878);
and U2497 (N_2497,N_1041,N_1319);
nor U2498 (N_2498,N_1123,N_1009);
or U2499 (N_2499,N_1778,N_1560);
or U2500 (N_2500,N_1482,N_1278);
xor U2501 (N_2501,N_1234,N_1644);
and U2502 (N_2502,N_1262,N_1015);
nor U2503 (N_2503,N_1958,N_1994);
xnor U2504 (N_2504,N_1238,N_1395);
xor U2505 (N_2505,N_1176,N_1703);
xnor U2506 (N_2506,N_1554,N_1534);
xor U2507 (N_2507,N_1484,N_1711);
nor U2508 (N_2508,N_1418,N_1733);
xnor U2509 (N_2509,N_1969,N_1517);
nor U2510 (N_2510,N_1710,N_1732);
nor U2511 (N_2511,N_1276,N_1845);
and U2512 (N_2512,N_1166,N_1705);
and U2513 (N_2513,N_1402,N_1941);
or U2514 (N_2514,N_1754,N_1608);
or U2515 (N_2515,N_1219,N_1080);
and U2516 (N_2516,N_1187,N_1793);
nor U2517 (N_2517,N_1425,N_1595);
or U2518 (N_2518,N_1847,N_1890);
nand U2519 (N_2519,N_1864,N_1506);
and U2520 (N_2520,N_1488,N_1950);
or U2521 (N_2521,N_1610,N_1474);
and U2522 (N_2522,N_1266,N_1098);
and U2523 (N_2523,N_1863,N_1891);
xnor U2524 (N_2524,N_1244,N_1043);
and U2525 (N_2525,N_1820,N_1138);
and U2526 (N_2526,N_1487,N_1444);
nor U2527 (N_2527,N_1485,N_1482);
and U2528 (N_2528,N_1091,N_1591);
and U2529 (N_2529,N_1548,N_1022);
and U2530 (N_2530,N_1560,N_1026);
nand U2531 (N_2531,N_1762,N_1606);
or U2532 (N_2532,N_1938,N_1317);
or U2533 (N_2533,N_1395,N_1495);
and U2534 (N_2534,N_1138,N_1969);
nor U2535 (N_2535,N_1392,N_1881);
nor U2536 (N_2536,N_1379,N_1465);
nor U2537 (N_2537,N_1919,N_1851);
and U2538 (N_2538,N_1177,N_1865);
or U2539 (N_2539,N_1406,N_1032);
nor U2540 (N_2540,N_1901,N_1376);
xnor U2541 (N_2541,N_1170,N_1083);
nor U2542 (N_2542,N_1483,N_1025);
xnor U2543 (N_2543,N_1121,N_1954);
and U2544 (N_2544,N_1465,N_1512);
and U2545 (N_2545,N_1118,N_1746);
nand U2546 (N_2546,N_1168,N_1803);
xnor U2547 (N_2547,N_1020,N_1491);
nor U2548 (N_2548,N_1046,N_1268);
and U2549 (N_2549,N_1885,N_1564);
nand U2550 (N_2550,N_1979,N_1389);
or U2551 (N_2551,N_1361,N_1943);
or U2552 (N_2552,N_1450,N_1887);
or U2553 (N_2553,N_1070,N_1145);
xor U2554 (N_2554,N_1230,N_1062);
xor U2555 (N_2555,N_1480,N_1281);
or U2556 (N_2556,N_1250,N_1120);
and U2557 (N_2557,N_1035,N_1350);
and U2558 (N_2558,N_1590,N_1153);
and U2559 (N_2559,N_1825,N_1925);
xor U2560 (N_2560,N_1267,N_1044);
and U2561 (N_2561,N_1151,N_1323);
xor U2562 (N_2562,N_1285,N_1752);
and U2563 (N_2563,N_1340,N_1972);
and U2564 (N_2564,N_1824,N_1411);
nand U2565 (N_2565,N_1391,N_1823);
xnor U2566 (N_2566,N_1075,N_1817);
xor U2567 (N_2567,N_1070,N_1283);
xnor U2568 (N_2568,N_1602,N_1610);
nand U2569 (N_2569,N_1707,N_1843);
xnor U2570 (N_2570,N_1539,N_1846);
xor U2571 (N_2571,N_1840,N_1516);
nand U2572 (N_2572,N_1558,N_1365);
or U2573 (N_2573,N_1524,N_1053);
xnor U2574 (N_2574,N_1640,N_1686);
nand U2575 (N_2575,N_1121,N_1863);
nor U2576 (N_2576,N_1823,N_1393);
and U2577 (N_2577,N_1156,N_1867);
nor U2578 (N_2578,N_1312,N_1945);
and U2579 (N_2579,N_1454,N_1523);
xor U2580 (N_2580,N_1239,N_1828);
and U2581 (N_2581,N_1533,N_1428);
and U2582 (N_2582,N_1416,N_1122);
and U2583 (N_2583,N_1766,N_1704);
and U2584 (N_2584,N_1564,N_1824);
nor U2585 (N_2585,N_1088,N_1037);
or U2586 (N_2586,N_1351,N_1703);
or U2587 (N_2587,N_1990,N_1717);
xor U2588 (N_2588,N_1875,N_1120);
nor U2589 (N_2589,N_1500,N_1818);
xnor U2590 (N_2590,N_1012,N_1493);
or U2591 (N_2591,N_1273,N_1676);
xnor U2592 (N_2592,N_1622,N_1015);
xnor U2593 (N_2593,N_1249,N_1812);
or U2594 (N_2594,N_1783,N_1427);
or U2595 (N_2595,N_1060,N_1604);
or U2596 (N_2596,N_1505,N_1394);
nor U2597 (N_2597,N_1616,N_1498);
nand U2598 (N_2598,N_1417,N_1955);
nor U2599 (N_2599,N_1702,N_1186);
nand U2600 (N_2600,N_1131,N_1465);
xor U2601 (N_2601,N_1917,N_1632);
nand U2602 (N_2602,N_1866,N_1387);
nor U2603 (N_2603,N_1693,N_1672);
and U2604 (N_2604,N_1557,N_1978);
nand U2605 (N_2605,N_1433,N_1607);
nor U2606 (N_2606,N_1292,N_1680);
nand U2607 (N_2607,N_1001,N_1650);
nor U2608 (N_2608,N_1329,N_1508);
xor U2609 (N_2609,N_1682,N_1167);
and U2610 (N_2610,N_1327,N_1360);
nand U2611 (N_2611,N_1559,N_1327);
nand U2612 (N_2612,N_1707,N_1637);
nand U2613 (N_2613,N_1517,N_1502);
nor U2614 (N_2614,N_1581,N_1988);
or U2615 (N_2615,N_1220,N_1242);
and U2616 (N_2616,N_1059,N_1315);
nor U2617 (N_2617,N_1528,N_1636);
and U2618 (N_2618,N_1016,N_1460);
nor U2619 (N_2619,N_1958,N_1178);
xor U2620 (N_2620,N_1902,N_1731);
nand U2621 (N_2621,N_1846,N_1930);
nand U2622 (N_2622,N_1686,N_1511);
nor U2623 (N_2623,N_1356,N_1674);
nand U2624 (N_2624,N_1272,N_1529);
and U2625 (N_2625,N_1742,N_1162);
nor U2626 (N_2626,N_1017,N_1011);
nor U2627 (N_2627,N_1756,N_1788);
xnor U2628 (N_2628,N_1305,N_1805);
nor U2629 (N_2629,N_1554,N_1760);
nand U2630 (N_2630,N_1481,N_1052);
xnor U2631 (N_2631,N_1565,N_1416);
nor U2632 (N_2632,N_1120,N_1343);
xor U2633 (N_2633,N_1548,N_1197);
xnor U2634 (N_2634,N_1478,N_1684);
and U2635 (N_2635,N_1723,N_1714);
xor U2636 (N_2636,N_1093,N_1742);
and U2637 (N_2637,N_1043,N_1986);
or U2638 (N_2638,N_1754,N_1269);
or U2639 (N_2639,N_1598,N_1333);
and U2640 (N_2640,N_1467,N_1218);
xnor U2641 (N_2641,N_1593,N_1178);
nand U2642 (N_2642,N_1395,N_1401);
nand U2643 (N_2643,N_1333,N_1951);
and U2644 (N_2644,N_1913,N_1632);
nor U2645 (N_2645,N_1355,N_1334);
or U2646 (N_2646,N_1130,N_1713);
nand U2647 (N_2647,N_1417,N_1452);
nor U2648 (N_2648,N_1163,N_1141);
xor U2649 (N_2649,N_1635,N_1981);
nand U2650 (N_2650,N_1132,N_1894);
and U2651 (N_2651,N_1495,N_1030);
nor U2652 (N_2652,N_1753,N_1804);
nor U2653 (N_2653,N_1616,N_1495);
and U2654 (N_2654,N_1243,N_1424);
nand U2655 (N_2655,N_1873,N_1433);
nand U2656 (N_2656,N_1313,N_1003);
and U2657 (N_2657,N_1111,N_1892);
nand U2658 (N_2658,N_1914,N_1835);
or U2659 (N_2659,N_1326,N_1313);
nor U2660 (N_2660,N_1802,N_1384);
xor U2661 (N_2661,N_1272,N_1188);
nor U2662 (N_2662,N_1148,N_1858);
nand U2663 (N_2663,N_1087,N_1113);
and U2664 (N_2664,N_1564,N_1286);
or U2665 (N_2665,N_1491,N_1492);
and U2666 (N_2666,N_1591,N_1018);
or U2667 (N_2667,N_1470,N_1827);
nand U2668 (N_2668,N_1868,N_1524);
nand U2669 (N_2669,N_1654,N_1348);
or U2670 (N_2670,N_1828,N_1125);
and U2671 (N_2671,N_1266,N_1675);
and U2672 (N_2672,N_1269,N_1724);
and U2673 (N_2673,N_1516,N_1763);
and U2674 (N_2674,N_1582,N_1269);
or U2675 (N_2675,N_1103,N_1438);
nor U2676 (N_2676,N_1081,N_1697);
xor U2677 (N_2677,N_1231,N_1293);
nor U2678 (N_2678,N_1177,N_1412);
xor U2679 (N_2679,N_1809,N_1000);
nor U2680 (N_2680,N_1268,N_1682);
nand U2681 (N_2681,N_1051,N_1615);
nand U2682 (N_2682,N_1161,N_1895);
xor U2683 (N_2683,N_1130,N_1886);
nand U2684 (N_2684,N_1199,N_1918);
or U2685 (N_2685,N_1031,N_1932);
nor U2686 (N_2686,N_1900,N_1643);
or U2687 (N_2687,N_1378,N_1563);
or U2688 (N_2688,N_1581,N_1869);
nor U2689 (N_2689,N_1995,N_1538);
xor U2690 (N_2690,N_1548,N_1655);
or U2691 (N_2691,N_1819,N_1253);
and U2692 (N_2692,N_1231,N_1817);
nand U2693 (N_2693,N_1597,N_1523);
nor U2694 (N_2694,N_1588,N_1028);
nor U2695 (N_2695,N_1249,N_1677);
xnor U2696 (N_2696,N_1048,N_1049);
xnor U2697 (N_2697,N_1757,N_1365);
or U2698 (N_2698,N_1865,N_1066);
nor U2699 (N_2699,N_1252,N_1629);
xor U2700 (N_2700,N_1964,N_1757);
nand U2701 (N_2701,N_1417,N_1554);
and U2702 (N_2702,N_1506,N_1796);
and U2703 (N_2703,N_1539,N_1006);
nand U2704 (N_2704,N_1582,N_1654);
xnor U2705 (N_2705,N_1647,N_1344);
xnor U2706 (N_2706,N_1524,N_1955);
and U2707 (N_2707,N_1655,N_1661);
nor U2708 (N_2708,N_1197,N_1513);
or U2709 (N_2709,N_1434,N_1216);
and U2710 (N_2710,N_1439,N_1402);
xor U2711 (N_2711,N_1311,N_1978);
xnor U2712 (N_2712,N_1607,N_1889);
or U2713 (N_2713,N_1070,N_1398);
or U2714 (N_2714,N_1477,N_1206);
nand U2715 (N_2715,N_1342,N_1264);
and U2716 (N_2716,N_1038,N_1978);
or U2717 (N_2717,N_1881,N_1398);
or U2718 (N_2718,N_1928,N_1913);
nor U2719 (N_2719,N_1730,N_1972);
nand U2720 (N_2720,N_1474,N_1524);
nor U2721 (N_2721,N_1986,N_1210);
or U2722 (N_2722,N_1893,N_1756);
and U2723 (N_2723,N_1862,N_1631);
nor U2724 (N_2724,N_1596,N_1039);
nor U2725 (N_2725,N_1725,N_1045);
xnor U2726 (N_2726,N_1965,N_1731);
or U2727 (N_2727,N_1468,N_1563);
and U2728 (N_2728,N_1221,N_1149);
xor U2729 (N_2729,N_1180,N_1619);
and U2730 (N_2730,N_1948,N_1952);
xnor U2731 (N_2731,N_1906,N_1902);
nor U2732 (N_2732,N_1423,N_1052);
xnor U2733 (N_2733,N_1551,N_1447);
and U2734 (N_2734,N_1909,N_1231);
xnor U2735 (N_2735,N_1485,N_1715);
and U2736 (N_2736,N_1448,N_1750);
nor U2737 (N_2737,N_1526,N_1349);
xor U2738 (N_2738,N_1304,N_1163);
xnor U2739 (N_2739,N_1881,N_1017);
xor U2740 (N_2740,N_1534,N_1895);
nand U2741 (N_2741,N_1878,N_1455);
nor U2742 (N_2742,N_1939,N_1842);
xnor U2743 (N_2743,N_1346,N_1570);
xor U2744 (N_2744,N_1287,N_1435);
nand U2745 (N_2745,N_1049,N_1653);
nand U2746 (N_2746,N_1384,N_1999);
and U2747 (N_2747,N_1754,N_1370);
xor U2748 (N_2748,N_1520,N_1038);
or U2749 (N_2749,N_1720,N_1485);
xor U2750 (N_2750,N_1173,N_1449);
nand U2751 (N_2751,N_1986,N_1445);
nor U2752 (N_2752,N_1365,N_1533);
and U2753 (N_2753,N_1734,N_1228);
nand U2754 (N_2754,N_1243,N_1907);
or U2755 (N_2755,N_1330,N_1168);
xnor U2756 (N_2756,N_1612,N_1526);
nor U2757 (N_2757,N_1310,N_1386);
and U2758 (N_2758,N_1612,N_1064);
nor U2759 (N_2759,N_1482,N_1267);
and U2760 (N_2760,N_1921,N_1486);
nand U2761 (N_2761,N_1553,N_1616);
nor U2762 (N_2762,N_1107,N_1477);
nor U2763 (N_2763,N_1136,N_1557);
xnor U2764 (N_2764,N_1744,N_1672);
nor U2765 (N_2765,N_1199,N_1978);
or U2766 (N_2766,N_1545,N_1280);
xnor U2767 (N_2767,N_1650,N_1981);
or U2768 (N_2768,N_1348,N_1005);
nand U2769 (N_2769,N_1262,N_1376);
xor U2770 (N_2770,N_1591,N_1194);
nor U2771 (N_2771,N_1485,N_1490);
or U2772 (N_2772,N_1789,N_1894);
nor U2773 (N_2773,N_1845,N_1248);
and U2774 (N_2774,N_1430,N_1272);
or U2775 (N_2775,N_1471,N_1503);
nand U2776 (N_2776,N_1792,N_1048);
or U2777 (N_2777,N_1976,N_1347);
and U2778 (N_2778,N_1606,N_1210);
nor U2779 (N_2779,N_1905,N_1141);
xnor U2780 (N_2780,N_1164,N_1217);
and U2781 (N_2781,N_1908,N_1409);
nand U2782 (N_2782,N_1097,N_1256);
nand U2783 (N_2783,N_1544,N_1566);
xnor U2784 (N_2784,N_1635,N_1559);
xor U2785 (N_2785,N_1166,N_1935);
nand U2786 (N_2786,N_1059,N_1531);
or U2787 (N_2787,N_1024,N_1351);
xnor U2788 (N_2788,N_1402,N_1199);
nand U2789 (N_2789,N_1407,N_1569);
and U2790 (N_2790,N_1845,N_1170);
and U2791 (N_2791,N_1075,N_1873);
nand U2792 (N_2792,N_1877,N_1954);
or U2793 (N_2793,N_1188,N_1860);
nor U2794 (N_2794,N_1799,N_1542);
nor U2795 (N_2795,N_1493,N_1195);
xnor U2796 (N_2796,N_1514,N_1290);
and U2797 (N_2797,N_1857,N_1413);
or U2798 (N_2798,N_1266,N_1180);
nand U2799 (N_2799,N_1329,N_1295);
or U2800 (N_2800,N_1135,N_1531);
nand U2801 (N_2801,N_1818,N_1035);
nand U2802 (N_2802,N_1720,N_1428);
and U2803 (N_2803,N_1917,N_1237);
and U2804 (N_2804,N_1095,N_1014);
nor U2805 (N_2805,N_1435,N_1970);
or U2806 (N_2806,N_1477,N_1480);
and U2807 (N_2807,N_1449,N_1481);
xor U2808 (N_2808,N_1688,N_1610);
and U2809 (N_2809,N_1068,N_1777);
and U2810 (N_2810,N_1129,N_1033);
nor U2811 (N_2811,N_1650,N_1318);
xor U2812 (N_2812,N_1832,N_1181);
and U2813 (N_2813,N_1452,N_1357);
nor U2814 (N_2814,N_1041,N_1703);
xor U2815 (N_2815,N_1393,N_1533);
and U2816 (N_2816,N_1571,N_1468);
xor U2817 (N_2817,N_1482,N_1096);
xnor U2818 (N_2818,N_1987,N_1304);
or U2819 (N_2819,N_1744,N_1566);
nor U2820 (N_2820,N_1046,N_1305);
nand U2821 (N_2821,N_1772,N_1152);
and U2822 (N_2822,N_1865,N_1986);
and U2823 (N_2823,N_1001,N_1901);
nor U2824 (N_2824,N_1755,N_1226);
nor U2825 (N_2825,N_1921,N_1720);
nor U2826 (N_2826,N_1692,N_1484);
and U2827 (N_2827,N_1692,N_1894);
nand U2828 (N_2828,N_1359,N_1366);
and U2829 (N_2829,N_1158,N_1395);
and U2830 (N_2830,N_1639,N_1298);
and U2831 (N_2831,N_1685,N_1177);
nand U2832 (N_2832,N_1105,N_1272);
and U2833 (N_2833,N_1546,N_1463);
nand U2834 (N_2834,N_1096,N_1442);
and U2835 (N_2835,N_1338,N_1485);
xor U2836 (N_2836,N_1703,N_1458);
or U2837 (N_2837,N_1333,N_1924);
or U2838 (N_2838,N_1623,N_1729);
nand U2839 (N_2839,N_1775,N_1894);
or U2840 (N_2840,N_1119,N_1640);
xor U2841 (N_2841,N_1889,N_1071);
nand U2842 (N_2842,N_1944,N_1408);
xnor U2843 (N_2843,N_1527,N_1896);
or U2844 (N_2844,N_1539,N_1116);
nor U2845 (N_2845,N_1738,N_1378);
nor U2846 (N_2846,N_1207,N_1606);
and U2847 (N_2847,N_1457,N_1385);
and U2848 (N_2848,N_1968,N_1285);
xnor U2849 (N_2849,N_1722,N_1092);
or U2850 (N_2850,N_1449,N_1913);
nor U2851 (N_2851,N_1994,N_1769);
and U2852 (N_2852,N_1073,N_1589);
or U2853 (N_2853,N_1271,N_1746);
xnor U2854 (N_2854,N_1498,N_1478);
xor U2855 (N_2855,N_1409,N_1130);
nand U2856 (N_2856,N_1881,N_1251);
and U2857 (N_2857,N_1039,N_1640);
xnor U2858 (N_2858,N_1983,N_1993);
and U2859 (N_2859,N_1294,N_1319);
or U2860 (N_2860,N_1754,N_1554);
nor U2861 (N_2861,N_1728,N_1844);
or U2862 (N_2862,N_1228,N_1175);
xnor U2863 (N_2863,N_1159,N_1481);
nor U2864 (N_2864,N_1085,N_1418);
xnor U2865 (N_2865,N_1385,N_1748);
and U2866 (N_2866,N_1074,N_1313);
nor U2867 (N_2867,N_1450,N_1032);
nor U2868 (N_2868,N_1825,N_1170);
xnor U2869 (N_2869,N_1436,N_1111);
and U2870 (N_2870,N_1563,N_1251);
and U2871 (N_2871,N_1171,N_1489);
nand U2872 (N_2872,N_1733,N_1652);
nand U2873 (N_2873,N_1732,N_1450);
or U2874 (N_2874,N_1296,N_1988);
nor U2875 (N_2875,N_1858,N_1102);
nor U2876 (N_2876,N_1054,N_1220);
or U2877 (N_2877,N_1284,N_1585);
or U2878 (N_2878,N_1190,N_1196);
or U2879 (N_2879,N_1770,N_1868);
nor U2880 (N_2880,N_1142,N_1812);
xor U2881 (N_2881,N_1076,N_1188);
or U2882 (N_2882,N_1702,N_1917);
nor U2883 (N_2883,N_1709,N_1003);
or U2884 (N_2884,N_1485,N_1429);
xnor U2885 (N_2885,N_1812,N_1388);
or U2886 (N_2886,N_1326,N_1001);
nand U2887 (N_2887,N_1891,N_1509);
nand U2888 (N_2888,N_1691,N_1951);
nand U2889 (N_2889,N_1642,N_1154);
nor U2890 (N_2890,N_1309,N_1363);
nor U2891 (N_2891,N_1017,N_1590);
nand U2892 (N_2892,N_1831,N_1624);
xnor U2893 (N_2893,N_1434,N_1581);
xnor U2894 (N_2894,N_1106,N_1811);
nor U2895 (N_2895,N_1782,N_1247);
nor U2896 (N_2896,N_1143,N_1583);
nand U2897 (N_2897,N_1841,N_1664);
nor U2898 (N_2898,N_1333,N_1482);
nor U2899 (N_2899,N_1713,N_1194);
nor U2900 (N_2900,N_1839,N_1801);
and U2901 (N_2901,N_1562,N_1712);
xnor U2902 (N_2902,N_1453,N_1832);
nor U2903 (N_2903,N_1859,N_1743);
nor U2904 (N_2904,N_1029,N_1590);
nor U2905 (N_2905,N_1378,N_1600);
and U2906 (N_2906,N_1609,N_1107);
nor U2907 (N_2907,N_1489,N_1167);
and U2908 (N_2908,N_1884,N_1228);
nor U2909 (N_2909,N_1947,N_1380);
and U2910 (N_2910,N_1838,N_1341);
nor U2911 (N_2911,N_1834,N_1223);
xor U2912 (N_2912,N_1566,N_1236);
nand U2913 (N_2913,N_1876,N_1091);
xnor U2914 (N_2914,N_1364,N_1007);
nor U2915 (N_2915,N_1727,N_1130);
xor U2916 (N_2916,N_1469,N_1418);
nor U2917 (N_2917,N_1221,N_1578);
or U2918 (N_2918,N_1925,N_1697);
xor U2919 (N_2919,N_1740,N_1932);
nor U2920 (N_2920,N_1456,N_1967);
or U2921 (N_2921,N_1468,N_1992);
xnor U2922 (N_2922,N_1484,N_1193);
nand U2923 (N_2923,N_1324,N_1343);
nor U2924 (N_2924,N_1510,N_1775);
and U2925 (N_2925,N_1228,N_1424);
nand U2926 (N_2926,N_1313,N_1995);
xnor U2927 (N_2927,N_1504,N_1110);
nand U2928 (N_2928,N_1646,N_1555);
and U2929 (N_2929,N_1965,N_1801);
nand U2930 (N_2930,N_1293,N_1334);
and U2931 (N_2931,N_1444,N_1453);
xnor U2932 (N_2932,N_1457,N_1119);
xnor U2933 (N_2933,N_1061,N_1657);
nor U2934 (N_2934,N_1435,N_1832);
nor U2935 (N_2935,N_1311,N_1982);
xor U2936 (N_2936,N_1111,N_1449);
and U2937 (N_2937,N_1842,N_1729);
xor U2938 (N_2938,N_1589,N_1829);
nand U2939 (N_2939,N_1210,N_1257);
nand U2940 (N_2940,N_1939,N_1358);
xnor U2941 (N_2941,N_1568,N_1435);
nand U2942 (N_2942,N_1023,N_1294);
and U2943 (N_2943,N_1276,N_1157);
nor U2944 (N_2944,N_1191,N_1247);
nor U2945 (N_2945,N_1437,N_1265);
or U2946 (N_2946,N_1498,N_1954);
xnor U2947 (N_2947,N_1056,N_1411);
or U2948 (N_2948,N_1299,N_1965);
nor U2949 (N_2949,N_1437,N_1755);
xnor U2950 (N_2950,N_1358,N_1649);
or U2951 (N_2951,N_1779,N_1551);
xnor U2952 (N_2952,N_1439,N_1492);
or U2953 (N_2953,N_1980,N_1550);
nand U2954 (N_2954,N_1487,N_1912);
nand U2955 (N_2955,N_1552,N_1371);
or U2956 (N_2956,N_1878,N_1561);
and U2957 (N_2957,N_1688,N_1214);
xnor U2958 (N_2958,N_1159,N_1520);
and U2959 (N_2959,N_1700,N_1315);
nand U2960 (N_2960,N_1466,N_1493);
and U2961 (N_2961,N_1818,N_1691);
or U2962 (N_2962,N_1330,N_1367);
or U2963 (N_2963,N_1123,N_1756);
xnor U2964 (N_2964,N_1071,N_1127);
and U2965 (N_2965,N_1620,N_1204);
nor U2966 (N_2966,N_1972,N_1002);
and U2967 (N_2967,N_1638,N_1294);
nor U2968 (N_2968,N_1933,N_1143);
or U2969 (N_2969,N_1942,N_1916);
xnor U2970 (N_2970,N_1127,N_1214);
xnor U2971 (N_2971,N_1089,N_1363);
or U2972 (N_2972,N_1135,N_1594);
or U2973 (N_2973,N_1614,N_1829);
nand U2974 (N_2974,N_1347,N_1288);
nand U2975 (N_2975,N_1626,N_1867);
and U2976 (N_2976,N_1123,N_1312);
nand U2977 (N_2977,N_1110,N_1832);
nand U2978 (N_2978,N_1368,N_1323);
or U2979 (N_2979,N_1530,N_1470);
or U2980 (N_2980,N_1489,N_1423);
nor U2981 (N_2981,N_1927,N_1418);
nor U2982 (N_2982,N_1201,N_1588);
xnor U2983 (N_2983,N_1205,N_1536);
or U2984 (N_2984,N_1738,N_1844);
or U2985 (N_2985,N_1544,N_1912);
xor U2986 (N_2986,N_1288,N_1599);
and U2987 (N_2987,N_1118,N_1942);
or U2988 (N_2988,N_1078,N_1851);
or U2989 (N_2989,N_1526,N_1267);
xnor U2990 (N_2990,N_1792,N_1064);
nor U2991 (N_2991,N_1122,N_1661);
and U2992 (N_2992,N_1355,N_1637);
xor U2993 (N_2993,N_1298,N_1286);
or U2994 (N_2994,N_1134,N_1557);
nand U2995 (N_2995,N_1855,N_1113);
and U2996 (N_2996,N_1085,N_1720);
nand U2997 (N_2997,N_1427,N_1668);
nor U2998 (N_2998,N_1091,N_1100);
or U2999 (N_2999,N_1981,N_1388);
xor U3000 (N_3000,N_2298,N_2909);
nor U3001 (N_3001,N_2226,N_2274);
nand U3002 (N_3002,N_2306,N_2839);
xnor U3003 (N_3003,N_2930,N_2905);
nand U3004 (N_3004,N_2138,N_2410);
and U3005 (N_3005,N_2822,N_2624);
nor U3006 (N_3006,N_2239,N_2510);
or U3007 (N_3007,N_2921,N_2857);
nor U3008 (N_3008,N_2545,N_2266);
nor U3009 (N_3009,N_2901,N_2892);
xor U3010 (N_3010,N_2371,N_2590);
or U3011 (N_3011,N_2279,N_2358);
and U3012 (N_3012,N_2094,N_2418);
xnor U3013 (N_3013,N_2990,N_2565);
and U3014 (N_3014,N_2446,N_2307);
nand U3015 (N_3015,N_2402,N_2005);
nor U3016 (N_3016,N_2170,N_2063);
nor U3017 (N_3017,N_2889,N_2696);
nor U3018 (N_3018,N_2638,N_2136);
xor U3019 (N_3019,N_2300,N_2182);
and U3020 (N_3020,N_2619,N_2475);
or U3021 (N_3021,N_2335,N_2232);
xnor U3022 (N_3022,N_2734,N_2776);
or U3023 (N_3023,N_2961,N_2100);
xor U3024 (N_3024,N_2960,N_2914);
nor U3025 (N_3025,N_2424,N_2327);
xor U3026 (N_3026,N_2713,N_2497);
nor U3027 (N_3027,N_2016,N_2724);
nor U3028 (N_3028,N_2052,N_2049);
xnor U3029 (N_3029,N_2487,N_2374);
xnor U3030 (N_3030,N_2150,N_2096);
nand U3031 (N_3031,N_2254,N_2476);
and U3032 (N_3032,N_2981,N_2467);
nand U3033 (N_3033,N_2012,N_2847);
and U3034 (N_3034,N_2527,N_2652);
nor U3035 (N_3035,N_2861,N_2086);
nor U3036 (N_3036,N_2163,N_2607);
and U3037 (N_3037,N_2025,N_2470);
or U3038 (N_3038,N_2645,N_2864);
nand U3039 (N_3039,N_2200,N_2074);
and U3040 (N_3040,N_2918,N_2657);
and U3041 (N_3041,N_2473,N_2591);
nor U3042 (N_3042,N_2422,N_2433);
or U3043 (N_3043,N_2739,N_2492);
nor U3044 (N_3044,N_2479,N_2931);
nand U3045 (N_3045,N_2099,N_2186);
xor U3046 (N_3046,N_2962,N_2378);
nand U3047 (N_3047,N_2210,N_2557);
xnor U3048 (N_3048,N_2660,N_2583);
nor U3049 (N_3049,N_2205,N_2423);
nor U3050 (N_3050,N_2983,N_2152);
and U3051 (N_3051,N_2750,N_2425);
nand U3052 (N_3052,N_2754,N_2634);
nand U3053 (N_3053,N_2332,N_2268);
or U3054 (N_3054,N_2593,N_2865);
and U3055 (N_3055,N_2117,N_2569);
nand U3056 (N_3056,N_2044,N_2048);
nand U3057 (N_3057,N_2993,N_2089);
and U3058 (N_3058,N_2903,N_2489);
xor U3059 (N_3059,N_2775,N_2870);
xor U3060 (N_3060,N_2040,N_2669);
or U3061 (N_3061,N_2340,N_2508);
xor U3062 (N_3062,N_2401,N_2855);
or U3063 (N_3063,N_2649,N_2718);
nand U3064 (N_3064,N_2004,N_2925);
xor U3065 (N_3065,N_2400,N_2391);
or U3066 (N_3066,N_2689,N_2168);
or U3067 (N_3067,N_2428,N_2585);
xnor U3068 (N_3068,N_2547,N_2404);
xnor U3069 (N_3069,N_2654,N_2625);
and U3070 (N_3070,N_2280,N_2042);
nor U3071 (N_3071,N_2966,N_2072);
or U3072 (N_3072,N_2132,N_2351);
xnor U3073 (N_3073,N_2618,N_2924);
nand U3074 (N_3074,N_2490,N_2802);
and U3075 (N_3075,N_2106,N_2256);
xnor U3076 (N_3076,N_2753,N_2301);
or U3077 (N_3077,N_2050,N_2453);
or U3078 (N_3078,N_2154,N_2166);
or U3079 (N_3079,N_2071,N_2933);
or U3080 (N_3080,N_2881,N_2955);
xor U3081 (N_3081,N_2631,N_2816);
nor U3082 (N_3082,N_2524,N_2509);
and U3083 (N_3083,N_2720,N_2749);
nand U3084 (N_3084,N_2697,N_2965);
xor U3085 (N_3085,N_2602,N_2584);
nor U3086 (N_3086,N_2110,N_2693);
nand U3087 (N_3087,N_2437,N_2751);
and U3088 (N_3088,N_2324,N_2195);
and U3089 (N_3089,N_2465,N_2513);
nor U3090 (N_3090,N_2493,N_2766);
and U3091 (N_3091,N_2491,N_2309);
nand U3092 (N_3092,N_2989,N_2915);
xnor U3093 (N_3093,N_2204,N_2843);
and U3094 (N_3094,N_2258,N_2045);
nand U3095 (N_3095,N_2502,N_2633);
or U3096 (N_3096,N_2611,N_2676);
and U3097 (N_3097,N_2623,N_2572);
nand U3098 (N_3098,N_2169,N_2640);
or U3099 (N_3099,N_2786,N_2999);
nand U3100 (N_3100,N_2281,N_2725);
nor U3101 (N_3101,N_2587,N_2002);
and U3102 (N_3102,N_2155,N_2243);
nor U3103 (N_3103,N_2825,N_2135);
nand U3104 (N_3104,N_2963,N_2177);
or U3105 (N_3105,N_2790,N_2367);
xor U3106 (N_3106,N_2819,N_2503);
xnor U3107 (N_3107,N_2833,N_2831);
nor U3108 (N_3108,N_2873,N_2273);
or U3109 (N_3109,N_2159,N_2726);
xor U3110 (N_3110,N_2255,N_2488);
or U3111 (N_3111,N_2167,N_2445);
nor U3112 (N_3112,N_2917,N_2597);
and U3113 (N_3113,N_2015,N_2685);
and U3114 (N_3114,N_2541,N_2321);
nor U3115 (N_3115,N_2091,N_2779);
and U3116 (N_3116,N_2039,N_2011);
or U3117 (N_3117,N_2573,N_2608);
nor U3118 (N_3118,N_2616,N_2807);
xnor U3119 (N_3119,N_2265,N_2518);
or U3120 (N_3120,N_2483,N_2020);
or U3121 (N_3121,N_2067,N_2439);
and U3122 (N_3122,N_2604,N_2793);
xnor U3123 (N_3123,N_2691,N_2187);
nand U3124 (N_3124,N_2871,N_2532);
nor U3125 (N_3125,N_2125,N_2403);
nand U3126 (N_3126,N_2577,N_2795);
nor U3127 (N_3127,N_2061,N_2784);
nor U3128 (N_3128,N_2956,N_2594);
xor U3129 (N_3129,N_2008,N_2471);
nand U3130 (N_3130,N_2904,N_2610);
and U3131 (N_3131,N_2114,N_2938);
nand U3132 (N_3132,N_2299,N_2712);
and U3133 (N_3133,N_2076,N_2636);
and U3134 (N_3134,N_2107,N_2009);
and U3135 (N_3135,N_2600,N_2863);
or U3136 (N_3136,N_2460,N_2088);
xnor U3137 (N_3137,N_2038,N_2389);
or U3138 (N_3138,N_2264,N_2026);
nor U3139 (N_3139,N_2525,N_2916);
or U3140 (N_3140,N_2308,N_2238);
nand U3141 (N_3141,N_2995,N_2910);
xnor U3142 (N_3142,N_2858,N_2350);
nor U3143 (N_3143,N_2520,N_2868);
nor U3144 (N_3144,N_2162,N_2627);
nand U3145 (N_3145,N_2116,N_2664);
xnor U3146 (N_3146,N_2124,N_2303);
or U3147 (N_3147,N_2586,N_2349);
xor U3148 (N_3148,N_2806,N_2755);
nor U3149 (N_3149,N_2874,N_2006);
or U3150 (N_3150,N_2253,N_2021);
nand U3151 (N_3151,N_2103,N_2193);
xor U3152 (N_3152,N_2810,N_2261);
nor U3153 (N_3153,N_2536,N_2059);
nor U3154 (N_3154,N_2115,N_2366);
or U3155 (N_3155,N_2282,N_2970);
and U3156 (N_3156,N_2051,N_2856);
or U3157 (N_3157,N_2835,N_2443);
or U3158 (N_3158,N_2478,N_2364);
xor U3159 (N_3159,N_2249,N_2284);
nor U3160 (N_3160,N_2706,N_2369);
nand U3161 (N_3161,N_2133,N_2537);
and U3162 (N_3162,N_2582,N_2058);
and U3163 (N_3163,N_2801,N_2529);
or U3164 (N_3164,N_2242,N_2733);
and U3165 (N_3165,N_2820,N_2411);
and U3166 (N_3166,N_2758,N_2211);
xnor U3167 (N_3167,N_2534,N_2377);
nand U3168 (N_3168,N_2511,N_2416);
nand U3169 (N_3169,N_2866,N_2945);
or U3170 (N_3170,N_2558,N_2546);
and U3171 (N_3171,N_2845,N_2296);
nor U3172 (N_3172,N_2053,N_2174);
and U3173 (N_3173,N_2405,N_2531);
nand U3174 (N_3174,N_2375,N_2196);
nand U3175 (N_3175,N_2480,N_2251);
and U3176 (N_3176,N_2932,N_2544);
or U3177 (N_3177,N_2578,N_2474);
and U3178 (N_3178,N_2207,N_2768);
or U3179 (N_3179,N_2900,N_2986);
and U3180 (N_3180,N_2683,N_2774);
xor U3181 (N_3181,N_2716,N_2974);
nor U3182 (N_3182,N_2208,N_2289);
and U3183 (N_3183,N_2944,N_2287);
nand U3184 (N_3184,N_2212,N_2003);
xnor U3185 (N_3185,N_2496,N_2730);
nand U3186 (N_3186,N_2879,N_2746);
nor U3187 (N_3187,N_2551,N_2538);
and U3188 (N_3188,N_2789,N_2799);
xnor U3189 (N_3189,N_2421,N_2681);
and U3190 (N_3190,N_2798,N_2151);
nor U3191 (N_3191,N_2482,N_2736);
xnor U3192 (N_3192,N_2247,N_2939);
and U3193 (N_3193,N_2523,N_2957);
or U3194 (N_3194,N_2760,N_2568);
and U3195 (N_3195,N_2846,N_2215);
nor U3196 (N_3196,N_2969,N_2535);
and U3197 (N_3197,N_2522,N_2782);
and U3198 (N_3198,N_2269,N_2899);
nand U3199 (N_3199,N_2838,N_2704);
and U3200 (N_3200,N_2397,N_2415);
and U3201 (N_3201,N_2895,N_2887);
or U3202 (N_3202,N_2761,N_2142);
nand U3203 (N_3203,N_2398,N_2064);
or U3204 (N_3204,N_2875,N_2022);
and U3205 (N_3205,N_2548,N_2507);
and U3206 (N_3206,N_2632,N_2457);
nor U3207 (N_3207,N_2054,N_2455);
nor U3208 (N_3208,N_2773,N_2700);
nor U3209 (N_3209,N_2000,N_2090);
nand U3210 (N_3210,N_2926,N_2348);
and U3211 (N_3211,N_2047,N_2562);
xnor U3212 (N_3212,N_2729,N_2352);
xnor U3213 (N_3213,N_2841,N_2339);
or U3214 (N_3214,N_2392,N_2036);
nand U3215 (N_3215,N_2844,N_2069);
xnor U3216 (N_3216,N_2996,N_2705);
or U3217 (N_3217,N_2601,N_2438);
xor U3218 (N_3218,N_2250,N_2313);
nor U3219 (N_3219,N_2842,N_2043);
xor U3220 (N_3220,N_2224,N_2164);
or U3221 (N_3221,N_2894,N_2338);
nand U3222 (N_3222,N_2414,N_2456);
nand U3223 (N_3223,N_2271,N_2030);
and U3224 (N_3224,N_2646,N_2236);
and U3225 (N_3225,N_2526,N_2252);
nor U3226 (N_3226,N_2721,N_2588);
xor U3227 (N_3227,N_2670,N_2027);
xor U3228 (N_3228,N_2095,N_2714);
nor U3229 (N_3229,N_2673,N_2417);
xnor U3230 (N_3230,N_2908,N_2862);
or U3231 (N_3231,N_2628,N_2336);
or U3232 (N_3232,N_2517,N_2715);
or U3233 (N_3233,N_2785,N_2185);
and U3234 (N_3234,N_2988,N_2080);
xor U3235 (N_3235,N_2183,N_2085);
xnor U3236 (N_3236,N_2466,N_2245);
and U3237 (N_3237,N_2958,N_2675);
nor U3238 (N_3238,N_2678,N_2630);
xor U3239 (N_3239,N_2898,N_2292);
nand U3240 (N_3240,N_2554,N_2141);
or U3241 (N_3241,N_2019,N_2598);
xnor U3242 (N_3242,N_2028,N_2987);
nor U3243 (N_3243,N_2145,N_2564);
xnor U3244 (N_3244,N_2276,N_2160);
and U3245 (N_3245,N_2221,N_2780);
nand U3246 (N_3246,N_2686,N_2635);
or U3247 (N_3247,N_2362,N_2123);
nor U3248 (N_3248,N_2500,N_2288);
xor U3249 (N_3249,N_2495,N_2614);
xor U3250 (N_3250,N_2199,N_2001);
xor U3251 (N_3251,N_2192,N_2555);
or U3252 (N_3252,N_2745,N_2070);
and U3253 (N_3253,N_2528,N_2728);
or U3254 (N_3254,N_2940,N_2740);
nand U3255 (N_3255,N_2821,N_2688);
nand U3256 (N_3256,N_2815,N_2129);
nor U3257 (N_3257,N_2621,N_2384);
or U3258 (N_3258,N_2943,N_2663);
or U3259 (N_3259,N_2952,N_2575);
nand U3260 (N_3260,N_2967,N_2007);
nand U3261 (N_3261,N_2581,N_2566);
xor U3262 (N_3262,N_2073,N_2744);
nand U3263 (N_3263,N_2923,N_2620);
and U3264 (N_3264,N_2161,N_2355);
xor U3265 (N_3265,N_2891,N_2771);
nand U3266 (N_3266,N_2248,N_2363);
nor U3267 (N_3267,N_2450,N_2927);
or U3268 (N_3268,N_2172,N_2148);
nand U3269 (N_3269,N_2451,N_2440);
nand U3270 (N_3270,N_2748,N_2119);
or U3271 (N_3271,N_2330,N_2719);
and U3272 (N_3272,N_2413,N_2655);
and U3273 (N_3273,N_2214,N_2318);
nand U3274 (N_3274,N_2334,N_2886);
nand U3275 (N_3275,N_2687,N_2512);
nand U3276 (N_3276,N_2180,N_2477);
nor U3277 (N_3277,N_2257,N_2329);
and U3278 (N_3278,N_2209,N_2122);
or U3279 (N_3279,N_2263,N_2501);
or U3280 (N_3280,N_2794,N_2390);
nand U3281 (N_3281,N_2702,N_2919);
nor U3282 (N_3282,N_2156,N_2406);
and U3283 (N_3283,N_2230,N_2677);
nand U3284 (N_3284,N_2033,N_2950);
nand U3285 (N_3285,N_2157,N_2108);
nand U3286 (N_3286,N_2354,N_2991);
and U3287 (N_3287,N_2882,N_2171);
and U3288 (N_3288,N_2742,N_2244);
or U3289 (N_3289,N_2060,N_2971);
or U3290 (N_3290,N_2143,N_2087);
nor U3291 (N_3291,N_2034,N_2765);
nor U3292 (N_3292,N_2922,N_2722);
and U3293 (N_3293,N_2459,N_2829);
nor U3294 (N_3294,N_2066,N_2018);
and U3295 (N_3295,N_2852,N_2641);
nor U3296 (N_3296,N_2752,N_2978);
nor U3297 (N_3297,N_2104,N_2817);
and U3298 (N_3298,N_2788,N_2068);
nand U3299 (N_3299,N_2189,N_2651);
nand U3300 (N_3300,N_2854,N_2710);
nand U3301 (N_3301,N_2840,N_2202);
or U3302 (N_3302,N_2304,N_2851);
xor U3303 (N_3303,N_2783,N_2827);
or U3304 (N_3304,N_2468,N_2648);
nand U3305 (N_3305,N_2747,N_2432);
or U3306 (N_3306,N_2331,N_2549);
nor U3307 (N_3307,N_2121,N_2738);
and U3308 (N_3308,N_2533,N_2302);
and U3309 (N_3309,N_2826,N_2658);
or U3310 (N_3310,N_2241,N_2982);
xnor U3311 (N_3311,N_2395,N_2360);
and U3312 (N_3312,N_2772,N_2599);
or U3313 (N_3313,N_2046,N_2310);
nand U3314 (N_3314,N_2035,N_2345);
xnor U3315 (N_3315,N_2128,N_2234);
xnor U3316 (N_3316,N_2396,N_2949);
or U3317 (N_3317,N_2290,N_2435);
or U3318 (N_3318,N_2286,N_2201);
nand U3319 (N_3319,N_2612,N_2326);
or U3320 (N_3320,N_2556,N_2579);
nor U3321 (N_3321,N_2356,N_2191);
and U3322 (N_3322,N_2092,N_2563);
nand U3323 (N_3323,N_2973,N_2928);
and U3324 (N_3324,N_2540,N_2105);
or U3325 (N_3325,N_2173,N_2013);
nand U3326 (N_3326,N_2550,N_2486);
or U3327 (N_3327,N_2278,N_2316);
or U3328 (N_3328,N_2385,N_2231);
and U3329 (N_3329,N_2869,N_2665);
and U3330 (N_3330,N_2792,N_2770);
nor U3331 (N_3331,N_2684,N_2997);
xnor U3332 (N_3332,N_2325,N_2498);
xnor U3333 (N_3333,N_2951,N_2149);
nand U3334 (N_3334,N_2229,N_2659);
and U3335 (N_3335,N_2464,N_2661);
and U3336 (N_3336,N_2181,N_2357);
or U3337 (N_3337,N_2368,N_2393);
nor U3338 (N_3338,N_2408,N_2101);
and U3339 (N_3339,N_2184,N_2275);
and U3340 (N_3340,N_2017,N_2860);
xnor U3341 (N_3341,N_2376,N_2014);
xnor U3342 (N_3342,N_2606,N_2031);
xor U3343 (N_3343,N_2897,N_2504);
nor U3344 (N_3344,N_2373,N_2305);
nor U3345 (N_3345,N_2796,N_2065);
nor U3346 (N_3346,N_2297,N_2041);
xor U3347 (N_3347,N_2694,N_2342);
nor U3348 (N_3348,N_2707,N_2291);
nand U3349 (N_3349,N_2270,N_2977);
and U3350 (N_3350,N_2893,N_2217);
or U3351 (N_3351,N_2672,N_2530);
nor U3352 (N_3352,N_2319,N_2823);
or U3353 (N_3353,N_2723,N_2797);
or U3354 (N_3354,N_2818,N_2920);
xor U3355 (N_3355,N_2223,N_2140);
xnor U3356 (N_3356,N_2260,N_2580);
nor U3357 (N_3357,N_2102,N_2222);
nor U3358 (N_3358,N_2442,N_2727);
xor U3359 (N_3359,N_2849,N_2711);
or U3360 (N_3360,N_2777,N_2539);
nand U3361 (N_3361,N_2589,N_2343);
and U3362 (N_3362,N_2936,N_2639);
xor U3363 (N_3363,N_2552,N_2394);
xor U3364 (N_3364,N_2165,N_2828);
nor U3365 (N_3365,N_2097,N_2285);
or U3366 (N_3366,N_2194,N_2848);
nand U3367 (N_3367,N_2188,N_2913);
and U3368 (N_3368,N_2671,N_2571);
or U3369 (N_3369,N_2998,N_2975);
nor U3370 (N_3370,N_2314,N_2429);
nor U3371 (N_3371,N_2344,N_2543);
and U3372 (N_3372,N_2937,N_2472);
nor U3373 (N_3373,N_2312,N_2246);
and U3374 (N_3374,N_2622,N_2494);
or U3375 (N_3375,N_2515,N_2227);
nand U3376 (N_3376,N_2505,N_2444);
nand U3377 (N_3377,N_2888,N_2656);
nor U3378 (N_3378,N_2032,N_2463);
nor U3379 (N_3379,N_2380,N_2062);
and U3380 (N_3380,N_2853,N_2240);
nand U3381 (N_3381,N_2735,N_2650);
or U3382 (N_3382,N_2653,N_2878);
and U3383 (N_3383,N_2272,N_2323);
nor U3384 (N_3384,N_2934,N_2462);
xnor U3385 (N_3385,N_2617,N_2809);
and U3386 (N_3386,N_2430,N_2832);
and U3387 (N_3387,N_2093,N_2521);
nor U3388 (N_3388,N_2233,N_2762);
or U3389 (N_3389,N_2322,N_2984);
nor U3390 (N_3390,N_2884,N_2056);
and U3391 (N_3391,N_2144,N_2979);
or U3392 (N_3392,N_2458,N_2461);
or U3393 (N_3393,N_2388,N_2057);
or U3394 (N_3394,N_2811,N_2109);
xnor U3395 (N_3395,N_2929,N_2499);
or U3396 (N_3396,N_2203,N_2347);
and U3397 (N_3397,N_2381,N_2346);
and U3398 (N_3398,N_2830,N_2448);
xor U3399 (N_3399,N_2759,N_2902);
and U3400 (N_3400,N_2426,N_2225);
nand U3401 (N_3401,N_2698,N_2077);
or U3402 (N_3402,N_2262,N_2146);
or U3403 (N_3403,N_2680,N_2972);
nand U3404 (N_3404,N_2359,N_2701);
and U3405 (N_3405,N_2592,N_2130);
and U3406 (N_3406,N_2791,N_2328);
xor U3407 (N_3407,N_2741,N_2912);
or U3408 (N_3408,N_2695,N_2337);
xor U3409 (N_3409,N_2075,N_2294);
or U3410 (N_3410,N_2519,N_2382);
nor U3411 (N_3411,N_2737,N_2703);
nand U3412 (N_3412,N_2023,N_2668);
and U3413 (N_3413,N_2213,N_2341);
or U3414 (N_3414,N_2506,N_2699);
xor U3415 (N_3415,N_2690,N_2948);
nand U3416 (N_3416,N_2235,N_2372);
or U3417 (N_3417,N_2662,N_2804);
nand U3418 (N_3418,N_2353,N_2743);
or U3419 (N_3419,N_2179,N_2436);
xnor U3420 (N_3420,N_2813,N_2370);
xnor U3421 (N_3421,N_2824,N_2609);
xor U3422 (N_3422,N_2876,N_2010);
xor U3423 (N_3423,N_2559,N_2808);
nor U3424 (N_3424,N_2709,N_2764);
xnor U3425 (N_3425,N_2126,N_2283);
nand U3426 (N_3426,N_2434,N_2576);
nor U3427 (N_3427,N_2431,N_2112);
and U3428 (N_3428,N_2137,N_2814);
and U3429 (N_3429,N_2427,N_2859);
nor U3430 (N_3430,N_2111,N_2935);
and U3431 (N_3431,N_2120,N_2980);
or U3432 (N_3432,N_2964,N_2365);
nand U3433 (N_3433,N_2731,N_2454);
and U3434 (N_3434,N_2647,N_2642);
xnor U3435 (N_3435,N_2667,N_2985);
or U3436 (N_3436,N_2781,N_2158);
nand U3437 (N_3437,N_2637,N_2293);
or U3438 (N_3438,N_2763,N_2867);
or U3439 (N_3439,N_2024,N_2147);
and U3440 (N_3440,N_2139,N_2767);
or U3441 (N_3441,N_2084,N_2834);
nand U3442 (N_3442,N_2644,N_2134);
nand U3443 (N_3443,N_2883,N_2947);
nand U3444 (N_3444,N_2769,N_2399);
and U3445 (N_3445,N_2872,N_2409);
and U3446 (N_3446,N_2954,N_2216);
and U3447 (N_3447,N_2055,N_2542);
nand U3448 (N_3448,N_2412,N_2447);
nor U3449 (N_3449,N_2469,N_2732);
xnor U3450 (N_3450,N_2946,N_2603);
nand U3451 (N_3451,N_2516,N_2386);
nor U3452 (N_3452,N_2311,N_2315);
and U3453 (N_3453,N_2570,N_2595);
nor U3454 (N_3454,N_2992,N_2837);
and U3455 (N_3455,N_2407,N_2198);
or U3456 (N_3456,N_2485,N_2452);
xnor U3457 (N_3457,N_2885,N_2953);
xnor U3458 (N_3458,N_2994,N_2850);
xnor U3459 (N_3459,N_2757,N_2220);
nand U3460 (N_3460,N_2277,N_2803);
and U3461 (N_3461,N_2596,N_2379);
or U3462 (N_3462,N_2514,N_2441);
xor U3463 (N_3463,N_2896,N_2419);
or U3464 (N_3464,N_2666,N_2228);
and U3465 (N_3465,N_2605,N_2081);
or U3466 (N_3466,N_2127,N_2387);
xnor U3467 (N_3467,N_2083,N_2037);
xnor U3468 (N_3468,N_2082,N_2237);
nor U3469 (N_3469,N_2449,N_2880);
and U3470 (N_3470,N_2259,N_2175);
nor U3471 (N_3471,N_2560,N_2484);
and U3472 (N_3472,N_2078,N_2643);
nand U3473 (N_3473,N_2629,N_2911);
and U3474 (N_3474,N_2567,N_2812);
xor U3475 (N_3475,N_2787,N_2333);
xor U3476 (N_3476,N_2178,N_2361);
and U3477 (N_3477,N_2190,N_2890);
and U3478 (N_3478,N_2613,N_2968);
nor U3479 (N_3479,N_2692,N_2079);
nand U3480 (N_3480,N_2717,N_2317);
nand U3481 (N_3481,N_2206,N_2942);
xnor U3482 (N_3482,N_2153,N_2197);
nor U3483 (N_3483,N_2113,N_2131);
nor U3484 (N_3484,N_2708,N_2098);
nand U3485 (N_3485,N_2877,N_2218);
and U3486 (N_3486,N_2756,N_2906);
xor U3487 (N_3487,N_2800,N_2626);
and U3488 (N_3488,N_2267,N_2574);
nand U3489 (N_3489,N_2805,N_2941);
nor U3490 (N_3490,N_2481,N_2778);
and U3491 (N_3491,N_2029,N_2219);
nand U3492 (N_3492,N_2959,N_2674);
nand U3493 (N_3493,N_2836,N_2320);
and U3494 (N_3494,N_2615,N_2295);
xor U3495 (N_3495,N_2383,N_2561);
nand U3496 (N_3496,N_2679,N_2420);
or U3497 (N_3497,N_2118,N_2976);
nand U3498 (N_3498,N_2553,N_2682);
and U3499 (N_3499,N_2907,N_2176);
and U3500 (N_3500,N_2644,N_2432);
or U3501 (N_3501,N_2015,N_2787);
xor U3502 (N_3502,N_2185,N_2985);
or U3503 (N_3503,N_2325,N_2381);
nand U3504 (N_3504,N_2339,N_2368);
nor U3505 (N_3505,N_2361,N_2780);
or U3506 (N_3506,N_2052,N_2339);
xnor U3507 (N_3507,N_2657,N_2073);
nor U3508 (N_3508,N_2782,N_2657);
xnor U3509 (N_3509,N_2074,N_2752);
nand U3510 (N_3510,N_2807,N_2130);
nand U3511 (N_3511,N_2521,N_2760);
or U3512 (N_3512,N_2363,N_2253);
xor U3513 (N_3513,N_2891,N_2682);
and U3514 (N_3514,N_2442,N_2668);
or U3515 (N_3515,N_2311,N_2951);
and U3516 (N_3516,N_2294,N_2108);
nand U3517 (N_3517,N_2136,N_2351);
nand U3518 (N_3518,N_2464,N_2021);
xnor U3519 (N_3519,N_2295,N_2301);
and U3520 (N_3520,N_2033,N_2963);
xnor U3521 (N_3521,N_2162,N_2245);
nand U3522 (N_3522,N_2447,N_2002);
and U3523 (N_3523,N_2733,N_2972);
nor U3524 (N_3524,N_2646,N_2229);
nand U3525 (N_3525,N_2968,N_2939);
nor U3526 (N_3526,N_2579,N_2125);
or U3527 (N_3527,N_2357,N_2802);
or U3528 (N_3528,N_2645,N_2200);
nand U3529 (N_3529,N_2203,N_2792);
nor U3530 (N_3530,N_2620,N_2372);
nand U3531 (N_3531,N_2884,N_2223);
and U3532 (N_3532,N_2368,N_2360);
nor U3533 (N_3533,N_2284,N_2814);
xnor U3534 (N_3534,N_2409,N_2640);
xor U3535 (N_3535,N_2350,N_2475);
nor U3536 (N_3536,N_2670,N_2137);
nor U3537 (N_3537,N_2374,N_2678);
xor U3538 (N_3538,N_2074,N_2392);
nor U3539 (N_3539,N_2536,N_2537);
nor U3540 (N_3540,N_2712,N_2501);
and U3541 (N_3541,N_2158,N_2837);
or U3542 (N_3542,N_2056,N_2402);
nor U3543 (N_3543,N_2325,N_2849);
and U3544 (N_3544,N_2599,N_2276);
nor U3545 (N_3545,N_2728,N_2226);
xnor U3546 (N_3546,N_2204,N_2676);
nand U3547 (N_3547,N_2111,N_2058);
nand U3548 (N_3548,N_2144,N_2903);
and U3549 (N_3549,N_2259,N_2440);
or U3550 (N_3550,N_2485,N_2226);
and U3551 (N_3551,N_2064,N_2754);
xor U3552 (N_3552,N_2727,N_2994);
nor U3553 (N_3553,N_2015,N_2359);
or U3554 (N_3554,N_2961,N_2735);
xnor U3555 (N_3555,N_2366,N_2529);
nand U3556 (N_3556,N_2689,N_2086);
nor U3557 (N_3557,N_2339,N_2538);
xor U3558 (N_3558,N_2265,N_2129);
nand U3559 (N_3559,N_2959,N_2942);
nor U3560 (N_3560,N_2006,N_2861);
xor U3561 (N_3561,N_2280,N_2463);
nor U3562 (N_3562,N_2751,N_2556);
or U3563 (N_3563,N_2390,N_2578);
and U3564 (N_3564,N_2887,N_2313);
xnor U3565 (N_3565,N_2246,N_2648);
and U3566 (N_3566,N_2283,N_2822);
nand U3567 (N_3567,N_2738,N_2293);
nor U3568 (N_3568,N_2726,N_2933);
and U3569 (N_3569,N_2880,N_2841);
or U3570 (N_3570,N_2289,N_2909);
or U3571 (N_3571,N_2846,N_2596);
nand U3572 (N_3572,N_2508,N_2633);
nor U3573 (N_3573,N_2410,N_2173);
or U3574 (N_3574,N_2338,N_2263);
nor U3575 (N_3575,N_2166,N_2176);
nand U3576 (N_3576,N_2063,N_2641);
or U3577 (N_3577,N_2977,N_2123);
xnor U3578 (N_3578,N_2101,N_2667);
or U3579 (N_3579,N_2036,N_2271);
xnor U3580 (N_3580,N_2936,N_2095);
nand U3581 (N_3581,N_2202,N_2897);
nand U3582 (N_3582,N_2611,N_2522);
nor U3583 (N_3583,N_2759,N_2072);
and U3584 (N_3584,N_2678,N_2121);
or U3585 (N_3585,N_2483,N_2977);
nand U3586 (N_3586,N_2608,N_2646);
and U3587 (N_3587,N_2721,N_2794);
nand U3588 (N_3588,N_2618,N_2063);
and U3589 (N_3589,N_2026,N_2605);
or U3590 (N_3590,N_2123,N_2508);
nor U3591 (N_3591,N_2635,N_2993);
nand U3592 (N_3592,N_2667,N_2751);
xnor U3593 (N_3593,N_2198,N_2348);
or U3594 (N_3594,N_2292,N_2728);
xnor U3595 (N_3595,N_2547,N_2855);
or U3596 (N_3596,N_2167,N_2981);
xor U3597 (N_3597,N_2293,N_2580);
or U3598 (N_3598,N_2753,N_2880);
nand U3599 (N_3599,N_2959,N_2136);
or U3600 (N_3600,N_2261,N_2705);
and U3601 (N_3601,N_2627,N_2896);
xor U3602 (N_3602,N_2252,N_2051);
and U3603 (N_3603,N_2691,N_2272);
xnor U3604 (N_3604,N_2627,N_2806);
and U3605 (N_3605,N_2603,N_2102);
and U3606 (N_3606,N_2079,N_2656);
nor U3607 (N_3607,N_2528,N_2843);
or U3608 (N_3608,N_2166,N_2629);
nor U3609 (N_3609,N_2648,N_2221);
and U3610 (N_3610,N_2969,N_2735);
nor U3611 (N_3611,N_2355,N_2797);
nor U3612 (N_3612,N_2734,N_2573);
nor U3613 (N_3613,N_2348,N_2302);
or U3614 (N_3614,N_2273,N_2794);
nor U3615 (N_3615,N_2137,N_2366);
nand U3616 (N_3616,N_2996,N_2889);
and U3617 (N_3617,N_2251,N_2484);
nand U3618 (N_3618,N_2861,N_2703);
nand U3619 (N_3619,N_2913,N_2813);
nor U3620 (N_3620,N_2706,N_2398);
nand U3621 (N_3621,N_2776,N_2109);
or U3622 (N_3622,N_2122,N_2124);
xor U3623 (N_3623,N_2661,N_2293);
nor U3624 (N_3624,N_2510,N_2210);
nand U3625 (N_3625,N_2787,N_2438);
nand U3626 (N_3626,N_2807,N_2767);
xor U3627 (N_3627,N_2314,N_2466);
xnor U3628 (N_3628,N_2395,N_2526);
nor U3629 (N_3629,N_2503,N_2708);
or U3630 (N_3630,N_2239,N_2723);
nor U3631 (N_3631,N_2050,N_2030);
nor U3632 (N_3632,N_2616,N_2400);
nor U3633 (N_3633,N_2253,N_2137);
xnor U3634 (N_3634,N_2926,N_2479);
nand U3635 (N_3635,N_2590,N_2278);
nor U3636 (N_3636,N_2702,N_2848);
or U3637 (N_3637,N_2974,N_2563);
nor U3638 (N_3638,N_2046,N_2883);
and U3639 (N_3639,N_2573,N_2551);
xor U3640 (N_3640,N_2842,N_2898);
nor U3641 (N_3641,N_2796,N_2403);
or U3642 (N_3642,N_2347,N_2448);
or U3643 (N_3643,N_2230,N_2234);
xor U3644 (N_3644,N_2611,N_2944);
nor U3645 (N_3645,N_2883,N_2695);
and U3646 (N_3646,N_2414,N_2520);
nand U3647 (N_3647,N_2249,N_2147);
nor U3648 (N_3648,N_2485,N_2091);
xor U3649 (N_3649,N_2454,N_2480);
xnor U3650 (N_3650,N_2490,N_2669);
nand U3651 (N_3651,N_2616,N_2612);
or U3652 (N_3652,N_2001,N_2721);
nand U3653 (N_3653,N_2439,N_2846);
xor U3654 (N_3654,N_2917,N_2277);
and U3655 (N_3655,N_2587,N_2934);
or U3656 (N_3656,N_2421,N_2052);
or U3657 (N_3657,N_2189,N_2749);
xnor U3658 (N_3658,N_2367,N_2266);
nor U3659 (N_3659,N_2103,N_2688);
nand U3660 (N_3660,N_2326,N_2647);
xnor U3661 (N_3661,N_2089,N_2062);
and U3662 (N_3662,N_2669,N_2639);
or U3663 (N_3663,N_2168,N_2954);
or U3664 (N_3664,N_2103,N_2837);
and U3665 (N_3665,N_2811,N_2846);
and U3666 (N_3666,N_2623,N_2958);
nand U3667 (N_3667,N_2602,N_2575);
xor U3668 (N_3668,N_2548,N_2257);
nor U3669 (N_3669,N_2742,N_2533);
or U3670 (N_3670,N_2544,N_2197);
nand U3671 (N_3671,N_2340,N_2706);
or U3672 (N_3672,N_2277,N_2139);
and U3673 (N_3673,N_2872,N_2871);
nand U3674 (N_3674,N_2193,N_2969);
nor U3675 (N_3675,N_2368,N_2776);
xnor U3676 (N_3676,N_2387,N_2064);
xnor U3677 (N_3677,N_2182,N_2832);
or U3678 (N_3678,N_2585,N_2786);
xnor U3679 (N_3679,N_2991,N_2374);
or U3680 (N_3680,N_2871,N_2595);
and U3681 (N_3681,N_2945,N_2548);
nor U3682 (N_3682,N_2870,N_2874);
or U3683 (N_3683,N_2206,N_2087);
or U3684 (N_3684,N_2476,N_2469);
nor U3685 (N_3685,N_2942,N_2748);
xnor U3686 (N_3686,N_2824,N_2677);
or U3687 (N_3687,N_2063,N_2662);
and U3688 (N_3688,N_2836,N_2983);
or U3689 (N_3689,N_2460,N_2296);
or U3690 (N_3690,N_2742,N_2104);
nand U3691 (N_3691,N_2080,N_2028);
nor U3692 (N_3692,N_2568,N_2877);
nor U3693 (N_3693,N_2640,N_2763);
and U3694 (N_3694,N_2641,N_2652);
nor U3695 (N_3695,N_2225,N_2986);
nand U3696 (N_3696,N_2133,N_2776);
xnor U3697 (N_3697,N_2445,N_2894);
nor U3698 (N_3698,N_2616,N_2961);
and U3699 (N_3699,N_2641,N_2840);
or U3700 (N_3700,N_2249,N_2198);
and U3701 (N_3701,N_2335,N_2188);
xnor U3702 (N_3702,N_2382,N_2839);
nor U3703 (N_3703,N_2258,N_2387);
nand U3704 (N_3704,N_2413,N_2773);
and U3705 (N_3705,N_2787,N_2665);
xor U3706 (N_3706,N_2863,N_2668);
xnor U3707 (N_3707,N_2446,N_2525);
nor U3708 (N_3708,N_2940,N_2588);
or U3709 (N_3709,N_2380,N_2566);
xnor U3710 (N_3710,N_2958,N_2720);
nor U3711 (N_3711,N_2607,N_2117);
and U3712 (N_3712,N_2936,N_2645);
nor U3713 (N_3713,N_2365,N_2798);
or U3714 (N_3714,N_2676,N_2094);
xor U3715 (N_3715,N_2018,N_2903);
xor U3716 (N_3716,N_2990,N_2369);
nor U3717 (N_3717,N_2953,N_2815);
nand U3718 (N_3718,N_2958,N_2549);
nand U3719 (N_3719,N_2402,N_2873);
nor U3720 (N_3720,N_2628,N_2047);
xnor U3721 (N_3721,N_2361,N_2956);
and U3722 (N_3722,N_2591,N_2545);
and U3723 (N_3723,N_2287,N_2285);
and U3724 (N_3724,N_2169,N_2244);
nor U3725 (N_3725,N_2381,N_2690);
nand U3726 (N_3726,N_2713,N_2984);
or U3727 (N_3727,N_2234,N_2846);
nand U3728 (N_3728,N_2783,N_2817);
or U3729 (N_3729,N_2557,N_2645);
nor U3730 (N_3730,N_2959,N_2536);
nand U3731 (N_3731,N_2403,N_2993);
nand U3732 (N_3732,N_2247,N_2851);
or U3733 (N_3733,N_2597,N_2448);
nand U3734 (N_3734,N_2206,N_2305);
nand U3735 (N_3735,N_2169,N_2321);
nand U3736 (N_3736,N_2202,N_2376);
nor U3737 (N_3737,N_2415,N_2953);
nand U3738 (N_3738,N_2635,N_2239);
or U3739 (N_3739,N_2800,N_2075);
nor U3740 (N_3740,N_2945,N_2623);
nand U3741 (N_3741,N_2831,N_2691);
and U3742 (N_3742,N_2707,N_2881);
nand U3743 (N_3743,N_2154,N_2197);
nand U3744 (N_3744,N_2708,N_2916);
and U3745 (N_3745,N_2853,N_2955);
nand U3746 (N_3746,N_2799,N_2565);
xor U3747 (N_3747,N_2272,N_2312);
and U3748 (N_3748,N_2994,N_2105);
nand U3749 (N_3749,N_2038,N_2338);
xnor U3750 (N_3750,N_2675,N_2914);
nor U3751 (N_3751,N_2349,N_2597);
nor U3752 (N_3752,N_2116,N_2684);
nor U3753 (N_3753,N_2740,N_2074);
nor U3754 (N_3754,N_2237,N_2350);
and U3755 (N_3755,N_2798,N_2795);
or U3756 (N_3756,N_2622,N_2733);
nor U3757 (N_3757,N_2341,N_2018);
nand U3758 (N_3758,N_2529,N_2260);
or U3759 (N_3759,N_2608,N_2680);
and U3760 (N_3760,N_2185,N_2227);
or U3761 (N_3761,N_2316,N_2181);
nor U3762 (N_3762,N_2008,N_2980);
nor U3763 (N_3763,N_2520,N_2682);
or U3764 (N_3764,N_2193,N_2392);
nor U3765 (N_3765,N_2726,N_2340);
and U3766 (N_3766,N_2216,N_2468);
or U3767 (N_3767,N_2425,N_2716);
nand U3768 (N_3768,N_2880,N_2131);
xnor U3769 (N_3769,N_2153,N_2547);
nand U3770 (N_3770,N_2439,N_2642);
or U3771 (N_3771,N_2412,N_2208);
nor U3772 (N_3772,N_2091,N_2186);
nand U3773 (N_3773,N_2457,N_2873);
nand U3774 (N_3774,N_2412,N_2165);
or U3775 (N_3775,N_2145,N_2822);
nor U3776 (N_3776,N_2616,N_2394);
or U3777 (N_3777,N_2824,N_2688);
and U3778 (N_3778,N_2737,N_2506);
nand U3779 (N_3779,N_2724,N_2033);
and U3780 (N_3780,N_2105,N_2640);
or U3781 (N_3781,N_2689,N_2830);
nand U3782 (N_3782,N_2231,N_2005);
and U3783 (N_3783,N_2573,N_2774);
nand U3784 (N_3784,N_2047,N_2832);
xor U3785 (N_3785,N_2717,N_2579);
nor U3786 (N_3786,N_2531,N_2228);
xor U3787 (N_3787,N_2387,N_2706);
and U3788 (N_3788,N_2612,N_2770);
or U3789 (N_3789,N_2031,N_2614);
nor U3790 (N_3790,N_2165,N_2639);
nand U3791 (N_3791,N_2044,N_2697);
and U3792 (N_3792,N_2305,N_2311);
or U3793 (N_3793,N_2268,N_2537);
and U3794 (N_3794,N_2910,N_2422);
nand U3795 (N_3795,N_2156,N_2482);
and U3796 (N_3796,N_2558,N_2970);
nor U3797 (N_3797,N_2889,N_2225);
or U3798 (N_3798,N_2499,N_2330);
xor U3799 (N_3799,N_2602,N_2142);
and U3800 (N_3800,N_2480,N_2092);
xor U3801 (N_3801,N_2210,N_2886);
nor U3802 (N_3802,N_2422,N_2658);
nand U3803 (N_3803,N_2410,N_2045);
xor U3804 (N_3804,N_2477,N_2704);
xor U3805 (N_3805,N_2189,N_2412);
nor U3806 (N_3806,N_2397,N_2996);
nor U3807 (N_3807,N_2984,N_2104);
xnor U3808 (N_3808,N_2602,N_2382);
nor U3809 (N_3809,N_2646,N_2858);
or U3810 (N_3810,N_2186,N_2633);
nand U3811 (N_3811,N_2026,N_2128);
nand U3812 (N_3812,N_2095,N_2153);
xor U3813 (N_3813,N_2462,N_2974);
nor U3814 (N_3814,N_2947,N_2814);
or U3815 (N_3815,N_2457,N_2785);
nand U3816 (N_3816,N_2495,N_2726);
and U3817 (N_3817,N_2971,N_2020);
xor U3818 (N_3818,N_2015,N_2683);
nor U3819 (N_3819,N_2511,N_2153);
or U3820 (N_3820,N_2798,N_2984);
nand U3821 (N_3821,N_2389,N_2229);
or U3822 (N_3822,N_2402,N_2071);
nor U3823 (N_3823,N_2414,N_2420);
nor U3824 (N_3824,N_2971,N_2212);
xor U3825 (N_3825,N_2844,N_2096);
nand U3826 (N_3826,N_2468,N_2685);
nand U3827 (N_3827,N_2864,N_2886);
nor U3828 (N_3828,N_2785,N_2199);
nand U3829 (N_3829,N_2489,N_2839);
and U3830 (N_3830,N_2776,N_2850);
and U3831 (N_3831,N_2088,N_2121);
nor U3832 (N_3832,N_2621,N_2491);
xnor U3833 (N_3833,N_2374,N_2288);
nand U3834 (N_3834,N_2587,N_2966);
xor U3835 (N_3835,N_2740,N_2208);
nand U3836 (N_3836,N_2656,N_2469);
or U3837 (N_3837,N_2595,N_2737);
xnor U3838 (N_3838,N_2384,N_2465);
and U3839 (N_3839,N_2268,N_2106);
nor U3840 (N_3840,N_2150,N_2058);
and U3841 (N_3841,N_2762,N_2042);
and U3842 (N_3842,N_2408,N_2421);
nor U3843 (N_3843,N_2366,N_2439);
or U3844 (N_3844,N_2073,N_2268);
and U3845 (N_3845,N_2429,N_2470);
xor U3846 (N_3846,N_2525,N_2397);
xor U3847 (N_3847,N_2644,N_2163);
or U3848 (N_3848,N_2261,N_2264);
nand U3849 (N_3849,N_2334,N_2425);
or U3850 (N_3850,N_2514,N_2861);
and U3851 (N_3851,N_2596,N_2501);
nand U3852 (N_3852,N_2901,N_2944);
xor U3853 (N_3853,N_2246,N_2127);
nor U3854 (N_3854,N_2999,N_2621);
and U3855 (N_3855,N_2292,N_2628);
nor U3856 (N_3856,N_2791,N_2894);
or U3857 (N_3857,N_2738,N_2330);
xor U3858 (N_3858,N_2395,N_2971);
or U3859 (N_3859,N_2947,N_2614);
nand U3860 (N_3860,N_2365,N_2741);
or U3861 (N_3861,N_2389,N_2536);
or U3862 (N_3862,N_2835,N_2051);
nand U3863 (N_3863,N_2937,N_2108);
and U3864 (N_3864,N_2692,N_2844);
nand U3865 (N_3865,N_2864,N_2621);
nand U3866 (N_3866,N_2488,N_2808);
nor U3867 (N_3867,N_2182,N_2240);
or U3868 (N_3868,N_2098,N_2160);
nand U3869 (N_3869,N_2957,N_2568);
or U3870 (N_3870,N_2657,N_2034);
and U3871 (N_3871,N_2602,N_2461);
or U3872 (N_3872,N_2170,N_2172);
nand U3873 (N_3873,N_2428,N_2111);
and U3874 (N_3874,N_2373,N_2771);
and U3875 (N_3875,N_2967,N_2113);
nand U3876 (N_3876,N_2160,N_2655);
and U3877 (N_3877,N_2010,N_2394);
xnor U3878 (N_3878,N_2301,N_2702);
or U3879 (N_3879,N_2114,N_2746);
nor U3880 (N_3880,N_2874,N_2079);
and U3881 (N_3881,N_2155,N_2441);
xnor U3882 (N_3882,N_2613,N_2170);
or U3883 (N_3883,N_2002,N_2112);
or U3884 (N_3884,N_2063,N_2070);
or U3885 (N_3885,N_2819,N_2987);
xnor U3886 (N_3886,N_2831,N_2859);
or U3887 (N_3887,N_2075,N_2187);
xor U3888 (N_3888,N_2918,N_2592);
xnor U3889 (N_3889,N_2329,N_2685);
nor U3890 (N_3890,N_2073,N_2127);
and U3891 (N_3891,N_2631,N_2241);
nor U3892 (N_3892,N_2267,N_2998);
nor U3893 (N_3893,N_2762,N_2349);
and U3894 (N_3894,N_2211,N_2782);
nor U3895 (N_3895,N_2661,N_2203);
and U3896 (N_3896,N_2283,N_2338);
xnor U3897 (N_3897,N_2883,N_2497);
and U3898 (N_3898,N_2031,N_2530);
or U3899 (N_3899,N_2733,N_2676);
nor U3900 (N_3900,N_2629,N_2393);
or U3901 (N_3901,N_2725,N_2801);
xor U3902 (N_3902,N_2184,N_2149);
and U3903 (N_3903,N_2149,N_2429);
and U3904 (N_3904,N_2349,N_2744);
nor U3905 (N_3905,N_2634,N_2308);
or U3906 (N_3906,N_2069,N_2922);
nand U3907 (N_3907,N_2633,N_2098);
nor U3908 (N_3908,N_2939,N_2316);
nand U3909 (N_3909,N_2883,N_2078);
or U3910 (N_3910,N_2297,N_2939);
nor U3911 (N_3911,N_2150,N_2916);
or U3912 (N_3912,N_2741,N_2277);
and U3913 (N_3913,N_2520,N_2040);
nand U3914 (N_3914,N_2553,N_2338);
and U3915 (N_3915,N_2066,N_2217);
nand U3916 (N_3916,N_2079,N_2535);
nor U3917 (N_3917,N_2204,N_2236);
or U3918 (N_3918,N_2495,N_2486);
nor U3919 (N_3919,N_2459,N_2959);
nand U3920 (N_3920,N_2202,N_2101);
xor U3921 (N_3921,N_2069,N_2960);
nor U3922 (N_3922,N_2651,N_2347);
nor U3923 (N_3923,N_2208,N_2593);
and U3924 (N_3924,N_2249,N_2431);
nand U3925 (N_3925,N_2405,N_2800);
or U3926 (N_3926,N_2487,N_2378);
xnor U3927 (N_3927,N_2808,N_2178);
or U3928 (N_3928,N_2992,N_2724);
or U3929 (N_3929,N_2048,N_2478);
nor U3930 (N_3930,N_2396,N_2163);
nor U3931 (N_3931,N_2711,N_2174);
or U3932 (N_3932,N_2516,N_2513);
nor U3933 (N_3933,N_2816,N_2760);
nor U3934 (N_3934,N_2610,N_2934);
and U3935 (N_3935,N_2229,N_2713);
nor U3936 (N_3936,N_2689,N_2863);
nor U3937 (N_3937,N_2366,N_2163);
nand U3938 (N_3938,N_2434,N_2085);
xor U3939 (N_3939,N_2861,N_2395);
or U3940 (N_3940,N_2275,N_2611);
or U3941 (N_3941,N_2157,N_2046);
xnor U3942 (N_3942,N_2157,N_2110);
or U3943 (N_3943,N_2387,N_2343);
xor U3944 (N_3944,N_2858,N_2876);
nor U3945 (N_3945,N_2527,N_2290);
xor U3946 (N_3946,N_2337,N_2347);
xor U3947 (N_3947,N_2182,N_2218);
nand U3948 (N_3948,N_2148,N_2774);
xnor U3949 (N_3949,N_2717,N_2968);
nor U3950 (N_3950,N_2701,N_2562);
nand U3951 (N_3951,N_2190,N_2779);
or U3952 (N_3952,N_2858,N_2759);
xor U3953 (N_3953,N_2244,N_2549);
or U3954 (N_3954,N_2596,N_2935);
xor U3955 (N_3955,N_2312,N_2616);
xnor U3956 (N_3956,N_2887,N_2181);
xor U3957 (N_3957,N_2282,N_2831);
nor U3958 (N_3958,N_2179,N_2095);
or U3959 (N_3959,N_2596,N_2480);
nor U3960 (N_3960,N_2997,N_2613);
or U3961 (N_3961,N_2480,N_2577);
or U3962 (N_3962,N_2203,N_2936);
nand U3963 (N_3963,N_2014,N_2368);
nor U3964 (N_3964,N_2898,N_2864);
nor U3965 (N_3965,N_2573,N_2061);
nand U3966 (N_3966,N_2671,N_2461);
and U3967 (N_3967,N_2790,N_2886);
or U3968 (N_3968,N_2504,N_2781);
nand U3969 (N_3969,N_2081,N_2957);
and U3970 (N_3970,N_2143,N_2681);
or U3971 (N_3971,N_2096,N_2498);
nor U3972 (N_3972,N_2243,N_2702);
xnor U3973 (N_3973,N_2640,N_2423);
and U3974 (N_3974,N_2227,N_2223);
nand U3975 (N_3975,N_2465,N_2871);
and U3976 (N_3976,N_2653,N_2296);
nand U3977 (N_3977,N_2171,N_2917);
xnor U3978 (N_3978,N_2038,N_2863);
nand U3979 (N_3979,N_2763,N_2824);
xor U3980 (N_3980,N_2524,N_2287);
and U3981 (N_3981,N_2338,N_2983);
and U3982 (N_3982,N_2382,N_2722);
and U3983 (N_3983,N_2635,N_2561);
xor U3984 (N_3984,N_2963,N_2553);
nand U3985 (N_3985,N_2485,N_2418);
and U3986 (N_3986,N_2897,N_2793);
or U3987 (N_3987,N_2358,N_2600);
nand U3988 (N_3988,N_2445,N_2318);
xnor U3989 (N_3989,N_2867,N_2551);
xor U3990 (N_3990,N_2513,N_2475);
xor U3991 (N_3991,N_2195,N_2468);
or U3992 (N_3992,N_2147,N_2890);
xnor U3993 (N_3993,N_2313,N_2875);
nand U3994 (N_3994,N_2264,N_2743);
and U3995 (N_3995,N_2979,N_2825);
nand U3996 (N_3996,N_2889,N_2810);
xor U3997 (N_3997,N_2113,N_2097);
nor U3998 (N_3998,N_2914,N_2458);
or U3999 (N_3999,N_2978,N_2833);
xor U4000 (N_4000,N_3782,N_3071);
nor U4001 (N_4001,N_3236,N_3392);
and U4002 (N_4002,N_3291,N_3325);
nand U4003 (N_4003,N_3832,N_3190);
nand U4004 (N_4004,N_3666,N_3356);
or U4005 (N_4005,N_3361,N_3111);
xnor U4006 (N_4006,N_3156,N_3309);
or U4007 (N_4007,N_3612,N_3448);
xnor U4008 (N_4008,N_3511,N_3495);
nor U4009 (N_4009,N_3372,N_3390);
xor U4010 (N_4010,N_3409,N_3130);
xnor U4011 (N_4011,N_3177,N_3858);
and U4012 (N_4012,N_3305,N_3730);
or U4013 (N_4013,N_3524,N_3061);
xnor U4014 (N_4014,N_3295,N_3327);
or U4015 (N_4015,N_3480,N_3971);
or U4016 (N_4016,N_3226,N_3041);
and U4017 (N_4017,N_3558,N_3207);
nand U4018 (N_4018,N_3687,N_3778);
xor U4019 (N_4019,N_3455,N_3319);
xor U4020 (N_4020,N_3642,N_3530);
and U4021 (N_4021,N_3186,N_3263);
or U4022 (N_4022,N_3636,N_3969);
and U4023 (N_4023,N_3216,N_3193);
nand U4024 (N_4024,N_3395,N_3746);
and U4025 (N_4025,N_3382,N_3124);
and U4026 (N_4026,N_3814,N_3673);
and U4027 (N_4027,N_3113,N_3279);
or U4028 (N_4028,N_3556,N_3913);
and U4029 (N_4029,N_3608,N_3710);
nor U4030 (N_4030,N_3398,N_3223);
xor U4031 (N_4031,N_3707,N_3030);
and U4032 (N_4032,N_3387,N_3788);
xnor U4033 (N_4033,N_3484,N_3087);
or U4034 (N_4034,N_3347,N_3627);
nor U4035 (N_4035,N_3683,N_3645);
or U4036 (N_4036,N_3354,N_3653);
nand U4037 (N_4037,N_3973,N_3581);
xor U4038 (N_4038,N_3447,N_3757);
nand U4039 (N_4039,N_3097,N_3020);
xnor U4040 (N_4040,N_3035,N_3888);
nand U4041 (N_4041,N_3574,N_3091);
nand U4042 (N_4042,N_3235,N_3275);
nor U4043 (N_4043,N_3902,N_3431);
nand U4044 (N_4044,N_3464,N_3460);
xor U4045 (N_4045,N_3210,N_3352);
or U4046 (N_4046,N_3977,N_3605);
xor U4047 (N_4047,N_3812,N_3432);
and U4048 (N_4048,N_3238,N_3801);
xor U4049 (N_4049,N_3592,N_3090);
or U4050 (N_4050,N_3478,N_3676);
nor U4051 (N_4051,N_3438,N_3895);
nand U4052 (N_4052,N_3657,N_3951);
nand U4053 (N_4053,N_3093,N_3928);
and U4054 (N_4054,N_3709,N_3648);
and U4055 (N_4055,N_3557,N_3878);
xnor U4056 (N_4056,N_3075,N_3215);
nor U4057 (N_4057,N_3899,N_3119);
nor U4058 (N_4058,N_3708,N_3531);
nor U4059 (N_4059,N_3150,N_3400);
nor U4060 (N_4060,N_3954,N_3500);
xor U4061 (N_4061,N_3363,N_3655);
or U4062 (N_4062,N_3674,N_3200);
nor U4063 (N_4063,N_3640,N_3346);
xor U4064 (N_4064,N_3461,N_3960);
or U4065 (N_4065,N_3544,N_3172);
nor U4066 (N_4066,N_3493,N_3918);
nor U4067 (N_4067,N_3519,N_3911);
nand U4068 (N_4068,N_3306,N_3934);
nand U4069 (N_4069,N_3294,N_3479);
nand U4070 (N_4070,N_3595,N_3976);
or U4071 (N_4071,N_3576,N_3842);
and U4072 (N_4072,N_3194,N_3208);
and U4073 (N_4073,N_3085,N_3807);
nand U4074 (N_4074,N_3649,N_3797);
xnor U4075 (N_4075,N_3611,N_3700);
and U4076 (N_4076,N_3885,N_3414);
nand U4077 (N_4077,N_3213,N_3566);
nor U4078 (N_4078,N_3009,N_3247);
xor U4079 (N_4079,N_3007,N_3261);
nand U4080 (N_4080,N_3441,N_3498);
and U4081 (N_4081,N_3251,N_3583);
and U4082 (N_4082,N_3317,N_3989);
xnor U4083 (N_4083,N_3830,N_3063);
xor U4084 (N_4084,N_3910,N_3561);
xor U4085 (N_4085,N_3927,N_3897);
or U4086 (N_4086,N_3922,N_3278);
or U4087 (N_4087,N_3887,N_3909);
xor U4088 (N_4088,N_3879,N_3121);
or U4089 (N_4089,N_3132,N_3394);
nor U4090 (N_4090,N_3517,N_3889);
or U4091 (N_4091,N_3522,N_3758);
xnor U4092 (N_4092,N_3670,N_3234);
and U4093 (N_4093,N_3793,N_3411);
or U4094 (N_4094,N_3751,N_3066);
nand U4095 (N_4095,N_3602,N_3729);
xor U4096 (N_4096,N_3362,N_3231);
xnor U4097 (N_4097,N_3330,N_3287);
or U4098 (N_4098,N_3140,N_3980);
nand U4099 (N_4099,N_3120,N_3932);
and U4100 (N_4100,N_3211,N_3735);
and U4101 (N_4101,N_3148,N_3512);
nand U4102 (N_4102,N_3964,N_3250);
and U4103 (N_4103,N_3665,N_3252);
or U4104 (N_4104,N_3074,N_3824);
or U4105 (N_4105,N_3123,N_3599);
and U4106 (N_4106,N_3738,N_3131);
xor U4107 (N_4107,N_3776,N_3127);
or U4108 (N_4108,N_3326,N_3714);
or U4109 (N_4109,N_3678,N_3525);
or U4110 (N_4110,N_3430,N_3863);
xnor U4111 (N_4111,N_3153,N_3384);
or U4112 (N_4112,N_3618,N_3301);
nand U4113 (N_4113,N_3024,N_3420);
nor U4114 (N_4114,N_3101,N_3022);
nor U4115 (N_4115,N_3129,N_3859);
nor U4116 (N_4116,N_3167,N_3136);
xnor U4117 (N_4117,N_3849,N_3871);
nor U4118 (N_4118,N_3957,N_3039);
nor U4119 (N_4119,N_3984,N_3926);
or U4120 (N_4120,N_3182,N_3571);
and U4121 (N_4121,N_3045,N_3332);
xnor U4122 (N_4122,N_3855,N_3056);
and U4123 (N_4123,N_3241,N_3718);
and U4124 (N_4124,N_3508,N_3552);
or U4125 (N_4125,N_3138,N_3952);
xnor U4126 (N_4126,N_3567,N_3310);
or U4127 (N_4127,N_3162,N_3701);
nor U4128 (N_4128,N_3819,N_3745);
xor U4129 (N_4129,N_3963,N_3497);
or U4130 (N_4130,N_3084,N_3168);
nand U4131 (N_4131,N_3891,N_3388);
xor U4132 (N_4132,N_3137,N_3262);
xor U4133 (N_4133,N_3134,N_3463);
nor U4134 (N_4134,N_3684,N_3652);
or U4135 (N_4135,N_3426,N_3117);
nand U4136 (N_4136,N_3660,N_3866);
nand U4137 (N_4137,N_3869,N_3610);
nand U4138 (N_4138,N_3949,N_3418);
nand U4139 (N_4139,N_3597,N_3465);
nand U4140 (N_4140,N_3505,N_3584);
or U4141 (N_4141,N_3769,N_3504);
or U4142 (N_4142,N_3816,N_3568);
xnor U4143 (N_4143,N_3154,N_3256);
or U4144 (N_4144,N_3621,N_3303);
nand U4145 (N_4145,N_3032,N_3429);
nor U4146 (N_4146,N_3661,N_3339);
or U4147 (N_4147,N_3916,N_3767);
and U4148 (N_4148,N_3092,N_3086);
xnor U4149 (N_4149,N_3001,N_3615);
xor U4150 (N_4150,N_3065,N_3875);
nand U4151 (N_4151,N_3450,N_3125);
or U4152 (N_4152,N_3986,N_3170);
nor U4153 (N_4153,N_3348,N_3004);
nor U4154 (N_4154,N_3218,N_3466);
or U4155 (N_4155,N_3536,N_3834);
nand U4156 (N_4156,N_3790,N_3983);
and U4157 (N_4157,N_3017,N_3861);
nand U4158 (N_4158,N_3375,N_3864);
and U4159 (N_4159,N_3658,N_3237);
nor U4160 (N_4160,N_3192,N_3482);
and U4161 (N_4161,N_3695,N_3492);
and U4162 (N_4162,N_3403,N_3694);
or U4163 (N_4163,N_3924,N_3853);
nand U4164 (N_4164,N_3224,N_3770);
or U4165 (N_4165,N_3644,N_3051);
nor U4166 (N_4166,N_3914,N_3060);
xnor U4167 (N_4167,N_3693,N_3232);
nor U4168 (N_4168,N_3178,N_3506);
nand U4169 (N_4169,N_3547,N_3662);
and U4170 (N_4170,N_3811,N_3639);
xor U4171 (N_4171,N_3635,N_3947);
nor U4172 (N_4172,N_3314,N_3015);
nor U4173 (N_4173,N_3548,N_3383);
and U4174 (N_4174,N_3641,N_3320);
xor U4175 (N_4175,N_3163,N_3365);
or U4176 (N_4176,N_3741,N_3318);
nand U4177 (N_4177,N_3052,N_3095);
xor U4178 (N_4178,N_3836,N_3115);
nor U4179 (N_4179,N_3139,N_3313);
nand U4180 (N_4180,N_3159,N_3764);
xor U4181 (N_4181,N_3302,N_3374);
and U4182 (N_4182,N_3946,N_3582);
xnor U4183 (N_4183,N_3685,N_3399);
xnor U4184 (N_4184,N_3355,N_3591);
or U4185 (N_4185,N_3002,N_3803);
nand U4186 (N_4186,N_3462,N_3854);
xor U4187 (N_4187,N_3029,N_3000);
nand U4188 (N_4188,N_3796,N_3994);
and U4189 (N_4189,N_3122,N_3072);
and U4190 (N_4190,N_3328,N_3189);
or U4191 (N_4191,N_3507,N_3634);
or U4192 (N_4192,N_3412,N_3533);
nor U4193 (N_4193,N_3931,N_3096);
and U4194 (N_4194,N_3098,N_3270);
xnor U4195 (N_4195,N_3335,N_3697);
and U4196 (N_4196,N_3290,N_3838);
and U4197 (N_4197,N_3623,N_3475);
and U4198 (N_4198,N_3702,N_3011);
xnor U4199 (N_4199,N_3083,N_3273);
xnor U4200 (N_4200,N_3883,N_3481);
nand U4201 (N_4201,N_3179,N_3972);
nand U4202 (N_4202,N_3164,N_3006);
or U4203 (N_4203,N_3712,N_3271);
or U4204 (N_4204,N_3619,N_3961);
or U4205 (N_4205,N_3529,N_3276);
nand U4206 (N_4206,N_3981,N_3152);
nor U4207 (N_4207,N_3021,N_3114);
or U4208 (N_4208,N_3606,N_3532);
and U4209 (N_4209,N_3862,N_3806);
nand U4210 (N_4210,N_3690,N_3212);
nor U4211 (N_4211,N_3467,N_3058);
or U4212 (N_4212,N_3732,N_3936);
or U4213 (N_4213,N_3755,N_3026);
or U4214 (N_4214,N_3047,N_3907);
and U4215 (N_4215,N_3825,N_3217);
or U4216 (N_4216,N_3471,N_3473);
xnor U4217 (N_4217,N_3109,N_3756);
nand U4218 (N_4218,N_3381,N_3711);
nand U4219 (N_4219,N_3754,N_3253);
nand U4220 (N_4220,N_3956,N_3600);
or U4221 (N_4221,N_3872,N_3285);
nand U4222 (N_4222,N_3818,N_3573);
xor U4223 (N_4223,N_3353,N_3935);
and U4224 (N_4224,N_3835,N_3637);
and U4225 (N_4225,N_3173,N_3716);
nor U4226 (N_4226,N_3799,N_3297);
and U4227 (N_4227,N_3203,N_3445);
nand U4228 (N_4228,N_3828,N_3982);
and U4229 (N_4229,N_3987,N_3706);
nor U4230 (N_4230,N_3366,N_3717);
and U4231 (N_4231,N_3242,N_3289);
or U4232 (N_4232,N_3555,N_3538);
xnor U4233 (N_4233,N_3100,N_3267);
or U4234 (N_4234,N_3128,N_3821);
nor U4235 (N_4235,N_3791,N_3991);
or U4236 (N_4236,N_3704,N_3449);
nand U4237 (N_4237,N_3542,N_3541);
and U4238 (N_4238,N_3043,N_3938);
nor U4239 (N_4239,N_3378,N_3917);
or U4240 (N_4240,N_3815,N_3359);
and U4241 (N_4241,N_3427,N_3283);
nor U4242 (N_4242,N_3196,N_3458);
nor U4243 (N_4243,N_3488,N_3616);
or U4244 (N_4244,N_3850,N_3787);
and U4245 (N_4245,N_3474,N_3440);
xnor U4246 (N_4246,N_3886,N_3199);
nor U4247 (N_4247,N_3698,N_3721);
and U4248 (N_4248,N_3865,N_3968);
and U4249 (N_4249,N_3201,N_3453);
nand U4250 (N_4250,N_3765,N_3880);
or U4251 (N_4251,N_3527,N_3421);
or U4252 (N_4252,N_3696,N_3733);
nand U4253 (N_4253,N_3244,N_3749);
xor U4254 (N_4254,N_3570,N_3185);
nor U4255 (N_4255,N_3176,N_3350);
and U4256 (N_4256,N_3943,N_3692);
nand U4257 (N_4257,N_3978,N_3559);
or U4258 (N_4258,N_3843,N_3993);
nand U4259 (N_4259,N_3013,N_3870);
and U4260 (N_4260,N_3174,N_3435);
nand U4261 (N_4261,N_3165,N_3245);
xnor U4262 (N_4262,N_3722,N_3903);
xor U4263 (N_4263,N_3079,N_3265);
and U4264 (N_4264,N_3456,N_3070);
or U4265 (N_4265,N_3802,N_3622);
xnor U4266 (N_4266,N_3293,N_3340);
or U4267 (N_4267,N_3341,N_3603);
xor U4268 (N_4268,N_3659,N_3161);
or U4269 (N_4269,N_3739,N_3929);
nand U4270 (N_4270,N_3331,N_3225);
xor U4271 (N_4271,N_3368,N_3728);
nor U4272 (N_4272,N_3997,N_3133);
nand U4273 (N_4273,N_3656,N_3781);
xnor U4274 (N_4274,N_3281,N_3679);
xor U4275 (N_4275,N_3624,N_3094);
xnor U4276 (N_4276,N_3147,N_3876);
nor U4277 (N_4277,N_3930,N_3089);
nand U4278 (N_4278,N_3628,N_3404);
xor U4279 (N_4279,N_3681,N_3151);
nand U4280 (N_4280,N_3672,N_3633);
nor U4281 (N_4281,N_3104,N_3428);
nor U4282 (N_4282,N_3425,N_3537);
nor U4283 (N_4283,N_3073,N_3405);
and U4284 (N_4284,N_3499,N_3436);
nand U4285 (N_4285,N_3112,N_3748);
or U4286 (N_4286,N_3280,N_3925);
nand U4287 (N_4287,N_3753,N_3059);
and U4288 (N_4288,N_3945,N_3491);
xnor U4289 (N_4289,N_3396,N_3025);
or U4290 (N_4290,N_3933,N_3338);
or U4291 (N_4291,N_3446,N_3496);
nor U4292 (N_4292,N_3423,N_3845);
nor U4293 (N_4293,N_3664,N_3078);
nor U4294 (N_4294,N_3406,N_3996);
and U4295 (N_4295,N_3175,N_3663);
and U4296 (N_4296,N_3577,N_3389);
nand U4297 (N_4297,N_3554,N_3364);
xor U4298 (N_4298,N_3324,N_3233);
or U4299 (N_4299,N_3743,N_3116);
and U4300 (N_4300,N_3740,N_3158);
nor U4301 (N_4301,N_3761,N_3485);
or U4302 (N_4302,N_3892,N_3286);
or U4303 (N_4303,N_3343,N_3483);
xor U4304 (N_4304,N_3311,N_3985);
nand U4305 (N_4305,N_3258,N_3638);
nor U4306 (N_4306,N_3171,N_3434);
and U4307 (N_4307,N_3629,N_3080);
or U4308 (N_4308,N_3012,N_3135);
and U4309 (N_4309,N_3470,N_3540);
and U4310 (N_4310,N_3713,N_3048);
xor U4311 (N_4311,N_3691,N_3546);
or U4312 (N_4312,N_3367,N_3974);
and U4313 (N_4313,N_3489,N_3780);
nand U4314 (N_4314,N_3268,N_3249);
xnor U4315 (N_4315,N_3771,N_3370);
nand U4316 (N_4316,N_3920,N_3523);
xor U4317 (N_4317,N_3562,N_3794);
nor U4318 (N_4318,N_3626,N_3565);
xor U4319 (N_4319,N_3774,N_3351);
xnor U4320 (N_4320,N_3514,N_3564);
nand U4321 (N_4321,N_3839,N_3654);
nor U4322 (N_4322,N_3786,N_3415);
and U4323 (N_4323,N_3940,N_3349);
or U4324 (N_4324,N_3316,N_3376);
nand U4325 (N_4325,N_3579,N_3601);
nor U4326 (N_4326,N_3358,N_3408);
or U4327 (N_4327,N_3593,N_3014);
nor U4328 (N_4328,N_3857,N_3155);
or U4329 (N_4329,N_3823,N_3220);
and U4330 (N_4330,N_3195,N_3939);
xor U4331 (N_4331,N_3468,N_3292);
nand U4332 (N_4332,N_3028,N_3742);
nor U4333 (N_4333,N_3912,N_3944);
or U4334 (N_4334,N_3360,N_3110);
nand U4335 (N_4335,N_3018,N_3345);
and U4336 (N_4336,N_3402,N_3334);
nand U4337 (N_4337,N_3336,N_3469);
nand U4338 (N_4338,N_3810,N_3841);
nand U4339 (N_4339,N_3008,N_3760);
and U4340 (N_4340,N_3037,N_3321);
nand U4341 (N_4341,N_3904,N_3424);
or U4342 (N_4342,N_3143,N_3342);
or U4343 (N_4343,N_3631,N_3221);
xor U4344 (N_4344,N_3900,N_3580);
or U4345 (N_4345,N_3766,N_3257);
nor U4346 (N_4346,N_3792,N_3181);
xnor U4347 (N_4347,N_3042,N_3490);
nand U4348 (N_4348,N_3569,N_3118);
nand U4349 (N_4349,N_3442,N_3894);
nand U4350 (N_4350,N_3979,N_3304);
nand U4351 (N_4351,N_3477,N_3784);
or U4352 (N_4352,N_3607,N_3369);
nand U4353 (N_4353,N_3759,N_3344);
nand U4354 (N_4354,N_3789,N_3397);
and U4355 (N_4355,N_3027,N_3202);
or U4356 (N_4356,N_3501,N_3723);
nor U4357 (N_4357,N_3590,N_3703);
or U4358 (N_4358,N_3046,N_3563);
nor U4359 (N_4359,N_3813,N_3534);
and U4360 (N_4360,N_3598,N_3433);
xnor U4361 (N_4361,N_3169,N_3827);
xor U4362 (N_4362,N_3543,N_3785);
xor U4363 (N_4363,N_3959,N_3053);
xor U4364 (N_4364,N_3617,N_3630);
nor U4365 (N_4365,N_3844,N_3166);
and U4366 (N_4366,N_3919,N_3572);
and U4367 (N_4367,N_3783,N_3243);
nor U4368 (N_4368,N_3588,N_3768);
nor U4369 (N_4369,N_3596,N_3105);
nor U4370 (N_4370,N_3609,N_3373);
and U4371 (N_4371,N_3259,N_3229);
nand U4372 (N_4372,N_3444,N_3209);
or U4373 (N_4373,N_3264,N_3724);
nand U4374 (N_4374,N_3647,N_3545);
and U4375 (N_4375,N_3103,N_3955);
nand U4376 (N_4376,N_3833,N_3874);
nand U4377 (N_4377,N_3064,N_3820);
nor U4378 (N_4378,N_3144,N_3575);
nand U4379 (N_4379,N_3898,N_3915);
xor U4380 (N_4380,N_3050,N_3081);
xnor U4381 (N_4381,N_3371,N_3068);
xnor U4382 (N_4382,N_3416,N_3551);
nand U4383 (N_4383,N_3266,N_3023);
nand U4384 (N_4384,N_3108,N_3705);
nand U4385 (N_4385,N_3476,N_3443);
and U4386 (N_4386,N_3230,N_3227);
and U4387 (N_4387,N_3298,N_3417);
nand U4388 (N_4388,N_3160,N_3107);
or U4389 (N_4389,N_3494,N_3808);
or U4390 (N_4390,N_3720,N_3183);
nand U4391 (N_4391,N_3950,N_3521);
and U4392 (N_4392,N_3272,N_3099);
nand U4393 (N_4393,N_3502,N_3868);
and U4394 (N_4394,N_3312,N_3995);
and U4395 (N_4395,N_3255,N_3401);
xor U4396 (N_4396,N_3419,N_3958);
xor U4397 (N_4397,N_3187,N_3604);
nand U4398 (N_4398,N_3386,N_3379);
and U4399 (N_4399,N_3049,N_3962);
and U4400 (N_4400,N_3437,N_3391);
xnor U4401 (N_4401,N_3675,N_3809);
nand U4402 (N_4402,N_3333,N_3539);
nor U4403 (N_4403,N_3549,N_3214);
nand U4404 (N_4404,N_3699,N_3804);
and U4405 (N_4405,N_3688,N_3965);
nor U4406 (N_4406,N_3667,N_3518);
nand U4407 (N_4407,N_3222,N_3614);
nand U4408 (N_4408,N_3680,N_3677);
nor U4409 (N_4409,N_3439,N_3747);
nor U4410 (N_4410,N_3848,N_3454);
xor U4411 (N_4411,N_3077,N_3385);
and U4412 (N_4412,N_3805,N_3323);
nor U4413 (N_4413,N_3003,N_3254);
nand U4414 (N_4414,N_3744,N_3998);
nand U4415 (N_4415,N_3413,N_3036);
or U4416 (N_4416,N_3239,N_3589);
nor U4417 (N_4417,N_3033,N_3487);
xor U4418 (N_4418,N_3831,N_3142);
or U4419 (N_4419,N_3750,N_3779);
or U4420 (N_4420,N_3288,N_3921);
nand U4421 (N_4421,N_3393,N_3906);
nor U4422 (N_4422,N_3777,N_3851);
nor U4423 (N_4423,N_3197,N_3513);
xnor U4424 (N_4424,N_3520,N_3860);
nor U4425 (N_4425,N_3451,N_3578);
or U4426 (N_4426,N_3205,N_3005);
xor U4427 (N_4427,N_3069,N_3516);
or U4428 (N_4428,N_3715,N_3184);
and U4429 (N_4429,N_3410,N_3669);
xor U4430 (N_4430,N_3550,N_3877);
or U4431 (N_4431,N_3795,N_3737);
nor U4432 (N_4432,N_3054,N_3299);
nand U4433 (N_4433,N_3204,N_3689);
or U4434 (N_4434,N_3646,N_3515);
xnor U4435 (N_4435,N_3322,N_3937);
and U4436 (N_4436,N_3031,N_3126);
and U4437 (N_4437,N_3826,N_3719);
and U4438 (N_4438,N_3731,N_3948);
nand U4439 (N_4439,N_3062,N_3248);
nand U4440 (N_4440,N_3308,N_3300);
and U4441 (N_4441,N_3736,N_3867);
and U4442 (N_4442,N_3613,N_3510);
nor U4443 (N_4443,N_3509,N_3503);
or U4444 (N_4444,N_3587,N_3188);
nor U4445 (N_4445,N_3157,N_3457);
nor U4446 (N_4446,N_3822,N_3725);
and U4447 (N_4447,N_3992,N_3852);
nand U4448 (N_4448,N_3422,N_3752);
and U4449 (N_4449,N_3274,N_3191);
and U4450 (N_4450,N_3970,N_3873);
nand U4451 (N_4451,N_3942,N_3219);
nand U4452 (N_4452,N_3727,N_3890);
nor U4453 (N_4453,N_3817,N_3010);
nand U4454 (N_4454,N_3553,N_3882);
xnor U4455 (N_4455,N_3452,N_3459);
or U4456 (N_4456,N_3620,N_3472);
and U4457 (N_4457,N_3038,N_3967);
and U4458 (N_4458,N_3180,N_3076);
or U4459 (N_4459,N_3145,N_3284);
nor U4460 (N_4460,N_3893,N_3668);
nand U4461 (N_4461,N_3019,N_3651);
and U4462 (N_4462,N_3040,N_3526);
or U4463 (N_4463,N_3632,N_3560);
nor U4464 (N_4464,N_3240,N_3277);
xnor U4465 (N_4465,N_3856,N_3198);
xor U4466 (N_4466,N_3763,N_3941);
xor U4467 (N_4467,N_3905,N_3034);
nor U4468 (N_4468,N_3228,N_3775);
nor U4469 (N_4469,N_3988,N_3141);
or U4470 (N_4470,N_3643,N_3528);
xnor U4471 (N_4471,N_3896,N_3269);
xnor U4472 (N_4472,N_3847,N_3057);
xnor U4473 (N_4473,N_3535,N_3486);
nor U4474 (N_4474,N_3975,N_3734);
nor U4475 (N_4475,N_3044,N_3106);
and U4476 (N_4476,N_3773,N_3686);
or U4477 (N_4477,N_3357,N_3246);
or U4478 (N_4478,N_3908,N_3594);
xor U4479 (N_4479,N_3102,N_3282);
nand U4480 (N_4480,N_3881,N_3650);
nor U4481 (N_4481,N_3923,N_3296);
nand U4482 (N_4482,N_3082,N_3884);
or U4483 (N_4483,N_3016,N_3671);
nor U4484 (N_4484,N_3772,N_3055);
nor U4485 (N_4485,N_3315,N_3337);
or U4486 (N_4486,N_3682,N_3800);
or U4487 (N_4487,N_3149,N_3586);
and U4488 (N_4488,N_3585,N_3966);
nand U4489 (N_4489,N_3377,N_3798);
and U4490 (N_4490,N_3260,N_3067);
or U4491 (N_4491,N_3762,N_3726);
xor U4492 (N_4492,N_3990,N_3840);
nand U4493 (N_4493,N_3146,N_3088);
nor U4494 (N_4494,N_3829,N_3329);
xnor U4495 (N_4495,N_3837,N_3206);
nor U4496 (N_4496,N_3846,N_3380);
xor U4497 (N_4497,N_3307,N_3953);
nor U4498 (N_4498,N_3625,N_3407);
and U4499 (N_4499,N_3999,N_3901);
xnor U4500 (N_4500,N_3364,N_3132);
or U4501 (N_4501,N_3540,N_3661);
or U4502 (N_4502,N_3978,N_3353);
or U4503 (N_4503,N_3821,N_3107);
or U4504 (N_4504,N_3287,N_3630);
and U4505 (N_4505,N_3868,N_3093);
nand U4506 (N_4506,N_3482,N_3208);
and U4507 (N_4507,N_3061,N_3715);
and U4508 (N_4508,N_3595,N_3858);
or U4509 (N_4509,N_3957,N_3977);
xor U4510 (N_4510,N_3919,N_3459);
xnor U4511 (N_4511,N_3098,N_3737);
nor U4512 (N_4512,N_3526,N_3025);
and U4513 (N_4513,N_3925,N_3024);
xor U4514 (N_4514,N_3847,N_3146);
xnor U4515 (N_4515,N_3444,N_3805);
nor U4516 (N_4516,N_3810,N_3144);
xor U4517 (N_4517,N_3528,N_3604);
nand U4518 (N_4518,N_3836,N_3204);
nand U4519 (N_4519,N_3051,N_3203);
nor U4520 (N_4520,N_3259,N_3363);
nand U4521 (N_4521,N_3594,N_3469);
or U4522 (N_4522,N_3831,N_3991);
or U4523 (N_4523,N_3313,N_3362);
nand U4524 (N_4524,N_3347,N_3940);
xnor U4525 (N_4525,N_3326,N_3217);
or U4526 (N_4526,N_3111,N_3426);
xnor U4527 (N_4527,N_3128,N_3033);
xnor U4528 (N_4528,N_3828,N_3336);
and U4529 (N_4529,N_3820,N_3637);
nand U4530 (N_4530,N_3530,N_3677);
nor U4531 (N_4531,N_3852,N_3416);
and U4532 (N_4532,N_3109,N_3425);
xnor U4533 (N_4533,N_3589,N_3775);
and U4534 (N_4534,N_3228,N_3477);
nor U4535 (N_4535,N_3994,N_3952);
and U4536 (N_4536,N_3682,N_3241);
nor U4537 (N_4537,N_3206,N_3829);
xnor U4538 (N_4538,N_3867,N_3473);
nand U4539 (N_4539,N_3151,N_3570);
and U4540 (N_4540,N_3230,N_3374);
and U4541 (N_4541,N_3162,N_3393);
xor U4542 (N_4542,N_3148,N_3395);
nor U4543 (N_4543,N_3097,N_3240);
or U4544 (N_4544,N_3214,N_3254);
nand U4545 (N_4545,N_3397,N_3135);
xnor U4546 (N_4546,N_3924,N_3326);
xor U4547 (N_4547,N_3198,N_3330);
xnor U4548 (N_4548,N_3702,N_3518);
xnor U4549 (N_4549,N_3066,N_3775);
nor U4550 (N_4550,N_3684,N_3337);
nor U4551 (N_4551,N_3073,N_3543);
xor U4552 (N_4552,N_3522,N_3295);
or U4553 (N_4553,N_3578,N_3645);
and U4554 (N_4554,N_3534,N_3006);
or U4555 (N_4555,N_3098,N_3458);
xor U4556 (N_4556,N_3552,N_3240);
nand U4557 (N_4557,N_3385,N_3347);
xor U4558 (N_4558,N_3194,N_3327);
and U4559 (N_4559,N_3269,N_3362);
and U4560 (N_4560,N_3693,N_3911);
nand U4561 (N_4561,N_3728,N_3954);
or U4562 (N_4562,N_3967,N_3135);
and U4563 (N_4563,N_3449,N_3293);
nand U4564 (N_4564,N_3301,N_3549);
nor U4565 (N_4565,N_3184,N_3201);
or U4566 (N_4566,N_3397,N_3571);
and U4567 (N_4567,N_3461,N_3908);
nor U4568 (N_4568,N_3859,N_3902);
xnor U4569 (N_4569,N_3912,N_3322);
nand U4570 (N_4570,N_3695,N_3560);
and U4571 (N_4571,N_3951,N_3445);
xnor U4572 (N_4572,N_3183,N_3819);
xnor U4573 (N_4573,N_3974,N_3487);
and U4574 (N_4574,N_3386,N_3909);
and U4575 (N_4575,N_3010,N_3936);
xnor U4576 (N_4576,N_3011,N_3755);
and U4577 (N_4577,N_3709,N_3007);
nand U4578 (N_4578,N_3038,N_3758);
xnor U4579 (N_4579,N_3055,N_3603);
nor U4580 (N_4580,N_3356,N_3769);
nor U4581 (N_4581,N_3937,N_3670);
xor U4582 (N_4582,N_3554,N_3546);
and U4583 (N_4583,N_3641,N_3387);
nor U4584 (N_4584,N_3077,N_3372);
nand U4585 (N_4585,N_3299,N_3635);
nand U4586 (N_4586,N_3422,N_3434);
xor U4587 (N_4587,N_3292,N_3287);
xnor U4588 (N_4588,N_3935,N_3085);
or U4589 (N_4589,N_3291,N_3553);
or U4590 (N_4590,N_3036,N_3932);
or U4591 (N_4591,N_3908,N_3759);
nor U4592 (N_4592,N_3437,N_3420);
or U4593 (N_4593,N_3345,N_3608);
nand U4594 (N_4594,N_3918,N_3062);
xor U4595 (N_4595,N_3196,N_3975);
xnor U4596 (N_4596,N_3649,N_3652);
nand U4597 (N_4597,N_3092,N_3858);
xnor U4598 (N_4598,N_3917,N_3692);
nand U4599 (N_4599,N_3557,N_3695);
xor U4600 (N_4600,N_3680,N_3771);
nor U4601 (N_4601,N_3028,N_3928);
nand U4602 (N_4602,N_3830,N_3734);
nor U4603 (N_4603,N_3011,N_3701);
or U4604 (N_4604,N_3813,N_3348);
nor U4605 (N_4605,N_3820,N_3365);
and U4606 (N_4606,N_3516,N_3118);
or U4607 (N_4607,N_3288,N_3354);
and U4608 (N_4608,N_3491,N_3004);
nor U4609 (N_4609,N_3078,N_3290);
nand U4610 (N_4610,N_3738,N_3262);
xnor U4611 (N_4611,N_3367,N_3818);
xor U4612 (N_4612,N_3113,N_3233);
nor U4613 (N_4613,N_3985,N_3629);
or U4614 (N_4614,N_3040,N_3510);
xnor U4615 (N_4615,N_3033,N_3130);
and U4616 (N_4616,N_3047,N_3271);
nor U4617 (N_4617,N_3987,N_3461);
nand U4618 (N_4618,N_3936,N_3662);
or U4619 (N_4619,N_3855,N_3876);
nor U4620 (N_4620,N_3588,N_3837);
nand U4621 (N_4621,N_3201,N_3385);
nand U4622 (N_4622,N_3883,N_3185);
and U4623 (N_4623,N_3784,N_3567);
and U4624 (N_4624,N_3682,N_3167);
and U4625 (N_4625,N_3996,N_3498);
xor U4626 (N_4626,N_3871,N_3719);
nand U4627 (N_4627,N_3368,N_3076);
or U4628 (N_4628,N_3723,N_3329);
and U4629 (N_4629,N_3754,N_3613);
and U4630 (N_4630,N_3906,N_3901);
xor U4631 (N_4631,N_3325,N_3562);
nor U4632 (N_4632,N_3750,N_3578);
and U4633 (N_4633,N_3312,N_3020);
nand U4634 (N_4634,N_3856,N_3620);
nor U4635 (N_4635,N_3121,N_3680);
nand U4636 (N_4636,N_3722,N_3009);
xor U4637 (N_4637,N_3002,N_3960);
or U4638 (N_4638,N_3595,N_3583);
and U4639 (N_4639,N_3555,N_3788);
nor U4640 (N_4640,N_3890,N_3290);
or U4641 (N_4641,N_3008,N_3868);
nor U4642 (N_4642,N_3765,N_3978);
nor U4643 (N_4643,N_3813,N_3002);
nor U4644 (N_4644,N_3743,N_3522);
nor U4645 (N_4645,N_3856,N_3593);
nor U4646 (N_4646,N_3328,N_3430);
or U4647 (N_4647,N_3068,N_3174);
nor U4648 (N_4648,N_3786,N_3445);
and U4649 (N_4649,N_3318,N_3903);
or U4650 (N_4650,N_3041,N_3261);
nand U4651 (N_4651,N_3411,N_3879);
xnor U4652 (N_4652,N_3596,N_3077);
or U4653 (N_4653,N_3507,N_3071);
nand U4654 (N_4654,N_3825,N_3868);
nand U4655 (N_4655,N_3919,N_3341);
and U4656 (N_4656,N_3914,N_3055);
nand U4657 (N_4657,N_3770,N_3301);
nand U4658 (N_4658,N_3972,N_3168);
and U4659 (N_4659,N_3560,N_3583);
xor U4660 (N_4660,N_3142,N_3684);
xnor U4661 (N_4661,N_3394,N_3081);
nor U4662 (N_4662,N_3499,N_3590);
xnor U4663 (N_4663,N_3501,N_3775);
and U4664 (N_4664,N_3330,N_3012);
and U4665 (N_4665,N_3762,N_3290);
nand U4666 (N_4666,N_3032,N_3979);
and U4667 (N_4667,N_3931,N_3437);
nand U4668 (N_4668,N_3047,N_3355);
nand U4669 (N_4669,N_3864,N_3380);
and U4670 (N_4670,N_3769,N_3475);
xor U4671 (N_4671,N_3981,N_3600);
xnor U4672 (N_4672,N_3006,N_3559);
xnor U4673 (N_4673,N_3478,N_3933);
xnor U4674 (N_4674,N_3243,N_3025);
xnor U4675 (N_4675,N_3017,N_3224);
nor U4676 (N_4676,N_3157,N_3063);
and U4677 (N_4677,N_3145,N_3759);
nor U4678 (N_4678,N_3714,N_3917);
nand U4679 (N_4679,N_3313,N_3566);
nand U4680 (N_4680,N_3127,N_3301);
or U4681 (N_4681,N_3261,N_3744);
and U4682 (N_4682,N_3792,N_3847);
nor U4683 (N_4683,N_3405,N_3246);
and U4684 (N_4684,N_3696,N_3616);
or U4685 (N_4685,N_3629,N_3075);
or U4686 (N_4686,N_3843,N_3940);
and U4687 (N_4687,N_3593,N_3752);
and U4688 (N_4688,N_3324,N_3612);
nand U4689 (N_4689,N_3568,N_3173);
and U4690 (N_4690,N_3717,N_3293);
nand U4691 (N_4691,N_3572,N_3030);
xor U4692 (N_4692,N_3836,N_3664);
nand U4693 (N_4693,N_3683,N_3047);
xnor U4694 (N_4694,N_3084,N_3654);
and U4695 (N_4695,N_3982,N_3890);
xnor U4696 (N_4696,N_3468,N_3682);
or U4697 (N_4697,N_3255,N_3073);
nand U4698 (N_4698,N_3953,N_3496);
and U4699 (N_4699,N_3270,N_3908);
nand U4700 (N_4700,N_3736,N_3279);
or U4701 (N_4701,N_3697,N_3470);
and U4702 (N_4702,N_3687,N_3681);
xnor U4703 (N_4703,N_3190,N_3333);
xor U4704 (N_4704,N_3723,N_3688);
nand U4705 (N_4705,N_3459,N_3651);
or U4706 (N_4706,N_3825,N_3689);
nand U4707 (N_4707,N_3959,N_3853);
or U4708 (N_4708,N_3366,N_3177);
nand U4709 (N_4709,N_3712,N_3190);
nand U4710 (N_4710,N_3497,N_3670);
nand U4711 (N_4711,N_3123,N_3975);
and U4712 (N_4712,N_3391,N_3031);
or U4713 (N_4713,N_3757,N_3400);
and U4714 (N_4714,N_3568,N_3706);
or U4715 (N_4715,N_3487,N_3464);
and U4716 (N_4716,N_3170,N_3547);
or U4717 (N_4717,N_3602,N_3779);
nor U4718 (N_4718,N_3180,N_3773);
nor U4719 (N_4719,N_3501,N_3828);
nand U4720 (N_4720,N_3549,N_3060);
nand U4721 (N_4721,N_3207,N_3990);
nand U4722 (N_4722,N_3603,N_3161);
or U4723 (N_4723,N_3804,N_3074);
xor U4724 (N_4724,N_3196,N_3525);
or U4725 (N_4725,N_3565,N_3155);
and U4726 (N_4726,N_3103,N_3959);
nor U4727 (N_4727,N_3564,N_3273);
and U4728 (N_4728,N_3857,N_3532);
xor U4729 (N_4729,N_3597,N_3813);
nor U4730 (N_4730,N_3350,N_3388);
or U4731 (N_4731,N_3188,N_3244);
and U4732 (N_4732,N_3568,N_3710);
or U4733 (N_4733,N_3901,N_3977);
nor U4734 (N_4734,N_3072,N_3102);
or U4735 (N_4735,N_3677,N_3381);
xor U4736 (N_4736,N_3757,N_3286);
xnor U4737 (N_4737,N_3849,N_3722);
nor U4738 (N_4738,N_3731,N_3261);
nor U4739 (N_4739,N_3580,N_3645);
or U4740 (N_4740,N_3779,N_3805);
or U4741 (N_4741,N_3515,N_3743);
and U4742 (N_4742,N_3686,N_3230);
xnor U4743 (N_4743,N_3277,N_3151);
nand U4744 (N_4744,N_3107,N_3052);
nor U4745 (N_4745,N_3777,N_3147);
and U4746 (N_4746,N_3383,N_3064);
nand U4747 (N_4747,N_3049,N_3294);
nor U4748 (N_4748,N_3926,N_3731);
or U4749 (N_4749,N_3477,N_3904);
nor U4750 (N_4750,N_3564,N_3602);
nand U4751 (N_4751,N_3825,N_3759);
xnor U4752 (N_4752,N_3988,N_3916);
or U4753 (N_4753,N_3811,N_3418);
nor U4754 (N_4754,N_3646,N_3393);
and U4755 (N_4755,N_3373,N_3126);
and U4756 (N_4756,N_3639,N_3162);
nand U4757 (N_4757,N_3157,N_3559);
or U4758 (N_4758,N_3982,N_3478);
xor U4759 (N_4759,N_3794,N_3527);
nor U4760 (N_4760,N_3106,N_3261);
xnor U4761 (N_4761,N_3676,N_3846);
xnor U4762 (N_4762,N_3349,N_3855);
and U4763 (N_4763,N_3019,N_3928);
and U4764 (N_4764,N_3284,N_3153);
or U4765 (N_4765,N_3214,N_3985);
or U4766 (N_4766,N_3262,N_3344);
nand U4767 (N_4767,N_3241,N_3631);
or U4768 (N_4768,N_3534,N_3234);
nor U4769 (N_4769,N_3009,N_3117);
nor U4770 (N_4770,N_3110,N_3774);
and U4771 (N_4771,N_3101,N_3957);
nor U4772 (N_4772,N_3897,N_3788);
nor U4773 (N_4773,N_3613,N_3390);
xor U4774 (N_4774,N_3551,N_3469);
xor U4775 (N_4775,N_3375,N_3329);
nand U4776 (N_4776,N_3382,N_3892);
nand U4777 (N_4777,N_3791,N_3391);
or U4778 (N_4778,N_3127,N_3467);
nor U4779 (N_4779,N_3146,N_3892);
nand U4780 (N_4780,N_3364,N_3685);
and U4781 (N_4781,N_3362,N_3684);
or U4782 (N_4782,N_3449,N_3709);
nand U4783 (N_4783,N_3424,N_3969);
xor U4784 (N_4784,N_3841,N_3183);
nor U4785 (N_4785,N_3987,N_3974);
nor U4786 (N_4786,N_3431,N_3794);
nand U4787 (N_4787,N_3452,N_3191);
nor U4788 (N_4788,N_3170,N_3246);
xnor U4789 (N_4789,N_3375,N_3430);
xnor U4790 (N_4790,N_3239,N_3702);
or U4791 (N_4791,N_3529,N_3497);
and U4792 (N_4792,N_3259,N_3169);
and U4793 (N_4793,N_3756,N_3188);
and U4794 (N_4794,N_3298,N_3437);
nor U4795 (N_4795,N_3100,N_3008);
nand U4796 (N_4796,N_3140,N_3202);
or U4797 (N_4797,N_3456,N_3276);
xnor U4798 (N_4798,N_3863,N_3824);
xor U4799 (N_4799,N_3083,N_3356);
xnor U4800 (N_4800,N_3542,N_3438);
or U4801 (N_4801,N_3709,N_3771);
nor U4802 (N_4802,N_3391,N_3986);
nand U4803 (N_4803,N_3199,N_3117);
nor U4804 (N_4804,N_3463,N_3200);
nand U4805 (N_4805,N_3425,N_3855);
xor U4806 (N_4806,N_3492,N_3474);
and U4807 (N_4807,N_3819,N_3471);
nand U4808 (N_4808,N_3843,N_3933);
nor U4809 (N_4809,N_3301,N_3530);
xor U4810 (N_4810,N_3571,N_3905);
and U4811 (N_4811,N_3726,N_3678);
or U4812 (N_4812,N_3593,N_3919);
xnor U4813 (N_4813,N_3975,N_3426);
nand U4814 (N_4814,N_3691,N_3982);
or U4815 (N_4815,N_3540,N_3736);
or U4816 (N_4816,N_3871,N_3259);
and U4817 (N_4817,N_3402,N_3475);
nand U4818 (N_4818,N_3268,N_3627);
xnor U4819 (N_4819,N_3266,N_3115);
or U4820 (N_4820,N_3789,N_3222);
and U4821 (N_4821,N_3828,N_3275);
or U4822 (N_4822,N_3979,N_3630);
xnor U4823 (N_4823,N_3652,N_3499);
nand U4824 (N_4824,N_3546,N_3653);
xor U4825 (N_4825,N_3439,N_3695);
xor U4826 (N_4826,N_3751,N_3908);
nand U4827 (N_4827,N_3672,N_3514);
nand U4828 (N_4828,N_3570,N_3395);
xor U4829 (N_4829,N_3054,N_3355);
nand U4830 (N_4830,N_3546,N_3069);
xnor U4831 (N_4831,N_3111,N_3225);
or U4832 (N_4832,N_3530,N_3449);
and U4833 (N_4833,N_3470,N_3002);
nand U4834 (N_4834,N_3012,N_3112);
nand U4835 (N_4835,N_3188,N_3931);
nand U4836 (N_4836,N_3404,N_3903);
or U4837 (N_4837,N_3221,N_3318);
and U4838 (N_4838,N_3309,N_3382);
xor U4839 (N_4839,N_3473,N_3273);
or U4840 (N_4840,N_3001,N_3211);
nand U4841 (N_4841,N_3374,N_3720);
nor U4842 (N_4842,N_3424,N_3736);
and U4843 (N_4843,N_3348,N_3173);
or U4844 (N_4844,N_3005,N_3318);
nand U4845 (N_4845,N_3729,N_3692);
nor U4846 (N_4846,N_3050,N_3676);
or U4847 (N_4847,N_3324,N_3465);
or U4848 (N_4848,N_3238,N_3487);
or U4849 (N_4849,N_3599,N_3946);
and U4850 (N_4850,N_3281,N_3875);
nand U4851 (N_4851,N_3972,N_3324);
xor U4852 (N_4852,N_3429,N_3687);
nor U4853 (N_4853,N_3401,N_3031);
xor U4854 (N_4854,N_3163,N_3573);
nand U4855 (N_4855,N_3295,N_3637);
nand U4856 (N_4856,N_3371,N_3221);
nand U4857 (N_4857,N_3182,N_3619);
nand U4858 (N_4858,N_3835,N_3327);
nor U4859 (N_4859,N_3695,N_3541);
or U4860 (N_4860,N_3657,N_3443);
nor U4861 (N_4861,N_3301,N_3423);
or U4862 (N_4862,N_3261,N_3732);
and U4863 (N_4863,N_3429,N_3394);
or U4864 (N_4864,N_3891,N_3386);
nor U4865 (N_4865,N_3397,N_3707);
nor U4866 (N_4866,N_3023,N_3215);
nor U4867 (N_4867,N_3235,N_3754);
and U4868 (N_4868,N_3358,N_3766);
and U4869 (N_4869,N_3679,N_3228);
xnor U4870 (N_4870,N_3929,N_3662);
and U4871 (N_4871,N_3543,N_3324);
nand U4872 (N_4872,N_3956,N_3091);
nand U4873 (N_4873,N_3765,N_3739);
or U4874 (N_4874,N_3805,N_3884);
and U4875 (N_4875,N_3388,N_3101);
and U4876 (N_4876,N_3557,N_3271);
or U4877 (N_4877,N_3770,N_3678);
and U4878 (N_4878,N_3559,N_3189);
and U4879 (N_4879,N_3213,N_3259);
xnor U4880 (N_4880,N_3501,N_3803);
and U4881 (N_4881,N_3491,N_3310);
xnor U4882 (N_4882,N_3081,N_3464);
xnor U4883 (N_4883,N_3092,N_3979);
nand U4884 (N_4884,N_3777,N_3784);
and U4885 (N_4885,N_3702,N_3635);
and U4886 (N_4886,N_3106,N_3181);
and U4887 (N_4887,N_3098,N_3005);
xnor U4888 (N_4888,N_3568,N_3835);
nor U4889 (N_4889,N_3652,N_3651);
and U4890 (N_4890,N_3164,N_3620);
nand U4891 (N_4891,N_3845,N_3957);
nand U4892 (N_4892,N_3365,N_3501);
xnor U4893 (N_4893,N_3879,N_3972);
nor U4894 (N_4894,N_3594,N_3635);
or U4895 (N_4895,N_3269,N_3557);
and U4896 (N_4896,N_3219,N_3515);
and U4897 (N_4897,N_3885,N_3942);
xnor U4898 (N_4898,N_3845,N_3962);
or U4899 (N_4899,N_3543,N_3342);
xnor U4900 (N_4900,N_3469,N_3738);
and U4901 (N_4901,N_3205,N_3321);
and U4902 (N_4902,N_3547,N_3761);
and U4903 (N_4903,N_3107,N_3980);
nand U4904 (N_4904,N_3184,N_3447);
nor U4905 (N_4905,N_3222,N_3176);
and U4906 (N_4906,N_3085,N_3828);
and U4907 (N_4907,N_3977,N_3198);
xor U4908 (N_4908,N_3205,N_3600);
nand U4909 (N_4909,N_3051,N_3271);
and U4910 (N_4910,N_3096,N_3875);
and U4911 (N_4911,N_3436,N_3780);
nand U4912 (N_4912,N_3949,N_3939);
nor U4913 (N_4913,N_3066,N_3984);
or U4914 (N_4914,N_3232,N_3300);
nor U4915 (N_4915,N_3956,N_3725);
and U4916 (N_4916,N_3947,N_3272);
nor U4917 (N_4917,N_3388,N_3479);
nor U4918 (N_4918,N_3231,N_3669);
nor U4919 (N_4919,N_3384,N_3676);
nor U4920 (N_4920,N_3270,N_3918);
and U4921 (N_4921,N_3554,N_3332);
xnor U4922 (N_4922,N_3650,N_3862);
xnor U4923 (N_4923,N_3996,N_3131);
and U4924 (N_4924,N_3154,N_3505);
nand U4925 (N_4925,N_3866,N_3968);
or U4926 (N_4926,N_3310,N_3208);
nand U4927 (N_4927,N_3928,N_3629);
or U4928 (N_4928,N_3892,N_3854);
nand U4929 (N_4929,N_3761,N_3140);
or U4930 (N_4930,N_3666,N_3404);
xnor U4931 (N_4931,N_3753,N_3369);
nor U4932 (N_4932,N_3812,N_3318);
and U4933 (N_4933,N_3768,N_3861);
xnor U4934 (N_4934,N_3146,N_3726);
xnor U4935 (N_4935,N_3255,N_3866);
nor U4936 (N_4936,N_3470,N_3402);
and U4937 (N_4937,N_3690,N_3976);
or U4938 (N_4938,N_3916,N_3669);
xnor U4939 (N_4939,N_3123,N_3220);
and U4940 (N_4940,N_3463,N_3902);
nand U4941 (N_4941,N_3985,N_3485);
nand U4942 (N_4942,N_3467,N_3887);
or U4943 (N_4943,N_3703,N_3575);
nor U4944 (N_4944,N_3816,N_3292);
or U4945 (N_4945,N_3282,N_3202);
xnor U4946 (N_4946,N_3925,N_3897);
nand U4947 (N_4947,N_3487,N_3934);
or U4948 (N_4948,N_3722,N_3150);
nor U4949 (N_4949,N_3703,N_3538);
nand U4950 (N_4950,N_3532,N_3728);
and U4951 (N_4951,N_3525,N_3886);
and U4952 (N_4952,N_3478,N_3756);
or U4953 (N_4953,N_3442,N_3317);
and U4954 (N_4954,N_3409,N_3493);
xnor U4955 (N_4955,N_3054,N_3927);
xor U4956 (N_4956,N_3718,N_3702);
and U4957 (N_4957,N_3950,N_3917);
or U4958 (N_4958,N_3051,N_3301);
and U4959 (N_4959,N_3763,N_3415);
and U4960 (N_4960,N_3690,N_3129);
and U4961 (N_4961,N_3366,N_3888);
xnor U4962 (N_4962,N_3196,N_3869);
or U4963 (N_4963,N_3503,N_3365);
nand U4964 (N_4964,N_3620,N_3779);
nor U4965 (N_4965,N_3276,N_3160);
xnor U4966 (N_4966,N_3347,N_3866);
nor U4967 (N_4967,N_3819,N_3837);
nor U4968 (N_4968,N_3145,N_3174);
xor U4969 (N_4969,N_3398,N_3725);
nor U4970 (N_4970,N_3718,N_3383);
nor U4971 (N_4971,N_3241,N_3841);
xnor U4972 (N_4972,N_3907,N_3027);
or U4973 (N_4973,N_3175,N_3153);
nand U4974 (N_4974,N_3654,N_3457);
xnor U4975 (N_4975,N_3118,N_3326);
and U4976 (N_4976,N_3489,N_3496);
or U4977 (N_4977,N_3836,N_3971);
or U4978 (N_4978,N_3170,N_3404);
or U4979 (N_4979,N_3319,N_3648);
xnor U4980 (N_4980,N_3206,N_3359);
or U4981 (N_4981,N_3241,N_3025);
xor U4982 (N_4982,N_3084,N_3837);
nand U4983 (N_4983,N_3957,N_3092);
or U4984 (N_4984,N_3574,N_3459);
nand U4985 (N_4985,N_3457,N_3048);
or U4986 (N_4986,N_3259,N_3043);
nand U4987 (N_4987,N_3021,N_3194);
nor U4988 (N_4988,N_3679,N_3437);
xor U4989 (N_4989,N_3651,N_3985);
nor U4990 (N_4990,N_3685,N_3693);
nor U4991 (N_4991,N_3385,N_3436);
or U4992 (N_4992,N_3224,N_3805);
nand U4993 (N_4993,N_3176,N_3932);
xnor U4994 (N_4994,N_3699,N_3957);
nor U4995 (N_4995,N_3083,N_3751);
xnor U4996 (N_4996,N_3562,N_3137);
or U4997 (N_4997,N_3805,N_3669);
xor U4998 (N_4998,N_3999,N_3182);
nand U4999 (N_4999,N_3971,N_3274);
nor U5000 (N_5000,N_4407,N_4850);
and U5001 (N_5001,N_4355,N_4833);
nand U5002 (N_5002,N_4964,N_4174);
or U5003 (N_5003,N_4820,N_4685);
nor U5004 (N_5004,N_4233,N_4341);
or U5005 (N_5005,N_4491,N_4943);
and U5006 (N_5006,N_4713,N_4516);
nor U5007 (N_5007,N_4780,N_4023);
and U5008 (N_5008,N_4972,N_4599);
nand U5009 (N_5009,N_4231,N_4667);
nor U5010 (N_5010,N_4771,N_4671);
or U5011 (N_5011,N_4888,N_4154);
xnor U5012 (N_5012,N_4077,N_4448);
and U5013 (N_5013,N_4922,N_4322);
nand U5014 (N_5014,N_4526,N_4996);
and U5015 (N_5015,N_4345,N_4364);
xnor U5016 (N_5016,N_4110,N_4249);
nor U5017 (N_5017,N_4803,N_4814);
xor U5018 (N_5018,N_4193,N_4417);
nand U5019 (N_5019,N_4575,N_4657);
nand U5020 (N_5020,N_4026,N_4409);
or U5021 (N_5021,N_4948,N_4973);
or U5022 (N_5022,N_4038,N_4477);
or U5023 (N_5023,N_4502,N_4604);
nor U5024 (N_5024,N_4111,N_4933);
xor U5025 (N_5025,N_4600,N_4378);
xnor U5026 (N_5026,N_4829,N_4646);
nand U5027 (N_5027,N_4944,N_4445);
or U5028 (N_5028,N_4936,N_4775);
xor U5029 (N_5029,N_4184,N_4428);
or U5030 (N_5030,N_4628,N_4505);
nand U5031 (N_5031,N_4558,N_4458);
nor U5032 (N_5032,N_4256,N_4028);
nor U5033 (N_5033,N_4762,N_4162);
and U5034 (N_5034,N_4275,N_4043);
or U5035 (N_5035,N_4224,N_4408);
nor U5036 (N_5036,N_4506,N_4267);
nor U5037 (N_5037,N_4166,N_4260);
xor U5038 (N_5038,N_4248,N_4885);
and U5039 (N_5039,N_4072,N_4858);
nor U5040 (N_5040,N_4237,N_4896);
xnor U5041 (N_5041,N_4606,N_4765);
nor U5042 (N_5042,N_4180,N_4298);
and U5043 (N_5043,N_4379,N_4801);
nand U5044 (N_5044,N_4659,N_4925);
xnor U5045 (N_5045,N_4995,N_4441);
and U5046 (N_5046,N_4677,N_4168);
xnor U5047 (N_5047,N_4681,N_4638);
and U5048 (N_5048,N_4728,N_4084);
nand U5049 (N_5049,N_4213,N_4917);
or U5050 (N_5050,N_4869,N_4702);
nor U5051 (N_5051,N_4965,N_4429);
and U5052 (N_5052,N_4641,N_4980);
nor U5053 (N_5053,N_4487,N_4239);
xor U5054 (N_5054,N_4562,N_4016);
xor U5055 (N_5055,N_4394,N_4294);
xor U5056 (N_5056,N_4454,N_4482);
xnor U5057 (N_5057,N_4284,N_4512);
or U5058 (N_5058,N_4089,N_4092);
and U5059 (N_5059,N_4879,N_4645);
and U5060 (N_5060,N_4555,N_4088);
nor U5061 (N_5061,N_4361,N_4986);
nor U5062 (N_5062,N_4344,N_4565);
nor U5063 (N_5063,N_4283,N_4150);
nor U5064 (N_5064,N_4992,N_4613);
nand U5065 (N_5065,N_4483,N_4019);
nand U5066 (N_5066,N_4205,N_4642);
or U5067 (N_5067,N_4350,N_4511);
nor U5068 (N_5068,N_4410,N_4603);
nand U5069 (N_5069,N_4247,N_4336);
and U5070 (N_5070,N_4549,N_4706);
or U5071 (N_5071,N_4363,N_4773);
and U5072 (N_5072,N_4020,N_4737);
nand U5073 (N_5073,N_4911,N_4392);
and U5074 (N_5074,N_4694,N_4954);
nor U5075 (N_5075,N_4889,N_4472);
or U5076 (N_5076,N_4831,N_4086);
xor U5077 (N_5077,N_4501,N_4824);
or U5078 (N_5078,N_4013,N_4580);
or U5079 (N_5079,N_4669,N_4532);
xnor U5080 (N_5080,N_4893,N_4805);
nor U5081 (N_5081,N_4509,N_4198);
nand U5082 (N_5082,N_4176,N_4591);
nand U5083 (N_5083,N_4756,N_4238);
nor U5084 (N_5084,N_4131,N_4348);
xnor U5085 (N_5085,N_4195,N_4229);
xnor U5086 (N_5086,N_4203,N_4949);
nor U5087 (N_5087,N_4513,N_4931);
xnor U5088 (N_5088,N_4956,N_4220);
nor U5089 (N_5089,N_4607,N_4999);
nand U5090 (N_5090,N_4116,N_4542);
nor U5091 (N_5091,N_4676,N_4630);
xnor U5092 (N_5092,N_4495,N_4418);
and U5093 (N_5093,N_4800,N_4264);
nor U5094 (N_5094,N_4990,N_4847);
xor U5095 (N_5095,N_4356,N_4304);
nand U5096 (N_5096,N_4844,N_4941);
xnor U5097 (N_5097,N_4700,N_4480);
nor U5098 (N_5098,N_4717,N_4290);
nor U5099 (N_5099,N_4867,N_4354);
nand U5100 (N_5100,N_4317,N_4411);
and U5101 (N_5101,N_4437,N_4967);
xnor U5102 (N_5102,N_4621,N_4056);
or U5103 (N_5103,N_4537,N_4962);
or U5104 (N_5104,N_4935,N_4842);
and U5105 (N_5105,N_4251,N_4870);
or U5106 (N_5106,N_4006,N_4293);
or U5107 (N_5107,N_4004,N_4873);
nand U5108 (N_5108,N_4795,N_4959);
or U5109 (N_5109,N_4309,N_4209);
xor U5110 (N_5110,N_4250,N_4178);
or U5111 (N_5111,N_4312,N_4924);
nor U5112 (N_5112,N_4170,N_4474);
xnor U5113 (N_5113,N_4612,N_4519);
and U5114 (N_5114,N_4779,N_4450);
nand U5115 (N_5115,N_4637,N_4105);
and U5116 (N_5116,N_4804,N_4617);
or U5117 (N_5117,N_4633,N_4988);
nor U5118 (N_5118,N_4464,N_4977);
and U5119 (N_5119,N_4834,N_4191);
and U5120 (N_5120,N_4045,N_4697);
and U5121 (N_5121,N_4871,N_4711);
nand U5122 (N_5122,N_4707,N_4119);
nor U5123 (N_5123,N_4399,N_4052);
xor U5124 (N_5124,N_4504,N_4648);
xnor U5125 (N_5125,N_4571,N_4329);
and U5126 (N_5126,N_4757,N_4259);
or U5127 (N_5127,N_4930,N_4579);
xnor U5128 (N_5128,N_4272,N_4823);
nor U5129 (N_5129,N_4414,N_4357);
or U5130 (N_5130,N_4211,N_4859);
or U5131 (N_5131,N_4003,N_4576);
nor U5132 (N_5132,N_4839,N_4186);
nor U5133 (N_5133,N_4066,N_4650);
or U5134 (N_5134,N_4287,N_4416);
or U5135 (N_5135,N_4337,N_4811);
or U5136 (N_5136,N_4330,N_4978);
xor U5137 (N_5137,N_4367,N_4601);
and U5138 (N_5138,N_4902,N_4432);
and U5139 (N_5139,N_4451,N_4950);
and U5140 (N_5140,N_4254,N_4622);
nor U5141 (N_5141,N_4567,N_4548);
and U5142 (N_5142,N_4975,N_4686);
nand U5143 (N_5143,N_4557,N_4522);
or U5144 (N_5144,N_4087,N_4449);
nand U5145 (N_5145,N_4524,N_4760);
or U5146 (N_5146,N_4720,N_4569);
xnor U5147 (N_5147,N_4369,N_4325);
or U5148 (N_5148,N_4794,N_4172);
and U5149 (N_5149,N_4303,N_4815);
xor U5150 (N_5150,N_4071,N_4321);
or U5151 (N_5151,N_4583,N_4360);
and U5152 (N_5152,N_4271,N_4435);
and U5153 (N_5153,N_4000,N_4382);
nor U5154 (N_5154,N_4358,N_4792);
xnor U5155 (N_5155,N_4733,N_4405);
or U5156 (N_5156,N_4588,N_4422);
or U5157 (N_5157,N_4320,N_4161);
and U5158 (N_5158,N_4770,N_4208);
nor U5159 (N_5159,N_4169,N_4029);
or U5160 (N_5160,N_4094,N_4050);
xnor U5161 (N_5161,N_4521,N_4277);
xor U5162 (N_5162,N_4966,N_4598);
nand U5163 (N_5163,N_4587,N_4400);
or U5164 (N_5164,N_4031,N_4171);
nor U5165 (N_5165,N_4920,N_4214);
nor U5166 (N_5166,N_4955,N_4476);
nor U5167 (N_5167,N_4164,N_4957);
and U5168 (N_5168,N_4307,N_4739);
nor U5169 (N_5169,N_4563,N_4235);
nor U5170 (N_5170,N_4974,N_4701);
nor U5171 (N_5171,N_4696,N_4826);
and U5172 (N_5172,N_4396,N_4373);
or U5173 (N_5173,N_4776,N_4488);
nand U5174 (N_5174,N_4910,N_4046);
and U5175 (N_5175,N_4255,N_4160);
nor U5176 (N_5176,N_4037,N_4009);
nor U5177 (N_5177,N_4022,N_4489);
nor U5178 (N_5178,N_4610,N_4627);
and U5179 (N_5179,N_4377,N_4712);
and U5180 (N_5180,N_4553,N_4715);
or U5181 (N_5181,N_4242,N_4691);
xnor U5182 (N_5182,N_4528,N_4543);
xor U5183 (N_5183,N_4723,N_4117);
nor U5184 (N_5184,N_4291,N_4245);
nand U5185 (N_5185,N_4793,N_4012);
nand U5186 (N_5186,N_4300,N_4616);
and U5187 (N_5187,N_4976,N_4215);
or U5188 (N_5188,N_4987,N_4136);
nand U5189 (N_5189,N_4219,N_4586);
nand U5190 (N_5190,N_4151,N_4081);
and U5191 (N_5191,N_4158,N_4297);
nor U5192 (N_5192,N_4280,N_4629);
nor U5193 (N_5193,N_4093,N_4845);
xnor U5194 (N_5194,N_4130,N_4692);
nor U5195 (N_5195,N_4313,N_4206);
and U5196 (N_5196,N_4651,N_4693);
nand U5197 (N_5197,N_4611,N_4518);
and U5198 (N_5198,N_4118,N_4490);
or U5199 (N_5199,N_4375,N_4822);
or U5200 (N_5200,N_4385,N_4527);
or U5201 (N_5201,N_4817,N_4547);
nor U5202 (N_5202,N_4787,N_4806);
nor U5203 (N_5203,N_4989,N_4097);
and U5204 (N_5204,N_4568,N_4661);
and U5205 (N_5205,N_4452,N_4199);
nand U5206 (N_5206,N_4718,N_4327);
nand U5207 (N_5207,N_4531,N_4467);
xnor U5208 (N_5208,N_4636,N_4295);
nand U5209 (N_5209,N_4324,N_4062);
nand U5210 (N_5210,N_4574,N_4241);
nand U5211 (N_5211,N_4554,N_4556);
nor U5212 (N_5212,N_4708,N_4391);
xor U5213 (N_5213,N_4892,N_4940);
or U5214 (N_5214,N_4729,N_4486);
xor U5215 (N_5215,N_4849,N_4866);
nand U5216 (N_5216,N_4863,N_4658);
xnor U5217 (N_5217,N_4926,N_4049);
xor U5218 (N_5218,N_4132,N_4194);
and U5219 (N_5219,N_4748,N_4106);
nor U5220 (N_5220,N_4011,N_4500);
xnor U5221 (N_5221,N_4481,N_4017);
xnor U5222 (N_5222,N_4761,N_4589);
xnor U5223 (N_5223,N_4109,N_4240);
nand U5224 (N_5224,N_4210,N_4424);
or U5225 (N_5225,N_4069,N_4063);
xor U5226 (N_5226,N_4840,N_4101);
and U5227 (N_5227,N_4631,N_4076);
nor U5228 (N_5228,N_4352,N_4852);
or U5229 (N_5229,N_4122,N_4114);
or U5230 (N_5230,N_4015,N_4632);
nand U5231 (N_5231,N_4510,N_4226);
nand U5232 (N_5232,N_4758,N_4520);
nand U5233 (N_5233,N_4121,N_4721);
xor U5234 (N_5234,N_4138,N_4541);
xor U5235 (N_5235,N_4937,N_4851);
nand U5236 (N_5236,N_4305,N_4891);
xnor U5237 (N_5237,N_4137,N_4014);
and U5238 (N_5238,N_4459,N_4402);
or U5239 (N_5239,N_4857,N_4942);
nand U5240 (N_5240,N_4872,N_4266);
or U5241 (N_5241,N_4230,N_4544);
xor U5242 (N_5242,N_4647,N_4460);
and U5243 (N_5243,N_4884,N_4623);
xor U5244 (N_5244,N_4783,N_4722);
nor U5245 (N_5245,N_4906,N_4912);
nand U5246 (N_5246,N_4279,N_4900);
or U5247 (N_5247,N_4427,N_4877);
and U5248 (N_5248,N_4156,N_4079);
nand U5249 (N_5249,N_4991,N_4660);
or U5250 (N_5250,N_4192,N_4024);
and U5251 (N_5251,N_4025,N_4484);
and U5252 (N_5252,N_4133,N_4807);
xnor U5253 (N_5253,N_4075,N_4351);
xnor U5254 (N_5254,N_4887,N_4703);
nand U5255 (N_5255,N_4881,N_4061);
and U5256 (N_5256,N_4243,N_4534);
or U5257 (N_5257,N_4430,N_4129);
nor U5258 (N_5258,N_4462,N_4535);
nand U5259 (N_5259,N_4919,N_4306);
or U5260 (N_5260,N_4340,N_4068);
or U5261 (N_5261,N_4578,N_4503);
and U5262 (N_5262,N_4932,N_4672);
or U5263 (N_5263,N_4998,N_4832);
or U5264 (N_5264,N_4767,N_4420);
and U5265 (N_5265,N_4876,N_4690);
and U5266 (N_5266,N_4618,N_4564);
nand U5267 (N_5267,N_4102,N_4818);
nand U5268 (N_5268,N_4673,N_4898);
nand U5269 (N_5269,N_4197,N_4257);
nand U5270 (N_5270,N_4639,N_4281);
and U5271 (N_5271,N_4552,N_4107);
and U5272 (N_5272,N_4401,N_4838);
nor U5273 (N_5273,N_4566,N_4590);
xnor U5274 (N_5274,N_4853,N_4752);
nor U5275 (N_5275,N_4057,N_4719);
or U5276 (N_5276,N_4615,N_4790);
nand U5277 (N_5277,N_4308,N_4497);
and U5278 (N_5278,N_4440,N_4395);
or U5279 (N_5279,N_4808,N_4246);
or U5280 (N_5280,N_4145,N_4799);
or U5281 (N_5281,N_4635,N_4453);
xnor U5282 (N_5282,N_4047,N_4584);
nand U5283 (N_5283,N_4750,N_4159);
and U5284 (N_5284,N_4143,N_4342);
nor U5285 (N_5285,N_4594,N_4423);
or U5286 (N_5286,N_4861,N_4812);
nor U5287 (N_5287,N_4680,N_4044);
nor U5288 (N_5288,N_4332,N_4821);
or U5289 (N_5289,N_4302,N_4163);
nand U5290 (N_5290,N_4916,N_4918);
or U5291 (N_5291,N_4412,N_4338);
xnor U5292 (N_5292,N_4095,N_4494);
nand U5293 (N_5293,N_4433,N_4883);
nand U5294 (N_5294,N_4749,N_4862);
and U5295 (N_5295,N_4945,N_4963);
or U5296 (N_5296,N_4727,N_4323);
and U5297 (N_5297,N_4655,N_4335);
nand U5298 (N_5298,N_4791,N_4514);
and U5299 (N_5299,N_4289,N_4099);
and U5300 (N_5300,N_4296,N_4856);
nand U5301 (N_5301,N_4263,N_4705);
xor U5302 (N_5302,N_4415,N_4921);
and U5303 (N_5303,N_4010,N_4292);
or U5304 (N_5304,N_4426,N_4843);
or U5305 (N_5305,N_4915,N_4529);
nor U5306 (N_5306,N_4777,N_4837);
or U5307 (N_5307,N_4666,N_4759);
xnor U5308 (N_5308,N_4536,N_4540);
and U5309 (N_5309,N_4983,N_4070);
nor U5310 (N_5310,N_4841,N_4596);
and U5311 (N_5311,N_4736,N_4042);
and U5312 (N_5312,N_4585,N_4624);
and U5313 (N_5313,N_4146,N_4388);
xor U5314 (N_5314,N_4581,N_4640);
and U5315 (N_5315,N_4390,N_4626);
nand U5316 (N_5316,N_4466,N_4286);
xnor U5317 (N_5317,N_4985,N_4326);
xnor U5318 (N_5318,N_4124,N_4784);
and U5319 (N_5319,N_4007,N_4316);
xor U5320 (N_5320,N_4142,N_4609);
nor U5321 (N_5321,N_4187,N_4679);
and U5322 (N_5322,N_4463,N_4570);
and U5323 (N_5323,N_4155,N_4059);
xor U5324 (N_5324,N_4764,N_4083);
xnor U5325 (N_5325,N_4112,N_4864);
nand U5326 (N_5326,N_4465,N_4836);
xnor U5327 (N_5327,N_4461,N_4381);
and U5328 (N_5328,N_4383,N_4714);
nor U5329 (N_5329,N_4969,N_4314);
xnor U5330 (N_5330,N_4034,N_4455);
and U5331 (N_5331,N_4258,N_4875);
xnor U5332 (N_5332,N_4301,N_4496);
and U5333 (N_5333,N_4809,N_4668);
nor U5334 (N_5334,N_4802,N_4997);
nor U5335 (N_5335,N_4123,N_4830);
xor U5336 (N_5336,N_4148,N_4927);
nand U5337 (N_5337,N_4582,N_4970);
xor U5338 (N_5338,N_4040,N_4055);
nand U5339 (N_5339,N_4436,N_4781);
nand U5340 (N_5340,N_4903,N_4868);
and U5341 (N_5341,N_4273,N_4048);
nand U5342 (N_5342,N_4678,N_4227);
xor U5343 (N_5343,N_4855,N_4656);
nand U5344 (N_5344,N_4152,N_4421);
xor U5345 (N_5345,N_4065,N_4183);
and U5346 (N_5346,N_4662,N_4030);
and U5347 (N_5347,N_4653,N_4090);
or U5348 (N_5348,N_4649,N_4595);
and U5349 (N_5349,N_4319,N_4001);
nand U5350 (N_5350,N_4766,N_4725);
or U5351 (N_5351,N_4054,N_4744);
and U5352 (N_5352,N_4082,N_4498);
nor U5353 (N_5353,N_4147,N_4053);
xor U5354 (N_5354,N_4201,N_4769);
or U5355 (N_5355,N_4431,N_4270);
nor U5356 (N_5356,N_4605,N_4370);
and U5357 (N_5357,N_4797,N_4128);
and U5358 (N_5358,N_4468,N_4202);
nor U5359 (N_5359,N_4865,N_4096);
nand U5360 (N_5360,N_4139,N_4127);
nor U5361 (N_5361,N_4036,N_4934);
nand U5362 (N_5362,N_4153,N_4874);
nand U5363 (N_5363,N_4157,N_4078);
nor U5364 (N_5364,N_4113,N_4288);
or U5365 (N_5365,N_4175,N_4825);
xnor U5366 (N_5366,N_4993,N_4643);
nor U5367 (N_5367,N_4904,N_4545);
xor U5368 (N_5368,N_4098,N_4982);
nor U5369 (N_5369,N_4994,N_4473);
nand U5370 (N_5370,N_4860,N_4366);
nor U5371 (N_5371,N_4878,N_4108);
xor U5372 (N_5372,N_4755,N_4644);
and U5373 (N_5373,N_4359,N_4960);
xor U5374 (N_5374,N_4939,N_4269);
and U5375 (N_5375,N_4508,N_4315);
and U5376 (N_5376,N_4827,N_4968);
or U5377 (N_5377,N_4561,N_4740);
nor U5378 (N_5378,N_4126,N_4334);
nand U5379 (N_5379,N_4614,N_4285);
and U5380 (N_5380,N_4785,N_4216);
or U5381 (N_5381,N_4716,N_4625);
or U5382 (N_5382,N_4493,N_4393);
nand U5383 (N_5383,N_4786,N_4371);
or U5384 (N_5384,N_4523,N_4167);
xnor U5385 (N_5385,N_4021,N_4173);
and U5386 (N_5386,N_4539,N_4782);
or U5387 (N_5387,N_4741,N_4559);
nor U5388 (N_5388,N_4346,N_4525);
nand U5389 (N_5389,N_4058,N_4731);
nand U5390 (N_5390,N_4828,N_4041);
nand U5391 (N_5391,N_4689,N_4406);
nor U5392 (N_5392,N_4438,N_4443);
and U5393 (N_5393,N_4261,N_4981);
nor U5394 (N_5394,N_4018,N_4204);
nor U5395 (N_5395,N_4745,N_4492);
or U5396 (N_5396,N_4515,N_4442);
nand U5397 (N_5397,N_4895,N_4665);
nand U5398 (N_5398,N_4909,N_4709);
and U5399 (N_5399,N_4517,N_4899);
xnor U5400 (N_5400,N_4747,N_4347);
nor U5401 (N_5401,N_4165,N_4276);
and U5402 (N_5402,N_4738,N_4135);
nor U5403 (N_5403,N_4002,N_4035);
and U5404 (N_5404,N_4188,N_4971);
or U5405 (N_5405,N_4343,N_4221);
and U5406 (N_5406,N_4282,N_4262);
nand U5407 (N_5407,N_4479,N_4951);
xor U5408 (N_5408,N_4311,N_4593);
and U5409 (N_5409,N_4947,N_4386);
xnor U5410 (N_5410,N_4880,N_4810);
nand U5411 (N_5411,N_4234,N_4404);
xnor U5412 (N_5412,N_4958,N_4365);
nor U5413 (N_5413,N_4546,N_4100);
nand U5414 (N_5414,N_4478,N_4372);
and U5415 (N_5415,N_4684,N_4200);
nand U5416 (N_5416,N_4675,N_4217);
nor U5417 (N_5417,N_4073,N_4961);
nor U5418 (N_5418,N_4890,N_4602);
xnor U5419 (N_5419,N_4835,N_4318);
or U5420 (N_5420,N_4274,N_4952);
nor U5421 (N_5421,N_4218,N_4039);
or U5422 (N_5422,N_4104,N_4953);
nand U5423 (N_5423,N_4688,N_4457);
or U5424 (N_5424,N_4236,N_4067);
nor U5425 (N_5425,N_4742,N_4470);
or U5426 (N_5426,N_4695,N_4140);
and U5427 (N_5427,N_4085,N_4670);
nor U5428 (N_5428,N_4819,N_4349);
or U5429 (N_5429,N_4222,N_4190);
nand U5430 (N_5430,N_4507,N_4439);
nor U5431 (N_5431,N_4333,N_4734);
nand U5432 (N_5432,N_4735,N_4005);
nand U5433 (N_5433,N_4223,N_4032);
or U5434 (N_5434,N_4149,N_4634);
xor U5435 (N_5435,N_4789,N_4091);
xor U5436 (N_5436,N_4120,N_4597);
and U5437 (N_5437,N_4710,N_4928);
xnor U5438 (N_5438,N_4654,N_4380);
or U5439 (N_5439,N_4403,N_4577);
or U5440 (N_5440,N_4746,N_4984);
xnor U5441 (N_5441,N_4704,N_4469);
nor U5442 (N_5442,N_4724,N_4652);
xnor U5443 (N_5443,N_4115,N_4027);
xnor U5444 (N_5444,N_4664,N_4929);
xor U5445 (N_5445,N_4572,N_4244);
and U5446 (N_5446,N_4620,N_4674);
or U5447 (N_5447,N_4447,N_4182);
xor U5448 (N_5448,N_4798,N_4232);
xor U5449 (N_5449,N_4753,N_4573);
nand U5450 (N_5450,N_4592,N_4726);
xnor U5451 (N_5451,N_4397,N_4339);
nor U5452 (N_5452,N_4751,N_4763);
xor U5453 (N_5453,N_4699,N_4471);
nor U5454 (N_5454,N_4475,N_4499);
or U5455 (N_5455,N_4908,N_4389);
and U5456 (N_5456,N_4196,N_4485);
xnor U5457 (N_5457,N_4754,N_4225);
and U5458 (N_5458,N_4368,N_4177);
or U5459 (N_5459,N_4252,N_4854);
nor U5460 (N_5460,N_4446,N_4778);
nand U5461 (N_5461,N_4398,N_4730);
nor U5462 (N_5462,N_4914,N_4268);
or U5463 (N_5463,N_4846,N_4560);
or U5464 (N_5464,N_4064,N_4444);
or U5465 (N_5465,N_4212,N_4331);
xnor U5466 (N_5466,N_4608,N_4253);
or U5467 (N_5467,N_4207,N_4743);
or U5468 (N_5468,N_4387,N_4683);
nor U5469 (N_5469,N_4144,N_4816);
nand U5470 (N_5470,N_4923,N_4901);
nand U5471 (N_5471,N_4310,N_4299);
or U5472 (N_5472,N_4768,N_4374);
nor U5473 (N_5473,N_4376,N_4103);
or U5474 (N_5474,N_4813,N_4080);
nor U5475 (N_5475,N_4179,N_4788);
nand U5476 (N_5476,N_4848,N_4796);
or U5477 (N_5477,N_4384,N_4774);
and U5478 (N_5478,N_4897,N_4619);
nor U5479 (N_5479,N_4362,N_4663);
nor U5480 (N_5480,N_4060,N_4134);
nand U5481 (N_5481,N_4979,N_4228);
or U5482 (N_5482,N_4682,N_4687);
nor U5483 (N_5483,N_4533,N_4141);
and U5484 (N_5484,N_4425,N_4353);
or U5485 (N_5485,N_4907,N_4278);
and U5486 (N_5486,N_4181,N_4698);
nor U5487 (N_5487,N_4074,N_4938);
and U5488 (N_5488,N_4033,N_4413);
and U5489 (N_5489,N_4550,N_4008);
nand U5490 (N_5490,N_4772,N_4419);
or U5491 (N_5491,N_4882,N_4946);
or U5492 (N_5492,N_4189,N_4328);
or U5493 (N_5493,N_4551,N_4051);
or U5494 (N_5494,N_4265,N_4913);
nand U5495 (N_5495,N_4125,N_4530);
xor U5496 (N_5496,N_4886,N_4185);
or U5497 (N_5497,N_4894,N_4434);
and U5498 (N_5498,N_4732,N_4456);
or U5499 (N_5499,N_4905,N_4538);
or U5500 (N_5500,N_4009,N_4610);
and U5501 (N_5501,N_4606,N_4237);
nand U5502 (N_5502,N_4619,N_4472);
nand U5503 (N_5503,N_4952,N_4418);
nand U5504 (N_5504,N_4782,N_4686);
nor U5505 (N_5505,N_4331,N_4831);
or U5506 (N_5506,N_4337,N_4001);
xnor U5507 (N_5507,N_4737,N_4128);
xor U5508 (N_5508,N_4188,N_4378);
or U5509 (N_5509,N_4734,N_4482);
nand U5510 (N_5510,N_4540,N_4443);
and U5511 (N_5511,N_4759,N_4936);
or U5512 (N_5512,N_4935,N_4162);
and U5513 (N_5513,N_4389,N_4139);
or U5514 (N_5514,N_4783,N_4978);
nor U5515 (N_5515,N_4363,N_4037);
or U5516 (N_5516,N_4830,N_4794);
and U5517 (N_5517,N_4167,N_4571);
xnor U5518 (N_5518,N_4773,N_4765);
nor U5519 (N_5519,N_4840,N_4302);
or U5520 (N_5520,N_4229,N_4790);
nand U5521 (N_5521,N_4454,N_4818);
nand U5522 (N_5522,N_4217,N_4633);
nand U5523 (N_5523,N_4611,N_4777);
or U5524 (N_5524,N_4214,N_4573);
nor U5525 (N_5525,N_4123,N_4178);
and U5526 (N_5526,N_4316,N_4563);
nor U5527 (N_5527,N_4668,N_4564);
and U5528 (N_5528,N_4967,N_4439);
and U5529 (N_5529,N_4036,N_4731);
nor U5530 (N_5530,N_4270,N_4039);
nand U5531 (N_5531,N_4179,N_4755);
nand U5532 (N_5532,N_4743,N_4213);
and U5533 (N_5533,N_4181,N_4710);
or U5534 (N_5534,N_4724,N_4920);
nand U5535 (N_5535,N_4024,N_4616);
xnor U5536 (N_5536,N_4798,N_4448);
and U5537 (N_5537,N_4126,N_4078);
nor U5538 (N_5538,N_4916,N_4831);
or U5539 (N_5539,N_4653,N_4093);
nand U5540 (N_5540,N_4098,N_4364);
nand U5541 (N_5541,N_4080,N_4406);
nor U5542 (N_5542,N_4186,N_4331);
nand U5543 (N_5543,N_4022,N_4534);
xnor U5544 (N_5544,N_4146,N_4253);
xor U5545 (N_5545,N_4850,N_4443);
nor U5546 (N_5546,N_4007,N_4061);
nand U5547 (N_5547,N_4050,N_4197);
nand U5548 (N_5548,N_4382,N_4311);
xor U5549 (N_5549,N_4726,N_4594);
nor U5550 (N_5550,N_4052,N_4849);
or U5551 (N_5551,N_4050,N_4112);
and U5552 (N_5552,N_4105,N_4601);
or U5553 (N_5553,N_4104,N_4211);
nand U5554 (N_5554,N_4383,N_4660);
nor U5555 (N_5555,N_4933,N_4652);
xor U5556 (N_5556,N_4173,N_4595);
and U5557 (N_5557,N_4524,N_4868);
or U5558 (N_5558,N_4522,N_4327);
xor U5559 (N_5559,N_4746,N_4303);
xnor U5560 (N_5560,N_4283,N_4380);
or U5561 (N_5561,N_4675,N_4743);
nor U5562 (N_5562,N_4702,N_4865);
nor U5563 (N_5563,N_4820,N_4565);
nand U5564 (N_5564,N_4428,N_4591);
nand U5565 (N_5565,N_4099,N_4827);
nor U5566 (N_5566,N_4655,N_4507);
or U5567 (N_5567,N_4665,N_4364);
and U5568 (N_5568,N_4315,N_4377);
xor U5569 (N_5569,N_4180,N_4592);
nand U5570 (N_5570,N_4834,N_4910);
xor U5571 (N_5571,N_4026,N_4627);
xor U5572 (N_5572,N_4917,N_4371);
nand U5573 (N_5573,N_4466,N_4549);
xor U5574 (N_5574,N_4807,N_4526);
and U5575 (N_5575,N_4238,N_4502);
or U5576 (N_5576,N_4452,N_4082);
or U5577 (N_5577,N_4498,N_4093);
or U5578 (N_5578,N_4850,N_4326);
nand U5579 (N_5579,N_4892,N_4352);
xnor U5580 (N_5580,N_4354,N_4532);
xor U5581 (N_5581,N_4829,N_4163);
and U5582 (N_5582,N_4679,N_4376);
and U5583 (N_5583,N_4728,N_4973);
or U5584 (N_5584,N_4544,N_4962);
nor U5585 (N_5585,N_4804,N_4181);
nand U5586 (N_5586,N_4564,N_4240);
or U5587 (N_5587,N_4054,N_4195);
or U5588 (N_5588,N_4589,N_4303);
and U5589 (N_5589,N_4714,N_4220);
xnor U5590 (N_5590,N_4320,N_4483);
nand U5591 (N_5591,N_4620,N_4320);
and U5592 (N_5592,N_4483,N_4718);
or U5593 (N_5593,N_4678,N_4687);
nand U5594 (N_5594,N_4462,N_4946);
nand U5595 (N_5595,N_4363,N_4067);
and U5596 (N_5596,N_4036,N_4380);
xor U5597 (N_5597,N_4222,N_4829);
and U5598 (N_5598,N_4833,N_4189);
nor U5599 (N_5599,N_4900,N_4784);
xnor U5600 (N_5600,N_4471,N_4682);
or U5601 (N_5601,N_4945,N_4410);
nand U5602 (N_5602,N_4598,N_4602);
nor U5603 (N_5603,N_4122,N_4893);
or U5604 (N_5604,N_4412,N_4433);
and U5605 (N_5605,N_4070,N_4663);
and U5606 (N_5606,N_4818,N_4623);
nor U5607 (N_5607,N_4091,N_4453);
or U5608 (N_5608,N_4437,N_4426);
nand U5609 (N_5609,N_4168,N_4447);
xnor U5610 (N_5610,N_4355,N_4088);
xor U5611 (N_5611,N_4917,N_4897);
or U5612 (N_5612,N_4996,N_4956);
nor U5613 (N_5613,N_4129,N_4102);
xnor U5614 (N_5614,N_4665,N_4102);
xor U5615 (N_5615,N_4833,N_4637);
or U5616 (N_5616,N_4276,N_4456);
nor U5617 (N_5617,N_4303,N_4468);
xor U5618 (N_5618,N_4947,N_4192);
and U5619 (N_5619,N_4081,N_4185);
and U5620 (N_5620,N_4086,N_4334);
nor U5621 (N_5621,N_4185,N_4102);
or U5622 (N_5622,N_4595,N_4910);
nand U5623 (N_5623,N_4598,N_4706);
nor U5624 (N_5624,N_4159,N_4027);
and U5625 (N_5625,N_4344,N_4102);
and U5626 (N_5626,N_4986,N_4770);
xor U5627 (N_5627,N_4406,N_4784);
xnor U5628 (N_5628,N_4244,N_4643);
xor U5629 (N_5629,N_4758,N_4793);
nand U5630 (N_5630,N_4740,N_4688);
or U5631 (N_5631,N_4837,N_4087);
nand U5632 (N_5632,N_4405,N_4457);
or U5633 (N_5633,N_4397,N_4935);
xnor U5634 (N_5634,N_4709,N_4659);
nor U5635 (N_5635,N_4859,N_4929);
or U5636 (N_5636,N_4217,N_4291);
nor U5637 (N_5637,N_4819,N_4479);
nor U5638 (N_5638,N_4611,N_4003);
nor U5639 (N_5639,N_4861,N_4964);
and U5640 (N_5640,N_4566,N_4816);
nor U5641 (N_5641,N_4267,N_4555);
nor U5642 (N_5642,N_4749,N_4152);
or U5643 (N_5643,N_4754,N_4668);
nor U5644 (N_5644,N_4197,N_4996);
or U5645 (N_5645,N_4203,N_4071);
nand U5646 (N_5646,N_4326,N_4530);
or U5647 (N_5647,N_4671,N_4982);
or U5648 (N_5648,N_4868,N_4323);
xnor U5649 (N_5649,N_4912,N_4682);
nand U5650 (N_5650,N_4325,N_4119);
and U5651 (N_5651,N_4199,N_4581);
nor U5652 (N_5652,N_4279,N_4664);
nand U5653 (N_5653,N_4703,N_4064);
nand U5654 (N_5654,N_4302,N_4389);
and U5655 (N_5655,N_4099,N_4901);
nor U5656 (N_5656,N_4714,N_4953);
or U5657 (N_5657,N_4306,N_4039);
nand U5658 (N_5658,N_4174,N_4187);
and U5659 (N_5659,N_4589,N_4032);
or U5660 (N_5660,N_4451,N_4551);
or U5661 (N_5661,N_4725,N_4967);
or U5662 (N_5662,N_4653,N_4319);
or U5663 (N_5663,N_4944,N_4669);
xnor U5664 (N_5664,N_4770,N_4684);
nor U5665 (N_5665,N_4697,N_4039);
or U5666 (N_5666,N_4931,N_4262);
nand U5667 (N_5667,N_4941,N_4975);
nor U5668 (N_5668,N_4125,N_4604);
nand U5669 (N_5669,N_4191,N_4889);
nor U5670 (N_5670,N_4411,N_4204);
nor U5671 (N_5671,N_4500,N_4648);
nand U5672 (N_5672,N_4879,N_4359);
xnor U5673 (N_5673,N_4171,N_4948);
and U5674 (N_5674,N_4084,N_4372);
and U5675 (N_5675,N_4241,N_4749);
xnor U5676 (N_5676,N_4163,N_4967);
nand U5677 (N_5677,N_4876,N_4571);
nor U5678 (N_5678,N_4466,N_4231);
and U5679 (N_5679,N_4485,N_4483);
nand U5680 (N_5680,N_4975,N_4293);
nand U5681 (N_5681,N_4791,N_4327);
or U5682 (N_5682,N_4560,N_4404);
nand U5683 (N_5683,N_4292,N_4766);
and U5684 (N_5684,N_4921,N_4416);
and U5685 (N_5685,N_4067,N_4621);
nand U5686 (N_5686,N_4651,N_4413);
nand U5687 (N_5687,N_4586,N_4319);
and U5688 (N_5688,N_4244,N_4506);
and U5689 (N_5689,N_4056,N_4315);
nand U5690 (N_5690,N_4143,N_4605);
or U5691 (N_5691,N_4527,N_4416);
or U5692 (N_5692,N_4126,N_4068);
nor U5693 (N_5693,N_4985,N_4852);
nor U5694 (N_5694,N_4178,N_4025);
and U5695 (N_5695,N_4612,N_4443);
or U5696 (N_5696,N_4106,N_4237);
or U5697 (N_5697,N_4205,N_4082);
xnor U5698 (N_5698,N_4190,N_4092);
nand U5699 (N_5699,N_4458,N_4621);
or U5700 (N_5700,N_4146,N_4731);
nor U5701 (N_5701,N_4351,N_4584);
or U5702 (N_5702,N_4821,N_4274);
and U5703 (N_5703,N_4870,N_4526);
nand U5704 (N_5704,N_4238,N_4779);
xor U5705 (N_5705,N_4636,N_4184);
xnor U5706 (N_5706,N_4810,N_4243);
or U5707 (N_5707,N_4559,N_4882);
and U5708 (N_5708,N_4260,N_4811);
xnor U5709 (N_5709,N_4030,N_4568);
xnor U5710 (N_5710,N_4883,N_4552);
or U5711 (N_5711,N_4832,N_4605);
nor U5712 (N_5712,N_4316,N_4583);
or U5713 (N_5713,N_4885,N_4453);
or U5714 (N_5714,N_4693,N_4550);
and U5715 (N_5715,N_4316,N_4815);
xor U5716 (N_5716,N_4340,N_4532);
and U5717 (N_5717,N_4562,N_4583);
nand U5718 (N_5718,N_4504,N_4242);
and U5719 (N_5719,N_4323,N_4922);
nor U5720 (N_5720,N_4287,N_4638);
nand U5721 (N_5721,N_4591,N_4317);
and U5722 (N_5722,N_4254,N_4958);
nor U5723 (N_5723,N_4332,N_4544);
or U5724 (N_5724,N_4164,N_4554);
and U5725 (N_5725,N_4569,N_4992);
and U5726 (N_5726,N_4112,N_4625);
xor U5727 (N_5727,N_4997,N_4781);
and U5728 (N_5728,N_4192,N_4095);
nor U5729 (N_5729,N_4320,N_4253);
xor U5730 (N_5730,N_4686,N_4044);
and U5731 (N_5731,N_4446,N_4271);
xnor U5732 (N_5732,N_4288,N_4149);
xnor U5733 (N_5733,N_4570,N_4220);
xor U5734 (N_5734,N_4560,N_4444);
nand U5735 (N_5735,N_4956,N_4307);
or U5736 (N_5736,N_4283,N_4924);
or U5737 (N_5737,N_4702,N_4779);
nor U5738 (N_5738,N_4745,N_4420);
xnor U5739 (N_5739,N_4870,N_4130);
and U5740 (N_5740,N_4322,N_4800);
nor U5741 (N_5741,N_4215,N_4286);
nor U5742 (N_5742,N_4333,N_4292);
or U5743 (N_5743,N_4203,N_4287);
and U5744 (N_5744,N_4978,N_4104);
xor U5745 (N_5745,N_4491,N_4605);
or U5746 (N_5746,N_4882,N_4425);
nand U5747 (N_5747,N_4064,N_4394);
nor U5748 (N_5748,N_4862,N_4229);
or U5749 (N_5749,N_4666,N_4050);
xnor U5750 (N_5750,N_4869,N_4197);
xor U5751 (N_5751,N_4320,N_4604);
or U5752 (N_5752,N_4763,N_4951);
nor U5753 (N_5753,N_4286,N_4064);
nor U5754 (N_5754,N_4757,N_4925);
nand U5755 (N_5755,N_4218,N_4199);
xor U5756 (N_5756,N_4694,N_4638);
xor U5757 (N_5757,N_4475,N_4611);
nor U5758 (N_5758,N_4387,N_4746);
or U5759 (N_5759,N_4663,N_4607);
xor U5760 (N_5760,N_4489,N_4759);
nor U5761 (N_5761,N_4656,N_4661);
and U5762 (N_5762,N_4412,N_4244);
nor U5763 (N_5763,N_4934,N_4912);
and U5764 (N_5764,N_4198,N_4346);
or U5765 (N_5765,N_4868,N_4779);
xor U5766 (N_5766,N_4298,N_4218);
and U5767 (N_5767,N_4643,N_4460);
and U5768 (N_5768,N_4130,N_4425);
and U5769 (N_5769,N_4634,N_4185);
or U5770 (N_5770,N_4540,N_4405);
nor U5771 (N_5771,N_4899,N_4698);
or U5772 (N_5772,N_4338,N_4848);
and U5773 (N_5773,N_4596,N_4606);
and U5774 (N_5774,N_4406,N_4071);
xnor U5775 (N_5775,N_4919,N_4196);
or U5776 (N_5776,N_4171,N_4153);
nor U5777 (N_5777,N_4237,N_4475);
nor U5778 (N_5778,N_4133,N_4954);
xnor U5779 (N_5779,N_4294,N_4970);
nand U5780 (N_5780,N_4970,N_4538);
or U5781 (N_5781,N_4496,N_4910);
nand U5782 (N_5782,N_4502,N_4328);
xor U5783 (N_5783,N_4459,N_4645);
or U5784 (N_5784,N_4876,N_4023);
or U5785 (N_5785,N_4434,N_4844);
nand U5786 (N_5786,N_4017,N_4611);
nand U5787 (N_5787,N_4761,N_4813);
xor U5788 (N_5788,N_4935,N_4138);
nor U5789 (N_5789,N_4051,N_4086);
xor U5790 (N_5790,N_4523,N_4274);
and U5791 (N_5791,N_4511,N_4185);
and U5792 (N_5792,N_4843,N_4044);
nor U5793 (N_5793,N_4420,N_4652);
nor U5794 (N_5794,N_4294,N_4160);
nand U5795 (N_5795,N_4220,N_4781);
or U5796 (N_5796,N_4488,N_4703);
nor U5797 (N_5797,N_4703,N_4753);
xor U5798 (N_5798,N_4959,N_4273);
or U5799 (N_5799,N_4304,N_4909);
or U5800 (N_5800,N_4991,N_4671);
or U5801 (N_5801,N_4999,N_4508);
nor U5802 (N_5802,N_4985,N_4736);
nand U5803 (N_5803,N_4044,N_4618);
xnor U5804 (N_5804,N_4894,N_4771);
and U5805 (N_5805,N_4952,N_4510);
nand U5806 (N_5806,N_4010,N_4861);
nor U5807 (N_5807,N_4390,N_4796);
or U5808 (N_5808,N_4625,N_4440);
xor U5809 (N_5809,N_4653,N_4734);
and U5810 (N_5810,N_4832,N_4425);
nand U5811 (N_5811,N_4337,N_4618);
xnor U5812 (N_5812,N_4218,N_4338);
xor U5813 (N_5813,N_4998,N_4601);
nand U5814 (N_5814,N_4351,N_4954);
nand U5815 (N_5815,N_4088,N_4126);
nand U5816 (N_5816,N_4187,N_4074);
nand U5817 (N_5817,N_4972,N_4860);
xor U5818 (N_5818,N_4632,N_4908);
nand U5819 (N_5819,N_4211,N_4187);
xor U5820 (N_5820,N_4030,N_4145);
nand U5821 (N_5821,N_4909,N_4168);
or U5822 (N_5822,N_4870,N_4651);
or U5823 (N_5823,N_4958,N_4049);
xor U5824 (N_5824,N_4326,N_4261);
or U5825 (N_5825,N_4449,N_4422);
nor U5826 (N_5826,N_4987,N_4296);
or U5827 (N_5827,N_4691,N_4295);
and U5828 (N_5828,N_4200,N_4440);
and U5829 (N_5829,N_4553,N_4941);
or U5830 (N_5830,N_4604,N_4744);
xor U5831 (N_5831,N_4980,N_4547);
xnor U5832 (N_5832,N_4352,N_4025);
or U5833 (N_5833,N_4697,N_4803);
nand U5834 (N_5834,N_4148,N_4854);
nand U5835 (N_5835,N_4256,N_4554);
and U5836 (N_5836,N_4114,N_4790);
xnor U5837 (N_5837,N_4586,N_4201);
nor U5838 (N_5838,N_4753,N_4093);
or U5839 (N_5839,N_4900,N_4478);
nand U5840 (N_5840,N_4325,N_4013);
nor U5841 (N_5841,N_4130,N_4477);
xnor U5842 (N_5842,N_4073,N_4786);
or U5843 (N_5843,N_4384,N_4125);
and U5844 (N_5844,N_4863,N_4033);
nand U5845 (N_5845,N_4872,N_4763);
xor U5846 (N_5846,N_4717,N_4534);
nand U5847 (N_5847,N_4169,N_4487);
nor U5848 (N_5848,N_4194,N_4788);
nor U5849 (N_5849,N_4517,N_4871);
or U5850 (N_5850,N_4111,N_4982);
nand U5851 (N_5851,N_4378,N_4667);
and U5852 (N_5852,N_4096,N_4848);
nand U5853 (N_5853,N_4923,N_4214);
and U5854 (N_5854,N_4549,N_4363);
nand U5855 (N_5855,N_4629,N_4257);
or U5856 (N_5856,N_4199,N_4941);
nor U5857 (N_5857,N_4006,N_4725);
nor U5858 (N_5858,N_4751,N_4902);
or U5859 (N_5859,N_4713,N_4155);
nand U5860 (N_5860,N_4840,N_4371);
nor U5861 (N_5861,N_4192,N_4128);
nand U5862 (N_5862,N_4331,N_4267);
or U5863 (N_5863,N_4637,N_4307);
or U5864 (N_5864,N_4686,N_4002);
nand U5865 (N_5865,N_4587,N_4439);
and U5866 (N_5866,N_4764,N_4916);
and U5867 (N_5867,N_4226,N_4289);
or U5868 (N_5868,N_4167,N_4391);
nor U5869 (N_5869,N_4025,N_4549);
nor U5870 (N_5870,N_4297,N_4083);
or U5871 (N_5871,N_4779,N_4947);
nor U5872 (N_5872,N_4675,N_4133);
xor U5873 (N_5873,N_4294,N_4180);
xor U5874 (N_5874,N_4887,N_4302);
xnor U5875 (N_5875,N_4484,N_4505);
nor U5876 (N_5876,N_4201,N_4810);
nand U5877 (N_5877,N_4347,N_4595);
xor U5878 (N_5878,N_4446,N_4943);
and U5879 (N_5879,N_4772,N_4465);
or U5880 (N_5880,N_4340,N_4639);
and U5881 (N_5881,N_4735,N_4440);
and U5882 (N_5882,N_4136,N_4803);
nand U5883 (N_5883,N_4346,N_4846);
nor U5884 (N_5884,N_4432,N_4883);
xor U5885 (N_5885,N_4847,N_4226);
xor U5886 (N_5886,N_4681,N_4383);
and U5887 (N_5887,N_4248,N_4432);
xnor U5888 (N_5888,N_4826,N_4258);
and U5889 (N_5889,N_4874,N_4279);
xor U5890 (N_5890,N_4946,N_4802);
or U5891 (N_5891,N_4398,N_4209);
xor U5892 (N_5892,N_4899,N_4855);
nor U5893 (N_5893,N_4488,N_4372);
or U5894 (N_5894,N_4135,N_4717);
nand U5895 (N_5895,N_4011,N_4157);
nor U5896 (N_5896,N_4150,N_4594);
or U5897 (N_5897,N_4140,N_4633);
or U5898 (N_5898,N_4838,N_4934);
or U5899 (N_5899,N_4028,N_4858);
nand U5900 (N_5900,N_4663,N_4940);
xnor U5901 (N_5901,N_4432,N_4465);
or U5902 (N_5902,N_4941,N_4760);
and U5903 (N_5903,N_4777,N_4018);
nor U5904 (N_5904,N_4623,N_4759);
xnor U5905 (N_5905,N_4960,N_4595);
nand U5906 (N_5906,N_4573,N_4519);
or U5907 (N_5907,N_4776,N_4638);
nor U5908 (N_5908,N_4750,N_4192);
nand U5909 (N_5909,N_4230,N_4939);
or U5910 (N_5910,N_4500,N_4054);
xor U5911 (N_5911,N_4052,N_4370);
xnor U5912 (N_5912,N_4004,N_4795);
and U5913 (N_5913,N_4492,N_4682);
or U5914 (N_5914,N_4992,N_4677);
nor U5915 (N_5915,N_4726,N_4056);
or U5916 (N_5916,N_4555,N_4718);
nor U5917 (N_5917,N_4431,N_4437);
nand U5918 (N_5918,N_4101,N_4596);
nor U5919 (N_5919,N_4174,N_4445);
nand U5920 (N_5920,N_4353,N_4355);
or U5921 (N_5921,N_4600,N_4305);
nor U5922 (N_5922,N_4777,N_4266);
xor U5923 (N_5923,N_4069,N_4578);
nand U5924 (N_5924,N_4900,N_4914);
or U5925 (N_5925,N_4778,N_4513);
and U5926 (N_5926,N_4300,N_4621);
nand U5927 (N_5927,N_4999,N_4616);
and U5928 (N_5928,N_4703,N_4072);
nand U5929 (N_5929,N_4041,N_4841);
and U5930 (N_5930,N_4207,N_4930);
nor U5931 (N_5931,N_4135,N_4915);
nor U5932 (N_5932,N_4237,N_4163);
or U5933 (N_5933,N_4666,N_4653);
or U5934 (N_5934,N_4440,N_4709);
and U5935 (N_5935,N_4030,N_4618);
nand U5936 (N_5936,N_4032,N_4396);
and U5937 (N_5937,N_4279,N_4716);
xor U5938 (N_5938,N_4610,N_4027);
nor U5939 (N_5939,N_4707,N_4520);
nand U5940 (N_5940,N_4298,N_4545);
xnor U5941 (N_5941,N_4202,N_4284);
xnor U5942 (N_5942,N_4215,N_4659);
or U5943 (N_5943,N_4017,N_4776);
xor U5944 (N_5944,N_4108,N_4853);
or U5945 (N_5945,N_4860,N_4290);
xnor U5946 (N_5946,N_4376,N_4711);
or U5947 (N_5947,N_4777,N_4674);
xnor U5948 (N_5948,N_4993,N_4553);
and U5949 (N_5949,N_4704,N_4667);
nand U5950 (N_5950,N_4249,N_4142);
nand U5951 (N_5951,N_4720,N_4843);
or U5952 (N_5952,N_4248,N_4509);
or U5953 (N_5953,N_4540,N_4628);
or U5954 (N_5954,N_4874,N_4394);
nor U5955 (N_5955,N_4907,N_4704);
nand U5956 (N_5956,N_4952,N_4106);
or U5957 (N_5957,N_4340,N_4911);
and U5958 (N_5958,N_4008,N_4415);
or U5959 (N_5959,N_4161,N_4958);
or U5960 (N_5960,N_4519,N_4089);
nand U5961 (N_5961,N_4333,N_4961);
or U5962 (N_5962,N_4495,N_4516);
nor U5963 (N_5963,N_4577,N_4991);
nor U5964 (N_5964,N_4085,N_4332);
xor U5965 (N_5965,N_4463,N_4082);
nand U5966 (N_5966,N_4923,N_4273);
and U5967 (N_5967,N_4067,N_4090);
and U5968 (N_5968,N_4639,N_4542);
and U5969 (N_5969,N_4950,N_4176);
xnor U5970 (N_5970,N_4096,N_4388);
and U5971 (N_5971,N_4100,N_4309);
nor U5972 (N_5972,N_4303,N_4345);
xnor U5973 (N_5973,N_4227,N_4671);
xor U5974 (N_5974,N_4527,N_4936);
nor U5975 (N_5975,N_4912,N_4913);
nand U5976 (N_5976,N_4476,N_4972);
xnor U5977 (N_5977,N_4932,N_4557);
nand U5978 (N_5978,N_4131,N_4014);
nor U5979 (N_5979,N_4342,N_4298);
xor U5980 (N_5980,N_4590,N_4370);
and U5981 (N_5981,N_4090,N_4045);
nor U5982 (N_5982,N_4076,N_4225);
or U5983 (N_5983,N_4772,N_4738);
and U5984 (N_5984,N_4671,N_4754);
and U5985 (N_5985,N_4901,N_4825);
xnor U5986 (N_5986,N_4569,N_4382);
nand U5987 (N_5987,N_4120,N_4881);
or U5988 (N_5988,N_4288,N_4048);
nor U5989 (N_5989,N_4702,N_4475);
or U5990 (N_5990,N_4642,N_4493);
nand U5991 (N_5991,N_4477,N_4661);
nand U5992 (N_5992,N_4212,N_4054);
nor U5993 (N_5993,N_4377,N_4199);
and U5994 (N_5994,N_4861,N_4255);
nand U5995 (N_5995,N_4085,N_4449);
or U5996 (N_5996,N_4251,N_4916);
and U5997 (N_5997,N_4485,N_4330);
nand U5998 (N_5998,N_4912,N_4004);
nand U5999 (N_5999,N_4344,N_4868);
or U6000 (N_6000,N_5895,N_5900);
nor U6001 (N_6001,N_5603,N_5310);
nand U6002 (N_6002,N_5845,N_5926);
and U6003 (N_6003,N_5316,N_5696);
xor U6004 (N_6004,N_5004,N_5920);
nand U6005 (N_6005,N_5114,N_5588);
nand U6006 (N_6006,N_5436,N_5681);
xor U6007 (N_6007,N_5279,N_5257);
nor U6008 (N_6008,N_5499,N_5647);
xnor U6009 (N_6009,N_5817,N_5465);
or U6010 (N_6010,N_5863,N_5783);
or U6011 (N_6011,N_5081,N_5698);
nor U6012 (N_6012,N_5077,N_5398);
nand U6013 (N_6013,N_5837,N_5195);
nor U6014 (N_6014,N_5220,N_5339);
or U6015 (N_6015,N_5556,N_5497);
or U6016 (N_6016,N_5215,N_5075);
and U6017 (N_6017,N_5251,N_5213);
or U6018 (N_6018,N_5986,N_5143);
and U6019 (N_6019,N_5534,N_5169);
nand U6020 (N_6020,N_5221,N_5611);
nor U6021 (N_6021,N_5604,N_5346);
and U6022 (N_6022,N_5761,N_5995);
nor U6023 (N_6023,N_5821,N_5537);
xor U6024 (N_6024,N_5123,N_5711);
or U6025 (N_6025,N_5917,N_5804);
nand U6026 (N_6026,N_5368,N_5846);
or U6027 (N_6027,N_5142,N_5483);
nor U6028 (N_6028,N_5126,N_5854);
or U6029 (N_6029,N_5601,N_5040);
xor U6030 (N_6030,N_5746,N_5009);
and U6031 (N_6031,N_5536,N_5966);
and U6032 (N_6032,N_5940,N_5472);
and U6033 (N_6033,N_5811,N_5411);
and U6034 (N_6034,N_5918,N_5296);
or U6035 (N_6035,N_5041,N_5700);
nor U6036 (N_6036,N_5883,N_5558);
or U6037 (N_6037,N_5214,N_5808);
or U6038 (N_6038,N_5978,N_5999);
nand U6039 (N_6039,N_5701,N_5802);
nor U6040 (N_6040,N_5862,N_5452);
and U6041 (N_6041,N_5450,N_5300);
and U6042 (N_6042,N_5638,N_5786);
and U6043 (N_6043,N_5847,N_5798);
and U6044 (N_6044,N_5779,N_5338);
xor U6045 (N_6045,N_5388,N_5417);
or U6046 (N_6046,N_5823,N_5822);
nor U6047 (N_6047,N_5873,N_5407);
or U6048 (N_6048,N_5810,N_5052);
and U6049 (N_6049,N_5107,N_5663);
xnor U6050 (N_6050,N_5096,N_5939);
nor U6051 (N_6051,N_5841,N_5113);
nor U6052 (N_6052,N_5757,N_5870);
or U6053 (N_6053,N_5580,N_5160);
or U6054 (N_6054,N_5139,N_5941);
or U6055 (N_6055,N_5649,N_5460);
and U6056 (N_6056,N_5894,N_5349);
xnor U6057 (N_6057,N_5959,N_5751);
xor U6058 (N_6058,N_5270,N_5172);
and U6059 (N_6059,N_5832,N_5797);
nand U6060 (N_6060,N_5197,N_5530);
or U6061 (N_6061,N_5313,N_5112);
or U6062 (N_6062,N_5108,N_5631);
or U6063 (N_6063,N_5931,N_5887);
nor U6064 (N_6064,N_5374,N_5188);
xnor U6065 (N_6065,N_5003,N_5692);
or U6066 (N_6066,N_5813,N_5651);
nor U6067 (N_6067,N_5366,N_5442);
xnor U6068 (N_6068,N_5294,N_5623);
nand U6069 (N_6069,N_5382,N_5741);
xnor U6070 (N_6070,N_5031,N_5955);
xnor U6071 (N_6071,N_5210,N_5979);
xnor U6072 (N_6072,N_5010,N_5515);
nand U6073 (N_6073,N_5519,N_5383);
nand U6074 (N_6074,N_5867,N_5104);
nor U6075 (N_6075,N_5250,N_5196);
xnor U6076 (N_6076,N_5618,N_5127);
and U6077 (N_6077,N_5731,N_5019);
and U6078 (N_6078,N_5414,N_5306);
nor U6079 (N_6079,N_5843,N_5889);
or U6080 (N_6080,N_5670,N_5275);
nor U6081 (N_6081,N_5375,N_5583);
nand U6082 (N_6082,N_5456,N_5401);
or U6083 (N_6083,N_5317,N_5790);
nor U6084 (N_6084,N_5975,N_5988);
xnor U6085 (N_6085,N_5860,N_5514);
nor U6086 (N_6086,N_5998,N_5945);
nor U6087 (N_6087,N_5770,N_5523);
or U6088 (N_6088,N_5679,N_5165);
xnor U6089 (N_6089,N_5470,N_5993);
nand U6090 (N_6090,N_5377,N_5181);
or U6091 (N_6091,N_5311,N_5384);
and U6092 (N_6092,N_5665,N_5906);
and U6093 (N_6093,N_5657,N_5147);
nand U6094 (N_6094,N_5690,N_5987);
nor U6095 (N_6095,N_5954,N_5639);
nand U6096 (N_6096,N_5260,N_5119);
and U6097 (N_6097,N_5570,N_5732);
or U6098 (N_6098,N_5239,N_5269);
xor U6099 (N_6099,N_5819,N_5881);
and U6100 (N_6100,N_5896,N_5866);
nor U6101 (N_6101,N_5989,N_5968);
nand U6102 (N_6102,N_5633,N_5569);
nor U6103 (N_6103,N_5551,N_5037);
or U6104 (N_6104,N_5001,N_5946);
xor U6105 (N_6105,N_5319,N_5793);
or U6106 (N_6106,N_5415,N_5496);
and U6107 (N_6107,N_5066,N_5237);
xnor U6108 (N_6108,N_5205,N_5029);
nand U6109 (N_6109,N_5400,N_5421);
nand U6110 (N_6110,N_5035,N_5303);
or U6111 (N_6111,N_5489,N_5728);
nor U6112 (N_6112,N_5632,N_5913);
and U6113 (N_6113,N_5501,N_5722);
nor U6114 (N_6114,N_5555,N_5297);
nor U6115 (N_6115,N_5760,N_5391);
nand U6116 (N_6116,N_5078,N_5535);
xor U6117 (N_6117,N_5613,N_5617);
and U6118 (N_6118,N_5348,N_5115);
and U6119 (N_6119,N_5737,N_5371);
nand U6120 (N_6120,N_5776,N_5805);
nor U6121 (N_6121,N_5413,N_5676);
or U6122 (N_6122,N_5587,N_5667);
xor U6123 (N_6123,N_5516,N_5991);
nor U6124 (N_6124,N_5405,N_5258);
xor U6125 (N_6125,N_5518,N_5595);
and U6126 (N_6126,N_5974,N_5340);
or U6127 (N_6127,N_5399,N_5193);
nand U6128 (N_6128,N_5246,N_5357);
or U6129 (N_6129,N_5106,N_5764);
nand U6130 (N_6130,N_5660,N_5645);
and U6131 (N_6131,N_5255,N_5390);
nand U6132 (N_6132,N_5017,N_5034);
or U6133 (N_6133,N_5186,N_5495);
and U6134 (N_6134,N_5949,N_5206);
nand U6135 (N_6135,N_5047,N_5980);
or U6136 (N_6136,N_5050,N_5884);
nor U6137 (N_6137,N_5185,N_5125);
nand U6138 (N_6138,N_5137,N_5345);
xor U6139 (N_6139,N_5434,N_5691);
and U6140 (N_6140,N_5743,N_5170);
xnor U6141 (N_6141,N_5902,N_5610);
and U6142 (N_6142,N_5528,N_5739);
or U6143 (N_6143,N_5953,N_5468);
nand U6144 (N_6144,N_5678,N_5506);
or U6145 (N_6145,N_5350,N_5818);
nand U6146 (N_6146,N_5164,N_5965);
xor U6147 (N_6147,N_5581,N_5292);
and U6148 (N_6148,N_5634,N_5437);
xor U6149 (N_6149,N_5135,N_5148);
and U6150 (N_6150,N_5560,N_5397);
xor U6151 (N_6151,N_5943,N_5763);
nor U6152 (N_6152,N_5136,N_5750);
or U6153 (N_6153,N_5834,N_5198);
and U6154 (N_6154,N_5262,N_5594);
or U6155 (N_6155,N_5543,N_5283);
nor U6156 (N_6156,N_5507,N_5203);
nor U6157 (N_6157,N_5836,N_5550);
or U6158 (N_6158,N_5418,N_5363);
nor U6159 (N_6159,N_5589,N_5559);
or U6160 (N_6160,N_5911,N_5592);
and U6161 (N_6161,N_5272,N_5539);
xnor U6162 (N_6162,N_5423,N_5608);
nor U6163 (N_6163,N_5074,N_5922);
xnor U6164 (N_6164,N_5322,N_5088);
xnor U6165 (N_6165,N_5504,N_5950);
nand U6166 (N_6166,N_5686,N_5295);
xor U6167 (N_6167,N_5175,N_5231);
nor U6168 (N_6168,N_5782,N_5430);
and U6169 (N_6169,N_5021,N_5276);
or U6170 (N_6170,N_5566,N_5178);
nand U6171 (N_6171,N_5500,N_5564);
nand U6172 (N_6172,N_5488,N_5030);
nand U6173 (N_6173,N_5593,N_5597);
or U6174 (N_6174,N_5409,N_5155);
nor U6175 (N_6175,N_5769,N_5444);
nand U6176 (N_6176,N_5724,N_5734);
and U6177 (N_6177,N_5312,N_5264);
and U6178 (N_6178,N_5152,N_5892);
or U6179 (N_6179,N_5331,N_5915);
and U6180 (N_6180,N_5109,N_5243);
xnor U6181 (N_6181,N_5253,N_5372);
xnor U6182 (N_6182,N_5806,N_5777);
or U6183 (N_6183,N_5302,N_5419);
nor U6184 (N_6184,N_5046,N_5194);
xor U6185 (N_6185,N_5752,N_5526);
xnor U6186 (N_6186,N_5969,N_5932);
nor U6187 (N_6187,N_5102,N_5266);
or U6188 (N_6188,N_5083,N_5352);
and U6189 (N_6189,N_5532,N_5199);
and U6190 (N_6190,N_5730,N_5869);
nand U6191 (N_6191,N_5183,N_5157);
xor U6192 (N_6192,N_5138,N_5598);
xor U6193 (N_6193,N_5621,N_5855);
nor U6194 (N_6194,N_5996,N_5005);
xor U6195 (N_6195,N_5674,N_5053);
xor U6196 (N_6196,N_5494,N_5983);
nand U6197 (N_6197,N_5154,N_5961);
nand U6198 (N_6198,N_5717,N_5548);
nor U6199 (N_6199,N_5838,N_5461);
nor U6200 (N_6200,N_5727,N_5685);
nand U6201 (N_6201,N_5641,N_5844);
nand U6202 (N_6202,N_5957,N_5872);
and U6203 (N_6203,N_5509,N_5803);
xor U6204 (N_6204,N_5874,N_5694);
nor U6205 (N_6205,N_5709,N_5935);
nor U6206 (N_6206,N_5238,N_5742);
nand U6207 (N_6207,N_5893,N_5006);
and U6208 (N_6208,N_5923,N_5947);
and U6209 (N_6209,N_5642,N_5187);
nor U6210 (N_6210,N_5775,N_5341);
or U6211 (N_6211,N_5067,N_5936);
or U6212 (N_6212,N_5023,N_5201);
and U6213 (N_6213,N_5567,N_5851);
nand U6214 (N_6214,N_5145,N_5058);
or U6215 (N_6215,N_5085,N_5982);
or U6216 (N_6216,N_5626,N_5192);
nor U6217 (N_6217,N_5481,N_5099);
and U6218 (N_6218,N_5156,N_5441);
or U6219 (N_6219,N_5619,N_5718);
and U6220 (N_6220,N_5479,N_5373);
nor U6221 (N_6221,N_5616,N_5908);
nor U6222 (N_6222,N_5308,N_5533);
nor U6223 (N_6223,N_5547,N_5609);
nand U6224 (N_6224,N_5379,N_5952);
and U6225 (N_6225,N_5778,N_5265);
or U6226 (N_6226,N_5985,N_5241);
nand U6227 (N_6227,N_5853,N_5655);
or U6228 (N_6228,N_5582,N_5141);
nand U6229 (N_6229,N_5630,N_5622);
and U6230 (N_6230,N_5353,N_5715);
nor U6231 (N_6231,N_5133,N_5242);
or U6232 (N_6232,N_5439,N_5219);
xnor U6233 (N_6233,N_5222,N_5247);
nor U6234 (N_6234,N_5217,N_5216);
or U6235 (N_6235,N_5044,N_5230);
nor U6236 (N_6236,N_5584,N_5487);
and U6237 (N_6237,N_5422,N_5174);
and U6238 (N_6238,N_5771,N_5403);
nor U6239 (N_6239,N_5815,N_5380);
nor U6240 (N_6240,N_5284,N_5024);
or U6241 (N_6241,N_5129,N_5110);
nor U6242 (N_6242,N_5705,N_5459);
xor U6243 (N_6243,N_5561,N_5381);
nand U6244 (N_6244,N_5552,N_5719);
xor U6245 (N_6245,N_5224,N_5944);
xnor U6246 (N_6246,N_5697,N_5288);
and U6247 (N_6247,N_5054,N_5271);
nand U6248 (N_6248,N_5850,N_5827);
or U6249 (N_6249,N_5877,N_5579);
or U6250 (N_6250,N_5791,N_5599);
nand U6251 (N_6251,N_5682,N_5412);
nand U6252 (N_6252,N_5189,N_5449);
nand U6253 (N_6253,N_5321,N_5848);
nor U6254 (N_6254,N_5725,N_5240);
xor U6255 (N_6255,N_5684,N_5045);
nand U6256 (N_6256,N_5491,N_5958);
xnor U6257 (N_6257,N_5209,N_5087);
xor U6258 (N_6258,N_5208,N_5659);
xnor U6259 (N_6259,N_5090,N_5669);
or U6260 (N_6260,N_5858,N_5000);
xnor U6261 (N_6261,N_5480,N_5886);
or U6262 (N_6262,N_5524,N_5788);
and U6263 (N_6263,N_5754,N_5573);
and U6264 (N_6264,N_5773,N_5432);
or U6265 (N_6265,N_5086,N_5478);
nand U6266 (N_6266,N_5182,N_5131);
and U6267 (N_6267,N_5934,N_5972);
nor U6268 (N_6268,N_5644,N_5464);
or U6269 (N_6269,N_5278,N_5320);
nand U6270 (N_6270,N_5702,N_5510);
and U6271 (N_6271,N_5956,N_5713);
and U6272 (N_6272,N_5520,N_5425);
nand U6273 (N_6273,N_5795,N_5544);
or U6274 (N_6274,N_5151,N_5749);
nor U6275 (N_6275,N_5748,N_5180);
nor U6276 (N_6276,N_5190,N_5904);
xor U6277 (N_6277,N_5726,N_5475);
xor U6278 (N_6278,N_5103,N_5080);
xor U6279 (N_6279,N_5720,N_5233);
nand U6280 (N_6280,N_5355,N_5211);
and U6281 (N_6281,N_5245,N_5059);
nand U6282 (N_6282,N_5868,N_5859);
xor U6283 (N_6283,N_5888,N_5281);
nand U6284 (N_6284,N_5508,N_5007);
xor U6285 (N_6285,N_5695,N_5072);
xnor U6286 (N_6286,N_5314,N_5490);
nand U6287 (N_6287,N_5878,N_5293);
nor U6288 (N_6288,N_5554,N_5429);
nand U6289 (N_6289,N_5824,N_5057);
nand U6290 (N_6290,N_5577,N_5140);
and U6291 (N_6291,N_5097,N_5254);
nor U6292 (N_6292,N_5885,N_5410);
xnor U6293 (N_6293,N_5063,N_5658);
nand U6294 (N_6294,N_5937,N_5903);
and U6295 (N_6295,N_5273,N_5636);
or U6296 (N_6296,N_5130,N_5228);
and U6297 (N_6297,N_5071,N_5435);
nor U6298 (N_6298,N_5919,N_5298);
xor U6299 (N_6299,N_5505,N_5688);
xnor U6300 (N_6300,N_5565,N_5683);
nand U6301 (N_6301,N_5916,N_5128);
nor U6302 (N_6302,N_5335,N_5122);
or U6303 (N_6303,N_5627,N_5714);
or U6304 (N_6304,N_5359,N_5234);
nand U6305 (N_6305,N_5799,N_5880);
and U6306 (N_6306,N_5328,N_5406);
nor U6307 (N_6307,N_5898,N_5068);
or U6308 (N_6308,N_5326,N_5531);
xor U6309 (N_6309,N_5899,N_5404);
xor U6310 (N_6310,N_5962,N_5092);
xnor U6311 (N_6311,N_5890,N_5901);
and U6312 (N_6312,N_5280,N_5365);
and U6313 (N_6313,N_5389,N_5291);
or U6314 (N_6314,N_5386,N_5984);
or U6315 (N_6315,N_5236,N_5875);
or U6316 (N_6316,N_5615,N_5132);
or U6317 (N_6317,N_5337,N_5891);
and U6318 (N_6318,N_5438,N_5376);
nor U6319 (N_6319,N_5166,N_5781);
nand U6320 (N_6320,N_5492,N_5716);
xnor U6321 (N_6321,N_5602,N_5814);
or U6322 (N_6322,N_5529,N_5557);
or U6323 (N_6323,N_5424,N_5218);
and U6324 (N_6324,N_5861,N_5008);
nand U6325 (N_6325,N_5290,N_5226);
nand U6326 (N_6326,N_5014,N_5025);
nor U6327 (N_6327,N_5816,N_5204);
and U6328 (N_6328,N_5084,N_5232);
or U6329 (N_6329,N_5740,N_5467);
or U6330 (N_6330,N_5267,N_5428);
and U6331 (N_6331,N_5789,N_5358);
xor U6332 (N_6332,N_5427,N_5022);
or U6333 (N_6333,N_5513,N_5787);
nor U6334 (N_6334,N_5333,N_5012);
or U6335 (N_6335,N_5990,N_5762);
nor U6336 (N_6336,N_5354,N_5876);
nor U6337 (N_6337,N_5336,N_5244);
nor U6338 (N_6338,N_5856,N_5994);
or U6339 (N_6339,N_5591,N_5235);
nand U6340 (N_6340,N_5049,N_5318);
xnor U6341 (N_6341,N_5277,N_5973);
or U6342 (N_6342,N_5699,N_5671);
nand U6343 (N_6343,N_5648,N_5706);
nor U6344 (N_6344,N_5062,N_5538);
xnor U6345 (N_6345,N_5451,N_5735);
nand U6346 (N_6346,N_5356,N_5402);
and U6347 (N_6347,N_5056,N_5252);
nor U6348 (N_6348,N_5738,N_5909);
or U6349 (N_6349,N_5307,N_5600);
nand U6350 (N_6350,N_5073,N_5522);
and U6351 (N_6351,N_5553,N_5677);
nand U6352 (N_6352,N_5563,N_5925);
nand U6353 (N_6353,N_5612,N_5879);
and U6354 (N_6354,N_5287,N_5723);
nand U6355 (N_6355,N_5202,N_5680);
xor U6356 (N_6356,N_5347,N_5360);
xnor U6357 (N_6357,N_5447,N_5042);
nor U6358 (N_6358,N_5094,N_5482);
nand U6359 (N_6359,N_5431,N_5650);
or U6360 (N_6360,N_5575,N_5159);
and U6361 (N_6361,N_5249,N_5079);
nand U6362 (N_6362,N_5330,N_5016);
or U6363 (N_6363,N_5800,N_5324);
or U6364 (N_6364,N_5091,N_5309);
nand U6365 (N_6365,N_5511,N_5652);
xor U6366 (N_6366,N_5392,N_5469);
nand U6367 (N_6367,N_5905,N_5020);
and U6368 (N_6368,N_5656,N_5334);
and U6369 (N_6369,N_5525,N_5687);
nand U6370 (N_6370,N_5289,N_5527);
or U6371 (N_6371,N_5614,N_5733);
or U6372 (N_6372,N_5766,N_5512);
xor U6373 (N_6373,N_5268,N_5301);
nand U6374 (N_6374,N_5394,N_5036);
or U6375 (N_6375,N_5585,N_5924);
and U6376 (N_6376,N_5486,N_5117);
nor U6377 (N_6377,N_5503,N_5013);
xnor U6378 (N_6378,N_5689,N_5546);
nor U6379 (N_6379,N_5158,N_5395);
nand U6380 (N_6380,N_5794,N_5455);
xnor U6381 (N_6381,N_5426,N_5664);
xnor U6382 (N_6382,N_5828,N_5493);
or U6383 (N_6383,N_5342,N_5369);
nor U6384 (N_6384,N_5545,N_5261);
or U6385 (N_6385,N_5625,N_5453);
xnor U6386 (N_6386,N_5286,N_5849);
nor U6387 (N_6387,N_5517,N_5171);
nand U6388 (N_6388,N_5105,N_5248);
and U6389 (N_6389,N_5606,N_5736);
nand U6390 (N_6390,N_5666,N_5223);
nor U6391 (N_6391,N_5329,N_5089);
nor U6392 (N_6392,N_5256,N_5484);
or U6393 (N_6393,N_5605,N_5011);
or U6394 (N_6394,N_5571,N_5938);
nand U6395 (N_6395,N_5144,N_5076);
nand U6396 (N_6396,N_5361,N_5176);
nand U6397 (N_6397,N_5095,N_5977);
xor U6398 (N_6398,N_5229,N_5440);
and U6399 (N_6399,N_5263,N_5864);
xnor U6400 (N_6400,N_5897,N_5445);
and U6401 (N_6401,N_5963,N_5976);
nor U6402 (N_6402,N_5929,N_5745);
or U6403 (N_6403,N_5082,N_5471);
nand U6404 (N_6404,N_5928,N_5408);
nor U6405 (N_6405,N_5367,N_5474);
nand U6406 (N_6406,N_5637,N_5807);
or U6407 (N_6407,N_5458,N_5729);
or U6408 (N_6408,N_5344,N_5712);
nand U6409 (N_6409,N_5704,N_5948);
nor U6410 (N_6410,N_5043,N_5462);
nand U6411 (N_6411,N_5362,N_5907);
nand U6412 (N_6412,N_5784,N_5032);
and U6413 (N_6413,N_5162,N_5967);
and U6414 (N_6414,N_5765,N_5852);
xnor U6415 (N_6415,N_5443,N_5672);
and U6416 (N_6416,N_5116,N_5590);
nand U6417 (N_6417,N_5673,N_5812);
nand U6418 (N_6418,N_5315,N_5753);
xor U6419 (N_6419,N_5039,N_5387);
or U6420 (N_6420,N_5351,N_5792);
and U6421 (N_6421,N_5146,N_5393);
nand U6422 (N_6422,N_5758,N_5572);
nor U6423 (N_6423,N_5149,N_5912);
nor U6424 (N_6424,N_5259,N_5343);
xnor U6425 (N_6425,N_5064,N_5780);
nor U6426 (N_6426,N_5646,N_5153);
xor U6427 (N_6427,N_5774,N_5997);
and U6428 (N_6428,N_5747,N_5981);
and U6429 (N_6429,N_5839,N_5018);
or U6430 (N_6430,N_5693,N_5454);
nand U6431 (N_6431,N_5274,N_5457);
or U6432 (N_6432,N_5930,N_5477);
xor U6433 (N_6433,N_5364,N_5173);
nor U6434 (N_6434,N_5596,N_5661);
nor U6435 (N_6435,N_5653,N_5721);
nor U6436 (N_6436,N_5755,N_5055);
nand U6437 (N_6437,N_5654,N_5829);
and U6438 (N_6438,N_5772,N_5675);
nand U6439 (N_6439,N_5038,N_5448);
nor U6440 (N_6440,N_5927,N_5285);
or U6441 (N_6441,N_5446,N_5433);
nor U6442 (N_6442,N_5325,N_5177);
and U6443 (N_6443,N_5970,N_5065);
or U6444 (N_6444,N_5942,N_5466);
nand U6445 (N_6445,N_5098,N_5420);
xor U6446 (N_6446,N_5502,N_5871);
nand U6447 (N_6447,N_5028,N_5212);
and U6448 (N_6448,N_5168,N_5826);
nand U6449 (N_6449,N_5620,N_5910);
xnor U6450 (N_6450,N_5282,N_5161);
nand U6451 (N_6451,N_5227,N_5992);
or U6452 (N_6452,N_5759,N_5586);
xnor U6453 (N_6453,N_5498,N_5323);
nor U6454 (N_6454,N_5184,N_5299);
and U6455 (N_6455,N_5703,N_5026);
nor U6456 (N_6456,N_5485,N_5207);
nand U6457 (N_6457,N_5370,N_5830);
and U6458 (N_6458,N_5416,N_5048);
nand U6459 (N_6459,N_5069,N_5578);
or U6460 (N_6460,N_5002,N_5396);
nand U6461 (N_6461,N_5820,N_5327);
nor U6462 (N_6462,N_5574,N_5027);
or U6463 (N_6463,N_5476,N_5629);
nand U6464 (N_6464,N_5120,N_5121);
xnor U6465 (N_6465,N_5960,N_5060);
xor U6466 (N_6466,N_5635,N_5576);
nor U6467 (N_6467,N_5840,N_5521);
nor U6468 (N_6468,N_5549,N_5015);
nand U6469 (N_6469,N_5708,N_5707);
xor U6470 (N_6470,N_5191,N_5796);
nor U6471 (N_6471,N_5179,N_5882);
xor U6472 (N_6472,N_5785,N_5541);
xor U6473 (N_6473,N_5835,N_5305);
nor U6474 (N_6474,N_5385,N_5225);
nand U6475 (N_6475,N_5767,N_5825);
or U6476 (N_6476,N_5756,N_5833);
and U6477 (N_6477,N_5857,N_5033);
nor U6478 (N_6478,N_5051,N_5163);
xnor U6479 (N_6479,N_5842,N_5865);
xor U6480 (N_6480,N_5951,N_5061);
nor U6481 (N_6481,N_5914,N_5662);
nand U6482 (N_6482,N_5473,N_5101);
and U6483 (N_6483,N_5562,N_5628);
xnor U6484 (N_6484,N_5921,N_5304);
nor U6485 (N_6485,N_5964,N_5200);
or U6486 (N_6486,N_5124,N_5542);
xor U6487 (N_6487,N_5768,N_5134);
nor U6488 (N_6488,N_5568,N_5100);
nand U6489 (N_6489,N_5643,N_5744);
nor U6490 (N_6490,N_5332,N_5150);
xor U6491 (N_6491,N_5118,N_5378);
and U6492 (N_6492,N_5809,N_5801);
and U6493 (N_6493,N_5463,N_5607);
and U6494 (N_6494,N_5710,N_5831);
xor U6495 (N_6495,N_5070,N_5971);
xor U6496 (N_6496,N_5640,N_5624);
nor U6497 (N_6497,N_5668,N_5540);
nor U6498 (N_6498,N_5111,N_5933);
nor U6499 (N_6499,N_5093,N_5167);
or U6500 (N_6500,N_5776,N_5179);
xnor U6501 (N_6501,N_5831,N_5133);
or U6502 (N_6502,N_5069,N_5007);
and U6503 (N_6503,N_5815,N_5817);
and U6504 (N_6504,N_5506,N_5601);
or U6505 (N_6505,N_5258,N_5205);
nor U6506 (N_6506,N_5729,N_5010);
xor U6507 (N_6507,N_5604,N_5498);
and U6508 (N_6508,N_5911,N_5212);
nand U6509 (N_6509,N_5584,N_5694);
nand U6510 (N_6510,N_5785,N_5261);
nor U6511 (N_6511,N_5771,N_5281);
nor U6512 (N_6512,N_5456,N_5682);
and U6513 (N_6513,N_5174,N_5539);
nand U6514 (N_6514,N_5279,N_5876);
nand U6515 (N_6515,N_5939,N_5712);
nor U6516 (N_6516,N_5700,N_5100);
and U6517 (N_6517,N_5586,N_5081);
and U6518 (N_6518,N_5552,N_5544);
nand U6519 (N_6519,N_5956,N_5817);
nand U6520 (N_6520,N_5645,N_5003);
nand U6521 (N_6521,N_5288,N_5715);
xor U6522 (N_6522,N_5228,N_5983);
nand U6523 (N_6523,N_5191,N_5000);
and U6524 (N_6524,N_5881,N_5471);
xnor U6525 (N_6525,N_5034,N_5418);
xnor U6526 (N_6526,N_5946,N_5338);
nor U6527 (N_6527,N_5041,N_5059);
and U6528 (N_6528,N_5058,N_5142);
nand U6529 (N_6529,N_5699,N_5683);
xnor U6530 (N_6530,N_5061,N_5306);
xor U6531 (N_6531,N_5449,N_5565);
nand U6532 (N_6532,N_5227,N_5869);
nor U6533 (N_6533,N_5015,N_5709);
and U6534 (N_6534,N_5350,N_5857);
nor U6535 (N_6535,N_5066,N_5718);
and U6536 (N_6536,N_5473,N_5474);
and U6537 (N_6537,N_5032,N_5430);
or U6538 (N_6538,N_5694,N_5534);
xor U6539 (N_6539,N_5152,N_5284);
xnor U6540 (N_6540,N_5023,N_5127);
and U6541 (N_6541,N_5014,N_5569);
nor U6542 (N_6542,N_5604,N_5295);
nand U6543 (N_6543,N_5156,N_5727);
nor U6544 (N_6544,N_5264,N_5191);
xnor U6545 (N_6545,N_5921,N_5680);
nor U6546 (N_6546,N_5110,N_5549);
nand U6547 (N_6547,N_5444,N_5805);
or U6548 (N_6548,N_5360,N_5418);
and U6549 (N_6549,N_5293,N_5988);
xnor U6550 (N_6550,N_5972,N_5892);
and U6551 (N_6551,N_5939,N_5906);
xor U6552 (N_6552,N_5643,N_5799);
nand U6553 (N_6553,N_5323,N_5435);
xnor U6554 (N_6554,N_5965,N_5709);
nand U6555 (N_6555,N_5174,N_5034);
nor U6556 (N_6556,N_5356,N_5853);
or U6557 (N_6557,N_5194,N_5657);
or U6558 (N_6558,N_5629,N_5135);
nor U6559 (N_6559,N_5076,N_5740);
xnor U6560 (N_6560,N_5483,N_5745);
nand U6561 (N_6561,N_5121,N_5449);
xnor U6562 (N_6562,N_5632,N_5607);
nor U6563 (N_6563,N_5520,N_5726);
nand U6564 (N_6564,N_5440,N_5910);
and U6565 (N_6565,N_5648,N_5036);
xnor U6566 (N_6566,N_5345,N_5944);
nand U6567 (N_6567,N_5622,N_5709);
or U6568 (N_6568,N_5410,N_5023);
or U6569 (N_6569,N_5579,N_5495);
nor U6570 (N_6570,N_5021,N_5414);
nor U6571 (N_6571,N_5561,N_5765);
and U6572 (N_6572,N_5692,N_5544);
nor U6573 (N_6573,N_5629,N_5372);
xor U6574 (N_6574,N_5666,N_5588);
nor U6575 (N_6575,N_5523,N_5544);
nand U6576 (N_6576,N_5750,N_5295);
or U6577 (N_6577,N_5411,N_5750);
nand U6578 (N_6578,N_5983,N_5244);
nand U6579 (N_6579,N_5895,N_5113);
nand U6580 (N_6580,N_5610,N_5782);
and U6581 (N_6581,N_5965,N_5322);
and U6582 (N_6582,N_5877,N_5020);
or U6583 (N_6583,N_5075,N_5717);
nand U6584 (N_6584,N_5800,N_5478);
nor U6585 (N_6585,N_5498,N_5320);
or U6586 (N_6586,N_5973,N_5096);
xnor U6587 (N_6587,N_5232,N_5537);
nor U6588 (N_6588,N_5214,N_5428);
or U6589 (N_6589,N_5427,N_5396);
or U6590 (N_6590,N_5849,N_5962);
or U6591 (N_6591,N_5708,N_5518);
xnor U6592 (N_6592,N_5815,N_5560);
xnor U6593 (N_6593,N_5478,N_5643);
nand U6594 (N_6594,N_5589,N_5852);
nand U6595 (N_6595,N_5234,N_5873);
nor U6596 (N_6596,N_5528,N_5524);
or U6597 (N_6597,N_5920,N_5838);
nor U6598 (N_6598,N_5343,N_5496);
or U6599 (N_6599,N_5827,N_5349);
or U6600 (N_6600,N_5488,N_5425);
xnor U6601 (N_6601,N_5284,N_5352);
or U6602 (N_6602,N_5253,N_5558);
or U6603 (N_6603,N_5605,N_5729);
nor U6604 (N_6604,N_5381,N_5712);
nor U6605 (N_6605,N_5220,N_5830);
and U6606 (N_6606,N_5005,N_5697);
nor U6607 (N_6607,N_5940,N_5294);
nand U6608 (N_6608,N_5400,N_5066);
or U6609 (N_6609,N_5232,N_5911);
and U6610 (N_6610,N_5278,N_5596);
and U6611 (N_6611,N_5735,N_5474);
nand U6612 (N_6612,N_5725,N_5318);
or U6613 (N_6613,N_5645,N_5707);
xor U6614 (N_6614,N_5747,N_5437);
and U6615 (N_6615,N_5081,N_5656);
nor U6616 (N_6616,N_5875,N_5940);
or U6617 (N_6617,N_5315,N_5502);
or U6618 (N_6618,N_5662,N_5949);
nor U6619 (N_6619,N_5273,N_5783);
nand U6620 (N_6620,N_5363,N_5197);
or U6621 (N_6621,N_5047,N_5777);
nand U6622 (N_6622,N_5595,N_5922);
xor U6623 (N_6623,N_5862,N_5272);
and U6624 (N_6624,N_5094,N_5917);
or U6625 (N_6625,N_5682,N_5226);
and U6626 (N_6626,N_5555,N_5927);
nor U6627 (N_6627,N_5197,N_5152);
nor U6628 (N_6628,N_5008,N_5771);
nor U6629 (N_6629,N_5434,N_5984);
nand U6630 (N_6630,N_5231,N_5460);
or U6631 (N_6631,N_5218,N_5530);
nor U6632 (N_6632,N_5274,N_5587);
nor U6633 (N_6633,N_5166,N_5585);
and U6634 (N_6634,N_5652,N_5741);
or U6635 (N_6635,N_5274,N_5103);
nor U6636 (N_6636,N_5524,N_5158);
and U6637 (N_6637,N_5430,N_5862);
or U6638 (N_6638,N_5139,N_5951);
xor U6639 (N_6639,N_5811,N_5007);
or U6640 (N_6640,N_5981,N_5662);
xor U6641 (N_6641,N_5458,N_5925);
and U6642 (N_6642,N_5057,N_5523);
or U6643 (N_6643,N_5235,N_5562);
or U6644 (N_6644,N_5086,N_5261);
nor U6645 (N_6645,N_5571,N_5819);
nor U6646 (N_6646,N_5317,N_5250);
xnor U6647 (N_6647,N_5867,N_5542);
nor U6648 (N_6648,N_5386,N_5301);
and U6649 (N_6649,N_5882,N_5056);
or U6650 (N_6650,N_5922,N_5877);
and U6651 (N_6651,N_5856,N_5728);
or U6652 (N_6652,N_5916,N_5527);
or U6653 (N_6653,N_5526,N_5756);
and U6654 (N_6654,N_5189,N_5254);
nor U6655 (N_6655,N_5665,N_5961);
or U6656 (N_6656,N_5826,N_5511);
xor U6657 (N_6657,N_5353,N_5817);
xor U6658 (N_6658,N_5535,N_5745);
nor U6659 (N_6659,N_5409,N_5328);
nor U6660 (N_6660,N_5407,N_5672);
nand U6661 (N_6661,N_5584,N_5585);
nand U6662 (N_6662,N_5138,N_5316);
nand U6663 (N_6663,N_5560,N_5174);
and U6664 (N_6664,N_5356,N_5935);
and U6665 (N_6665,N_5452,N_5715);
or U6666 (N_6666,N_5095,N_5433);
nand U6667 (N_6667,N_5910,N_5811);
nand U6668 (N_6668,N_5296,N_5092);
and U6669 (N_6669,N_5624,N_5697);
nand U6670 (N_6670,N_5294,N_5688);
xor U6671 (N_6671,N_5117,N_5746);
nor U6672 (N_6672,N_5109,N_5526);
and U6673 (N_6673,N_5086,N_5810);
nand U6674 (N_6674,N_5941,N_5447);
xor U6675 (N_6675,N_5923,N_5326);
and U6676 (N_6676,N_5670,N_5106);
xor U6677 (N_6677,N_5817,N_5303);
or U6678 (N_6678,N_5606,N_5763);
and U6679 (N_6679,N_5929,N_5774);
nand U6680 (N_6680,N_5539,N_5820);
nand U6681 (N_6681,N_5679,N_5214);
xnor U6682 (N_6682,N_5599,N_5220);
or U6683 (N_6683,N_5396,N_5480);
nand U6684 (N_6684,N_5836,N_5241);
and U6685 (N_6685,N_5030,N_5954);
nor U6686 (N_6686,N_5878,N_5934);
or U6687 (N_6687,N_5831,N_5322);
nor U6688 (N_6688,N_5795,N_5730);
xor U6689 (N_6689,N_5543,N_5198);
and U6690 (N_6690,N_5243,N_5530);
and U6691 (N_6691,N_5742,N_5035);
nand U6692 (N_6692,N_5000,N_5022);
or U6693 (N_6693,N_5614,N_5047);
nor U6694 (N_6694,N_5972,N_5359);
nor U6695 (N_6695,N_5147,N_5664);
xnor U6696 (N_6696,N_5703,N_5795);
nor U6697 (N_6697,N_5932,N_5876);
nor U6698 (N_6698,N_5381,N_5882);
nand U6699 (N_6699,N_5246,N_5347);
and U6700 (N_6700,N_5174,N_5985);
nand U6701 (N_6701,N_5166,N_5233);
nand U6702 (N_6702,N_5809,N_5510);
nand U6703 (N_6703,N_5895,N_5691);
or U6704 (N_6704,N_5173,N_5715);
nand U6705 (N_6705,N_5662,N_5845);
and U6706 (N_6706,N_5527,N_5595);
xor U6707 (N_6707,N_5908,N_5623);
and U6708 (N_6708,N_5725,N_5192);
or U6709 (N_6709,N_5646,N_5599);
or U6710 (N_6710,N_5918,N_5815);
nand U6711 (N_6711,N_5590,N_5218);
xor U6712 (N_6712,N_5915,N_5116);
nor U6713 (N_6713,N_5177,N_5818);
and U6714 (N_6714,N_5327,N_5895);
or U6715 (N_6715,N_5860,N_5878);
or U6716 (N_6716,N_5622,N_5737);
nand U6717 (N_6717,N_5052,N_5870);
and U6718 (N_6718,N_5304,N_5983);
and U6719 (N_6719,N_5447,N_5126);
nor U6720 (N_6720,N_5912,N_5497);
and U6721 (N_6721,N_5926,N_5581);
nand U6722 (N_6722,N_5097,N_5757);
and U6723 (N_6723,N_5513,N_5909);
xor U6724 (N_6724,N_5254,N_5224);
xnor U6725 (N_6725,N_5734,N_5927);
or U6726 (N_6726,N_5020,N_5042);
xnor U6727 (N_6727,N_5703,N_5459);
or U6728 (N_6728,N_5603,N_5772);
or U6729 (N_6729,N_5481,N_5896);
nand U6730 (N_6730,N_5733,N_5553);
or U6731 (N_6731,N_5589,N_5616);
and U6732 (N_6732,N_5467,N_5580);
nand U6733 (N_6733,N_5678,N_5749);
nand U6734 (N_6734,N_5262,N_5743);
and U6735 (N_6735,N_5131,N_5000);
nand U6736 (N_6736,N_5569,N_5235);
xor U6737 (N_6737,N_5809,N_5460);
or U6738 (N_6738,N_5667,N_5227);
or U6739 (N_6739,N_5373,N_5131);
nand U6740 (N_6740,N_5691,N_5502);
and U6741 (N_6741,N_5304,N_5409);
xor U6742 (N_6742,N_5297,N_5598);
nand U6743 (N_6743,N_5304,N_5183);
nor U6744 (N_6744,N_5416,N_5875);
nor U6745 (N_6745,N_5816,N_5804);
and U6746 (N_6746,N_5818,N_5629);
nand U6747 (N_6747,N_5546,N_5916);
nand U6748 (N_6748,N_5436,N_5035);
and U6749 (N_6749,N_5690,N_5909);
and U6750 (N_6750,N_5280,N_5001);
xor U6751 (N_6751,N_5216,N_5720);
nand U6752 (N_6752,N_5225,N_5339);
or U6753 (N_6753,N_5455,N_5043);
or U6754 (N_6754,N_5231,N_5523);
xnor U6755 (N_6755,N_5283,N_5591);
nor U6756 (N_6756,N_5718,N_5730);
nor U6757 (N_6757,N_5430,N_5527);
nand U6758 (N_6758,N_5592,N_5074);
nand U6759 (N_6759,N_5918,N_5907);
and U6760 (N_6760,N_5310,N_5891);
or U6761 (N_6761,N_5631,N_5080);
nor U6762 (N_6762,N_5782,N_5401);
nand U6763 (N_6763,N_5958,N_5781);
and U6764 (N_6764,N_5444,N_5185);
xnor U6765 (N_6765,N_5894,N_5642);
and U6766 (N_6766,N_5397,N_5012);
or U6767 (N_6767,N_5270,N_5811);
nand U6768 (N_6768,N_5306,N_5016);
nor U6769 (N_6769,N_5706,N_5393);
and U6770 (N_6770,N_5653,N_5602);
nand U6771 (N_6771,N_5293,N_5850);
or U6772 (N_6772,N_5696,N_5347);
and U6773 (N_6773,N_5750,N_5438);
nand U6774 (N_6774,N_5696,N_5587);
xnor U6775 (N_6775,N_5659,N_5845);
and U6776 (N_6776,N_5992,N_5852);
or U6777 (N_6777,N_5928,N_5635);
xnor U6778 (N_6778,N_5910,N_5797);
nand U6779 (N_6779,N_5627,N_5147);
nand U6780 (N_6780,N_5408,N_5481);
nand U6781 (N_6781,N_5505,N_5908);
and U6782 (N_6782,N_5365,N_5167);
or U6783 (N_6783,N_5035,N_5163);
or U6784 (N_6784,N_5008,N_5775);
xnor U6785 (N_6785,N_5788,N_5848);
xnor U6786 (N_6786,N_5055,N_5135);
or U6787 (N_6787,N_5012,N_5774);
nand U6788 (N_6788,N_5950,N_5633);
xnor U6789 (N_6789,N_5240,N_5548);
xor U6790 (N_6790,N_5960,N_5801);
nor U6791 (N_6791,N_5444,N_5973);
nand U6792 (N_6792,N_5050,N_5003);
nand U6793 (N_6793,N_5027,N_5642);
nand U6794 (N_6794,N_5576,N_5370);
nand U6795 (N_6795,N_5156,N_5256);
nor U6796 (N_6796,N_5928,N_5280);
xnor U6797 (N_6797,N_5121,N_5165);
or U6798 (N_6798,N_5797,N_5976);
nor U6799 (N_6799,N_5556,N_5524);
nor U6800 (N_6800,N_5659,N_5590);
xnor U6801 (N_6801,N_5824,N_5362);
and U6802 (N_6802,N_5430,N_5861);
or U6803 (N_6803,N_5847,N_5281);
or U6804 (N_6804,N_5738,N_5542);
nand U6805 (N_6805,N_5602,N_5315);
xor U6806 (N_6806,N_5504,N_5483);
and U6807 (N_6807,N_5709,N_5961);
or U6808 (N_6808,N_5646,N_5015);
and U6809 (N_6809,N_5811,N_5452);
nand U6810 (N_6810,N_5989,N_5855);
or U6811 (N_6811,N_5116,N_5837);
and U6812 (N_6812,N_5492,N_5944);
nand U6813 (N_6813,N_5497,N_5673);
or U6814 (N_6814,N_5486,N_5082);
nand U6815 (N_6815,N_5105,N_5517);
xnor U6816 (N_6816,N_5108,N_5690);
and U6817 (N_6817,N_5734,N_5019);
and U6818 (N_6818,N_5985,N_5678);
or U6819 (N_6819,N_5686,N_5693);
or U6820 (N_6820,N_5770,N_5020);
nand U6821 (N_6821,N_5609,N_5191);
or U6822 (N_6822,N_5488,N_5024);
nand U6823 (N_6823,N_5142,N_5435);
nor U6824 (N_6824,N_5430,N_5454);
nor U6825 (N_6825,N_5896,N_5564);
nand U6826 (N_6826,N_5690,N_5978);
nor U6827 (N_6827,N_5835,N_5529);
nand U6828 (N_6828,N_5819,N_5500);
nand U6829 (N_6829,N_5883,N_5651);
nand U6830 (N_6830,N_5960,N_5101);
xor U6831 (N_6831,N_5194,N_5638);
nor U6832 (N_6832,N_5289,N_5629);
xor U6833 (N_6833,N_5486,N_5654);
nand U6834 (N_6834,N_5371,N_5618);
or U6835 (N_6835,N_5734,N_5567);
and U6836 (N_6836,N_5606,N_5256);
nor U6837 (N_6837,N_5469,N_5529);
xnor U6838 (N_6838,N_5852,N_5542);
xnor U6839 (N_6839,N_5513,N_5297);
and U6840 (N_6840,N_5304,N_5973);
nand U6841 (N_6841,N_5533,N_5317);
nand U6842 (N_6842,N_5909,N_5047);
and U6843 (N_6843,N_5643,N_5185);
or U6844 (N_6844,N_5104,N_5078);
nor U6845 (N_6845,N_5695,N_5499);
and U6846 (N_6846,N_5154,N_5482);
or U6847 (N_6847,N_5234,N_5303);
and U6848 (N_6848,N_5621,N_5648);
nand U6849 (N_6849,N_5802,N_5920);
xor U6850 (N_6850,N_5611,N_5792);
or U6851 (N_6851,N_5203,N_5807);
or U6852 (N_6852,N_5281,N_5593);
xor U6853 (N_6853,N_5191,N_5184);
xnor U6854 (N_6854,N_5928,N_5511);
nand U6855 (N_6855,N_5307,N_5567);
xnor U6856 (N_6856,N_5433,N_5511);
nor U6857 (N_6857,N_5592,N_5323);
or U6858 (N_6858,N_5486,N_5837);
xnor U6859 (N_6859,N_5122,N_5251);
nand U6860 (N_6860,N_5940,N_5122);
nand U6861 (N_6861,N_5892,N_5675);
nor U6862 (N_6862,N_5356,N_5229);
nor U6863 (N_6863,N_5785,N_5204);
xor U6864 (N_6864,N_5383,N_5858);
xor U6865 (N_6865,N_5622,N_5784);
or U6866 (N_6866,N_5976,N_5026);
and U6867 (N_6867,N_5315,N_5891);
nor U6868 (N_6868,N_5811,N_5356);
or U6869 (N_6869,N_5792,N_5769);
nand U6870 (N_6870,N_5389,N_5729);
or U6871 (N_6871,N_5177,N_5271);
nand U6872 (N_6872,N_5239,N_5146);
xnor U6873 (N_6873,N_5917,N_5414);
nand U6874 (N_6874,N_5125,N_5328);
nand U6875 (N_6875,N_5637,N_5971);
nand U6876 (N_6876,N_5227,N_5832);
nand U6877 (N_6877,N_5037,N_5522);
xnor U6878 (N_6878,N_5229,N_5644);
and U6879 (N_6879,N_5620,N_5887);
nand U6880 (N_6880,N_5558,N_5086);
or U6881 (N_6881,N_5704,N_5035);
or U6882 (N_6882,N_5406,N_5094);
nand U6883 (N_6883,N_5716,N_5348);
and U6884 (N_6884,N_5681,N_5369);
xnor U6885 (N_6885,N_5468,N_5164);
nor U6886 (N_6886,N_5962,N_5281);
or U6887 (N_6887,N_5449,N_5045);
nor U6888 (N_6888,N_5954,N_5824);
nand U6889 (N_6889,N_5861,N_5800);
nand U6890 (N_6890,N_5174,N_5755);
nand U6891 (N_6891,N_5634,N_5787);
and U6892 (N_6892,N_5470,N_5456);
and U6893 (N_6893,N_5687,N_5154);
nand U6894 (N_6894,N_5969,N_5259);
xor U6895 (N_6895,N_5872,N_5208);
or U6896 (N_6896,N_5554,N_5458);
and U6897 (N_6897,N_5641,N_5346);
nor U6898 (N_6898,N_5055,N_5392);
nor U6899 (N_6899,N_5651,N_5406);
and U6900 (N_6900,N_5413,N_5593);
and U6901 (N_6901,N_5246,N_5327);
and U6902 (N_6902,N_5847,N_5536);
or U6903 (N_6903,N_5442,N_5646);
nand U6904 (N_6904,N_5094,N_5924);
and U6905 (N_6905,N_5737,N_5013);
or U6906 (N_6906,N_5313,N_5850);
nand U6907 (N_6907,N_5846,N_5412);
nor U6908 (N_6908,N_5797,N_5834);
and U6909 (N_6909,N_5723,N_5702);
and U6910 (N_6910,N_5765,N_5476);
nand U6911 (N_6911,N_5601,N_5152);
nand U6912 (N_6912,N_5587,N_5336);
xor U6913 (N_6913,N_5599,N_5688);
or U6914 (N_6914,N_5471,N_5696);
or U6915 (N_6915,N_5048,N_5708);
nor U6916 (N_6916,N_5375,N_5026);
nor U6917 (N_6917,N_5490,N_5450);
nand U6918 (N_6918,N_5283,N_5267);
or U6919 (N_6919,N_5070,N_5716);
nor U6920 (N_6920,N_5715,N_5386);
nor U6921 (N_6921,N_5020,N_5740);
or U6922 (N_6922,N_5803,N_5253);
and U6923 (N_6923,N_5535,N_5474);
and U6924 (N_6924,N_5839,N_5003);
nor U6925 (N_6925,N_5482,N_5815);
or U6926 (N_6926,N_5727,N_5770);
or U6927 (N_6927,N_5583,N_5758);
and U6928 (N_6928,N_5404,N_5302);
and U6929 (N_6929,N_5998,N_5044);
or U6930 (N_6930,N_5784,N_5490);
or U6931 (N_6931,N_5645,N_5087);
nor U6932 (N_6932,N_5115,N_5790);
and U6933 (N_6933,N_5821,N_5786);
or U6934 (N_6934,N_5332,N_5957);
and U6935 (N_6935,N_5114,N_5013);
or U6936 (N_6936,N_5464,N_5954);
nor U6937 (N_6937,N_5426,N_5939);
xor U6938 (N_6938,N_5232,N_5801);
nand U6939 (N_6939,N_5104,N_5453);
or U6940 (N_6940,N_5354,N_5441);
and U6941 (N_6941,N_5440,N_5435);
or U6942 (N_6942,N_5126,N_5365);
or U6943 (N_6943,N_5138,N_5629);
or U6944 (N_6944,N_5720,N_5204);
and U6945 (N_6945,N_5902,N_5630);
xnor U6946 (N_6946,N_5788,N_5859);
nor U6947 (N_6947,N_5173,N_5880);
nor U6948 (N_6948,N_5302,N_5548);
nand U6949 (N_6949,N_5282,N_5992);
nand U6950 (N_6950,N_5564,N_5991);
nand U6951 (N_6951,N_5161,N_5520);
nor U6952 (N_6952,N_5998,N_5942);
or U6953 (N_6953,N_5958,N_5186);
nor U6954 (N_6954,N_5583,N_5030);
and U6955 (N_6955,N_5116,N_5694);
and U6956 (N_6956,N_5653,N_5773);
and U6957 (N_6957,N_5162,N_5937);
nor U6958 (N_6958,N_5285,N_5255);
xor U6959 (N_6959,N_5210,N_5192);
and U6960 (N_6960,N_5139,N_5394);
xnor U6961 (N_6961,N_5376,N_5385);
xor U6962 (N_6962,N_5224,N_5239);
xnor U6963 (N_6963,N_5248,N_5882);
or U6964 (N_6964,N_5800,N_5169);
xor U6965 (N_6965,N_5279,N_5124);
xnor U6966 (N_6966,N_5203,N_5909);
xor U6967 (N_6967,N_5224,N_5255);
nor U6968 (N_6968,N_5679,N_5004);
or U6969 (N_6969,N_5636,N_5805);
nor U6970 (N_6970,N_5258,N_5415);
xor U6971 (N_6971,N_5660,N_5701);
nor U6972 (N_6972,N_5786,N_5557);
nand U6973 (N_6973,N_5748,N_5816);
xnor U6974 (N_6974,N_5030,N_5282);
nand U6975 (N_6975,N_5294,N_5608);
and U6976 (N_6976,N_5192,N_5792);
or U6977 (N_6977,N_5328,N_5585);
xnor U6978 (N_6978,N_5735,N_5688);
or U6979 (N_6979,N_5836,N_5841);
or U6980 (N_6980,N_5027,N_5306);
nor U6981 (N_6981,N_5164,N_5714);
and U6982 (N_6982,N_5974,N_5830);
and U6983 (N_6983,N_5925,N_5780);
xor U6984 (N_6984,N_5769,N_5111);
nor U6985 (N_6985,N_5634,N_5338);
nand U6986 (N_6986,N_5483,N_5562);
nand U6987 (N_6987,N_5709,N_5029);
or U6988 (N_6988,N_5958,N_5631);
and U6989 (N_6989,N_5086,N_5063);
nand U6990 (N_6990,N_5663,N_5850);
nor U6991 (N_6991,N_5408,N_5575);
or U6992 (N_6992,N_5739,N_5485);
xor U6993 (N_6993,N_5003,N_5099);
or U6994 (N_6994,N_5812,N_5386);
xnor U6995 (N_6995,N_5387,N_5800);
or U6996 (N_6996,N_5826,N_5142);
xor U6997 (N_6997,N_5379,N_5942);
and U6998 (N_6998,N_5441,N_5429);
and U6999 (N_6999,N_5937,N_5472);
nor U7000 (N_7000,N_6063,N_6195);
or U7001 (N_7001,N_6363,N_6813);
and U7002 (N_7002,N_6208,N_6588);
xor U7003 (N_7003,N_6962,N_6656);
or U7004 (N_7004,N_6372,N_6302);
or U7005 (N_7005,N_6470,N_6469);
and U7006 (N_7006,N_6895,N_6238);
nand U7007 (N_7007,N_6095,N_6938);
or U7008 (N_7008,N_6601,N_6537);
nand U7009 (N_7009,N_6915,N_6262);
xnor U7010 (N_7010,N_6657,N_6904);
xnor U7011 (N_7011,N_6531,N_6647);
or U7012 (N_7012,N_6825,N_6655);
or U7013 (N_7013,N_6663,N_6041);
and U7014 (N_7014,N_6031,N_6753);
nand U7015 (N_7015,N_6722,N_6923);
and U7016 (N_7016,N_6040,N_6506);
xnor U7017 (N_7017,N_6687,N_6336);
nor U7018 (N_7018,N_6475,N_6178);
xor U7019 (N_7019,N_6077,N_6089);
nand U7020 (N_7020,N_6815,N_6201);
xnor U7021 (N_7021,N_6673,N_6582);
and U7022 (N_7022,N_6439,N_6155);
nand U7023 (N_7023,N_6350,N_6256);
nand U7024 (N_7024,N_6411,N_6198);
and U7025 (N_7025,N_6203,N_6718);
and U7026 (N_7026,N_6886,N_6342);
and U7027 (N_7027,N_6274,N_6227);
and U7028 (N_7028,N_6567,N_6260);
nor U7029 (N_7029,N_6770,N_6480);
nor U7030 (N_7030,N_6574,N_6510);
nor U7031 (N_7031,N_6925,N_6635);
nor U7032 (N_7032,N_6829,N_6528);
nand U7033 (N_7033,N_6140,N_6586);
xnor U7034 (N_7034,N_6267,N_6228);
nor U7035 (N_7035,N_6045,N_6512);
nor U7036 (N_7036,N_6503,N_6892);
or U7037 (N_7037,N_6836,N_6787);
and U7038 (N_7038,N_6988,N_6028);
nand U7039 (N_7039,N_6812,N_6622);
or U7040 (N_7040,N_6278,N_6774);
or U7041 (N_7041,N_6175,N_6446);
xnor U7042 (N_7042,N_6630,N_6616);
xor U7043 (N_7043,N_6711,N_6735);
or U7044 (N_7044,N_6253,N_6550);
and U7045 (N_7045,N_6468,N_6569);
nor U7046 (N_7046,N_6896,N_6597);
nor U7047 (N_7047,N_6265,N_6857);
nor U7048 (N_7048,N_6998,N_6641);
nand U7049 (N_7049,N_6014,N_6897);
xor U7050 (N_7050,N_6951,N_6078);
nor U7051 (N_7051,N_6621,N_6946);
and U7052 (N_7052,N_6183,N_6057);
nor U7053 (N_7053,N_6778,N_6414);
or U7054 (N_7054,N_6375,N_6610);
nand U7055 (N_7055,N_6181,N_6147);
and U7056 (N_7056,N_6810,N_6392);
xor U7057 (N_7057,N_6868,N_6947);
or U7058 (N_7058,N_6488,N_6395);
or U7059 (N_7059,N_6076,N_6800);
xnor U7060 (N_7060,N_6455,N_6403);
or U7061 (N_7061,N_6313,N_6384);
xnor U7062 (N_7062,N_6235,N_6158);
and U7063 (N_7063,N_6995,N_6786);
xor U7064 (N_7064,N_6990,N_6294);
xor U7065 (N_7065,N_6715,N_6087);
xnor U7066 (N_7066,N_6276,N_6166);
nor U7067 (N_7067,N_6339,N_6481);
nor U7068 (N_7068,N_6308,N_6628);
xor U7069 (N_7069,N_6594,N_6590);
and U7070 (N_7070,N_6581,N_6879);
and U7071 (N_7071,N_6548,N_6913);
or U7072 (N_7072,N_6798,N_6280);
and U7073 (N_7073,N_6357,N_6871);
nor U7074 (N_7074,N_6324,N_6376);
xor U7075 (N_7075,N_6640,N_6981);
nand U7076 (N_7076,N_6092,N_6551);
xor U7077 (N_7077,N_6237,N_6501);
or U7078 (N_7078,N_6524,N_6286);
or U7079 (N_7079,N_6856,N_6434);
nor U7080 (N_7080,N_6606,N_6881);
nand U7081 (N_7081,N_6240,N_6568);
nor U7082 (N_7082,N_6114,N_6404);
and U7083 (N_7083,N_6373,N_6002);
nand U7084 (N_7084,N_6138,N_6213);
nand U7085 (N_7085,N_6499,N_6162);
nor U7086 (N_7086,N_6333,N_6710);
and U7087 (N_7087,N_6298,N_6843);
xor U7088 (N_7088,N_6393,N_6659);
nand U7089 (N_7089,N_6257,N_6607);
xor U7090 (N_7090,N_6254,N_6973);
and U7091 (N_7091,N_6697,N_6218);
xnor U7092 (N_7092,N_6458,N_6361);
and U7093 (N_7093,N_6232,N_6269);
nor U7094 (N_7094,N_6391,N_6413);
nor U7095 (N_7095,N_6565,N_6685);
or U7096 (N_7096,N_6771,N_6169);
or U7097 (N_7097,N_6937,N_6523);
or U7098 (N_7098,N_6609,N_6936);
nor U7099 (N_7099,N_6129,N_6943);
nand U7100 (N_7100,N_6241,N_6894);
nand U7101 (N_7101,N_6561,N_6136);
and U7102 (N_7102,N_6526,N_6865);
xor U7103 (N_7103,N_6194,N_6992);
xor U7104 (N_7104,N_6563,N_6553);
and U7105 (N_7105,N_6277,N_6049);
nor U7106 (N_7106,N_6126,N_6473);
xnor U7107 (N_7107,N_6354,N_6281);
nand U7108 (N_7108,N_6495,N_6975);
nand U7109 (N_7109,N_6017,N_6611);
or U7110 (N_7110,N_6584,N_6381);
or U7111 (N_7111,N_6182,N_6855);
and U7112 (N_7112,N_6750,N_6283);
and U7113 (N_7113,N_6364,N_6128);
xor U7114 (N_7114,N_6795,N_6156);
nand U7115 (N_7115,N_6779,N_6030);
and U7116 (N_7116,N_6793,N_6074);
and U7117 (N_7117,N_6084,N_6599);
xor U7118 (N_7118,N_6759,N_6461);
nor U7119 (N_7119,N_6081,N_6234);
nor U7120 (N_7120,N_6767,N_6820);
nand U7121 (N_7121,N_6848,N_6131);
or U7122 (N_7122,N_6487,N_6683);
or U7123 (N_7123,N_6852,N_6916);
nor U7124 (N_7124,N_6982,N_6742);
or U7125 (N_7125,N_6696,N_6775);
and U7126 (N_7126,N_6486,N_6766);
xnor U7127 (N_7127,N_6451,N_6681);
nand U7128 (N_7128,N_6080,N_6824);
nand U7129 (N_7129,N_6679,N_6427);
or U7130 (N_7130,N_6589,N_6070);
or U7131 (N_7131,N_6500,N_6006);
nor U7132 (N_7132,N_6456,N_6934);
or U7133 (N_7133,N_6629,N_6170);
nor U7134 (N_7134,N_6612,N_6782);
or U7135 (N_7135,N_6874,N_6728);
nor U7136 (N_7136,N_6119,N_6001);
or U7137 (N_7137,N_6559,N_6867);
nand U7138 (N_7138,N_6579,N_6387);
nor U7139 (N_7139,N_6890,N_6036);
and U7140 (N_7140,N_6008,N_6214);
nor U7141 (N_7141,N_6303,N_6618);
or U7142 (N_7142,N_6039,N_6514);
nor U7143 (N_7143,N_6408,N_6991);
nand U7144 (N_7144,N_6496,N_6004);
xnor U7145 (N_7145,N_6244,N_6910);
and U7146 (N_7146,N_6048,N_6519);
or U7147 (N_7147,N_6359,N_6167);
nand U7148 (N_7148,N_6211,N_6652);
nor U7149 (N_7149,N_6306,N_6318);
or U7150 (N_7150,N_6709,N_6191);
xnor U7151 (N_7151,N_6661,N_6570);
or U7152 (N_7152,N_6189,N_6250);
xnor U7153 (N_7153,N_6249,N_6365);
nor U7154 (N_7154,N_6963,N_6907);
or U7155 (N_7155,N_6018,N_6534);
xnor U7156 (N_7156,N_6533,N_6026);
and U7157 (N_7157,N_6111,N_6204);
nor U7158 (N_7158,N_6769,N_6580);
nand U7159 (N_7159,N_6419,N_6754);
or U7160 (N_7160,N_6639,N_6511);
xor U7161 (N_7161,N_6627,N_6719);
nor U7162 (N_7162,N_6329,N_6012);
and U7163 (N_7163,N_6987,N_6113);
xnor U7164 (N_7164,N_6341,N_6704);
and U7165 (N_7165,N_6478,N_6958);
nor U7166 (N_7166,N_6802,N_6840);
nor U7167 (N_7167,N_6816,N_6604);
xor U7168 (N_7168,N_6690,N_6513);
xor U7169 (N_7169,N_6634,N_6420);
xor U7170 (N_7170,N_6956,N_6423);
nor U7171 (N_7171,N_6142,N_6109);
xor U7172 (N_7172,N_6636,N_6864);
or U7173 (N_7173,N_6994,N_6110);
xor U7174 (N_7174,N_6643,N_6343);
and U7175 (N_7175,N_6424,N_6686);
nor U7176 (N_7176,N_6216,N_6858);
and U7177 (N_7177,N_6396,N_6493);
or U7178 (N_7178,N_6876,N_6530);
or U7179 (N_7179,N_6471,N_6974);
or U7180 (N_7180,N_6304,N_6436);
or U7181 (N_7181,N_6356,N_6190);
and U7182 (N_7182,N_6872,N_6841);
nor U7183 (N_7183,N_6970,N_6729);
and U7184 (N_7184,N_6781,N_6650);
or U7185 (N_7185,N_6337,N_6645);
nor U7186 (N_7186,N_6431,N_6023);
and U7187 (N_7187,N_6139,N_6877);
and U7188 (N_7188,N_6326,N_6052);
nand U7189 (N_7189,N_6355,N_6319);
nand U7190 (N_7190,N_6115,N_6527);
or U7191 (N_7191,N_6732,N_6462);
or U7192 (N_7192,N_6703,N_6112);
or U7193 (N_7193,N_6418,N_6300);
and U7194 (N_7194,N_6555,N_6159);
nand U7195 (N_7195,N_6442,N_6233);
or U7196 (N_7196,N_6021,N_6091);
or U7197 (N_7197,N_6993,N_6926);
and U7198 (N_7198,N_6849,N_6801);
nor U7199 (N_7199,N_6171,N_6971);
xor U7200 (N_7200,N_6747,N_6508);
nor U7201 (N_7201,N_6549,N_6046);
or U7202 (N_7202,N_6061,N_6415);
xnor U7203 (N_7203,N_6573,N_6425);
nor U7204 (N_7204,N_6058,N_6295);
nand U7205 (N_7205,N_6176,N_6056);
nand U7206 (N_7206,N_6430,N_6215);
nor U7207 (N_7207,N_6029,N_6906);
xnor U7208 (N_7208,N_6050,N_6094);
nor U7209 (N_7209,N_6741,N_6331);
nand U7210 (N_7210,N_6044,N_6505);
nand U7211 (N_7211,N_6490,N_6299);
nor U7212 (N_7212,N_6544,N_6389);
or U7213 (N_7213,N_6474,N_6831);
xor U7214 (N_7214,N_6422,N_6059);
xnor U7215 (N_7215,N_6323,N_6691);
and U7216 (N_7216,N_6726,N_6448);
nand U7217 (N_7217,N_6585,N_6309);
xor U7218 (N_7218,N_6417,N_6051);
nor U7219 (N_7219,N_6117,N_6082);
and U7220 (N_7220,N_6931,N_6121);
xor U7221 (N_7221,N_6577,N_6949);
and U7222 (N_7222,N_6399,N_6637);
nand U7223 (N_7223,N_6953,N_6477);
xnor U7224 (N_7224,N_6445,N_6273);
nand U7225 (N_7225,N_6416,N_6713);
and U7226 (N_7226,N_6187,N_6327);
or U7227 (N_7227,N_6217,N_6177);
or U7228 (N_7228,N_6509,N_6065);
and U7229 (N_7229,N_6792,N_6658);
nor U7230 (N_7230,N_6521,N_6349);
or U7231 (N_7231,N_6557,N_6385);
nor U7232 (N_7232,N_6624,N_6406);
xor U7233 (N_7233,N_6020,N_6055);
nor U7234 (N_7234,N_6866,N_6619);
nor U7235 (N_7235,N_6307,N_6435);
and U7236 (N_7236,N_6928,N_6933);
and U7237 (N_7237,N_6772,N_6572);
or U7238 (N_7238,N_6738,N_6598);
nand U7239 (N_7239,N_6914,N_6447);
and U7240 (N_7240,N_6251,N_6540);
nand U7241 (N_7241,N_6891,N_6246);
and U7242 (N_7242,N_6777,N_6097);
nor U7243 (N_7243,N_6737,N_6623);
xnor U7244 (N_7244,N_6067,N_6053);
or U7245 (N_7245,N_6522,N_6107);
nor U7246 (N_7246,N_6224,N_6518);
and U7247 (N_7247,N_6483,N_6702);
xnor U7248 (N_7248,N_6543,N_6003);
and U7249 (N_7249,N_6185,N_6912);
xor U7250 (N_7250,N_6733,N_6893);
or U7251 (N_7251,N_6672,N_6730);
or U7252 (N_7252,N_6721,N_6734);
nor U7253 (N_7253,N_6744,N_6748);
and U7254 (N_7254,N_6380,N_6444);
xnor U7255 (N_7255,N_6297,N_6438);
and U7256 (N_7256,N_6264,N_6498);
nor U7257 (N_7257,N_6132,N_6985);
or U7258 (N_7258,N_6908,N_6068);
or U7259 (N_7259,N_6714,N_6644);
nand U7260 (N_7260,N_6328,N_6860);
nand U7261 (N_7261,N_6016,N_6646);
nor U7262 (N_7262,N_6986,N_6861);
nand U7263 (N_7263,N_6976,N_6492);
and U7264 (N_7264,N_6862,N_6388);
and U7265 (N_7265,N_6806,N_6402);
nor U7266 (N_7266,N_6199,N_6207);
nand U7267 (N_7267,N_6037,N_6450);
or U7268 (N_7268,N_6072,N_6838);
and U7269 (N_7269,N_6999,N_6465);
nor U7270 (N_7270,N_6608,N_6948);
or U7271 (N_7271,N_6823,N_6371);
nor U7272 (N_7272,N_6547,N_6821);
or U7273 (N_7273,N_6157,N_6315);
xnor U7274 (N_7274,N_6071,N_6268);
nor U7275 (N_7275,N_6965,N_6614);
nor U7276 (N_7276,N_6684,N_6252);
or U7277 (N_7277,N_6977,N_6520);
nand U7278 (N_7278,N_6123,N_6751);
xnor U7279 (N_7279,N_6773,N_6620);
and U7280 (N_7280,N_6909,N_6311);
xor U7281 (N_7281,N_6542,N_6613);
or U7282 (N_7282,N_6209,N_6124);
or U7283 (N_7283,N_6366,N_6961);
nand U7284 (N_7284,N_6920,N_6151);
nor U7285 (N_7285,N_6803,N_6595);
xnor U7286 (N_7286,N_6847,N_6727);
xnor U7287 (N_7287,N_6900,N_6674);
or U7288 (N_7288,N_6134,N_6212);
nand U7289 (N_7289,N_6453,N_6869);
or U7290 (N_7290,N_6822,N_6790);
or U7291 (N_7291,N_6022,N_6287);
xor U7292 (N_7292,N_6193,N_6924);
and U7293 (N_7293,N_6541,N_6880);
and U7294 (N_7294,N_6103,N_6226);
nand U7295 (N_7295,N_6332,N_6148);
xnor U7296 (N_7296,N_6873,N_6762);
nor U7297 (N_7297,N_6064,N_6270);
and U7298 (N_7298,N_6675,N_6116);
xor U7299 (N_7299,N_6489,N_6069);
nor U7300 (N_7300,N_6504,N_6625);
and U7301 (N_7301,N_6789,N_6038);
or U7302 (N_7302,N_6693,N_6130);
xnor U7303 (N_7303,N_6811,N_6707);
xor U7304 (N_7304,N_6085,N_6688);
or U7305 (N_7305,N_6494,N_6818);
nand U7306 (N_7306,N_6255,N_6261);
and U7307 (N_7307,N_6168,N_6348);
or U7308 (N_7308,N_6780,N_6412);
xnor U7309 (N_7309,N_6667,N_6186);
nand U7310 (N_7310,N_6460,N_6596);
nand U7311 (N_7311,N_6804,N_6334);
and U7312 (N_7312,N_6027,N_6073);
and U7313 (N_7313,N_6671,N_6282);
or U7314 (N_7314,N_6141,N_6043);
or U7315 (N_7315,N_6996,N_6137);
and U7316 (N_7316,N_6854,N_6576);
nor U7317 (N_7317,N_6668,N_6593);
and U7318 (N_7318,N_6353,N_6377);
nand U7319 (N_7319,N_6653,N_6160);
nand U7320 (N_7320,N_6740,N_6791);
or U7321 (N_7321,N_6428,N_6788);
nand U7322 (N_7322,N_6409,N_6062);
and U7323 (N_7323,N_6086,N_6784);
and U7324 (N_7324,N_6013,N_6694);
or U7325 (N_7325,N_6516,N_6535);
xnor U7326 (N_7326,N_6497,N_6223);
or U7327 (N_7327,N_6150,N_6546);
xor U7328 (N_7328,N_6197,N_6670);
nand U7329 (N_7329,N_6314,N_6785);
or U7330 (N_7330,N_6720,N_6983);
nor U7331 (N_7331,N_6352,N_6905);
nand U7332 (N_7332,N_6827,N_6479);
or U7333 (N_7333,N_6903,N_6347);
or U7334 (N_7334,N_6154,N_6248);
or U7335 (N_7335,N_6292,N_6382);
and U7336 (N_7336,N_6545,N_6699);
and U7337 (N_7337,N_6410,N_6960);
nand U7338 (N_7338,N_6184,N_6033);
xor U7339 (N_7339,N_6401,N_6096);
nor U7340 (N_7340,N_6529,N_6370);
nand U7341 (N_7341,N_6809,N_6870);
or U7342 (N_7342,N_6745,N_6532);
nand U7343 (N_7343,N_6899,N_6457);
nand U7344 (N_7344,N_6919,N_6592);
nand U7345 (N_7345,N_6725,N_6664);
and U7346 (N_7346,N_6556,N_6321);
xor U7347 (N_7347,N_6941,N_6739);
and U7348 (N_7348,N_6901,N_6105);
and U7349 (N_7349,N_6144,N_6898);
nand U7350 (N_7350,N_6236,N_6942);
xor U7351 (N_7351,N_6221,N_6560);
or U7352 (N_7352,N_6290,N_6649);
nor U7353 (N_7353,N_6682,N_6379);
and U7354 (N_7354,N_6259,N_6472);
or U7355 (N_7355,N_6258,N_6485);
or U7356 (N_7356,N_6918,N_6717);
and U7357 (N_7357,N_6000,N_6152);
or U7358 (N_7358,N_6817,N_6954);
nand U7359 (N_7359,N_6997,N_6188);
nor U7360 (N_7360,N_6108,N_6397);
nand U7361 (N_7361,N_6638,N_6689);
nor U7362 (N_7362,N_6320,N_6692);
nand U7363 (N_7363,N_6239,N_6205);
or U7364 (N_7364,N_6174,N_6440);
and U7365 (N_7365,N_6764,N_6932);
xnor U7366 (N_7366,N_6398,N_6515);
nor U7367 (N_7367,N_6887,N_6957);
or U7368 (N_7368,N_6826,N_6626);
and U7369 (N_7369,N_6564,N_6575);
and U7370 (N_7370,N_6225,N_6940);
nor U7371 (N_7371,N_6875,N_6980);
or U7372 (N_7372,N_6676,N_6952);
nor U7373 (N_7373,N_6602,N_6301);
nand U7374 (N_7374,N_6369,N_6145);
xnor U7375 (N_7375,N_6210,N_6878);
or U7376 (N_7376,N_6093,N_6964);
nand U7377 (N_7377,N_6830,N_6677);
xor U7378 (N_7378,N_6378,N_6390);
xor U7379 (N_7379,N_6796,N_6367);
xnor U7380 (N_7380,N_6202,N_6405);
and U7381 (N_7381,N_6752,N_6133);
nor U7382 (N_7382,N_6010,N_6834);
xor U7383 (N_7383,N_6066,N_6749);
xor U7384 (N_7384,N_6322,N_6009);
and U7385 (N_7385,N_6288,N_6968);
and U7386 (N_7386,N_6959,N_6853);
nor U7387 (N_7387,N_6578,N_6426);
and U7388 (N_7388,N_6678,N_6192);
nor U7389 (N_7389,N_6945,N_6180);
xnor U7390 (N_7390,N_6007,N_6605);
and U7391 (N_7391,N_6716,N_6206);
xnor U7392 (N_7392,N_6955,N_6507);
and U7393 (N_7393,N_6746,N_6705);
or U7394 (N_7394,N_6024,N_6833);
and U7395 (N_7395,N_6648,N_6927);
nand U7396 (N_7396,N_6502,N_6344);
or U7397 (N_7397,N_6536,N_6034);
and U7398 (N_7398,N_6966,N_6911);
and U7399 (N_7399,N_6464,N_6433);
or U7400 (N_7400,N_6083,N_6368);
xnor U7401 (N_7401,N_6837,N_6374);
nand U7402 (N_7402,N_6229,N_6701);
or U7403 (N_7403,N_6079,N_6090);
nand U7404 (N_7404,N_6386,N_6902);
nor U7405 (N_7405,N_6122,N_6101);
and U7406 (N_7406,N_6617,N_6756);
nand U7407 (N_7407,N_6651,N_6432);
nand U7408 (N_7408,N_6296,N_6275);
or U7409 (N_7409,N_6757,N_6100);
or U7410 (N_7410,N_6102,N_6054);
nor U7411 (N_7411,N_6755,N_6763);
nor U7412 (N_7412,N_6761,N_6042);
nor U7413 (N_7413,N_6165,N_6466);
xnor U7414 (N_7414,N_6736,N_6317);
nor U7415 (N_7415,N_6340,N_6950);
xnor U7416 (N_7416,N_6346,N_6885);
and U7417 (N_7417,N_6441,N_6172);
nand U7418 (N_7418,N_6088,N_6120);
nand U7419 (N_7419,N_6768,N_6179);
nand U7420 (N_7420,N_6539,N_6247);
nor U7421 (N_7421,N_6305,N_6978);
and U7422 (N_7422,N_6285,N_6989);
xnor U7423 (N_7423,N_6452,N_6099);
nor U7424 (N_7424,N_6312,N_6149);
nor U7425 (N_7425,N_6325,N_6538);
nand U7426 (N_7426,N_6799,N_6743);
nor U7427 (N_7427,N_6633,N_6035);
or U7428 (N_7428,N_6525,N_6631);
xnor U7429 (N_7429,N_6272,N_6015);
or U7430 (N_7430,N_6330,N_6929);
or U7431 (N_7431,N_6723,N_6118);
and U7432 (N_7432,N_6846,N_6125);
nand U7433 (N_7433,N_6143,N_6163);
or U7434 (N_7434,N_6698,N_6459);
or U7435 (N_7435,N_6047,N_6844);
or U7436 (N_7436,N_6362,N_6922);
nand U7437 (N_7437,N_6394,N_6917);
nor U7438 (N_7438,N_6443,N_6695);
nand U7439 (N_7439,N_6266,N_6491);
nand U7440 (N_7440,N_6808,N_6984);
nor U7441 (N_7441,N_6562,N_6517);
or U7442 (N_7442,N_6807,N_6383);
nor U7443 (N_7443,N_6888,N_6127);
nand U7444 (N_7444,N_6429,N_6828);
xnor U7445 (N_7445,N_6712,N_6421);
or U7446 (N_7446,N_6760,N_6603);
and U7447 (N_7447,N_6284,N_6600);
or U7448 (N_7448,N_6245,N_6776);
nand U7449 (N_7449,N_6407,N_6583);
and U7450 (N_7450,N_6642,N_6935);
nor U7451 (N_7451,N_6164,N_6075);
nand U7452 (N_7452,N_6098,N_6289);
or U7453 (N_7453,N_6969,N_6231);
or U7454 (N_7454,N_6851,N_6338);
xnor U7455 (N_7455,N_6554,N_6591);
xnor U7456 (N_7456,N_6161,N_6484);
or U7457 (N_7457,N_6863,N_6883);
nor U7458 (N_7458,N_6351,N_6222);
nand U7459 (N_7459,N_6032,N_6930);
and U7460 (N_7460,N_6680,N_6797);
and U7461 (N_7461,N_6400,N_6967);
and U7462 (N_7462,N_6106,N_6850);
nand U7463 (N_7463,N_6454,N_6310);
xnor U7464 (N_7464,N_6814,N_6842);
nand U7465 (N_7465,N_6566,N_6263);
nand U7466 (N_7466,N_6884,N_6832);
and U7467 (N_7467,N_6291,N_6558);
nand U7468 (N_7468,N_6921,N_6662);
xnor U7469 (N_7469,N_6660,N_6845);
or U7470 (N_7470,N_6019,N_6316);
or U7471 (N_7471,N_6708,N_6449);
nor U7472 (N_7472,N_6242,N_6783);
or U7473 (N_7473,N_6345,N_6437);
xor U7474 (N_7474,N_6200,N_6665);
or U7475 (N_7475,N_6615,N_6173);
and U7476 (N_7476,N_6243,N_6104);
nand U7477 (N_7477,N_6654,N_6005);
nor U7478 (N_7478,N_6146,N_6135);
xor U7479 (N_7479,N_6025,N_6463);
nor U7480 (N_7480,N_6939,N_6360);
nor U7481 (N_7481,N_6972,N_6279);
xor U7482 (N_7482,N_6700,N_6060);
xor U7483 (N_7483,N_6724,N_6835);
nor U7484 (N_7484,N_6666,N_6358);
nand U7485 (N_7485,N_6230,N_6552);
nor U7486 (N_7486,N_6669,N_6476);
or U7487 (N_7487,N_6587,N_6882);
nor U7488 (N_7488,N_6196,N_6731);
xnor U7489 (N_7489,N_6011,N_6706);
nor U7490 (N_7490,N_6632,N_6482);
xnor U7491 (N_7491,N_6571,N_6467);
nor U7492 (N_7492,N_6839,N_6335);
and U7493 (N_7493,N_6219,N_6805);
nand U7494 (N_7494,N_6220,N_6794);
xor U7495 (N_7495,N_6153,N_6819);
nor U7496 (N_7496,N_6271,N_6889);
nor U7497 (N_7497,N_6859,N_6758);
xnor U7498 (N_7498,N_6979,N_6765);
nor U7499 (N_7499,N_6944,N_6293);
xor U7500 (N_7500,N_6088,N_6793);
nand U7501 (N_7501,N_6823,N_6391);
xor U7502 (N_7502,N_6443,N_6103);
xor U7503 (N_7503,N_6023,N_6840);
nor U7504 (N_7504,N_6865,N_6593);
or U7505 (N_7505,N_6831,N_6667);
nand U7506 (N_7506,N_6021,N_6191);
nand U7507 (N_7507,N_6704,N_6108);
nand U7508 (N_7508,N_6108,N_6637);
or U7509 (N_7509,N_6747,N_6724);
nand U7510 (N_7510,N_6552,N_6044);
nor U7511 (N_7511,N_6139,N_6595);
xor U7512 (N_7512,N_6821,N_6239);
nor U7513 (N_7513,N_6474,N_6367);
nor U7514 (N_7514,N_6517,N_6540);
xor U7515 (N_7515,N_6815,N_6110);
nand U7516 (N_7516,N_6914,N_6719);
xnor U7517 (N_7517,N_6780,N_6487);
nand U7518 (N_7518,N_6785,N_6882);
and U7519 (N_7519,N_6723,N_6036);
or U7520 (N_7520,N_6415,N_6050);
xor U7521 (N_7521,N_6591,N_6441);
nor U7522 (N_7522,N_6791,N_6739);
or U7523 (N_7523,N_6825,N_6907);
or U7524 (N_7524,N_6025,N_6039);
nor U7525 (N_7525,N_6034,N_6686);
or U7526 (N_7526,N_6380,N_6054);
nand U7527 (N_7527,N_6121,N_6656);
or U7528 (N_7528,N_6332,N_6135);
and U7529 (N_7529,N_6658,N_6463);
xnor U7530 (N_7530,N_6363,N_6021);
xor U7531 (N_7531,N_6592,N_6705);
xor U7532 (N_7532,N_6620,N_6489);
nor U7533 (N_7533,N_6830,N_6596);
nor U7534 (N_7534,N_6867,N_6619);
and U7535 (N_7535,N_6237,N_6392);
nand U7536 (N_7536,N_6619,N_6922);
nand U7537 (N_7537,N_6467,N_6805);
xnor U7538 (N_7538,N_6056,N_6520);
nor U7539 (N_7539,N_6215,N_6975);
xnor U7540 (N_7540,N_6182,N_6510);
nor U7541 (N_7541,N_6476,N_6633);
nand U7542 (N_7542,N_6037,N_6435);
xor U7543 (N_7543,N_6191,N_6076);
and U7544 (N_7544,N_6219,N_6767);
xor U7545 (N_7545,N_6899,N_6322);
nand U7546 (N_7546,N_6778,N_6108);
nand U7547 (N_7547,N_6248,N_6364);
and U7548 (N_7548,N_6388,N_6337);
and U7549 (N_7549,N_6552,N_6161);
nand U7550 (N_7550,N_6675,N_6303);
and U7551 (N_7551,N_6274,N_6942);
nand U7552 (N_7552,N_6835,N_6211);
and U7553 (N_7553,N_6267,N_6908);
or U7554 (N_7554,N_6423,N_6156);
or U7555 (N_7555,N_6182,N_6489);
nand U7556 (N_7556,N_6551,N_6807);
and U7557 (N_7557,N_6674,N_6039);
nand U7558 (N_7558,N_6741,N_6784);
or U7559 (N_7559,N_6275,N_6255);
nand U7560 (N_7560,N_6690,N_6571);
nor U7561 (N_7561,N_6859,N_6229);
nand U7562 (N_7562,N_6802,N_6866);
nor U7563 (N_7563,N_6464,N_6073);
or U7564 (N_7564,N_6143,N_6797);
or U7565 (N_7565,N_6169,N_6836);
or U7566 (N_7566,N_6543,N_6501);
nand U7567 (N_7567,N_6201,N_6795);
and U7568 (N_7568,N_6056,N_6884);
xnor U7569 (N_7569,N_6949,N_6026);
nor U7570 (N_7570,N_6586,N_6024);
nand U7571 (N_7571,N_6995,N_6157);
xnor U7572 (N_7572,N_6120,N_6312);
or U7573 (N_7573,N_6079,N_6626);
nand U7574 (N_7574,N_6698,N_6322);
nand U7575 (N_7575,N_6281,N_6777);
or U7576 (N_7576,N_6146,N_6789);
and U7577 (N_7577,N_6465,N_6218);
and U7578 (N_7578,N_6483,N_6942);
xnor U7579 (N_7579,N_6229,N_6255);
nor U7580 (N_7580,N_6061,N_6943);
xnor U7581 (N_7581,N_6163,N_6761);
or U7582 (N_7582,N_6090,N_6356);
or U7583 (N_7583,N_6475,N_6337);
or U7584 (N_7584,N_6734,N_6387);
nor U7585 (N_7585,N_6544,N_6999);
xor U7586 (N_7586,N_6636,N_6360);
xor U7587 (N_7587,N_6661,N_6874);
nor U7588 (N_7588,N_6423,N_6036);
nand U7589 (N_7589,N_6430,N_6103);
nand U7590 (N_7590,N_6468,N_6748);
nor U7591 (N_7591,N_6976,N_6422);
nor U7592 (N_7592,N_6087,N_6951);
nand U7593 (N_7593,N_6556,N_6417);
nor U7594 (N_7594,N_6041,N_6981);
xor U7595 (N_7595,N_6615,N_6792);
xnor U7596 (N_7596,N_6866,N_6272);
nand U7597 (N_7597,N_6034,N_6210);
nor U7598 (N_7598,N_6314,N_6866);
and U7599 (N_7599,N_6587,N_6438);
and U7600 (N_7600,N_6968,N_6785);
nor U7601 (N_7601,N_6564,N_6609);
and U7602 (N_7602,N_6013,N_6077);
or U7603 (N_7603,N_6342,N_6740);
and U7604 (N_7604,N_6466,N_6966);
or U7605 (N_7605,N_6335,N_6504);
or U7606 (N_7606,N_6606,N_6450);
xnor U7607 (N_7607,N_6752,N_6713);
nor U7608 (N_7608,N_6209,N_6550);
or U7609 (N_7609,N_6668,N_6874);
nand U7610 (N_7610,N_6768,N_6124);
and U7611 (N_7611,N_6993,N_6729);
xor U7612 (N_7612,N_6690,N_6793);
or U7613 (N_7613,N_6047,N_6060);
xnor U7614 (N_7614,N_6209,N_6580);
nand U7615 (N_7615,N_6331,N_6939);
or U7616 (N_7616,N_6725,N_6676);
nor U7617 (N_7617,N_6778,N_6291);
or U7618 (N_7618,N_6992,N_6957);
nor U7619 (N_7619,N_6101,N_6933);
or U7620 (N_7620,N_6283,N_6322);
nor U7621 (N_7621,N_6398,N_6452);
nor U7622 (N_7622,N_6109,N_6775);
nand U7623 (N_7623,N_6596,N_6638);
or U7624 (N_7624,N_6914,N_6403);
or U7625 (N_7625,N_6600,N_6614);
and U7626 (N_7626,N_6135,N_6742);
or U7627 (N_7627,N_6659,N_6143);
nand U7628 (N_7628,N_6425,N_6358);
and U7629 (N_7629,N_6449,N_6444);
or U7630 (N_7630,N_6335,N_6880);
or U7631 (N_7631,N_6663,N_6656);
nor U7632 (N_7632,N_6533,N_6170);
nor U7633 (N_7633,N_6734,N_6753);
nor U7634 (N_7634,N_6075,N_6796);
nand U7635 (N_7635,N_6738,N_6247);
nand U7636 (N_7636,N_6713,N_6860);
or U7637 (N_7637,N_6190,N_6084);
or U7638 (N_7638,N_6969,N_6476);
or U7639 (N_7639,N_6799,N_6068);
xnor U7640 (N_7640,N_6576,N_6521);
or U7641 (N_7641,N_6212,N_6417);
xnor U7642 (N_7642,N_6334,N_6972);
and U7643 (N_7643,N_6665,N_6947);
and U7644 (N_7644,N_6364,N_6760);
xor U7645 (N_7645,N_6010,N_6620);
and U7646 (N_7646,N_6220,N_6176);
nor U7647 (N_7647,N_6476,N_6948);
and U7648 (N_7648,N_6819,N_6649);
or U7649 (N_7649,N_6366,N_6923);
nor U7650 (N_7650,N_6837,N_6349);
xor U7651 (N_7651,N_6955,N_6797);
and U7652 (N_7652,N_6763,N_6483);
and U7653 (N_7653,N_6038,N_6568);
nor U7654 (N_7654,N_6499,N_6867);
nand U7655 (N_7655,N_6687,N_6255);
nand U7656 (N_7656,N_6066,N_6129);
nand U7657 (N_7657,N_6312,N_6574);
nand U7658 (N_7658,N_6690,N_6315);
and U7659 (N_7659,N_6968,N_6513);
xor U7660 (N_7660,N_6667,N_6878);
nor U7661 (N_7661,N_6537,N_6765);
and U7662 (N_7662,N_6700,N_6416);
and U7663 (N_7663,N_6019,N_6175);
or U7664 (N_7664,N_6274,N_6415);
or U7665 (N_7665,N_6356,N_6140);
nand U7666 (N_7666,N_6821,N_6173);
nor U7667 (N_7667,N_6824,N_6071);
nand U7668 (N_7668,N_6843,N_6861);
xnor U7669 (N_7669,N_6916,N_6895);
nor U7670 (N_7670,N_6948,N_6623);
and U7671 (N_7671,N_6894,N_6589);
and U7672 (N_7672,N_6552,N_6100);
nor U7673 (N_7673,N_6436,N_6229);
xor U7674 (N_7674,N_6380,N_6639);
xnor U7675 (N_7675,N_6572,N_6187);
xnor U7676 (N_7676,N_6677,N_6469);
nor U7677 (N_7677,N_6084,N_6311);
and U7678 (N_7678,N_6552,N_6857);
nor U7679 (N_7679,N_6835,N_6127);
and U7680 (N_7680,N_6711,N_6576);
nor U7681 (N_7681,N_6680,N_6757);
or U7682 (N_7682,N_6717,N_6888);
nor U7683 (N_7683,N_6607,N_6350);
or U7684 (N_7684,N_6063,N_6815);
xnor U7685 (N_7685,N_6708,N_6929);
xnor U7686 (N_7686,N_6632,N_6102);
xor U7687 (N_7687,N_6914,N_6550);
and U7688 (N_7688,N_6260,N_6592);
nor U7689 (N_7689,N_6246,N_6928);
or U7690 (N_7690,N_6496,N_6437);
nor U7691 (N_7691,N_6691,N_6139);
or U7692 (N_7692,N_6031,N_6745);
or U7693 (N_7693,N_6139,N_6028);
nor U7694 (N_7694,N_6442,N_6155);
and U7695 (N_7695,N_6616,N_6936);
or U7696 (N_7696,N_6996,N_6314);
or U7697 (N_7697,N_6511,N_6971);
nand U7698 (N_7698,N_6717,N_6015);
nor U7699 (N_7699,N_6601,N_6339);
xor U7700 (N_7700,N_6806,N_6457);
nand U7701 (N_7701,N_6841,N_6849);
and U7702 (N_7702,N_6588,N_6116);
nor U7703 (N_7703,N_6793,N_6591);
nand U7704 (N_7704,N_6386,N_6611);
and U7705 (N_7705,N_6866,N_6424);
nor U7706 (N_7706,N_6212,N_6286);
nand U7707 (N_7707,N_6266,N_6291);
nor U7708 (N_7708,N_6176,N_6609);
xnor U7709 (N_7709,N_6559,N_6307);
nand U7710 (N_7710,N_6761,N_6535);
xnor U7711 (N_7711,N_6753,N_6865);
nor U7712 (N_7712,N_6385,N_6087);
and U7713 (N_7713,N_6187,N_6616);
and U7714 (N_7714,N_6198,N_6483);
xor U7715 (N_7715,N_6213,N_6621);
nor U7716 (N_7716,N_6887,N_6006);
nand U7717 (N_7717,N_6737,N_6659);
nor U7718 (N_7718,N_6739,N_6081);
nand U7719 (N_7719,N_6371,N_6457);
nand U7720 (N_7720,N_6070,N_6376);
xor U7721 (N_7721,N_6443,N_6116);
and U7722 (N_7722,N_6529,N_6349);
nor U7723 (N_7723,N_6249,N_6386);
and U7724 (N_7724,N_6967,N_6845);
nor U7725 (N_7725,N_6548,N_6511);
nor U7726 (N_7726,N_6947,N_6719);
xor U7727 (N_7727,N_6812,N_6379);
nand U7728 (N_7728,N_6510,N_6220);
nand U7729 (N_7729,N_6292,N_6704);
or U7730 (N_7730,N_6701,N_6466);
nor U7731 (N_7731,N_6501,N_6037);
nand U7732 (N_7732,N_6376,N_6789);
nand U7733 (N_7733,N_6295,N_6620);
and U7734 (N_7734,N_6312,N_6964);
xnor U7735 (N_7735,N_6938,N_6975);
or U7736 (N_7736,N_6476,N_6327);
and U7737 (N_7737,N_6734,N_6761);
and U7738 (N_7738,N_6168,N_6889);
xnor U7739 (N_7739,N_6460,N_6217);
xnor U7740 (N_7740,N_6893,N_6209);
nor U7741 (N_7741,N_6595,N_6601);
or U7742 (N_7742,N_6963,N_6645);
xor U7743 (N_7743,N_6650,N_6290);
nand U7744 (N_7744,N_6012,N_6979);
or U7745 (N_7745,N_6652,N_6866);
nor U7746 (N_7746,N_6086,N_6581);
or U7747 (N_7747,N_6878,N_6068);
xnor U7748 (N_7748,N_6001,N_6002);
nor U7749 (N_7749,N_6362,N_6515);
and U7750 (N_7750,N_6500,N_6861);
xor U7751 (N_7751,N_6002,N_6149);
and U7752 (N_7752,N_6429,N_6932);
xor U7753 (N_7753,N_6640,N_6786);
or U7754 (N_7754,N_6525,N_6013);
nand U7755 (N_7755,N_6625,N_6896);
xor U7756 (N_7756,N_6419,N_6606);
nand U7757 (N_7757,N_6607,N_6094);
nand U7758 (N_7758,N_6358,N_6294);
xnor U7759 (N_7759,N_6845,N_6592);
and U7760 (N_7760,N_6088,N_6894);
nand U7761 (N_7761,N_6435,N_6369);
and U7762 (N_7762,N_6399,N_6295);
nand U7763 (N_7763,N_6228,N_6080);
or U7764 (N_7764,N_6811,N_6788);
nand U7765 (N_7765,N_6618,N_6278);
and U7766 (N_7766,N_6656,N_6088);
and U7767 (N_7767,N_6689,N_6827);
and U7768 (N_7768,N_6010,N_6830);
nor U7769 (N_7769,N_6972,N_6965);
and U7770 (N_7770,N_6051,N_6238);
nor U7771 (N_7771,N_6944,N_6223);
or U7772 (N_7772,N_6519,N_6643);
or U7773 (N_7773,N_6325,N_6843);
or U7774 (N_7774,N_6715,N_6130);
xnor U7775 (N_7775,N_6510,N_6897);
and U7776 (N_7776,N_6783,N_6326);
and U7777 (N_7777,N_6718,N_6863);
and U7778 (N_7778,N_6672,N_6237);
nor U7779 (N_7779,N_6293,N_6010);
xor U7780 (N_7780,N_6528,N_6474);
xnor U7781 (N_7781,N_6190,N_6536);
nor U7782 (N_7782,N_6597,N_6288);
nor U7783 (N_7783,N_6745,N_6215);
nand U7784 (N_7784,N_6116,N_6359);
xnor U7785 (N_7785,N_6788,N_6786);
xor U7786 (N_7786,N_6407,N_6728);
or U7787 (N_7787,N_6703,N_6290);
nor U7788 (N_7788,N_6321,N_6562);
xor U7789 (N_7789,N_6304,N_6038);
and U7790 (N_7790,N_6431,N_6689);
nor U7791 (N_7791,N_6135,N_6075);
or U7792 (N_7792,N_6082,N_6496);
nand U7793 (N_7793,N_6099,N_6262);
xor U7794 (N_7794,N_6480,N_6866);
nor U7795 (N_7795,N_6018,N_6779);
xnor U7796 (N_7796,N_6734,N_6670);
and U7797 (N_7797,N_6191,N_6620);
nor U7798 (N_7798,N_6166,N_6698);
nor U7799 (N_7799,N_6557,N_6246);
nand U7800 (N_7800,N_6899,N_6394);
xnor U7801 (N_7801,N_6954,N_6627);
nor U7802 (N_7802,N_6382,N_6013);
xnor U7803 (N_7803,N_6763,N_6730);
or U7804 (N_7804,N_6912,N_6285);
and U7805 (N_7805,N_6535,N_6252);
or U7806 (N_7806,N_6205,N_6121);
or U7807 (N_7807,N_6682,N_6070);
and U7808 (N_7808,N_6149,N_6256);
and U7809 (N_7809,N_6112,N_6977);
nor U7810 (N_7810,N_6113,N_6824);
or U7811 (N_7811,N_6440,N_6725);
nand U7812 (N_7812,N_6655,N_6007);
nand U7813 (N_7813,N_6882,N_6503);
nor U7814 (N_7814,N_6768,N_6573);
or U7815 (N_7815,N_6140,N_6060);
and U7816 (N_7816,N_6893,N_6088);
nor U7817 (N_7817,N_6747,N_6395);
or U7818 (N_7818,N_6365,N_6876);
nor U7819 (N_7819,N_6201,N_6092);
nor U7820 (N_7820,N_6957,N_6165);
nand U7821 (N_7821,N_6457,N_6262);
nand U7822 (N_7822,N_6823,N_6038);
xor U7823 (N_7823,N_6042,N_6030);
xnor U7824 (N_7824,N_6146,N_6624);
or U7825 (N_7825,N_6662,N_6655);
or U7826 (N_7826,N_6495,N_6617);
nand U7827 (N_7827,N_6715,N_6871);
xnor U7828 (N_7828,N_6953,N_6908);
nor U7829 (N_7829,N_6553,N_6033);
nand U7830 (N_7830,N_6608,N_6056);
nand U7831 (N_7831,N_6680,N_6238);
nor U7832 (N_7832,N_6120,N_6668);
nand U7833 (N_7833,N_6881,N_6946);
and U7834 (N_7834,N_6623,N_6272);
nor U7835 (N_7835,N_6094,N_6587);
xnor U7836 (N_7836,N_6219,N_6778);
nor U7837 (N_7837,N_6656,N_6393);
xor U7838 (N_7838,N_6471,N_6285);
nand U7839 (N_7839,N_6235,N_6714);
nor U7840 (N_7840,N_6044,N_6416);
or U7841 (N_7841,N_6873,N_6280);
xor U7842 (N_7842,N_6608,N_6048);
and U7843 (N_7843,N_6539,N_6189);
nor U7844 (N_7844,N_6217,N_6445);
or U7845 (N_7845,N_6863,N_6346);
nor U7846 (N_7846,N_6058,N_6976);
nand U7847 (N_7847,N_6303,N_6502);
xor U7848 (N_7848,N_6122,N_6900);
nand U7849 (N_7849,N_6710,N_6216);
nand U7850 (N_7850,N_6545,N_6626);
or U7851 (N_7851,N_6644,N_6400);
and U7852 (N_7852,N_6190,N_6573);
xnor U7853 (N_7853,N_6132,N_6476);
and U7854 (N_7854,N_6063,N_6277);
xor U7855 (N_7855,N_6593,N_6523);
xor U7856 (N_7856,N_6352,N_6099);
or U7857 (N_7857,N_6921,N_6055);
nor U7858 (N_7858,N_6643,N_6627);
nand U7859 (N_7859,N_6252,N_6514);
xor U7860 (N_7860,N_6554,N_6828);
and U7861 (N_7861,N_6932,N_6292);
nand U7862 (N_7862,N_6258,N_6775);
nand U7863 (N_7863,N_6037,N_6279);
nand U7864 (N_7864,N_6198,N_6643);
xnor U7865 (N_7865,N_6041,N_6050);
or U7866 (N_7866,N_6854,N_6728);
and U7867 (N_7867,N_6915,N_6870);
or U7868 (N_7868,N_6178,N_6680);
nand U7869 (N_7869,N_6757,N_6838);
nand U7870 (N_7870,N_6386,N_6861);
nor U7871 (N_7871,N_6801,N_6308);
or U7872 (N_7872,N_6300,N_6677);
or U7873 (N_7873,N_6167,N_6255);
or U7874 (N_7874,N_6991,N_6329);
xnor U7875 (N_7875,N_6794,N_6847);
or U7876 (N_7876,N_6285,N_6520);
and U7877 (N_7877,N_6748,N_6199);
nand U7878 (N_7878,N_6848,N_6044);
and U7879 (N_7879,N_6407,N_6841);
nand U7880 (N_7880,N_6747,N_6340);
or U7881 (N_7881,N_6190,N_6575);
xnor U7882 (N_7882,N_6307,N_6076);
xor U7883 (N_7883,N_6808,N_6188);
and U7884 (N_7884,N_6797,N_6840);
xor U7885 (N_7885,N_6279,N_6903);
nand U7886 (N_7886,N_6747,N_6153);
or U7887 (N_7887,N_6790,N_6910);
or U7888 (N_7888,N_6985,N_6678);
nor U7889 (N_7889,N_6479,N_6484);
or U7890 (N_7890,N_6009,N_6204);
or U7891 (N_7891,N_6103,N_6980);
nor U7892 (N_7892,N_6833,N_6318);
xnor U7893 (N_7893,N_6451,N_6033);
nor U7894 (N_7894,N_6273,N_6766);
nor U7895 (N_7895,N_6312,N_6048);
or U7896 (N_7896,N_6934,N_6938);
xnor U7897 (N_7897,N_6613,N_6747);
or U7898 (N_7898,N_6084,N_6544);
or U7899 (N_7899,N_6406,N_6701);
xnor U7900 (N_7900,N_6594,N_6245);
xor U7901 (N_7901,N_6846,N_6669);
nand U7902 (N_7902,N_6118,N_6340);
and U7903 (N_7903,N_6921,N_6146);
nand U7904 (N_7904,N_6636,N_6790);
nor U7905 (N_7905,N_6120,N_6950);
nand U7906 (N_7906,N_6223,N_6762);
or U7907 (N_7907,N_6263,N_6389);
nand U7908 (N_7908,N_6653,N_6619);
nand U7909 (N_7909,N_6737,N_6608);
nand U7910 (N_7910,N_6184,N_6738);
xor U7911 (N_7911,N_6704,N_6701);
or U7912 (N_7912,N_6703,N_6103);
and U7913 (N_7913,N_6718,N_6656);
nand U7914 (N_7914,N_6055,N_6818);
nand U7915 (N_7915,N_6604,N_6793);
nor U7916 (N_7916,N_6030,N_6080);
nand U7917 (N_7917,N_6060,N_6902);
or U7918 (N_7918,N_6626,N_6426);
nor U7919 (N_7919,N_6111,N_6229);
nor U7920 (N_7920,N_6048,N_6907);
nand U7921 (N_7921,N_6231,N_6025);
nand U7922 (N_7922,N_6571,N_6168);
and U7923 (N_7923,N_6542,N_6578);
nand U7924 (N_7924,N_6166,N_6011);
and U7925 (N_7925,N_6254,N_6491);
nand U7926 (N_7926,N_6687,N_6744);
nand U7927 (N_7927,N_6956,N_6374);
and U7928 (N_7928,N_6122,N_6185);
nor U7929 (N_7929,N_6965,N_6735);
xnor U7930 (N_7930,N_6428,N_6638);
nand U7931 (N_7931,N_6380,N_6227);
nor U7932 (N_7932,N_6983,N_6595);
nor U7933 (N_7933,N_6699,N_6202);
and U7934 (N_7934,N_6372,N_6191);
or U7935 (N_7935,N_6135,N_6940);
nor U7936 (N_7936,N_6900,N_6785);
nand U7937 (N_7937,N_6021,N_6259);
xor U7938 (N_7938,N_6970,N_6480);
nor U7939 (N_7939,N_6751,N_6042);
or U7940 (N_7940,N_6100,N_6429);
xnor U7941 (N_7941,N_6310,N_6234);
nand U7942 (N_7942,N_6526,N_6772);
xor U7943 (N_7943,N_6672,N_6155);
nand U7944 (N_7944,N_6409,N_6859);
xor U7945 (N_7945,N_6713,N_6553);
nand U7946 (N_7946,N_6438,N_6704);
and U7947 (N_7947,N_6309,N_6426);
nand U7948 (N_7948,N_6123,N_6537);
or U7949 (N_7949,N_6197,N_6530);
or U7950 (N_7950,N_6833,N_6411);
nand U7951 (N_7951,N_6414,N_6080);
nor U7952 (N_7952,N_6552,N_6070);
and U7953 (N_7953,N_6726,N_6441);
and U7954 (N_7954,N_6686,N_6299);
and U7955 (N_7955,N_6594,N_6191);
and U7956 (N_7956,N_6588,N_6883);
or U7957 (N_7957,N_6196,N_6458);
nand U7958 (N_7958,N_6070,N_6403);
and U7959 (N_7959,N_6933,N_6302);
or U7960 (N_7960,N_6703,N_6794);
xnor U7961 (N_7961,N_6521,N_6331);
xor U7962 (N_7962,N_6230,N_6033);
nor U7963 (N_7963,N_6284,N_6571);
nor U7964 (N_7964,N_6368,N_6762);
or U7965 (N_7965,N_6532,N_6383);
or U7966 (N_7966,N_6129,N_6034);
xnor U7967 (N_7967,N_6868,N_6790);
nand U7968 (N_7968,N_6161,N_6685);
xnor U7969 (N_7969,N_6520,N_6001);
and U7970 (N_7970,N_6776,N_6174);
and U7971 (N_7971,N_6926,N_6247);
or U7972 (N_7972,N_6721,N_6538);
and U7973 (N_7973,N_6882,N_6429);
nor U7974 (N_7974,N_6317,N_6250);
nor U7975 (N_7975,N_6234,N_6110);
nand U7976 (N_7976,N_6697,N_6839);
nor U7977 (N_7977,N_6586,N_6806);
nor U7978 (N_7978,N_6783,N_6683);
and U7979 (N_7979,N_6925,N_6234);
nor U7980 (N_7980,N_6987,N_6641);
xor U7981 (N_7981,N_6845,N_6516);
nor U7982 (N_7982,N_6769,N_6812);
or U7983 (N_7983,N_6849,N_6912);
nor U7984 (N_7984,N_6881,N_6634);
or U7985 (N_7985,N_6719,N_6310);
xor U7986 (N_7986,N_6372,N_6255);
and U7987 (N_7987,N_6603,N_6662);
and U7988 (N_7988,N_6021,N_6721);
and U7989 (N_7989,N_6933,N_6766);
xnor U7990 (N_7990,N_6223,N_6697);
xnor U7991 (N_7991,N_6125,N_6146);
and U7992 (N_7992,N_6017,N_6740);
xnor U7993 (N_7993,N_6876,N_6721);
or U7994 (N_7994,N_6188,N_6468);
and U7995 (N_7995,N_6277,N_6478);
or U7996 (N_7996,N_6291,N_6195);
or U7997 (N_7997,N_6436,N_6163);
and U7998 (N_7998,N_6470,N_6274);
or U7999 (N_7999,N_6030,N_6871);
or U8000 (N_8000,N_7726,N_7085);
or U8001 (N_8001,N_7820,N_7801);
nor U8002 (N_8002,N_7523,N_7078);
nand U8003 (N_8003,N_7843,N_7217);
and U8004 (N_8004,N_7895,N_7572);
and U8005 (N_8005,N_7839,N_7877);
nor U8006 (N_8006,N_7677,N_7267);
and U8007 (N_8007,N_7077,N_7794);
or U8008 (N_8008,N_7351,N_7832);
nand U8009 (N_8009,N_7674,N_7384);
xor U8010 (N_8010,N_7395,N_7744);
nor U8011 (N_8011,N_7380,N_7630);
xnor U8012 (N_8012,N_7368,N_7706);
nor U8013 (N_8013,N_7927,N_7885);
nand U8014 (N_8014,N_7062,N_7902);
or U8015 (N_8015,N_7250,N_7819);
or U8016 (N_8016,N_7005,N_7458);
and U8017 (N_8017,N_7957,N_7886);
and U8018 (N_8018,N_7404,N_7101);
or U8019 (N_8019,N_7683,N_7029);
nor U8020 (N_8020,N_7076,N_7386);
or U8021 (N_8021,N_7610,N_7342);
and U8022 (N_8022,N_7598,N_7130);
or U8023 (N_8023,N_7714,N_7031);
xnor U8024 (N_8024,N_7498,N_7797);
and U8025 (N_8025,N_7387,N_7583);
xor U8026 (N_8026,N_7012,N_7139);
nand U8027 (N_8027,N_7441,N_7360);
nor U8028 (N_8028,N_7204,N_7298);
nor U8029 (N_8029,N_7481,N_7708);
xor U8030 (N_8030,N_7492,N_7923);
and U8031 (N_8031,N_7858,N_7881);
or U8032 (N_8032,N_7716,N_7975);
xor U8033 (N_8033,N_7277,N_7397);
nand U8034 (N_8034,N_7324,N_7475);
nand U8035 (N_8035,N_7179,N_7039);
or U8036 (N_8036,N_7308,N_7450);
and U8037 (N_8037,N_7034,N_7753);
nand U8038 (N_8038,N_7868,N_7695);
or U8039 (N_8039,N_7383,N_7017);
xor U8040 (N_8040,N_7268,N_7741);
and U8041 (N_8041,N_7999,N_7749);
and U8042 (N_8042,N_7206,N_7325);
and U8043 (N_8043,N_7149,N_7912);
xnor U8044 (N_8044,N_7331,N_7917);
nand U8045 (N_8045,N_7542,N_7200);
and U8046 (N_8046,N_7611,N_7157);
nor U8047 (N_8047,N_7913,N_7785);
and U8048 (N_8048,N_7246,N_7056);
nand U8049 (N_8049,N_7619,N_7265);
or U8050 (N_8050,N_7191,N_7466);
nand U8051 (N_8051,N_7903,N_7549);
nor U8052 (N_8052,N_7335,N_7847);
or U8053 (N_8053,N_7873,N_7033);
or U8054 (N_8054,N_7750,N_7929);
and U8055 (N_8055,N_7815,N_7291);
nand U8056 (N_8056,N_7586,N_7676);
or U8057 (N_8057,N_7374,N_7208);
or U8058 (N_8058,N_7399,N_7125);
nand U8059 (N_8059,N_7252,N_7192);
nor U8060 (N_8060,N_7436,N_7216);
nand U8061 (N_8061,N_7552,N_7494);
nand U8062 (N_8062,N_7457,N_7071);
xor U8063 (N_8063,N_7168,N_7569);
or U8064 (N_8064,N_7953,N_7963);
nor U8065 (N_8065,N_7045,N_7535);
or U8066 (N_8066,N_7231,N_7269);
nor U8067 (N_8067,N_7348,N_7205);
nand U8068 (N_8068,N_7508,N_7057);
or U8069 (N_8069,N_7640,N_7911);
xnor U8070 (N_8070,N_7106,N_7745);
nor U8071 (N_8071,N_7233,N_7339);
xnor U8072 (N_8072,N_7122,N_7852);
and U8073 (N_8073,N_7987,N_7218);
and U8074 (N_8074,N_7402,N_7748);
nor U8075 (N_8075,N_7701,N_7067);
nand U8076 (N_8076,N_7789,N_7996);
nor U8077 (N_8077,N_7560,N_7124);
xnor U8078 (N_8078,N_7937,N_7771);
and U8079 (N_8079,N_7792,N_7530);
nand U8080 (N_8080,N_7228,N_7439);
nand U8081 (N_8081,N_7018,N_7720);
nor U8082 (N_8082,N_7734,N_7696);
or U8083 (N_8083,N_7440,N_7155);
nand U8084 (N_8084,N_7871,N_7609);
xnor U8085 (N_8085,N_7964,N_7471);
xor U8086 (N_8086,N_7737,N_7555);
nor U8087 (N_8087,N_7952,N_7775);
xor U8088 (N_8088,N_7697,N_7392);
xnor U8089 (N_8089,N_7958,N_7703);
and U8090 (N_8090,N_7922,N_7317);
xnor U8091 (N_8091,N_7562,N_7137);
xor U8092 (N_8092,N_7866,N_7756);
xor U8093 (N_8093,N_7517,N_7261);
xor U8094 (N_8094,N_7694,N_7491);
nor U8095 (N_8095,N_7988,N_7768);
xor U8096 (N_8096,N_7730,N_7140);
or U8097 (N_8097,N_7110,N_7008);
nand U8098 (N_8098,N_7307,N_7480);
and U8099 (N_8099,N_7512,N_7593);
nand U8100 (N_8100,N_7333,N_7415);
xor U8101 (N_8101,N_7486,N_7002);
and U8102 (N_8102,N_7181,N_7025);
nor U8103 (N_8103,N_7459,N_7582);
or U8104 (N_8104,N_7263,N_7778);
xnor U8105 (N_8105,N_7490,N_7617);
nor U8106 (N_8106,N_7303,N_7295);
or U8107 (N_8107,N_7310,N_7717);
and U8108 (N_8108,N_7722,N_7275);
nor U8109 (N_8109,N_7976,N_7270);
xor U8110 (N_8110,N_7563,N_7770);
nor U8111 (N_8111,N_7152,N_7190);
and U8112 (N_8112,N_7294,N_7534);
or U8113 (N_8113,N_7069,N_7980);
nor U8114 (N_8114,N_7243,N_7575);
nand U8115 (N_8115,N_7763,N_7272);
xor U8116 (N_8116,N_7848,N_7973);
or U8117 (N_8117,N_7812,N_7669);
xor U8118 (N_8118,N_7513,N_7121);
nor U8119 (N_8119,N_7428,N_7639);
or U8120 (N_8120,N_7514,N_7213);
nand U8121 (N_8121,N_7764,N_7391);
nor U8122 (N_8122,N_7736,N_7478);
and U8123 (N_8123,N_7707,N_7482);
xor U8124 (N_8124,N_7581,N_7890);
or U8125 (N_8125,N_7189,N_7460);
or U8126 (N_8126,N_7648,N_7553);
xnor U8127 (N_8127,N_7548,N_7100);
and U8128 (N_8128,N_7974,N_7787);
nand U8129 (N_8129,N_7188,N_7223);
nand U8130 (N_8130,N_7052,N_7529);
xnor U8131 (N_8131,N_7398,N_7063);
xor U8132 (N_8132,N_7524,N_7762);
xnor U8133 (N_8133,N_7343,N_7961);
or U8134 (N_8134,N_7808,N_7431);
xor U8135 (N_8135,N_7306,N_7526);
nor U8136 (N_8136,N_7334,N_7813);
or U8137 (N_8137,N_7326,N_7350);
nand U8138 (N_8138,N_7951,N_7729);
nor U8139 (N_8139,N_7418,N_7144);
or U8140 (N_8140,N_7414,N_7662);
and U8141 (N_8141,N_7977,N_7625);
and U8142 (N_8142,N_7919,N_7219);
xnor U8143 (N_8143,N_7477,N_7599);
nand U8144 (N_8144,N_7081,N_7469);
xnor U8145 (N_8145,N_7665,N_7914);
or U8146 (N_8146,N_7153,N_7358);
nor U8147 (N_8147,N_7255,N_7165);
and U8148 (N_8148,N_7821,N_7557);
and U8149 (N_8149,N_7993,N_7313);
nor U8150 (N_8150,N_7184,N_7282);
or U8151 (N_8151,N_7273,N_7158);
nand U8152 (N_8152,N_7401,N_7271);
nor U8153 (N_8153,N_7288,N_7518);
xnor U8154 (N_8154,N_7758,N_7869);
and U8155 (N_8155,N_7680,N_7826);
xnor U8156 (N_8156,N_7042,N_7875);
nand U8157 (N_8157,N_7073,N_7783);
and U8158 (N_8158,N_7891,N_7698);
xor U8159 (N_8159,N_7989,N_7286);
xor U8160 (N_8160,N_7765,N_7114);
and U8161 (N_8161,N_7969,N_7613);
xor U8162 (N_8162,N_7962,N_7527);
xnor U8163 (N_8163,N_7520,N_7661);
and U8164 (N_8164,N_7882,N_7585);
and U8165 (N_8165,N_7925,N_7878);
nand U8166 (N_8166,N_7773,N_7405);
nor U8167 (N_8167,N_7488,N_7690);
or U8168 (N_8168,N_7984,N_7107);
nor U8169 (N_8169,N_7222,N_7315);
and U8170 (N_8170,N_7788,N_7910);
xor U8171 (N_8171,N_7811,N_7187);
and U8172 (N_8172,N_7502,N_7510);
nand U8173 (N_8173,N_7171,N_7851);
or U8174 (N_8174,N_7452,N_7242);
and U8175 (N_8175,N_7629,N_7983);
and U8176 (N_8176,N_7994,N_7944);
and U8177 (N_8177,N_7943,N_7833);
nand U8178 (N_8178,N_7175,N_7506);
and U8179 (N_8179,N_7934,N_7505);
or U8180 (N_8180,N_7151,N_7389);
and U8181 (N_8181,N_7332,N_7058);
xnor U8182 (N_8182,N_7115,N_7390);
nand U8183 (N_8183,N_7864,N_7026);
nor U8184 (N_8184,N_7899,N_7237);
nand U8185 (N_8185,N_7090,N_7007);
and U8186 (N_8186,N_7825,N_7793);
or U8187 (N_8187,N_7670,N_7373);
nand U8188 (N_8188,N_7096,N_7254);
and U8189 (N_8189,N_7860,N_7127);
nor U8190 (N_8190,N_7713,N_7900);
and U8191 (N_8191,N_7060,N_7564);
xor U8192 (N_8192,N_7176,N_7435);
xnor U8193 (N_8193,N_7461,N_7699);
xnor U8194 (N_8194,N_7644,N_7330);
and U8195 (N_8195,N_7495,N_7221);
nor U8196 (N_8196,N_7889,N_7940);
nor U8197 (N_8197,N_7658,N_7309);
nor U8198 (N_8198,N_7497,N_7499);
xor U8199 (N_8199,N_7632,N_7606);
xor U8200 (N_8200,N_7588,N_7232);
and U8201 (N_8201,N_7182,N_7620);
nor U8202 (N_8202,N_7378,N_7388);
xnor U8203 (N_8203,N_7604,N_7827);
or U8204 (N_8204,N_7584,N_7337);
or U8205 (N_8205,N_7064,N_7627);
and U8206 (N_8206,N_7509,N_7098);
nor U8207 (N_8207,N_7016,N_7183);
xor U8208 (N_8208,N_7382,N_7995);
nand U8209 (N_8209,N_7249,N_7049);
nand U8210 (N_8210,N_7769,N_7830);
xor U8211 (N_8211,N_7936,N_7394);
nor U8212 (N_8212,N_7804,N_7372);
nand U8213 (N_8213,N_7280,N_7111);
and U8214 (N_8214,N_7960,N_7215);
nand U8215 (N_8215,N_7809,N_7614);
or U8216 (N_8216,N_7352,N_7199);
or U8217 (N_8217,N_7577,N_7766);
xor U8218 (N_8218,N_7319,N_7074);
nand U8219 (N_8219,N_7318,N_7659);
nand U8220 (N_8220,N_7321,N_7455);
nor U8221 (N_8221,N_7412,N_7657);
nand U8222 (N_8222,N_7207,N_7301);
or U8223 (N_8223,N_7863,N_7979);
nor U8224 (N_8224,N_7915,N_7304);
xor U8225 (N_8225,N_7939,N_7533);
or U8226 (N_8226,N_7180,N_7230);
and U8227 (N_8227,N_7022,N_7251);
and U8228 (N_8228,N_7791,N_7129);
and U8229 (N_8229,N_7814,N_7733);
and U8230 (N_8230,N_7992,N_7592);
or U8231 (N_8231,N_7278,N_7143);
xor U8232 (N_8232,N_7705,N_7366);
nor U8233 (N_8233,N_7501,N_7244);
xor U8234 (N_8234,N_7772,N_7986);
nor U8235 (N_8235,N_7311,N_7550);
nor U8236 (N_8236,N_7369,N_7041);
and U8237 (N_8237,N_7340,N_7551);
nand U8238 (N_8238,N_7715,N_7879);
nand U8239 (N_8239,N_7693,N_7567);
nor U8240 (N_8240,N_7872,N_7160);
nand U8241 (N_8241,N_7645,N_7924);
nand U8242 (N_8242,N_7603,N_7123);
nor U8243 (N_8243,N_7897,N_7195);
xnor U8244 (N_8244,N_7021,N_7220);
nor U8245 (N_8245,N_7921,N_7624);
nor U8246 (N_8246,N_7673,N_7036);
and U8247 (N_8247,N_7245,N_7709);
nand U8248 (N_8248,N_7214,N_7344);
or U8249 (N_8249,N_7449,N_7009);
xnor U8250 (N_8250,N_7774,N_7982);
nor U8251 (N_8251,N_7971,N_7818);
nand U8252 (N_8252,N_7167,N_7883);
and U8253 (N_8253,N_7253,N_7561);
nor U8254 (N_8254,N_7727,N_7210);
nor U8255 (N_8255,N_7105,N_7884);
or U8256 (N_8256,N_7568,N_7238);
nand U8257 (N_8257,N_7044,N_7487);
and U8258 (N_8258,N_7597,N_7136);
nor U8259 (N_8259,N_7692,N_7430);
xnor U8260 (N_8260,N_7972,N_7462);
and U8261 (N_8261,N_7299,N_7032);
xnor U8262 (N_8262,N_7359,N_7615);
xor U8263 (N_8263,N_7867,N_7393);
nand U8264 (N_8264,N_7746,N_7362);
and U8265 (N_8265,N_7587,N_7618);
nand U8266 (N_8266,N_7667,N_7711);
xnor U8267 (N_8267,N_7112,N_7361);
xnor U8268 (N_8268,N_7410,N_7892);
nand U8269 (N_8269,N_7844,N_7916);
or U8270 (N_8270,N_7666,N_7345);
nand U8271 (N_8271,N_7859,N_7001);
nor U8272 (N_8272,N_7134,N_7400);
nand U8273 (N_8273,N_7651,N_7145);
or U8274 (N_8274,N_7159,N_7447);
or U8275 (N_8275,N_7636,N_7522);
and U8276 (N_8276,N_7576,N_7235);
xnor U8277 (N_8277,N_7464,N_7968);
nand U8278 (N_8278,N_7285,N_7652);
and U8279 (N_8279,N_7099,N_7600);
nor U8280 (N_8280,N_7327,N_7546);
nor U8281 (N_8281,N_7807,N_7194);
xor U8282 (N_8282,N_7836,N_7193);
or U8283 (N_8283,N_7685,N_7898);
and U8284 (N_8284,N_7967,N_7102);
and U8285 (N_8285,N_7837,N_7164);
or U8286 (N_8286,N_7876,N_7850);
nor U8287 (N_8287,N_7767,N_7817);
nor U8288 (N_8288,N_7671,N_7132);
nand U8289 (N_8289,N_7409,N_7484);
or U8290 (N_8290,N_7038,N_7258);
nand U8291 (N_8291,N_7959,N_7754);
and U8292 (N_8292,N_7816,N_7453);
xor U8293 (N_8293,N_7248,N_7646);
nor U8294 (N_8294,N_7856,N_7020);
and U8295 (N_8295,N_7565,N_7476);
and U8296 (N_8296,N_7236,N_7663);
xor U8297 (N_8297,N_7095,N_7831);
xor U8298 (N_8298,N_7050,N_7949);
and U8299 (N_8299,N_7945,N_7721);
nand U8300 (N_8300,N_7880,N_7647);
and U8301 (N_8301,N_7451,N_7283);
and U8302 (N_8302,N_7197,N_7829);
nor U8303 (N_8303,N_7838,N_7907);
xor U8304 (N_8304,N_7473,N_7966);
xnor U8305 (N_8305,N_7950,N_7810);
nand U8306 (N_8306,N_7948,N_7170);
or U8307 (N_8307,N_7147,N_7589);
nor U8308 (N_8308,N_7483,N_7376);
and U8309 (N_8309,N_7545,N_7874);
xor U8310 (N_8310,N_7634,N_7084);
or U8311 (N_8311,N_7446,N_7905);
xnor U8312 (N_8312,N_7528,N_7421);
nor U8313 (N_8313,N_7347,N_7594);
and U8314 (N_8314,N_7672,N_7718);
and U8315 (N_8315,N_7855,N_7346);
nor U8316 (N_8316,N_7048,N_7638);
nand U8317 (N_8317,N_7805,N_7760);
or U8318 (N_8318,N_7011,N_7454);
nor U8319 (N_8319,N_7314,N_7631);
xnor U8320 (N_8320,N_7297,N_7686);
nor U8321 (N_8321,N_7616,N_7336);
nor U8322 (N_8322,N_7920,N_7234);
nor U8323 (N_8323,N_7169,N_7840);
nand U8324 (N_8324,N_7547,N_7229);
or U8325 (N_8325,N_7621,N_7465);
and U8326 (N_8326,N_7803,N_7637);
nor U8327 (N_8327,N_7558,N_7172);
nor U8328 (N_8328,N_7946,N_7539);
and U8329 (N_8329,N_7928,N_7456);
xor U8330 (N_8330,N_7355,N_7846);
or U8331 (N_8331,N_7479,N_7679);
nand U8332 (N_8332,N_7841,N_7654);
nand U8333 (N_8333,N_7135,N_7823);
nor U8334 (N_8334,N_7908,N_7531);
or U8335 (N_8335,N_7128,N_7862);
xor U8336 (N_8336,N_7516,N_7612);
nor U8337 (N_8337,N_7515,N_7688);
xor U8338 (N_8338,N_7186,N_7093);
nor U8339 (N_8339,N_7279,N_7626);
or U8340 (N_8340,N_7027,N_7938);
nor U8341 (N_8341,N_7417,N_7998);
xnor U8342 (N_8342,N_7070,N_7381);
nor U8343 (N_8343,N_7434,N_7544);
nor U8344 (N_8344,N_7728,N_7668);
or U8345 (N_8345,N_7131,N_7198);
nor U8346 (N_8346,N_7740,N_7725);
or U8347 (N_8347,N_7622,N_7857);
and U8348 (N_8348,N_7166,N_7341);
nor U8349 (N_8349,N_7595,N_7861);
nand U8350 (N_8350,N_7853,N_7735);
nor U8351 (N_8351,N_7842,N_7500);
nand U8352 (N_8352,N_7256,N_7023);
nor U8353 (N_8353,N_7757,N_7795);
nand U8354 (N_8354,N_7083,N_7849);
xnor U8355 (N_8355,N_7328,N_7030);
and U8356 (N_8356,N_7240,N_7904);
xnor U8357 (N_8357,N_7396,N_7338);
nor U8358 (N_8358,N_7655,N_7930);
nor U8359 (N_8359,N_7257,N_7448);
or U8360 (N_8360,N_7554,N_7424);
or U8361 (N_8361,N_7092,N_7426);
xnor U8362 (N_8362,N_7724,N_7227);
or U8363 (N_8363,N_7296,N_7004);
or U8364 (N_8364,N_7574,N_7541);
nor U8365 (N_8365,N_7259,N_7543);
or U8366 (N_8366,N_7075,N_7174);
xor U8367 (N_8367,N_7161,N_7623);
and U8368 (N_8368,N_7407,N_7997);
xor U8369 (N_8369,N_7028,N_7463);
xor U8370 (N_8370,N_7802,N_7828);
xor U8371 (N_8371,N_7377,N_7935);
nand U8372 (N_8372,N_7365,N_7888);
or U8373 (N_8373,N_7054,N_7065);
nand U8374 (N_8374,N_7053,N_7293);
and U8375 (N_8375,N_7202,N_7747);
xnor U8376 (N_8376,N_7519,N_7474);
nand U8377 (N_8377,N_7035,N_7422);
nor U8378 (N_8378,N_7931,N_7941);
and U8379 (N_8379,N_7579,N_7211);
and U8380 (N_8380,N_7413,N_7322);
nor U8381 (N_8381,N_7173,N_7097);
or U8382 (N_8382,N_7643,N_7423);
nand U8383 (N_8383,N_7538,N_7349);
and U8384 (N_8384,N_7371,N_7738);
nor U8385 (N_8385,N_7357,N_7700);
nand U8386 (N_8386,N_7682,N_7154);
nand U8387 (N_8387,N_7089,N_7601);
nor U8388 (N_8388,N_7786,N_7894);
xnor U8389 (N_8389,N_7420,N_7429);
and U8390 (N_8390,N_7470,N_7024);
nand U8391 (N_8391,N_7743,N_7316);
and U8392 (N_8392,N_7103,N_7824);
nand U8393 (N_8393,N_7675,N_7780);
nor U8394 (N_8394,N_7068,N_7443);
nand U8395 (N_8395,N_7909,N_7117);
xor U8396 (N_8396,N_7965,N_7119);
xor U8397 (N_8397,N_7723,N_7467);
and U8398 (N_8398,N_7425,N_7990);
nor U8399 (N_8399,N_7893,N_7047);
or U8400 (N_8400,N_7088,N_7710);
or U8401 (N_8401,N_7266,N_7329);
xnor U8402 (N_8402,N_7570,N_7241);
xnor U8403 (N_8403,N_7689,N_7777);
or U8404 (N_8404,N_7691,N_7403);
nand U8405 (N_8405,N_7302,N_7353);
nand U8406 (N_8406,N_7408,N_7226);
nor U8407 (N_8407,N_7416,N_7203);
xnor U8408 (N_8408,N_7751,N_7664);
and U8409 (N_8409,N_7146,N_7870);
and U8410 (N_8410,N_7761,N_7356);
nor U8411 (N_8411,N_7163,N_7608);
nor U8412 (N_8412,N_7537,N_7442);
xor U8413 (N_8413,N_7472,N_7865);
and U8414 (N_8414,N_7385,N_7156);
or U8415 (N_8415,N_7684,N_7731);
and U8416 (N_8416,N_7901,N_7605);
nand U8417 (N_8417,N_7061,N_7755);
nor U8418 (N_8418,N_7013,N_7051);
nor U8419 (N_8419,N_7732,N_7046);
and U8420 (N_8420,N_7521,N_7066);
nand U8421 (N_8421,N_7918,N_7970);
xnor U8422 (N_8422,N_7784,N_7578);
and U8423 (N_8423,N_7759,N_7906);
xor U8424 (N_8424,N_7704,N_7320);
xor U8425 (N_8425,N_7580,N_7468);
or U8426 (N_8426,N_7411,N_7043);
nor U8427 (N_8427,N_7126,N_7274);
and U8428 (N_8428,N_7437,N_7800);
or U8429 (N_8429,N_7419,N_7292);
nor U8430 (N_8430,N_7822,N_7926);
or U8431 (N_8431,N_7712,N_7590);
or U8432 (N_8432,N_7224,N_7000);
or U8433 (N_8433,N_7438,N_7942);
xor U8434 (N_8434,N_7656,N_7489);
nand U8435 (N_8435,N_7086,N_7742);
nand U8436 (N_8436,N_7300,N_7504);
nor U8437 (N_8437,N_7375,N_7427);
and U8438 (N_8438,N_7596,N_7010);
xor U8439 (N_8439,N_7933,N_7239);
nand U8440 (N_8440,N_7082,N_7991);
xnor U8441 (N_8441,N_7503,N_7635);
or U8442 (N_8442,N_7080,N_7887);
xor U8443 (N_8443,N_7525,N_7536);
nand U8444 (N_8444,N_7602,N_7641);
and U8445 (N_8445,N_7094,N_7806);
and U8446 (N_8446,N_7116,N_7896);
and U8447 (N_8447,N_7109,N_7354);
or U8448 (N_8448,N_7003,N_7019);
nand U8449 (N_8449,N_7854,N_7370);
or U8450 (N_8450,N_7281,N_7571);
or U8451 (N_8451,N_7954,N_7798);
or U8452 (N_8452,N_7178,N_7719);
or U8453 (N_8453,N_7932,N_7573);
xnor U8454 (N_8454,N_7150,N_7782);
and U8455 (N_8455,N_7978,N_7262);
and U8456 (N_8456,N_7196,N_7055);
nor U8457 (N_8457,N_7108,N_7790);
xnor U8458 (N_8458,N_7532,N_7290);
and U8459 (N_8459,N_7087,N_7485);
or U8460 (N_8460,N_7493,N_7113);
and U8461 (N_8461,N_7653,N_7649);
nand U8462 (N_8462,N_7834,N_7776);
and U8463 (N_8463,N_7264,N_7642);
and U8464 (N_8464,N_7591,N_7059);
or U8465 (N_8465,N_7702,N_7540);
nand U8466 (N_8466,N_7289,N_7496);
nand U8467 (N_8467,N_7015,N_7660);
or U8468 (N_8468,N_7118,N_7364);
nand U8469 (N_8469,N_7091,N_7367);
or U8470 (N_8470,N_7445,N_7287);
and U8471 (N_8471,N_7037,N_7379);
xnor U8472 (N_8472,N_7177,N_7138);
xnor U8473 (N_8473,N_7305,N_7955);
and U8474 (N_8474,N_7628,N_7981);
and U8475 (N_8475,N_7566,N_7444);
nand U8476 (N_8476,N_7752,N_7507);
and U8477 (N_8477,N_7014,N_7678);
xnor U8478 (N_8478,N_7739,N_7209);
nand U8479 (N_8479,N_7040,N_7323);
and U8480 (N_8480,N_7796,N_7633);
and U8481 (N_8481,N_7072,N_7276);
and U8482 (N_8482,N_7559,N_7148);
xor U8483 (N_8483,N_7835,N_7433);
and U8484 (N_8484,N_7650,N_7284);
nand U8485 (N_8485,N_7185,N_7006);
nand U8486 (N_8486,N_7947,N_7779);
nor U8487 (N_8487,N_7247,N_7406);
nand U8488 (N_8488,N_7363,N_7201);
nand U8489 (N_8489,N_7781,N_7162);
nand U8490 (N_8490,N_7556,N_7681);
nor U8491 (N_8491,N_7212,N_7985);
nor U8492 (N_8492,N_7607,N_7142);
or U8493 (N_8493,N_7079,N_7799);
nor U8494 (N_8494,N_7260,N_7511);
nand U8495 (N_8495,N_7312,N_7432);
or U8496 (N_8496,N_7845,N_7956);
nor U8497 (N_8497,N_7141,N_7104);
xnor U8498 (N_8498,N_7133,N_7687);
or U8499 (N_8499,N_7225,N_7120);
and U8500 (N_8500,N_7564,N_7137);
and U8501 (N_8501,N_7908,N_7775);
xor U8502 (N_8502,N_7793,N_7527);
and U8503 (N_8503,N_7282,N_7846);
or U8504 (N_8504,N_7603,N_7643);
or U8505 (N_8505,N_7792,N_7952);
or U8506 (N_8506,N_7000,N_7328);
or U8507 (N_8507,N_7612,N_7463);
and U8508 (N_8508,N_7180,N_7213);
nand U8509 (N_8509,N_7157,N_7615);
and U8510 (N_8510,N_7557,N_7569);
nand U8511 (N_8511,N_7124,N_7101);
nor U8512 (N_8512,N_7460,N_7400);
nand U8513 (N_8513,N_7651,N_7617);
and U8514 (N_8514,N_7054,N_7602);
and U8515 (N_8515,N_7682,N_7105);
xnor U8516 (N_8516,N_7374,N_7122);
nand U8517 (N_8517,N_7712,N_7735);
or U8518 (N_8518,N_7260,N_7282);
nand U8519 (N_8519,N_7339,N_7297);
or U8520 (N_8520,N_7971,N_7430);
nor U8521 (N_8521,N_7045,N_7185);
and U8522 (N_8522,N_7059,N_7541);
xor U8523 (N_8523,N_7448,N_7411);
nor U8524 (N_8524,N_7933,N_7056);
or U8525 (N_8525,N_7858,N_7788);
and U8526 (N_8526,N_7433,N_7696);
and U8527 (N_8527,N_7518,N_7219);
xor U8528 (N_8528,N_7502,N_7094);
and U8529 (N_8529,N_7967,N_7270);
xnor U8530 (N_8530,N_7253,N_7322);
or U8531 (N_8531,N_7970,N_7734);
xor U8532 (N_8532,N_7237,N_7784);
xnor U8533 (N_8533,N_7199,N_7709);
and U8534 (N_8534,N_7960,N_7648);
xnor U8535 (N_8535,N_7685,N_7962);
xor U8536 (N_8536,N_7228,N_7513);
or U8537 (N_8537,N_7448,N_7546);
xor U8538 (N_8538,N_7307,N_7908);
and U8539 (N_8539,N_7612,N_7388);
and U8540 (N_8540,N_7491,N_7759);
and U8541 (N_8541,N_7049,N_7366);
or U8542 (N_8542,N_7102,N_7395);
and U8543 (N_8543,N_7952,N_7687);
nand U8544 (N_8544,N_7210,N_7311);
xor U8545 (N_8545,N_7527,N_7693);
xor U8546 (N_8546,N_7896,N_7636);
or U8547 (N_8547,N_7085,N_7781);
or U8548 (N_8548,N_7887,N_7143);
or U8549 (N_8549,N_7495,N_7881);
nor U8550 (N_8550,N_7520,N_7614);
and U8551 (N_8551,N_7791,N_7765);
nor U8552 (N_8552,N_7681,N_7784);
or U8553 (N_8553,N_7350,N_7701);
nand U8554 (N_8554,N_7669,N_7507);
or U8555 (N_8555,N_7354,N_7204);
nand U8556 (N_8556,N_7766,N_7267);
nor U8557 (N_8557,N_7337,N_7565);
and U8558 (N_8558,N_7450,N_7883);
nor U8559 (N_8559,N_7840,N_7124);
or U8560 (N_8560,N_7972,N_7083);
nor U8561 (N_8561,N_7937,N_7788);
or U8562 (N_8562,N_7599,N_7551);
nor U8563 (N_8563,N_7455,N_7731);
or U8564 (N_8564,N_7704,N_7947);
nand U8565 (N_8565,N_7684,N_7210);
and U8566 (N_8566,N_7935,N_7013);
and U8567 (N_8567,N_7941,N_7692);
and U8568 (N_8568,N_7237,N_7435);
or U8569 (N_8569,N_7560,N_7313);
nor U8570 (N_8570,N_7148,N_7170);
nor U8571 (N_8571,N_7568,N_7925);
or U8572 (N_8572,N_7628,N_7783);
nand U8573 (N_8573,N_7858,N_7892);
xor U8574 (N_8574,N_7071,N_7163);
xor U8575 (N_8575,N_7062,N_7504);
xor U8576 (N_8576,N_7016,N_7495);
nor U8577 (N_8577,N_7220,N_7004);
nand U8578 (N_8578,N_7411,N_7945);
nand U8579 (N_8579,N_7291,N_7644);
or U8580 (N_8580,N_7775,N_7282);
xor U8581 (N_8581,N_7241,N_7986);
nor U8582 (N_8582,N_7594,N_7992);
and U8583 (N_8583,N_7970,N_7345);
xnor U8584 (N_8584,N_7046,N_7357);
and U8585 (N_8585,N_7661,N_7415);
and U8586 (N_8586,N_7192,N_7330);
or U8587 (N_8587,N_7758,N_7054);
and U8588 (N_8588,N_7033,N_7767);
xnor U8589 (N_8589,N_7076,N_7500);
or U8590 (N_8590,N_7806,N_7620);
xor U8591 (N_8591,N_7945,N_7703);
and U8592 (N_8592,N_7844,N_7449);
nand U8593 (N_8593,N_7465,N_7848);
and U8594 (N_8594,N_7303,N_7168);
xnor U8595 (N_8595,N_7286,N_7547);
and U8596 (N_8596,N_7652,N_7790);
nor U8597 (N_8597,N_7037,N_7005);
nor U8598 (N_8598,N_7079,N_7048);
and U8599 (N_8599,N_7900,N_7495);
nor U8600 (N_8600,N_7356,N_7603);
and U8601 (N_8601,N_7497,N_7977);
xor U8602 (N_8602,N_7623,N_7218);
xor U8603 (N_8603,N_7088,N_7000);
nand U8604 (N_8604,N_7617,N_7132);
xnor U8605 (N_8605,N_7630,N_7810);
or U8606 (N_8606,N_7575,N_7938);
nor U8607 (N_8607,N_7033,N_7405);
and U8608 (N_8608,N_7513,N_7899);
xnor U8609 (N_8609,N_7874,N_7045);
or U8610 (N_8610,N_7135,N_7205);
or U8611 (N_8611,N_7470,N_7990);
and U8612 (N_8612,N_7110,N_7611);
and U8613 (N_8613,N_7660,N_7265);
xnor U8614 (N_8614,N_7903,N_7466);
nor U8615 (N_8615,N_7947,N_7419);
and U8616 (N_8616,N_7835,N_7442);
xnor U8617 (N_8617,N_7158,N_7770);
and U8618 (N_8618,N_7212,N_7714);
or U8619 (N_8619,N_7358,N_7570);
and U8620 (N_8620,N_7394,N_7716);
or U8621 (N_8621,N_7641,N_7937);
or U8622 (N_8622,N_7620,N_7024);
nor U8623 (N_8623,N_7391,N_7587);
nand U8624 (N_8624,N_7769,N_7068);
nor U8625 (N_8625,N_7004,N_7077);
xor U8626 (N_8626,N_7947,N_7715);
xnor U8627 (N_8627,N_7557,N_7930);
nand U8628 (N_8628,N_7008,N_7069);
nand U8629 (N_8629,N_7744,N_7352);
and U8630 (N_8630,N_7731,N_7305);
nor U8631 (N_8631,N_7204,N_7640);
nor U8632 (N_8632,N_7908,N_7978);
or U8633 (N_8633,N_7484,N_7972);
and U8634 (N_8634,N_7332,N_7262);
xnor U8635 (N_8635,N_7061,N_7902);
xnor U8636 (N_8636,N_7951,N_7127);
or U8637 (N_8637,N_7376,N_7823);
nor U8638 (N_8638,N_7038,N_7287);
nand U8639 (N_8639,N_7699,N_7501);
nand U8640 (N_8640,N_7735,N_7541);
nand U8641 (N_8641,N_7638,N_7687);
nor U8642 (N_8642,N_7375,N_7405);
nor U8643 (N_8643,N_7418,N_7237);
nor U8644 (N_8644,N_7342,N_7810);
and U8645 (N_8645,N_7717,N_7642);
nand U8646 (N_8646,N_7159,N_7705);
nand U8647 (N_8647,N_7289,N_7486);
or U8648 (N_8648,N_7987,N_7969);
nand U8649 (N_8649,N_7728,N_7975);
nor U8650 (N_8650,N_7630,N_7765);
or U8651 (N_8651,N_7722,N_7626);
or U8652 (N_8652,N_7457,N_7546);
and U8653 (N_8653,N_7819,N_7758);
xor U8654 (N_8654,N_7682,N_7716);
and U8655 (N_8655,N_7169,N_7178);
or U8656 (N_8656,N_7679,N_7552);
nor U8657 (N_8657,N_7078,N_7268);
nor U8658 (N_8658,N_7687,N_7965);
xor U8659 (N_8659,N_7553,N_7560);
or U8660 (N_8660,N_7581,N_7564);
nor U8661 (N_8661,N_7050,N_7066);
or U8662 (N_8662,N_7097,N_7690);
xor U8663 (N_8663,N_7221,N_7438);
and U8664 (N_8664,N_7770,N_7511);
xnor U8665 (N_8665,N_7804,N_7167);
nand U8666 (N_8666,N_7436,N_7341);
or U8667 (N_8667,N_7454,N_7567);
nor U8668 (N_8668,N_7146,N_7423);
and U8669 (N_8669,N_7193,N_7761);
and U8670 (N_8670,N_7301,N_7104);
xnor U8671 (N_8671,N_7058,N_7633);
or U8672 (N_8672,N_7351,N_7664);
nor U8673 (N_8673,N_7948,N_7406);
nand U8674 (N_8674,N_7617,N_7079);
nand U8675 (N_8675,N_7461,N_7051);
or U8676 (N_8676,N_7382,N_7410);
or U8677 (N_8677,N_7336,N_7630);
nand U8678 (N_8678,N_7475,N_7741);
and U8679 (N_8679,N_7615,N_7167);
nor U8680 (N_8680,N_7954,N_7782);
nor U8681 (N_8681,N_7414,N_7994);
or U8682 (N_8682,N_7040,N_7107);
and U8683 (N_8683,N_7647,N_7473);
nand U8684 (N_8684,N_7520,N_7358);
or U8685 (N_8685,N_7315,N_7463);
nor U8686 (N_8686,N_7884,N_7395);
xor U8687 (N_8687,N_7853,N_7400);
or U8688 (N_8688,N_7992,N_7103);
xor U8689 (N_8689,N_7347,N_7542);
nand U8690 (N_8690,N_7673,N_7898);
or U8691 (N_8691,N_7106,N_7170);
nand U8692 (N_8692,N_7934,N_7254);
or U8693 (N_8693,N_7285,N_7255);
xnor U8694 (N_8694,N_7838,N_7115);
nand U8695 (N_8695,N_7968,N_7276);
nand U8696 (N_8696,N_7193,N_7629);
and U8697 (N_8697,N_7352,N_7431);
xnor U8698 (N_8698,N_7723,N_7494);
or U8699 (N_8699,N_7446,N_7857);
and U8700 (N_8700,N_7745,N_7685);
nor U8701 (N_8701,N_7294,N_7021);
or U8702 (N_8702,N_7145,N_7299);
or U8703 (N_8703,N_7834,N_7684);
nand U8704 (N_8704,N_7377,N_7961);
xor U8705 (N_8705,N_7371,N_7431);
nand U8706 (N_8706,N_7168,N_7477);
nand U8707 (N_8707,N_7583,N_7517);
nor U8708 (N_8708,N_7719,N_7068);
or U8709 (N_8709,N_7200,N_7440);
nand U8710 (N_8710,N_7771,N_7041);
nand U8711 (N_8711,N_7294,N_7945);
or U8712 (N_8712,N_7658,N_7295);
nor U8713 (N_8713,N_7596,N_7233);
nand U8714 (N_8714,N_7326,N_7884);
nand U8715 (N_8715,N_7473,N_7366);
or U8716 (N_8716,N_7114,N_7211);
nand U8717 (N_8717,N_7688,N_7347);
and U8718 (N_8718,N_7136,N_7801);
nor U8719 (N_8719,N_7718,N_7095);
and U8720 (N_8720,N_7319,N_7599);
or U8721 (N_8721,N_7973,N_7346);
or U8722 (N_8722,N_7486,N_7617);
or U8723 (N_8723,N_7617,N_7623);
or U8724 (N_8724,N_7629,N_7360);
or U8725 (N_8725,N_7899,N_7047);
nand U8726 (N_8726,N_7219,N_7227);
nor U8727 (N_8727,N_7194,N_7109);
or U8728 (N_8728,N_7556,N_7534);
and U8729 (N_8729,N_7466,N_7908);
nand U8730 (N_8730,N_7219,N_7511);
nand U8731 (N_8731,N_7143,N_7685);
or U8732 (N_8732,N_7140,N_7321);
and U8733 (N_8733,N_7205,N_7570);
or U8734 (N_8734,N_7032,N_7393);
nor U8735 (N_8735,N_7160,N_7833);
xnor U8736 (N_8736,N_7084,N_7737);
and U8737 (N_8737,N_7833,N_7695);
nand U8738 (N_8738,N_7845,N_7918);
xnor U8739 (N_8739,N_7622,N_7849);
xor U8740 (N_8740,N_7847,N_7864);
nand U8741 (N_8741,N_7190,N_7048);
xnor U8742 (N_8742,N_7878,N_7657);
or U8743 (N_8743,N_7632,N_7072);
xor U8744 (N_8744,N_7049,N_7706);
nor U8745 (N_8745,N_7462,N_7156);
nand U8746 (N_8746,N_7928,N_7378);
and U8747 (N_8747,N_7257,N_7495);
or U8748 (N_8748,N_7098,N_7947);
and U8749 (N_8749,N_7624,N_7702);
nand U8750 (N_8750,N_7448,N_7321);
and U8751 (N_8751,N_7685,N_7168);
nor U8752 (N_8752,N_7907,N_7226);
xor U8753 (N_8753,N_7718,N_7833);
xnor U8754 (N_8754,N_7012,N_7665);
and U8755 (N_8755,N_7171,N_7472);
nand U8756 (N_8756,N_7074,N_7647);
and U8757 (N_8757,N_7939,N_7762);
xnor U8758 (N_8758,N_7811,N_7114);
or U8759 (N_8759,N_7951,N_7562);
nor U8760 (N_8760,N_7561,N_7211);
nand U8761 (N_8761,N_7935,N_7433);
and U8762 (N_8762,N_7235,N_7664);
xnor U8763 (N_8763,N_7325,N_7954);
nor U8764 (N_8764,N_7950,N_7110);
nand U8765 (N_8765,N_7882,N_7888);
nor U8766 (N_8766,N_7678,N_7729);
nor U8767 (N_8767,N_7223,N_7459);
and U8768 (N_8768,N_7017,N_7675);
nand U8769 (N_8769,N_7964,N_7853);
and U8770 (N_8770,N_7141,N_7662);
or U8771 (N_8771,N_7540,N_7137);
nand U8772 (N_8772,N_7082,N_7332);
nor U8773 (N_8773,N_7795,N_7696);
xor U8774 (N_8774,N_7454,N_7418);
nand U8775 (N_8775,N_7969,N_7337);
and U8776 (N_8776,N_7791,N_7704);
and U8777 (N_8777,N_7184,N_7229);
and U8778 (N_8778,N_7329,N_7181);
nand U8779 (N_8779,N_7462,N_7308);
xnor U8780 (N_8780,N_7067,N_7112);
or U8781 (N_8781,N_7543,N_7793);
nor U8782 (N_8782,N_7350,N_7002);
nor U8783 (N_8783,N_7219,N_7717);
and U8784 (N_8784,N_7145,N_7207);
nand U8785 (N_8785,N_7101,N_7719);
nand U8786 (N_8786,N_7067,N_7012);
xor U8787 (N_8787,N_7261,N_7380);
nand U8788 (N_8788,N_7684,N_7347);
and U8789 (N_8789,N_7907,N_7157);
nand U8790 (N_8790,N_7073,N_7205);
or U8791 (N_8791,N_7838,N_7949);
xnor U8792 (N_8792,N_7986,N_7899);
nand U8793 (N_8793,N_7118,N_7475);
xnor U8794 (N_8794,N_7319,N_7447);
nand U8795 (N_8795,N_7810,N_7927);
or U8796 (N_8796,N_7309,N_7523);
xor U8797 (N_8797,N_7180,N_7614);
nor U8798 (N_8798,N_7218,N_7611);
nand U8799 (N_8799,N_7995,N_7708);
nor U8800 (N_8800,N_7979,N_7964);
or U8801 (N_8801,N_7406,N_7565);
nand U8802 (N_8802,N_7842,N_7063);
nand U8803 (N_8803,N_7146,N_7800);
nand U8804 (N_8804,N_7271,N_7755);
or U8805 (N_8805,N_7520,N_7386);
nand U8806 (N_8806,N_7123,N_7631);
xor U8807 (N_8807,N_7776,N_7742);
and U8808 (N_8808,N_7165,N_7224);
xor U8809 (N_8809,N_7267,N_7392);
nor U8810 (N_8810,N_7880,N_7891);
nor U8811 (N_8811,N_7694,N_7262);
or U8812 (N_8812,N_7197,N_7415);
or U8813 (N_8813,N_7484,N_7001);
and U8814 (N_8814,N_7056,N_7550);
or U8815 (N_8815,N_7945,N_7441);
nand U8816 (N_8816,N_7755,N_7659);
nand U8817 (N_8817,N_7579,N_7392);
or U8818 (N_8818,N_7850,N_7786);
and U8819 (N_8819,N_7984,N_7730);
nand U8820 (N_8820,N_7144,N_7986);
xnor U8821 (N_8821,N_7534,N_7376);
nand U8822 (N_8822,N_7926,N_7141);
nand U8823 (N_8823,N_7389,N_7771);
nand U8824 (N_8824,N_7281,N_7775);
or U8825 (N_8825,N_7622,N_7311);
nor U8826 (N_8826,N_7258,N_7133);
nand U8827 (N_8827,N_7182,N_7778);
and U8828 (N_8828,N_7913,N_7274);
xnor U8829 (N_8829,N_7368,N_7698);
or U8830 (N_8830,N_7348,N_7284);
nand U8831 (N_8831,N_7941,N_7780);
and U8832 (N_8832,N_7509,N_7978);
and U8833 (N_8833,N_7752,N_7305);
nand U8834 (N_8834,N_7359,N_7260);
xor U8835 (N_8835,N_7444,N_7653);
or U8836 (N_8836,N_7159,N_7472);
nor U8837 (N_8837,N_7842,N_7615);
and U8838 (N_8838,N_7120,N_7735);
and U8839 (N_8839,N_7572,N_7283);
and U8840 (N_8840,N_7332,N_7804);
nand U8841 (N_8841,N_7824,N_7494);
or U8842 (N_8842,N_7854,N_7702);
nor U8843 (N_8843,N_7476,N_7179);
nor U8844 (N_8844,N_7621,N_7315);
nor U8845 (N_8845,N_7186,N_7269);
xor U8846 (N_8846,N_7045,N_7032);
and U8847 (N_8847,N_7525,N_7195);
nor U8848 (N_8848,N_7694,N_7226);
nand U8849 (N_8849,N_7937,N_7666);
nand U8850 (N_8850,N_7756,N_7957);
xnor U8851 (N_8851,N_7734,N_7639);
and U8852 (N_8852,N_7826,N_7464);
nand U8853 (N_8853,N_7316,N_7286);
and U8854 (N_8854,N_7818,N_7461);
xor U8855 (N_8855,N_7146,N_7814);
and U8856 (N_8856,N_7710,N_7157);
xor U8857 (N_8857,N_7203,N_7894);
xnor U8858 (N_8858,N_7448,N_7463);
nand U8859 (N_8859,N_7519,N_7622);
xor U8860 (N_8860,N_7546,N_7203);
nor U8861 (N_8861,N_7755,N_7786);
nor U8862 (N_8862,N_7083,N_7260);
xor U8863 (N_8863,N_7269,N_7580);
or U8864 (N_8864,N_7644,N_7251);
nor U8865 (N_8865,N_7660,N_7720);
nor U8866 (N_8866,N_7502,N_7079);
or U8867 (N_8867,N_7847,N_7745);
nand U8868 (N_8868,N_7439,N_7844);
nand U8869 (N_8869,N_7661,N_7017);
xnor U8870 (N_8870,N_7824,N_7198);
xnor U8871 (N_8871,N_7561,N_7604);
or U8872 (N_8872,N_7126,N_7020);
or U8873 (N_8873,N_7370,N_7502);
xor U8874 (N_8874,N_7916,N_7547);
xor U8875 (N_8875,N_7974,N_7139);
nor U8876 (N_8876,N_7751,N_7757);
nand U8877 (N_8877,N_7266,N_7395);
nand U8878 (N_8878,N_7721,N_7296);
and U8879 (N_8879,N_7126,N_7141);
nand U8880 (N_8880,N_7714,N_7236);
and U8881 (N_8881,N_7948,N_7423);
nand U8882 (N_8882,N_7810,N_7943);
nand U8883 (N_8883,N_7257,N_7992);
nor U8884 (N_8884,N_7399,N_7368);
or U8885 (N_8885,N_7738,N_7900);
nand U8886 (N_8886,N_7302,N_7402);
or U8887 (N_8887,N_7774,N_7738);
and U8888 (N_8888,N_7862,N_7104);
nor U8889 (N_8889,N_7453,N_7867);
and U8890 (N_8890,N_7350,N_7643);
or U8891 (N_8891,N_7213,N_7906);
xnor U8892 (N_8892,N_7754,N_7780);
xor U8893 (N_8893,N_7559,N_7912);
nor U8894 (N_8894,N_7327,N_7443);
xor U8895 (N_8895,N_7492,N_7915);
xnor U8896 (N_8896,N_7658,N_7853);
nor U8897 (N_8897,N_7381,N_7955);
nor U8898 (N_8898,N_7766,N_7301);
nor U8899 (N_8899,N_7251,N_7005);
or U8900 (N_8900,N_7251,N_7259);
nand U8901 (N_8901,N_7946,N_7422);
or U8902 (N_8902,N_7199,N_7864);
nand U8903 (N_8903,N_7474,N_7247);
and U8904 (N_8904,N_7223,N_7452);
nor U8905 (N_8905,N_7916,N_7223);
and U8906 (N_8906,N_7922,N_7141);
or U8907 (N_8907,N_7337,N_7594);
xnor U8908 (N_8908,N_7271,N_7121);
or U8909 (N_8909,N_7792,N_7421);
xor U8910 (N_8910,N_7431,N_7817);
xnor U8911 (N_8911,N_7540,N_7264);
or U8912 (N_8912,N_7309,N_7971);
and U8913 (N_8913,N_7081,N_7485);
or U8914 (N_8914,N_7334,N_7603);
xnor U8915 (N_8915,N_7883,N_7041);
nor U8916 (N_8916,N_7776,N_7731);
xnor U8917 (N_8917,N_7773,N_7297);
nor U8918 (N_8918,N_7306,N_7978);
nand U8919 (N_8919,N_7032,N_7891);
and U8920 (N_8920,N_7279,N_7537);
and U8921 (N_8921,N_7654,N_7919);
nand U8922 (N_8922,N_7002,N_7990);
and U8923 (N_8923,N_7268,N_7852);
or U8924 (N_8924,N_7872,N_7400);
and U8925 (N_8925,N_7334,N_7384);
xor U8926 (N_8926,N_7925,N_7088);
nand U8927 (N_8927,N_7485,N_7634);
xor U8928 (N_8928,N_7981,N_7322);
xor U8929 (N_8929,N_7698,N_7324);
nor U8930 (N_8930,N_7799,N_7826);
nand U8931 (N_8931,N_7097,N_7494);
and U8932 (N_8932,N_7928,N_7009);
nand U8933 (N_8933,N_7910,N_7271);
nand U8934 (N_8934,N_7071,N_7682);
nor U8935 (N_8935,N_7950,N_7343);
xor U8936 (N_8936,N_7220,N_7694);
nor U8937 (N_8937,N_7965,N_7398);
nand U8938 (N_8938,N_7232,N_7225);
nand U8939 (N_8939,N_7534,N_7761);
and U8940 (N_8940,N_7679,N_7396);
nand U8941 (N_8941,N_7954,N_7741);
nand U8942 (N_8942,N_7910,N_7027);
xor U8943 (N_8943,N_7364,N_7803);
nor U8944 (N_8944,N_7112,N_7660);
nor U8945 (N_8945,N_7066,N_7944);
nor U8946 (N_8946,N_7559,N_7908);
nand U8947 (N_8947,N_7655,N_7066);
and U8948 (N_8948,N_7538,N_7684);
xnor U8949 (N_8949,N_7951,N_7561);
xnor U8950 (N_8950,N_7099,N_7722);
and U8951 (N_8951,N_7587,N_7510);
or U8952 (N_8952,N_7080,N_7915);
and U8953 (N_8953,N_7239,N_7483);
or U8954 (N_8954,N_7518,N_7725);
xnor U8955 (N_8955,N_7109,N_7446);
and U8956 (N_8956,N_7229,N_7655);
and U8957 (N_8957,N_7004,N_7065);
or U8958 (N_8958,N_7150,N_7672);
nand U8959 (N_8959,N_7584,N_7638);
xor U8960 (N_8960,N_7404,N_7703);
and U8961 (N_8961,N_7597,N_7899);
nor U8962 (N_8962,N_7767,N_7202);
and U8963 (N_8963,N_7337,N_7181);
and U8964 (N_8964,N_7293,N_7794);
xnor U8965 (N_8965,N_7794,N_7060);
nand U8966 (N_8966,N_7971,N_7950);
nor U8967 (N_8967,N_7256,N_7117);
nand U8968 (N_8968,N_7083,N_7962);
nor U8969 (N_8969,N_7239,N_7667);
and U8970 (N_8970,N_7858,N_7259);
nand U8971 (N_8971,N_7554,N_7453);
xor U8972 (N_8972,N_7038,N_7218);
xnor U8973 (N_8973,N_7538,N_7818);
nor U8974 (N_8974,N_7790,N_7863);
or U8975 (N_8975,N_7991,N_7448);
nand U8976 (N_8976,N_7373,N_7630);
xnor U8977 (N_8977,N_7254,N_7490);
xnor U8978 (N_8978,N_7443,N_7032);
or U8979 (N_8979,N_7734,N_7918);
nor U8980 (N_8980,N_7074,N_7947);
nand U8981 (N_8981,N_7949,N_7830);
or U8982 (N_8982,N_7389,N_7709);
xor U8983 (N_8983,N_7937,N_7145);
and U8984 (N_8984,N_7541,N_7956);
xnor U8985 (N_8985,N_7726,N_7711);
nor U8986 (N_8986,N_7761,N_7859);
nand U8987 (N_8987,N_7617,N_7070);
and U8988 (N_8988,N_7855,N_7338);
xnor U8989 (N_8989,N_7259,N_7525);
nand U8990 (N_8990,N_7983,N_7728);
or U8991 (N_8991,N_7570,N_7914);
nand U8992 (N_8992,N_7733,N_7137);
xor U8993 (N_8993,N_7101,N_7762);
nand U8994 (N_8994,N_7412,N_7348);
nand U8995 (N_8995,N_7717,N_7452);
nand U8996 (N_8996,N_7328,N_7802);
nor U8997 (N_8997,N_7630,N_7391);
nand U8998 (N_8998,N_7070,N_7675);
nor U8999 (N_8999,N_7375,N_7551);
and U9000 (N_9000,N_8655,N_8549);
nor U9001 (N_9001,N_8315,N_8845);
nor U9002 (N_9002,N_8042,N_8821);
nor U9003 (N_9003,N_8388,N_8959);
nand U9004 (N_9004,N_8202,N_8383);
and U9005 (N_9005,N_8810,N_8634);
or U9006 (N_9006,N_8924,N_8505);
nand U9007 (N_9007,N_8559,N_8840);
and U9008 (N_9008,N_8292,N_8771);
and U9009 (N_9009,N_8744,N_8417);
nand U9010 (N_9010,N_8266,N_8467);
nor U9011 (N_9011,N_8367,N_8408);
nor U9012 (N_9012,N_8158,N_8069);
or U9013 (N_9013,N_8349,N_8950);
or U9014 (N_9014,N_8874,N_8426);
xnor U9015 (N_9015,N_8486,N_8766);
and U9016 (N_9016,N_8477,N_8431);
or U9017 (N_9017,N_8329,N_8418);
xnor U9018 (N_9018,N_8360,N_8747);
and U9019 (N_9019,N_8446,N_8900);
or U9020 (N_9020,N_8003,N_8304);
nor U9021 (N_9021,N_8673,N_8465);
or U9022 (N_9022,N_8974,N_8098);
nand U9023 (N_9023,N_8853,N_8931);
nor U9024 (N_9024,N_8822,N_8186);
and U9025 (N_9025,N_8863,N_8200);
nand U9026 (N_9026,N_8272,N_8730);
nor U9027 (N_9027,N_8935,N_8632);
or U9028 (N_9028,N_8541,N_8084);
nand U9029 (N_9029,N_8251,N_8770);
or U9030 (N_9030,N_8263,N_8926);
and U9031 (N_9031,N_8111,N_8313);
or U9032 (N_9032,N_8048,N_8796);
xnor U9033 (N_9033,N_8011,N_8547);
or U9034 (N_9034,N_8018,N_8551);
nand U9035 (N_9035,N_8583,N_8658);
xor U9036 (N_9036,N_8455,N_8737);
nand U9037 (N_9037,N_8289,N_8253);
nor U9038 (N_9038,N_8414,N_8219);
and U9039 (N_9039,N_8957,N_8882);
nand U9040 (N_9040,N_8654,N_8509);
nand U9041 (N_9041,N_8090,N_8904);
or U9042 (N_9042,N_8270,N_8144);
and U9043 (N_9043,N_8193,N_8682);
nand U9044 (N_9044,N_8601,N_8185);
nor U9045 (N_9045,N_8085,N_8861);
xnor U9046 (N_9046,N_8035,N_8110);
nand U9047 (N_9047,N_8476,N_8621);
nor U9048 (N_9048,N_8793,N_8996);
and U9049 (N_9049,N_8390,N_8459);
or U9050 (N_9050,N_8079,N_8045);
nor U9051 (N_9051,N_8819,N_8841);
and U9052 (N_9052,N_8129,N_8762);
xnor U9053 (N_9053,N_8539,N_8320);
nand U9054 (N_9054,N_8948,N_8553);
nor U9055 (N_9055,N_8433,N_8576);
or U9056 (N_9056,N_8855,N_8648);
and U9057 (N_9057,N_8457,N_8005);
nand U9058 (N_9058,N_8319,N_8076);
nor U9059 (N_9059,N_8914,N_8293);
nor U9060 (N_9060,N_8680,N_8103);
nand U9061 (N_9061,N_8578,N_8381);
and U9062 (N_9062,N_8517,N_8141);
nand U9063 (N_9063,N_8019,N_8759);
xor U9064 (N_9064,N_8557,N_8925);
nand U9065 (N_9065,N_8222,N_8000);
xnor U9066 (N_9066,N_8617,N_8975);
nor U9067 (N_9067,N_8223,N_8120);
and U9068 (N_9068,N_8432,N_8366);
nand U9069 (N_9069,N_8218,N_8732);
or U9070 (N_9070,N_8661,N_8310);
xnor U9071 (N_9071,N_8858,N_8579);
xnor U9072 (N_9072,N_8735,N_8561);
and U9073 (N_9073,N_8269,N_8083);
or U9074 (N_9074,N_8848,N_8058);
and U9075 (N_9075,N_8512,N_8183);
nand U9076 (N_9076,N_8958,N_8402);
and U9077 (N_9077,N_8976,N_8365);
nor U9078 (N_9078,N_8754,N_8462);
nand U9079 (N_9079,N_8247,N_8811);
and U9080 (N_9080,N_8154,N_8729);
or U9081 (N_9081,N_8839,N_8258);
or U9082 (N_9082,N_8241,N_8679);
or U9083 (N_9083,N_8441,N_8898);
or U9084 (N_9084,N_8394,N_8142);
and U9085 (N_9085,N_8884,N_8508);
or U9086 (N_9086,N_8693,N_8635);
or U9087 (N_9087,N_8677,N_8734);
xnor U9088 (N_9088,N_8830,N_8104);
xnor U9089 (N_9089,N_8236,N_8833);
or U9090 (N_9090,N_8943,N_8808);
or U9091 (N_9091,N_8453,N_8343);
nand U9092 (N_9092,N_8697,N_8955);
nand U9093 (N_9093,N_8472,N_8335);
and U9094 (N_9094,N_8502,N_8212);
xnor U9095 (N_9095,N_8751,N_8739);
and U9096 (N_9096,N_8540,N_8178);
nor U9097 (N_9097,N_8772,N_8849);
and U9098 (N_9098,N_8448,N_8043);
and U9099 (N_9099,N_8930,N_8741);
or U9100 (N_9100,N_8887,N_8073);
or U9101 (N_9101,N_8731,N_8618);
or U9102 (N_9102,N_8125,N_8061);
xor U9103 (N_9103,N_8750,N_8067);
xor U9104 (N_9104,N_8988,N_8716);
and U9105 (N_9105,N_8143,N_8702);
or U9106 (N_9106,N_8795,N_8938);
and U9107 (N_9107,N_8978,N_8020);
or U9108 (N_9108,N_8967,N_8317);
and U9109 (N_9109,N_8445,N_8851);
nand U9110 (N_9110,N_8769,N_8657);
xnor U9111 (N_9111,N_8574,N_8033);
or U9112 (N_9112,N_8286,N_8917);
nor U9113 (N_9113,N_8006,N_8603);
and U9114 (N_9114,N_8554,N_8646);
xnor U9115 (N_9115,N_8893,N_8080);
or U9116 (N_9116,N_8789,N_8639);
nor U9117 (N_9117,N_8375,N_8086);
nand U9118 (N_9118,N_8806,N_8447);
xnor U9119 (N_9119,N_8867,N_8273);
or U9120 (N_9120,N_8026,N_8382);
and U9121 (N_9121,N_8131,N_8520);
and U9122 (N_9122,N_8609,N_8591);
nand U9123 (N_9123,N_8587,N_8350);
and U9124 (N_9124,N_8815,N_8303);
and U9125 (N_9125,N_8667,N_8225);
nor U9126 (N_9126,N_8279,N_8473);
and U9127 (N_9127,N_8624,N_8514);
and U9128 (N_9128,N_8182,N_8555);
or U9129 (N_9129,N_8719,N_8036);
nor U9130 (N_9130,N_8786,N_8485);
xnor U9131 (N_9131,N_8596,N_8107);
and U9132 (N_9132,N_8545,N_8101);
nor U9133 (N_9133,N_8281,N_8153);
nand U9134 (N_9134,N_8507,N_8877);
or U9135 (N_9135,N_8009,N_8985);
and U9136 (N_9136,N_8322,N_8074);
and U9137 (N_9137,N_8314,N_8167);
nand U9138 (N_9138,N_8643,N_8044);
or U9139 (N_9139,N_8029,N_8162);
and U9140 (N_9140,N_8865,N_8892);
or U9141 (N_9141,N_8179,N_8911);
xnor U9142 (N_9142,N_8929,N_8450);
xnor U9143 (N_9143,N_8704,N_8136);
and U9144 (N_9144,N_8715,N_8664);
nor U9145 (N_9145,N_8072,N_8788);
nand U9146 (N_9146,N_8169,N_8238);
nand U9147 (N_9147,N_8740,N_8267);
or U9148 (N_9148,N_8933,N_8638);
xnor U9149 (N_9149,N_8565,N_8548);
xor U9150 (N_9150,N_8568,N_8790);
nor U9151 (N_9151,N_8296,N_8049);
xor U9152 (N_9152,N_8246,N_8971);
nand U9153 (N_9153,N_8259,N_8387);
nand U9154 (N_9154,N_8922,N_8139);
nor U9155 (N_9155,N_8669,N_8207);
and U9156 (N_9156,N_8665,N_8653);
nor U9157 (N_9157,N_8767,N_8905);
xor U9158 (N_9158,N_8992,N_8582);
and U9159 (N_9159,N_8093,N_8916);
nor U9160 (N_9160,N_8331,N_8452);
xnor U9161 (N_9161,N_8660,N_8965);
xnor U9162 (N_9162,N_8599,N_8172);
nor U9163 (N_9163,N_8017,N_8945);
xnor U9164 (N_9164,N_8023,N_8175);
xor U9165 (N_9165,N_8411,N_8969);
nor U9166 (N_9166,N_8434,N_8336);
or U9167 (N_9167,N_8829,N_8340);
xor U9168 (N_9168,N_8990,N_8530);
or U9169 (N_9169,N_8590,N_8358);
nand U9170 (N_9170,N_8287,N_8250);
nand U9171 (N_9171,N_8002,N_8210);
xor U9172 (N_9172,N_8181,N_8245);
xor U9173 (N_9173,N_8818,N_8598);
or U9174 (N_9174,N_8531,N_8135);
and U9175 (N_9175,N_8866,N_8393);
nand U9176 (N_9176,N_8326,N_8312);
and U9177 (N_9177,N_8989,N_8252);
nor U9178 (N_9178,N_8161,N_8150);
xor U9179 (N_9179,N_8297,N_8337);
nand U9180 (N_9180,N_8413,N_8610);
and U9181 (N_9181,N_8055,N_8435);
or U9182 (N_9182,N_8717,N_8666);
and U9183 (N_9183,N_8616,N_8500);
nor U9184 (N_9184,N_8983,N_8984);
or U9185 (N_9185,N_8956,N_8600);
or U9186 (N_9186,N_8742,N_8470);
or U9187 (N_9187,N_8763,N_8592);
xnor U9188 (N_9188,N_8012,N_8152);
nor U9189 (N_9189,N_8968,N_8440);
nor U9190 (N_9190,N_8577,N_8112);
nor U9191 (N_9191,N_8588,N_8961);
and U9192 (N_9192,N_8379,N_8323);
nand U9193 (N_9193,N_8464,N_8195);
xnor U9194 (N_9194,N_8886,N_8890);
and U9195 (N_9195,N_8306,N_8092);
nor U9196 (N_9196,N_8949,N_8525);
nor U9197 (N_9197,N_8928,N_8755);
and U9198 (N_9198,N_8235,N_8628);
nor U9199 (N_9199,N_8897,N_8506);
xnor U9200 (N_9200,N_8982,N_8234);
xor U9201 (N_9201,N_8403,N_8163);
or U9202 (N_9202,N_8145,N_8690);
and U9203 (N_9203,N_8889,N_8451);
xnor U9204 (N_9204,N_8825,N_8007);
and U9205 (N_9205,N_8176,N_8998);
nand U9206 (N_9206,N_8149,N_8558);
nand U9207 (N_9207,N_8799,N_8567);
or U9208 (N_9208,N_8339,N_8856);
xor U9209 (N_9209,N_8781,N_8670);
nor U9210 (N_9210,N_8116,N_8436);
nor U9211 (N_9211,N_8255,N_8230);
and U9212 (N_9212,N_8108,N_8995);
and U9213 (N_9213,N_8311,N_8407);
nor U9214 (N_9214,N_8993,N_8140);
nor U9215 (N_9215,N_8761,N_8484);
xnor U9216 (N_9216,N_8333,N_8787);
xnor U9217 (N_9217,N_8096,N_8089);
and U9218 (N_9218,N_8792,N_8901);
nor U9219 (N_9219,N_8416,N_8777);
nand U9220 (N_9220,N_8823,N_8663);
or U9221 (N_9221,N_8947,N_8529);
xnor U9222 (N_9222,N_8695,N_8205);
nor U9223 (N_9223,N_8121,N_8834);
nand U9224 (N_9224,N_8208,N_8535);
nor U9225 (N_9225,N_8233,N_8981);
nor U9226 (N_9226,N_8156,N_8921);
or U9227 (N_9227,N_8791,N_8994);
nor U9228 (N_9228,N_8564,N_8878);
or U9229 (N_9229,N_8391,N_8174);
or U9230 (N_9230,N_8052,N_8952);
xor U9231 (N_9231,N_8873,N_8997);
or U9232 (N_9232,N_8720,N_8868);
and U9233 (N_9233,N_8030,N_8875);
and U9234 (N_9234,N_8124,N_8626);
nand U9235 (N_9235,N_8261,N_8423);
xor U9236 (N_9236,N_8608,N_8062);
nand U9237 (N_9237,N_8429,N_8907);
and U9238 (N_9238,N_8262,N_8113);
and U9239 (N_9239,N_8344,N_8619);
or U9240 (N_9240,N_8516,N_8078);
and U9241 (N_9241,N_8797,N_8571);
nor U9242 (N_9242,N_8209,N_8039);
xnor U9243 (N_9243,N_8854,N_8271);
xor U9244 (N_9244,N_8710,N_8798);
xor U9245 (N_9245,N_8134,N_8275);
nor U9246 (N_9246,N_8521,N_8338);
nand U9247 (N_9247,N_8649,N_8395);
nor U9248 (N_9248,N_8040,N_8920);
nand U9249 (N_9249,N_8180,N_8910);
and U9250 (N_9250,N_8479,N_8082);
or U9251 (N_9251,N_8016,N_8686);
or U9252 (N_9252,N_8902,N_8494);
or U9253 (N_9253,N_8392,N_8065);
nor U9254 (N_9254,N_8115,N_8187);
nor U9255 (N_9255,N_8063,N_8895);
or U9256 (N_9256,N_8515,N_8779);
and U9257 (N_9257,N_8492,N_8325);
nand U9258 (N_9258,N_8231,N_8691);
or U9259 (N_9259,N_8157,N_8227);
and U9260 (N_9260,N_8964,N_8188);
xnor U9261 (N_9261,N_8192,N_8427);
or U9262 (N_9262,N_8449,N_8249);
xor U9263 (N_9263,N_8242,N_8166);
nand U9264 (N_9264,N_8733,N_8087);
nand U9265 (N_9265,N_8370,N_8217);
nor U9266 (N_9266,N_8454,N_8784);
nand U9267 (N_9267,N_8243,N_8405);
nand U9268 (N_9268,N_8444,N_8357);
nor U9269 (N_9269,N_8378,N_8102);
nand U9270 (N_9270,N_8501,N_8363);
xnor U9271 (N_9271,N_8345,N_8780);
nor U9272 (N_9272,N_8847,N_8756);
or U9273 (N_9273,N_8305,N_8004);
and U9274 (N_9274,N_8400,N_8294);
nand U9275 (N_9275,N_8346,N_8630);
nor U9276 (N_9276,N_8291,N_8586);
nor U9277 (N_9277,N_8528,N_8936);
or U9278 (N_9278,N_8511,N_8031);
xnor U9279 (N_9279,N_8652,N_8778);
xnor U9280 (N_9280,N_8420,N_8064);
or U9281 (N_9281,N_8024,N_8972);
xor U9282 (N_9282,N_8355,N_8836);
and U9283 (N_9283,N_8300,N_8773);
and U9284 (N_9284,N_8199,N_8354);
nor U9285 (N_9285,N_8700,N_8694);
or U9286 (N_9286,N_8721,N_8838);
nor U9287 (N_9287,N_8748,N_8097);
nand U9288 (N_9288,N_8672,N_8524);
and U9289 (N_9289,N_8569,N_8196);
and U9290 (N_9290,N_8268,N_8475);
xor U9291 (N_9291,N_8912,N_8216);
and U9292 (N_9292,N_8859,N_8490);
nor U9293 (N_9293,N_8119,N_8683);
nor U9294 (N_9294,N_8523,N_8862);
nor U9295 (N_9295,N_8832,N_8749);
or U9296 (N_9296,N_8842,N_8321);
or U9297 (N_9297,N_8232,N_8527);
or U9298 (N_9298,N_8348,N_8605);
and U9299 (N_9299,N_8668,N_8692);
and U9300 (N_9300,N_8099,N_8510);
or U9301 (N_9301,N_8059,N_8909);
xor U9302 (N_9302,N_8341,N_8977);
and U9303 (N_9303,N_8334,N_8768);
xor U9304 (N_9304,N_8896,N_8491);
nand U9305 (N_9305,N_8412,N_8155);
nor U9306 (N_9306,N_8211,N_8659);
and U9307 (N_9307,N_8533,N_8709);
and U9308 (N_9308,N_8633,N_8960);
and U9309 (N_9309,N_8128,N_8330);
nand U9310 (N_9310,N_8194,N_8913);
nor U9311 (N_9311,N_8264,N_8359);
nand U9312 (N_9312,N_8637,N_8147);
or U9313 (N_9313,N_8021,N_8206);
nor U9314 (N_9314,N_8594,N_8151);
xnor U9315 (N_9315,N_8871,N_8148);
xnor U9316 (N_9316,N_8973,N_8274);
nand U9317 (N_9317,N_8708,N_8308);
xor U9318 (N_9318,N_8932,N_8718);
nor U9319 (N_9319,N_8642,N_8425);
or U9320 (N_9320,N_8309,N_8437);
nand U9321 (N_9321,N_8572,N_8927);
xor U9322 (N_9322,N_8595,N_8872);
nand U9323 (N_9323,N_8474,N_8220);
and U9324 (N_9324,N_8037,N_8864);
and U9325 (N_9325,N_8999,N_8712);
and U9326 (N_9326,N_8372,N_8229);
or U9327 (N_9327,N_8891,N_8239);
or U9328 (N_9328,N_8461,N_8614);
xor U9329 (N_9329,N_8537,N_8597);
xor U9330 (N_9330,N_8644,N_8689);
xnor U9331 (N_9331,N_8068,N_8100);
nor U9332 (N_9332,N_8575,N_8438);
or U9333 (N_9333,N_8463,N_8738);
nor U9334 (N_9334,N_8805,N_8226);
nand U9335 (N_9335,N_8589,N_8204);
and U9336 (N_9336,N_8585,N_8640);
nand U9337 (N_9337,N_8368,N_8481);
nand U9338 (N_9338,N_8177,N_8880);
or U9339 (N_9339,N_8809,N_8852);
and U9340 (N_9340,N_8028,N_8816);
or U9341 (N_9341,N_8881,N_8662);
nor U9342 (N_9342,N_8915,N_8295);
xor U9343 (N_9343,N_8351,N_8937);
nand U9344 (N_9344,N_8794,N_8288);
nor U9345 (N_9345,N_8894,N_8979);
and U9346 (N_9346,N_8352,N_8497);
nand U9347 (N_9347,N_8197,N_8631);
and U9348 (N_9348,N_8800,N_8482);
and U9349 (N_9349,N_8705,N_8404);
and U9350 (N_9350,N_8615,N_8409);
nand U9351 (N_9351,N_8522,N_8347);
nor U9352 (N_9352,N_8146,N_8504);
nand U9353 (N_9353,N_8728,N_8278);
nor U9354 (N_9354,N_8137,N_8132);
nand U9355 (N_9355,N_8094,N_8460);
nand U9356 (N_9356,N_8106,N_8168);
or U9357 (N_9357,N_8318,N_8953);
nand U9358 (N_9358,N_8707,N_8298);
and U9359 (N_9359,N_8812,N_8041);
nor U9360 (N_9360,N_8428,N_8191);
xnor U9361 (N_9361,N_8641,N_8681);
or U9362 (N_9362,N_8396,N_8560);
nor U9363 (N_9363,N_8857,N_8138);
nand U9364 (N_9364,N_8443,N_8127);
xor U9365 (N_9365,N_8478,N_8038);
nand U9366 (N_9366,N_8034,N_8277);
and U9367 (N_9367,N_8688,N_8803);
and U9368 (N_9368,N_8991,N_8488);
and U9369 (N_9369,N_8421,N_8493);
or U9370 (N_9370,N_8081,N_8386);
nand U9371 (N_9371,N_8398,N_8051);
xor U9372 (N_9372,N_8962,N_8332);
nand U9373 (N_9373,N_8760,N_8114);
and U9374 (N_9374,N_8552,N_8046);
nand U9375 (N_9375,N_8536,N_8057);
xnor U9376 (N_9376,N_8570,N_8843);
xnor U9377 (N_9377,N_8160,N_8870);
or U9378 (N_9378,N_8060,N_8951);
nand U9379 (N_9379,N_8471,N_8397);
or U9380 (N_9380,N_8257,N_8703);
and U9381 (N_9381,N_8419,N_8944);
nand U9382 (N_9382,N_8783,N_8774);
nor U9383 (N_9383,N_8757,N_8986);
and U9384 (N_9384,N_8939,N_8526);
xor U9385 (N_9385,N_8837,N_8091);
and U9386 (N_9386,N_8899,N_8980);
nand U9387 (N_9387,N_8817,N_8356);
xor U9388 (N_9388,N_8676,N_8280);
nand U9389 (N_9389,N_8743,N_8723);
or U9390 (N_9390,N_8963,N_8224);
nand U9391 (N_9391,N_8650,N_8105);
and U9392 (N_9392,N_8027,N_8165);
or U9393 (N_9393,N_8807,N_8130);
nor U9394 (N_9394,N_8054,N_8290);
xnor U9395 (N_9395,N_8353,N_8301);
nor U9396 (N_9396,N_8503,N_8458);
and U9397 (N_9397,N_8254,N_8946);
nor U9398 (N_9398,N_8835,N_8256);
xnor U9399 (N_9399,N_8285,N_8342);
nor U9400 (N_9400,N_8307,N_8070);
xor U9401 (N_9401,N_8543,N_8625);
nor U9402 (N_9402,N_8215,N_8629);
and U9403 (N_9403,N_8422,N_8623);
or U9404 (N_9404,N_8954,N_8469);
nor U9405 (N_9405,N_8934,N_8373);
or U9406 (N_9406,N_8265,N_8888);
xor U9407 (N_9407,N_8237,N_8430);
nor U9408 (N_9408,N_8627,N_8785);
or U9409 (N_9409,N_8327,N_8814);
nor U9410 (N_9410,N_8903,N_8328);
xor U9411 (N_9411,N_8032,N_8844);
or U9412 (N_9412,N_8415,N_8088);
nand U9413 (N_9413,N_8942,N_8713);
and U9414 (N_9414,N_8651,N_8611);
or U9415 (N_9415,N_8613,N_8544);
xnor U9416 (N_9416,N_8056,N_8389);
nor U9417 (N_9417,N_8198,N_8109);
or U9418 (N_9418,N_8612,N_8213);
or U9419 (N_9419,N_8189,N_8678);
nor U9420 (N_9420,N_8828,N_8736);
or U9421 (N_9421,N_8752,N_8802);
or U9422 (N_9422,N_8699,N_8483);
nand U9423 (N_9423,N_8410,N_8276);
nand U9424 (N_9424,N_8015,N_8362);
and U9425 (N_9425,N_8987,N_8302);
and U9426 (N_9426,N_8745,N_8201);
xor U9427 (N_9427,N_8159,N_8401);
nor U9428 (N_9428,N_8804,N_8518);
nand U9429 (N_9429,N_8371,N_8684);
nand U9430 (N_9430,N_8385,N_8919);
nand U9431 (N_9431,N_8519,N_8499);
xnor U9432 (N_9432,N_8593,N_8820);
and U9433 (N_9433,N_8123,N_8746);
or U9434 (N_9434,N_8701,N_8826);
xnor U9435 (N_9435,N_8622,N_8260);
and U9436 (N_9436,N_8831,N_8671);
and U9437 (N_9437,N_8966,N_8620);
nor U9438 (N_9438,N_8283,N_8456);
nand U9439 (N_9439,N_8636,N_8824);
xor U9440 (N_9440,N_8918,N_8047);
or U9441 (N_9441,N_8581,N_8184);
xor U9442 (N_9442,N_8566,N_8133);
and U9443 (N_9443,N_8722,N_8282);
or U9444 (N_9444,N_8758,N_8645);
xnor U9445 (N_9445,N_8361,N_8126);
nand U9446 (N_9446,N_8468,N_8923);
nor U9447 (N_9447,N_8606,N_8495);
nand U9448 (N_9448,N_8496,N_8013);
and U9449 (N_9449,N_8066,N_8244);
or U9450 (N_9450,N_8753,N_8675);
xor U9451 (N_9451,N_8480,N_8377);
nand U9452 (N_9452,N_8487,N_8376);
or U9453 (N_9453,N_8075,N_8764);
and U9454 (N_9454,N_8542,N_8221);
or U9455 (N_9455,N_8846,N_8656);
xnor U9456 (N_9456,N_8173,N_8299);
xnor U9457 (N_9457,N_8685,N_8022);
or U9458 (N_9458,N_8498,N_8850);
nand U9459 (N_9459,N_8813,N_8876);
and U9460 (N_9460,N_8726,N_8696);
or U9461 (N_9461,N_8240,N_8324);
xnor U9462 (N_9462,N_8556,N_8513);
nor U9463 (N_9463,N_8970,N_8010);
nand U9464 (N_9464,N_8364,N_8214);
and U9465 (N_9465,N_8190,N_8727);
nand U9466 (N_9466,N_8647,N_8775);
or U9467 (N_9467,N_8706,N_8489);
and U9468 (N_9468,N_8071,N_8118);
nor U9469 (N_9469,N_8001,N_8008);
or U9470 (N_9470,N_8885,N_8380);
xnor U9471 (N_9471,N_8801,N_8604);
or U9472 (N_9472,N_8095,N_8532);
and U9473 (N_9473,N_8711,N_8765);
nand U9474 (N_9474,N_8687,N_8584);
or U9475 (N_9475,N_8284,N_8050);
or U9476 (N_9476,N_8117,N_8724);
xnor U9477 (N_9477,N_8908,N_8025);
or U9478 (N_9478,N_8442,N_8369);
nor U9479 (N_9479,N_8883,N_8316);
and U9480 (N_9480,N_8203,N_8698);
xnor U9481 (N_9481,N_8170,N_8122);
nand U9482 (N_9482,N_8538,N_8782);
xnor U9483 (N_9483,N_8550,N_8053);
nor U9484 (N_9484,N_8228,N_8573);
nor U9485 (N_9485,N_8406,N_8860);
or U9486 (N_9486,N_8014,N_8580);
nand U9487 (N_9487,N_8534,N_8607);
or U9488 (N_9488,N_8171,N_8563);
xor U9489 (N_9489,N_8384,N_8602);
and U9490 (N_9490,N_8248,N_8869);
xnor U9491 (N_9491,N_8674,N_8776);
nand U9492 (N_9492,N_8940,N_8562);
nand U9493 (N_9493,N_8906,N_8827);
and U9494 (N_9494,N_8374,N_8941);
nand U9495 (N_9495,N_8077,N_8424);
and U9496 (N_9496,N_8164,N_8399);
xnor U9497 (N_9497,N_8879,N_8714);
and U9498 (N_9498,N_8725,N_8439);
or U9499 (N_9499,N_8466,N_8546);
or U9500 (N_9500,N_8427,N_8608);
or U9501 (N_9501,N_8042,N_8522);
nand U9502 (N_9502,N_8357,N_8041);
nor U9503 (N_9503,N_8778,N_8395);
and U9504 (N_9504,N_8514,N_8887);
xnor U9505 (N_9505,N_8289,N_8688);
or U9506 (N_9506,N_8692,N_8709);
or U9507 (N_9507,N_8972,N_8462);
nand U9508 (N_9508,N_8045,N_8832);
and U9509 (N_9509,N_8306,N_8399);
nand U9510 (N_9510,N_8400,N_8075);
and U9511 (N_9511,N_8548,N_8780);
or U9512 (N_9512,N_8083,N_8685);
or U9513 (N_9513,N_8179,N_8925);
xnor U9514 (N_9514,N_8822,N_8047);
nor U9515 (N_9515,N_8033,N_8078);
and U9516 (N_9516,N_8857,N_8664);
nor U9517 (N_9517,N_8031,N_8668);
nand U9518 (N_9518,N_8255,N_8102);
and U9519 (N_9519,N_8103,N_8452);
nand U9520 (N_9520,N_8866,N_8357);
nor U9521 (N_9521,N_8173,N_8499);
and U9522 (N_9522,N_8007,N_8432);
or U9523 (N_9523,N_8248,N_8901);
xnor U9524 (N_9524,N_8832,N_8528);
or U9525 (N_9525,N_8235,N_8352);
or U9526 (N_9526,N_8605,N_8937);
nand U9527 (N_9527,N_8116,N_8704);
nand U9528 (N_9528,N_8085,N_8285);
xnor U9529 (N_9529,N_8081,N_8314);
nand U9530 (N_9530,N_8840,N_8154);
and U9531 (N_9531,N_8374,N_8618);
nor U9532 (N_9532,N_8536,N_8966);
nand U9533 (N_9533,N_8095,N_8968);
nand U9534 (N_9534,N_8320,N_8776);
nor U9535 (N_9535,N_8910,N_8087);
and U9536 (N_9536,N_8884,N_8554);
or U9537 (N_9537,N_8898,N_8646);
or U9538 (N_9538,N_8871,N_8612);
nor U9539 (N_9539,N_8167,N_8143);
and U9540 (N_9540,N_8001,N_8880);
nand U9541 (N_9541,N_8721,N_8449);
xnor U9542 (N_9542,N_8938,N_8259);
nand U9543 (N_9543,N_8566,N_8783);
nor U9544 (N_9544,N_8798,N_8479);
nor U9545 (N_9545,N_8555,N_8928);
or U9546 (N_9546,N_8917,N_8841);
and U9547 (N_9547,N_8092,N_8395);
or U9548 (N_9548,N_8512,N_8298);
nand U9549 (N_9549,N_8982,N_8966);
nand U9550 (N_9550,N_8992,N_8859);
or U9551 (N_9551,N_8243,N_8167);
or U9552 (N_9552,N_8192,N_8909);
nor U9553 (N_9553,N_8154,N_8831);
or U9554 (N_9554,N_8923,N_8570);
nand U9555 (N_9555,N_8175,N_8289);
or U9556 (N_9556,N_8365,N_8564);
xor U9557 (N_9557,N_8064,N_8154);
xnor U9558 (N_9558,N_8986,N_8917);
or U9559 (N_9559,N_8590,N_8564);
and U9560 (N_9560,N_8850,N_8736);
and U9561 (N_9561,N_8105,N_8925);
nor U9562 (N_9562,N_8258,N_8601);
nor U9563 (N_9563,N_8087,N_8895);
nand U9564 (N_9564,N_8214,N_8183);
nand U9565 (N_9565,N_8884,N_8590);
or U9566 (N_9566,N_8979,N_8348);
and U9567 (N_9567,N_8060,N_8818);
xnor U9568 (N_9568,N_8502,N_8823);
nor U9569 (N_9569,N_8937,N_8544);
or U9570 (N_9570,N_8899,N_8318);
and U9571 (N_9571,N_8651,N_8140);
xnor U9572 (N_9572,N_8379,N_8344);
and U9573 (N_9573,N_8128,N_8275);
or U9574 (N_9574,N_8920,N_8426);
and U9575 (N_9575,N_8207,N_8347);
or U9576 (N_9576,N_8901,N_8562);
or U9577 (N_9577,N_8315,N_8246);
nand U9578 (N_9578,N_8634,N_8024);
nand U9579 (N_9579,N_8255,N_8262);
nand U9580 (N_9580,N_8320,N_8376);
nand U9581 (N_9581,N_8853,N_8483);
and U9582 (N_9582,N_8334,N_8682);
nand U9583 (N_9583,N_8433,N_8255);
and U9584 (N_9584,N_8938,N_8401);
and U9585 (N_9585,N_8807,N_8826);
nor U9586 (N_9586,N_8561,N_8935);
nor U9587 (N_9587,N_8068,N_8767);
nand U9588 (N_9588,N_8195,N_8926);
nor U9589 (N_9589,N_8609,N_8729);
and U9590 (N_9590,N_8827,N_8203);
nor U9591 (N_9591,N_8251,N_8558);
or U9592 (N_9592,N_8353,N_8605);
xor U9593 (N_9593,N_8043,N_8168);
xor U9594 (N_9594,N_8568,N_8917);
nor U9595 (N_9595,N_8285,N_8395);
or U9596 (N_9596,N_8992,N_8936);
and U9597 (N_9597,N_8444,N_8923);
xnor U9598 (N_9598,N_8682,N_8813);
or U9599 (N_9599,N_8147,N_8109);
or U9600 (N_9600,N_8018,N_8803);
xor U9601 (N_9601,N_8444,N_8875);
xnor U9602 (N_9602,N_8006,N_8504);
xor U9603 (N_9603,N_8373,N_8362);
or U9604 (N_9604,N_8943,N_8940);
and U9605 (N_9605,N_8079,N_8706);
or U9606 (N_9606,N_8264,N_8828);
or U9607 (N_9607,N_8702,N_8085);
nor U9608 (N_9608,N_8437,N_8459);
xor U9609 (N_9609,N_8235,N_8415);
or U9610 (N_9610,N_8855,N_8408);
xnor U9611 (N_9611,N_8900,N_8646);
nor U9612 (N_9612,N_8867,N_8282);
or U9613 (N_9613,N_8814,N_8104);
or U9614 (N_9614,N_8869,N_8946);
or U9615 (N_9615,N_8319,N_8054);
nand U9616 (N_9616,N_8723,N_8289);
nor U9617 (N_9617,N_8272,N_8432);
nand U9618 (N_9618,N_8379,N_8703);
or U9619 (N_9619,N_8505,N_8623);
xnor U9620 (N_9620,N_8138,N_8108);
nor U9621 (N_9621,N_8481,N_8473);
nand U9622 (N_9622,N_8054,N_8761);
nor U9623 (N_9623,N_8057,N_8316);
nor U9624 (N_9624,N_8235,N_8735);
nand U9625 (N_9625,N_8360,N_8965);
or U9626 (N_9626,N_8250,N_8780);
xor U9627 (N_9627,N_8311,N_8352);
xor U9628 (N_9628,N_8201,N_8952);
and U9629 (N_9629,N_8092,N_8299);
and U9630 (N_9630,N_8974,N_8742);
and U9631 (N_9631,N_8043,N_8312);
xor U9632 (N_9632,N_8230,N_8305);
or U9633 (N_9633,N_8178,N_8364);
or U9634 (N_9634,N_8491,N_8300);
nor U9635 (N_9635,N_8908,N_8156);
nor U9636 (N_9636,N_8908,N_8416);
and U9637 (N_9637,N_8640,N_8429);
and U9638 (N_9638,N_8082,N_8718);
and U9639 (N_9639,N_8666,N_8294);
xor U9640 (N_9640,N_8769,N_8620);
nor U9641 (N_9641,N_8516,N_8446);
xor U9642 (N_9642,N_8515,N_8332);
or U9643 (N_9643,N_8690,N_8210);
xor U9644 (N_9644,N_8494,N_8436);
or U9645 (N_9645,N_8133,N_8727);
nand U9646 (N_9646,N_8452,N_8338);
and U9647 (N_9647,N_8643,N_8307);
nand U9648 (N_9648,N_8309,N_8217);
xnor U9649 (N_9649,N_8435,N_8708);
nand U9650 (N_9650,N_8053,N_8149);
xor U9651 (N_9651,N_8669,N_8023);
and U9652 (N_9652,N_8563,N_8396);
nor U9653 (N_9653,N_8534,N_8442);
or U9654 (N_9654,N_8798,N_8109);
xnor U9655 (N_9655,N_8292,N_8664);
and U9656 (N_9656,N_8222,N_8763);
nor U9657 (N_9657,N_8367,N_8143);
and U9658 (N_9658,N_8514,N_8977);
nor U9659 (N_9659,N_8897,N_8820);
nor U9660 (N_9660,N_8724,N_8197);
nand U9661 (N_9661,N_8613,N_8169);
nand U9662 (N_9662,N_8944,N_8404);
and U9663 (N_9663,N_8976,N_8709);
nor U9664 (N_9664,N_8529,N_8792);
or U9665 (N_9665,N_8031,N_8117);
or U9666 (N_9666,N_8672,N_8650);
or U9667 (N_9667,N_8215,N_8068);
nor U9668 (N_9668,N_8570,N_8447);
and U9669 (N_9669,N_8349,N_8164);
and U9670 (N_9670,N_8878,N_8324);
xnor U9671 (N_9671,N_8736,N_8915);
and U9672 (N_9672,N_8786,N_8339);
nand U9673 (N_9673,N_8164,N_8291);
xnor U9674 (N_9674,N_8705,N_8988);
nand U9675 (N_9675,N_8474,N_8470);
nand U9676 (N_9676,N_8177,N_8150);
xnor U9677 (N_9677,N_8580,N_8071);
nor U9678 (N_9678,N_8238,N_8347);
or U9679 (N_9679,N_8410,N_8910);
or U9680 (N_9680,N_8275,N_8201);
and U9681 (N_9681,N_8053,N_8922);
xnor U9682 (N_9682,N_8038,N_8618);
and U9683 (N_9683,N_8137,N_8112);
nand U9684 (N_9684,N_8184,N_8443);
or U9685 (N_9685,N_8925,N_8562);
and U9686 (N_9686,N_8147,N_8612);
and U9687 (N_9687,N_8991,N_8076);
and U9688 (N_9688,N_8946,N_8329);
and U9689 (N_9689,N_8420,N_8258);
and U9690 (N_9690,N_8016,N_8212);
and U9691 (N_9691,N_8638,N_8162);
xnor U9692 (N_9692,N_8232,N_8298);
nor U9693 (N_9693,N_8349,N_8793);
xnor U9694 (N_9694,N_8922,N_8137);
xor U9695 (N_9695,N_8451,N_8619);
nor U9696 (N_9696,N_8802,N_8731);
or U9697 (N_9697,N_8771,N_8230);
and U9698 (N_9698,N_8844,N_8370);
nand U9699 (N_9699,N_8290,N_8451);
xnor U9700 (N_9700,N_8985,N_8590);
xor U9701 (N_9701,N_8589,N_8506);
xor U9702 (N_9702,N_8181,N_8871);
or U9703 (N_9703,N_8639,N_8798);
and U9704 (N_9704,N_8497,N_8541);
nor U9705 (N_9705,N_8532,N_8338);
and U9706 (N_9706,N_8850,N_8313);
or U9707 (N_9707,N_8585,N_8838);
xor U9708 (N_9708,N_8173,N_8092);
and U9709 (N_9709,N_8422,N_8350);
and U9710 (N_9710,N_8460,N_8301);
nand U9711 (N_9711,N_8180,N_8589);
nor U9712 (N_9712,N_8619,N_8041);
xnor U9713 (N_9713,N_8707,N_8524);
nor U9714 (N_9714,N_8289,N_8998);
nand U9715 (N_9715,N_8977,N_8923);
nand U9716 (N_9716,N_8462,N_8987);
nor U9717 (N_9717,N_8045,N_8906);
xnor U9718 (N_9718,N_8744,N_8328);
and U9719 (N_9719,N_8097,N_8597);
nand U9720 (N_9720,N_8614,N_8832);
and U9721 (N_9721,N_8376,N_8491);
nand U9722 (N_9722,N_8670,N_8160);
nand U9723 (N_9723,N_8971,N_8654);
nor U9724 (N_9724,N_8714,N_8100);
xor U9725 (N_9725,N_8660,N_8110);
or U9726 (N_9726,N_8063,N_8267);
or U9727 (N_9727,N_8559,N_8321);
nand U9728 (N_9728,N_8764,N_8427);
nor U9729 (N_9729,N_8709,N_8937);
and U9730 (N_9730,N_8263,N_8212);
nor U9731 (N_9731,N_8080,N_8744);
and U9732 (N_9732,N_8813,N_8736);
and U9733 (N_9733,N_8762,N_8322);
and U9734 (N_9734,N_8482,N_8124);
and U9735 (N_9735,N_8503,N_8897);
nor U9736 (N_9736,N_8960,N_8844);
xor U9737 (N_9737,N_8641,N_8376);
nor U9738 (N_9738,N_8569,N_8704);
nor U9739 (N_9739,N_8438,N_8731);
and U9740 (N_9740,N_8268,N_8091);
nand U9741 (N_9741,N_8108,N_8050);
or U9742 (N_9742,N_8209,N_8617);
and U9743 (N_9743,N_8783,N_8961);
or U9744 (N_9744,N_8269,N_8337);
or U9745 (N_9745,N_8433,N_8245);
or U9746 (N_9746,N_8770,N_8476);
nand U9747 (N_9747,N_8633,N_8132);
nand U9748 (N_9748,N_8798,N_8586);
nand U9749 (N_9749,N_8536,N_8457);
xnor U9750 (N_9750,N_8757,N_8714);
or U9751 (N_9751,N_8747,N_8632);
and U9752 (N_9752,N_8575,N_8843);
nor U9753 (N_9753,N_8161,N_8098);
nand U9754 (N_9754,N_8425,N_8555);
nor U9755 (N_9755,N_8855,N_8025);
and U9756 (N_9756,N_8293,N_8945);
xnor U9757 (N_9757,N_8391,N_8553);
xnor U9758 (N_9758,N_8648,N_8545);
xnor U9759 (N_9759,N_8394,N_8027);
or U9760 (N_9760,N_8517,N_8646);
xor U9761 (N_9761,N_8531,N_8600);
and U9762 (N_9762,N_8172,N_8142);
nor U9763 (N_9763,N_8983,N_8018);
or U9764 (N_9764,N_8949,N_8340);
and U9765 (N_9765,N_8865,N_8665);
or U9766 (N_9766,N_8678,N_8463);
and U9767 (N_9767,N_8375,N_8390);
xor U9768 (N_9768,N_8595,N_8337);
nand U9769 (N_9769,N_8165,N_8542);
nand U9770 (N_9770,N_8201,N_8199);
xor U9771 (N_9771,N_8075,N_8984);
and U9772 (N_9772,N_8113,N_8532);
or U9773 (N_9773,N_8529,N_8924);
nor U9774 (N_9774,N_8405,N_8190);
or U9775 (N_9775,N_8070,N_8645);
nor U9776 (N_9776,N_8915,N_8698);
nand U9777 (N_9777,N_8973,N_8553);
and U9778 (N_9778,N_8203,N_8719);
xor U9779 (N_9779,N_8753,N_8917);
and U9780 (N_9780,N_8787,N_8105);
or U9781 (N_9781,N_8782,N_8903);
and U9782 (N_9782,N_8541,N_8008);
nor U9783 (N_9783,N_8219,N_8573);
xnor U9784 (N_9784,N_8527,N_8914);
or U9785 (N_9785,N_8781,N_8800);
xnor U9786 (N_9786,N_8118,N_8846);
nand U9787 (N_9787,N_8514,N_8589);
or U9788 (N_9788,N_8810,N_8230);
or U9789 (N_9789,N_8666,N_8220);
xor U9790 (N_9790,N_8026,N_8839);
and U9791 (N_9791,N_8281,N_8526);
xnor U9792 (N_9792,N_8060,N_8372);
and U9793 (N_9793,N_8025,N_8876);
nand U9794 (N_9794,N_8962,N_8997);
and U9795 (N_9795,N_8897,N_8808);
or U9796 (N_9796,N_8673,N_8378);
or U9797 (N_9797,N_8858,N_8846);
nor U9798 (N_9798,N_8953,N_8425);
nand U9799 (N_9799,N_8507,N_8551);
and U9800 (N_9800,N_8858,N_8617);
nand U9801 (N_9801,N_8919,N_8461);
nand U9802 (N_9802,N_8062,N_8657);
xor U9803 (N_9803,N_8763,N_8501);
xor U9804 (N_9804,N_8018,N_8386);
nand U9805 (N_9805,N_8629,N_8143);
nor U9806 (N_9806,N_8328,N_8782);
nand U9807 (N_9807,N_8820,N_8296);
or U9808 (N_9808,N_8550,N_8207);
or U9809 (N_9809,N_8457,N_8733);
nand U9810 (N_9810,N_8137,N_8927);
xor U9811 (N_9811,N_8117,N_8910);
or U9812 (N_9812,N_8722,N_8728);
xor U9813 (N_9813,N_8511,N_8527);
and U9814 (N_9814,N_8722,N_8276);
or U9815 (N_9815,N_8679,N_8209);
nand U9816 (N_9816,N_8736,N_8866);
nor U9817 (N_9817,N_8305,N_8899);
and U9818 (N_9818,N_8572,N_8782);
or U9819 (N_9819,N_8012,N_8617);
nor U9820 (N_9820,N_8935,N_8459);
nor U9821 (N_9821,N_8715,N_8944);
xnor U9822 (N_9822,N_8407,N_8013);
nand U9823 (N_9823,N_8142,N_8916);
xor U9824 (N_9824,N_8800,N_8034);
and U9825 (N_9825,N_8225,N_8806);
or U9826 (N_9826,N_8955,N_8722);
nand U9827 (N_9827,N_8756,N_8520);
and U9828 (N_9828,N_8699,N_8421);
and U9829 (N_9829,N_8107,N_8070);
xnor U9830 (N_9830,N_8074,N_8014);
or U9831 (N_9831,N_8071,N_8005);
nor U9832 (N_9832,N_8595,N_8827);
xnor U9833 (N_9833,N_8745,N_8360);
nand U9834 (N_9834,N_8544,N_8612);
xor U9835 (N_9835,N_8037,N_8557);
nand U9836 (N_9836,N_8534,N_8830);
nand U9837 (N_9837,N_8845,N_8434);
and U9838 (N_9838,N_8944,N_8175);
xnor U9839 (N_9839,N_8189,N_8519);
xnor U9840 (N_9840,N_8507,N_8618);
nor U9841 (N_9841,N_8597,N_8819);
xor U9842 (N_9842,N_8418,N_8783);
xnor U9843 (N_9843,N_8070,N_8050);
or U9844 (N_9844,N_8823,N_8335);
nand U9845 (N_9845,N_8989,N_8664);
and U9846 (N_9846,N_8677,N_8743);
nand U9847 (N_9847,N_8527,N_8313);
nor U9848 (N_9848,N_8913,N_8298);
xor U9849 (N_9849,N_8428,N_8348);
or U9850 (N_9850,N_8508,N_8752);
xor U9851 (N_9851,N_8705,N_8780);
nor U9852 (N_9852,N_8683,N_8638);
xor U9853 (N_9853,N_8778,N_8316);
xor U9854 (N_9854,N_8054,N_8715);
nor U9855 (N_9855,N_8663,N_8487);
and U9856 (N_9856,N_8354,N_8002);
nor U9857 (N_9857,N_8608,N_8422);
nor U9858 (N_9858,N_8747,N_8160);
nand U9859 (N_9859,N_8153,N_8211);
xnor U9860 (N_9860,N_8177,N_8113);
or U9861 (N_9861,N_8497,N_8672);
or U9862 (N_9862,N_8427,N_8220);
xnor U9863 (N_9863,N_8169,N_8028);
or U9864 (N_9864,N_8955,N_8643);
nand U9865 (N_9865,N_8253,N_8904);
nor U9866 (N_9866,N_8575,N_8933);
nand U9867 (N_9867,N_8626,N_8341);
xnor U9868 (N_9868,N_8990,N_8340);
nand U9869 (N_9869,N_8700,N_8226);
xnor U9870 (N_9870,N_8507,N_8142);
nand U9871 (N_9871,N_8146,N_8300);
or U9872 (N_9872,N_8204,N_8702);
nand U9873 (N_9873,N_8348,N_8476);
and U9874 (N_9874,N_8410,N_8533);
nor U9875 (N_9875,N_8830,N_8068);
xnor U9876 (N_9876,N_8645,N_8513);
xor U9877 (N_9877,N_8974,N_8042);
nand U9878 (N_9878,N_8027,N_8535);
nand U9879 (N_9879,N_8200,N_8203);
and U9880 (N_9880,N_8376,N_8646);
nand U9881 (N_9881,N_8770,N_8396);
or U9882 (N_9882,N_8356,N_8357);
nand U9883 (N_9883,N_8404,N_8784);
nand U9884 (N_9884,N_8862,N_8156);
or U9885 (N_9885,N_8172,N_8357);
xnor U9886 (N_9886,N_8494,N_8988);
nor U9887 (N_9887,N_8402,N_8471);
nand U9888 (N_9888,N_8109,N_8695);
nor U9889 (N_9889,N_8674,N_8077);
nand U9890 (N_9890,N_8190,N_8373);
nor U9891 (N_9891,N_8483,N_8705);
xor U9892 (N_9892,N_8945,N_8205);
nand U9893 (N_9893,N_8422,N_8156);
xnor U9894 (N_9894,N_8417,N_8359);
and U9895 (N_9895,N_8672,N_8009);
nor U9896 (N_9896,N_8914,N_8067);
nand U9897 (N_9897,N_8916,N_8099);
or U9898 (N_9898,N_8373,N_8133);
and U9899 (N_9899,N_8644,N_8308);
and U9900 (N_9900,N_8001,N_8840);
nor U9901 (N_9901,N_8599,N_8498);
nand U9902 (N_9902,N_8626,N_8706);
nand U9903 (N_9903,N_8846,N_8370);
or U9904 (N_9904,N_8586,N_8112);
and U9905 (N_9905,N_8589,N_8298);
and U9906 (N_9906,N_8013,N_8079);
or U9907 (N_9907,N_8156,N_8875);
or U9908 (N_9908,N_8575,N_8358);
nand U9909 (N_9909,N_8686,N_8520);
xnor U9910 (N_9910,N_8031,N_8378);
xnor U9911 (N_9911,N_8999,N_8242);
nand U9912 (N_9912,N_8482,N_8012);
nor U9913 (N_9913,N_8673,N_8747);
xnor U9914 (N_9914,N_8701,N_8024);
nor U9915 (N_9915,N_8398,N_8659);
xnor U9916 (N_9916,N_8464,N_8942);
xor U9917 (N_9917,N_8800,N_8278);
nand U9918 (N_9918,N_8940,N_8082);
or U9919 (N_9919,N_8690,N_8591);
nor U9920 (N_9920,N_8035,N_8730);
xnor U9921 (N_9921,N_8563,N_8179);
nand U9922 (N_9922,N_8712,N_8885);
or U9923 (N_9923,N_8387,N_8879);
and U9924 (N_9924,N_8167,N_8165);
or U9925 (N_9925,N_8495,N_8569);
nand U9926 (N_9926,N_8389,N_8270);
nand U9927 (N_9927,N_8686,N_8750);
nand U9928 (N_9928,N_8457,N_8128);
or U9929 (N_9929,N_8495,N_8492);
nor U9930 (N_9930,N_8942,N_8683);
or U9931 (N_9931,N_8721,N_8911);
nor U9932 (N_9932,N_8581,N_8505);
nand U9933 (N_9933,N_8591,N_8400);
nand U9934 (N_9934,N_8122,N_8459);
nand U9935 (N_9935,N_8744,N_8460);
xnor U9936 (N_9936,N_8159,N_8730);
nor U9937 (N_9937,N_8469,N_8412);
xor U9938 (N_9938,N_8359,N_8396);
xor U9939 (N_9939,N_8024,N_8303);
and U9940 (N_9940,N_8774,N_8925);
or U9941 (N_9941,N_8837,N_8802);
nand U9942 (N_9942,N_8767,N_8988);
or U9943 (N_9943,N_8855,N_8574);
or U9944 (N_9944,N_8890,N_8648);
or U9945 (N_9945,N_8067,N_8635);
nand U9946 (N_9946,N_8232,N_8624);
or U9947 (N_9947,N_8020,N_8113);
and U9948 (N_9948,N_8991,N_8112);
nand U9949 (N_9949,N_8817,N_8537);
and U9950 (N_9950,N_8282,N_8726);
and U9951 (N_9951,N_8468,N_8734);
nand U9952 (N_9952,N_8649,N_8681);
xnor U9953 (N_9953,N_8730,N_8853);
or U9954 (N_9954,N_8002,N_8249);
and U9955 (N_9955,N_8089,N_8113);
nor U9956 (N_9956,N_8752,N_8575);
nand U9957 (N_9957,N_8065,N_8165);
nor U9958 (N_9958,N_8998,N_8910);
or U9959 (N_9959,N_8821,N_8262);
or U9960 (N_9960,N_8037,N_8969);
or U9961 (N_9961,N_8037,N_8267);
or U9962 (N_9962,N_8631,N_8047);
nand U9963 (N_9963,N_8979,N_8372);
nor U9964 (N_9964,N_8583,N_8793);
nor U9965 (N_9965,N_8844,N_8616);
xor U9966 (N_9966,N_8462,N_8297);
nor U9967 (N_9967,N_8041,N_8241);
nor U9968 (N_9968,N_8822,N_8572);
nand U9969 (N_9969,N_8678,N_8697);
or U9970 (N_9970,N_8860,N_8876);
or U9971 (N_9971,N_8680,N_8242);
xnor U9972 (N_9972,N_8578,N_8627);
or U9973 (N_9973,N_8817,N_8564);
and U9974 (N_9974,N_8163,N_8914);
and U9975 (N_9975,N_8833,N_8974);
nor U9976 (N_9976,N_8137,N_8492);
nor U9977 (N_9977,N_8259,N_8189);
or U9978 (N_9978,N_8226,N_8880);
nor U9979 (N_9979,N_8294,N_8958);
and U9980 (N_9980,N_8236,N_8349);
or U9981 (N_9981,N_8486,N_8431);
and U9982 (N_9982,N_8851,N_8059);
and U9983 (N_9983,N_8807,N_8264);
nand U9984 (N_9984,N_8631,N_8950);
or U9985 (N_9985,N_8315,N_8277);
nor U9986 (N_9986,N_8846,N_8263);
nand U9987 (N_9987,N_8304,N_8722);
and U9988 (N_9988,N_8464,N_8412);
xor U9989 (N_9989,N_8408,N_8415);
nor U9990 (N_9990,N_8414,N_8696);
or U9991 (N_9991,N_8399,N_8257);
nor U9992 (N_9992,N_8101,N_8508);
nand U9993 (N_9993,N_8663,N_8740);
and U9994 (N_9994,N_8924,N_8242);
or U9995 (N_9995,N_8974,N_8989);
nand U9996 (N_9996,N_8621,N_8075);
and U9997 (N_9997,N_8386,N_8759);
xor U9998 (N_9998,N_8142,N_8098);
nand U9999 (N_9999,N_8293,N_8960);
nand U10000 (N_10000,N_9646,N_9807);
nand U10001 (N_10001,N_9344,N_9564);
xor U10002 (N_10002,N_9282,N_9215);
or U10003 (N_10003,N_9079,N_9500);
xor U10004 (N_10004,N_9896,N_9303);
xor U10005 (N_10005,N_9703,N_9680);
and U10006 (N_10006,N_9613,N_9793);
and U10007 (N_10007,N_9112,N_9236);
and U10008 (N_10008,N_9558,N_9374);
xnor U10009 (N_10009,N_9962,N_9573);
and U10010 (N_10010,N_9822,N_9651);
or U10011 (N_10011,N_9944,N_9032);
or U10012 (N_10012,N_9562,N_9679);
or U10013 (N_10013,N_9263,N_9586);
nor U10014 (N_10014,N_9144,N_9729);
nor U10015 (N_10015,N_9191,N_9714);
xor U10016 (N_10016,N_9231,N_9183);
nand U10017 (N_10017,N_9991,N_9406);
xor U10018 (N_10018,N_9290,N_9918);
nor U10019 (N_10019,N_9635,N_9375);
nand U10020 (N_10020,N_9545,N_9170);
nand U10021 (N_10021,N_9181,N_9435);
nand U10022 (N_10022,N_9213,N_9849);
xor U10023 (N_10023,N_9972,N_9983);
or U10024 (N_10024,N_9782,N_9491);
xnor U10025 (N_10025,N_9077,N_9682);
or U10026 (N_10026,N_9838,N_9654);
and U10027 (N_10027,N_9411,N_9018);
xnor U10028 (N_10028,N_9168,N_9592);
or U10029 (N_10029,N_9625,N_9865);
or U10030 (N_10030,N_9088,N_9816);
xnor U10031 (N_10031,N_9949,N_9410);
nand U10032 (N_10032,N_9866,N_9605);
or U10033 (N_10033,N_9804,N_9467);
xor U10034 (N_10034,N_9463,N_9421);
and U10035 (N_10035,N_9489,N_9315);
or U10036 (N_10036,N_9953,N_9081);
nor U10037 (N_10037,N_9888,N_9496);
and U10038 (N_10038,N_9292,N_9832);
or U10039 (N_10039,N_9709,N_9102);
and U10040 (N_10040,N_9200,N_9905);
nor U10041 (N_10041,N_9770,N_9967);
nor U10042 (N_10042,N_9204,N_9543);
xnor U10043 (N_10043,N_9890,N_9920);
xor U10044 (N_10044,N_9990,N_9055);
nor U10045 (N_10045,N_9726,N_9644);
xor U10046 (N_10046,N_9945,N_9935);
nor U10047 (N_10047,N_9692,N_9280);
nor U10048 (N_10048,N_9356,N_9447);
or U10049 (N_10049,N_9606,N_9764);
xor U10050 (N_10050,N_9187,N_9777);
xor U10051 (N_10051,N_9350,N_9796);
and U10052 (N_10052,N_9567,N_9520);
or U10053 (N_10053,N_9129,N_9359);
xnor U10054 (N_10054,N_9425,N_9718);
nor U10055 (N_10055,N_9169,N_9085);
nand U10056 (N_10056,N_9330,N_9148);
nand U10057 (N_10057,N_9874,N_9391);
nor U10058 (N_10058,N_9660,N_9551);
or U10059 (N_10059,N_9759,N_9221);
nor U10060 (N_10060,N_9050,N_9255);
nand U10061 (N_10061,N_9639,N_9994);
or U10062 (N_10062,N_9369,N_9891);
xor U10063 (N_10063,N_9041,N_9474);
xor U10064 (N_10064,N_9408,N_9560);
or U10065 (N_10065,N_9647,N_9358);
xnor U10066 (N_10066,N_9960,N_9700);
or U10067 (N_10067,N_9048,N_9748);
nand U10068 (N_10068,N_9033,N_9017);
or U10069 (N_10069,N_9532,N_9583);
xor U10070 (N_10070,N_9951,N_9071);
nor U10071 (N_10071,N_9593,N_9347);
nand U10072 (N_10072,N_9548,N_9024);
nor U10073 (N_10073,N_9863,N_9514);
nor U10074 (N_10074,N_9284,N_9407);
or U10075 (N_10075,N_9109,N_9602);
and U10076 (N_10076,N_9300,N_9878);
nor U10077 (N_10077,N_9192,N_9083);
xor U10078 (N_10078,N_9604,N_9846);
and U10079 (N_10079,N_9264,N_9328);
nor U10080 (N_10080,N_9368,N_9027);
or U10081 (N_10081,N_9853,N_9964);
nor U10082 (N_10082,N_9513,N_9941);
xnor U10083 (N_10083,N_9008,N_9094);
and U10084 (N_10084,N_9788,N_9022);
xor U10085 (N_10085,N_9295,N_9565);
and U10086 (N_10086,N_9974,N_9291);
xnor U10087 (N_10087,N_9011,N_9332);
nor U10088 (N_10088,N_9707,N_9780);
nor U10089 (N_10089,N_9909,N_9057);
nor U10090 (N_10090,N_9663,N_9334);
or U10091 (N_10091,N_9245,N_9981);
nand U10092 (N_10092,N_9355,N_9069);
nor U10093 (N_10093,N_9582,N_9311);
xnor U10094 (N_10094,N_9076,N_9308);
nor U10095 (N_10095,N_9727,N_9519);
and U10096 (N_10096,N_9855,N_9000);
xor U10097 (N_10097,N_9823,N_9986);
or U10098 (N_10098,N_9938,N_9847);
nand U10099 (N_10099,N_9133,N_9082);
and U10100 (N_10100,N_9667,N_9320);
nand U10101 (N_10101,N_9572,N_9090);
or U10102 (N_10102,N_9120,N_9316);
nand U10103 (N_10103,N_9268,N_9304);
nand U10104 (N_10104,N_9526,N_9252);
xor U10105 (N_10105,N_9488,N_9220);
nor U10106 (N_10106,N_9237,N_9821);
nor U10107 (N_10107,N_9553,N_9769);
nor U10108 (N_10108,N_9314,N_9508);
or U10109 (N_10109,N_9060,N_9697);
or U10110 (N_10110,N_9756,N_9059);
xor U10111 (N_10111,N_9190,N_9323);
nor U10112 (N_10112,N_9546,N_9193);
or U10113 (N_10113,N_9498,N_9265);
or U10114 (N_10114,N_9261,N_9418);
or U10115 (N_10115,N_9121,N_9705);
and U10116 (N_10116,N_9720,N_9885);
nor U10117 (N_10117,N_9776,N_9899);
xor U10118 (N_10118,N_9742,N_9465);
xnor U10119 (N_10119,N_9023,N_9266);
nor U10120 (N_10120,N_9642,N_9256);
nand U10121 (N_10121,N_9157,N_9063);
or U10122 (N_10122,N_9638,N_9387);
and U10123 (N_10123,N_9214,N_9341);
or U10124 (N_10124,N_9445,N_9458);
or U10125 (N_10125,N_9078,N_9342);
and U10126 (N_10126,N_9665,N_9515);
xor U10127 (N_10127,N_9829,N_9814);
or U10128 (N_10128,N_9616,N_9812);
and U10129 (N_10129,N_9750,N_9650);
and U10130 (N_10130,N_9373,N_9395);
or U10131 (N_10131,N_9414,N_9452);
xnor U10132 (N_10132,N_9149,N_9158);
and U10133 (N_10133,N_9980,N_9224);
or U10134 (N_10134,N_9774,N_9331);
nand U10135 (N_10135,N_9004,N_9757);
xnor U10136 (N_10136,N_9744,N_9765);
xor U10137 (N_10137,N_9862,N_9724);
or U10138 (N_10138,N_9946,N_9108);
and U10139 (N_10139,N_9669,N_9441);
or U10140 (N_10140,N_9629,N_9758);
nor U10141 (N_10141,N_9695,N_9906);
or U10142 (N_10142,N_9730,N_9423);
nand U10143 (N_10143,N_9791,N_9424);
xnor U10144 (N_10144,N_9831,N_9449);
or U10145 (N_10145,N_9388,N_9633);
and U10146 (N_10146,N_9529,N_9167);
nor U10147 (N_10147,N_9509,N_9523);
or U10148 (N_10148,N_9539,N_9163);
or U10149 (N_10149,N_9596,N_9417);
or U10150 (N_10150,N_9688,N_9289);
or U10151 (N_10151,N_9074,N_9335);
or U10152 (N_10152,N_9656,N_9916);
or U10153 (N_10153,N_9184,N_9015);
nor U10154 (N_10154,N_9099,N_9666);
xor U10155 (N_10155,N_9794,N_9195);
or U10156 (N_10156,N_9338,N_9239);
and U10157 (N_10157,N_9883,N_9908);
xor U10158 (N_10158,N_9851,N_9670);
xor U10159 (N_10159,N_9913,N_9249);
nand U10160 (N_10160,N_9615,N_9684);
nand U10161 (N_10161,N_9432,N_9399);
or U10162 (N_10162,N_9881,N_9557);
and U10163 (N_10163,N_9456,N_9766);
or U10164 (N_10164,N_9106,N_9242);
nor U10165 (N_10165,N_9232,N_9171);
nand U10166 (N_10166,N_9732,N_9608);
or U10167 (N_10167,N_9741,N_9947);
nor U10168 (N_10168,N_9547,N_9678);
and U10169 (N_10169,N_9747,N_9911);
or U10170 (N_10170,N_9603,N_9561);
and U10171 (N_10171,N_9366,N_9227);
and U10172 (N_10172,N_9536,N_9578);
and U10173 (N_10173,N_9258,N_9113);
xnor U10174 (N_10174,N_9609,N_9333);
nor U10175 (N_10175,N_9510,N_9965);
xor U10176 (N_10176,N_9858,N_9226);
nor U10177 (N_10177,N_9689,N_9749);
or U10178 (N_10178,N_9324,N_9844);
nand U10179 (N_10179,N_9124,N_9092);
nand U10180 (N_10180,N_9542,N_9143);
xor U10181 (N_10181,N_9156,N_9497);
nand U10182 (N_10182,N_9571,N_9882);
and U10183 (N_10183,N_9690,N_9437);
nand U10184 (N_10184,N_9999,N_9351);
nand U10185 (N_10185,N_9468,N_9626);
nand U10186 (N_10186,N_9979,N_9618);
or U10187 (N_10187,N_9172,N_9492);
xnor U10188 (N_10188,N_9243,N_9940);
nand U10189 (N_10189,N_9767,N_9118);
or U10190 (N_10190,N_9820,N_9025);
or U10191 (N_10191,N_9957,N_9763);
or U10192 (N_10192,N_9378,N_9202);
nor U10193 (N_10193,N_9924,N_9969);
or U10194 (N_10194,N_9073,N_9768);
nand U10195 (N_10195,N_9131,N_9146);
nor U10196 (N_10196,N_9904,N_9459);
and U10197 (N_10197,N_9309,N_9483);
nor U10198 (N_10198,N_9661,N_9577);
xnor U10199 (N_10199,N_9599,N_9716);
and U10200 (N_10200,N_9907,N_9065);
or U10201 (N_10201,N_9563,N_9628);
nand U10202 (N_10202,N_9939,N_9702);
xor U10203 (N_10203,N_9222,N_9783);
and U10204 (N_10204,N_9116,N_9089);
and U10205 (N_10205,N_9559,N_9385);
nand U10206 (N_10206,N_9096,N_9062);
nand U10207 (N_10207,N_9588,N_9932);
and U10208 (N_10208,N_9275,N_9186);
nor U10209 (N_10209,N_9166,N_9481);
xnor U10210 (N_10210,N_9367,N_9868);
nor U10211 (N_10211,N_9589,N_9634);
xnor U10212 (N_10212,N_9693,N_9495);
xor U10213 (N_10213,N_9860,N_9310);
nor U10214 (N_10214,N_9686,N_9180);
or U10215 (N_10215,N_9100,N_9648);
nand U10216 (N_10216,N_9627,N_9392);
and U10217 (N_10217,N_9987,N_9789);
xnor U10218 (N_10218,N_9067,N_9360);
xor U10219 (N_10219,N_9594,N_9030);
and U10220 (N_10220,N_9451,N_9457);
nor U10221 (N_10221,N_9105,N_9054);
xor U10222 (N_10222,N_9218,N_9929);
or U10223 (N_10223,N_9824,N_9499);
and U10224 (N_10224,N_9552,N_9927);
nor U10225 (N_10225,N_9046,N_9098);
or U10226 (N_10226,N_9671,N_9349);
nand U10227 (N_10227,N_9438,N_9401);
xnor U10228 (N_10228,N_9995,N_9029);
xor U10229 (N_10229,N_9296,N_9541);
nand U10230 (N_10230,N_9294,N_9655);
or U10231 (N_10231,N_9436,N_9028);
xor U10232 (N_10232,N_9659,N_9569);
xnor U10233 (N_10233,N_9576,N_9760);
and U10234 (N_10234,N_9892,N_9478);
xnor U10235 (N_10235,N_9472,N_9313);
xor U10236 (N_10236,N_9502,N_9982);
or U10237 (N_10237,N_9177,N_9450);
and U10238 (N_10238,N_9856,N_9630);
xnor U10239 (N_10239,N_9959,N_9555);
or U10240 (N_10240,N_9731,N_9601);
and U10241 (N_10241,N_9412,N_9792);
and U10242 (N_10242,N_9127,N_9955);
or U10243 (N_10243,N_9128,N_9640);
and U10244 (N_10244,N_9002,N_9799);
nor U10245 (N_10245,N_9694,N_9574);
and U10246 (N_10246,N_9696,N_9404);
nand U10247 (N_10247,N_9591,N_9476);
or U10248 (N_10248,N_9598,N_9524);
xor U10249 (N_10249,N_9234,N_9636);
xnor U10250 (N_10250,N_9318,N_9466);
nor U10251 (N_10251,N_9016,N_9993);
nor U10252 (N_10252,N_9042,N_9197);
nand U10253 (N_10253,N_9762,N_9135);
nand U10254 (N_10254,N_9403,N_9897);
nor U10255 (N_10255,N_9830,N_9400);
nor U10256 (N_10256,N_9097,N_9178);
or U10257 (N_10257,N_9317,N_9056);
nor U10258 (N_10258,N_9440,N_9117);
and U10259 (N_10259,N_9841,N_9875);
nand U10260 (N_10260,N_9611,N_9525);
nor U10261 (N_10261,N_9087,N_9337);
xnor U10262 (N_10262,N_9738,N_9068);
and U10263 (N_10263,N_9619,N_9066);
or U10264 (N_10264,N_9867,N_9988);
nand U10265 (N_10265,N_9754,N_9072);
nand U10266 (N_10266,N_9211,N_9001);
nand U10267 (N_10267,N_9162,N_9464);
and U10268 (N_10268,N_9173,N_9610);
or U10269 (N_10269,N_9138,N_9958);
xor U10270 (N_10270,N_9871,N_9902);
nor U10271 (N_10271,N_9251,N_9479);
nand U10272 (N_10272,N_9322,N_9299);
nand U10273 (N_10273,N_9521,N_9685);
nand U10274 (N_10274,N_9722,N_9036);
and U10275 (N_10275,N_9926,N_9522);
nor U10276 (N_10276,N_9683,N_9165);
and U10277 (N_10277,N_9119,N_9394);
and U10278 (N_10278,N_9454,N_9198);
or U10279 (N_10279,N_9475,N_9708);
nor U10280 (N_10280,N_9880,N_9954);
and U10281 (N_10281,N_9486,N_9271);
or U10282 (N_10282,N_9091,N_9934);
and U10283 (N_10283,N_9922,N_9809);
nor U10284 (N_10284,N_9267,N_9274);
xnor U10285 (N_10285,N_9687,N_9409);
nand U10286 (N_10286,N_9053,N_9453);
nand U10287 (N_10287,N_9061,N_9019);
and U10288 (N_10288,N_9051,N_9527);
or U10289 (N_10289,N_9533,N_9182);
xor U10290 (N_10290,N_9781,N_9710);
nor U10291 (N_10291,N_9327,N_9740);
xnor U10292 (N_10292,N_9728,N_9364);
xor U10293 (N_10293,N_9413,N_9370);
nor U10294 (N_10294,N_9624,N_9006);
nor U10295 (N_10295,N_9622,N_9446);
nand U10296 (N_10296,N_9581,N_9674);
xor U10297 (N_10297,N_9223,N_9806);
and U10298 (N_10298,N_9086,N_9701);
or U10299 (N_10299,N_9269,N_9787);
or U10300 (N_10300,N_9746,N_9970);
and U10301 (N_10301,N_9971,N_9857);
nand U10302 (N_10302,N_9039,N_9383);
xnor U10303 (N_10303,N_9281,N_9339);
nand U10304 (N_10304,N_9805,N_9933);
nor U10305 (N_10305,N_9925,N_9978);
nor U10306 (N_10306,N_9530,N_9228);
nand U10307 (N_10307,N_9931,N_9672);
nor U10308 (N_10308,N_9270,N_9745);
xnor U10309 (N_10309,N_9505,N_9026);
or U10310 (N_10310,N_9321,N_9325);
and U10311 (N_10311,N_9996,N_9817);
xnor U10312 (N_10312,N_9645,N_9312);
nand U10313 (N_10313,N_9715,N_9595);
and U10314 (N_10314,N_9235,N_9159);
nor U10315 (N_10315,N_9216,N_9164);
nor U10316 (N_10316,N_9285,N_9585);
or U10317 (N_10317,N_9699,N_9879);
xnor U10318 (N_10318,N_9047,N_9556);
nor U10319 (N_10319,N_9772,N_9021);
and U10320 (N_10320,N_9590,N_9713);
and U10321 (N_10321,N_9652,N_9307);
xnor U10322 (N_10322,N_9207,N_9405);
nor U10323 (N_10323,N_9176,N_9203);
nor U10324 (N_10324,N_9393,N_9554);
or U10325 (N_10325,N_9043,N_9901);
nor U10326 (N_10326,N_9210,N_9676);
and U10327 (N_10327,N_9535,N_9379);
and U10328 (N_10328,N_9910,N_9504);
xor U10329 (N_10329,N_9151,N_9653);
nand U10330 (N_10330,N_9123,N_9587);
and U10331 (N_10331,N_9319,N_9431);
nor U10332 (N_10332,N_9798,N_9376);
xor U10333 (N_10333,N_9381,N_9487);
nand U10334 (N_10334,N_9196,N_9761);
nand U10335 (N_10335,N_9735,N_9390);
and U10336 (N_10336,N_9775,N_9637);
nand U10337 (N_10337,N_9473,N_9260);
nand U10338 (N_10338,N_9828,N_9386);
and U10339 (N_10339,N_9607,N_9305);
or U10340 (N_10340,N_9448,N_9973);
nor U10341 (N_10341,N_9900,N_9155);
nand U10342 (N_10342,N_9247,N_9273);
nor U10343 (N_10343,N_9471,N_9912);
nand U10344 (N_10344,N_9442,N_9826);
nand U10345 (N_10345,N_9430,N_9272);
or U10346 (N_10346,N_9943,N_9600);
and U10347 (N_10347,N_9717,N_9737);
xnor U10348 (N_10348,N_9175,N_9219);
and U10349 (N_10349,N_9597,N_9813);
xnor U10350 (N_10350,N_9836,N_9711);
xor U10351 (N_10351,N_9917,N_9877);
nor U10352 (N_10352,N_9540,N_9005);
or U10353 (N_10353,N_9632,N_9125);
nand U10354 (N_10354,N_9104,N_9889);
nor U10355 (N_10355,N_9070,N_9064);
xnor U10356 (N_10356,N_9840,N_9518);
or U10357 (N_10357,N_9095,N_9107);
xor U10358 (N_10358,N_9803,N_9287);
and U10359 (N_10359,N_9614,N_9278);
and U10360 (N_10360,N_9426,N_9101);
or U10361 (N_10361,N_9340,N_9254);
nor U10362 (N_10362,N_9966,N_9968);
xor U10363 (N_10363,N_9205,N_9773);
nand U10364 (N_10364,N_9516,N_9277);
xor U10365 (N_10365,N_9537,N_9549);
nor U10366 (N_10366,N_9049,N_9903);
nand U10367 (N_10367,N_9253,N_9733);
nor U10368 (N_10368,N_9462,N_9930);
nor U10369 (N_10369,N_9725,N_9801);
nand U10370 (N_10370,N_9003,N_9677);
or U10371 (N_10371,N_9861,N_9736);
nand U10372 (N_10372,N_9887,N_9876);
or U10373 (N_10373,N_9810,N_9503);
or U10374 (N_10374,N_9045,N_9914);
xnor U10375 (N_10375,N_9477,N_9415);
nor U10376 (N_10376,N_9839,N_9326);
nor U10377 (N_10377,N_9837,N_9185);
nand U10378 (N_10378,N_9869,N_9461);
xor U10379 (N_10379,N_9921,N_9818);
xor U10380 (N_10380,N_9052,N_9229);
or U10381 (N_10381,N_9977,N_9819);
nor U10382 (N_10382,N_9361,N_9825);
xnor U10383 (N_10383,N_9579,N_9115);
nor U10384 (N_10384,N_9620,N_9649);
nor U10385 (N_10385,N_9298,N_9217);
and U10386 (N_10386,N_9140,N_9194);
nor U10387 (N_10387,N_9136,N_9811);
nand U10388 (N_10388,N_9534,N_9485);
or U10389 (N_10389,N_9575,N_9110);
xor U10390 (N_10390,N_9434,N_9852);
nor U10391 (N_10391,N_9712,N_9948);
nor U10392 (N_10392,N_9942,N_9544);
nand U10393 (N_10393,N_9833,N_9150);
and U10394 (N_10394,N_9528,N_9126);
xnor U10395 (N_10395,N_9363,N_9035);
nand U10396 (N_10396,N_9835,N_9842);
nand U10397 (N_10397,N_9362,N_9283);
or U10398 (N_10398,N_9698,N_9402);
xor U10399 (N_10399,N_9240,N_9631);
nand U10400 (N_10400,N_9241,N_9512);
nand U10401 (N_10401,N_9179,N_9511);
nor U10402 (N_10402,N_9797,N_9779);
or U10403 (N_10403,N_9137,N_9134);
and U10404 (N_10404,N_9785,N_9984);
and U10405 (N_10405,N_9482,N_9377);
nand U10406 (N_10406,N_9201,N_9854);
nand U10407 (N_10407,N_9443,N_9668);
nor U10408 (N_10408,N_9188,N_9494);
xnor U10409 (N_10409,N_9859,N_9427);
or U10410 (N_10410,N_9800,N_9952);
xor U10411 (N_10411,N_9936,N_9790);
nand U10412 (N_10412,N_9416,N_9623);
xnor U10413 (N_10413,N_9673,N_9306);
nor U10414 (N_10414,N_9843,N_9989);
and U10415 (N_10415,N_9396,N_9531);
or U10416 (N_10416,N_9225,N_9484);
nor U10417 (N_10417,N_9570,N_9233);
nand U10418 (N_10418,N_9297,N_9132);
xor U10419 (N_10419,N_9238,N_9915);
nor U10420 (N_10420,N_9020,N_9354);
nand U10421 (N_10421,N_9142,N_9657);
nand U10422 (N_10422,N_9230,N_9075);
and U10423 (N_10423,N_9139,N_9044);
and U10424 (N_10424,N_9460,N_9037);
xor U10425 (N_10425,N_9444,N_9428);
xnor U10426 (N_10426,N_9345,N_9658);
nor U10427 (N_10427,N_9568,N_9739);
or U10428 (N_10428,N_9147,N_9898);
nor U10429 (N_10429,N_9886,N_9084);
nand U10430 (N_10430,N_9009,N_9808);
and U10431 (N_10431,N_9279,N_9919);
xnor U10432 (N_10432,N_9013,N_9894);
xor U10433 (N_10433,N_9950,N_9584);
and U10434 (N_10434,N_9493,N_9038);
or U10435 (N_10435,N_9975,N_9439);
nand U10436 (N_10436,N_9870,N_9161);
xor U10437 (N_10437,N_9336,N_9751);
xor U10438 (N_10438,N_9681,N_9371);
nand U10439 (N_10439,N_9506,N_9276);
nand U10440 (N_10440,N_9103,N_9145);
or U10441 (N_10441,N_9997,N_9470);
nand U10442 (N_10442,N_9058,N_9617);
nand U10443 (N_10443,N_9286,N_9641);
and U10444 (N_10444,N_9937,N_9141);
or U10445 (N_10445,N_9093,N_9420);
xor U10446 (N_10446,N_9998,N_9248);
and U10447 (N_10447,N_9014,N_9834);
or U10448 (N_10448,N_9827,N_9246);
xor U10449 (N_10449,N_9154,N_9455);
xor U10450 (N_10450,N_9398,N_9382);
xor U10451 (N_10451,N_9538,N_9963);
nand U10452 (N_10452,N_9786,N_9244);
xnor U10453 (N_10453,N_9872,N_9643);
and U10454 (N_10454,N_9348,N_9153);
and U10455 (N_10455,N_9288,N_9490);
nand U10456 (N_10456,N_9753,N_9864);
nor U10457 (N_10457,N_9419,N_9357);
nor U10458 (N_10458,N_9734,N_9704);
xor U10459 (N_10459,N_9721,N_9848);
and U10460 (N_10460,N_9985,N_9329);
xnor U10461 (N_10461,N_9302,N_9114);
and U10462 (N_10462,N_9884,N_9422);
nor U10463 (N_10463,N_9259,N_9893);
xnor U10464 (N_10464,N_9480,N_9353);
nor U10465 (N_10465,N_9621,N_9691);
and U10466 (N_10466,N_9152,N_9992);
and U10467 (N_10467,N_9080,N_9293);
nor U10468 (N_10468,N_9815,N_9384);
or U10469 (N_10469,N_9845,N_9160);
nor U10470 (N_10470,N_9778,N_9010);
or U10471 (N_10471,N_9743,N_9873);
xnor U10472 (N_10472,N_9566,N_9664);
xnor U10473 (N_10473,N_9365,N_9397);
or U10474 (N_10474,N_9612,N_9928);
and U10475 (N_10475,N_9262,N_9372);
and U10476 (N_10476,N_9034,N_9675);
nor U10477 (N_10477,N_9122,N_9209);
and U10478 (N_10478,N_9040,N_9189);
xnor U10479 (N_10479,N_9517,N_9802);
and U10480 (N_10480,N_9662,N_9343);
nand U10481 (N_10481,N_9352,N_9433);
nor U10482 (N_10482,N_9550,N_9795);
xnor U10483 (N_10483,N_9752,N_9007);
nor U10484 (N_10484,N_9206,N_9755);
or U10485 (N_10485,N_9130,N_9212);
nand U10486 (N_10486,N_9895,N_9784);
and U10487 (N_10487,N_9961,N_9301);
nand U10488 (N_10488,N_9257,N_9956);
nor U10489 (N_10489,N_9111,N_9719);
and U10490 (N_10490,N_9923,N_9346);
and U10491 (N_10491,N_9250,N_9771);
or U10492 (N_10492,N_9706,N_9976);
xor U10493 (N_10493,N_9031,N_9850);
nor U10494 (N_10494,N_9507,N_9469);
and U10495 (N_10495,N_9174,N_9580);
nand U10496 (N_10496,N_9208,N_9012);
and U10497 (N_10497,N_9501,N_9380);
or U10498 (N_10498,N_9199,N_9429);
or U10499 (N_10499,N_9389,N_9723);
or U10500 (N_10500,N_9417,N_9102);
nand U10501 (N_10501,N_9327,N_9714);
nand U10502 (N_10502,N_9632,N_9651);
or U10503 (N_10503,N_9829,N_9344);
xnor U10504 (N_10504,N_9783,N_9724);
nor U10505 (N_10505,N_9618,N_9063);
and U10506 (N_10506,N_9306,N_9807);
and U10507 (N_10507,N_9086,N_9829);
xnor U10508 (N_10508,N_9074,N_9055);
nor U10509 (N_10509,N_9128,N_9969);
or U10510 (N_10510,N_9356,N_9588);
nand U10511 (N_10511,N_9892,N_9064);
or U10512 (N_10512,N_9487,N_9393);
xnor U10513 (N_10513,N_9267,N_9452);
and U10514 (N_10514,N_9045,N_9227);
xor U10515 (N_10515,N_9979,N_9765);
and U10516 (N_10516,N_9177,N_9857);
xor U10517 (N_10517,N_9450,N_9503);
or U10518 (N_10518,N_9528,N_9584);
xor U10519 (N_10519,N_9690,N_9538);
xnor U10520 (N_10520,N_9438,N_9945);
xnor U10521 (N_10521,N_9853,N_9351);
xnor U10522 (N_10522,N_9360,N_9309);
nand U10523 (N_10523,N_9690,N_9796);
and U10524 (N_10524,N_9904,N_9450);
nor U10525 (N_10525,N_9038,N_9043);
or U10526 (N_10526,N_9174,N_9648);
or U10527 (N_10527,N_9231,N_9277);
xnor U10528 (N_10528,N_9624,N_9807);
nand U10529 (N_10529,N_9049,N_9584);
or U10530 (N_10530,N_9382,N_9262);
nor U10531 (N_10531,N_9202,N_9098);
or U10532 (N_10532,N_9167,N_9624);
nor U10533 (N_10533,N_9746,N_9229);
xor U10534 (N_10534,N_9058,N_9424);
or U10535 (N_10535,N_9422,N_9309);
nor U10536 (N_10536,N_9650,N_9134);
and U10537 (N_10537,N_9862,N_9036);
and U10538 (N_10538,N_9036,N_9951);
nor U10539 (N_10539,N_9499,N_9603);
or U10540 (N_10540,N_9132,N_9325);
nor U10541 (N_10541,N_9521,N_9812);
xnor U10542 (N_10542,N_9380,N_9506);
or U10543 (N_10543,N_9191,N_9056);
nand U10544 (N_10544,N_9399,N_9614);
nand U10545 (N_10545,N_9246,N_9665);
xor U10546 (N_10546,N_9463,N_9418);
xnor U10547 (N_10547,N_9812,N_9121);
nor U10548 (N_10548,N_9057,N_9300);
nor U10549 (N_10549,N_9302,N_9605);
and U10550 (N_10550,N_9197,N_9032);
xor U10551 (N_10551,N_9723,N_9495);
or U10552 (N_10552,N_9814,N_9994);
or U10553 (N_10553,N_9655,N_9272);
or U10554 (N_10554,N_9524,N_9148);
or U10555 (N_10555,N_9876,N_9927);
and U10556 (N_10556,N_9244,N_9258);
or U10557 (N_10557,N_9247,N_9042);
nor U10558 (N_10558,N_9782,N_9389);
or U10559 (N_10559,N_9611,N_9012);
nor U10560 (N_10560,N_9047,N_9743);
xor U10561 (N_10561,N_9331,N_9798);
xnor U10562 (N_10562,N_9529,N_9719);
or U10563 (N_10563,N_9756,N_9298);
xnor U10564 (N_10564,N_9298,N_9728);
or U10565 (N_10565,N_9878,N_9170);
nand U10566 (N_10566,N_9323,N_9157);
or U10567 (N_10567,N_9499,N_9596);
and U10568 (N_10568,N_9649,N_9460);
xor U10569 (N_10569,N_9304,N_9218);
xnor U10570 (N_10570,N_9248,N_9391);
or U10571 (N_10571,N_9602,N_9553);
xnor U10572 (N_10572,N_9626,N_9874);
nand U10573 (N_10573,N_9413,N_9674);
xnor U10574 (N_10574,N_9995,N_9862);
and U10575 (N_10575,N_9282,N_9408);
nor U10576 (N_10576,N_9829,N_9992);
nand U10577 (N_10577,N_9703,N_9141);
nand U10578 (N_10578,N_9899,N_9038);
nand U10579 (N_10579,N_9127,N_9549);
xor U10580 (N_10580,N_9319,N_9564);
and U10581 (N_10581,N_9297,N_9521);
xor U10582 (N_10582,N_9988,N_9490);
xor U10583 (N_10583,N_9024,N_9105);
and U10584 (N_10584,N_9340,N_9578);
nand U10585 (N_10585,N_9493,N_9587);
or U10586 (N_10586,N_9518,N_9236);
nand U10587 (N_10587,N_9805,N_9744);
or U10588 (N_10588,N_9706,N_9175);
or U10589 (N_10589,N_9437,N_9675);
and U10590 (N_10590,N_9233,N_9810);
nand U10591 (N_10591,N_9007,N_9524);
or U10592 (N_10592,N_9203,N_9107);
and U10593 (N_10593,N_9172,N_9668);
nor U10594 (N_10594,N_9221,N_9888);
nand U10595 (N_10595,N_9067,N_9703);
or U10596 (N_10596,N_9014,N_9040);
xor U10597 (N_10597,N_9001,N_9174);
nand U10598 (N_10598,N_9699,N_9906);
nand U10599 (N_10599,N_9255,N_9302);
nor U10600 (N_10600,N_9442,N_9767);
nor U10601 (N_10601,N_9121,N_9106);
xor U10602 (N_10602,N_9127,N_9045);
and U10603 (N_10603,N_9070,N_9804);
nor U10604 (N_10604,N_9061,N_9860);
and U10605 (N_10605,N_9936,N_9199);
or U10606 (N_10606,N_9410,N_9486);
nand U10607 (N_10607,N_9171,N_9383);
or U10608 (N_10608,N_9013,N_9483);
nor U10609 (N_10609,N_9203,N_9782);
or U10610 (N_10610,N_9181,N_9532);
and U10611 (N_10611,N_9912,N_9035);
xor U10612 (N_10612,N_9149,N_9585);
or U10613 (N_10613,N_9101,N_9114);
xor U10614 (N_10614,N_9215,N_9430);
or U10615 (N_10615,N_9056,N_9732);
xnor U10616 (N_10616,N_9353,N_9915);
nor U10617 (N_10617,N_9936,N_9461);
and U10618 (N_10618,N_9190,N_9317);
nor U10619 (N_10619,N_9104,N_9903);
nor U10620 (N_10620,N_9122,N_9070);
and U10621 (N_10621,N_9226,N_9774);
nand U10622 (N_10622,N_9632,N_9748);
and U10623 (N_10623,N_9303,N_9788);
and U10624 (N_10624,N_9621,N_9792);
or U10625 (N_10625,N_9645,N_9977);
nor U10626 (N_10626,N_9174,N_9481);
xor U10627 (N_10627,N_9386,N_9757);
xor U10628 (N_10628,N_9700,N_9808);
nor U10629 (N_10629,N_9497,N_9762);
xor U10630 (N_10630,N_9614,N_9974);
xor U10631 (N_10631,N_9455,N_9941);
nor U10632 (N_10632,N_9084,N_9616);
nand U10633 (N_10633,N_9462,N_9583);
and U10634 (N_10634,N_9300,N_9354);
xor U10635 (N_10635,N_9608,N_9024);
or U10636 (N_10636,N_9969,N_9387);
nand U10637 (N_10637,N_9487,N_9311);
and U10638 (N_10638,N_9237,N_9348);
and U10639 (N_10639,N_9515,N_9643);
and U10640 (N_10640,N_9891,N_9355);
nor U10641 (N_10641,N_9227,N_9148);
and U10642 (N_10642,N_9646,N_9094);
xnor U10643 (N_10643,N_9020,N_9837);
nand U10644 (N_10644,N_9693,N_9157);
or U10645 (N_10645,N_9151,N_9563);
nand U10646 (N_10646,N_9701,N_9259);
nor U10647 (N_10647,N_9107,N_9506);
xnor U10648 (N_10648,N_9575,N_9605);
xnor U10649 (N_10649,N_9051,N_9726);
nand U10650 (N_10650,N_9342,N_9412);
nor U10651 (N_10651,N_9203,N_9091);
and U10652 (N_10652,N_9886,N_9960);
xor U10653 (N_10653,N_9434,N_9794);
xor U10654 (N_10654,N_9825,N_9226);
and U10655 (N_10655,N_9970,N_9198);
and U10656 (N_10656,N_9110,N_9178);
nor U10657 (N_10657,N_9252,N_9197);
and U10658 (N_10658,N_9755,N_9380);
or U10659 (N_10659,N_9881,N_9874);
nor U10660 (N_10660,N_9326,N_9149);
nor U10661 (N_10661,N_9548,N_9385);
nor U10662 (N_10662,N_9569,N_9425);
or U10663 (N_10663,N_9707,N_9367);
nand U10664 (N_10664,N_9579,N_9027);
or U10665 (N_10665,N_9923,N_9653);
nand U10666 (N_10666,N_9388,N_9279);
nor U10667 (N_10667,N_9544,N_9766);
xnor U10668 (N_10668,N_9215,N_9507);
and U10669 (N_10669,N_9849,N_9781);
nand U10670 (N_10670,N_9092,N_9057);
and U10671 (N_10671,N_9945,N_9884);
nand U10672 (N_10672,N_9011,N_9743);
xor U10673 (N_10673,N_9253,N_9001);
xnor U10674 (N_10674,N_9836,N_9237);
xor U10675 (N_10675,N_9872,N_9867);
nand U10676 (N_10676,N_9681,N_9020);
nand U10677 (N_10677,N_9610,N_9424);
or U10678 (N_10678,N_9729,N_9940);
nand U10679 (N_10679,N_9958,N_9501);
nor U10680 (N_10680,N_9035,N_9127);
nand U10681 (N_10681,N_9617,N_9915);
xor U10682 (N_10682,N_9921,N_9032);
xor U10683 (N_10683,N_9627,N_9343);
xnor U10684 (N_10684,N_9307,N_9989);
nand U10685 (N_10685,N_9965,N_9162);
and U10686 (N_10686,N_9868,N_9885);
or U10687 (N_10687,N_9488,N_9674);
and U10688 (N_10688,N_9609,N_9497);
nand U10689 (N_10689,N_9556,N_9371);
xnor U10690 (N_10690,N_9048,N_9040);
xnor U10691 (N_10691,N_9711,N_9555);
nand U10692 (N_10692,N_9270,N_9110);
and U10693 (N_10693,N_9467,N_9922);
and U10694 (N_10694,N_9496,N_9265);
nor U10695 (N_10695,N_9399,N_9993);
nand U10696 (N_10696,N_9098,N_9078);
nand U10697 (N_10697,N_9718,N_9115);
and U10698 (N_10698,N_9364,N_9273);
xor U10699 (N_10699,N_9079,N_9067);
xnor U10700 (N_10700,N_9734,N_9377);
nand U10701 (N_10701,N_9754,N_9958);
or U10702 (N_10702,N_9531,N_9110);
nand U10703 (N_10703,N_9576,N_9732);
xnor U10704 (N_10704,N_9009,N_9221);
nand U10705 (N_10705,N_9199,N_9298);
nand U10706 (N_10706,N_9297,N_9985);
or U10707 (N_10707,N_9982,N_9730);
or U10708 (N_10708,N_9286,N_9102);
xnor U10709 (N_10709,N_9450,N_9905);
nand U10710 (N_10710,N_9775,N_9328);
xnor U10711 (N_10711,N_9627,N_9933);
xor U10712 (N_10712,N_9510,N_9533);
nor U10713 (N_10713,N_9094,N_9201);
or U10714 (N_10714,N_9752,N_9385);
nand U10715 (N_10715,N_9690,N_9294);
and U10716 (N_10716,N_9768,N_9845);
nor U10717 (N_10717,N_9409,N_9566);
xor U10718 (N_10718,N_9793,N_9338);
or U10719 (N_10719,N_9517,N_9413);
nand U10720 (N_10720,N_9549,N_9228);
xnor U10721 (N_10721,N_9254,N_9324);
nor U10722 (N_10722,N_9548,N_9677);
or U10723 (N_10723,N_9767,N_9235);
xnor U10724 (N_10724,N_9368,N_9221);
nor U10725 (N_10725,N_9082,N_9267);
and U10726 (N_10726,N_9580,N_9162);
nand U10727 (N_10727,N_9124,N_9823);
nand U10728 (N_10728,N_9321,N_9097);
xnor U10729 (N_10729,N_9197,N_9810);
or U10730 (N_10730,N_9908,N_9532);
and U10731 (N_10731,N_9604,N_9751);
or U10732 (N_10732,N_9761,N_9639);
or U10733 (N_10733,N_9420,N_9692);
xnor U10734 (N_10734,N_9967,N_9813);
or U10735 (N_10735,N_9185,N_9317);
xor U10736 (N_10736,N_9172,N_9763);
nor U10737 (N_10737,N_9566,N_9013);
and U10738 (N_10738,N_9373,N_9790);
or U10739 (N_10739,N_9625,N_9845);
nand U10740 (N_10740,N_9113,N_9927);
and U10741 (N_10741,N_9454,N_9666);
xnor U10742 (N_10742,N_9738,N_9648);
and U10743 (N_10743,N_9695,N_9374);
or U10744 (N_10744,N_9207,N_9631);
nor U10745 (N_10745,N_9684,N_9777);
and U10746 (N_10746,N_9236,N_9874);
and U10747 (N_10747,N_9994,N_9002);
and U10748 (N_10748,N_9525,N_9549);
xnor U10749 (N_10749,N_9485,N_9748);
or U10750 (N_10750,N_9997,N_9394);
xor U10751 (N_10751,N_9001,N_9267);
xnor U10752 (N_10752,N_9379,N_9216);
or U10753 (N_10753,N_9323,N_9116);
and U10754 (N_10754,N_9138,N_9313);
and U10755 (N_10755,N_9699,N_9799);
xor U10756 (N_10756,N_9352,N_9967);
or U10757 (N_10757,N_9038,N_9655);
xor U10758 (N_10758,N_9336,N_9815);
nor U10759 (N_10759,N_9320,N_9576);
nand U10760 (N_10760,N_9051,N_9848);
and U10761 (N_10761,N_9069,N_9755);
nand U10762 (N_10762,N_9398,N_9191);
xor U10763 (N_10763,N_9609,N_9094);
nand U10764 (N_10764,N_9677,N_9543);
nor U10765 (N_10765,N_9433,N_9519);
or U10766 (N_10766,N_9433,N_9096);
xnor U10767 (N_10767,N_9733,N_9070);
or U10768 (N_10768,N_9830,N_9808);
and U10769 (N_10769,N_9829,N_9105);
or U10770 (N_10770,N_9741,N_9300);
xor U10771 (N_10771,N_9887,N_9967);
xor U10772 (N_10772,N_9411,N_9040);
or U10773 (N_10773,N_9168,N_9327);
or U10774 (N_10774,N_9283,N_9215);
nor U10775 (N_10775,N_9478,N_9151);
nor U10776 (N_10776,N_9183,N_9948);
xor U10777 (N_10777,N_9872,N_9333);
and U10778 (N_10778,N_9076,N_9560);
nand U10779 (N_10779,N_9033,N_9311);
and U10780 (N_10780,N_9833,N_9199);
nor U10781 (N_10781,N_9587,N_9786);
or U10782 (N_10782,N_9705,N_9134);
xnor U10783 (N_10783,N_9968,N_9144);
nand U10784 (N_10784,N_9884,N_9358);
and U10785 (N_10785,N_9027,N_9040);
xor U10786 (N_10786,N_9804,N_9150);
xnor U10787 (N_10787,N_9912,N_9301);
xnor U10788 (N_10788,N_9853,N_9383);
nor U10789 (N_10789,N_9638,N_9407);
or U10790 (N_10790,N_9676,N_9059);
or U10791 (N_10791,N_9120,N_9713);
xor U10792 (N_10792,N_9293,N_9956);
or U10793 (N_10793,N_9357,N_9751);
and U10794 (N_10794,N_9163,N_9150);
xnor U10795 (N_10795,N_9201,N_9952);
nand U10796 (N_10796,N_9153,N_9076);
nor U10797 (N_10797,N_9600,N_9489);
and U10798 (N_10798,N_9569,N_9760);
nor U10799 (N_10799,N_9449,N_9462);
or U10800 (N_10800,N_9462,N_9962);
and U10801 (N_10801,N_9540,N_9901);
or U10802 (N_10802,N_9509,N_9793);
nand U10803 (N_10803,N_9330,N_9940);
xnor U10804 (N_10804,N_9478,N_9931);
and U10805 (N_10805,N_9425,N_9964);
nor U10806 (N_10806,N_9589,N_9256);
nand U10807 (N_10807,N_9675,N_9964);
and U10808 (N_10808,N_9834,N_9303);
or U10809 (N_10809,N_9699,N_9574);
nand U10810 (N_10810,N_9433,N_9467);
or U10811 (N_10811,N_9625,N_9136);
or U10812 (N_10812,N_9287,N_9277);
or U10813 (N_10813,N_9514,N_9755);
nand U10814 (N_10814,N_9275,N_9195);
xnor U10815 (N_10815,N_9856,N_9108);
and U10816 (N_10816,N_9443,N_9724);
or U10817 (N_10817,N_9600,N_9840);
and U10818 (N_10818,N_9931,N_9791);
and U10819 (N_10819,N_9186,N_9939);
nand U10820 (N_10820,N_9245,N_9219);
or U10821 (N_10821,N_9661,N_9608);
nor U10822 (N_10822,N_9247,N_9737);
nor U10823 (N_10823,N_9007,N_9221);
or U10824 (N_10824,N_9936,N_9131);
xor U10825 (N_10825,N_9234,N_9892);
nand U10826 (N_10826,N_9416,N_9574);
nor U10827 (N_10827,N_9225,N_9964);
xnor U10828 (N_10828,N_9640,N_9257);
xor U10829 (N_10829,N_9306,N_9933);
nand U10830 (N_10830,N_9748,N_9976);
and U10831 (N_10831,N_9561,N_9140);
or U10832 (N_10832,N_9487,N_9728);
and U10833 (N_10833,N_9286,N_9937);
nor U10834 (N_10834,N_9296,N_9830);
nor U10835 (N_10835,N_9779,N_9869);
or U10836 (N_10836,N_9853,N_9214);
nor U10837 (N_10837,N_9735,N_9268);
or U10838 (N_10838,N_9917,N_9210);
or U10839 (N_10839,N_9675,N_9905);
and U10840 (N_10840,N_9073,N_9924);
nor U10841 (N_10841,N_9560,N_9184);
and U10842 (N_10842,N_9179,N_9967);
nand U10843 (N_10843,N_9450,N_9388);
nor U10844 (N_10844,N_9462,N_9133);
xor U10845 (N_10845,N_9822,N_9968);
nor U10846 (N_10846,N_9425,N_9292);
or U10847 (N_10847,N_9623,N_9597);
and U10848 (N_10848,N_9201,N_9203);
or U10849 (N_10849,N_9648,N_9792);
nand U10850 (N_10850,N_9811,N_9698);
or U10851 (N_10851,N_9951,N_9642);
xnor U10852 (N_10852,N_9193,N_9845);
or U10853 (N_10853,N_9251,N_9112);
nand U10854 (N_10854,N_9981,N_9165);
nand U10855 (N_10855,N_9293,N_9738);
and U10856 (N_10856,N_9082,N_9278);
nand U10857 (N_10857,N_9576,N_9175);
or U10858 (N_10858,N_9815,N_9978);
nand U10859 (N_10859,N_9364,N_9470);
xor U10860 (N_10860,N_9655,N_9118);
xnor U10861 (N_10861,N_9466,N_9424);
and U10862 (N_10862,N_9589,N_9798);
nor U10863 (N_10863,N_9150,N_9281);
or U10864 (N_10864,N_9589,N_9543);
nand U10865 (N_10865,N_9245,N_9976);
nand U10866 (N_10866,N_9056,N_9720);
nand U10867 (N_10867,N_9513,N_9731);
xor U10868 (N_10868,N_9796,N_9457);
or U10869 (N_10869,N_9072,N_9230);
and U10870 (N_10870,N_9095,N_9710);
and U10871 (N_10871,N_9569,N_9829);
xnor U10872 (N_10872,N_9103,N_9244);
and U10873 (N_10873,N_9198,N_9665);
and U10874 (N_10874,N_9611,N_9756);
nor U10875 (N_10875,N_9543,N_9839);
and U10876 (N_10876,N_9073,N_9199);
and U10877 (N_10877,N_9975,N_9769);
and U10878 (N_10878,N_9062,N_9064);
nand U10879 (N_10879,N_9335,N_9788);
nand U10880 (N_10880,N_9517,N_9023);
or U10881 (N_10881,N_9753,N_9212);
xor U10882 (N_10882,N_9480,N_9157);
or U10883 (N_10883,N_9033,N_9014);
or U10884 (N_10884,N_9963,N_9434);
nand U10885 (N_10885,N_9625,N_9262);
nor U10886 (N_10886,N_9419,N_9491);
or U10887 (N_10887,N_9798,N_9512);
xnor U10888 (N_10888,N_9147,N_9139);
xnor U10889 (N_10889,N_9755,N_9608);
nand U10890 (N_10890,N_9587,N_9863);
xor U10891 (N_10891,N_9628,N_9456);
nand U10892 (N_10892,N_9499,N_9094);
and U10893 (N_10893,N_9357,N_9471);
and U10894 (N_10894,N_9034,N_9266);
nand U10895 (N_10895,N_9582,N_9401);
nand U10896 (N_10896,N_9254,N_9148);
nand U10897 (N_10897,N_9736,N_9123);
and U10898 (N_10898,N_9176,N_9632);
and U10899 (N_10899,N_9292,N_9766);
nand U10900 (N_10900,N_9434,N_9609);
xnor U10901 (N_10901,N_9472,N_9246);
nor U10902 (N_10902,N_9134,N_9057);
nor U10903 (N_10903,N_9247,N_9016);
or U10904 (N_10904,N_9184,N_9391);
and U10905 (N_10905,N_9493,N_9459);
and U10906 (N_10906,N_9110,N_9698);
nand U10907 (N_10907,N_9314,N_9244);
nand U10908 (N_10908,N_9822,N_9914);
nor U10909 (N_10909,N_9185,N_9157);
or U10910 (N_10910,N_9475,N_9526);
and U10911 (N_10911,N_9413,N_9341);
or U10912 (N_10912,N_9238,N_9257);
and U10913 (N_10913,N_9247,N_9219);
xor U10914 (N_10914,N_9712,N_9717);
or U10915 (N_10915,N_9470,N_9457);
xnor U10916 (N_10916,N_9554,N_9071);
or U10917 (N_10917,N_9061,N_9752);
nor U10918 (N_10918,N_9754,N_9105);
xnor U10919 (N_10919,N_9697,N_9290);
nor U10920 (N_10920,N_9197,N_9825);
nand U10921 (N_10921,N_9019,N_9832);
and U10922 (N_10922,N_9527,N_9286);
nand U10923 (N_10923,N_9931,N_9611);
and U10924 (N_10924,N_9059,N_9615);
or U10925 (N_10925,N_9372,N_9830);
nand U10926 (N_10926,N_9970,N_9234);
nor U10927 (N_10927,N_9756,N_9837);
or U10928 (N_10928,N_9519,N_9021);
xnor U10929 (N_10929,N_9931,N_9318);
nand U10930 (N_10930,N_9534,N_9203);
nor U10931 (N_10931,N_9820,N_9127);
nor U10932 (N_10932,N_9228,N_9781);
and U10933 (N_10933,N_9503,N_9250);
or U10934 (N_10934,N_9276,N_9024);
nor U10935 (N_10935,N_9796,N_9738);
or U10936 (N_10936,N_9565,N_9073);
nand U10937 (N_10937,N_9944,N_9840);
nand U10938 (N_10938,N_9060,N_9679);
and U10939 (N_10939,N_9732,N_9684);
and U10940 (N_10940,N_9066,N_9749);
nor U10941 (N_10941,N_9040,N_9993);
or U10942 (N_10942,N_9042,N_9048);
or U10943 (N_10943,N_9842,N_9841);
and U10944 (N_10944,N_9035,N_9174);
nor U10945 (N_10945,N_9456,N_9144);
nor U10946 (N_10946,N_9336,N_9419);
nand U10947 (N_10947,N_9266,N_9482);
nand U10948 (N_10948,N_9260,N_9638);
nor U10949 (N_10949,N_9018,N_9945);
xor U10950 (N_10950,N_9918,N_9993);
nand U10951 (N_10951,N_9725,N_9852);
nor U10952 (N_10952,N_9252,N_9453);
nand U10953 (N_10953,N_9583,N_9610);
xor U10954 (N_10954,N_9248,N_9476);
nand U10955 (N_10955,N_9818,N_9363);
xnor U10956 (N_10956,N_9590,N_9642);
or U10957 (N_10957,N_9536,N_9716);
and U10958 (N_10958,N_9489,N_9612);
nor U10959 (N_10959,N_9399,N_9599);
nor U10960 (N_10960,N_9484,N_9183);
or U10961 (N_10961,N_9042,N_9995);
nand U10962 (N_10962,N_9405,N_9055);
and U10963 (N_10963,N_9354,N_9924);
and U10964 (N_10964,N_9362,N_9196);
and U10965 (N_10965,N_9322,N_9780);
xor U10966 (N_10966,N_9680,N_9544);
xnor U10967 (N_10967,N_9603,N_9766);
nor U10968 (N_10968,N_9703,N_9321);
xor U10969 (N_10969,N_9096,N_9353);
nor U10970 (N_10970,N_9531,N_9357);
nand U10971 (N_10971,N_9662,N_9358);
nor U10972 (N_10972,N_9791,N_9667);
xnor U10973 (N_10973,N_9204,N_9753);
xor U10974 (N_10974,N_9998,N_9974);
and U10975 (N_10975,N_9231,N_9591);
nand U10976 (N_10976,N_9188,N_9502);
xnor U10977 (N_10977,N_9003,N_9379);
or U10978 (N_10978,N_9900,N_9651);
nor U10979 (N_10979,N_9863,N_9890);
nor U10980 (N_10980,N_9428,N_9767);
and U10981 (N_10981,N_9100,N_9375);
nand U10982 (N_10982,N_9260,N_9529);
nor U10983 (N_10983,N_9713,N_9325);
and U10984 (N_10984,N_9203,N_9348);
and U10985 (N_10985,N_9454,N_9121);
xor U10986 (N_10986,N_9429,N_9788);
nand U10987 (N_10987,N_9723,N_9290);
nor U10988 (N_10988,N_9308,N_9441);
nand U10989 (N_10989,N_9240,N_9270);
nand U10990 (N_10990,N_9630,N_9270);
xnor U10991 (N_10991,N_9093,N_9673);
and U10992 (N_10992,N_9162,N_9560);
nor U10993 (N_10993,N_9846,N_9607);
nor U10994 (N_10994,N_9305,N_9956);
or U10995 (N_10995,N_9735,N_9677);
nand U10996 (N_10996,N_9494,N_9176);
xnor U10997 (N_10997,N_9555,N_9726);
and U10998 (N_10998,N_9495,N_9751);
nand U10999 (N_10999,N_9353,N_9294);
or U11000 (N_11000,N_10843,N_10164);
nand U11001 (N_11001,N_10799,N_10154);
nand U11002 (N_11002,N_10294,N_10071);
xor U11003 (N_11003,N_10900,N_10017);
nand U11004 (N_11004,N_10642,N_10142);
nand U11005 (N_11005,N_10611,N_10863);
or U11006 (N_11006,N_10834,N_10997);
or U11007 (N_11007,N_10480,N_10203);
or U11008 (N_11008,N_10947,N_10449);
or U11009 (N_11009,N_10955,N_10521);
or U11010 (N_11010,N_10807,N_10297);
or U11011 (N_11011,N_10924,N_10332);
xnor U11012 (N_11012,N_10585,N_10308);
and U11013 (N_11013,N_10353,N_10706);
xor U11014 (N_11014,N_10695,N_10437);
or U11015 (N_11015,N_10571,N_10870);
and U11016 (N_11016,N_10321,N_10392);
nand U11017 (N_11017,N_10043,N_10214);
or U11018 (N_11018,N_10994,N_10599);
nor U11019 (N_11019,N_10177,N_10737);
xnor U11020 (N_11020,N_10731,N_10016);
and U11021 (N_11021,N_10696,N_10701);
or U11022 (N_11022,N_10830,N_10772);
nand U11023 (N_11023,N_10451,N_10476);
or U11024 (N_11024,N_10271,N_10378);
or U11025 (N_11025,N_10121,N_10605);
nor U11026 (N_11026,N_10042,N_10583);
nor U11027 (N_11027,N_10926,N_10036);
or U11028 (N_11028,N_10816,N_10329);
or U11029 (N_11029,N_10064,N_10893);
xor U11030 (N_11030,N_10335,N_10769);
xor U11031 (N_11031,N_10953,N_10151);
and U11032 (N_11032,N_10587,N_10442);
nand U11033 (N_11033,N_10986,N_10676);
xor U11034 (N_11034,N_10768,N_10199);
xor U11035 (N_11035,N_10699,N_10651);
and U11036 (N_11036,N_10591,N_10938);
nor U11037 (N_11037,N_10349,N_10508);
or U11038 (N_11038,N_10977,N_10812);
xnor U11039 (N_11039,N_10631,N_10312);
and U11040 (N_11040,N_10359,N_10922);
and U11041 (N_11041,N_10111,N_10311);
and U11042 (N_11042,N_10325,N_10894);
xor U11043 (N_11043,N_10813,N_10336);
xor U11044 (N_11044,N_10510,N_10837);
nand U11045 (N_11045,N_10693,N_10190);
and U11046 (N_11046,N_10298,N_10879);
or U11047 (N_11047,N_10009,N_10469);
or U11048 (N_11048,N_10103,N_10943);
nand U11049 (N_11049,N_10512,N_10310);
and U11050 (N_11050,N_10145,N_10345);
and U11051 (N_11051,N_10160,N_10999);
and U11052 (N_11052,N_10233,N_10193);
xnor U11053 (N_11053,N_10805,N_10496);
xor U11054 (N_11054,N_10598,N_10020);
xor U11055 (N_11055,N_10270,N_10448);
nand U11056 (N_11056,N_10109,N_10840);
nor U11057 (N_11057,N_10369,N_10169);
xnor U11058 (N_11058,N_10608,N_10101);
nand U11059 (N_11059,N_10096,N_10950);
and U11060 (N_11060,N_10860,N_10523);
xor U11061 (N_11061,N_10562,N_10283);
nand U11062 (N_11062,N_10492,N_10134);
nor U11063 (N_11063,N_10590,N_10739);
nand U11064 (N_11064,N_10440,N_10291);
nor U11065 (N_11065,N_10525,N_10722);
nor U11066 (N_11066,N_10761,N_10129);
or U11067 (N_11067,N_10886,N_10005);
nor U11068 (N_11068,N_10856,N_10973);
nor U11069 (N_11069,N_10342,N_10880);
nor U11070 (N_11070,N_10896,N_10023);
and U11071 (N_11071,N_10503,N_10954);
or U11072 (N_11072,N_10668,N_10589);
and U11073 (N_11073,N_10721,N_10106);
nor U11074 (N_11074,N_10213,N_10466);
nor U11075 (N_11075,N_10839,N_10889);
and U11076 (N_11076,N_10531,N_10912);
nand U11077 (N_11077,N_10559,N_10010);
xor U11078 (N_11078,N_10427,N_10343);
nor U11079 (N_11079,N_10965,N_10753);
nand U11080 (N_11080,N_10018,N_10666);
nor U11081 (N_11081,N_10268,N_10906);
and U11082 (N_11082,N_10654,N_10350);
and U11083 (N_11083,N_10620,N_10781);
nand U11084 (N_11084,N_10675,N_10618);
and U11085 (N_11085,N_10218,N_10749);
and U11086 (N_11086,N_10588,N_10502);
xnor U11087 (N_11087,N_10550,N_10905);
nand U11088 (N_11088,N_10689,N_10150);
and U11089 (N_11089,N_10832,N_10174);
or U11090 (N_11090,N_10789,N_10405);
and U11091 (N_11091,N_10993,N_10022);
nand U11092 (N_11092,N_10411,N_10286);
nor U11093 (N_11093,N_10798,N_10691);
xor U11094 (N_11094,N_10755,N_10093);
or U11095 (N_11095,N_10518,N_10563);
nand U11096 (N_11096,N_10173,N_10714);
xnor U11097 (N_11097,N_10102,N_10113);
and U11098 (N_11098,N_10300,N_10711);
and U11099 (N_11099,N_10226,N_10517);
or U11100 (N_11100,N_10210,N_10777);
or U11101 (N_11101,N_10034,N_10060);
and U11102 (N_11102,N_10680,N_10478);
xnor U11103 (N_11103,N_10388,N_10119);
xnor U11104 (N_11104,N_10149,N_10454);
or U11105 (N_11105,N_10963,N_10494);
xnor U11106 (N_11106,N_10771,N_10658);
or U11107 (N_11107,N_10648,N_10600);
nand U11108 (N_11108,N_10338,N_10672);
or U11109 (N_11109,N_10187,N_10800);
nand U11110 (N_11110,N_10415,N_10385);
nand U11111 (N_11111,N_10086,N_10495);
or U11112 (N_11112,N_10989,N_10844);
and U11113 (N_11113,N_10797,N_10864);
nand U11114 (N_11114,N_10975,N_10483);
and U11115 (N_11115,N_10551,N_10417);
nor U11116 (N_11116,N_10972,N_10913);
nand U11117 (N_11117,N_10625,N_10626);
xor U11118 (N_11118,N_10374,N_10100);
xnor U11119 (N_11119,N_10747,N_10969);
and U11120 (N_11120,N_10110,N_10726);
nor U11121 (N_11121,N_10540,N_10524);
and U11122 (N_11122,N_10192,N_10386);
nor U11123 (N_11123,N_10914,N_10541);
and U11124 (N_11124,N_10700,N_10614);
nand U11125 (N_11125,N_10384,N_10290);
nor U11126 (N_11126,N_10108,N_10802);
xnor U11127 (N_11127,N_10104,N_10376);
and U11128 (N_11128,N_10944,N_10253);
nand U11129 (N_11129,N_10581,N_10996);
nor U11130 (N_11130,N_10015,N_10804);
nand U11131 (N_11131,N_10489,N_10849);
nand U11132 (N_11132,N_10008,N_10673);
xnor U11133 (N_11133,N_10046,N_10464);
nor U11134 (N_11134,N_10021,N_10828);
nor U11135 (N_11135,N_10227,N_10001);
nand U11136 (N_11136,N_10764,N_10951);
nand U11137 (N_11137,N_10340,N_10661);
xor U11138 (N_11138,N_10252,N_10992);
nand U11139 (N_11139,N_10171,N_10179);
xnor U11140 (N_11140,N_10133,N_10081);
nand U11141 (N_11141,N_10299,N_10940);
nand U11142 (N_11142,N_10868,N_10729);
nand U11143 (N_11143,N_10430,N_10130);
or U11144 (N_11144,N_10967,N_10982);
nor U11145 (N_11145,N_10740,N_10189);
or U11146 (N_11146,N_10665,N_10602);
or U11147 (N_11147,N_10289,N_10098);
nand U11148 (N_11148,N_10296,N_10330);
nand U11149 (N_11149,N_10754,N_10097);
xor U11150 (N_11150,N_10678,N_10413);
nand U11151 (N_11151,N_10644,N_10621);
nor U11152 (N_11152,N_10534,N_10617);
nor U11153 (N_11153,N_10748,N_10208);
and U11154 (N_11154,N_10249,N_10202);
and U11155 (N_11155,N_10120,N_10535);
or U11156 (N_11156,N_10075,N_10244);
nor U11157 (N_11157,N_10653,N_10301);
nor U11158 (N_11158,N_10669,N_10640);
or U11159 (N_11159,N_10791,N_10318);
nand U11160 (N_11160,N_10037,N_10707);
and U11161 (N_11161,N_10934,N_10235);
nor U11162 (N_11162,N_10012,N_10334);
and U11163 (N_11163,N_10632,N_10875);
nor U11164 (N_11164,N_10593,N_10782);
or U11165 (N_11165,N_10776,N_10434);
nor U11166 (N_11166,N_10462,N_10265);
nor U11167 (N_11167,N_10509,N_10423);
xor U11168 (N_11168,N_10724,N_10794);
and U11169 (N_11169,N_10452,N_10135);
nand U11170 (N_11170,N_10333,N_10543);
nor U11171 (N_11171,N_10567,N_10881);
or U11172 (N_11172,N_10780,N_10854);
xor U11173 (N_11173,N_10988,N_10536);
and U11174 (N_11174,N_10850,N_10395);
xnor U11175 (N_11175,N_10056,N_10878);
or U11176 (N_11176,N_10116,N_10767);
nand U11177 (N_11177,N_10146,N_10115);
nor U11178 (N_11178,N_10916,N_10744);
and U11179 (N_11179,N_10885,N_10928);
nor U11180 (N_11180,N_10811,N_10984);
nand U11181 (N_11181,N_10090,N_10515);
nand U11182 (N_11182,N_10806,N_10014);
nor U11183 (N_11183,N_10643,N_10738);
and U11184 (N_11184,N_10705,N_10507);
nor U11185 (N_11185,N_10792,N_10309);
and U11186 (N_11186,N_10428,N_10156);
and U11187 (N_11187,N_10178,N_10078);
xnor U11188 (N_11188,N_10138,N_10117);
nor U11189 (N_11189,N_10931,N_10266);
and U11190 (N_11190,N_10118,N_10401);
or U11191 (N_11191,N_10319,N_10929);
xor U11192 (N_11192,N_10751,N_10939);
nand U11193 (N_11193,N_10114,N_10026);
xnor U11194 (N_11194,N_10513,N_10399);
or U11195 (N_11195,N_10964,N_10242);
xor U11196 (N_11196,N_10718,N_10438);
xor U11197 (N_11197,N_10228,N_10728);
nor U11198 (N_11198,N_10439,N_10609);
or U11199 (N_11199,N_10315,N_10267);
or U11200 (N_11200,N_10158,N_10381);
xnor U11201 (N_11201,N_10396,N_10067);
and U11202 (N_11202,N_10364,N_10168);
and U11203 (N_11203,N_10710,N_10491);
or U11204 (N_11204,N_10196,N_10897);
nand U11205 (N_11205,N_10546,N_10820);
and U11206 (N_11206,N_10433,N_10959);
nor U11207 (N_11207,N_10279,N_10263);
nand U11208 (N_11208,N_10835,N_10241);
xor U11209 (N_11209,N_10592,N_10481);
nand U11210 (N_11210,N_10899,N_10978);
xor U11211 (N_11211,N_10645,N_10520);
nand U11212 (N_11212,N_10247,N_10412);
nor U11213 (N_11213,N_10057,N_10601);
and U11214 (N_11214,N_10474,N_10424);
nor U11215 (N_11215,N_10076,N_10264);
nand U11216 (N_11216,N_10091,N_10248);
xor U11217 (N_11217,N_10918,N_10105);
xor U11218 (N_11218,N_10087,N_10923);
nand U11219 (N_11219,N_10061,N_10441);
nor U11220 (N_11220,N_10514,N_10161);
nor U11221 (N_11221,N_10882,N_10936);
or U11222 (N_11222,N_10341,N_10597);
or U11223 (N_11223,N_10649,N_10468);
nand U11224 (N_11224,N_10829,N_10372);
xor U11225 (N_11225,N_10742,N_10371);
and U11226 (N_11226,N_10634,N_10063);
nand U11227 (N_11227,N_10783,N_10450);
xnor U11228 (N_11228,N_10095,N_10663);
and U11229 (N_11229,N_10047,N_10407);
nor U11230 (N_11230,N_10089,N_10222);
or U11231 (N_11231,N_10741,N_10259);
nand U11232 (N_11232,N_10183,N_10453);
xnor U11233 (N_11233,N_10209,N_10305);
and U11234 (N_11234,N_10092,N_10556);
nand U11235 (N_11235,N_10671,N_10207);
or U11236 (N_11236,N_10823,N_10282);
xnor U11237 (N_11237,N_10200,N_10980);
and U11238 (N_11238,N_10770,N_10313);
and U11239 (N_11239,N_10532,N_10809);
nand U11240 (N_11240,N_10960,N_10888);
xnor U11241 (N_11241,N_10258,N_10231);
and U11242 (N_11242,N_10205,N_10933);
nor U11243 (N_11243,N_10758,N_10516);
nor U11244 (N_11244,N_10303,N_10763);
xnor U11245 (N_11245,N_10172,N_10927);
nor U11246 (N_11246,N_10292,N_10373);
and U11247 (N_11247,N_10773,N_10136);
or U11248 (N_11248,N_10493,N_10659);
xor U11249 (N_11249,N_10482,N_10697);
nand U11250 (N_11250,N_10394,N_10143);
xnor U11251 (N_11251,N_10025,N_10638);
nand U11252 (N_11252,N_10237,N_10871);
xor U11253 (N_11253,N_10197,N_10733);
and U11254 (N_11254,N_10945,N_10793);
xnor U11255 (N_11255,N_10656,N_10243);
or U11256 (N_11256,N_10387,N_10606);
nor U11257 (N_11257,N_10817,N_10486);
nor U11258 (N_11258,N_10575,N_10861);
nand U11259 (N_11259,N_10628,N_10530);
or U11260 (N_11260,N_10487,N_10377);
nand U11261 (N_11261,N_10088,N_10094);
xor U11262 (N_11262,N_10326,N_10790);
or U11263 (N_11263,N_10528,N_10968);
xor U11264 (N_11264,N_10351,N_10317);
nand U11265 (N_11265,N_10162,N_10957);
nand U11266 (N_11266,N_10688,N_10485);
nor U11267 (N_11267,N_10278,N_10261);
and U11268 (N_11268,N_10892,N_10447);
nor U11269 (N_11269,N_10414,N_10498);
nand U11270 (N_11270,N_10255,N_10785);
nand U11271 (N_11271,N_10778,N_10028);
nand U11272 (N_11272,N_10112,N_10526);
and U11273 (N_11273,N_10375,N_10033);
and U11274 (N_11274,N_10041,N_10504);
xnor U11275 (N_11275,N_10490,N_10690);
and U11276 (N_11276,N_10736,N_10538);
or U11277 (N_11277,N_10288,N_10052);
and U11278 (N_11278,N_10038,N_10324);
nand U11279 (N_11279,N_10470,N_10971);
nand U11280 (N_11280,N_10555,N_10560);
nand U11281 (N_11281,N_10362,N_10409);
and U11282 (N_11282,N_10527,N_10035);
nor U11283 (N_11283,N_10836,N_10873);
xor U11284 (N_11284,N_10683,N_10435);
and U11285 (N_11285,N_10465,N_10070);
xor U11286 (N_11286,N_10182,N_10361);
and U11287 (N_11287,N_10212,N_10910);
and U11288 (N_11288,N_10219,N_10962);
nand U11289 (N_11289,N_10459,N_10181);
or U11290 (N_11290,N_10667,N_10568);
and U11291 (N_11291,N_10920,N_10692);
and U11292 (N_11292,N_10354,N_10838);
xor U11293 (N_11293,N_10223,N_10629);
nor U11294 (N_11294,N_10446,N_10185);
nand U11295 (N_11295,N_10131,N_10687);
or U11296 (N_11296,N_10921,N_10698);
nand U11297 (N_11297,N_10304,N_10307);
and U11298 (N_11298,N_10819,N_10007);
xor U11299 (N_11299,N_10272,N_10082);
or U11300 (N_11300,N_10735,N_10674);
or U11301 (N_11301,N_10031,N_10876);
xnor U11302 (N_11302,N_10273,N_10884);
or U11303 (N_11303,N_10029,N_10883);
nor U11304 (N_11304,N_10670,N_10765);
nand U11305 (N_11305,N_10937,N_10544);
nand U11306 (N_11306,N_10463,N_10725);
and U11307 (N_11307,N_10347,N_10677);
or U11308 (N_11308,N_10908,N_10281);
or U11309 (N_11309,N_10467,N_10574);
and U11310 (N_11310,N_10402,N_10635);
nand U11311 (N_11311,N_10256,N_10979);
and U11312 (N_11312,N_10217,N_10746);
nor U11313 (N_11313,N_10011,N_10397);
xnor U11314 (N_11314,N_10859,N_10175);
and U11315 (N_11315,N_10280,N_10821);
xnor U11316 (N_11316,N_10952,N_10365);
and U11317 (N_11317,N_10080,N_10814);
and U11318 (N_11318,N_10444,N_10681);
or U11319 (N_11319,N_10858,N_10229);
or U11320 (N_11320,N_10853,N_10363);
xor U11321 (N_11321,N_10458,N_10084);
nor U11322 (N_11322,N_10529,N_10477);
nor U11323 (N_11323,N_10573,N_10901);
or U11324 (N_11324,N_10732,N_10930);
nor U11325 (N_11325,N_10719,N_10511);
xnor U11326 (N_11326,N_10852,N_10251);
nand U11327 (N_11327,N_10519,N_10079);
and U11328 (N_11328,N_10557,N_10584);
or U11329 (N_11329,N_10500,N_10195);
nor U11330 (N_11330,N_10942,N_10366);
or U11331 (N_11331,N_10276,N_10622);
or U11332 (N_11332,N_10069,N_10225);
nor U11333 (N_11333,N_10215,N_10624);
and U11334 (N_11334,N_10039,N_10501);
or U11335 (N_11335,N_10269,N_10866);
nand U11336 (N_11336,N_10077,N_10024);
or U11337 (N_11337,N_10633,N_10406);
xnor U11338 (N_11338,N_10027,N_10472);
and U11339 (N_11339,N_10577,N_10542);
nor U11340 (N_11340,N_10576,N_10637);
or U11341 (N_11341,N_10730,N_10295);
nor U11342 (N_11342,N_10322,N_10966);
xnor U11343 (N_11343,N_10236,N_10339);
nand U11344 (N_11344,N_10337,N_10049);
and U11345 (N_11345,N_10419,N_10533);
or U11346 (N_11346,N_10431,N_10976);
xnor U11347 (N_11347,N_10141,N_10646);
or U11348 (N_11348,N_10457,N_10380);
or U11349 (N_11349,N_10006,N_10085);
nand U11350 (N_11350,N_10824,N_10682);
and U11351 (N_11351,N_10499,N_10262);
nand U11352 (N_11352,N_10221,N_10422);
or U11353 (N_11353,N_10679,N_10198);
xor U11354 (N_11354,N_10473,N_10561);
nor U11355 (N_11355,N_10147,N_10961);
and U11356 (N_11356,N_10055,N_10211);
nor U11357 (N_11357,N_10685,N_10872);
nand U11358 (N_11358,N_10355,N_10660);
nor U11359 (N_11359,N_10990,N_10246);
or U11360 (N_11360,N_10619,N_10564);
xor U11361 (N_11361,N_10987,N_10408);
and U11362 (N_11362,N_10352,N_10774);
and U11363 (N_11363,N_10314,N_10566);
or U11364 (N_11364,N_10904,N_10915);
and U11365 (N_11365,N_10702,N_10716);
nand U11366 (N_11366,N_10847,N_10549);
nor U11367 (N_11367,N_10383,N_10615);
or U11368 (N_11368,N_10356,N_10302);
nor U11369 (N_11369,N_10331,N_10013);
or U11370 (N_11370,N_10254,N_10461);
xnor U11371 (N_11371,N_10919,N_10786);
nand U11372 (N_11372,N_10416,N_10074);
and U11373 (N_11373,N_10357,N_10652);
or U11374 (N_11374,N_10862,N_10429);
and U11375 (N_11375,N_10909,N_10613);
xor U11376 (N_11376,N_10059,N_10180);
and U11377 (N_11377,N_10194,N_10157);
and U11378 (N_11378,N_10639,N_10848);
and U11379 (N_11379,N_10623,N_10443);
and U11380 (N_11380,N_10616,N_10795);
or U11381 (N_11381,N_10044,N_10432);
nor U11382 (N_11382,N_10970,N_10418);
nor U11383 (N_11383,N_10066,N_10857);
or U11384 (N_11384,N_10801,N_10506);
nand U11385 (N_11385,N_10610,N_10285);
or U11386 (N_11386,N_10803,N_10991);
nand U11387 (N_11387,N_10323,N_10019);
xor U11388 (N_11388,N_10787,N_10650);
and U11389 (N_11389,N_10144,N_10715);
nand U11390 (N_11390,N_10275,N_10456);
nand U11391 (N_11391,N_10420,N_10902);
and U11392 (N_11392,N_10045,N_10004);
nor U11393 (N_11393,N_10911,N_10686);
and U11394 (N_11394,N_10974,N_10316);
nor U11395 (N_11395,N_10895,N_10410);
xor U11396 (N_11396,N_10287,N_10328);
nand U11397 (N_11397,N_10981,N_10713);
nor U11398 (N_11398,N_10717,N_10400);
or U11399 (N_11399,N_10708,N_10891);
nor U11400 (N_11400,N_10831,N_10917);
xnor U11401 (N_11401,N_10122,N_10580);
and U11402 (N_11402,N_10166,N_10107);
xnor U11403 (N_11403,N_10065,N_10826);
nand U11404 (N_11404,N_10238,N_10139);
nor U11405 (N_11405,N_10346,N_10148);
nand U11406 (N_11406,N_10240,N_10204);
or U11407 (N_11407,N_10949,N_10126);
xnor U11408 (N_11408,N_10865,N_10578);
nor U11409 (N_11409,N_10709,N_10393);
nand U11410 (N_11410,N_10054,N_10260);
or U11411 (N_11411,N_10995,N_10779);
or U11412 (N_11412,N_10867,N_10050);
xor U11413 (N_11413,N_10522,N_10191);
nor U11414 (N_11414,N_10554,N_10201);
or U11415 (N_11415,N_10186,N_10946);
xor U11416 (N_11416,N_10941,N_10762);
nor U11417 (N_11417,N_10775,N_10907);
nand U11418 (N_11418,N_10426,N_10596);
xnor U11419 (N_11419,N_10985,N_10842);
and U11420 (N_11420,N_10760,N_10603);
xor U11421 (N_11421,N_10796,N_10460);
xnor U11422 (N_11422,N_10404,N_10391);
nand U11423 (N_11423,N_10887,N_10390);
xnor U11424 (N_11424,N_10948,N_10704);
nand U11425 (N_11425,N_10630,N_10664);
or U11426 (N_11426,N_10935,N_10403);
xnor U11427 (N_11427,N_10000,N_10586);
or U11428 (N_11428,N_10818,N_10368);
and U11429 (N_11429,N_10163,N_10245);
nor U11430 (N_11430,N_10833,N_10072);
nor U11431 (N_11431,N_10032,N_10184);
or U11432 (N_11432,N_10306,N_10703);
nor U11433 (N_11433,N_10565,N_10505);
nand U11434 (N_11434,N_10723,N_10165);
nor U11435 (N_11435,N_10132,N_10277);
nor U11436 (N_11436,N_10898,N_10745);
xor U11437 (N_11437,N_10479,N_10436);
xor U11438 (N_11438,N_10152,N_10983);
or U11439 (N_11439,N_10455,N_10360);
or U11440 (N_11440,N_10788,N_10140);
xnor U11441 (N_11441,N_10636,N_10320);
xor U11442 (N_11442,N_10874,N_10572);
or U11443 (N_11443,N_10815,N_10155);
nand U11444 (N_11444,N_10827,N_10595);
and U11445 (N_11445,N_10003,N_10475);
or U11446 (N_11446,N_10284,N_10224);
nor U11447 (N_11447,N_10484,N_10250);
nand U11448 (N_11448,N_10727,N_10851);
or U11449 (N_11449,N_10053,N_10206);
nand U11450 (N_11450,N_10159,N_10752);
nor U11451 (N_11451,N_10684,N_10073);
xor U11452 (N_11452,N_10220,N_10825);
and U11453 (N_11453,N_10757,N_10846);
or U11454 (N_11454,N_10612,N_10124);
and U11455 (N_11455,N_10750,N_10570);
and U11456 (N_11456,N_10421,N_10998);
nand U11457 (N_11457,N_10030,N_10358);
nand U11458 (N_11458,N_10932,N_10547);
nor U11459 (N_11459,N_10170,N_10137);
or U11460 (N_11460,N_10845,N_10232);
nand U11461 (N_11461,N_10657,N_10176);
and U11462 (N_11462,N_10058,N_10497);
nor U11463 (N_11463,N_10379,N_10062);
xor U11464 (N_11464,N_10784,N_10367);
or U11465 (N_11465,N_10127,N_10293);
xnor U11466 (N_11466,N_10167,N_10558);
nand U11467 (N_11467,N_10641,N_10582);
xnor U11468 (N_11468,N_10048,N_10627);
and U11469 (N_11469,N_10239,N_10370);
xnor U11470 (N_11470,N_10445,N_10734);
xnor U11471 (N_11471,N_10822,N_10545);
and U11472 (N_11472,N_10123,N_10537);
or U11473 (N_11473,N_10552,N_10234);
or U11474 (N_11474,N_10655,N_10128);
xor U11475 (N_11475,N_10068,N_10002);
or U11476 (N_11476,N_10099,N_10389);
xnor U11477 (N_11477,N_10810,N_10759);
xor U11478 (N_11478,N_10230,N_10040);
or U11479 (N_11479,N_10051,N_10216);
and U11480 (N_11480,N_10855,N_10125);
nor U11481 (N_11481,N_10153,N_10756);
and U11482 (N_11482,N_10548,N_10594);
xnor U11483 (N_11483,N_10647,N_10720);
xnor U11484 (N_11484,N_10257,N_10553);
and U11485 (N_11485,N_10327,N_10743);
or U11486 (N_11486,N_10604,N_10869);
xnor U11487 (N_11487,N_10877,N_10958);
xnor U11488 (N_11488,N_10712,N_10344);
nor U11489 (N_11489,N_10569,N_10662);
nand U11490 (N_11490,N_10471,N_10766);
and U11491 (N_11491,N_10607,N_10274);
and U11492 (N_11492,N_10083,N_10808);
or U11493 (N_11493,N_10488,N_10398);
nand U11494 (N_11494,N_10348,N_10579);
or U11495 (N_11495,N_10903,N_10841);
nand U11496 (N_11496,N_10539,N_10890);
xor U11497 (N_11497,N_10382,N_10425);
or U11498 (N_11498,N_10188,N_10925);
or U11499 (N_11499,N_10694,N_10956);
or U11500 (N_11500,N_10082,N_10722);
xnor U11501 (N_11501,N_10889,N_10707);
and U11502 (N_11502,N_10035,N_10244);
or U11503 (N_11503,N_10274,N_10072);
nor U11504 (N_11504,N_10560,N_10256);
nor U11505 (N_11505,N_10073,N_10121);
and U11506 (N_11506,N_10583,N_10045);
or U11507 (N_11507,N_10910,N_10621);
nor U11508 (N_11508,N_10035,N_10117);
nor U11509 (N_11509,N_10552,N_10499);
xor U11510 (N_11510,N_10041,N_10858);
xnor U11511 (N_11511,N_10919,N_10489);
or U11512 (N_11512,N_10784,N_10077);
or U11513 (N_11513,N_10472,N_10610);
and U11514 (N_11514,N_10194,N_10474);
or U11515 (N_11515,N_10612,N_10789);
xor U11516 (N_11516,N_10436,N_10216);
and U11517 (N_11517,N_10944,N_10441);
nand U11518 (N_11518,N_10184,N_10675);
xor U11519 (N_11519,N_10890,N_10140);
xor U11520 (N_11520,N_10278,N_10295);
or U11521 (N_11521,N_10488,N_10422);
and U11522 (N_11522,N_10510,N_10322);
xnor U11523 (N_11523,N_10691,N_10654);
nor U11524 (N_11524,N_10165,N_10778);
xor U11525 (N_11525,N_10068,N_10565);
and U11526 (N_11526,N_10264,N_10030);
nand U11527 (N_11527,N_10062,N_10614);
nand U11528 (N_11528,N_10751,N_10016);
or U11529 (N_11529,N_10872,N_10340);
nor U11530 (N_11530,N_10185,N_10093);
nand U11531 (N_11531,N_10523,N_10971);
or U11532 (N_11532,N_10086,N_10518);
or U11533 (N_11533,N_10113,N_10143);
and U11534 (N_11534,N_10813,N_10351);
nand U11535 (N_11535,N_10178,N_10942);
nor U11536 (N_11536,N_10804,N_10625);
nor U11537 (N_11537,N_10836,N_10469);
or U11538 (N_11538,N_10366,N_10419);
nand U11539 (N_11539,N_10348,N_10884);
xor U11540 (N_11540,N_10406,N_10767);
and U11541 (N_11541,N_10724,N_10083);
or U11542 (N_11542,N_10638,N_10445);
nand U11543 (N_11543,N_10434,N_10570);
xor U11544 (N_11544,N_10488,N_10980);
nand U11545 (N_11545,N_10269,N_10785);
and U11546 (N_11546,N_10564,N_10459);
nor U11547 (N_11547,N_10383,N_10123);
or U11548 (N_11548,N_10551,N_10964);
nand U11549 (N_11549,N_10831,N_10453);
or U11550 (N_11550,N_10859,N_10756);
xor U11551 (N_11551,N_10857,N_10383);
and U11552 (N_11552,N_10559,N_10300);
or U11553 (N_11553,N_10719,N_10289);
and U11554 (N_11554,N_10850,N_10857);
xnor U11555 (N_11555,N_10849,N_10437);
or U11556 (N_11556,N_10798,N_10690);
nand U11557 (N_11557,N_10105,N_10645);
nand U11558 (N_11558,N_10641,N_10213);
and U11559 (N_11559,N_10476,N_10315);
nand U11560 (N_11560,N_10764,N_10571);
nor U11561 (N_11561,N_10699,N_10800);
nand U11562 (N_11562,N_10727,N_10974);
nor U11563 (N_11563,N_10916,N_10991);
nand U11564 (N_11564,N_10757,N_10604);
nand U11565 (N_11565,N_10937,N_10611);
and U11566 (N_11566,N_10139,N_10041);
nor U11567 (N_11567,N_10706,N_10636);
xor U11568 (N_11568,N_10890,N_10449);
nor U11569 (N_11569,N_10724,N_10194);
xnor U11570 (N_11570,N_10325,N_10725);
xor U11571 (N_11571,N_10065,N_10035);
and U11572 (N_11572,N_10486,N_10848);
and U11573 (N_11573,N_10811,N_10467);
and U11574 (N_11574,N_10659,N_10409);
nor U11575 (N_11575,N_10932,N_10127);
or U11576 (N_11576,N_10587,N_10260);
or U11577 (N_11577,N_10701,N_10758);
or U11578 (N_11578,N_10067,N_10870);
nor U11579 (N_11579,N_10305,N_10980);
nor U11580 (N_11580,N_10495,N_10501);
nand U11581 (N_11581,N_10892,N_10041);
nor U11582 (N_11582,N_10141,N_10418);
nand U11583 (N_11583,N_10649,N_10590);
nand U11584 (N_11584,N_10844,N_10708);
nor U11585 (N_11585,N_10462,N_10835);
nand U11586 (N_11586,N_10941,N_10266);
nand U11587 (N_11587,N_10420,N_10364);
nand U11588 (N_11588,N_10449,N_10818);
nor U11589 (N_11589,N_10073,N_10817);
and U11590 (N_11590,N_10150,N_10215);
xnor U11591 (N_11591,N_10300,N_10836);
or U11592 (N_11592,N_10896,N_10724);
nor U11593 (N_11593,N_10447,N_10430);
and U11594 (N_11594,N_10445,N_10686);
xnor U11595 (N_11595,N_10196,N_10668);
or U11596 (N_11596,N_10990,N_10868);
xor U11597 (N_11597,N_10111,N_10176);
or U11598 (N_11598,N_10366,N_10206);
and U11599 (N_11599,N_10616,N_10820);
xnor U11600 (N_11600,N_10671,N_10810);
xnor U11601 (N_11601,N_10781,N_10733);
and U11602 (N_11602,N_10924,N_10098);
and U11603 (N_11603,N_10574,N_10739);
nor U11604 (N_11604,N_10983,N_10359);
nor U11605 (N_11605,N_10023,N_10350);
and U11606 (N_11606,N_10202,N_10514);
and U11607 (N_11607,N_10901,N_10881);
or U11608 (N_11608,N_10187,N_10441);
xor U11609 (N_11609,N_10503,N_10363);
xor U11610 (N_11610,N_10289,N_10248);
and U11611 (N_11611,N_10928,N_10076);
or U11612 (N_11612,N_10248,N_10565);
and U11613 (N_11613,N_10720,N_10941);
and U11614 (N_11614,N_10681,N_10087);
nor U11615 (N_11615,N_10262,N_10475);
or U11616 (N_11616,N_10828,N_10190);
nand U11617 (N_11617,N_10188,N_10672);
nand U11618 (N_11618,N_10832,N_10284);
nand U11619 (N_11619,N_10541,N_10431);
or U11620 (N_11620,N_10196,N_10217);
or U11621 (N_11621,N_10482,N_10884);
xor U11622 (N_11622,N_10698,N_10450);
nand U11623 (N_11623,N_10674,N_10707);
nor U11624 (N_11624,N_10589,N_10924);
nand U11625 (N_11625,N_10776,N_10345);
nand U11626 (N_11626,N_10161,N_10208);
nor U11627 (N_11627,N_10716,N_10782);
nand U11628 (N_11628,N_10115,N_10855);
and U11629 (N_11629,N_10410,N_10575);
nand U11630 (N_11630,N_10264,N_10746);
nand U11631 (N_11631,N_10600,N_10634);
or U11632 (N_11632,N_10048,N_10803);
and U11633 (N_11633,N_10996,N_10466);
nand U11634 (N_11634,N_10992,N_10706);
nand U11635 (N_11635,N_10483,N_10225);
or U11636 (N_11636,N_10081,N_10430);
or U11637 (N_11637,N_10160,N_10730);
or U11638 (N_11638,N_10884,N_10798);
and U11639 (N_11639,N_10269,N_10389);
nor U11640 (N_11640,N_10723,N_10465);
xnor U11641 (N_11641,N_10098,N_10813);
xor U11642 (N_11642,N_10168,N_10855);
nand U11643 (N_11643,N_10371,N_10471);
and U11644 (N_11644,N_10355,N_10330);
nand U11645 (N_11645,N_10660,N_10760);
nor U11646 (N_11646,N_10235,N_10006);
xnor U11647 (N_11647,N_10238,N_10593);
nand U11648 (N_11648,N_10382,N_10112);
nand U11649 (N_11649,N_10659,N_10735);
nor U11650 (N_11650,N_10169,N_10007);
and U11651 (N_11651,N_10723,N_10677);
xnor U11652 (N_11652,N_10912,N_10012);
nor U11653 (N_11653,N_10722,N_10046);
or U11654 (N_11654,N_10449,N_10136);
nor U11655 (N_11655,N_10814,N_10214);
or U11656 (N_11656,N_10070,N_10036);
and U11657 (N_11657,N_10051,N_10586);
and U11658 (N_11658,N_10423,N_10743);
xor U11659 (N_11659,N_10338,N_10852);
or U11660 (N_11660,N_10826,N_10536);
xor U11661 (N_11661,N_10793,N_10546);
and U11662 (N_11662,N_10927,N_10162);
or U11663 (N_11663,N_10995,N_10902);
or U11664 (N_11664,N_10385,N_10617);
or U11665 (N_11665,N_10238,N_10638);
nand U11666 (N_11666,N_10459,N_10589);
nor U11667 (N_11667,N_10857,N_10601);
or U11668 (N_11668,N_10983,N_10292);
nand U11669 (N_11669,N_10886,N_10374);
nand U11670 (N_11670,N_10232,N_10203);
xor U11671 (N_11671,N_10583,N_10248);
and U11672 (N_11672,N_10050,N_10956);
xnor U11673 (N_11673,N_10573,N_10819);
xnor U11674 (N_11674,N_10063,N_10073);
nand U11675 (N_11675,N_10076,N_10881);
or U11676 (N_11676,N_10514,N_10267);
nand U11677 (N_11677,N_10496,N_10923);
and U11678 (N_11678,N_10580,N_10379);
nor U11679 (N_11679,N_10653,N_10676);
and U11680 (N_11680,N_10753,N_10996);
or U11681 (N_11681,N_10001,N_10127);
or U11682 (N_11682,N_10745,N_10842);
xor U11683 (N_11683,N_10333,N_10074);
nor U11684 (N_11684,N_10646,N_10743);
nand U11685 (N_11685,N_10712,N_10822);
nor U11686 (N_11686,N_10594,N_10376);
xnor U11687 (N_11687,N_10629,N_10213);
and U11688 (N_11688,N_10524,N_10660);
and U11689 (N_11689,N_10346,N_10386);
xnor U11690 (N_11690,N_10089,N_10659);
xnor U11691 (N_11691,N_10860,N_10066);
or U11692 (N_11692,N_10476,N_10493);
xor U11693 (N_11693,N_10253,N_10942);
xor U11694 (N_11694,N_10510,N_10209);
xor U11695 (N_11695,N_10115,N_10040);
nand U11696 (N_11696,N_10356,N_10382);
nor U11697 (N_11697,N_10276,N_10345);
or U11698 (N_11698,N_10236,N_10011);
nor U11699 (N_11699,N_10837,N_10060);
nand U11700 (N_11700,N_10480,N_10997);
nand U11701 (N_11701,N_10583,N_10404);
xor U11702 (N_11702,N_10887,N_10205);
nor U11703 (N_11703,N_10674,N_10101);
and U11704 (N_11704,N_10780,N_10478);
and U11705 (N_11705,N_10863,N_10900);
and U11706 (N_11706,N_10346,N_10432);
xnor U11707 (N_11707,N_10853,N_10214);
or U11708 (N_11708,N_10505,N_10303);
and U11709 (N_11709,N_10695,N_10328);
nor U11710 (N_11710,N_10409,N_10376);
nand U11711 (N_11711,N_10792,N_10832);
and U11712 (N_11712,N_10570,N_10860);
or U11713 (N_11713,N_10148,N_10184);
and U11714 (N_11714,N_10849,N_10645);
and U11715 (N_11715,N_10980,N_10609);
and U11716 (N_11716,N_10342,N_10241);
nand U11717 (N_11717,N_10744,N_10419);
and U11718 (N_11718,N_10642,N_10131);
or U11719 (N_11719,N_10762,N_10133);
nor U11720 (N_11720,N_10321,N_10975);
and U11721 (N_11721,N_10019,N_10448);
and U11722 (N_11722,N_10618,N_10776);
nor U11723 (N_11723,N_10790,N_10867);
xor U11724 (N_11724,N_10206,N_10975);
and U11725 (N_11725,N_10546,N_10421);
xnor U11726 (N_11726,N_10720,N_10746);
and U11727 (N_11727,N_10134,N_10226);
nor U11728 (N_11728,N_10190,N_10994);
and U11729 (N_11729,N_10011,N_10663);
nor U11730 (N_11730,N_10132,N_10983);
nor U11731 (N_11731,N_10701,N_10007);
nand U11732 (N_11732,N_10163,N_10823);
nand U11733 (N_11733,N_10191,N_10293);
or U11734 (N_11734,N_10905,N_10839);
nor U11735 (N_11735,N_10076,N_10630);
nand U11736 (N_11736,N_10828,N_10791);
nand U11737 (N_11737,N_10886,N_10864);
and U11738 (N_11738,N_10823,N_10013);
and U11739 (N_11739,N_10923,N_10187);
nor U11740 (N_11740,N_10239,N_10146);
nor U11741 (N_11741,N_10707,N_10709);
and U11742 (N_11742,N_10439,N_10918);
or U11743 (N_11743,N_10043,N_10011);
nand U11744 (N_11744,N_10162,N_10524);
nor U11745 (N_11745,N_10156,N_10213);
and U11746 (N_11746,N_10185,N_10528);
xor U11747 (N_11747,N_10611,N_10032);
nor U11748 (N_11748,N_10090,N_10829);
xnor U11749 (N_11749,N_10781,N_10259);
and U11750 (N_11750,N_10146,N_10955);
nand U11751 (N_11751,N_10802,N_10694);
nand U11752 (N_11752,N_10881,N_10011);
or U11753 (N_11753,N_10084,N_10642);
and U11754 (N_11754,N_10643,N_10268);
nand U11755 (N_11755,N_10948,N_10029);
nor U11756 (N_11756,N_10247,N_10264);
and U11757 (N_11757,N_10082,N_10053);
nand U11758 (N_11758,N_10969,N_10843);
xor U11759 (N_11759,N_10853,N_10090);
or U11760 (N_11760,N_10399,N_10174);
and U11761 (N_11761,N_10456,N_10822);
xnor U11762 (N_11762,N_10008,N_10034);
nor U11763 (N_11763,N_10234,N_10788);
nor U11764 (N_11764,N_10052,N_10313);
or U11765 (N_11765,N_10970,N_10497);
nor U11766 (N_11766,N_10069,N_10295);
nand U11767 (N_11767,N_10539,N_10530);
xor U11768 (N_11768,N_10354,N_10226);
nor U11769 (N_11769,N_10274,N_10108);
and U11770 (N_11770,N_10864,N_10889);
xor U11771 (N_11771,N_10400,N_10505);
or U11772 (N_11772,N_10540,N_10500);
or U11773 (N_11773,N_10032,N_10839);
or U11774 (N_11774,N_10048,N_10461);
or U11775 (N_11775,N_10129,N_10687);
and U11776 (N_11776,N_10180,N_10491);
nor U11777 (N_11777,N_10848,N_10028);
or U11778 (N_11778,N_10296,N_10329);
xor U11779 (N_11779,N_10004,N_10357);
nor U11780 (N_11780,N_10141,N_10178);
xor U11781 (N_11781,N_10688,N_10213);
nor U11782 (N_11782,N_10815,N_10399);
and U11783 (N_11783,N_10690,N_10349);
nand U11784 (N_11784,N_10754,N_10780);
and U11785 (N_11785,N_10211,N_10873);
or U11786 (N_11786,N_10047,N_10060);
nand U11787 (N_11787,N_10850,N_10324);
nand U11788 (N_11788,N_10091,N_10596);
and U11789 (N_11789,N_10735,N_10309);
nor U11790 (N_11790,N_10138,N_10763);
xor U11791 (N_11791,N_10340,N_10043);
and U11792 (N_11792,N_10812,N_10482);
and U11793 (N_11793,N_10513,N_10201);
nand U11794 (N_11794,N_10577,N_10583);
and U11795 (N_11795,N_10589,N_10150);
nor U11796 (N_11796,N_10062,N_10207);
nor U11797 (N_11797,N_10388,N_10080);
nor U11798 (N_11798,N_10335,N_10665);
xnor U11799 (N_11799,N_10273,N_10685);
xnor U11800 (N_11800,N_10961,N_10893);
nand U11801 (N_11801,N_10351,N_10849);
nand U11802 (N_11802,N_10786,N_10312);
nor U11803 (N_11803,N_10997,N_10620);
xor U11804 (N_11804,N_10936,N_10728);
and U11805 (N_11805,N_10015,N_10174);
nor U11806 (N_11806,N_10736,N_10693);
nor U11807 (N_11807,N_10181,N_10997);
nor U11808 (N_11808,N_10086,N_10905);
and U11809 (N_11809,N_10618,N_10125);
nand U11810 (N_11810,N_10836,N_10257);
or U11811 (N_11811,N_10260,N_10266);
xnor U11812 (N_11812,N_10214,N_10358);
nand U11813 (N_11813,N_10787,N_10928);
nand U11814 (N_11814,N_10387,N_10119);
nand U11815 (N_11815,N_10208,N_10979);
or U11816 (N_11816,N_10315,N_10935);
nor U11817 (N_11817,N_10350,N_10715);
and U11818 (N_11818,N_10033,N_10258);
xor U11819 (N_11819,N_10523,N_10967);
or U11820 (N_11820,N_10456,N_10361);
xor U11821 (N_11821,N_10388,N_10832);
nand U11822 (N_11822,N_10441,N_10815);
and U11823 (N_11823,N_10693,N_10556);
xor U11824 (N_11824,N_10136,N_10966);
nor U11825 (N_11825,N_10440,N_10507);
nand U11826 (N_11826,N_10830,N_10028);
nor U11827 (N_11827,N_10167,N_10567);
and U11828 (N_11828,N_10019,N_10722);
nor U11829 (N_11829,N_10556,N_10772);
or U11830 (N_11830,N_10206,N_10964);
nor U11831 (N_11831,N_10836,N_10474);
or U11832 (N_11832,N_10344,N_10188);
or U11833 (N_11833,N_10265,N_10026);
nand U11834 (N_11834,N_10141,N_10506);
or U11835 (N_11835,N_10291,N_10513);
nor U11836 (N_11836,N_10537,N_10632);
or U11837 (N_11837,N_10496,N_10576);
xnor U11838 (N_11838,N_10545,N_10567);
nor U11839 (N_11839,N_10575,N_10323);
nor U11840 (N_11840,N_10581,N_10988);
nand U11841 (N_11841,N_10051,N_10133);
and U11842 (N_11842,N_10664,N_10163);
or U11843 (N_11843,N_10550,N_10157);
nand U11844 (N_11844,N_10304,N_10953);
nand U11845 (N_11845,N_10949,N_10276);
xor U11846 (N_11846,N_10520,N_10008);
nand U11847 (N_11847,N_10189,N_10856);
nand U11848 (N_11848,N_10347,N_10193);
nor U11849 (N_11849,N_10266,N_10241);
and U11850 (N_11850,N_10376,N_10665);
nand U11851 (N_11851,N_10347,N_10971);
xnor U11852 (N_11852,N_10397,N_10258);
or U11853 (N_11853,N_10539,N_10281);
nor U11854 (N_11854,N_10948,N_10581);
xor U11855 (N_11855,N_10950,N_10172);
and U11856 (N_11856,N_10162,N_10236);
xnor U11857 (N_11857,N_10677,N_10027);
nand U11858 (N_11858,N_10399,N_10318);
or U11859 (N_11859,N_10929,N_10228);
nor U11860 (N_11860,N_10488,N_10430);
nand U11861 (N_11861,N_10778,N_10148);
or U11862 (N_11862,N_10373,N_10382);
nand U11863 (N_11863,N_10953,N_10549);
or U11864 (N_11864,N_10114,N_10994);
or U11865 (N_11865,N_10112,N_10362);
and U11866 (N_11866,N_10918,N_10780);
nor U11867 (N_11867,N_10929,N_10245);
or U11868 (N_11868,N_10952,N_10518);
and U11869 (N_11869,N_10534,N_10426);
xor U11870 (N_11870,N_10492,N_10561);
nor U11871 (N_11871,N_10887,N_10350);
and U11872 (N_11872,N_10518,N_10832);
and U11873 (N_11873,N_10041,N_10324);
xor U11874 (N_11874,N_10273,N_10375);
xor U11875 (N_11875,N_10528,N_10660);
or U11876 (N_11876,N_10778,N_10306);
xnor U11877 (N_11877,N_10576,N_10600);
or U11878 (N_11878,N_10328,N_10251);
nand U11879 (N_11879,N_10638,N_10913);
and U11880 (N_11880,N_10265,N_10523);
nand U11881 (N_11881,N_10670,N_10745);
xor U11882 (N_11882,N_10141,N_10949);
xor U11883 (N_11883,N_10619,N_10730);
nand U11884 (N_11884,N_10414,N_10070);
or U11885 (N_11885,N_10772,N_10971);
and U11886 (N_11886,N_10204,N_10763);
nand U11887 (N_11887,N_10291,N_10709);
and U11888 (N_11888,N_10335,N_10987);
nor U11889 (N_11889,N_10262,N_10188);
xor U11890 (N_11890,N_10546,N_10985);
and U11891 (N_11891,N_10773,N_10214);
xor U11892 (N_11892,N_10410,N_10025);
nand U11893 (N_11893,N_10167,N_10111);
or U11894 (N_11894,N_10489,N_10992);
nor U11895 (N_11895,N_10344,N_10152);
or U11896 (N_11896,N_10484,N_10188);
nor U11897 (N_11897,N_10515,N_10773);
xnor U11898 (N_11898,N_10513,N_10972);
nand U11899 (N_11899,N_10393,N_10155);
xnor U11900 (N_11900,N_10710,N_10073);
nor U11901 (N_11901,N_10383,N_10559);
nor U11902 (N_11902,N_10430,N_10225);
or U11903 (N_11903,N_10848,N_10162);
nor U11904 (N_11904,N_10265,N_10111);
and U11905 (N_11905,N_10892,N_10552);
and U11906 (N_11906,N_10581,N_10179);
xnor U11907 (N_11907,N_10380,N_10207);
and U11908 (N_11908,N_10951,N_10663);
nand U11909 (N_11909,N_10008,N_10916);
nand U11910 (N_11910,N_10810,N_10458);
nand U11911 (N_11911,N_10011,N_10355);
nor U11912 (N_11912,N_10054,N_10015);
xor U11913 (N_11913,N_10855,N_10294);
xnor U11914 (N_11914,N_10088,N_10980);
nor U11915 (N_11915,N_10838,N_10769);
xnor U11916 (N_11916,N_10735,N_10996);
or U11917 (N_11917,N_10360,N_10138);
nand U11918 (N_11918,N_10657,N_10461);
nor U11919 (N_11919,N_10612,N_10467);
nand U11920 (N_11920,N_10330,N_10920);
and U11921 (N_11921,N_10556,N_10178);
or U11922 (N_11922,N_10144,N_10070);
or U11923 (N_11923,N_10462,N_10990);
xnor U11924 (N_11924,N_10749,N_10491);
and U11925 (N_11925,N_10340,N_10402);
nand U11926 (N_11926,N_10750,N_10605);
or U11927 (N_11927,N_10008,N_10971);
xor U11928 (N_11928,N_10235,N_10019);
nor U11929 (N_11929,N_10538,N_10362);
nand U11930 (N_11930,N_10049,N_10275);
nand U11931 (N_11931,N_10513,N_10707);
or U11932 (N_11932,N_10805,N_10284);
nand U11933 (N_11933,N_10818,N_10946);
nand U11934 (N_11934,N_10774,N_10522);
nand U11935 (N_11935,N_10584,N_10077);
nor U11936 (N_11936,N_10583,N_10770);
or U11937 (N_11937,N_10487,N_10189);
or U11938 (N_11938,N_10176,N_10362);
or U11939 (N_11939,N_10779,N_10212);
nor U11940 (N_11940,N_10863,N_10753);
xor U11941 (N_11941,N_10050,N_10244);
nor U11942 (N_11942,N_10042,N_10732);
nor U11943 (N_11943,N_10485,N_10039);
or U11944 (N_11944,N_10724,N_10485);
or U11945 (N_11945,N_10594,N_10092);
or U11946 (N_11946,N_10329,N_10562);
or U11947 (N_11947,N_10384,N_10312);
xor U11948 (N_11948,N_10543,N_10776);
and U11949 (N_11949,N_10792,N_10185);
xor U11950 (N_11950,N_10216,N_10212);
nor U11951 (N_11951,N_10238,N_10768);
nand U11952 (N_11952,N_10791,N_10106);
or U11953 (N_11953,N_10512,N_10737);
nand U11954 (N_11954,N_10342,N_10810);
nor U11955 (N_11955,N_10477,N_10075);
and U11956 (N_11956,N_10031,N_10621);
and U11957 (N_11957,N_10996,N_10420);
nor U11958 (N_11958,N_10031,N_10280);
and U11959 (N_11959,N_10301,N_10281);
or U11960 (N_11960,N_10812,N_10342);
and U11961 (N_11961,N_10764,N_10859);
xor U11962 (N_11962,N_10712,N_10956);
nor U11963 (N_11963,N_10695,N_10735);
nor U11964 (N_11964,N_10674,N_10279);
or U11965 (N_11965,N_10251,N_10392);
nand U11966 (N_11966,N_10308,N_10917);
and U11967 (N_11967,N_10445,N_10391);
and U11968 (N_11968,N_10902,N_10164);
xor U11969 (N_11969,N_10398,N_10298);
nand U11970 (N_11970,N_10791,N_10896);
xor U11971 (N_11971,N_10007,N_10724);
nand U11972 (N_11972,N_10642,N_10583);
nor U11973 (N_11973,N_10114,N_10665);
xor U11974 (N_11974,N_10515,N_10731);
or U11975 (N_11975,N_10801,N_10381);
and U11976 (N_11976,N_10142,N_10846);
and U11977 (N_11977,N_10265,N_10461);
and U11978 (N_11978,N_10326,N_10883);
xnor U11979 (N_11979,N_10044,N_10950);
nor U11980 (N_11980,N_10746,N_10239);
and U11981 (N_11981,N_10207,N_10310);
xor U11982 (N_11982,N_10067,N_10307);
or U11983 (N_11983,N_10823,N_10576);
xor U11984 (N_11984,N_10024,N_10882);
and U11985 (N_11985,N_10527,N_10898);
nand U11986 (N_11986,N_10797,N_10765);
nand U11987 (N_11987,N_10789,N_10575);
and U11988 (N_11988,N_10879,N_10607);
and U11989 (N_11989,N_10768,N_10863);
nand U11990 (N_11990,N_10249,N_10102);
or U11991 (N_11991,N_10564,N_10608);
nor U11992 (N_11992,N_10417,N_10387);
nor U11993 (N_11993,N_10645,N_10387);
or U11994 (N_11994,N_10972,N_10103);
and U11995 (N_11995,N_10467,N_10327);
nand U11996 (N_11996,N_10633,N_10048);
nor U11997 (N_11997,N_10610,N_10314);
and U11998 (N_11998,N_10212,N_10949);
nor U11999 (N_11999,N_10076,N_10903);
and U12000 (N_12000,N_11574,N_11326);
and U12001 (N_12001,N_11414,N_11290);
xnor U12002 (N_12002,N_11753,N_11083);
nor U12003 (N_12003,N_11171,N_11208);
xor U12004 (N_12004,N_11277,N_11148);
nand U12005 (N_12005,N_11296,N_11346);
xnor U12006 (N_12006,N_11144,N_11614);
nand U12007 (N_12007,N_11065,N_11402);
nor U12008 (N_12008,N_11023,N_11983);
and U12009 (N_12009,N_11192,N_11300);
nor U12010 (N_12010,N_11980,N_11339);
xnor U12011 (N_12011,N_11348,N_11123);
nand U12012 (N_12012,N_11774,N_11587);
nand U12013 (N_12013,N_11447,N_11384);
or U12014 (N_12014,N_11316,N_11270);
or U12015 (N_12015,N_11230,N_11837);
nand U12016 (N_12016,N_11871,N_11040);
nor U12017 (N_12017,N_11498,N_11616);
xnor U12018 (N_12018,N_11762,N_11379);
xnor U12019 (N_12019,N_11454,N_11882);
or U12020 (N_12020,N_11780,N_11553);
nor U12021 (N_12021,N_11904,N_11131);
or U12022 (N_12022,N_11631,N_11404);
nand U12023 (N_12023,N_11403,N_11480);
nor U12024 (N_12024,N_11242,N_11071);
xor U12025 (N_12025,N_11645,N_11347);
nor U12026 (N_12026,N_11662,N_11199);
nand U12027 (N_12027,N_11126,N_11118);
xnor U12028 (N_12028,N_11568,N_11485);
or U12029 (N_12029,N_11566,N_11995);
nand U12030 (N_12030,N_11976,N_11799);
and U12031 (N_12031,N_11164,N_11530);
nor U12032 (N_12032,N_11932,N_11944);
nor U12033 (N_12033,N_11500,N_11696);
or U12034 (N_12034,N_11150,N_11763);
nor U12035 (N_12035,N_11926,N_11730);
and U12036 (N_12036,N_11028,N_11222);
xnor U12037 (N_12037,N_11656,N_11761);
or U12038 (N_12038,N_11130,N_11786);
nand U12039 (N_12039,N_11293,N_11271);
or U12040 (N_12040,N_11973,N_11335);
nor U12041 (N_12041,N_11776,N_11667);
nand U12042 (N_12042,N_11410,N_11582);
nand U12043 (N_12043,N_11729,N_11968);
or U12044 (N_12044,N_11427,N_11033);
or U12045 (N_12045,N_11019,N_11930);
nand U12046 (N_12046,N_11865,N_11201);
xnor U12047 (N_12047,N_11420,N_11193);
nand U12048 (N_12048,N_11880,N_11987);
and U12049 (N_12049,N_11200,N_11330);
nor U12050 (N_12050,N_11001,N_11704);
and U12051 (N_12051,N_11375,N_11114);
xor U12052 (N_12052,N_11358,N_11579);
nor U12053 (N_12053,N_11555,N_11756);
nand U12054 (N_12054,N_11661,N_11409);
nor U12055 (N_12055,N_11266,N_11363);
and U12056 (N_12056,N_11655,N_11642);
or U12057 (N_12057,N_11298,N_11121);
or U12058 (N_12058,N_11511,N_11985);
nand U12059 (N_12059,N_11981,N_11589);
xor U12060 (N_12060,N_11212,N_11840);
nor U12061 (N_12061,N_11571,N_11769);
xor U12062 (N_12062,N_11946,N_11997);
nor U12063 (N_12063,N_11135,N_11960);
xor U12064 (N_12064,N_11595,N_11464);
and U12065 (N_12065,N_11401,N_11214);
nor U12066 (N_12066,N_11385,N_11344);
nand U12067 (N_12067,N_11000,N_11870);
nor U12068 (N_12068,N_11721,N_11496);
nor U12069 (N_12069,N_11959,N_11659);
nor U12070 (N_12070,N_11239,N_11815);
or U12071 (N_12071,N_11322,N_11458);
and U12072 (N_12072,N_11842,N_11180);
nand U12073 (N_12073,N_11607,N_11216);
or U12074 (N_12074,N_11390,N_11974);
and U12075 (N_12075,N_11791,N_11839);
xnor U12076 (N_12076,N_11361,N_11098);
nor U12077 (N_12077,N_11591,N_11279);
nand U12078 (N_12078,N_11026,N_11552);
or U12079 (N_12079,N_11156,N_11615);
xor U12080 (N_12080,N_11042,N_11734);
nand U12081 (N_12081,N_11988,N_11736);
and U12082 (N_12082,N_11233,N_11707);
or U12083 (N_12083,N_11912,N_11080);
xor U12084 (N_12084,N_11773,N_11084);
xor U12085 (N_12085,N_11720,N_11977);
nor U12086 (N_12086,N_11641,N_11334);
or U12087 (N_12087,N_11961,N_11337);
xor U12088 (N_12088,N_11889,N_11857);
nor U12089 (N_12089,N_11524,N_11030);
nor U12090 (N_12090,N_11971,N_11577);
nand U12091 (N_12091,N_11318,N_11453);
xor U12092 (N_12092,N_11243,N_11754);
and U12093 (N_12093,N_11886,N_11057);
nor U12094 (N_12094,N_11867,N_11543);
nor U12095 (N_12095,N_11149,N_11016);
nor U12096 (N_12096,N_11223,N_11509);
and U12097 (N_12097,N_11991,N_11519);
and U12098 (N_12098,N_11964,N_11855);
and U12099 (N_12099,N_11706,N_11950);
xor U12100 (N_12100,N_11660,N_11467);
xor U12101 (N_12101,N_11482,N_11982);
nor U12102 (N_12102,N_11787,N_11039);
nand U12103 (N_12103,N_11087,N_11120);
nand U12104 (N_12104,N_11712,N_11072);
xor U12105 (N_12105,N_11701,N_11268);
nand U12106 (N_12106,N_11620,N_11702);
nand U12107 (N_12107,N_11726,N_11218);
and U12108 (N_12108,N_11184,N_11476);
nand U12109 (N_12109,N_11021,N_11628);
nand U12110 (N_12110,N_11690,N_11877);
nor U12111 (N_12111,N_11378,N_11020);
and U12112 (N_12112,N_11014,N_11638);
nand U12113 (N_12113,N_11928,N_11847);
nor U12114 (N_12114,N_11481,N_11473);
xnor U12115 (N_12115,N_11554,N_11737);
nand U12116 (N_12116,N_11433,N_11687);
nor U12117 (N_12117,N_11250,N_11175);
nand U12118 (N_12118,N_11731,N_11317);
or U12119 (N_12119,N_11226,N_11611);
nand U12120 (N_12120,N_11833,N_11795);
and U12121 (N_12121,N_11813,N_11399);
xor U12122 (N_12122,N_11510,N_11297);
nor U12123 (N_12123,N_11863,N_11394);
xnor U12124 (N_12124,N_11542,N_11006);
xnor U12125 (N_12125,N_11958,N_11758);
and U12126 (N_12126,N_11292,N_11342);
xor U12127 (N_12127,N_11527,N_11247);
nand U12128 (N_12128,N_11206,N_11858);
or U12129 (N_12129,N_11508,N_11122);
xor U12130 (N_12130,N_11419,N_11516);
nor U12131 (N_12131,N_11597,N_11738);
nor U12132 (N_12132,N_11281,N_11058);
nor U12133 (N_12133,N_11933,N_11967);
and U12134 (N_12134,N_11418,N_11260);
xor U12135 (N_12135,N_11760,N_11764);
nand U12136 (N_12136,N_11691,N_11008);
nor U12137 (N_12137,N_11949,N_11700);
xor U12138 (N_12138,N_11142,N_11003);
nor U12139 (N_12139,N_11015,N_11190);
nand U12140 (N_12140,N_11658,N_11816);
nand U12141 (N_12141,N_11416,N_11986);
xor U12142 (N_12142,N_11106,N_11422);
or U12143 (N_12143,N_11470,N_11565);
and U12144 (N_12144,N_11392,N_11942);
xor U12145 (N_12145,N_11103,N_11562);
nor U12146 (N_12146,N_11538,N_11365);
and U12147 (N_12147,N_11274,N_11531);
xor U12148 (N_12148,N_11695,N_11407);
nand U12149 (N_12149,N_11452,N_11547);
and U12150 (N_12150,N_11803,N_11514);
nor U12151 (N_12151,N_11793,N_11829);
or U12152 (N_12152,N_11817,N_11520);
or U12153 (N_12153,N_11862,N_11424);
nor U12154 (N_12154,N_11188,N_11777);
and U12155 (N_12155,N_11137,N_11475);
nor U12156 (N_12156,N_11966,N_11380);
nand U12157 (N_12157,N_11640,N_11619);
and U12158 (N_12158,N_11692,N_11772);
and U12159 (N_12159,N_11902,N_11059);
xor U12160 (N_12160,N_11654,N_11258);
nand U12161 (N_12161,N_11366,N_11421);
nor U12162 (N_12162,N_11256,N_11569);
nor U12163 (N_12163,N_11234,N_11609);
nor U12164 (N_12164,N_11309,N_11903);
nand U12165 (N_12165,N_11826,N_11602);
or U12166 (N_12166,N_11089,N_11489);
nor U12167 (N_12167,N_11082,N_11618);
and U12168 (N_12168,N_11592,N_11727);
nand U12169 (N_12169,N_11127,N_11096);
nand U12170 (N_12170,N_11189,N_11693);
xnor U12171 (N_12171,N_11885,N_11672);
nand U12172 (N_12172,N_11545,N_11231);
or U12173 (N_12173,N_11580,N_11617);
xnor U12174 (N_12174,N_11905,N_11235);
xnor U12175 (N_12175,N_11417,N_11610);
nand U12176 (N_12176,N_11431,N_11170);
or U12177 (N_12177,N_11504,N_11451);
nor U12178 (N_12178,N_11755,N_11133);
and U12179 (N_12179,N_11722,N_11283);
nor U12180 (N_12180,N_11563,N_11539);
xor U12181 (N_12181,N_11415,N_11457);
xor U12182 (N_12182,N_11989,N_11836);
or U12183 (N_12183,N_11713,N_11675);
xnor U12184 (N_12184,N_11469,N_11110);
and U12185 (N_12185,N_11099,N_11918);
and U12186 (N_12186,N_11934,N_11368);
xor U12187 (N_12187,N_11748,N_11370);
and U12188 (N_12188,N_11733,N_11167);
or U12189 (N_12189,N_11732,N_11939);
nor U12190 (N_12190,N_11820,N_11446);
nand U12191 (N_12191,N_11129,N_11338);
xor U12192 (N_12192,N_11109,N_11558);
nor U12193 (N_12193,N_11113,N_11472);
nand U12194 (N_12194,N_11411,N_11389);
nand U12195 (N_12195,N_11800,N_11124);
xor U12196 (N_12196,N_11490,N_11305);
xor U12197 (N_12197,N_11246,N_11581);
and U12198 (N_12198,N_11479,N_11864);
nand U12199 (N_12199,N_11350,N_11507);
nand U12200 (N_12200,N_11328,N_11079);
nand U12201 (N_12201,N_11158,N_11078);
xor U12202 (N_12202,N_11278,N_11797);
and U12203 (N_12203,N_11757,N_11116);
nor U12204 (N_12204,N_11187,N_11854);
or U12205 (N_12205,N_11186,N_11845);
nor U12206 (N_12206,N_11025,N_11567);
and U12207 (N_12207,N_11302,N_11630);
nand U12208 (N_12208,N_11360,N_11887);
xnor U12209 (N_12209,N_11273,N_11583);
nand U12210 (N_12210,N_11502,N_11573);
xor U12211 (N_12211,N_11790,N_11801);
nor U12212 (N_12212,N_11998,N_11821);
xnor U12213 (N_12213,N_11436,N_11090);
xnor U12214 (N_12214,N_11697,N_11670);
nor U12215 (N_12215,N_11698,N_11978);
or U12216 (N_12216,N_11049,N_11515);
nand U12217 (N_12217,N_11907,N_11434);
nor U12218 (N_12218,N_11248,N_11115);
nand U12219 (N_12219,N_11924,N_11911);
nor U12220 (N_12220,N_11413,N_11092);
and U12221 (N_12221,N_11004,N_11210);
and U12222 (N_12222,N_11371,N_11564);
and U12223 (N_12223,N_11285,N_11051);
nor U12224 (N_12224,N_11428,N_11232);
nand U12225 (N_12225,N_11532,N_11091);
nor U12226 (N_12226,N_11612,N_11228);
nand U12227 (N_12227,N_11657,N_11606);
nand U12228 (N_12228,N_11276,N_11299);
or U12229 (N_12229,N_11941,N_11750);
nand U12230 (N_12230,N_11220,N_11443);
and U12231 (N_12231,N_11017,N_11398);
xnor U12232 (N_12232,N_11493,N_11173);
and U12233 (N_12233,N_11994,N_11779);
nor U12234 (N_12234,N_11892,N_11373);
xnor U12235 (N_12235,N_11391,N_11537);
or U12236 (N_12236,N_11824,N_11007);
or U12237 (N_12237,N_11364,N_11157);
or U12238 (N_12238,N_11102,N_11805);
nor U12239 (N_12239,N_11310,N_11975);
or U12240 (N_12240,N_11831,N_11094);
or U12241 (N_12241,N_11703,N_11681);
nor U12242 (N_12242,N_11354,N_11775);
or U12243 (N_12243,N_11352,N_11533);
nand U12244 (N_12244,N_11637,N_11341);
or U12245 (N_12245,N_11425,N_11455);
or U12246 (N_12246,N_11717,N_11688);
and U12247 (N_12247,N_11913,N_11217);
or U12248 (N_12248,N_11497,N_11202);
nand U12249 (N_12249,N_11584,N_11965);
xnor U12250 (N_12250,N_11107,N_11355);
or U12251 (N_12251,N_11860,N_11888);
or U12252 (N_12252,N_11408,N_11321);
nor U12253 (N_12253,N_11719,N_11312);
and U12254 (N_12254,N_11183,N_11644);
or U12255 (N_12255,N_11062,N_11287);
nor U12256 (N_12256,N_11957,N_11244);
xor U12257 (N_12257,N_11909,N_11623);
xor U12258 (N_12258,N_11128,N_11073);
xnor U12259 (N_12259,N_11935,N_11255);
nor U12260 (N_12260,N_11570,N_11848);
xnor U12261 (N_12261,N_11132,N_11807);
nand U12262 (N_12262,N_11396,N_11176);
or U12263 (N_12263,N_11027,N_11329);
nand U12264 (N_12264,N_11916,N_11383);
or U12265 (N_12265,N_11055,N_11604);
nand U12266 (N_12266,N_11856,N_11809);
or U12267 (N_12267,N_11557,N_11125);
and U12268 (N_12268,N_11593,N_11471);
nor U12269 (N_12269,N_11353,N_11046);
nand U12270 (N_12270,N_11747,N_11869);
and U12271 (N_12271,N_11075,N_11134);
or U12272 (N_12272,N_11307,N_11561);
xor U12273 (N_12273,N_11922,N_11386);
xor U12274 (N_12274,N_11632,N_11314);
nand U12275 (N_12275,N_11685,N_11303);
nand U12276 (N_12276,N_11331,N_11600);
xnor U12277 (N_12277,N_11884,N_11653);
xnor U12278 (N_12278,N_11311,N_11362);
and U12279 (N_12279,N_11254,N_11548);
nor U12280 (N_12280,N_11919,N_11518);
xor U12281 (N_12281,N_11034,N_11136);
xnor U12282 (N_12282,N_11229,N_11387);
and U12283 (N_12283,N_11621,N_11647);
xnor U12284 (N_12284,N_11716,N_11851);
or U12285 (N_12285,N_11324,N_11032);
xnor U12286 (N_12286,N_11172,N_11970);
xor U12287 (N_12287,N_11241,N_11859);
xor U12288 (N_12288,N_11332,N_11723);
nor U12289 (N_12289,N_11327,N_11474);
xnor U12290 (N_12290,N_11048,N_11449);
xor U12291 (N_12291,N_11576,N_11501);
nor U12292 (N_12292,N_11100,N_11900);
nand U12293 (N_12293,N_11556,N_11203);
nand U12294 (N_12294,N_11728,N_11683);
or U12295 (N_12295,N_11639,N_11890);
xnor U12296 (N_12296,N_11437,N_11767);
nor U12297 (N_12297,N_11969,N_11450);
and U12298 (N_12298,N_11225,N_11286);
or U12299 (N_12299,N_11992,N_11038);
or U12300 (N_12300,N_11036,N_11677);
nand U12301 (N_12301,N_11770,N_11765);
and U12302 (N_12302,N_11468,N_11929);
xor U12303 (N_12303,N_11705,N_11104);
nor U12304 (N_12304,N_11323,N_11112);
xor U12305 (N_12305,N_11506,N_11315);
nand U12306 (N_12306,N_11633,N_11798);
and U12307 (N_12307,N_11282,N_11560);
nand U12308 (N_12308,N_11393,N_11466);
and U12309 (N_12309,N_11938,N_11671);
nand U12310 (N_12310,N_11893,N_11465);
xor U12311 (N_12311,N_11117,N_11359);
nand U12312 (N_12312,N_11435,N_11674);
and U12313 (N_12313,N_11304,N_11517);
nor U12314 (N_12314,N_11406,N_11914);
xor U12315 (N_12315,N_11525,N_11009);
and U12316 (N_12316,N_11979,N_11605);
nand U12317 (N_12317,N_11990,N_11669);
nand U12318 (N_12318,N_11955,N_11138);
xor U12319 (N_12319,N_11146,N_11010);
nor U12320 (N_12320,N_11682,N_11325);
xor U12321 (N_12321,N_11054,N_11784);
and U12322 (N_12322,N_11711,N_11588);
or U12323 (N_12323,N_11011,N_11252);
nand U12324 (N_12324,N_11503,N_11781);
or U12325 (N_12325,N_11262,N_11578);
nor U12326 (N_12326,N_11908,N_11650);
nor U12327 (N_12327,N_11219,N_11745);
nand U12328 (N_12328,N_11207,N_11369);
and U12329 (N_12329,N_11710,N_11740);
xor U12330 (N_12330,N_11830,N_11012);
nor U12331 (N_12331,N_11676,N_11374);
and U12332 (N_12332,N_11636,N_11744);
nand U12333 (N_12333,N_11625,N_11838);
nor U12334 (N_12334,N_11603,N_11185);
xnor U12335 (N_12335,N_11742,N_11541);
nor U12336 (N_12336,N_11843,N_11161);
and U12337 (N_12337,N_11461,N_11269);
or U12338 (N_12338,N_11061,N_11725);
and U12339 (N_12339,N_11253,N_11868);
or U12340 (N_12340,N_11491,N_11601);
and U12341 (N_12341,N_11095,N_11195);
nand U12342 (N_12342,N_11267,N_11288);
nand U12343 (N_12343,N_11648,N_11812);
or U12344 (N_12344,N_11108,N_11984);
nor U12345 (N_12345,N_11251,N_11818);
nand U12346 (N_12346,N_11846,N_11351);
nor U12347 (N_12347,N_11213,N_11943);
and U12348 (N_12348,N_11412,N_11035);
xor U12349 (N_12349,N_11689,N_11724);
nor U12350 (N_12350,N_11512,N_11444);
or U12351 (N_12351,N_11272,N_11849);
xor U12352 (N_12352,N_11626,N_11897);
or U12353 (N_12353,N_11739,N_11484);
nand U12354 (N_12354,N_11684,N_11013);
xor U12355 (N_12355,N_11629,N_11694);
nor U12356 (N_12356,N_11405,N_11395);
and U12357 (N_12357,N_11499,N_11521);
nand U12358 (N_12358,N_11295,N_11111);
nor U12359 (N_12359,N_11177,N_11896);
nand U12360 (N_12360,N_11819,N_11627);
and U12361 (N_12361,N_11093,N_11381);
or U12362 (N_12362,N_11492,N_11624);
or U12363 (N_12363,N_11037,N_11536);
nor U12364 (N_12364,N_11487,N_11320);
and U12365 (N_12365,N_11852,N_11333);
and U12366 (N_12366,N_11044,N_11486);
nor U12367 (N_12367,N_11196,N_11261);
nand U12368 (N_12368,N_11768,N_11382);
and U12369 (N_12369,N_11162,N_11160);
or U12370 (N_12370,N_11613,N_11460);
and U12371 (N_12371,N_11179,N_11962);
nor U12372 (N_12372,N_11047,N_11679);
nand U12373 (N_12373,N_11069,N_11792);
or U12374 (N_12374,N_11154,N_11634);
or U12375 (N_12375,N_11463,N_11878);
nand U12376 (N_12376,N_11349,N_11590);
nand U12377 (N_12377,N_11372,N_11874);
or U12378 (N_12378,N_11822,N_11459);
or U12379 (N_12379,N_11445,N_11649);
nor U12380 (N_12380,N_11952,N_11249);
xor U12381 (N_12381,N_11528,N_11191);
and U12382 (N_12382,N_11551,N_11081);
xnor U12383 (N_12383,N_11477,N_11766);
or U12384 (N_12384,N_11174,N_11280);
or U12385 (N_12385,N_11238,N_11544);
xnor U12386 (N_12386,N_11635,N_11686);
nor U12387 (N_12387,N_11357,N_11070);
and U12388 (N_12388,N_11945,N_11523);
xnor U12389 (N_12389,N_11743,N_11917);
xor U12390 (N_12390,N_11204,N_11906);
xnor U12391 (N_12391,N_11876,N_11529);
xnor U12392 (N_12392,N_11439,N_11088);
nor U12393 (N_12393,N_11708,N_11872);
and U12394 (N_12394,N_11925,N_11522);
nand U12395 (N_12395,N_11844,N_11221);
and U12396 (N_12396,N_11651,N_11963);
and U12397 (N_12397,N_11198,N_11294);
xor U12398 (N_12398,N_11211,N_11153);
or U12399 (N_12399,N_11056,N_11841);
nor U12400 (N_12400,N_11953,N_11972);
nor U12401 (N_12401,N_11931,N_11151);
xor U12402 (N_12402,N_11746,N_11598);
and U12403 (N_12403,N_11478,N_11834);
nor U12404 (N_12404,N_11018,N_11181);
nand U12405 (N_12405,N_11308,N_11002);
and U12406 (N_12406,N_11060,N_11827);
and U12407 (N_12407,N_11388,N_11993);
or U12408 (N_12408,N_11168,N_11076);
xnor U12409 (N_12409,N_11147,N_11263);
xor U12410 (N_12410,N_11927,N_11540);
and U12411 (N_12411,N_11665,N_11343);
or U12412 (N_12412,N_11883,N_11031);
nand U12413 (N_12413,N_11194,N_11064);
nor U12414 (N_12414,N_11257,N_11715);
xnor U12415 (N_12415,N_11549,N_11430);
nand U12416 (N_12416,N_11067,N_11178);
xor U12417 (N_12417,N_11789,N_11714);
xor U12418 (N_12418,N_11513,N_11954);
nor U12419 (N_12419,N_11879,N_11948);
and U12420 (N_12420,N_11155,N_11891);
xor U12421 (N_12421,N_11999,N_11397);
and U12422 (N_12422,N_11456,N_11227);
nand U12423 (N_12423,N_11377,N_11442);
and U12424 (N_12424,N_11426,N_11356);
nand U12425 (N_12425,N_11313,N_11245);
nand U12426 (N_12426,N_11159,N_11101);
xor U12427 (N_12427,N_11825,N_11275);
nor U12428 (N_12428,N_11041,N_11236);
nor U12429 (N_12429,N_11759,N_11205);
or U12430 (N_12430,N_11483,N_11495);
and U12431 (N_12431,N_11599,N_11169);
and U12432 (N_12432,N_11345,N_11749);
nand U12433 (N_12433,N_11259,N_11423);
nand U12434 (N_12434,N_11646,N_11488);
or U12435 (N_12435,N_11673,N_11086);
xor U12436 (N_12436,N_11119,N_11505);
nand U12437 (N_12437,N_11105,N_11319);
or U12438 (N_12438,N_11853,N_11145);
nor U12439 (N_12439,N_11264,N_11828);
nand U12440 (N_12440,N_11050,N_11141);
nand U12441 (N_12441,N_11866,N_11546);
and U12442 (N_12442,N_11718,N_11622);
and U12443 (N_12443,N_11996,N_11778);
and U12444 (N_12444,N_11209,N_11899);
and U12445 (N_12445,N_11265,N_11921);
and U12446 (N_12446,N_11240,N_11139);
xor U12447 (N_12447,N_11284,N_11910);
or U12448 (N_12448,N_11771,N_11794);
nand U12449 (N_12449,N_11940,N_11166);
xor U12450 (N_12450,N_11875,N_11752);
or U12451 (N_12451,N_11663,N_11894);
xnor U12452 (N_12452,N_11895,N_11596);
nor U12453 (N_12453,N_11143,N_11215);
nand U12454 (N_12454,N_11559,N_11400);
or U12455 (N_12455,N_11575,N_11898);
nor U12456 (N_12456,N_11526,N_11448);
nor U12457 (N_12457,N_11811,N_11237);
nand U12458 (N_12458,N_11005,N_11751);
nand U12459 (N_12459,N_11594,N_11045);
xor U12460 (N_12460,N_11783,N_11097);
xor U12461 (N_12461,N_11956,N_11785);
and U12462 (N_12462,N_11861,N_11814);
and U12463 (N_12463,N_11668,N_11915);
nand U12464 (N_12464,N_11741,N_11022);
and U12465 (N_12465,N_11462,N_11666);
xnor U12466 (N_12466,N_11336,N_11951);
nor U12467 (N_12467,N_11306,N_11832);
xor U12468 (N_12468,N_11152,N_11053);
xnor U12469 (N_12469,N_11936,N_11802);
or U12470 (N_12470,N_11163,N_11782);
nor U12471 (N_12471,N_11534,N_11224);
nor U12472 (N_12472,N_11550,N_11881);
nor U12473 (N_12473,N_11835,N_11140);
and U12474 (N_12474,N_11901,N_11438);
nor U12475 (N_12475,N_11586,N_11029);
or U12476 (N_12476,N_11796,N_11923);
and U12477 (N_12477,N_11085,N_11804);
nor U12478 (N_12478,N_11585,N_11806);
and U12479 (N_12479,N_11165,N_11494);
and U12480 (N_12480,N_11664,N_11074);
and U12481 (N_12481,N_11810,N_11788);
xor U12482 (N_12482,N_11024,N_11699);
xor U12483 (N_12483,N_11652,N_11920);
nand U12484 (N_12484,N_11052,N_11043);
nor U12485 (N_12485,N_11873,N_11678);
nor U12486 (N_12486,N_11441,N_11535);
nor U12487 (N_12487,N_11289,N_11077);
nand U12488 (N_12488,N_11735,N_11301);
xnor U12489 (N_12489,N_11608,N_11440);
nand U12490 (N_12490,N_11367,N_11808);
nand U12491 (N_12491,N_11066,N_11643);
xor U12492 (N_12492,N_11182,N_11937);
or U12493 (N_12493,N_11197,N_11947);
nand U12494 (N_12494,N_11709,N_11850);
or U12495 (N_12495,N_11291,N_11572);
xnor U12496 (N_12496,N_11680,N_11068);
nor U12497 (N_12497,N_11432,N_11340);
or U12498 (N_12498,N_11823,N_11063);
and U12499 (N_12499,N_11429,N_11376);
and U12500 (N_12500,N_11507,N_11590);
nand U12501 (N_12501,N_11468,N_11337);
nand U12502 (N_12502,N_11818,N_11699);
xor U12503 (N_12503,N_11917,N_11429);
or U12504 (N_12504,N_11961,N_11949);
xnor U12505 (N_12505,N_11273,N_11913);
and U12506 (N_12506,N_11642,N_11698);
xor U12507 (N_12507,N_11326,N_11843);
or U12508 (N_12508,N_11306,N_11304);
nor U12509 (N_12509,N_11056,N_11688);
or U12510 (N_12510,N_11159,N_11154);
xor U12511 (N_12511,N_11165,N_11719);
nor U12512 (N_12512,N_11734,N_11405);
nor U12513 (N_12513,N_11264,N_11347);
and U12514 (N_12514,N_11467,N_11728);
nand U12515 (N_12515,N_11486,N_11375);
xor U12516 (N_12516,N_11275,N_11223);
xor U12517 (N_12517,N_11079,N_11250);
nor U12518 (N_12518,N_11162,N_11888);
or U12519 (N_12519,N_11404,N_11863);
and U12520 (N_12520,N_11996,N_11625);
and U12521 (N_12521,N_11100,N_11133);
and U12522 (N_12522,N_11290,N_11122);
or U12523 (N_12523,N_11946,N_11934);
and U12524 (N_12524,N_11713,N_11479);
or U12525 (N_12525,N_11274,N_11896);
nor U12526 (N_12526,N_11965,N_11867);
xnor U12527 (N_12527,N_11406,N_11869);
or U12528 (N_12528,N_11925,N_11266);
nand U12529 (N_12529,N_11860,N_11641);
nor U12530 (N_12530,N_11087,N_11576);
nor U12531 (N_12531,N_11577,N_11918);
nor U12532 (N_12532,N_11547,N_11026);
or U12533 (N_12533,N_11172,N_11784);
nor U12534 (N_12534,N_11737,N_11629);
nor U12535 (N_12535,N_11311,N_11823);
nor U12536 (N_12536,N_11767,N_11818);
xor U12537 (N_12537,N_11001,N_11657);
or U12538 (N_12538,N_11734,N_11000);
nand U12539 (N_12539,N_11073,N_11380);
xor U12540 (N_12540,N_11003,N_11100);
nand U12541 (N_12541,N_11166,N_11325);
nor U12542 (N_12542,N_11042,N_11897);
nand U12543 (N_12543,N_11579,N_11759);
and U12544 (N_12544,N_11786,N_11513);
and U12545 (N_12545,N_11332,N_11752);
nor U12546 (N_12546,N_11130,N_11306);
xor U12547 (N_12547,N_11496,N_11268);
nor U12548 (N_12548,N_11994,N_11709);
xnor U12549 (N_12549,N_11750,N_11949);
nand U12550 (N_12550,N_11630,N_11602);
nand U12551 (N_12551,N_11768,N_11817);
and U12552 (N_12552,N_11225,N_11269);
and U12553 (N_12553,N_11660,N_11517);
or U12554 (N_12554,N_11443,N_11224);
nand U12555 (N_12555,N_11067,N_11060);
and U12556 (N_12556,N_11501,N_11198);
xor U12557 (N_12557,N_11433,N_11172);
xnor U12558 (N_12558,N_11148,N_11963);
nor U12559 (N_12559,N_11838,N_11557);
nand U12560 (N_12560,N_11935,N_11633);
or U12561 (N_12561,N_11613,N_11872);
nand U12562 (N_12562,N_11248,N_11703);
or U12563 (N_12563,N_11902,N_11201);
nand U12564 (N_12564,N_11098,N_11945);
or U12565 (N_12565,N_11117,N_11980);
or U12566 (N_12566,N_11397,N_11055);
nand U12567 (N_12567,N_11001,N_11133);
nand U12568 (N_12568,N_11484,N_11374);
nand U12569 (N_12569,N_11972,N_11304);
xnor U12570 (N_12570,N_11506,N_11254);
and U12571 (N_12571,N_11768,N_11904);
nand U12572 (N_12572,N_11169,N_11503);
nor U12573 (N_12573,N_11082,N_11210);
nor U12574 (N_12574,N_11262,N_11293);
and U12575 (N_12575,N_11235,N_11944);
nand U12576 (N_12576,N_11348,N_11231);
and U12577 (N_12577,N_11380,N_11580);
nor U12578 (N_12578,N_11834,N_11856);
and U12579 (N_12579,N_11574,N_11009);
nand U12580 (N_12580,N_11057,N_11808);
and U12581 (N_12581,N_11973,N_11076);
nor U12582 (N_12582,N_11323,N_11580);
nand U12583 (N_12583,N_11394,N_11425);
nor U12584 (N_12584,N_11999,N_11421);
nand U12585 (N_12585,N_11175,N_11636);
xnor U12586 (N_12586,N_11278,N_11117);
nor U12587 (N_12587,N_11423,N_11691);
xnor U12588 (N_12588,N_11334,N_11610);
nor U12589 (N_12589,N_11849,N_11634);
xor U12590 (N_12590,N_11487,N_11152);
nor U12591 (N_12591,N_11833,N_11166);
and U12592 (N_12592,N_11831,N_11723);
xnor U12593 (N_12593,N_11646,N_11734);
nand U12594 (N_12594,N_11830,N_11522);
or U12595 (N_12595,N_11733,N_11286);
nand U12596 (N_12596,N_11972,N_11802);
nor U12597 (N_12597,N_11608,N_11780);
or U12598 (N_12598,N_11567,N_11548);
xor U12599 (N_12599,N_11599,N_11916);
or U12600 (N_12600,N_11378,N_11821);
xor U12601 (N_12601,N_11730,N_11552);
nor U12602 (N_12602,N_11060,N_11692);
nand U12603 (N_12603,N_11031,N_11729);
or U12604 (N_12604,N_11080,N_11943);
or U12605 (N_12605,N_11956,N_11541);
and U12606 (N_12606,N_11082,N_11790);
nor U12607 (N_12607,N_11634,N_11069);
xnor U12608 (N_12608,N_11151,N_11163);
nand U12609 (N_12609,N_11497,N_11663);
nand U12610 (N_12610,N_11090,N_11897);
and U12611 (N_12611,N_11089,N_11886);
nor U12612 (N_12612,N_11514,N_11652);
xor U12613 (N_12613,N_11700,N_11473);
nor U12614 (N_12614,N_11993,N_11434);
nand U12615 (N_12615,N_11641,N_11423);
and U12616 (N_12616,N_11982,N_11851);
nor U12617 (N_12617,N_11234,N_11113);
and U12618 (N_12618,N_11932,N_11697);
and U12619 (N_12619,N_11383,N_11283);
nor U12620 (N_12620,N_11155,N_11011);
nor U12621 (N_12621,N_11183,N_11939);
nor U12622 (N_12622,N_11726,N_11938);
or U12623 (N_12623,N_11447,N_11035);
and U12624 (N_12624,N_11489,N_11301);
or U12625 (N_12625,N_11866,N_11178);
and U12626 (N_12626,N_11825,N_11077);
and U12627 (N_12627,N_11472,N_11842);
and U12628 (N_12628,N_11966,N_11671);
nand U12629 (N_12629,N_11135,N_11170);
or U12630 (N_12630,N_11067,N_11235);
nor U12631 (N_12631,N_11434,N_11575);
xor U12632 (N_12632,N_11624,N_11071);
or U12633 (N_12633,N_11511,N_11168);
or U12634 (N_12634,N_11199,N_11718);
nand U12635 (N_12635,N_11804,N_11262);
nand U12636 (N_12636,N_11021,N_11260);
xnor U12637 (N_12637,N_11202,N_11939);
and U12638 (N_12638,N_11935,N_11917);
and U12639 (N_12639,N_11788,N_11360);
nand U12640 (N_12640,N_11193,N_11979);
nor U12641 (N_12641,N_11919,N_11480);
xnor U12642 (N_12642,N_11455,N_11305);
nand U12643 (N_12643,N_11986,N_11256);
nor U12644 (N_12644,N_11439,N_11651);
xnor U12645 (N_12645,N_11720,N_11294);
nand U12646 (N_12646,N_11820,N_11398);
or U12647 (N_12647,N_11924,N_11767);
xor U12648 (N_12648,N_11262,N_11292);
and U12649 (N_12649,N_11100,N_11749);
or U12650 (N_12650,N_11192,N_11506);
xnor U12651 (N_12651,N_11931,N_11158);
or U12652 (N_12652,N_11544,N_11298);
xor U12653 (N_12653,N_11702,N_11965);
xor U12654 (N_12654,N_11532,N_11376);
nand U12655 (N_12655,N_11380,N_11121);
xor U12656 (N_12656,N_11391,N_11775);
nor U12657 (N_12657,N_11668,N_11731);
or U12658 (N_12658,N_11539,N_11842);
nand U12659 (N_12659,N_11574,N_11633);
or U12660 (N_12660,N_11142,N_11679);
nor U12661 (N_12661,N_11705,N_11503);
nor U12662 (N_12662,N_11515,N_11217);
xor U12663 (N_12663,N_11182,N_11796);
and U12664 (N_12664,N_11586,N_11523);
and U12665 (N_12665,N_11172,N_11055);
or U12666 (N_12666,N_11001,N_11947);
nor U12667 (N_12667,N_11925,N_11840);
xnor U12668 (N_12668,N_11647,N_11952);
xnor U12669 (N_12669,N_11063,N_11179);
xnor U12670 (N_12670,N_11428,N_11644);
xor U12671 (N_12671,N_11213,N_11043);
or U12672 (N_12672,N_11020,N_11337);
or U12673 (N_12673,N_11488,N_11873);
or U12674 (N_12674,N_11735,N_11083);
nor U12675 (N_12675,N_11620,N_11974);
xnor U12676 (N_12676,N_11458,N_11451);
and U12677 (N_12677,N_11863,N_11731);
xnor U12678 (N_12678,N_11182,N_11493);
nand U12679 (N_12679,N_11281,N_11596);
or U12680 (N_12680,N_11051,N_11410);
nand U12681 (N_12681,N_11124,N_11074);
and U12682 (N_12682,N_11998,N_11117);
and U12683 (N_12683,N_11759,N_11245);
xnor U12684 (N_12684,N_11697,N_11975);
and U12685 (N_12685,N_11147,N_11886);
xnor U12686 (N_12686,N_11657,N_11854);
nand U12687 (N_12687,N_11512,N_11740);
nand U12688 (N_12688,N_11590,N_11671);
xnor U12689 (N_12689,N_11980,N_11741);
or U12690 (N_12690,N_11740,N_11283);
or U12691 (N_12691,N_11541,N_11299);
nand U12692 (N_12692,N_11035,N_11026);
or U12693 (N_12693,N_11559,N_11622);
nor U12694 (N_12694,N_11200,N_11210);
xnor U12695 (N_12695,N_11860,N_11718);
or U12696 (N_12696,N_11406,N_11870);
or U12697 (N_12697,N_11787,N_11043);
and U12698 (N_12698,N_11236,N_11203);
xor U12699 (N_12699,N_11257,N_11433);
or U12700 (N_12700,N_11901,N_11559);
or U12701 (N_12701,N_11053,N_11162);
or U12702 (N_12702,N_11294,N_11269);
nor U12703 (N_12703,N_11012,N_11443);
nor U12704 (N_12704,N_11192,N_11605);
and U12705 (N_12705,N_11207,N_11609);
and U12706 (N_12706,N_11231,N_11162);
nor U12707 (N_12707,N_11819,N_11267);
or U12708 (N_12708,N_11058,N_11663);
nand U12709 (N_12709,N_11934,N_11187);
nor U12710 (N_12710,N_11578,N_11701);
xor U12711 (N_12711,N_11587,N_11755);
nand U12712 (N_12712,N_11472,N_11765);
or U12713 (N_12713,N_11154,N_11863);
nor U12714 (N_12714,N_11914,N_11021);
nand U12715 (N_12715,N_11687,N_11836);
nand U12716 (N_12716,N_11597,N_11324);
nor U12717 (N_12717,N_11616,N_11334);
nor U12718 (N_12718,N_11328,N_11037);
nand U12719 (N_12719,N_11101,N_11347);
nor U12720 (N_12720,N_11617,N_11210);
nand U12721 (N_12721,N_11586,N_11934);
and U12722 (N_12722,N_11154,N_11354);
nor U12723 (N_12723,N_11218,N_11190);
nand U12724 (N_12724,N_11079,N_11605);
nor U12725 (N_12725,N_11215,N_11338);
nor U12726 (N_12726,N_11625,N_11874);
or U12727 (N_12727,N_11173,N_11803);
xor U12728 (N_12728,N_11644,N_11856);
and U12729 (N_12729,N_11674,N_11398);
xnor U12730 (N_12730,N_11497,N_11397);
nand U12731 (N_12731,N_11990,N_11417);
and U12732 (N_12732,N_11863,N_11153);
nor U12733 (N_12733,N_11726,N_11545);
nor U12734 (N_12734,N_11710,N_11845);
and U12735 (N_12735,N_11738,N_11113);
nor U12736 (N_12736,N_11488,N_11198);
nor U12737 (N_12737,N_11587,N_11841);
nand U12738 (N_12738,N_11203,N_11541);
or U12739 (N_12739,N_11214,N_11544);
and U12740 (N_12740,N_11532,N_11469);
nand U12741 (N_12741,N_11528,N_11550);
nor U12742 (N_12742,N_11727,N_11559);
nand U12743 (N_12743,N_11114,N_11799);
or U12744 (N_12744,N_11199,N_11405);
and U12745 (N_12745,N_11771,N_11344);
or U12746 (N_12746,N_11971,N_11617);
xnor U12747 (N_12747,N_11367,N_11303);
nor U12748 (N_12748,N_11649,N_11965);
or U12749 (N_12749,N_11116,N_11823);
nor U12750 (N_12750,N_11856,N_11559);
nand U12751 (N_12751,N_11749,N_11476);
nand U12752 (N_12752,N_11514,N_11224);
or U12753 (N_12753,N_11817,N_11621);
nand U12754 (N_12754,N_11436,N_11729);
nand U12755 (N_12755,N_11730,N_11811);
xnor U12756 (N_12756,N_11570,N_11986);
or U12757 (N_12757,N_11357,N_11555);
and U12758 (N_12758,N_11629,N_11036);
xnor U12759 (N_12759,N_11047,N_11834);
nand U12760 (N_12760,N_11484,N_11162);
nor U12761 (N_12761,N_11809,N_11197);
nor U12762 (N_12762,N_11522,N_11405);
xor U12763 (N_12763,N_11922,N_11890);
and U12764 (N_12764,N_11256,N_11797);
xnor U12765 (N_12765,N_11440,N_11080);
or U12766 (N_12766,N_11028,N_11369);
xor U12767 (N_12767,N_11848,N_11652);
nand U12768 (N_12768,N_11749,N_11084);
nor U12769 (N_12769,N_11261,N_11864);
xor U12770 (N_12770,N_11473,N_11646);
or U12771 (N_12771,N_11093,N_11359);
nor U12772 (N_12772,N_11552,N_11160);
nor U12773 (N_12773,N_11006,N_11207);
xor U12774 (N_12774,N_11089,N_11040);
nand U12775 (N_12775,N_11355,N_11077);
xor U12776 (N_12776,N_11823,N_11441);
nand U12777 (N_12777,N_11011,N_11395);
xor U12778 (N_12778,N_11792,N_11680);
nor U12779 (N_12779,N_11867,N_11223);
or U12780 (N_12780,N_11384,N_11958);
and U12781 (N_12781,N_11467,N_11260);
and U12782 (N_12782,N_11750,N_11422);
and U12783 (N_12783,N_11695,N_11730);
and U12784 (N_12784,N_11629,N_11906);
xor U12785 (N_12785,N_11809,N_11125);
or U12786 (N_12786,N_11020,N_11865);
or U12787 (N_12787,N_11261,N_11918);
and U12788 (N_12788,N_11316,N_11619);
nand U12789 (N_12789,N_11481,N_11590);
and U12790 (N_12790,N_11119,N_11350);
and U12791 (N_12791,N_11469,N_11260);
and U12792 (N_12792,N_11528,N_11773);
nor U12793 (N_12793,N_11281,N_11731);
nor U12794 (N_12794,N_11687,N_11909);
or U12795 (N_12795,N_11970,N_11345);
xnor U12796 (N_12796,N_11066,N_11351);
and U12797 (N_12797,N_11774,N_11794);
and U12798 (N_12798,N_11032,N_11163);
xnor U12799 (N_12799,N_11566,N_11354);
nand U12800 (N_12800,N_11393,N_11825);
or U12801 (N_12801,N_11729,N_11366);
nand U12802 (N_12802,N_11646,N_11587);
or U12803 (N_12803,N_11908,N_11049);
xnor U12804 (N_12804,N_11494,N_11604);
xor U12805 (N_12805,N_11391,N_11944);
and U12806 (N_12806,N_11425,N_11445);
xor U12807 (N_12807,N_11325,N_11812);
and U12808 (N_12808,N_11476,N_11513);
nand U12809 (N_12809,N_11850,N_11482);
or U12810 (N_12810,N_11479,N_11277);
xor U12811 (N_12811,N_11567,N_11596);
or U12812 (N_12812,N_11930,N_11633);
nand U12813 (N_12813,N_11626,N_11825);
nand U12814 (N_12814,N_11602,N_11229);
or U12815 (N_12815,N_11733,N_11035);
xor U12816 (N_12816,N_11155,N_11580);
nand U12817 (N_12817,N_11458,N_11516);
xnor U12818 (N_12818,N_11894,N_11183);
nor U12819 (N_12819,N_11612,N_11241);
nor U12820 (N_12820,N_11556,N_11682);
or U12821 (N_12821,N_11799,N_11736);
xor U12822 (N_12822,N_11920,N_11907);
and U12823 (N_12823,N_11354,N_11584);
or U12824 (N_12824,N_11722,N_11357);
and U12825 (N_12825,N_11896,N_11837);
or U12826 (N_12826,N_11930,N_11912);
nand U12827 (N_12827,N_11677,N_11859);
xnor U12828 (N_12828,N_11159,N_11625);
nand U12829 (N_12829,N_11552,N_11439);
and U12830 (N_12830,N_11815,N_11041);
or U12831 (N_12831,N_11891,N_11836);
or U12832 (N_12832,N_11113,N_11432);
and U12833 (N_12833,N_11735,N_11674);
xor U12834 (N_12834,N_11680,N_11020);
xor U12835 (N_12835,N_11510,N_11191);
nand U12836 (N_12836,N_11760,N_11068);
and U12837 (N_12837,N_11691,N_11895);
or U12838 (N_12838,N_11662,N_11924);
xor U12839 (N_12839,N_11573,N_11759);
or U12840 (N_12840,N_11974,N_11292);
nand U12841 (N_12841,N_11742,N_11949);
xnor U12842 (N_12842,N_11515,N_11828);
xnor U12843 (N_12843,N_11737,N_11856);
nor U12844 (N_12844,N_11197,N_11983);
xnor U12845 (N_12845,N_11533,N_11444);
and U12846 (N_12846,N_11726,N_11506);
and U12847 (N_12847,N_11366,N_11167);
or U12848 (N_12848,N_11126,N_11779);
nor U12849 (N_12849,N_11974,N_11509);
xnor U12850 (N_12850,N_11898,N_11762);
nand U12851 (N_12851,N_11479,N_11783);
or U12852 (N_12852,N_11837,N_11271);
nor U12853 (N_12853,N_11029,N_11792);
nand U12854 (N_12854,N_11995,N_11246);
nand U12855 (N_12855,N_11258,N_11438);
and U12856 (N_12856,N_11993,N_11540);
nand U12857 (N_12857,N_11000,N_11746);
xnor U12858 (N_12858,N_11821,N_11876);
nor U12859 (N_12859,N_11970,N_11868);
or U12860 (N_12860,N_11093,N_11725);
xor U12861 (N_12861,N_11787,N_11475);
or U12862 (N_12862,N_11951,N_11581);
and U12863 (N_12863,N_11912,N_11314);
nor U12864 (N_12864,N_11297,N_11643);
or U12865 (N_12865,N_11378,N_11059);
nor U12866 (N_12866,N_11368,N_11110);
nand U12867 (N_12867,N_11287,N_11458);
or U12868 (N_12868,N_11742,N_11789);
xor U12869 (N_12869,N_11749,N_11855);
nand U12870 (N_12870,N_11761,N_11782);
nor U12871 (N_12871,N_11799,N_11422);
nand U12872 (N_12872,N_11859,N_11022);
or U12873 (N_12873,N_11544,N_11575);
or U12874 (N_12874,N_11528,N_11285);
nand U12875 (N_12875,N_11104,N_11500);
or U12876 (N_12876,N_11851,N_11915);
and U12877 (N_12877,N_11532,N_11148);
or U12878 (N_12878,N_11931,N_11480);
or U12879 (N_12879,N_11568,N_11532);
or U12880 (N_12880,N_11258,N_11210);
nor U12881 (N_12881,N_11452,N_11190);
and U12882 (N_12882,N_11350,N_11369);
and U12883 (N_12883,N_11389,N_11229);
nand U12884 (N_12884,N_11958,N_11170);
xor U12885 (N_12885,N_11176,N_11135);
nand U12886 (N_12886,N_11284,N_11325);
and U12887 (N_12887,N_11324,N_11921);
and U12888 (N_12888,N_11284,N_11823);
nand U12889 (N_12889,N_11846,N_11655);
and U12890 (N_12890,N_11248,N_11364);
and U12891 (N_12891,N_11526,N_11324);
or U12892 (N_12892,N_11991,N_11941);
xnor U12893 (N_12893,N_11779,N_11372);
xnor U12894 (N_12894,N_11264,N_11070);
nor U12895 (N_12895,N_11348,N_11785);
nand U12896 (N_12896,N_11249,N_11230);
nand U12897 (N_12897,N_11110,N_11307);
and U12898 (N_12898,N_11256,N_11798);
xor U12899 (N_12899,N_11942,N_11105);
nand U12900 (N_12900,N_11331,N_11563);
or U12901 (N_12901,N_11785,N_11668);
xnor U12902 (N_12902,N_11029,N_11498);
and U12903 (N_12903,N_11980,N_11892);
xor U12904 (N_12904,N_11421,N_11247);
or U12905 (N_12905,N_11995,N_11356);
xor U12906 (N_12906,N_11301,N_11896);
nor U12907 (N_12907,N_11657,N_11010);
or U12908 (N_12908,N_11321,N_11563);
or U12909 (N_12909,N_11263,N_11800);
and U12910 (N_12910,N_11990,N_11069);
xor U12911 (N_12911,N_11132,N_11554);
or U12912 (N_12912,N_11309,N_11476);
xnor U12913 (N_12913,N_11561,N_11425);
xor U12914 (N_12914,N_11022,N_11075);
nand U12915 (N_12915,N_11152,N_11369);
xor U12916 (N_12916,N_11319,N_11101);
and U12917 (N_12917,N_11396,N_11939);
xor U12918 (N_12918,N_11380,N_11222);
xor U12919 (N_12919,N_11228,N_11268);
xnor U12920 (N_12920,N_11263,N_11900);
nor U12921 (N_12921,N_11858,N_11779);
nor U12922 (N_12922,N_11399,N_11964);
and U12923 (N_12923,N_11742,N_11507);
or U12924 (N_12924,N_11509,N_11292);
xnor U12925 (N_12925,N_11534,N_11558);
nor U12926 (N_12926,N_11821,N_11781);
and U12927 (N_12927,N_11200,N_11074);
nor U12928 (N_12928,N_11014,N_11554);
nor U12929 (N_12929,N_11084,N_11579);
xnor U12930 (N_12930,N_11624,N_11692);
nand U12931 (N_12931,N_11505,N_11634);
nor U12932 (N_12932,N_11388,N_11191);
and U12933 (N_12933,N_11898,N_11954);
xnor U12934 (N_12934,N_11969,N_11271);
and U12935 (N_12935,N_11187,N_11308);
xnor U12936 (N_12936,N_11305,N_11763);
nand U12937 (N_12937,N_11507,N_11392);
xor U12938 (N_12938,N_11121,N_11948);
nor U12939 (N_12939,N_11313,N_11923);
nand U12940 (N_12940,N_11971,N_11740);
nand U12941 (N_12941,N_11452,N_11260);
nor U12942 (N_12942,N_11448,N_11479);
nor U12943 (N_12943,N_11493,N_11541);
or U12944 (N_12944,N_11215,N_11571);
nand U12945 (N_12945,N_11914,N_11249);
or U12946 (N_12946,N_11676,N_11381);
nor U12947 (N_12947,N_11425,N_11674);
or U12948 (N_12948,N_11600,N_11440);
nand U12949 (N_12949,N_11254,N_11352);
and U12950 (N_12950,N_11421,N_11840);
and U12951 (N_12951,N_11180,N_11862);
xor U12952 (N_12952,N_11306,N_11802);
nand U12953 (N_12953,N_11316,N_11786);
xor U12954 (N_12954,N_11120,N_11180);
or U12955 (N_12955,N_11468,N_11141);
and U12956 (N_12956,N_11013,N_11604);
and U12957 (N_12957,N_11853,N_11389);
nor U12958 (N_12958,N_11443,N_11125);
nand U12959 (N_12959,N_11055,N_11010);
and U12960 (N_12960,N_11358,N_11932);
and U12961 (N_12961,N_11610,N_11548);
nand U12962 (N_12962,N_11676,N_11500);
and U12963 (N_12963,N_11657,N_11969);
nand U12964 (N_12964,N_11506,N_11408);
nand U12965 (N_12965,N_11250,N_11226);
nor U12966 (N_12966,N_11027,N_11468);
and U12967 (N_12967,N_11370,N_11547);
or U12968 (N_12968,N_11697,N_11202);
nand U12969 (N_12969,N_11924,N_11160);
nand U12970 (N_12970,N_11813,N_11177);
xor U12971 (N_12971,N_11096,N_11374);
nand U12972 (N_12972,N_11134,N_11854);
or U12973 (N_12973,N_11438,N_11388);
nor U12974 (N_12974,N_11646,N_11708);
xnor U12975 (N_12975,N_11901,N_11132);
nor U12976 (N_12976,N_11099,N_11566);
nand U12977 (N_12977,N_11125,N_11211);
or U12978 (N_12978,N_11790,N_11862);
or U12979 (N_12979,N_11008,N_11562);
nand U12980 (N_12980,N_11529,N_11923);
nand U12981 (N_12981,N_11179,N_11197);
xnor U12982 (N_12982,N_11431,N_11905);
nand U12983 (N_12983,N_11093,N_11654);
xnor U12984 (N_12984,N_11617,N_11236);
xor U12985 (N_12985,N_11706,N_11762);
nand U12986 (N_12986,N_11156,N_11554);
and U12987 (N_12987,N_11279,N_11071);
and U12988 (N_12988,N_11211,N_11033);
nor U12989 (N_12989,N_11763,N_11787);
or U12990 (N_12990,N_11825,N_11336);
xnor U12991 (N_12991,N_11062,N_11521);
nor U12992 (N_12992,N_11572,N_11848);
nor U12993 (N_12993,N_11688,N_11085);
nand U12994 (N_12994,N_11129,N_11523);
nor U12995 (N_12995,N_11282,N_11475);
xnor U12996 (N_12996,N_11075,N_11742);
and U12997 (N_12997,N_11141,N_11582);
nor U12998 (N_12998,N_11753,N_11467);
xnor U12999 (N_12999,N_11725,N_11133);
xnor U13000 (N_13000,N_12079,N_12719);
nor U13001 (N_13001,N_12289,N_12152);
nor U13002 (N_13002,N_12860,N_12498);
xnor U13003 (N_13003,N_12159,N_12125);
nor U13004 (N_13004,N_12076,N_12505);
or U13005 (N_13005,N_12809,N_12984);
or U13006 (N_13006,N_12989,N_12141);
nor U13007 (N_13007,N_12452,N_12928);
or U13008 (N_13008,N_12113,N_12016);
and U13009 (N_13009,N_12904,N_12344);
or U13010 (N_13010,N_12957,N_12708);
nand U13011 (N_13011,N_12441,N_12245);
nand U13012 (N_13012,N_12670,N_12582);
xnor U13013 (N_13013,N_12836,N_12976);
and U13014 (N_13014,N_12037,N_12974);
xor U13015 (N_13015,N_12891,N_12806);
and U13016 (N_13016,N_12581,N_12338);
or U13017 (N_13017,N_12286,N_12366);
nand U13018 (N_13018,N_12645,N_12996);
xor U13019 (N_13019,N_12927,N_12442);
or U13020 (N_13020,N_12922,N_12781);
nand U13021 (N_13021,N_12252,N_12480);
xor U13022 (N_13022,N_12193,N_12693);
nand U13023 (N_13023,N_12622,N_12959);
and U13024 (N_13024,N_12937,N_12466);
nor U13025 (N_13025,N_12364,N_12729);
nand U13026 (N_13026,N_12420,N_12698);
nor U13027 (N_13027,N_12817,N_12110);
nor U13028 (N_13028,N_12147,N_12206);
or U13029 (N_13029,N_12491,N_12811);
xnor U13030 (N_13030,N_12356,N_12852);
nand U13031 (N_13031,N_12393,N_12512);
nand U13032 (N_13032,N_12888,N_12561);
nor U13033 (N_13033,N_12238,N_12856);
and U13034 (N_13034,N_12142,N_12676);
nand U13035 (N_13035,N_12686,N_12285);
and U13036 (N_13036,N_12691,N_12301);
and U13037 (N_13037,N_12926,N_12935);
nand U13038 (N_13038,N_12536,N_12662);
xor U13039 (N_13039,N_12094,N_12555);
nor U13040 (N_13040,N_12703,N_12369);
or U13041 (N_13041,N_12287,N_12796);
xor U13042 (N_13042,N_12062,N_12256);
and U13043 (N_13043,N_12760,N_12557);
nor U13044 (N_13044,N_12235,N_12661);
nor U13045 (N_13045,N_12523,N_12887);
or U13046 (N_13046,N_12669,N_12089);
and U13047 (N_13047,N_12962,N_12799);
nand U13048 (N_13048,N_12222,N_12036);
xnor U13049 (N_13049,N_12297,N_12422);
nor U13050 (N_13050,N_12969,N_12590);
xnor U13051 (N_13051,N_12058,N_12880);
xnor U13052 (N_13052,N_12299,N_12403);
xnor U13053 (N_13053,N_12990,N_12783);
xor U13054 (N_13054,N_12934,N_12718);
nor U13055 (N_13055,N_12390,N_12451);
nand U13056 (N_13056,N_12644,N_12368);
xnor U13057 (N_13057,N_12334,N_12471);
nor U13058 (N_13058,N_12524,N_12597);
xnor U13059 (N_13059,N_12343,N_12738);
nand U13060 (N_13060,N_12093,N_12564);
and U13061 (N_13061,N_12643,N_12361);
nor U13062 (N_13062,N_12731,N_12956);
and U13063 (N_13063,N_12855,N_12988);
nand U13064 (N_13064,N_12346,N_12653);
nand U13065 (N_13065,N_12033,N_12247);
and U13066 (N_13066,N_12170,N_12814);
nor U13067 (N_13067,N_12525,N_12109);
nor U13068 (N_13068,N_12423,N_12960);
nand U13069 (N_13069,N_12586,N_12825);
and U13070 (N_13070,N_12396,N_12885);
or U13071 (N_13071,N_12298,N_12756);
and U13072 (N_13072,N_12948,N_12627);
nor U13073 (N_13073,N_12223,N_12503);
xor U13074 (N_13074,N_12857,N_12474);
xnor U13075 (N_13075,N_12112,N_12114);
and U13076 (N_13076,N_12635,N_12476);
xor U13077 (N_13077,N_12791,N_12030);
nand U13078 (N_13078,N_12310,N_12117);
nand U13079 (N_13079,N_12761,N_12201);
or U13080 (N_13080,N_12164,N_12993);
nand U13081 (N_13081,N_12336,N_12242);
and U13082 (N_13082,N_12602,N_12100);
and U13083 (N_13083,N_12895,N_12973);
nand U13084 (N_13084,N_12626,N_12961);
or U13085 (N_13085,N_12402,N_12596);
nand U13086 (N_13086,N_12140,N_12508);
or U13087 (N_13087,N_12878,N_12459);
nor U13088 (N_13088,N_12004,N_12842);
or U13089 (N_13089,N_12646,N_12680);
nor U13090 (N_13090,N_12057,N_12700);
or U13091 (N_13091,N_12210,N_12306);
nor U13092 (N_13092,N_12690,N_12376);
nor U13093 (N_13093,N_12283,N_12429);
and U13094 (N_13094,N_12069,N_12560);
nor U13095 (N_13095,N_12194,N_12950);
or U13096 (N_13096,N_12843,N_12636);
or U13097 (N_13097,N_12634,N_12565);
and U13098 (N_13098,N_12707,N_12331);
xor U13099 (N_13099,N_12870,N_12540);
xor U13100 (N_13100,N_12056,N_12481);
nor U13101 (N_13101,N_12103,N_12949);
or U13102 (N_13102,N_12915,N_12231);
and U13103 (N_13103,N_12244,N_12207);
nor U13104 (N_13104,N_12320,N_12573);
nor U13105 (N_13105,N_12556,N_12454);
or U13106 (N_13106,N_12348,N_12131);
nor U13107 (N_13107,N_12335,N_12903);
nand U13108 (N_13108,N_12136,N_12877);
xnor U13109 (N_13109,N_12884,N_12945);
and U13110 (N_13110,N_12191,N_12464);
nand U13111 (N_13111,N_12721,N_12006);
nand U13112 (N_13112,N_12651,N_12132);
and U13113 (N_13113,N_12516,N_12835);
nor U13114 (N_13114,N_12327,N_12763);
xor U13115 (N_13115,N_12266,N_12415);
nor U13116 (N_13116,N_12660,N_12215);
nand U13117 (N_13117,N_12041,N_12453);
nand U13118 (N_13118,N_12279,N_12702);
nor U13119 (N_13119,N_12541,N_12165);
nand U13120 (N_13120,N_12351,N_12527);
nor U13121 (N_13121,N_12668,N_12224);
and U13122 (N_13122,N_12126,N_12407);
nand U13123 (N_13123,N_12359,N_12437);
nor U13124 (N_13124,N_12149,N_12324);
nor U13125 (N_13125,N_12576,N_12406);
nand U13126 (N_13126,N_12939,N_12086);
or U13127 (N_13127,N_12625,N_12765);
or U13128 (N_13128,N_12019,N_12241);
and U13129 (N_13129,N_12052,N_12001);
and U13130 (N_13130,N_12637,N_12360);
and U13131 (N_13131,N_12965,N_12387);
nor U13132 (N_13132,N_12380,N_12188);
nor U13133 (N_13133,N_12462,N_12704);
and U13134 (N_13134,N_12987,N_12239);
or U13135 (N_13135,N_12353,N_12196);
xor U13136 (N_13136,N_12205,N_12233);
xnor U13137 (N_13137,N_12190,N_12155);
nor U13138 (N_13138,N_12031,N_12492);
xnor U13139 (N_13139,N_12658,N_12410);
or U13140 (N_13140,N_12168,N_12873);
nand U13141 (N_13141,N_12829,N_12593);
xor U13142 (N_13142,N_12468,N_12539);
and U13143 (N_13143,N_12101,N_12605);
or U13144 (N_13144,N_12942,N_12896);
nand U13145 (N_13145,N_12946,N_12938);
nor U13146 (N_13146,N_12604,N_12513);
xor U13147 (N_13147,N_12897,N_12902);
and U13148 (N_13148,N_12489,N_12179);
xnor U13149 (N_13149,N_12259,N_12010);
and U13150 (N_13150,N_12439,N_12862);
nand U13151 (N_13151,N_12517,N_12807);
or U13152 (N_13152,N_12281,N_12055);
xor U13153 (N_13153,N_12479,N_12349);
or U13154 (N_13154,N_12409,N_12345);
and U13155 (N_13155,N_12156,N_12773);
or U13156 (N_13156,N_12612,N_12167);
or U13157 (N_13157,N_12780,N_12104);
or U13158 (N_13158,N_12032,N_12044);
xor U13159 (N_13159,N_12379,N_12929);
or U13160 (N_13160,N_12124,N_12532);
xor U13161 (N_13161,N_12998,N_12146);
or U13162 (N_13162,N_12659,N_12405);
nand U13163 (N_13163,N_12908,N_12186);
or U13164 (N_13164,N_12788,N_12600);
nor U13165 (N_13165,N_12826,N_12743);
or U13166 (N_13166,N_12518,N_12200);
nor U13167 (N_13167,N_12683,N_12907);
or U13168 (N_13168,N_12863,N_12434);
xnor U13169 (N_13169,N_12572,N_12568);
nand U13170 (N_13170,N_12175,N_12083);
or U13171 (N_13171,N_12633,N_12108);
nor U13172 (N_13172,N_12262,N_12701);
nor U13173 (N_13173,N_12717,N_12821);
or U13174 (N_13174,N_12663,N_12786);
nand U13175 (N_13175,N_12129,N_12975);
xor U13176 (N_13176,N_12801,N_12138);
nand U13177 (N_13177,N_12574,N_12070);
nor U13178 (N_13178,N_12447,N_12502);
and U13179 (N_13179,N_12347,N_12292);
and U13180 (N_13180,N_12805,N_12931);
nor U13181 (N_13181,N_12158,N_12071);
xnor U13182 (N_13182,N_12894,N_12048);
nor U13183 (N_13183,N_12162,N_12288);
or U13184 (N_13184,N_12460,N_12543);
nor U13185 (N_13185,N_12559,N_12367);
or U13186 (N_13186,N_12810,N_12787);
or U13187 (N_13187,N_12529,N_12936);
xor U13188 (N_13188,N_12566,N_12853);
and U13189 (N_13189,N_12257,N_12332);
and U13190 (N_13190,N_12672,N_12463);
or U13191 (N_13191,N_12461,N_12326);
nand U13192 (N_13192,N_12906,N_12377);
and U13193 (N_13193,N_12024,N_12594);
and U13194 (N_13194,N_12585,N_12027);
nor U13195 (N_13195,N_12449,N_12228);
or U13196 (N_13196,N_12900,N_12013);
nand U13197 (N_13197,N_12876,N_12715);
nand U13198 (N_13198,N_12771,N_12312);
and U13199 (N_13199,N_12264,N_12679);
and U13200 (N_13200,N_12025,N_12999);
or U13201 (N_13201,N_12355,N_12792);
and U13202 (N_13202,N_12802,N_12638);
or U13203 (N_13203,N_12198,N_12340);
nor U13204 (N_13204,N_12029,N_12838);
or U13205 (N_13205,N_12723,N_12022);
nor U13206 (N_13206,N_12064,N_12414);
nor U13207 (N_13207,N_12384,N_12121);
xor U13208 (N_13208,N_12383,N_12665);
xor U13209 (N_13209,N_12265,N_12397);
nor U13210 (N_13210,N_12169,N_12157);
xor U13211 (N_13211,N_12542,N_12373);
or U13212 (N_13212,N_12953,N_12833);
or U13213 (N_13213,N_12074,N_12766);
nor U13214 (N_13214,N_12095,N_12506);
and U13215 (N_13215,N_12674,N_12308);
or U13216 (N_13216,N_12457,N_12304);
nand U13217 (N_13217,N_12722,N_12710);
or U13218 (N_13218,N_12749,N_12184);
or U13219 (N_13219,N_12899,N_12769);
nor U13220 (N_13220,N_12219,N_12319);
nor U13221 (N_13221,N_12160,N_12746);
nand U13222 (N_13222,N_12274,N_12667);
and U13223 (N_13223,N_12485,N_12350);
or U13224 (N_13224,N_12753,N_12757);
nand U13225 (N_13225,N_12671,N_12930);
nand U13226 (N_13226,N_12418,N_12699);
or U13227 (N_13227,N_12519,N_12772);
nor U13228 (N_13228,N_12066,N_12128);
or U13229 (N_13229,N_12830,N_12762);
nor U13230 (N_13230,N_12912,N_12531);
nand U13231 (N_13231,N_12394,N_12425);
xnor U13232 (N_13232,N_12214,N_12150);
and U13233 (N_13233,N_12216,N_12681);
or U13234 (N_13234,N_12005,N_12692);
or U13235 (N_13235,N_12867,N_12195);
nand U13236 (N_13236,N_12624,N_12575);
nor U13237 (N_13237,N_12161,N_12225);
or U13238 (N_13238,N_12261,N_12433);
xnor U13239 (N_13239,N_12918,N_12980);
nor U13240 (N_13240,N_12774,N_12866);
and U13241 (N_13241,N_12972,N_12598);
nand U13242 (N_13242,N_12284,N_12143);
xnor U13243 (N_13243,N_12212,N_12477);
nand U13244 (N_13244,N_12028,N_12061);
or U13245 (N_13245,N_12985,N_12511);
xor U13246 (N_13246,N_12091,N_12096);
nand U13247 (N_13247,N_12197,N_12515);
or U13248 (N_13248,N_12226,N_12291);
nand U13249 (N_13249,N_12554,N_12372);
and U13250 (N_13250,N_12923,N_12417);
or U13251 (N_13251,N_12977,N_12535);
nand U13252 (N_13252,N_12750,N_12253);
or U13253 (N_13253,N_12116,N_12127);
or U13254 (N_13254,N_12174,N_12323);
nor U13255 (N_13255,N_12530,N_12778);
and U13256 (N_13256,N_12145,N_12794);
xor U13257 (N_13257,N_12090,N_12173);
xnor U13258 (N_13258,N_12917,N_12726);
xor U13259 (N_13259,N_12854,N_12398);
nor U13260 (N_13260,N_12898,N_12828);
and U13261 (N_13261,N_12371,N_12545);
nor U13262 (N_13262,N_12490,N_12849);
and U13263 (N_13263,N_12381,N_12657);
nor U13264 (N_13264,N_12591,N_12522);
nand U13265 (N_13265,N_12642,N_12111);
xnor U13266 (N_13266,N_12483,N_12421);
and U13267 (N_13267,N_12411,N_12322);
nor U13268 (N_13268,N_12712,N_12088);
and U13269 (N_13269,N_12603,N_12049);
and U13270 (N_13270,N_12208,N_12469);
xor U13271 (N_13271,N_12337,N_12130);
or U13272 (N_13272,N_12997,N_12435);
xnor U13273 (N_13273,N_12621,N_12694);
and U13274 (N_13274,N_12648,N_12845);
nand U13275 (N_13275,N_12800,N_12916);
nor U13276 (N_13276,N_12249,N_12171);
nor U13277 (N_13277,N_12709,N_12213);
nor U13278 (N_13278,N_12438,N_12578);
nand U13279 (N_13279,N_12592,N_12352);
or U13280 (N_13280,N_12290,N_12725);
xnor U13281 (N_13281,N_12488,N_12448);
nor U13282 (N_13282,N_12549,N_12300);
xnor U13283 (N_13283,N_12611,N_12385);
nand U13284 (N_13284,N_12209,N_12248);
nand U13285 (N_13285,N_12775,N_12436);
nor U13286 (N_13286,N_12747,N_12092);
nand U13287 (N_13287,N_12952,N_12135);
or U13288 (N_13288,N_12046,N_12105);
xor U13289 (N_13289,N_12258,N_12045);
or U13290 (N_13290,N_12487,N_12793);
and U13291 (N_13291,N_12097,N_12795);
xor U13292 (N_13292,N_12307,N_12232);
and U13293 (N_13293,N_12220,N_12589);
or U13294 (N_13294,N_12631,N_12706);
and U13295 (N_13295,N_12909,N_12958);
nand U13296 (N_13296,N_12619,N_12047);
nor U13297 (N_13297,N_12311,N_12951);
or U13298 (N_13298,N_12744,N_12510);
nor U13299 (N_13299,N_12697,N_12813);
xnor U13300 (N_13300,N_12859,N_12832);
nand U13301 (N_13301,N_12705,N_12440);
and U13302 (N_13302,N_12017,N_12363);
and U13303 (N_13303,N_12192,N_12106);
nor U13304 (N_13304,N_12085,N_12728);
and U13305 (N_13305,N_12779,N_12737);
and U13306 (N_13306,N_12251,N_12272);
xor U13307 (N_13307,N_12260,N_12970);
nor U13308 (N_13308,N_12325,N_12243);
nand U13309 (N_13309,N_12647,N_12185);
nand U13310 (N_13310,N_12831,N_12341);
nor U13311 (N_13311,N_12467,N_12655);
nor U13312 (N_13312,N_12014,N_12533);
or U13313 (N_13313,N_12741,N_12782);
or U13314 (N_13314,N_12869,N_12015);
nor U13315 (N_13315,N_12544,N_12270);
nor U13316 (N_13316,N_12925,N_12333);
nor U13317 (N_13317,N_12230,N_12803);
xor U13318 (N_13318,N_12754,N_12202);
nor U13319 (N_13319,N_12494,N_12507);
and U13320 (N_13320,N_12764,N_12401);
and U13321 (N_13321,N_12267,N_12607);
nor U13322 (N_13322,N_12892,N_12458);
xor U13323 (N_13323,N_12893,N_12082);
nand U13324 (N_13324,N_12455,N_12520);
nand U13325 (N_13325,N_12358,N_12685);
nand U13326 (N_13326,N_12837,N_12614);
xor U13327 (N_13327,N_12370,N_12183);
xnor U13328 (N_13328,N_12995,N_12848);
and U13329 (N_13329,N_12812,N_12724);
xor U13330 (N_13330,N_12182,N_12504);
and U13331 (N_13331,N_12313,N_12180);
nor U13332 (N_13332,N_12497,N_12296);
nand U13333 (N_13333,N_12039,N_12971);
or U13334 (N_13334,N_12742,N_12865);
xnor U13335 (N_13335,N_12321,N_12020);
xor U13336 (N_13336,N_12354,N_12427);
or U13337 (N_13337,N_12992,N_12472);
or U13338 (N_13338,N_12547,N_12294);
xor U13339 (N_13339,N_12172,N_12255);
xor U13340 (N_13340,N_12268,N_12315);
xor U13341 (N_13341,N_12979,N_12546);
and U13342 (N_13342,N_12919,N_12739);
nor U13343 (N_13343,N_12587,N_12227);
or U13344 (N_13344,N_12473,N_12968);
nand U13345 (N_13345,N_12932,N_12389);
nand U13346 (N_13346,N_12601,N_12770);
or U13347 (N_13347,N_12714,N_12632);
nand U13348 (N_13348,N_12820,N_12000);
xor U13349 (N_13349,N_12617,N_12615);
nand U13350 (N_13350,N_12577,N_12514);
xnor U13351 (N_13351,N_12727,N_12850);
or U13352 (N_13352,N_12616,N_12879);
and U13353 (N_13353,N_12176,N_12456);
xnor U13354 (N_13354,N_12318,N_12551);
xnor U13355 (N_13355,N_12501,N_12933);
xor U13356 (N_13356,N_12177,N_12081);
or U13357 (N_13357,N_12122,N_12982);
nor U13358 (N_13358,N_12077,N_12720);
nor U13359 (N_13359,N_12317,N_12009);
or U13360 (N_13360,N_12834,N_12840);
nor U13361 (N_13361,N_12018,N_12964);
or U13362 (N_13362,N_12711,N_12280);
or U13363 (N_13363,N_12940,N_12078);
or U13364 (N_13364,N_12102,N_12944);
nor U13365 (N_13365,N_12388,N_12804);
nand U13366 (N_13366,N_12021,N_12736);
and U13367 (N_13367,N_12986,N_12151);
or U13368 (N_13368,N_12966,N_12963);
xnor U13369 (N_13369,N_12400,N_12839);
xor U13370 (N_13370,N_12861,N_12858);
or U13371 (N_13371,N_12630,N_12273);
xor U13372 (N_13372,N_12562,N_12868);
xnor U13373 (N_13373,N_12579,N_12675);
xnor U13374 (N_13374,N_12716,N_12302);
and U13375 (N_13375,N_12654,N_12528);
and U13376 (N_13376,N_12446,N_12606);
nand U13377 (N_13377,N_12073,N_12098);
nor U13378 (N_13378,N_12818,N_12534);
and U13379 (N_13379,N_12827,N_12689);
nor U13380 (N_13380,N_12303,N_12943);
or U13381 (N_13381,N_12583,N_12470);
and U13382 (N_13382,N_12687,N_12901);
or U13383 (N_13383,N_12844,N_12847);
nor U13384 (N_13384,N_12254,N_12588);
and U13385 (N_13385,N_12684,N_12475);
nor U13386 (N_13386,N_12002,N_12875);
nand U13387 (N_13387,N_12914,N_12570);
nand U13388 (N_13388,N_12666,N_12595);
nand U13389 (N_13389,N_12234,N_12042);
or U13390 (N_13390,N_12465,N_12392);
nand U13391 (N_13391,N_12067,N_12493);
xnor U13392 (N_13392,N_12053,N_12060);
xnor U13393 (N_13393,N_12424,N_12011);
nand U13394 (N_13394,N_12735,N_12629);
or U13395 (N_13395,N_12211,N_12395);
and U13396 (N_13396,N_12329,N_12790);
nand U13397 (N_13397,N_12552,N_12163);
and U13398 (N_13398,N_12187,N_12733);
and U13399 (N_13399,N_12822,N_12293);
nand U13400 (N_13400,N_12537,N_12732);
nand U13401 (N_13401,N_12841,N_12416);
nor U13402 (N_13402,N_12050,N_12330);
nor U13403 (N_13403,N_12250,N_12107);
and U13404 (N_13404,N_12713,N_12295);
or U13405 (N_13405,N_12955,N_12751);
and U13406 (N_13406,N_12623,N_12526);
nor U13407 (N_13407,N_12075,N_12026);
nor U13408 (N_13408,N_12189,N_12412);
nor U13409 (N_13409,N_12375,N_12874);
or U13410 (N_13410,N_12784,N_12759);
nor U13411 (N_13411,N_12084,N_12580);
xor U13412 (N_13412,N_12316,N_12034);
nor U13413 (N_13413,N_12362,N_12881);
xor U13414 (N_13414,N_12639,N_12003);
xor U13415 (N_13415,N_12450,N_12240);
nor U13416 (N_13416,N_12563,N_12740);
nand U13417 (N_13417,N_12521,N_12824);
nand U13418 (N_13418,N_12305,N_12567);
nand U13419 (N_13419,N_12134,N_12099);
or U13420 (N_13420,N_12133,N_12063);
nand U13421 (N_13421,N_12144,N_12991);
and U13422 (N_13422,N_12426,N_12314);
or U13423 (N_13423,N_12652,N_12263);
or U13424 (N_13424,N_12408,N_12278);
and U13425 (N_13425,N_12068,N_12148);
xnor U13426 (N_13426,N_12342,N_12910);
nor U13427 (N_13427,N_12921,N_12038);
and U13428 (N_13428,N_12571,N_12040);
or U13429 (N_13429,N_12748,N_12846);
xnor U13430 (N_13430,N_12123,N_12823);
xor U13431 (N_13431,N_12277,N_12432);
nand U13432 (N_13432,N_12178,N_12509);
nor U13433 (N_13433,N_12886,N_12166);
xnor U13434 (N_13434,N_12628,N_12382);
xnor U13435 (N_13435,N_12391,N_12609);
nor U13436 (N_13436,N_12941,N_12229);
or U13437 (N_13437,N_12688,N_12767);
nand U13438 (N_13438,N_12808,N_12023);
or U13439 (N_13439,N_12798,N_12610);
and U13440 (N_13440,N_12237,N_12374);
or U13441 (N_13441,N_12569,N_12889);
nand U13442 (N_13442,N_12153,N_12484);
nor U13443 (N_13443,N_12478,N_12486);
xor U13444 (N_13444,N_12677,N_12905);
xor U13445 (N_13445,N_12443,N_12983);
and U13446 (N_13446,N_12217,N_12872);
and U13447 (N_13447,N_12399,N_12550);
or U13448 (N_13448,N_12978,N_12640);
nor U13449 (N_13449,N_12994,N_12012);
and U13450 (N_13450,N_12553,N_12065);
and U13451 (N_13451,N_12620,N_12678);
nand U13452 (N_13452,N_12339,N_12815);
nand U13453 (N_13453,N_12007,N_12496);
xor U13454 (N_13454,N_12181,N_12378);
nand U13455 (N_13455,N_12797,N_12043);
nand U13456 (N_13456,N_12682,N_12920);
and U13457 (N_13457,N_12981,N_12137);
nand U13458 (N_13458,N_12271,N_12584);
or U13459 (N_13459,N_12499,N_12618);
nor U13460 (N_13460,N_12752,N_12199);
nand U13461 (N_13461,N_12275,N_12967);
and U13462 (N_13462,N_12120,N_12115);
xor U13463 (N_13463,N_12882,N_12673);
nand U13464 (N_13464,N_12696,N_12282);
or U13465 (N_13465,N_12816,N_12883);
nand U13466 (N_13466,N_12819,N_12154);
and U13467 (N_13467,N_12613,N_12419);
xor U13468 (N_13468,N_12413,N_12954);
nor U13469 (N_13469,N_12404,N_12864);
nand U13470 (N_13470,N_12871,N_12495);
and U13471 (N_13471,N_12059,N_12236);
nand U13472 (N_13472,N_12309,N_12758);
xor U13473 (N_13473,N_12851,N_12548);
nor U13474 (N_13474,N_12269,N_12789);
nand U13475 (N_13475,N_12664,N_12649);
xor U13476 (N_13476,N_12246,N_12080);
nand U13477 (N_13477,N_12087,N_12734);
xnor U13478 (N_13478,N_12924,N_12538);
or U13479 (N_13479,N_12203,N_12913);
or U13480 (N_13480,N_12695,N_12482);
nor U13481 (N_13481,N_12386,N_12776);
xnor U13482 (N_13482,N_12221,N_12139);
nor U13483 (N_13483,N_12730,N_12785);
nor U13484 (N_13484,N_12428,N_12072);
and U13485 (N_13485,N_12890,N_12911);
nor U13486 (N_13486,N_12947,N_12755);
nand U13487 (N_13487,N_12430,N_12599);
nor U13488 (N_13488,N_12118,N_12608);
xnor U13489 (N_13489,N_12650,N_12035);
nor U13490 (N_13490,N_12218,N_12276);
and U13491 (N_13491,N_12445,N_12558);
nor U13492 (N_13492,N_12365,N_12357);
nand U13493 (N_13493,N_12777,N_12328);
nand U13494 (N_13494,N_12768,N_12656);
and U13495 (N_13495,N_12500,N_12051);
and U13496 (N_13496,N_12641,N_12204);
nor U13497 (N_13497,N_12054,N_12745);
nand U13498 (N_13498,N_12119,N_12008);
nor U13499 (N_13499,N_12431,N_12444);
or U13500 (N_13500,N_12072,N_12283);
and U13501 (N_13501,N_12826,N_12716);
or U13502 (N_13502,N_12708,N_12522);
nor U13503 (N_13503,N_12378,N_12472);
nor U13504 (N_13504,N_12190,N_12074);
xnor U13505 (N_13505,N_12324,N_12056);
and U13506 (N_13506,N_12576,N_12896);
nand U13507 (N_13507,N_12066,N_12305);
and U13508 (N_13508,N_12783,N_12907);
nand U13509 (N_13509,N_12053,N_12911);
and U13510 (N_13510,N_12480,N_12166);
xnor U13511 (N_13511,N_12456,N_12295);
nor U13512 (N_13512,N_12070,N_12883);
and U13513 (N_13513,N_12495,N_12863);
nor U13514 (N_13514,N_12493,N_12050);
nand U13515 (N_13515,N_12861,N_12327);
nor U13516 (N_13516,N_12950,N_12348);
nand U13517 (N_13517,N_12574,N_12346);
or U13518 (N_13518,N_12515,N_12570);
nand U13519 (N_13519,N_12280,N_12687);
nand U13520 (N_13520,N_12422,N_12402);
or U13521 (N_13521,N_12388,N_12356);
and U13522 (N_13522,N_12341,N_12793);
xor U13523 (N_13523,N_12925,N_12904);
nor U13524 (N_13524,N_12038,N_12623);
nor U13525 (N_13525,N_12576,N_12710);
and U13526 (N_13526,N_12669,N_12580);
xnor U13527 (N_13527,N_12188,N_12789);
nor U13528 (N_13528,N_12953,N_12375);
xor U13529 (N_13529,N_12506,N_12454);
nor U13530 (N_13530,N_12860,N_12746);
xor U13531 (N_13531,N_12289,N_12593);
nand U13532 (N_13532,N_12052,N_12002);
xor U13533 (N_13533,N_12932,N_12709);
and U13534 (N_13534,N_12348,N_12024);
xor U13535 (N_13535,N_12636,N_12133);
or U13536 (N_13536,N_12652,N_12778);
nand U13537 (N_13537,N_12136,N_12979);
xor U13538 (N_13538,N_12520,N_12884);
xor U13539 (N_13539,N_12423,N_12091);
and U13540 (N_13540,N_12023,N_12446);
and U13541 (N_13541,N_12355,N_12441);
or U13542 (N_13542,N_12207,N_12092);
nand U13543 (N_13543,N_12529,N_12389);
or U13544 (N_13544,N_12166,N_12497);
nor U13545 (N_13545,N_12023,N_12332);
or U13546 (N_13546,N_12813,N_12826);
xnor U13547 (N_13547,N_12796,N_12012);
nand U13548 (N_13548,N_12980,N_12582);
nor U13549 (N_13549,N_12814,N_12885);
and U13550 (N_13550,N_12472,N_12078);
xnor U13551 (N_13551,N_12435,N_12585);
nor U13552 (N_13552,N_12980,N_12894);
xor U13553 (N_13553,N_12515,N_12502);
nand U13554 (N_13554,N_12775,N_12562);
or U13555 (N_13555,N_12792,N_12238);
xor U13556 (N_13556,N_12006,N_12493);
and U13557 (N_13557,N_12396,N_12110);
nor U13558 (N_13558,N_12987,N_12829);
or U13559 (N_13559,N_12426,N_12463);
xnor U13560 (N_13560,N_12011,N_12484);
or U13561 (N_13561,N_12404,N_12111);
and U13562 (N_13562,N_12886,N_12413);
xor U13563 (N_13563,N_12564,N_12578);
xor U13564 (N_13564,N_12590,N_12305);
nand U13565 (N_13565,N_12499,N_12749);
nand U13566 (N_13566,N_12547,N_12143);
or U13567 (N_13567,N_12880,N_12227);
nand U13568 (N_13568,N_12597,N_12916);
xnor U13569 (N_13569,N_12833,N_12135);
nor U13570 (N_13570,N_12879,N_12925);
xor U13571 (N_13571,N_12487,N_12596);
xor U13572 (N_13572,N_12513,N_12534);
or U13573 (N_13573,N_12287,N_12235);
nor U13574 (N_13574,N_12705,N_12936);
xnor U13575 (N_13575,N_12608,N_12864);
or U13576 (N_13576,N_12785,N_12240);
nand U13577 (N_13577,N_12419,N_12650);
or U13578 (N_13578,N_12522,N_12186);
nor U13579 (N_13579,N_12075,N_12260);
nor U13580 (N_13580,N_12748,N_12521);
or U13581 (N_13581,N_12054,N_12644);
xor U13582 (N_13582,N_12649,N_12327);
nor U13583 (N_13583,N_12993,N_12239);
and U13584 (N_13584,N_12972,N_12759);
nand U13585 (N_13585,N_12210,N_12428);
or U13586 (N_13586,N_12185,N_12722);
nor U13587 (N_13587,N_12509,N_12819);
nor U13588 (N_13588,N_12052,N_12324);
nand U13589 (N_13589,N_12182,N_12678);
nand U13590 (N_13590,N_12658,N_12834);
and U13591 (N_13591,N_12990,N_12317);
or U13592 (N_13592,N_12840,N_12592);
or U13593 (N_13593,N_12598,N_12389);
or U13594 (N_13594,N_12096,N_12937);
nor U13595 (N_13595,N_12240,N_12653);
xnor U13596 (N_13596,N_12690,N_12393);
or U13597 (N_13597,N_12395,N_12766);
or U13598 (N_13598,N_12859,N_12160);
or U13599 (N_13599,N_12610,N_12614);
nand U13600 (N_13600,N_12615,N_12266);
xnor U13601 (N_13601,N_12349,N_12500);
nand U13602 (N_13602,N_12016,N_12806);
and U13603 (N_13603,N_12636,N_12182);
nand U13604 (N_13604,N_12755,N_12176);
or U13605 (N_13605,N_12535,N_12055);
xor U13606 (N_13606,N_12291,N_12249);
and U13607 (N_13607,N_12614,N_12602);
and U13608 (N_13608,N_12291,N_12755);
nand U13609 (N_13609,N_12315,N_12291);
nor U13610 (N_13610,N_12310,N_12875);
nor U13611 (N_13611,N_12722,N_12083);
nor U13612 (N_13612,N_12941,N_12082);
xnor U13613 (N_13613,N_12578,N_12508);
xnor U13614 (N_13614,N_12010,N_12413);
and U13615 (N_13615,N_12216,N_12632);
nor U13616 (N_13616,N_12213,N_12918);
nand U13617 (N_13617,N_12643,N_12930);
or U13618 (N_13618,N_12344,N_12485);
or U13619 (N_13619,N_12108,N_12586);
nor U13620 (N_13620,N_12104,N_12038);
xor U13621 (N_13621,N_12469,N_12095);
and U13622 (N_13622,N_12824,N_12958);
or U13623 (N_13623,N_12116,N_12531);
nand U13624 (N_13624,N_12497,N_12304);
nand U13625 (N_13625,N_12705,N_12550);
xnor U13626 (N_13626,N_12287,N_12099);
or U13627 (N_13627,N_12355,N_12864);
nand U13628 (N_13628,N_12509,N_12719);
xnor U13629 (N_13629,N_12018,N_12293);
and U13630 (N_13630,N_12467,N_12614);
and U13631 (N_13631,N_12512,N_12000);
xnor U13632 (N_13632,N_12382,N_12177);
nand U13633 (N_13633,N_12971,N_12759);
xnor U13634 (N_13634,N_12916,N_12363);
and U13635 (N_13635,N_12953,N_12220);
nor U13636 (N_13636,N_12068,N_12825);
xnor U13637 (N_13637,N_12114,N_12471);
and U13638 (N_13638,N_12177,N_12272);
nand U13639 (N_13639,N_12738,N_12877);
xnor U13640 (N_13640,N_12755,N_12592);
or U13641 (N_13641,N_12759,N_12801);
xnor U13642 (N_13642,N_12710,N_12657);
or U13643 (N_13643,N_12877,N_12461);
xor U13644 (N_13644,N_12694,N_12448);
nand U13645 (N_13645,N_12581,N_12705);
nor U13646 (N_13646,N_12635,N_12646);
nor U13647 (N_13647,N_12169,N_12070);
xnor U13648 (N_13648,N_12144,N_12528);
xnor U13649 (N_13649,N_12689,N_12504);
xor U13650 (N_13650,N_12877,N_12043);
xor U13651 (N_13651,N_12118,N_12053);
nor U13652 (N_13652,N_12706,N_12930);
nand U13653 (N_13653,N_12815,N_12688);
nand U13654 (N_13654,N_12732,N_12766);
nand U13655 (N_13655,N_12790,N_12617);
xnor U13656 (N_13656,N_12604,N_12090);
or U13657 (N_13657,N_12551,N_12471);
and U13658 (N_13658,N_12572,N_12866);
xor U13659 (N_13659,N_12883,N_12417);
xnor U13660 (N_13660,N_12247,N_12085);
nand U13661 (N_13661,N_12970,N_12759);
or U13662 (N_13662,N_12734,N_12809);
xnor U13663 (N_13663,N_12589,N_12207);
nand U13664 (N_13664,N_12841,N_12353);
and U13665 (N_13665,N_12204,N_12821);
nor U13666 (N_13666,N_12767,N_12217);
nand U13667 (N_13667,N_12430,N_12957);
and U13668 (N_13668,N_12411,N_12859);
nand U13669 (N_13669,N_12703,N_12511);
and U13670 (N_13670,N_12299,N_12644);
nand U13671 (N_13671,N_12479,N_12480);
or U13672 (N_13672,N_12838,N_12073);
or U13673 (N_13673,N_12583,N_12721);
nand U13674 (N_13674,N_12406,N_12204);
or U13675 (N_13675,N_12602,N_12907);
or U13676 (N_13676,N_12826,N_12585);
xnor U13677 (N_13677,N_12626,N_12121);
xnor U13678 (N_13678,N_12679,N_12021);
and U13679 (N_13679,N_12651,N_12638);
nor U13680 (N_13680,N_12134,N_12833);
nand U13681 (N_13681,N_12764,N_12335);
xnor U13682 (N_13682,N_12808,N_12182);
or U13683 (N_13683,N_12997,N_12741);
and U13684 (N_13684,N_12200,N_12346);
nor U13685 (N_13685,N_12068,N_12141);
xor U13686 (N_13686,N_12864,N_12577);
nand U13687 (N_13687,N_12940,N_12013);
xnor U13688 (N_13688,N_12531,N_12827);
nand U13689 (N_13689,N_12967,N_12802);
or U13690 (N_13690,N_12094,N_12158);
and U13691 (N_13691,N_12365,N_12754);
and U13692 (N_13692,N_12576,N_12910);
xnor U13693 (N_13693,N_12501,N_12205);
nor U13694 (N_13694,N_12955,N_12972);
or U13695 (N_13695,N_12572,N_12015);
nand U13696 (N_13696,N_12993,N_12506);
and U13697 (N_13697,N_12435,N_12215);
nor U13698 (N_13698,N_12985,N_12393);
and U13699 (N_13699,N_12488,N_12228);
nor U13700 (N_13700,N_12274,N_12775);
nand U13701 (N_13701,N_12476,N_12897);
or U13702 (N_13702,N_12298,N_12763);
or U13703 (N_13703,N_12838,N_12645);
or U13704 (N_13704,N_12039,N_12579);
nor U13705 (N_13705,N_12512,N_12231);
nor U13706 (N_13706,N_12559,N_12615);
nand U13707 (N_13707,N_12346,N_12839);
nor U13708 (N_13708,N_12393,N_12923);
nor U13709 (N_13709,N_12977,N_12069);
or U13710 (N_13710,N_12339,N_12414);
nor U13711 (N_13711,N_12918,N_12444);
nand U13712 (N_13712,N_12372,N_12906);
nor U13713 (N_13713,N_12336,N_12508);
nor U13714 (N_13714,N_12321,N_12941);
or U13715 (N_13715,N_12931,N_12083);
or U13716 (N_13716,N_12585,N_12420);
and U13717 (N_13717,N_12990,N_12598);
xnor U13718 (N_13718,N_12554,N_12168);
nor U13719 (N_13719,N_12868,N_12885);
nor U13720 (N_13720,N_12996,N_12668);
nor U13721 (N_13721,N_12098,N_12807);
xnor U13722 (N_13722,N_12575,N_12660);
and U13723 (N_13723,N_12886,N_12253);
nand U13724 (N_13724,N_12373,N_12075);
nand U13725 (N_13725,N_12171,N_12101);
or U13726 (N_13726,N_12489,N_12682);
nor U13727 (N_13727,N_12284,N_12668);
or U13728 (N_13728,N_12239,N_12278);
nor U13729 (N_13729,N_12219,N_12179);
nand U13730 (N_13730,N_12401,N_12282);
nand U13731 (N_13731,N_12369,N_12497);
xnor U13732 (N_13732,N_12371,N_12246);
and U13733 (N_13733,N_12310,N_12657);
or U13734 (N_13734,N_12340,N_12353);
xnor U13735 (N_13735,N_12489,N_12290);
or U13736 (N_13736,N_12073,N_12170);
and U13737 (N_13737,N_12712,N_12670);
and U13738 (N_13738,N_12764,N_12552);
and U13739 (N_13739,N_12554,N_12714);
xor U13740 (N_13740,N_12495,N_12385);
xnor U13741 (N_13741,N_12696,N_12649);
and U13742 (N_13742,N_12305,N_12527);
nand U13743 (N_13743,N_12606,N_12316);
and U13744 (N_13744,N_12056,N_12390);
xor U13745 (N_13745,N_12524,N_12505);
and U13746 (N_13746,N_12989,N_12811);
nor U13747 (N_13747,N_12407,N_12837);
nor U13748 (N_13748,N_12940,N_12694);
nor U13749 (N_13749,N_12577,N_12771);
or U13750 (N_13750,N_12636,N_12725);
or U13751 (N_13751,N_12528,N_12793);
nor U13752 (N_13752,N_12035,N_12763);
nor U13753 (N_13753,N_12791,N_12651);
or U13754 (N_13754,N_12274,N_12654);
nand U13755 (N_13755,N_12677,N_12417);
nand U13756 (N_13756,N_12498,N_12288);
xor U13757 (N_13757,N_12642,N_12689);
nand U13758 (N_13758,N_12389,N_12181);
and U13759 (N_13759,N_12683,N_12886);
and U13760 (N_13760,N_12923,N_12209);
and U13761 (N_13761,N_12082,N_12764);
nand U13762 (N_13762,N_12148,N_12130);
nor U13763 (N_13763,N_12962,N_12260);
and U13764 (N_13764,N_12422,N_12272);
nor U13765 (N_13765,N_12932,N_12707);
nor U13766 (N_13766,N_12735,N_12145);
nor U13767 (N_13767,N_12054,N_12607);
nor U13768 (N_13768,N_12853,N_12581);
nor U13769 (N_13769,N_12510,N_12402);
and U13770 (N_13770,N_12100,N_12135);
nand U13771 (N_13771,N_12657,N_12935);
nor U13772 (N_13772,N_12154,N_12459);
or U13773 (N_13773,N_12254,N_12553);
and U13774 (N_13774,N_12825,N_12186);
nor U13775 (N_13775,N_12892,N_12333);
nand U13776 (N_13776,N_12810,N_12560);
nand U13777 (N_13777,N_12302,N_12306);
nand U13778 (N_13778,N_12005,N_12949);
nand U13779 (N_13779,N_12499,N_12835);
or U13780 (N_13780,N_12948,N_12947);
xor U13781 (N_13781,N_12537,N_12784);
xor U13782 (N_13782,N_12439,N_12283);
xnor U13783 (N_13783,N_12605,N_12110);
nand U13784 (N_13784,N_12858,N_12835);
or U13785 (N_13785,N_12225,N_12327);
nand U13786 (N_13786,N_12338,N_12813);
nand U13787 (N_13787,N_12231,N_12236);
nand U13788 (N_13788,N_12357,N_12429);
nor U13789 (N_13789,N_12361,N_12459);
and U13790 (N_13790,N_12618,N_12213);
nor U13791 (N_13791,N_12663,N_12316);
nor U13792 (N_13792,N_12025,N_12707);
nand U13793 (N_13793,N_12228,N_12411);
nor U13794 (N_13794,N_12719,N_12897);
or U13795 (N_13795,N_12452,N_12838);
and U13796 (N_13796,N_12569,N_12943);
nor U13797 (N_13797,N_12304,N_12259);
and U13798 (N_13798,N_12762,N_12010);
nand U13799 (N_13799,N_12563,N_12730);
and U13800 (N_13800,N_12208,N_12559);
or U13801 (N_13801,N_12091,N_12723);
and U13802 (N_13802,N_12685,N_12108);
and U13803 (N_13803,N_12256,N_12517);
or U13804 (N_13804,N_12107,N_12660);
xnor U13805 (N_13805,N_12020,N_12596);
nand U13806 (N_13806,N_12910,N_12147);
and U13807 (N_13807,N_12560,N_12350);
xnor U13808 (N_13808,N_12650,N_12568);
or U13809 (N_13809,N_12404,N_12134);
or U13810 (N_13810,N_12268,N_12694);
or U13811 (N_13811,N_12465,N_12019);
and U13812 (N_13812,N_12521,N_12330);
nand U13813 (N_13813,N_12780,N_12082);
nor U13814 (N_13814,N_12981,N_12991);
nand U13815 (N_13815,N_12439,N_12462);
nor U13816 (N_13816,N_12526,N_12041);
xor U13817 (N_13817,N_12306,N_12640);
or U13818 (N_13818,N_12829,N_12159);
and U13819 (N_13819,N_12428,N_12708);
nand U13820 (N_13820,N_12103,N_12658);
and U13821 (N_13821,N_12923,N_12467);
nor U13822 (N_13822,N_12941,N_12002);
nor U13823 (N_13823,N_12448,N_12139);
nand U13824 (N_13824,N_12263,N_12480);
nor U13825 (N_13825,N_12882,N_12574);
nand U13826 (N_13826,N_12639,N_12907);
xnor U13827 (N_13827,N_12948,N_12292);
or U13828 (N_13828,N_12055,N_12553);
nand U13829 (N_13829,N_12950,N_12028);
and U13830 (N_13830,N_12046,N_12897);
xor U13831 (N_13831,N_12007,N_12658);
xnor U13832 (N_13832,N_12091,N_12336);
xor U13833 (N_13833,N_12337,N_12825);
xor U13834 (N_13834,N_12524,N_12908);
nand U13835 (N_13835,N_12399,N_12276);
nor U13836 (N_13836,N_12714,N_12253);
nand U13837 (N_13837,N_12559,N_12638);
or U13838 (N_13838,N_12726,N_12542);
nor U13839 (N_13839,N_12785,N_12597);
xor U13840 (N_13840,N_12141,N_12000);
nand U13841 (N_13841,N_12830,N_12188);
and U13842 (N_13842,N_12337,N_12908);
and U13843 (N_13843,N_12095,N_12719);
and U13844 (N_13844,N_12797,N_12943);
and U13845 (N_13845,N_12940,N_12126);
nor U13846 (N_13846,N_12712,N_12110);
or U13847 (N_13847,N_12850,N_12915);
xnor U13848 (N_13848,N_12615,N_12308);
nor U13849 (N_13849,N_12851,N_12425);
or U13850 (N_13850,N_12936,N_12064);
nor U13851 (N_13851,N_12959,N_12361);
nand U13852 (N_13852,N_12519,N_12928);
or U13853 (N_13853,N_12195,N_12873);
nand U13854 (N_13854,N_12096,N_12216);
xor U13855 (N_13855,N_12420,N_12920);
xnor U13856 (N_13856,N_12514,N_12169);
nand U13857 (N_13857,N_12274,N_12102);
nand U13858 (N_13858,N_12806,N_12298);
xnor U13859 (N_13859,N_12223,N_12814);
or U13860 (N_13860,N_12430,N_12397);
nor U13861 (N_13861,N_12875,N_12213);
and U13862 (N_13862,N_12656,N_12494);
xor U13863 (N_13863,N_12857,N_12225);
or U13864 (N_13864,N_12890,N_12434);
nor U13865 (N_13865,N_12050,N_12523);
and U13866 (N_13866,N_12166,N_12108);
xnor U13867 (N_13867,N_12672,N_12364);
xor U13868 (N_13868,N_12832,N_12593);
xor U13869 (N_13869,N_12801,N_12013);
nand U13870 (N_13870,N_12390,N_12585);
or U13871 (N_13871,N_12273,N_12083);
or U13872 (N_13872,N_12782,N_12167);
xnor U13873 (N_13873,N_12636,N_12528);
and U13874 (N_13874,N_12847,N_12092);
and U13875 (N_13875,N_12513,N_12307);
or U13876 (N_13876,N_12245,N_12083);
nor U13877 (N_13877,N_12040,N_12993);
and U13878 (N_13878,N_12915,N_12772);
or U13879 (N_13879,N_12963,N_12479);
or U13880 (N_13880,N_12594,N_12691);
or U13881 (N_13881,N_12983,N_12536);
or U13882 (N_13882,N_12498,N_12786);
nor U13883 (N_13883,N_12536,N_12136);
or U13884 (N_13884,N_12393,N_12223);
nor U13885 (N_13885,N_12232,N_12929);
or U13886 (N_13886,N_12578,N_12309);
nor U13887 (N_13887,N_12802,N_12444);
xnor U13888 (N_13888,N_12958,N_12275);
nand U13889 (N_13889,N_12030,N_12949);
xnor U13890 (N_13890,N_12049,N_12682);
nand U13891 (N_13891,N_12660,N_12391);
nor U13892 (N_13892,N_12918,N_12338);
nand U13893 (N_13893,N_12666,N_12970);
nor U13894 (N_13894,N_12049,N_12470);
xnor U13895 (N_13895,N_12340,N_12343);
and U13896 (N_13896,N_12997,N_12254);
nor U13897 (N_13897,N_12491,N_12994);
xor U13898 (N_13898,N_12313,N_12575);
and U13899 (N_13899,N_12911,N_12719);
or U13900 (N_13900,N_12034,N_12285);
or U13901 (N_13901,N_12119,N_12481);
nand U13902 (N_13902,N_12415,N_12273);
xor U13903 (N_13903,N_12685,N_12676);
xor U13904 (N_13904,N_12108,N_12191);
nor U13905 (N_13905,N_12753,N_12545);
or U13906 (N_13906,N_12359,N_12676);
nand U13907 (N_13907,N_12167,N_12848);
nand U13908 (N_13908,N_12646,N_12963);
nor U13909 (N_13909,N_12009,N_12924);
or U13910 (N_13910,N_12745,N_12473);
and U13911 (N_13911,N_12274,N_12664);
nor U13912 (N_13912,N_12316,N_12895);
nand U13913 (N_13913,N_12754,N_12481);
xor U13914 (N_13914,N_12577,N_12637);
nand U13915 (N_13915,N_12855,N_12522);
nand U13916 (N_13916,N_12737,N_12530);
xor U13917 (N_13917,N_12602,N_12987);
xnor U13918 (N_13918,N_12188,N_12349);
nand U13919 (N_13919,N_12928,N_12140);
nor U13920 (N_13920,N_12319,N_12682);
xnor U13921 (N_13921,N_12398,N_12439);
or U13922 (N_13922,N_12394,N_12990);
nor U13923 (N_13923,N_12800,N_12168);
or U13924 (N_13924,N_12383,N_12582);
nand U13925 (N_13925,N_12012,N_12508);
nand U13926 (N_13926,N_12611,N_12570);
nand U13927 (N_13927,N_12706,N_12453);
xnor U13928 (N_13928,N_12913,N_12583);
nand U13929 (N_13929,N_12690,N_12276);
nor U13930 (N_13930,N_12833,N_12938);
or U13931 (N_13931,N_12478,N_12825);
and U13932 (N_13932,N_12442,N_12796);
and U13933 (N_13933,N_12570,N_12144);
xor U13934 (N_13934,N_12042,N_12248);
xor U13935 (N_13935,N_12749,N_12047);
nor U13936 (N_13936,N_12136,N_12278);
or U13937 (N_13937,N_12351,N_12561);
or U13938 (N_13938,N_12251,N_12402);
and U13939 (N_13939,N_12262,N_12738);
nor U13940 (N_13940,N_12487,N_12115);
and U13941 (N_13941,N_12514,N_12444);
and U13942 (N_13942,N_12034,N_12738);
and U13943 (N_13943,N_12248,N_12235);
and U13944 (N_13944,N_12613,N_12727);
nand U13945 (N_13945,N_12033,N_12582);
nand U13946 (N_13946,N_12361,N_12225);
nor U13947 (N_13947,N_12012,N_12875);
and U13948 (N_13948,N_12948,N_12151);
nor U13949 (N_13949,N_12174,N_12583);
and U13950 (N_13950,N_12403,N_12231);
nor U13951 (N_13951,N_12700,N_12751);
nand U13952 (N_13952,N_12620,N_12417);
and U13953 (N_13953,N_12585,N_12479);
nand U13954 (N_13954,N_12289,N_12874);
and U13955 (N_13955,N_12023,N_12424);
nand U13956 (N_13956,N_12727,N_12381);
nor U13957 (N_13957,N_12250,N_12941);
or U13958 (N_13958,N_12156,N_12377);
nor U13959 (N_13959,N_12038,N_12358);
xor U13960 (N_13960,N_12464,N_12515);
nor U13961 (N_13961,N_12008,N_12866);
nor U13962 (N_13962,N_12523,N_12554);
xnor U13963 (N_13963,N_12701,N_12144);
nand U13964 (N_13964,N_12936,N_12608);
xor U13965 (N_13965,N_12941,N_12722);
and U13966 (N_13966,N_12390,N_12379);
xor U13967 (N_13967,N_12078,N_12377);
xnor U13968 (N_13968,N_12735,N_12680);
nand U13969 (N_13969,N_12530,N_12732);
or U13970 (N_13970,N_12527,N_12252);
and U13971 (N_13971,N_12603,N_12240);
xor U13972 (N_13972,N_12993,N_12009);
nor U13973 (N_13973,N_12209,N_12436);
nand U13974 (N_13974,N_12913,N_12136);
nor U13975 (N_13975,N_12037,N_12660);
or U13976 (N_13976,N_12534,N_12439);
nand U13977 (N_13977,N_12814,N_12317);
nor U13978 (N_13978,N_12518,N_12429);
or U13979 (N_13979,N_12857,N_12396);
or U13980 (N_13980,N_12830,N_12260);
or U13981 (N_13981,N_12678,N_12954);
or U13982 (N_13982,N_12695,N_12663);
or U13983 (N_13983,N_12778,N_12322);
or U13984 (N_13984,N_12087,N_12292);
nor U13985 (N_13985,N_12299,N_12713);
nand U13986 (N_13986,N_12937,N_12987);
and U13987 (N_13987,N_12891,N_12950);
nor U13988 (N_13988,N_12445,N_12850);
nand U13989 (N_13989,N_12228,N_12262);
or U13990 (N_13990,N_12317,N_12205);
nor U13991 (N_13991,N_12175,N_12886);
or U13992 (N_13992,N_12320,N_12793);
xnor U13993 (N_13993,N_12101,N_12272);
nor U13994 (N_13994,N_12323,N_12024);
or U13995 (N_13995,N_12351,N_12590);
xnor U13996 (N_13996,N_12833,N_12782);
and U13997 (N_13997,N_12246,N_12810);
nand U13998 (N_13998,N_12091,N_12655);
xnor U13999 (N_13999,N_12450,N_12774);
and U14000 (N_14000,N_13232,N_13243);
and U14001 (N_14001,N_13931,N_13131);
or U14002 (N_14002,N_13135,N_13364);
nor U14003 (N_14003,N_13320,N_13404);
xor U14004 (N_14004,N_13401,N_13659);
nor U14005 (N_14005,N_13610,N_13115);
nor U14006 (N_14006,N_13923,N_13684);
or U14007 (N_14007,N_13379,N_13191);
and U14008 (N_14008,N_13428,N_13479);
or U14009 (N_14009,N_13443,N_13454);
nor U14010 (N_14010,N_13398,N_13621);
or U14011 (N_14011,N_13526,N_13468);
and U14012 (N_14012,N_13969,N_13742);
nor U14013 (N_14013,N_13590,N_13868);
nand U14014 (N_14014,N_13861,N_13540);
nor U14015 (N_14015,N_13520,N_13215);
and U14016 (N_14016,N_13903,N_13780);
nand U14017 (N_14017,N_13709,N_13460);
nor U14018 (N_14018,N_13328,N_13300);
and U14019 (N_14019,N_13285,N_13718);
and U14020 (N_14020,N_13832,N_13862);
or U14021 (N_14021,N_13272,N_13360);
nor U14022 (N_14022,N_13871,N_13252);
and U14023 (N_14023,N_13563,N_13533);
or U14024 (N_14024,N_13933,N_13095);
nor U14025 (N_14025,N_13568,N_13966);
or U14026 (N_14026,N_13086,N_13865);
or U14027 (N_14027,N_13519,N_13508);
nor U14028 (N_14028,N_13333,N_13151);
nor U14029 (N_14029,N_13196,N_13651);
nor U14030 (N_14030,N_13828,N_13737);
xor U14031 (N_14031,N_13623,N_13376);
nand U14032 (N_14032,N_13751,N_13426);
or U14033 (N_14033,N_13672,N_13525);
nor U14034 (N_14034,N_13775,N_13658);
nor U14035 (N_14035,N_13943,N_13466);
and U14036 (N_14036,N_13004,N_13318);
nand U14037 (N_14037,N_13820,N_13986);
nand U14038 (N_14038,N_13522,N_13815);
xor U14039 (N_14039,N_13819,N_13909);
or U14040 (N_14040,N_13993,N_13101);
nand U14041 (N_14041,N_13298,N_13812);
nand U14042 (N_14042,N_13773,N_13158);
or U14043 (N_14043,N_13889,N_13039);
and U14044 (N_14044,N_13805,N_13884);
and U14045 (N_14045,N_13997,N_13268);
xnor U14046 (N_14046,N_13160,N_13792);
nand U14047 (N_14047,N_13925,N_13237);
nand U14048 (N_14048,N_13384,N_13410);
nor U14049 (N_14049,N_13210,N_13098);
and U14050 (N_14050,N_13313,N_13995);
nand U14051 (N_14051,N_13484,N_13053);
xnor U14052 (N_14052,N_13938,N_13059);
xor U14053 (N_14053,N_13319,N_13735);
nor U14054 (N_14054,N_13412,N_13302);
xor U14055 (N_14055,N_13743,N_13589);
nor U14056 (N_14056,N_13014,N_13717);
nand U14057 (N_14057,N_13619,N_13885);
xnor U14058 (N_14058,N_13130,N_13570);
nand U14059 (N_14059,N_13397,N_13114);
nand U14060 (N_14060,N_13099,N_13470);
nor U14061 (N_14061,N_13258,N_13498);
nor U14062 (N_14062,N_13827,N_13758);
nand U14063 (N_14063,N_13070,N_13557);
xor U14064 (N_14064,N_13297,N_13048);
xnor U14065 (N_14065,N_13680,N_13779);
nor U14066 (N_14066,N_13389,N_13976);
xnor U14067 (N_14067,N_13963,N_13283);
and U14068 (N_14068,N_13399,N_13562);
nor U14069 (N_14069,N_13878,N_13908);
or U14070 (N_14070,N_13181,N_13808);
nor U14071 (N_14071,N_13441,N_13572);
and U14072 (N_14072,N_13173,N_13795);
or U14073 (N_14073,N_13852,N_13016);
nand U14074 (N_14074,N_13536,N_13281);
nand U14075 (N_14075,N_13712,N_13670);
nand U14076 (N_14076,N_13287,N_13388);
nor U14077 (N_14077,N_13632,N_13643);
or U14078 (N_14078,N_13834,N_13661);
nor U14079 (N_14079,N_13574,N_13041);
nand U14080 (N_14080,N_13509,N_13683);
and U14081 (N_14081,N_13853,N_13161);
xor U14082 (N_14082,N_13125,N_13618);
or U14083 (N_14083,N_13825,N_13940);
nor U14084 (N_14084,N_13662,N_13061);
and U14085 (N_14085,N_13087,N_13080);
xor U14086 (N_14086,N_13420,N_13761);
xnor U14087 (N_14087,N_13981,N_13065);
or U14088 (N_14088,N_13624,N_13797);
nand U14089 (N_14089,N_13549,N_13387);
xor U14090 (N_14090,N_13858,N_13178);
or U14091 (N_14091,N_13935,N_13156);
nor U14092 (N_14092,N_13481,N_13524);
or U14093 (N_14093,N_13992,N_13596);
nor U14094 (N_14094,N_13107,N_13576);
nor U14095 (N_14095,N_13749,N_13924);
nor U14096 (N_14096,N_13382,N_13840);
and U14097 (N_14097,N_13959,N_13111);
xnor U14098 (N_14098,N_13888,N_13301);
xor U14099 (N_14099,N_13127,N_13257);
nor U14100 (N_14100,N_13042,N_13594);
nor U14101 (N_14101,N_13582,N_13807);
xor U14102 (N_14102,N_13902,N_13406);
and U14103 (N_14103,N_13571,N_13702);
and U14104 (N_14104,N_13506,N_13162);
nand U14105 (N_14105,N_13091,N_13960);
nor U14106 (N_14106,N_13078,N_13906);
nor U14107 (N_14107,N_13607,N_13036);
nor U14108 (N_14108,N_13645,N_13710);
and U14109 (N_14109,N_13421,N_13493);
or U14110 (N_14110,N_13803,N_13821);
or U14111 (N_14111,N_13381,N_13011);
nor U14112 (N_14112,N_13879,N_13788);
nand U14113 (N_14113,N_13308,N_13566);
nor U14114 (N_14114,N_13961,N_13018);
nor U14115 (N_14115,N_13510,N_13128);
or U14116 (N_14116,N_13979,N_13598);
xnor U14117 (N_14117,N_13244,N_13748);
and U14118 (N_14118,N_13818,N_13891);
nor U14119 (N_14119,N_13372,N_13019);
and U14120 (N_14120,N_13869,N_13642);
nand U14121 (N_14121,N_13093,N_13250);
xnor U14122 (N_14122,N_13882,N_13505);
or U14123 (N_14123,N_13072,N_13263);
and U14124 (N_14124,N_13309,N_13793);
nor U14125 (N_14125,N_13289,N_13330);
or U14126 (N_14126,N_13267,N_13535);
nand U14127 (N_14127,N_13760,N_13343);
nor U14128 (N_14128,N_13660,N_13732);
nand U14129 (N_14129,N_13770,N_13189);
and U14130 (N_14130,N_13789,N_13299);
nor U14131 (N_14131,N_13031,N_13425);
nor U14132 (N_14132,N_13523,N_13024);
or U14133 (N_14133,N_13546,N_13787);
nand U14134 (N_14134,N_13687,N_13198);
nand U14135 (N_14135,N_13886,N_13154);
and U14136 (N_14136,N_13930,N_13242);
or U14137 (N_14137,N_13491,N_13895);
xnor U14138 (N_14138,N_13634,N_13715);
and U14139 (N_14139,N_13591,N_13140);
nand U14140 (N_14140,N_13214,N_13306);
nor U14141 (N_14141,N_13430,N_13476);
or U14142 (N_14142,N_13141,N_13184);
or U14143 (N_14143,N_13463,N_13192);
nor U14144 (N_14144,N_13144,N_13530);
nor U14145 (N_14145,N_13073,N_13152);
or U14146 (N_14146,N_13276,N_13143);
and U14147 (N_14147,N_13734,N_13553);
nor U14148 (N_14148,N_13007,N_13423);
or U14149 (N_14149,N_13385,N_13456);
and U14150 (N_14150,N_13056,N_13714);
nand U14151 (N_14151,N_13068,N_13545);
nor U14152 (N_14152,N_13612,N_13097);
nand U14153 (N_14153,N_13453,N_13337);
or U14154 (N_14154,N_13835,N_13855);
nor U14155 (N_14155,N_13544,N_13394);
nor U14156 (N_14156,N_13405,N_13890);
xor U14157 (N_14157,N_13916,N_13987);
xor U14158 (N_14158,N_13691,N_13123);
or U14159 (N_14159,N_13824,N_13222);
and U14160 (N_14160,N_13677,N_13926);
xor U14161 (N_14161,N_13846,N_13839);
and U14162 (N_14162,N_13164,N_13977);
nand U14163 (N_14163,N_13230,N_13640);
nor U14164 (N_14164,N_13802,N_13555);
nor U14165 (N_14165,N_13109,N_13754);
and U14166 (N_14166,N_13648,N_13904);
nor U14167 (N_14167,N_13418,N_13548);
nand U14168 (N_14168,N_13870,N_13175);
and U14169 (N_14169,N_13062,N_13325);
or U14170 (N_14170,N_13488,N_13312);
nor U14171 (N_14171,N_13928,N_13696);
nand U14172 (N_14172,N_13573,N_13336);
nand U14173 (N_14173,N_13608,N_13338);
and U14174 (N_14174,N_13124,N_13217);
nand U14175 (N_14175,N_13705,N_13501);
nor U14176 (N_14176,N_13438,N_13772);
or U14177 (N_14177,N_13293,N_13584);
and U14178 (N_14178,N_13370,N_13875);
or U14179 (N_14179,N_13752,N_13502);
or U14180 (N_14180,N_13729,N_13850);
or U14181 (N_14181,N_13583,N_13390);
or U14182 (N_14182,N_13255,N_13517);
nor U14183 (N_14183,N_13409,N_13915);
or U14184 (N_14184,N_13616,N_13681);
xnor U14185 (N_14185,N_13918,N_13414);
or U14186 (N_14186,N_13764,N_13686);
nand U14187 (N_14187,N_13881,N_13528);
or U14188 (N_14188,N_13431,N_13894);
or U14189 (N_14189,N_13203,N_13781);
or U14190 (N_14190,N_13166,N_13323);
nor U14191 (N_14191,N_13006,N_13471);
nor U14192 (N_14192,N_13311,N_13708);
nor U14193 (N_14193,N_13380,N_13830);
nand U14194 (N_14194,N_13235,N_13613);
xor U14195 (N_14195,N_13733,N_13221);
nand U14196 (N_14196,N_13282,N_13633);
nand U14197 (N_14197,N_13701,N_13231);
xor U14198 (N_14198,N_13331,N_13190);
nor U14199 (N_14199,N_13201,N_13603);
or U14200 (N_14200,N_13393,N_13810);
and U14201 (N_14201,N_13182,N_13942);
nand U14202 (N_14202,N_13165,N_13483);
nor U14203 (N_14203,N_13216,N_13100);
xor U14204 (N_14204,N_13756,N_13265);
xnor U14205 (N_14205,N_13503,N_13679);
xor U14206 (N_14206,N_13635,N_13037);
or U14207 (N_14207,N_13082,N_13782);
and U14208 (N_14208,N_13447,N_13174);
and U14209 (N_14209,N_13266,N_13066);
and U14210 (N_14210,N_13801,N_13900);
and U14211 (N_14211,N_13450,N_13615);
nor U14212 (N_14212,N_13713,N_13515);
xnor U14213 (N_14213,N_13259,N_13464);
nand U14214 (N_14214,N_13090,N_13038);
nand U14215 (N_14215,N_13315,N_13367);
nand U14216 (N_14216,N_13249,N_13002);
and U14217 (N_14217,N_13046,N_13602);
and U14218 (N_14218,N_13075,N_13774);
xor U14219 (N_14219,N_13595,N_13085);
nor U14220 (N_14220,N_13740,N_13205);
and U14221 (N_14221,N_13759,N_13776);
nor U14222 (N_14222,N_13883,N_13836);
nor U14223 (N_14223,N_13543,N_13278);
xor U14224 (N_14224,N_13113,N_13357);
or U14225 (N_14225,N_13348,N_13392);
and U14226 (N_14226,N_13371,N_13951);
or U14227 (N_14227,N_13446,N_13682);
and U14228 (N_14228,N_13866,N_13044);
nand U14229 (N_14229,N_13726,N_13207);
and U14230 (N_14230,N_13295,N_13294);
or U14231 (N_14231,N_13587,N_13110);
and U14232 (N_14232,N_13863,N_13907);
and U14233 (N_14233,N_13722,N_13092);
nor U14234 (N_14234,N_13877,N_13697);
or U14235 (N_14235,N_13363,N_13274);
xor U14236 (N_14236,N_13204,N_13199);
or U14237 (N_14237,N_13206,N_13512);
and U14238 (N_14238,N_13170,N_13247);
or U14239 (N_14239,N_13334,N_13218);
nor U14240 (N_14240,N_13020,N_13332);
or U14241 (N_14241,N_13939,N_13153);
nor U14242 (N_14242,N_13197,N_13148);
or U14243 (N_14243,N_13213,N_13864);
nor U14244 (N_14244,N_13690,N_13800);
or U14245 (N_14245,N_13529,N_13996);
nor U14246 (N_14246,N_13435,N_13238);
and U14247 (N_14247,N_13872,N_13671);
and U14248 (N_14248,N_13054,N_13826);
xor U14249 (N_14249,N_13180,N_13606);
and U14250 (N_14250,N_13983,N_13703);
nor U14251 (N_14251,N_13187,N_13271);
nor U14252 (N_14252,N_13458,N_13035);
and U14253 (N_14253,N_13188,N_13669);
or U14254 (N_14254,N_13347,N_13777);
nor U14255 (N_14255,N_13822,N_13246);
and U14256 (N_14256,N_13952,N_13552);
and U14257 (N_14257,N_13351,N_13134);
nand U14258 (N_14258,N_13556,N_13550);
nand U14259 (N_14259,N_13208,N_13429);
and U14260 (N_14260,N_13688,N_13896);
nor U14261 (N_14261,N_13785,N_13771);
nor U14262 (N_14262,N_13728,N_13927);
and U14263 (N_14263,N_13946,N_13914);
and U14264 (N_14264,N_13142,N_13531);
or U14265 (N_14265,N_13767,N_13083);
xnor U14266 (N_14266,N_13920,N_13514);
nand U14267 (N_14267,N_13636,N_13487);
and U14268 (N_14268,N_13224,N_13383);
or U14269 (N_14269,N_13984,N_13980);
nand U14270 (N_14270,N_13848,N_13432);
xnor U14271 (N_14271,N_13999,N_13179);
xnor U14272 (N_14272,N_13245,N_13617);
nor U14273 (N_14273,N_13234,N_13211);
or U14274 (N_14274,N_13396,N_13547);
nand U14275 (N_14275,N_13029,N_13833);
or U14276 (N_14276,N_13736,N_13604);
nand U14277 (N_14277,N_13159,N_13727);
nand U14278 (N_14278,N_13240,N_13354);
xor U14279 (N_14279,N_13051,N_13622);
and U14280 (N_14280,N_13757,N_13851);
or U14281 (N_14281,N_13639,N_13474);
nand U14282 (N_14282,N_13724,N_13001);
nand U14283 (N_14283,N_13490,N_13079);
or U14284 (N_14284,N_13108,N_13579);
nor U14285 (N_14285,N_13813,N_13597);
xor U14286 (N_14286,N_13350,N_13798);
nand U14287 (N_14287,N_13442,N_13630);
and U14288 (N_14288,N_13588,N_13374);
nand U14289 (N_14289,N_13386,N_13436);
or U14290 (N_14290,N_13459,N_13316);
or U14291 (N_14291,N_13327,N_13653);
xnor U14292 (N_14292,N_13322,N_13880);
xnor U14293 (N_14293,N_13060,N_13559);
and U14294 (N_14294,N_13112,N_13032);
and U14295 (N_14295,N_13921,N_13058);
nor U14296 (N_14296,N_13183,N_13227);
nand U14297 (N_14297,N_13953,N_13893);
or U14298 (N_14298,N_13693,N_13857);
xnor U14299 (N_14299,N_13711,N_13071);
xnor U14300 (N_14300,N_13473,N_13292);
and U14301 (N_14301,N_13185,N_13346);
or U14302 (N_14302,N_13565,N_13150);
or U14303 (N_14303,N_13991,N_13403);
xnor U14304 (N_14304,N_13467,N_13650);
and U14305 (N_14305,N_13477,N_13149);
nand U14306 (N_14306,N_13202,N_13769);
xnor U14307 (N_14307,N_13972,N_13537);
or U14308 (N_14308,N_13362,N_13146);
nor U14309 (N_14309,N_13783,N_13273);
xor U14310 (N_14310,N_13129,N_13569);
or U14311 (N_14311,N_13700,N_13804);
nand U14312 (N_14312,N_13495,N_13122);
nor U14313 (N_14313,N_13950,N_13168);
nor U14314 (N_14314,N_13692,N_13500);
or U14315 (N_14315,N_13241,N_13133);
nor U14316 (N_14316,N_13567,N_13716);
xor U14317 (N_14317,N_13796,N_13448);
xnor U14318 (N_14318,N_13219,N_13668);
nand U14319 (N_14319,N_13874,N_13076);
nand U14320 (N_14320,N_13469,N_13694);
and U14321 (N_14321,N_13551,N_13970);
nor U14322 (N_14322,N_13407,N_13497);
nor U14323 (N_14323,N_13578,N_13982);
or U14324 (N_14324,N_13167,N_13262);
and U14325 (N_14325,N_13369,N_13867);
nand U14326 (N_14326,N_13492,N_13317);
or U14327 (N_14327,N_13286,N_13366);
and U14328 (N_14328,N_13947,N_13532);
nor U14329 (N_14329,N_13419,N_13067);
xor U14330 (N_14330,N_13955,N_13345);
nor U14331 (N_14331,N_13675,N_13934);
and U14332 (N_14332,N_13744,N_13088);
xor U14333 (N_14333,N_13462,N_13000);
xnor U14334 (N_14334,N_13009,N_13676);
nor U14335 (N_14335,N_13195,N_13706);
or U14336 (N_14336,N_13978,N_13342);
xnor U14337 (N_14337,N_13905,N_13937);
nor U14338 (N_14338,N_13849,N_13010);
xnor U14339 (N_14339,N_13814,N_13898);
and U14340 (N_14340,N_13220,N_13593);
nor U14341 (N_14341,N_13964,N_13339);
nor U14342 (N_14342,N_13956,N_13022);
or U14343 (N_14343,N_13324,N_13280);
and U14344 (N_14344,N_13200,N_13538);
nor U14345 (N_14345,N_13120,N_13081);
xor U14346 (N_14346,N_13784,N_13599);
xor U14347 (N_14347,N_13015,N_13269);
nor U14348 (N_14348,N_13028,N_13239);
nor U14349 (N_14349,N_13541,N_13177);
nor U14350 (N_14350,N_13228,N_13626);
and U14351 (N_14351,N_13030,N_13457);
or U14352 (N_14352,N_13845,N_13912);
nor U14353 (N_14353,N_13816,N_13911);
xor U14354 (N_14354,N_13747,N_13652);
xnor U14355 (N_14355,N_13138,N_13719);
xor U14356 (N_14356,N_13288,N_13254);
nor U14357 (N_14357,N_13725,N_13155);
or U14358 (N_14358,N_13077,N_13194);
xor U14359 (N_14359,N_13439,N_13766);
nand U14360 (N_14360,N_13415,N_13577);
xnor U14361 (N_14361,N_13609,N_13416);
or U14362 (N_14362,N_13627,N_13695);
or U14363 (N_14363,N_13145,N_13434);
or U14364 (N_14364,N_13856,N_13985);
and U14365 (N_14365,N_13395,N_13012);
nand U14366 (N_14366,N_13063,N_13307);
or U14367 (N_14367,N_13496,N_13365);
nor U14368 (N_14368,N_13482,N_13990);
and U14369 (N_14369,N_13945,N_13600);
nor U14370 (N_14370,N_13860,N_13975);
or U14371 (N_14371,N_13356,N_13417);
nand U14372 (N_14372,N_13017,N_13794);
nor U14373 (N_14373,N_13741,N_13817);
xor U14374 (N_14374,N_13229,N_13023);
nor U14375 (N_14375,N_13738,N_13910);
xnor U14376 (N_14376,N_13994,N_13507);
nor U14377 (N_14377,N_13455,N_13629);
nor U14378 (N_14378,N_13137,N_13136);
nand U14379 (N_14379,N_13251,N_13437);
xnor U14380 (N_14380,N_13005,N_13806);
or U14381 (N_14381,N_13261,N_13326);
or U14382 (N_14382,N_13043,N_13791);
xor U14383 (N_14383,N_13433,N_13226);
nand U14384 (N_14384,N_13637,N_13290);
and U14385 (N_14385,N_13040,N_13971);
or U14386 (N_14386,N_13919,N_13413);
and U14387 (N_14387,N_13277,N_13126);
nand U14388 (N_14388,N_13663,N_13303);
and U14389 (N_14389,N_13361,N_13516);
nand U14390 (N_14390,N_13103,N_13049);
xnor U14391 (N_14391,N_13586,N_13768);
xor U14392 (N_14392,N_13698,N_13223);
xor U14393 (N_14393,N_13799,N_13304);
or U14394 (N_14394,N_13892,N_13378);
xnor U14395 (N_14395,N_13045,N_13233);
nand U14396 (N_14396,N_13341,N_13270);
xor U14397 (N_14397,N_13723,N_13033);
xnor U14398 (N_14398,N_13753,N_13605);
nor U14399 (N_14399,N_13314,N_13451);
nand U14400 (N_14400,N_13638,N_13352);
xor U14401 (N_14401,N_13968,N_13932);
nand U14402 (N_14402,N_13485,N_13678);
xnor U14403 (N_14403,N_13400,N_13034);
and U14404 (N_14404,N_13873,N_13518);
nand U14405 (N_14405,N_13534,N_13344);
and U14406 (N_14406,N_13132,N_13922);
or U14407 (N_14407,N_13193,N_13611);
xnor U14408 (N_14408,N_13452,N_13656);
or U14409 (N_14409,N_13831,N_13008);
nor U14410 (N_14410,N_13209,N_13117);
nand U14411 (N_14411,N_13628,N_13765);
or U14412 (N_14412,N_13842,N_13465);
and U14413 (N_14413,N_13854,N_13998);
nand U14414 (N_14414,N_13913,N_13897);
nor U14415 (N_14415,N_13105,N_13340);
nand U14416 (N_14416,N_13731,N_13424);
and U14417 (N_14417,N_13472,N_13929);
and U14418 (N_14418,N_13657,N_13585);
nand U14419 (N_14419,N_13762,N_13260);
or U14420 (N_14420,N_13564,N_13427);
nor U14421 (N_14421,N_13561,N_13475);
nor U14422 (N_14422,N_13284,N_13704);
xor U14423 (N_14423,N_13358,N_13989);
nand U14424 (N_14424,N_13157,N_13368);
nor U14425 (N_14425,N_13655,N_13844);
nor U14426 (N_14426,N_13186,N_13026);
or U14427 (N_14427,N_13958,N_13377);
xnor U14428 (N_14428,N_13335,N_13355);
nand U14429 (N_14429,N_13411,N_13236);
or U14430 (N_14430,N_13592,N_13746);
xor U14431 (N_14431,N_13169,N_13027);
xor U14432 (N_14432,N_13375,N_13121);
or U14433 (N_14433,N_13391,N_13494);
xor U14434 (N_14434,N_13253,N_13601);
or U14435 (N_14435,N_13664,N_13809);
xnor U14436 (N_14436,N_13422,N_13461);
xnor U14437 (N_14437,N_13449,N_13305);
or U14438 (N_14438,N_13790,N_13876);
nor U14439 (N_14439,N_13838,N_13673);
nor U14440 (N_14440,N_13847,N_13139);
nand U14441 (N_14441,N_13118,N_13859);
nand U14442 (N_14442,N_13147,N_13811);
and U14443 (N_14443,N_13094,N_13013);
xor U14444 (N_14444,N_13580,N_13649);
and U14445 (N_14445,N_13402,N_13967);
and U14446 (N_14446,N_13665,N_13954);
nand U14447 (N_14447,N_13256,N_13685);
nor U14448 (N_14448,N_13069,N_13349);
nand U14449 (N_14449,N_13620,N_13212);
or U14450 (N_14450,N_13843,N_13965);
nor U14451 (N_14451,N_13225,N_13641);
nand U14452 (N_14452,N_13089,N_13944);
nor U14453 (N_14453,N_13321,N_13296);
nand U14454 (N_14454,N_13310,N_13106);
nor U14455 (N_14455,N_13064,N_13291);
or U14456 (N_14456,N_13521,N_13763);
and U14457 (N_14457,N_13899,N_13050);
nand U14458 (N_14458,N_13096,N_13554);
nand U14459 (N_14459,N_13674,N_13988);
nand U14460 (N_14460,N_13558,N_13074);
or U14461 (N_14461,N_13575,N_13445);
nand U14462 (N_14462,N_13666,N_13499);
and U14463 (N_14463,N_13539,N_13699);
nor U14464 (N_14464,N_13480,N_13973);
nor U14465 (N_14465,N_13755,N_13279);
nand U14466 (N_14466,N_13511,N_13948);
and U14467 (N_14467,N_13614,N_13778);
nand U14468 (N_14468,N_13329,N_13936);
and U14469 (N_14469,N_13084,N_13730);
nand U14470 (N_14470,N_13631,N_13025);
or U14471 (N_14471,N_13841,N_13052);
and U14472 (N_14472,N_13823,N_13172);
nand U14473 (N_14473,N_13962,N_13102);
xor U14474 (N_14474,N_13957,N_13542);
nand U14475 (N_14475,N_13644,N_13003);
xor U14476 (N_14476,N_13707,N_13513);
nand U14477 (N_14477,N_13489,N_13047);
nor U14478 (N_14478,N_13408,N_13901);
nor U14479 (N_14479,N_13647,N_13264);
xnor U14480 (N_14480,N_13104,N_13654);
nand U14481 (N_14481,N_13055,N_13353);
xnor U14482 (N_14482,N_13440,N_13119);
or U14483 (N_14483,N_13829,N_13667);
or U14484 (N_14484,N_13373,N_13176);
xor U14485 (N_14485,N_13275,N_13887);
xor U14486 (N_14486,N_13750,N_13745);
nor U14487 (N_14487,N_13837,N_13721);
or U14488 (N_14488,N_13057,N_13478);
or U14489 (N_14489,N_13486,N_13917);
nand U14490 (N_14490,N_13116,N_13689);
or U14491 (N_14491,N_13444,N_13581);
nor U14492 (N_14492,N_13646,N_13504);
nor U14493 (N_14493,N_13560,N_13949);
or U14494 (N_14494,N_13163,N_13720);
nand U14495 (N_14495,N_13248,N_13739);
nor U14496 (N_14496,N_13941,N_13359);
and U14497 (N_14497,N_13974,N_13625);
xnor U14498 (N_14498,N_13786,N_13527);
or U14499 (N_14499,N_13021,N_13171);
nor U14500 (N_14500,N_13445,N_13531);
nor U14501 (N_14501,N_13637,N_13360);
or U14502 (N_14502,N_13485,N_13891);
nor U14503 (N_14503,N_13899,N_13369);
or U14504 (N_14504,N_13415,N_13354);
nand U14505 (N_14505,N_13203,N_13624);
xor U14506 (N_14506,N_13181,N_13682);
nor U14507 (N_14507,N_13496,N_13678);
nor U14508 (N_14508,N_13361,N_13520);
nand U14509 (N_14509,N_13840,N_13014);
or U14510 (N_14510,N_13147,N_13904);
or U14511 (N_14511,N_13913,N_13270);
xnor U14512 (N_14512,N_13314,N_13537);
xnor U14513 (N_14513,N_13125,N_13290);
xor U14514 (N_14514,N_13434,N_13838);
nor U14515 (N_14515,N_13987,N_13564);
and U14516 (N_14516,N_13758,N_13655);
and U14517 (N_14517,N_13646,N_13118);
and U14518 (N_14518,N_13552,N_13537);
xnor U14519 (N_14519,N_13097,N_13483);
and U14520 (N_14520,N_13742,N_13108);
or U14521 (N_14521,N_13991,N_13158);
and U14522 (N_14522,N_13661,N_13647);
xnor U14523 (N_14523,N_13780,N_13913);
or U14524 (N_14524,N_13959,N_13741);
nand U14525 (N_14525,N_13584,N_13699);
xor U14526 (N_14526,N_13034,N_13085);
or U14527 (N_14527,N_13855,N_13388);
or U14528 (N_14528,N_13866,N_13519);
and U14529 (N_14529,N_13780,N_13760);
or U14530 (N_14530,N_13118,N_13315);
nor U14531 (N_14531,N_13486,N_13866);
nand U14532 (N_14532,N_13268,N_13544);
or U14533 (N_14533,N_13966,N_13185);
and U14534 (N_14534,N_13610,N_13888);
nor U14535 (N_14535,N_13076,N_13052);
or U14536 (N_14536,N_13362,N_13289);
or U14537 (N_14537,N_13385,N_13714);
and U14538 (N_14538,N_13765,N_13037);
xnor U14539 (N_14539,N_13585,N_13441);
or U14540 (N_14540,N_13641,N_13972);
nand U14541 (N_14541,N_13615,N_13098);
nor U14542 (N_14542,N_13376,N_13986);
nand U14543 (N_14543,N_13401,N_13463);
nor U14544 (N_14544,N_13215,N_13389);
or U14545 (N_14545,N_13025,N_13502);
xor U14546 (N_14546,N_13112,N_13810);
nand U14547 (N_14547,N_13139,N_13904);
and U14548 (N_14548,N_13723,N_13697);
xnor U14549 (N_14549,N_13905,N_13768);
and U14550 (N_14550,N_13812,N_13210);
and U14551 (N_14551,N_13502,N_13268);
xor U14552 (N_14552,N_13517,N_13734);
nor U14553 (N_14553,N_13026,N_13878);
and U14554 (N_14554,N_13404,N_13555);
or U14555 (N_14555,N_13902,N_13130);
and U14556 (N_14556,N_13596,N_13644);
nor U14557 (N_14557,N_13888,N_13587);
nand U14558 (N_14558,N_13847,N_13716);
nand U14559 (N_14559,N_13447,N_13806);
nand U14560 (N_14560,N_13979,N_13146);
nor U14561 (N_14561,N_13183,N_13189);
xnor U14562 (N_14562,N_13636,N_13804);
xnor U14563 (N_14563,N_13126,N_13181);
nand U14564 (N_14564,N_13236,N_13177);
nor U14565 (N_14565,N_13568,N_13745);
nand U14566 (N_14566,N_13806,N_13122);
nand U14567 (N_14567,N_13623,N_13530);
and U14568 (N_14568,N_13721,N_13604);
xnor U14569 (N_14569,N_13985,N_13611);
nor U14570 (N_14570,N_13080,N_13256);
and U14571 (N_14571,N_13537,N_13943);
or U14572 (N_14572,N_13961,N_13108);
or U14573 (N_14573,N_13870,N_13288);
nor U14574 (N_14574,N_13206,N_13167);
and U14575 (N_14575,N_13573,N_13410);
nor U14576 (N_14576,N_13050,N_13897);
xnor U14577 (N_14577,N_13585,N_13991);
or U14578 (N_14578,N_13184,N_13423);
nor U14579 (N_14579,N_13775,N_13066);
nand U14580 (N_14580,N_13335,N_13623);
or U14581 (N_14581,N_13764,N_13025);
or U14582 (N_14582,N_13728,N_13316);
and U14583 (N_14583,N_13278,N_13164);
or U14584 (N_14584,N_13220,N_13889);
nor U14585 (N_14585,N_13145,N_13647);
xnor U14586 (N_14586,N_13496,N_13644);
nor U14587 (N_14587,N_13413,N_13753);
nand U14588 (N_14588,N_13039,N_13886);
nor U14589 (N_14589,N_13693,N_13449);
nor U14590 (N_14590,N_13891,N_13480);
nor U14591 (N_14591,N_13215,N_13091);
xor U14592 (N_14592,N_13821,N_13879);
nor U14593 (N_14593,N_13302,N_13618);
and U14594 (N_14594,N_13675,N_13464);
xnor U14595 (N_14595,N_13317,N_13927);
or U14596 (N_14596,N_13608,N_13146);
xnor U14597 (N_14597,N_13617,N_13863);
xor U14598 (N_14598,N_13464,N_13083);
or U14599 (N_14599,N_13277,N_13377);
nor U14600 (N_14600,N_13337,N_13571);
nand U14601 (N_14601,N_13402,N_13098);
nor U14602 (N_14602,N_13710,N_13739);
xnor U14603 (N_14603,N_13853,N_13736);
or U14604 (N_14604,N_13193,N_13607);
nand U14605 (N_14605,N_13591,N_13432);
nor U14606 (N_14606,N_13362,N_13751);
or U14607 (N_14607,N_13081,N_13258);
and U14608 (N_14608,N_13180,N_13260);
and U14609 (N_14609,N_13884,N_13094);
xnor U14610 (N_14610,N_13714,N_13183);
or U14611 (N_14611,N_13114,N_13102);
nor U14612 (N_14612,N_13779,N_13224);
xnor U14613 (N_14613,N_13075,N_13696);
or U14614 (N_14614,N_13010,N_13966);
or U14615 (N_14615,N_13379,N_13076);
nand U14616 (N_14616,N_13882,N_13312);
and U14617 (N_14617,N_13326,N_13350);
nor U14618 (N_14618,N_13285,N_13032);
nand U14619 (N_14619,N_13366,N_13712);
nor U14620 (N_14620,N_13312,N_13371);
or U14621 (N_14621,N_13547,N_13520);
nand U14622 (N_14622,N_13830,N_13878);
xnor U14623 (N_14623,N_13730,N_13106);
or U14624 (N_14624,N_13598,N_13223);
xnor U14625 (N_14625,N_13530,N_13270);
or U14626 (N_14626,N_13614,N_13741);
or U14627 (N_14627,N_13351,N_13641);
and U14628 (N_14628,N_13156,N_13800);
or U14629 (N_14629,N_13168,N_13895);
and U14630 (N_14630,N_13246,N_13342);
nand U14631 (N_14631,N_13905,N_13098);
and U14632 (N_14632,N_13545,N_13394);
nand U14633 (N_14633,N_13253,N_13468);
nor U14634 (N_14634,N_13937,N_13371);
xor U14635 (N_14635,N_13040,N_13723);
and U14636 (N_14636,N_13458,N_13526);
nor U14637 (N_14637,N_13769,N_13155);
or U14638 (N_14638,N_13241,N_13790);
and U14639 (N_14639,N_13868,N_13333);
and U14640 (N_14640,N_13890,N_13230);
xor U14641 (N_14641,N_13924,N_13878);
nand U14642 (N_14642,N_13792,N_13737);
or U14643 (N_14643,N_13496,N_13169);
and U14644 (N_14644,N_13247,N_13252);
nor U14645 (N_14645,N_13904,N_13029);
xnor U14646 (N_14646,N_13788,N_13903);
nor U14647 (N_14647,N_13435,N_13630);
nor U14648 (N_14648,N_13157,N_13209);
nand U14649 (N_14649,N_13166,N_13109);
nor U14650 (N_14650,N_13093,N_13122);
or U14651 (N_14651,N_13657,N_13779);
or U14652 (N_14652,N_13881,N_13005);
and U14653 (N_14653,N_13356,N_13988);
nand U14654 (N_14654,N_13776,N_13992);
nor U14655 (N_14655,N_13555,N_13894);
nand U14656 (N_14656,N_13014,N_13124);
nor U14657 (N_14657,N_13186,N_13316);
xnor U14658 (N_14658,N_13573,N_13510);
and U14659 (N_14659,N_13358,N_13825);
nand U14660 (N_14660,N_13126,N_13906);
nor U14661 (N_14661,N_13150,N_13847);
nand U14662 (N_14662,N_13113,N_13822);
xnor U14663 (N_14663,N_13618,N_13732);
and U14664 (N_14664,N_13536,N_13128);
nand U14665 (N_14665,N_13810,N_13883);
nand U14666 (N_14666,N_13011,N_13494);
or U14667 (N_14667,N_13537,N_13882);
nand U14668 (N_14668,N_13175,N_13948);
nor U14669 (N_14669,N_13306,N_13695);
nand U14670 (N_14670,N_13551,N_13898);
and U14671 (N_14671,N_13633,N_13169);
nor U14672 (N_14672,N_13234,N_13628);
or U14673 (N_14673,N_13333,N_13440);
or U14674 (N_14674,N_13116,N_13702);
or U14675 (N_14675,N_13543,N_13364);
nor U14676 (N_14676,N_13294,N_13536);
and U14677 (N_14677,N_13700,N_13803);
and U14678 (N_14678,N_13055,N_13870);
and U14679 (N_14679,N_13413,N_13669);
nand U14680 (N_14680,N_13659,N_13557);
nand U14681 (N_14681,N_13037,N_13771);
nor U14682 (N_14682,N_13198,N_13808);
xnor U14683 (N_14683,N_13895,N_13709);
xor U14684 (N_14684,N_13047,N_13469);
or U14685 (N_14685,N_13558,N_13372);
nand U14686 (N_14686,N_13400,N_13448);
nor U14687 (N_14687,N_13103,N_13516);
or U14688 (N_14688,N_13743,N_13552);
xnor U14689 (N_14689,N_13158,N_13384);
xnor U14690 (N_14690,N_13292,N_13998);
or U14691 (N_14691,N_13568,N_13900);
and U14692 (N_14692,N_13333,N_13040);
nor U14693 (N_14693,N_13084,N_13346);
xor U14694 (N_14694,N_13749,N_13695);
or U14695 (N_14695,N_13025,N_13527);
or U14696 (N_14696,N_13653,N_13726);
nor U14697 (N_14697,N_13751,N_13470);
xnor U14698 (N_14698,N_13708,N_13429);
xnor U14699 (N_14699,N_13315,N_13374);
nand U14700 (N_14700,N_13093,N_13267);
and U14701 (N_14701,N_13979,N_13070);
xor U14702 (N_14702,N_13628,N_13499);
nand U14703 (N_14703,N_13171,N_13148);
xor U14704 (N_14704,N_13667,N_13014);
and U14705 (N_14705,N_13626,N_13099);
nand U14706 (N_14706,N_13350,N_13402);
and U14707 (N_14707,N_13909,N_13231);
and U14708 (N_14708,N_13478,N_13746);
nor U14709 (N_14709,N_13967,N_13253);
xnor U14710 (N_14710,N_13611,N_13570);
and U14711 (N_14711,N_13943,N_13215);
xor U14712 (N_14712,N_13414,N_13608);
and U14713 (N_14713,N_13241,N_13259);
and U14714 (N_14714,N_13608,N_13104);
and U14715 (N_14715,N_13767,N_13700);
nand U14716 (N_14716,N_13605,N_13944);
xnor U14717 (N_14717,N_13974,N_13293);
xor U14718 (N_14718,N_13144,N_13848);
nor U14719 (N_14719,N_13983,N_13922);
and U14720 (N_14720,N_13218,N_13427);
or U14721 (N_14721,N_13691,N_13954);
nand U14722 (N_14722,N_13023,N_13777);
nand U14723 (N_14723,N_13629,N_13505);
nand U14724 (N_14724,N_13808,N_13336);
xnor U14725 (N_14725,N_13310,N_13318);
nor U14726 (N_14726,N_13209,N_13127);
nand U14727 (N_14727,N_13010,N_13240);
xor U14728 (N_14728,N_13495,N_13179);
or U14729 (N_14729,N_13872,N_13000);
or U14730 (N_14730,N_13509,N_13589);
xnor U14731 (N_14731,N_13836,N_13660);
xnor U14732 (N_14732,N_13424,N_13627);
nor U14733 (N_14733,N_13352,N_13699);
nor U14734 (N_14734,N_13453,N_13361);
and U14735 (N_14735,N_13537,N_13864);
nor U14736 (N_14736,N_13226,N_13963);
nor U14737 (N_14737,N_13492,N_13988);
and U14738 (N_14738,N_13658,N_13582);
nor U14739 (N_14739,N_13016,N_13703);
and U14740 (N_14740,N_13939,N_13894);
or U14741 (N_14741,N_13142,N_13472);
and U14742 (N_14742,N_13940,N_13089);
nand U14743 (N_14743,N_13043,N_13194);
xnor U14744 (N_14744,N_13258,N_13190);
nand U14745 (N_14745,N_13911,N_13966);
or U14746 (N_14746,N_13737,N_13578);
and U14747 (N_14747,N_13371,N_13083);
or U14748 (N_14748,N_13437,N_13607);
and U14749 (N_14749,N_13850,N_13930);
xnor U14750 (N_14750,N_13923,N_13218);
nor U14751 (N_14751,N_13782,N_13483);
nor U14752 (N_14752,N_13593,N_13353);
nor U14753 (N_14753,N_13176,N_13769);
nand U14754 (N_14754,N_13184,N_13257);
nor U14755 (N_14755,N_13536,N_13095);
or U14756 (N_14756,N_13693,N_13884);
or U14757 (N_14757,N_13763,N_13753);
nand U14758 (N_14758,N_13033,N_13058);
or U14759 (N_14759,N_13063,N_13925);
xor U14760 (N_14760,N_13526,N_13500);
or U14761 (N_14761,N_13051,N_13461);
and U14762 (N_14762,N_13929,N_13696);
nand U14763 (N_14763,N_13839,N_13478);
or U14764 (N_14764,N_13192,N_13054);
nor U14765 (N_14765,N_13303,N_13367);
nor U14766 (N_14766,N_13816,N_13818);
nand U14767 (N_14767,N_13425,N_13263);
and U14768 (N_14768,N_13757,N_13010);
and U14769 (N_14769,N_13609,N_13633);
xnor U14770 (N_14770,N_13434,N_13897);
and U14771 (N_14771,N_13392,N_13736);
and U14772 (N_14772,N_13220,N_13254);
nand U14773 (N_14773,N_13964,N_13591);
xnor U14774 (N_14774,N_13434,N_13407);
or U14775 (N_14775,N_13421,N_13243);
and U14776 (N_14776,N_13899,N_13477);
or U14777 (N_14777,N_13016,N_13290);
nand U14778 (N_14778,N_13003,N_13494);
and U14779 (N_14779,N_13188,N_13819);
nand U14780 (N_14780,N_13174,N_13817);
or U14781 (N_14781,N_13417,N_13015);
xor U14782 (N_14782,N_13724,N_13946);
nor U14783 (N_14783,N_13536,N_13269);
or U14784 (N_14784,N_13380,N_13509);
nor U14785 (N_14785,N_13966,N_13069);
and U14786 (N_14786,N_13003,N_13646);
and U14787 (N_14787,N_13199,N_13468);
xor U14788 (N_14788,N_13082,N_13622);
xor U14789 (N_14789,N_13339,N_13469);
or U14790 (N_14790,N_13188,N_13695);
xor U14791 (N_14791,N_13570,N_13626);
nand U14792 (N_14792,N_13545,N_13992);
nor U14793 (N_14793,N_13118,N_13604);
or U14794 (N_14794,N_13211,N_13939);
nor U14795 (N_14795,N_13095,N_13038);
nor U14796 (N_14796,N_13085,N_13678);
nand U14797 (N_14797,N_13851,N_13272);
xor U14798 (N_14798,N_13136,N_13209);
nor U14799 (N_14799,N_13758,N_13545);
or U14800 (N_14800,N_13249,N_13829);
or U14801 (N_14801,N_13343,N_13682);
and U14802 (N_14802,N_13215,N_13879);
nand U14803 (N_14803,N_13590,N_13735);
xor U14804 (N_14804,N_13059,N_13173);
nand U14805 (N_14805,N_13270,N_13285);
or U14806 (N_14806,N_13607,N_13113);
and U14807 (N_14807,N_13588,N_13462);
nand U14808 (N_14808,N_13050,N_13110);
or U14809 (N_14809,N_13766,N_13851);
and U14810 (N_14810,N_13037,N_13093);
and U14811 (N_14811,N_13408,N_13697);
nand U14812 (N_14812,N_13172,N_13438);
nor U14813 (N_14813,N_13302,N_13344);
or U14814 (N_14814,N_13055,N_13307);
nand U14815 (N_14815,N_13660,N_13924);
nand U14816 (N_14816,N_13296,N_13745);
nand U14817 (N_14817,N_13544,N_13004);
xor U14818 (N_14818,N_13834,N_13579);
nand U14819 (N_14819,N_13861,N_13176);
xnor U14820 (N_14820,N_13329,N_13357);
nand U14821 (N_14821,N_13000,N_13610);
or U14822 (N_14822,N_13730,N_13138);
xor U14823 (N_14823,N_13382,N_13444);
nor U14824 (N_14824,N_13678,N_13693);
or U14825 (N_14825,N_13703,N_13491);
nand U14826 (N_14826,N_13411,N_13111);
nor U14827 (N_14827,N_13975,N_13539);
nand U14828 (N_14828,N_13438,N_13859);
xnor U14829 (N_14829,N_13493,N_13435);
nand U14830 (N_14830,N_13768,N_13116);
or U14831 (N_14831,N_13483,N_13448);
and U14832 (N_14832,N_13461,N_13270);
nor U14833 (N_14833,N_13793,N_13819);
xor U14834 (N_14834,N_13363,N_13024);
nor U14835 (N_14835,N_13322,N_13474);
and U14836 (N_14836,N_13468,N_13556);
nor U14837 (N_14837,N_13401,N_13452);
or U14838 (N_14838,N_13095,N_13378);
and U14839 (N_14839,N_13618,N_13149);
nand U14840 (N_14840,N_13131,N_13924);
nor U14841 (N_14841,N_13773,N_13951);
or U14842 (N_14842,N_13755,N_13951);
nand U14843 (N_14843,N_13301,N_13045);
nor U14844 (N_14844,N_13016,N_13366);
nand U14845 (N_14845,N_13369,N_13313);
nand U14846 (N_14846,N_13091,N_13011);
or U14847 (N_14847,N_13807,N_13584);
xor U14848 (N_14848,N_13717,N_13811);
or U14849 (N_14849,N_13202,N_13219);
and U14850 (N_14850,N_13384,N_13195);
or U14851 (N_14851,N_13603,N_13218);
or U14852 (N_14852,N_13965,N_13232);
or U14853 (N_14853,N_13101,N_13350);
or U14854 (N_14854,N_13860,N_13372);
nor U14855 (N_14855,N_13208,N_13392);
nor U14856 (N_14856,N_13199,N_13015);
nor U14857 (N_14857,N_13031,N_13178);
nor U14858 (N_14858,N_13008,N_13848);
nor U14859 (N_14859,N_13277,N_13508);
nor U14860 (N_14860,N_13175,N_13761);
nand U14861 (N_14861,N_13302,N_13542);
xnor U14862 (N_14862,N_13020,N_13695);
nor U14863 (N_14863,N_13315,N_13122);
or U14864 (N_14864,N_13294,N_13918);
xnor U14865 (N_14865,N_13809,N_13131);
xor U14866 (N_14866,N_13228,N_13763);
or U14867 (N_14867,N_13134,N_13617);
or U14868 (N_14868,N_13412,N_13976);
or U14869 (N_14869,N_13610,N_13826);
nor U14870 (N_14870,N_13664,N_13285);
xor U14871 (N_14871,N_13474,N_13248);
or U14872 (N_14872,N_13702,N_13440);
nand U14873 (N_14873,N_13311,N_13307);
nand U14874 (N_14874,N_13545,N_13983);
nand U14875 (N_14875,N_13310,N_13817);
or U14876 (N_14876,N_13663,N_13409);
xor U14877 (N_14877,N_13675,N_13195);
and U14878 (N_14878,N_13185,N_13857);
or U14879 (N_14879,N_13781,N_13538);
nand U14880 (N_14880,N_13731,N_13410);
nand U14881 (N_14881,N_13433,N_13862);
or U14882 (N_14882,N_13844,N_13928);
nor U14883 (N_14883,N_13424,N_13905);
and U14884 (N_14884,N_13452,N_13939);
and U14885 (N_14885,N_13686,N_13835);
or U14886 (N_14886,N_13056,N_13112);
and U14887 (N_14887,N_13971,N_13460);
nand U14888 (N_14888,N_13262,N_13585);
and U14889 (N_14889,N_13794,N_13049);
nand U14890 (N_14890,N_13878,N_13986);
or U14891 (N_14891,N_13460,N_13086);
nand U14892 (N_14892,N_13489,N_13175);
and U14893 (N_14893,N_13501,N_13465);
xor U14894 (N_14894,N_13883,N_13749);
nor U14895 (N_14895,N_13044,N_13404);
and U14896 (N_14896,N_13074,N_13011);
nor U14897 (N_14897,N_13384,N_13838);
xnor U14898 (N_14898,N_13899,N_13859);
xnor U14899 (N_14899,N_13866,N_13959);
nand U14900 (N_14900,N_13252,N_13406);
and U14901 (N_14901,N_13915,N_13444);
xor U14902 (N_14902,N_13403,N_13762);
xnor U14903 (N_14903,N_13742,N_13349);
and U14904 (N_14904,N_13780,N_13805);
nand U14905 (N_14905,N_13593,N_13543);
nor U14906 (N_14906,N_13982,N_13440);
nand U14907 (N_14907,N_13559,N_13532);
and U14908 (N_14908,N_13575,N_13647);
or U14909 (N_14909,N_13494,N_13080);
xnor U14910 (N_14910,N_13882,N_13610);
or U14911 (N_14911,N_13498,N_13418);
and U14912 (N_14912,N_13803,N_13333);
and U14913 (N_14913,N_13736,N_13187);
xor U14914 (N_14914,N_13246,N_13431);
or U14915 (N_14915,N_13460,N_13084);
xor U14916 (N_14916,N_13961,N_13826);
and U14917 (N_14917,N_13802,N_13687);
nor U14918 (N_14918,N_13277,N_13425);
or U14919 (N_14919,N_13293,N_13993);
and U14920 (N_14920,N_13472,N_13841);
nand U14921 (N_14921,N_13812,N_13954);
nor U14922 (N_14922,N_13085,N_13963);
nor U14923 (N_14923,N_13419,N_13226);
nand U14924 (N_14924,N_13983,N_13087);
nor U14925 (N_14925,N_13860,N_13690);
xnor U14926 (N_14926,N_13734,N_13467);
nand U14927 (N_14927,N_13787,N_13967);
xor U14928 (N_14928,N_13182,N_13475);
nor U14929 (N_14929,N_13721,N_13062);
and U14930 (N_14930,N_13443,N_13560);
or U14931 (N_14931,N_13583,N_13926);
or U14932 (N_14932,N_13431,N_13667);
nand U14933 (N_14933,N_13850,N_13915);
and U14934 (N_14934,N_13776,N_13180);
nand U14935 (N_14935,N_13717,N_13188);
xor U14936 (N_14936,N_13634,N_13800);
or U14937 (N_14937,N_13434,N_13465);
nand U14938 (N_14938,N_13064,N_13903);
nand U14939 (N_14939,N_13562,N_13242);
and U14940 (N_14940,N_13259,N_13545);
and U14941 (N_14941,N_13472,N_13763);
xor U14942 (N_14942,N_13646,N_13514);
nor U14943 (N_14943,N_13868,N_13386);
and U14944 (N_14944,N_13015,N_13682);
nor U14945 (N_14945,N_13783,N_13448);
and U14946 (N_14946,N_13553,N_13448);
or U14947 (N_14947,N_13586,N_13934);
nand U14948 (N_14948,N_13876,N_13065);
xnor U14949 (N_14949,N_13362,N_13951);
and U14950 (N_14950,N_13477,N_13067);
nand U14951 (N_14951,N_13568,N_13362);
and U14952 (N_14952,N_13804,N_13076);
nand U14953 (N_14953,N_13439,N_13800);
nand U14954 (N_14954,N_13869,N_13973);
and U14955 (N_14955,N_13749,N_13425);
nand U14956 (N_14956,N_13655,N_13112);
nor U14957 (N_14957,N_13264,N_13589);
nand U14958 (N_14958,N_13404,N_13856);
nor U14959 (N_14959,N_13382,N_13790);
or U14960 (N_14960,N_13473,N_13815);
xor U14961 (N_14961,N_13156,N_13200);
xnor U14962 (N_14962,N_13778,N_13303);
xnor U14963 (N_14963,N_13802,N_13071);
or U14964 (N_14964,N_13757,N_13080);
and U14965 (N_14965,N_13953,N_13142);
xnor U14966 (N_14966,N_13915,N_13496);
xnor U14967 (N_14967,N_13433,N_13734);
and U14968 (N_14968,N_13540,N_13453);
and U14969 (N_14969,N_13231,N_13092);
nor U14970 (N_14970,N_13534,N_13199);
nand U14971 (N_14971,N_13325,N_13237);
or U14972 (N_14972,N_13090,N_13802);
nand U14973 (N_14973,N_13932,N_13105);
or U14974 (N_14974,N_13997,N_13037);
or U14975 (N_14975,N_13569,N_13955);
and U14976 (N_14976,N_13671,N_13830);
and U14977 (N_14977,N_13327,N_13667);
or U14978 (N_14978,N_13284,N_13183);
or U14979 (N_14979,N_13541,N_13470);
nand U14980 (N_14980,N_13425,N_13159);
nor U14981 (N_14981,N_13954,N_13530);
or U14982 (N_14982,N_13129,N_13202);
xnor U14983 (N_14983,N_13985,N_13164);
nor U14984 (N_14984,N_13203,N_13633);
nand U14985 (N_14985,N_13498,N_13641);
xnor U14986 (N_14986,N_13769,N_13160);
or U14987 (N_14987,N_13782,N_13202);
and U14988 (N_14988,N_13570,N_13660);
xor U14989 (N_14989,N_13246,N_13243);
xnor U14990 (N_14990,N_13380,N_13852);
nand U14991 (N_14991,N_13630,N_13290);
nand U14992 (N_14992,N_13558,N_13466);
xor U14993 (N_14993,N_13780,N_13731);
or U14994 (N_14994,N_13719,N_13049);
or U14995 (N_14995,N_13354,N_13246);
nand U14996 (N_14996,N_13296,N_13114);
and U14997 (N_14997,N_13411,N_13903);
and U14998 (N_14998,N_13786,N_13497);
nand U14999 (N_14999,N_13704,N_13130);
and U15000 (N_15000,N_14792,N_14391);
xnor U15001 (N_15001,N_14971,N_14742);
and U15002 (N_15002,N_14621,N_14817);
nand U15003 (N_15003,N_14046,N_14016);
xnor U15004 (N_15004,N_14463,N_14900);
or U15005 (N_15005,N_14869,N_14289);
or U15006 (N_15006,N_14944,N_14131);
nor U15007 (N_15007,N_14117,N_14829);
nand U15008 (N_15008,N_14074,N_14411);
or U15009 (N_15009,N_14425,N_14753);
or U15010 (N_15010,N_14632,N_14918);
nor U15011 (N_15011,N_14053,N_14033);
or U15012 (N_15012,N_14433,N_14447);
xor U15013 (N_15013,N_14325,N_14474);
nor U15014 (N_15014,N_14269,N_14484);
nor U15015 (N_15015,N_14775,N_14594);
nor U15016 (N_15016,N_14418,N_14049);
and U15017 (N_15017,N_14809,N_14334);
and U15018 (N_15018,N_14952,N_14977);
and U15019 (N_15019,N_14277,N_14747);
or U15020 (N_15020,N_14109,N_14966);
and U15021 (N_15021,N_14057,N_14300);
or U15022 (N_15022,N_14865,N_14328);
nor U15023 (N_15023,N_14066,N_14663);
or U15024 (N_15024,N_14828,N_14667);
or U15025 (N_15025,N_14954,N_14853);
xor U15026 (N_15026,N_14628,N_14424);
xnor U15027 (N_15027,N_14989,N_14387);
nor U15028 (N_15028,N_14707,N_14654);
and U15029 (N_15029,N_14563,N_14575);
or U15030 (N_15030,N_14647,N_14838);
xnor U15031 (N_15031,N_14266,N_14452);
or U15032 (N_15032,N_14555,N_14513);
nor U15033 (N_15033,N_14741,N_14642);
nand U15034 (N_15034,N_14686,N_14991);
or U15035 (N_15035,N_14363,N_14261);
xnor U15036 (N_15036,N_14012,N_14490);
nand U15037 (N_15037,N_14920,N_14777);
and U15038 (N_15038,N_14728,N_14623);
xor U15039 (N_15039,N_14483,N_14950);
xnor U15040 (N_15040,N_14034,N_14441);
nor U15041 (N_15041,N_14079,N_14460);
nor U15042 (N_15042,N_14357,N_14873);
nand U15043 (N_15043,N_14048,N_14912);
and U15044 (N_15044,N_14037,N_14588);
or U15045 (N_15045,N_14488,N_14251);
or U15046 (N_15046,N_14038,N_14616);
and U15047 (N_15047,N_14135,N_14153);
xnor U15048 (N_15048,N_14604,N_14705);
nor U15049 (N_15049,N_14671,N_14749);
nand U15050 (N_15050,N_14400,N_14171);
nor U15051 (N_15051,N_14726,N_14580);
and U15052 (N_15052,N_14938,N_14745);
xor U15053 (N_15053,N_14003,N_14635);
xor U15054 (N_15054,N_14946,N_14147);
or U15055 (N_15055,N_14779,N_14470);
nor U15056 (N_15056,N_14720,N_14849);
xnor U15057 (N_15057,N_14509,N_14381);
nor U15058 (N_15058,N_14192,N_14414);
or U15059 (N_15059,N_14141,N_14395);
nor U15060 (N_15060,N_14190,N_14816);
and U15061 (N_15061,N_14760,N_14498);
nand U15062 (N_15062,N_14091,N_14032);
or U15063 (N_15063,N_14113,N_14926);
and U15064 (N_15064,N_14910,N_14886);
or U15065 (N_15065,N_14606,N_14984);
xnor U15066 (N_15066,N_14690,N_14687);
or U15067 (N_15067,N_14499,N_14557);
or U15068 (N_15068,N_14370,N_14618);
xnor U15069 (N_15069,N_14754,N_14818);
nand U15070 (N_15070,N_14010,N_14567);
nor U15071 (N_15071,N_14265,N_14321);
nand U15072 (N_15072,N_14800,N_14443);
xor U15073 (N_15073,N_14273,N_14652);
nand U15074 (N_15074,N_14689,N_14566);
nand U15075 (N_15075,N_14413,N_14633);
nand U15076 (N_15076,N_14442,N_14683);
xnor U15077 (N_15077,N_14009,N_14175);
xnor U15078 (N_15078,N_14547,N_14234);
and U15079 (N_15079,N_14721,N_14660);
and U15080 (N_15080,N_14485,N_14408);
or U15081 (N_15081,N_14364,N_14911);
nor U15082 (N_15082,N_14256,N_14231);
nand U15083 (N_15083,N_14008,N_14894);
xor U15084 (N_15084,N_14199,N_14957);
or U15085 (N_15085,N_14020,N_14319);
or U15086 (N_15086,N_14570,N_14170);
or U15087 (N_15087,N_14959,N_14326);
xnor U15088 (N_15088,N_14812,N_14907);
nand U15089 (N_15089,N_14786,N_14898);
and U15090 (N_15090,N_14311,N_14719);
xor U15091 (N_15091,N_14552,N_14784);
xnor U15092 (N_15092,N_14358,N_14206);
or U15093 (N_15093,N_14711,N_14612);
xnor U15094 (N_15094,N_14748,N_14309);
nand U15095 (N_15095,N_14027,N_14842);
nand U15096 (N_15096,N_14505,N_14982);
and U15097 (N_15097,N_14708,N_14921);
nand U15098 (N_15098,N_14051,N_14180);
and U15099 (N_15099,N_14675,N_14859);
nor U15100 (N_15100,N_14427,N_14415);
xnor U15101 (N_15101,N_14850,N_14148);
nor U15102 (N_15102,N_14821,N_14600);
nand U15103 (N_15103,N_14614,N_14333);
xor U15104 (N_15104,N_14876,N_14718);
nor U15105 (N_15105,N_14783,N_14220);
xor U15106 (N_15106,N_14672,N_14094);
nand U15107 (N_15107,N_14039,N_14198);
or U15108 (N_15108,N_14116,N_14359);
or U15109 (N_15109,N_14088,N_14528);
xnor U15110 (N_15110,N_14889,N_14511);
nor U15111 (N_15111,N_14815,N_14152);
xor U15112 (N_15112,N_14764,N_14794);
and U15113 (N_15113,N_14713,N_14845);
nor U15114 (N_15114,N_14024,N_14789);
nor U15115 (N_15115,N_14343,N_14223);
xor U15116 (N_15116,N_14322,N_14473);
nor U15117 (N_15117,N_14626,N_14909);
nor U15118 (N_15118,N_14704,N_14044);
and U15119 (N_15119,N_14183,N_14942);
and U15120 (N_15120,N_14331,N_14021);
xor U15121 (N_15121,N_14924,N_14578);
nand U15122 (N_15122,N_14130,N_14430);
xnor U15123 (N_15123,N_14242,N_14479);
xnor U15124 (N_15124,N_14860,N_14142);
xnor U15125 (N_15125,N_14734,N_14426);
or U15126 (N_15126,N_14362,N_14112);
xor U15127 (N_15127,N_14423,N_14390);
and U15128 (N_15128,N_14492,N_14061);
nor U15129 (N_15129,N_14194,N_14268);
nor U15130 (N_15130,N_14138,N_14820);
nand U15131 (N_15131,N_14673,N_14215);
nand U15132 (N_15132,N_14005,N_14915);
and U15133 (N_15133,N_14560,N_14438);
nand U15134 (N_15134,N_14840,N_14735);
and U15135 (N_15135,N_14512,N_14132);
or U15136 (N_15136,N_14429,N_14670);
and U15137 (N_15137,N_14646,N_14729);
and U15138 (N_15138,N_14879,N_14365);
or U15139 (N_15139,N_14939,N_14375);
nand U15140 (N_15140,N_14149,N_14136);
xnor U15141 (N_15141,N_14315,N_14213);
and U15142 (N_15142,N_14467,N_14680);
or U15143 (N_15143,N_14875,N_14863);
nand U15144 (N_15144,N_14056,N_14267);
xor U15145 (N_15145,N_14504,N_14384);
nand U15146 (N_15146,N_14593,N_14161);
xor U15147 (N_15147,N_14653,N_14761);
nand U15148 (N_15148,N_14461,N_14124);
and U15149 (N_15149,N_14550,N_14030);
or U15150 (N_15150,N_14996,N_14824);
or U15151 (N_15151,N_14545,N_14637);
nor U15152 (N_15152,N_14436,N_14145);
nand U15153 (N_15153,N_14848,N_14409);
or U15154 (N_15154,N_14595,N_14627);
nand U15155 (N_15155,N_14105,N_14613);
nand U15156 (N_15156,N_14209,N_14019);
nand U15157 (N_15157,N_14958,N_14770);
nor U15158 (N_15158,N_14174,N_14000);
nand U15159 (N_15159,N_14531,N_14001);
nand U15160 (N_15160,N_14072,N_14975);
nor U15161 (N_15161,N_14538,N_14189);
nor U15162 (N_15162,N_14520,N_14655);
and U15163 (N_15163,N_14477,N_14323);
and U15164 (N_15164,N_14118,N_14134);
xor U15165 (N_15165,N_14086,N_14247);
nand U15166 (N_15166,N_14967,N_14868);
and U15167 (N_15167,N_14211,N_14458);
xor U15168 (N_15168,N_14568,N_14313);
nand U15169 (N_15169,N_14043,N_14296);
xor U15170 (N_15170,N_14543,N_14533);
xor U15171 (N_15171,N_14345,N_14867);
xnor U15172 (N_15172,N_14597,N_14389);
xnor U15173 (N_15173,N_14649,N_14858);
nand U15174 (N_15174,N_14293,N_14986);
xnor U15175 (N_15175,N_14254,N_14440);
xnor U15176 (N_15176,N_14973,N_14767);
nor U15177 (N_15177,N_14350,N_14796);
nand U15178 (N_15178,N_14709,N_14523);
nand U15179 (N_15179,N_14640,N_14486);
xnor U15180 (N_15180,N_14941,N_14259);
xnor U15181 (N_15181,N_14607,N_14814);
nor U15182 (N_15182,N_14236,N_14237);
nand U15183 (N_15183,N_14746,N_14913);
nor U15184 (N_15184,N_14298,N_14249);
xnor U15185 (N_15185,N_14377,N_14449);
or U15186 (N_15186,N_14327,N_14255);
xor U15187 (N_15187,N_14457,N_14158);
nand U15188 (N_15188,N_14224,N_14144);
xor U15189 (N_15189,N_14897,N_14356);
nand U15190 (N_15190,N_14445,N_14835);
nand U15191 (N_15191,N_14217,N_14026);
and U15192 (N_15192,N_14896,N_14968);
and U15193 (N_15193,N_14862,N_14081);
or U15194 (N_15194,N_14608,N_14064);
nand U15195 (N_15195,N_14526,N_14195);
and U15196 (N_15196,N_14229,N_14733);
nand U15197 (N_15197,N_14063,N_14870);
xnor U15198 (N_15198,N_14830,N_14861);
and U15199 (N_15199,N_14222,N_14062);
xnor U15200 (N_15200,N_14955,N_14856);
or U15201 (N_15201,N_14453,N_14541);
xor U15202 (N_15202,N_14806,N_14448);
nand U15203 (N_15203,N_14114,N_14421);
xor U15204 (N_15204,N_14787,N_14407);
xnor U15205 (N_15205,N_14714,N_14258);
nor U15206 (N_15206,N_14609,N_14855);
or U15207 (N_15207,N_14994,N_14422);
xor U15208 (N_15208,N_14636,N_14839);
nor U15209 (N_15209,N_14083,N_14354);
xor U15210 (N_15210,N_14188,N_14451);
and U15211 (N_15211,N_14154,N_14791);
and U15212 (N_15212,N_14219,N_14585);
or U15213 (N_15213,N_14751,N_14097);
xor U15214 (N_15214,N_14750,N_14042);
nor U15215 (N_15215,N_14584,N_14330);
xor U15216 (N_15216,N_14664,N_14871);
nor U15217 (N_15217,N_14240,N_14157);
nand U15218 (N_15218,N_14306,N_14890);
xnor U15219 (N_15219,N_14774,N_14515);
xnor U15220 (N_15220,N_14065,N_14352);
and U15221 (N_15221,N_14272,N_14693);
nor U15222 (N_15222,N_14122,N_14290);
nor U15223 (N_15223,N_14998,N_14374);
or U15224 (N_15224,N_14163,N_14797);
xnor U15225 (N_15225,N_14241,N_14684);
xor U15226 (N_15226,N_14006,N_14630);
and U15227 (N_15227,N_14983,N_14762);
xor U15228 (N_15228,N_14727,N_14736);
and U15229 (N_15229,N_14759,N_14179);
nand U15230 (N_15230,N_14119,N_14233);
and U15231 (N_15231,N_14877,N_14549);
nand U15232 (N_15232,N_14444,N_14216);
xor U15233 (N_15233,N_14054,N_14823);
and U15234 (N_15234,N_14763,N_14833);
or U15235 (N_15235,N_14099,N_14253);
xnor U15236 (N_15236,N_14537,N_14715);
nor U15237 (N_15237,N_14115,N_14238);
nor U15238 (N_15238,N_14018,N_14120);
nor U15239 (N_15239,N_14454,N_14586);
xor U15240 (N_15240,N_14502,N_14874);
nand U15241 (N_15241,N_14945,N_14699);
nor U15242 (N_15242,N_14620,N_14257);
or U15243 (N_15243,N_14070,N_14286);
and U15244 (N_15244,N_14678,N_14104);
nor U15245 (N_15245,N_14469,N_14069);
and U15246 (N_15246,N_14111,N_14214);
xor U15247 (N_15247,N_14810,N_14353);
nor U15248 (N_15248,N_14262,N_14535);
xor U15249 (N_15249,N_14013,N_14022);
nor U15250 (N_15250,N_14697,N_14156);
nor U15251 (N_15251,N_14773,N_14923);
nand U15252 (N_15252,N_14698,N_14891);
or U15253 (N_15253,N_14128,N_14274);
xor U15254 (N_15254,N_14221,N_14965);
xor U15255 (N_15255,N_14948,N_14639);
nor U15256 (N_15256,N_14527,N_14819);
xnor U15257 (N_15257,N_14101,N_14831);
nand U15258 (N_15258,N_14121,N_14431);
and U15259 (N_15259,N_14371,N_14299);
and U15260 (N_15260,N_14940,N_14494);
nand U15261 (N_15261,N_14218,N_14386);
or U15262 (N_15262,N_14701,N_14361);
and U15263 (N_15263,N_14902,N_14169);
xnor U15264 (N_15264,N_14795,N_14596);
or U15265 (N_15265,N_14947,N_14881);
xnor U15266 (N_15266,N_14790,N_14651);
and U15267 (N_15267,N_14521,N_14349);
or U15268 (N_15268,N_14464,N_14250);
or U15269 (N_15269,N_14695,N_14312);
and U15270 (N_15270,N_14432,N_14963);
nand U15271 (N_15271,N_14446,N_14914);
xnor U15272 (N_15272,N_14826,N_14025);
xor U15273 (N_15273,N_14045,N_14532);
and U15274 (N_15274,N_14674,N_14602);
nand U15275 (N_15275,N_14808,N_14661);
xor U15276 (N_15276,N_14813,N_14956);
xor U15277 (N_15277,N_14320,N_14805);
xor U15278 (N_15278,N_14936,N_14015);
nor U15279 (N_15279,N_14688,N_14125);
and U15280 (N_15280,N_14228,N_14872);
and U15281 (N_15281,N_14631,N_14100);
and U15282 (N_15282,N_14029,N_14518);
xnor U15283 (N_15283,N_14793,N_14080);
xor U15284 (N_15284,N_14197,N_14851);
nor U15285 (N_15285,N_14590,N_14302);
xnor U15286 (N_15286,N_14722,N_14574);
xnor U15287 (N_15287,N_14768,N_14893);
nor U15288 (N_15288,N_14373,N_14428);
xor U15289 (N_15289,N_14577,N_14476);
nand U15290 (N_15290,N_14629,N_14934);
or U15291 (N_15291,N_14282,N_14332);
or U15292 (N_15292,N_14951,N_14329);
or U15293 (N_15293,N_14530,N_14093);
and U15294 (N_15294,N_14781,N_14730);
nand U15295 (N_15295,N_14960,N_14050);
nor U15296 (N_15296,N_14102,N_14324);
and U15297 (N_15297,N_14191,N_14992);
xor U15298 (N_15298,N_14976,N_14202);
xor U15299 (N_15299,N_14243,N_14772);
nor U15300 (N_15300,N_14304,N_14090);
nand U15301 (N_15301,N_14717,N_14227);
nor U15302 (N_15302,N_14852,N_14935);
nand U15303 (N_15303,N_14558,N_14316);
nand U15304 (N_15304,N_14677,N_14303);
or U15305 (N_15305,N_14599,N_14465);
xnor U15306 (N_15306,N_14766,N_14487);
nand U15307 (N_15307,N_14943,N_14662);
and U15308 (N_15308,N_14880,N_14514);
xor U15309 (N_15309,N_14318,N_14919);
nand U15310 (N_15310,N_14798,N_14825);
or U15311 (N_15311,N_14737,N_14917);
and U15312 (N_15312,N_14634,N_14703);
nand U15313 (N_15313,N_14011,N_14929);
xor U15314 (N_15314,N_14193,N_14073);
nand U15315 (N_15315,N_14712,N_14028);
and U15316 (N_15316,N_14185,N_14583);
or U15317 (N_15317,N_14276,N_14827);
nand U15318 (N_15318,N_14744,N_14162);
nor U15319 (N_15319,N_14164,N_14841);
nand U15320 (N_15320,N_14506,N_14650);
nor U15321 (N_15321,N_14140,N_14949);
or U15322 (N_15322,N_14559,N_14284);
nand U15323 (N_15323,N_14204,N_14696);
and U15324 (N_15324,N_14866,N_14546);
nor U15325 (N_15325,N_14776,N_14239);
xor U15326 (N_15326,N_14360,N_14419);
nand U15327 (N_15327,N_14397,N_14648);
or U15328 (N_15328,N_14103,N_14380);
nor U15329 (N_15329,N_14769,N_14420);
or U15330 (N_15330,N_14534,N_14404);
and U15331 (N_15331,N_14450,N_14058);
and U15332 (N_15332,N_14295,N_14669);
or U15333 (N_15333,N_14200,N_14723);
xor U15334 (N_15334,N_14378,N_14539);
nor U15335 (N_15335,N_14710,N_14969);
nand U15336 (N_15336,N_14916,N_14610);
nand U15337 (N_15337,N_14822,N_14905);
xnor U15338 (N_15338,N_14087,N_14060);
xor U15339 (N_15339,N_14439,N_14196);
nand U15340 (N_15340,N_14475,N_14096);
nand U15341 (N_15341,N_14366,N_14937);
nor U15342 (N_15342,N_14638,N_14681);
xnor U15343 (N_15343,N_14167,N_14287);
nand U15344 (N_15344,N_14564,N_14462);
xnor U15345 (N_15345,N_14172,N_14270);
nand U15346 (N_15346,N_14355,N_14988);
nor U15347 (N_15347,N_14592,N_14335);
nand U15348 (N_15348,N_14582,N_14587);
and U15349 (N_15349,N_14930,N_14572);
or U15350 (N_15350,N_14401,N_14981);
or U15351 (N_15351,N_14732,N_14706);
nand U15352 (N_15352,N_14139,N_14495);
nand U15353 (N_15353,N_14317,N_14883);
or U15354 (N_15354,N_14106,N_14092);
nand U15355 (N_15355,N_14676,N_14336);
nor U15356 (N_15356,N_14186,N_14887);
or U15357 (N_15357,N_14055,N_14398);
xor U15358 (N_15358,N_14110,N_14974);
and U15359 (N_15359,N_14553,N_14187);
and U15360 (N_15360,N_14788,N_14641);
or U15361 (N_15361,N_14579,N_14964);
or U15362 (N_15362,N_14244,N_14589);
xor U15363 (N_15363,N_14619,N_14344);
nand U15364 (N_15364,N_14603,N_14410);
xor U15365 (N_15365,N_14544,N_14288);
and U15366 (N_15366,N_14123,N_14962);
xnor U15367 (N_15367,N_14052,N_14888);
and U15368 (N_15368,N_14466,N_14098);
nand U15369 (N_15369,N_14645,N_14248);
nand U15370 (N_15370,N_14071,N_14529);
nand U15371 (N_15371,N_14246,N_14245);
nand U15372 (N_15372,N_14468,N_14383);
nor U15373 (N_15373,N_14904,N_14455);
xnor U15374 (N_15374,N_14382,N_14496);
and U15375 (N_15375,N_14803,N_14548);
and U15376 (N_15376,N_14508,N_14659);
and U15377 (N_15377,N_14456,N_14931);
nand U15378 (N_15378,N_14203,N_14075);
nand U15379 (N_15379,N_14725,N_14665);
nor U15380 (N_15380,N_14997,N_14666);
or U15381 (N_15381,N_14576,N_14507);
xor U15382 (N_15382,N_14656,N_14752);
or U15383 (N_15383,N_14581,N_14892);
nand U15384 (N_15384,N_14510,N_14014);
or U15385 (N_15385,N_14348,N_14536);
nor U15386 (N_15386,N_14405,N_14108);
nand U15387 (N_15387,N_14459,N_14230);
xor U15388 (N_15388,N_14847,N_14078);
and U15389 (N_15389,N_14757,N_14205);
nor U15390 (N_15390,N_14107,N_14396);
nand U15391 (N_15391,N_14041,N_14899);
xnor U15392 (N_15392,N_14503,N_14392);
and U15393 (N_15393,N_14184,N_14127);
and U15394 (N_15394,N_14077,N_14497);
and U15395 (N_15395,N_14758,N_14208);
and U15396 (N_15396,N_14150,N_14658);
nand U15397 (N_15397,N_14271,N_14301);
or U15398 (N_15398,N_14482,N_14685);
or U15399 (N_15399,N_14980,N_14857);
or U15400 (N_15400,N_14307,N_14137);
nor U15401 (N_15401,N_14035,N_14480);
and U15402 (N_15402,N_14500,N_14226);
nand U15403 (N_15403,N_14999,N_14165);
xor U15404 (N_15404,N_14782,N_14970);
or U15405 (N_15405,N_14906,N_14095);
nor U15406 (N_15406,N_14882,N_14151);
xnor U15407 (N_15407,N_14756,N_14854);
xnor U15408 (N_15408,N_14406,N_14995);
nand U15409 (N_15409,N_14489,N_14601);
xnor U15410 (N_15410,N_14160,N_14878);
xor U15411 (N_15411,N_14644,N_14181);
nand U15412 (N_15412,N_14337,N_14700);
or U15413 (N_15413,N_14394,N_14385);
or U15414 (N_15414,N_14281,N_14972);
nand U15415 (N_15415,N_14040,N_14624);
xnor U15416 (N_15416,N_14341,N_14031);
nand U15417 (N_15417,N_14369,N_14801);
nor U15418 (N_15418,N_14622,N_14168);
nor U15419 (N_15419,N_14285,N_14993);
and U15420 (N_15420,N_14264,N_14403);
nor U15421 (N_15421,N_14368,N_14067);
xnor U15422 (N_15422,N_14133,N_14339);
nand U15423 (N_15423,N_14085,N_14778);
nor U15424 (N_15424,N_14235,N_14279);
and U15425 (N_15425,N_14551,N_14351);
or U15426 (N_15426,N_14927,N_14657);
or U15427 (N_15427,N_14278,N_14979);
xor U15428 (N_15428,N_14182,N_14617);
xor U15429 (N_15429,N_14844,N_14166);
nand U15430 (N_15430,N_14089,N_14084);
nor U15431 (N_15431,N_14478,N_14901);
or U15432 (N_15432,N_14625,N_14212);
xor U15433 (N_15433,N_14292,N_14922);
xnor U15434 (N_15434,N_14047,N_14275);
and U15435 (N_15435,N_14481,N_14517);
xnor U15436 (N_15436,N_14399,N_14305);
nand U15437 (N_15437,N_14724,N_14210);
and U15438 (N_15438,N_14598,N_14280);
or U15439 (N_15439,N_14985,N_14565);
nor U15440 (N_15440,N_14561,N_14260);
nand U15441 (N_15441,N_14694,N_14605);
or U15442 (N_15442,N_14283,N_14771);
nand U15443 (N_15443,N_14802,N_14519);
and U15444 (N_15444,N_14691,N_14524);
or U15445 (N_15445,N_14679,N_14417);
or U15446 (N_15446,N_14412,N_14864);
or U15447 (N_15447,N_14785,N_14832);
nand U15448 (N_15448,N_14346,N_14068);
and U15449 (N_15449,N_14740,N_14562);
nor U15450 (N_15450,N_14082,N_14836);
nor U15451 (N_15451,N_14928,N_14347);
nor U15452 (N_15452,N_14232,N_14908);
or U15453 (N_15453,N_14525,N_14961);
nand U15454 (N_15454,N_14739,N_14702);
nand U15455 (N_15455,N_14978,N_14491);
nand U15456 (N_15456,N_14126,N_14903);
nor U15457 (N_15457,N_14493,N_14434);
or U15458 (N_15458,N_14990,N_14799);
nand U15459 (N_15459,N_14501,N_14176);
nor U15460 (N_15460,N_14143,N_14252);
or U15461 (N_15461,N_14437,N_14554);
and U15462 (N_15462,N_14291,N_14367);
xor U15463 (N_15463,N_14129,N_14340);
nand U15464 (N_15464,N_14059,N_14884);
nand U15465 (N_15465,N_14178,N_14843);
or U15466 (N_15466,N_14542,N_14402);
nor U15467 (N_15467,N_14591,N_14522);
or U15468 (N_15468,N_14573,N_14004);
or U15469 (N_15469,N_14207,N_14846);
or U15470 (N_15470,N_14173,N_14435);
nand U15471 (N_15471,N_14297,N_14668);
and U15472 (N_15472,N_14155,N_14885);
nor U15473 (N_15473,N_14310,N_14731);
nor U15474 (N_15474,N_14643,N_14263);
or U15475 (N_15475,N_14615,N_14516);
xor U15476 (N_15476,N_14556,N_14017);
or U15477 (N_15477,N_14932,N_14804);
nor U15478 (N_15478,N_14225,N_14540);
nand U15479 (N_15479,N_14780,N_14611);
nand U15480 (N_15480,N_14372,N_14388);
or U15481 (N_15481,N_14953,N_14023);
or U15482 (N_15482,N_14471,N_14834);
or U15483 (N_15483,N_14692,N_14755);
nor U15484 (N_15484,N_14765,N_14338);
or U15485 (N_15485,N_14569,N_14895);
or U15486 (N_15486,N_14294,N_14007);
and U15487 (N_15487,N_14177,N_14314);
nor U15488 (N_15488,N_14146,N_14308);
nor U15489 (N_15489,N_14807,N_14376);
and U15490 (N_15490,N_14811,N_14987);
or U15491 (N_15491,N_14002,N_14416);
nor U15492 (N_15492,N_14379,N_14201);
and U15493 (N_15493,N_14076,N_14933);
and U15494 (N_15494,N_14837,N_14716);
nand U15495 (N_15495,N_14571,N_14159);
and U15496 (N_15496,N_14342,N_14393);
nand U15497 (N_15497,N_14738,N_14472);
or U15498 (N_15498,N_14682,N_14743);
nor U15499 (N_15499,N_14036,N_14925);
nor U15500 (N_15500,N_14552,N_14220);
and U15501 (N_15501,N_14085,N_14557);
or U15502 (N_15502,N_14270,N_14645);
nand U15503 (N_15503,N_14704,N_14078);
and U15504 (N_15504,N_14662,N_14876);
or U15505 (N_15505,N_14860,N_14688);
or U15506 (N_15506,N_14687,N_14836);
or U15507 (N_15507,N_14073,N_14713);
xor U15508 (N_15508,N_14318,N_14045);
nor U15509 (N_15509,N_14734,N_14126);
and U15510 (N_15510,N_14439,N_14609);
xor U15511 (N_15511,N_14025,N_14442);
or U15512 (N_15512,N_14315,N_14973);
or U15513 (N_15513,N_14944,N_14783);
nor U15514 (N_15514,N_14130,N_14593);
xor U15515 (N_15515,N_14480,N_14905);
nor U15516 (N_15516,N_14821,N_14396);
xnor U15517 (N_15517,N_14627,N_14420);
and U15518 (N_15518,N_14318,N_14738);
xnor U15519 (N_15519,N_14420,N_14505);
nand U15520 (N_15520,N_14553,N_14411);
nand U15521 (N_15521,N_14913,N_14527);
and U15522 (N_15522,N_14903,N_14828);
or U15523 (N_15523,N_14570,N_14863);
or U15524 (N_15524,N_14283,N_14998);
or U15525 (N_15525,N_14179,N_14624);
nor U15526 (N_15526,N_14569,N_14060);
xnor U15527 (N_15527,N_14352,N_14542);
and U15528 (N_15528,N_14002,N_14934);
nand U15529 (N_15529,N_14725,N_14104);
and U15530 (N_15530,N_14950,N_14231);
nand U15531 (N_15531,N_14660,N_14291);
or U15532 (N_15532,N_14937,N_14534);
nor U15533 (N_15533,N_14142,N_14147);
nand U15534 (N_15534,N_14719,N_14483);
nand U15535 (N_15535,N_14747,N_14964);
and U15536 (N_15536,N_14786,N_14100);
and U15537 (N_15537,N_14935,N_14500);
xnor U15538 (N_15538,N_14410,N_14670);
and U15539 (N_15539,N_14160,N_14243);
and U15540 (N_15540,N_14394,N_14607);
xnor U15541 (N_15541,N_14200,N_14338);
xnor U15542 (N_15542,N_14334,N_14211);
nand U15543 (N_15543,N_14479,N_14835);
or U15544 (N_15544,N_14792,N_14946);
or U15545 (N_15545,N_14941,N_14515);
or U15546 (N_15546,N_14690,N_14620);
and U15547 (N_15547,N_14807,N_14588);
xor U15548 (N_15548,N_14125,N_14814);
xor U15549 (N_15549,N_14970,N_14203);
xor U15550 (N_15550,N_14020,N_14834);
and U15551 (N_15551,N_14901,N_14583);
nor U15552 (N_15552,N_14617,N_14162);
xor U15553 (N_15553,N_14040,N_14392);
or U15554 (N_15554,N_14752,N_14998);
xnor U15555 (N_15555,N_14331,N_14379);
xor U15556 (N_15556,N_14201,N_14866);
nor U15557 (N_15557,N_14565,N_14127);
xnor U15558 (N_15558,N_14627,N_14293);
and U15559 (N_15559,N_14319,N_14700);
nor U15560 (N_15560,N_14121,N_14808);
xnor U15561 (N_15561,N_14155,N_14751);
or U15562 (N_15562,N_14872,N_14758);
nor U15563 (N_15563,N_14505,N_14272);
xnor U15564 (N_15564,N_14605,N_14212);
or U15565 (N_15565,N_14846,N_14564);
xor U15566 (N_15566,N_14875,N_14865);
nor U15567 (N_15567,N_14537,N_14445);
or U15568 (N_15568,N_14686,N_14169);
and U15569 (N_15569,N_14825,N_14179);
and U15570 (N_15570,N_14867,N_14224);
and U15571 (N_15571,N_14165,N_14005);
nor U15572 (N_15572,N_14286,N_14176);
nand U15573 (N_15573,N_14260,N_14476);
or U15574 (N_15574,N_14357,N_14966);
or U15575 (N_15575,N_14744,N_14062);
and U15576 (N_15576,N_14779,N_14745);
nor U15577 (N_15577,N_14146,N_14545);
xnor U15578 (N_15578,N_14553,N_14603);
nor U15579 (N_15579,N_14828,N_14617);
and U15580 (N_15580,N_14344,N_14049);
nand U15581 (N_15581,N_14353,N_14424);
xor U15582 (N_15582,N_14393,N_14357);
xnor U15583 (N_15583,N_14336,N_14066);
xor U15584 (N_15584,N_14501,N_14209);
xor U15585 (N_15585,N_14560,N_14959);
nand U15586 (N_15586,N_14938,N_14791);
nand U15587 (N_15587,N_14552,N_14662);
nor U15588 (N_15588,N_14095,N_14503);
nor U15589 (N_15589,N_14018,N_14913);
and U15590 (N_15590,N_14454,N_14710);
and U15591 (N_15591,N_14610,N_14724);
nor U15592 (N_15592,N_14182,N_14845);
nand U15593 (N_15593,N_14164,N_14550);
nor U15594 (N_15594,N_14460,N_14927);
xnor U15595 (N_15595,N_14820,N_14853);
nor U15596 (N_15596,N_14127,N_14719);
xnor U15597 (N_15597,N_14431,N_14484);
or U15598 (N_15598,N_14424,N_14309);
or U15599 (N_15599,N_14377,N_14166);
nand U15600 (N_15600,N_14866,N_14902);
xor U15601 (N_15601,N_14975,N_14244);
or U15602 (N_15602,N_14874,N_14632);
or U15603 (N_15603,N_14034,N_14445);
nor U15604 (N_15604,N_14581,N_14172);
and U15605 (N_15605,N_14868,N_14290);
nor U15606 (N_15606,N_14773,N_14173);
or U15607 (N_15607,N_14049,N_14638);
or U15608 (N_15608,N_14427,N_14241);
nand U15609 (N_15609,N_14904,N_14127);
and U15610 (N_15610,N_14443,N_14356);
xnor U15611 (N_15611,N_14903,N_14240);
or U15612 (N_15612,N_14730,N_14020);
nand U15613 (N_15613,N_14984,N_14824);
nor U15614 (N_15614,N_14595,N_14824);
nor U15615 (N_15615,N_14914,N_14440);
nor U15616 (N_15616,N_14026,N_14846);
or U15617 (N_15617,N_14931,N_14520);
or U15618 (N_15618,N_14624,N_14643);
xor U15619 (N_15619,N_14659,N_14183);
or U15620 (N_15620,N_14173,N_14467);
nand U15621 (N_15621,N_14947,N_14621);
xor U15622 (N_15622,N_14189,N_14579);
nor U15623 (N_15623,N_14750,N_14709);
nor U15624 (N_15624,N_14151,N_14246);
nor U15625 (N_15625,N_14543,N_14117);
or U15626 (N_15626,N_14807,N_14141);
and U15627 (N_15627,N_14859,N_14178);
nand U15628 (N_15628,N_14877,N_14810);
xor U15629 (N_15629,N_14869,N_14359);
nand U15630 (N_15630,N_14772,N_14009);
or U15631 (N_15631,N_14365,N_14296);
nor U15632 (N_15632,N_14649,N_14842);
and U15633 (N_15633,N_14542,N_14948);
nand U15634 (N_15634,N_14565,N_14474);
xor U15635 (N_15635,N_14880,N_14011);
nor U15636 (N_15636,N_14017,N_14752);
nand U15637 (N_15637,N_14458,N_14288);
xnor U15638 (N_15638,N_14764,N_14453);
nand U15639 (N_15639,N_14545,N_14262);
or U15640 (N_15640,N_14065,N_14273);
nor U15641 (N_15641,N_14373,N_14397);
or U15642 (N_15642,N_14881,N_14581);
xor U15643 (N_15643,N_14824,N_14425);
nand U15644 (N_15644,N_14640,N_14543);
nor U15645 (N_15645,N_14769,N_14068);
xor U15646 (N_15646,N_14976,N_14320);
xnor U15647 (N_15647,N_14147,N_14916);
and U15648 (N_15648,N_14507,N_14845);
xnor U15649 (N_15649,N_14770,N_14020);
nand U15650 (N_15650,N_14319,N_14530);
and U15651 (N_15651,N_14979,N_14699);
and U15652 (N_15652,N_14793,N_14075);
nor U15653 (N_15653,N_14763,N_14481);
or U15654 (N_15654,N_14611,N_14034);
nand U15655 (N_15655,N_14216,N_14356);
xnor U15656 (N_15656,N_14080,N_14521);
nand U15657 (N_15657,N_14998,N_14648);
xnor U15658 (N_15658,N_14961,N_14347);
xor U15659 (N_15659,N_14151,N_14617);
xor U15660 (N_15660,N_14181,N_14794);
nand U15661 (N_15661,N_14897,N_14714);
xnor U15662 (N_15662,N_14305,N_14556);
xnor U15663 (N_15663,N_14312,N_14958);
or U15664 (N_15664,N_14880,N_14332);
xnor U15665 (N_15665,N_14933,N_14384);
or U15666 (N_15666,N_14976,N_14188);
nand U15667 (N_15667,N_14097,N_14855);
nand U15668 (N_15668,N_14690,N_14136);
or U15669 (N_15669,N_14668,N_14214);
nand U15670 (N_15670,N_14072,N_14096);
or U15671 (N_15671,N_14067,N_14667);
or U15672 (N_15672,N_14017,N_14142);
or U15673 (N_15673,N_14133,N_14080);
or U15674 (N_15674,N_14225,N_14439);
xnor U15675 (N_15675,N_14761,N_14779);
nor U15676 (N_15676,N_14050,N_14237);
xnor U15677 (N_15677,N_14014,N_14313);
or U15678 (N_15678,N_14521,N_14451);
nor U15679 (N_15679,N_14371,N_14263);
xnor U15680 (N_15680,N_14543,N_14307);
xor U15681 (N_15681,N_14565,N_14235);
xnor U15682 (N_15682,N_14452,N_14506);
or U15683 (N_15683,N_14131,N_14117);
and U15684 (N_15684,N_14236,N_14868);
nor U15685 (N_15685,N_14102,N_14511);
and U15686 (N_15686,N_14360,N_14212);
xnor U15687 (N_15687,N_14816,N_14157);
or U15688 (N_15688,N_14269,N_14093);
nor U15689 (N_15689,N_14904,N_14117);
or U15690 (N_15690,N_14975,N_14456);
nor U15691 (N_15691,N_14924,N_14826);
nor U15692 (N_15692,N_14667,N_14578);
nand U15693 (N_15693,N_14265,N_14304);
xnor U15694 (N_15694,N_14360,N_14920);
xnor U15695 (N_15695,N_14973,N_14551);
or U15696 (N_15696,N_14352,N_14899);
nand U15697 (N_15697,N_14257,N_14443);
and U15698 (N_15698,N_14312,N_14987);
and U15699 (N_15699,N_14042,N_14486);
nor U15700 (N_15700,N_14103,N_14234);
nor U15701 (N_15701,N_14089,N_14951);
nand U15702 (N_15702,N_14437,N_14118);
nand U15703 (N_15703,N_14225,N_14049);
and U15704 (N_15704,N_14001,N_14586);
or U15705 (N_15705,N_14996,N_14513);
nor U15706 (N_15706,N_14336,N_14027);
xnor U15707 (N_15707,N_14540,N_14647);
xor U15708 (N_15708,N_14443,N_14084);
nor U15709 (N_15709,N_14763,N_14987);
nor U15710 (N_15710,N_14763,N_14747);
and U15711 (N_15711,N_14954,N_14002);
and U15712 (N_15712,N_14468,N_14323);
and U15713 (N_15713,N_14626,N_14125);
nor U15714 (N_15714,N_14206,N_14661);
xor U15715 (N_15715,N_14051,N_14945);
nand U15716 (N_15716,N_14608,N_14591);
nand U15717 (N_15717,N_14943,N_14084);
xor U15718 (N_15718,N_14330,N_14756);
nand U15719 (N_15719,N_14403,N_14901);
or U15720 (N_15720,N_14217,N_14522);
nor U15721 (N_15721,N_14732,N_14898);
nand U15722 (N_15722,N_14358,N_14195);
nor U15723 (N_15723,N_14189,N_14094);
xor U15724 (N_15724,N_14268,N_14197);
nor U15725 (N_15725,N_14744,N_14522);
or U15726 (N_15726,N_14125,N_14182);
nor U15727 (N_15727,N_14643,N_14374);
nor U15728 (N_15728,N_14033,N_14970);
nand U15729 (N_15729,N_14510,N_14892);
nor U15730 (N_15730,N_14365,N_14122);
or U15731 (N_15731,N_14612,N_14205);
or U15732 (N_15732,N_14717,N_14530);
xnor U15733 (N_15733,N_14892,N_14585);
nand U15734 (N_15734,N_14219,N_14445);
nor U15735 (N_15735,N_14497,N_14126);
nand U15736 (N_15736,N_14102,N_14700);
nand U15737 (N_15737,N_14494,N_14720);
nor U15738 (N_15738,N_14490,N_14839);
and U15739 (N_15739,N_14409,N_14271);
xor U15740 (N_15740,N_14658,N_14895);
nand U15741 (N_15741,N_14033,N_14427);
or U15742 (N_15742,N_14146,N_14658);
or U15743 (N_15743,N_14530,N_14251);
nor U15744 (N_15744,N_14485,N_14105);
nor U15745 (N_15745,N_14539,N_14131);
nor U15746 (N_15746,N_14743,N_14827);
xor U15747 (N_15747,N_14213,N_14732);
and U15748 (N_15748,N_14079,N_14034);
nor U15749 (N_15749,N_14537,N_14629);
xor U15750 (N_15750,N_14982,N_14917);
nand U15751 (N_15751,N_14407,N_14143);
nand U15752 (N_15752,N_14867,N_14658);
nand U15753 (N_15753,N_14620,N_14054);
or U15754 (N_15754,N_14128,N_14101);
nand U15755 (N_15755,N_14593,N_14421);
nand U15756 (N_15756,N_14776,N_14573);
and U15757 (N_15757,N_14198,N_14760);
nor U15758 (N_15758,N_14193,N_14361);
nand U15759 (N_15759,N_14685,N_14887);
nand U15760 (N_15760,N_14386,N_14646);
nand U15761 (N_15761,N_14611,N_14745);
and U15762 (N_15762,N_14867,N_14833);
or U15763 (N_15763,N_14721,N_14713);
nor U15764 (N_15764,N_14628,N_14509);
xnor U15765 (N_15765,N_14510,N_14838);
nor U15766 (N_15766,N_14487,N_14330);
nor U15767 (N_15767,N_14539,N_14641);
nand U15768 (N_15768,N_14632,N_14697);
and U15769 (N_15769,N_14257,N_14896);
and U15770 (N_15770,N_14417,N_14654);
xor U15771 (N_15771,N_14937,N_14066);
or U15772 (N_15772,N_14148,N_14796);
nor U15773 (N_15773,N_14416,N_14946);
nor U15774 (N_15774,N_14241,N_14951);
xor U15775 (N_15775,N_14328,N_14768);
nor U15776 (N_15776,N_14000,N_14201);
nand U15777 (N_15777,N_14739,N_14873);
nor U15778 (N_15778,N_14148,N_14280);
and U15779 (N_15779,N_14528,N_14493);
nor U15780 (N_15780,N_14653,N_14588);
or U15781 (N_15781,N_14913,N_14837);
and U15782 (N_15782,N_14063,N_14173);
and U15783 (N_15783,N_14146,N_14870);
nor U15784 (N_15784,N_14591,N_14878);
nor U15785 (N_15785,N_14861,N_14477);
or U15786 (N_15786,N_14325,N_14632);
and U15787 (N_15787,N_14255,N_14093);
nor U15788 (N_15788,N_14769,N_14854);
nor U15789 (N_15789,N_14875,N_14947);
nor U15790 (N_15790,N_14871,N_14242);
nor U15791 (N_15791,N_14900,N_14931);
or U15792 (N_15792,N_14755,N_14189);
and U15793 (N_15793,N_14502,N_14289);
or U15794 (N_15794,N_14150,N_14885);
nand U15795 (N_15795,N_14780,N_14075);
or U15796 (N_15796,N_14553,N_14175);
nor U15797 (N_15797,N_14001,N_14785);
nand U15798 (N_15798,N_14254,N_14613);
and U15799 (N_15799,N_14771,N_14452);
and U15800 (N_15800,N_14709,N_14672);
xor U15801 (N_15801,N_14118,N_14719);
nor U15802 (N_15802,N_14019,N_14300);
nor U15803 (N_15803,N_14302,N_14374);
and U15804 (N_15804,N_14846,N_14762);
or U15805 (N_15805,N_14105,N_14592);
and U15806 (N_15806,N_14582,N_14398);
and U15807 (N_15807,N_14295,N_14119);
xor U15808 (N_15808,N_14201,N_14220);
nand U15809 (N_15809,N_14708,N_14544);
or U15810 (N_15810,N_14391,N_14388);
xnor U15811 (N_15811,N_14446,N_14889);
and U15812 (N_15812,N_14001,N_14657);
nand U15813 (N_15813,N_14318,N_14882);
and U15814 (N_15814,N_14370,N_14922);
xnor U15815 (N_15815,N_14497,N_14014);
or U15816 (N_15816,N_14640,N_14156);
nor U15817 (N_15817,N_14459,N_14104);
or U15818 (N_15818,N_14536,N_14116);
nand U15819 (N_15819,N_14427,N_14317);
nor U15820 (N_15820,N_14994,N_14219);
xor U15821 (N_15821,N_14679,N_14806);
nor U15822 (N_15822,N_14488,N_14482);
nor U15823 (N_15823,N_14174,N_14223);
nand U15824 (N_15824,N_14253,N_14396);
nor U15825 (N_15825,N_14295,N_14118);
or U15826 (N_15826,N_14033,N_14000);
nand U15827 (N_15827,N_14543,N_14360);
nor U15828 (N_15828,N_14277,N_14982);
nor U15829 (N_15829,N_14281,N_14951);
nor U15830 (N_15830,N_14845,N_14552);
or U15831 (N_15831,N_14413,N_14537);
nand U15832 (N_15832,N_14372,N_14926);
nor U15833 (N_15833,N_14643,N_14503);
xor U15834 (N_15834,N_14429,N_14400);
nand U15835 (N_15835,N_14531,N_14955);
xnor U15836 (N_15836,N_14827,N_14712);
and U15837 (N_15837,N_14672,N_14902);
xnor U15838 (N_15838,N_14426,N_14065);
nand U15839 (N_15839,N_14123,N_14904);
or U15840 (N_15840,N_14584,N_14128);
and U15841 (N_15841,N_14129,N_14100);
and U15842 (N_15842,N_14420,N_14839);
nor U15843 (N_15843,N_14483,N_14729);
and U15844 (N_15844,N_14772,N_14625);
or U15845 (N_15845,N_14945,N_14329);
and U15846 (N_15846,N_14057,N_14442);
and U15847 (N_15847,N_14169,N_14680);
and U15848 (N_15848,N_14472,N_14573);
and U15849 (N_15849,N_14670,N_14734);
and U15850 (N_15850,N_14902,N_14319);
or U15851 (N_15851,N_14071,N_14595);
or U15852 (N_15852,N_14637,N_14019);
or U15853 (N_15853,N_14093,N_14515);
or U15854 (N_15854,N_14769,N_14198);
nor U15855 (N_15855,N_14458,N_14480);
xnor U15856 (N_15856,N_14730,N_14852);
xnor U15857 (N_15857,N_14774,N_14072);
nor U15858 (N_15858,N_14735,N_14921);
nand U15859 (N_15859,N_14238,N_14908);
and U15860 (N_15860,N_14936,N_14786);
xor U15861 (N_15861,N_14742,N_14702);
xor U15862 (N_15862,N_14400,N_14624);
or U15863 (N_15863,N_14500,N_14964);
or U15864 (N_15864,N_14287,N_14759);
nor U15865 (N_15865,N_14913,N_14567);
nor U15866 (N_15866,N_14698,N_14479);
and U15867 (N_15867,N_14211,N_14196);
nand U15868 (N_15868,N_14012,N_14092);
nand U15869 (N_15869,N_14537,N_14615);
xnor U15870 (N_15870,N_14591,N_14447);
nor U15871 (N_15871,N_14292,N_14195);
or U15872 (N_15872,N_14112,N_14009);
nor U15873 (N_15873,N_14441,N_14850);
xnor U15874 (N_15874,N_14862,N_14972);
nor U15875 (N_15875,N_14505,N_14388);
and U15876 (N_15876,N_14276,N_14332);
xnor U15877 (N_15877,N_14150,N_14450);
nand U15878 (N_15878,N_14623,N_14709);
nand U15879 (N_15879,N_14209,N_14184);
nor U15880 (N_15880,N_14479,N_14467);
nor U15881 (N_15881,N_14632,N_14292);
nand U15882 (N_15882,N_14487,N_14705);
xnor U15883 (N_15883,N_14052,N_14991);
nand U15884 (N_15884,N_14587,N_14183);
xor U15885 (N_15885,N_14267,N_14276);
and U15886 (N_15886,N_14473,N_14634);
xor U15887 (N_15887,N_14183,N_14422);
and U15888 (N_15888,N_14323,N_14811);
xnor U15889 (N_15889,N_14850,N_14668);
and U15890 (N_15890,N_14824,N_14758);
nor U15891 (N_15891,N_14165,N_14194);
or U15892 (N_15892,N_14837,N_14068);
nor U15893 (N_15893,N_14959,N_14212);
and U15894 (N_15894,N_14367,N_14679);
xnor U15895 (N_15895,N_14424,N_14701);
and U15896 (N_15896,N_14667,N_14537);
nand U15897 (N_15897,N_14503,N_14617);
xnor U15898 (N_15898,N_14232,N_14336);
nand U15899 (N_15899,N_14776,N_14334);
nand U15900 (N_15900,N_14971,N_14956);
and U15901 (N_15901,N_14542,N_14342);
xnor U15902 (N_15902,N_14057,N_14053);
nand U15903 (N_15903,N_14776,N_14887);
or U15904 (N_15904,N_14319,N_14006);
and U15905 (N_15905,N_14843,N_14816);
nand U15906 (N_15906,N_14982,N_14478);
nand U15907 (N_15907,N_14271,N_14071);
or U15908 (N_15908,N_14344,N_14976);
nand U15909 (N_15909,N_14826,N_14591);
nand U15910 (N_15910,N_14134,N_14852);
nor U15911 (N_15911,N_14094,N_14891);
xor U15912 (N_15912,N_14691,N_14959);
nor U15913 (N_15913,N_14385,N_14067);
or U15914 (N_15914,N_14462,N_14891);
nand U15915 (N_15915,N_14787,N_14710);
xnor U15916 (N_15916,N_14524,N_14613);
nand U15917 (N_15917,N_14596,N_14890);
nor U15918 (N_15918,N_14335,N_14049);
nand U15919 (N_15919,N_14444,N_14312);
and U15920 (N_15920,N_14199,N_14598);
nand U15921 (N_15921,N_14318,N_14877);
and U15922 (N_15922,N_14562,N_14297);
xor U15923 (N_15923,N_14922,N_14642);
xnor U15924 (N_15924,N_14446,N_14581);
nand U15925 (N_15925,N_14287,N_14922);
and U15926 (N_15926,N_14468,N_14969);
nor U15927 (N_15927,N_14321,N_14627);
nor U15928 (N_15928,N_14255,N_14787);
xnor U15929 (N_15929,N_14212,N_14966);
nand U15930 (N_15930,N_14451,N_14969);
or U15931 (N_15931,N_14692,N_14222);
xnor U15932 (N_15932,N_14037,N_14736);
nand U15933 (N_15933,N_14000,N_14907);
nor U15934 (N_15934,N_14583,N_14146);
and U15935 (N_15935,N_14478,N_14824);
and U15936 (N_15936,N_14620,N_14267);
and U15937 (N_15937,N_14664,N_14486);
or U15938 (N_15938,N_14507,N_14108);
xnor U15939 (N_15939,N_14743,N_14716);
xnor U15940 (N_15940,N_14747,N_14281);
or U15941 (N_15941,N_14246,N_14338);
nor U15942 (N_15942,N_14811,N_14598);
xor U15943 (N_15943,N_14217,N_14617);
nor U15944 (N_15944,N_14953,N_14995);
nand U15945 (N_15945,N_14815,N_14578);
nor U15946 (N_15946,N_14054,N_14393);
or U15947 (N_15947,N_14670,N_14287);
nand U15948 (N_15948,N_14456,N_14637);
and U15949 (N_15949,N_14631,N_14817);
xor U15950 (N_15950,N_14594,N_14335);
xor U15951 (N_15951,N_14879,N_14651);
and U15952 (N_15952,N_14116,N_14897);
or U15953 (N_15953,N_14922,N_14570);
and U15954 (N_15954,N_14134,N_14835);
nor U15955 (N_15955,N_14868,N_14323);
nand U15956 (N_15956,N_14559,N_14102);
nand U15957 (N_15957,N_14410,N_14862);
or U15958 (N_15958,N_14858,N_14668);
or U15959 (N_15959,N_14781,N_14670);
and U15960 (N_15960,N_14570,N_14055);
xor U15961 (N_15961,N_14458,N_14902);
or U15962 (N_15962,N_14427,N_14904);
nand U15963 (N_15963,N_14815,N_14456);
or U15964 (N_15964,N_14204,N_14551);
and U15965 (N_15965,N_14453,N_14357);
nor U15966 (N_15966,N_14963,N_14353);
or U15967 (N_15967,N_14104,N_14573);
and U15968 (N_15968,N_14636,N_14794);
or U15969 (N_15969,N_14468,N_14194);
nor U15970 (N_15970,N_14833,N_14799);
or U15971 (N_15971,N_14769,N_14426);
or U15972 (N_15972,N_14488,N_14862);
and U15973 (N_15973,N_14847,N_14860);
or U15974 (N_15974,N_14604,N_14387);
xor U15975 (N_15975,N_14154,N_14410);
nor U15976 (N_15976,N_14009,N_14767);
or U15977 (N_15977,N_14095,N_14978);
or U15978 (N_15978,N_14567,N_14544);
xor U15979 (N_15979,N_14584,N_14277);
and U15980 (N_15980,N_14807,N_14026);
nor U15981 (N_15981,N_14476,N_14129);
nor U15982 (N_15982,N_14662,N_14534);
nor U15983 (N_15983,N_14866,N_14527);
xor U15984 (N_15984,N_14192,N_14962);
or U15985 (N_15985,N_14733,N_14643);
or U15986 (N_15986,N_14328,N_14257);
nand U15987 (N_15987,N_14812,N_14716);
or U15988 (N_15988,N_14486,N_14593);
and U15989 (N_15989,N_14435,N_14381);
or U15990 (N_15990,N_14439,N_14315);
nor U15991 (N_15991,N_14985,N_14607);
nor U15992 (N_15992,N_14969,N_14773);
nand U15993 (N_15993,N_14307,N_14969);
or U15994 (N_15994,N_14689,N_14488);
nand U15995 (N_15995,N_14719,N_14534);
and U15996 (N_15996,N_14860,N_14261);
nor U15997 (N_15997,N_14305,N_14488);
nor U15998 (N_15998,N_14945,N_14312);
nor U15999 (N_15999,N_14894,N_14820);
xnor U16000 (N_16000,N_15177,N_15259);
or U16001 (N_16001,N_15161,N_15239);
and U16002 (N_16002,N_15783,N_15215);
nor U16003 (N_16003,N_15713,N_15701);
or U16004 (N_16004,N_15753,N_15875);
nand U16005 (N_16005,N_15399,N_15101);
xnor U16006 (N_16006,N_15078,N_15842);
xor U16007 (N_16007,N_15360,N_15932);
nand U16008 (N_16008,N_15722,N_15036);
xor U16009 (N_16009,N_15396,N_15838);
nor U16010 (N_16010,N_15376,N_15410);
or U16011 (N_16011,N_15047,N_15939);
xor U16012 (N_16012,N_15976,N_15618);
or U16013 (N_16013,N_15346,N_15216);
nor U16014 (N_16014,N_15121,N_15823);
and U16015 (N_16015,N_15180,N_15416);
nand U16016 (N_16016,N_15240,N_15365);
nor U16017 (N_16017,N_15420,N_15579);
nor U16018 (N_16018,N_15706,N_15107);
and U16019 (N_16019,N_15651,N_15633);
nor U16020 (N_16020,N_15985,N_15150);
or U16021 (N_16021,N_15717,N_15250);
or U16022 (N_16022,N_15805,N_15544);
or U16023 (N_16023,N_15917,N_15265);
nand U16024 (N_16024,N_15637,N_15244);
or U16025 (N_16025,N_15248,N_15507);
nand U16026 (N_16026,N_15820,N_15666);
xor U16027 (N_16027,N_15219,N_15948);
or U16028 (N_16028,N_15252,N_15667);
or U16029 (N_16029,N_15311,N_15147);
or U16030 (N_16030,N_15950,N_15208);
and U16031 (N_16031,N_15214,N_15891);
nand U16032 (N_16032,N_15258,N_15608);
and U16033 (N_16033,N_15980,N_15961);
or U16034 (N_16034,N_15334,N_15692);
and U16035 (N_16035,N_15482,N_15058);
and U16036 (N_16036,N_15890,N_15880);
and U16037 (N_16037,N_15297,N_15750);
or U16038 (N_16038,N_15262,N_15131);
or U16039 (N_16039,N_15357,N_15638);
xor U16040 (N_16040,N_15430,N_15644);
and U16041 (N_16041,N_15495,N_15963);
nor U16042 (N_16042,N_15818,N_15893);
or U16043 (N_16043,N_15515,N_15234);
or U16044 (N_16044,N_15417,N_15743);
xnor U16045 (N_16045,N_15740,N_15777);
nor U16046 (N_16046,N_15347,N_15140);
and U16047 (N_16047,N_15075,N_15746);
nor U16048 (N_16048,N_15151,N_15433);
and U16049 (N_16049,N_15729,N_15862);
nand U16050 (N_16050,N_15469,N_15968);
and U16051 (N_16051,N_15703,N_15737);
nand U16052 (N_16052,N_15098,N_15723);
xor U16053 (N_16053,N_15388,N_15478);
xor U16054 (N_16054,N_15028,N_15756);
or U16055 (N_16055,N_15764,N_15871);
and U16056 (N_16056,N_15866,N_15460);
xor U16057 (N_16057,N_15125,N_15174);
xnor U16058 (N_16058,N_15711,N_15268);
nand U16059 (N_16059,N_15906,N_15336);
and U16060 (N_16060,N_15189,N_15872);
or U16061 (N_16061,N_15129,N_15484);
or U16062 (N_16062,N_15829,N_15959);
nand U16063 (N_16063,N_15074,N_15690);
nand U16064 (N_16064,N_15069,N_15669);
and U16065 (N_16065,N_15439,N_15839);
or U16066 (N_16066,N_15795,N_15953);
nand U16067 (N_16067,N_15598,N_15739);
xnor U16068 (N_16068,N_15732,N_15518);
or U16069 (N_16069,N_15779,N_15468);
xor U16070 (N_16070,N_15951,N_15942);
nand U16071 (N_16071,N_15883,N_15264);
or U16072 (N_16072,N_15015,N_15626);
and U16073 (N_16073,N_15628,N_15869);
and U16074 (N_16074,N_15558,N_15878);
nor U16075 (N_16075,N_15397,N_15176);
or U16076 (N_16076,N_15513,N_15170);
nand U16077 (N_16077,N_15619,N_15896);
or U16078 (N_16078,N_15909,N_15904);
xor U16079 (N_16079,N_15441,N_15418);
xnor U16080 (N_16080,N_15974,N_15242);
nor U16081 (N_16081,N_15575,N_15494);
xor U16082 (N_16082,N_15096,N_15424);
or U16083 (N_16083,N_15286,N_15162);
nand U16084 (N_16084,N_15745,N_15782);
xor U16085 (N_16085,N_15367,N_15362);
nor U16086 (N_16086,N_15926,N_15724);
xnor U16087 (N_16087,N_15304,N_15063);
nor U16088 (N_16088,N_15230,N_15382);
and U16089 (N_16089,N_15033,N_15762);
nand U16090 (N_16090,N_15555,N_15971);
nand U16091 (N_16091,N_15960,N_15733);
xnor U16092 (N_16092,N_15895,N_15500);
or U16093 (N_16093,N_15962,N_15812);
and U16094 (N_16094,N_15719,N_15175);
and U16095 (N_16095,N_15414,N_15492);
nand U16096 (N_16096,N_15340,N_15901);
or U16097 (N_16097,N_15664,N_15663);
or U16098 (N_16098,N_15094,N_15255);
nand U16099 (N_16099,N_15543,N_15999);
nor U16100 (N_16100,N_15765,N_15315);
or U16101 (N_16101,N_15952,N_15919);
nand U16102 (N_16102,N_15137,N_15594);
or U16103 (N_16103,N_15372,N_15538);
nand U16104 (N_16104,N_15899,N_15532);
nor U16105 (N_16105,N_15828,N_15580);
xnor U16106 (N_16106,N_15530,N_15688);
nand U16107 (N_16107,N_15696,N_15653);
nor U16108 (N_16108,N_15755,N_15674);
nand U16109 (N_16109,N_15200,N_15834);
nor U16110 (N_16110,N_15203,N_15730);
or U16111 (N_16111,N_15165,N_15973);
or U16112 (N_16112,N_15757,N_15395);
nand U16113 (N_16113,N_15389,N_15726);
nor U16114 (N_16114,N_15727,N_15853);
nor U16115 (N_16115,N_15569,N_15025);
xnor U16116 (N_16116,N_15991,N_15790);
and U16117 (N_16117,N_15712,N_15012);
and U16118 (N_16118,N_15049,N_15659);
nand U16119 (N_16119,N_15027,N_15865);
and U16120 (N_16120,N_15997,N_15648);
or U16121 (N_16121,N_15381,N_15789);
xor U16122 (N_16122,N_15572,N_15198);
xnor U16123 (N_16123,N_15285,N_15288);
nor U16124 (N_16124,N_15550,N_15741);
nand U16125 (N_16125,N_15132,N_15990);
xor U16126 (N_16126,N_15934,N_15053);
or U16127 (N_16127,N_15052,N_15531);
nor U16128 (N_16128,N_15989,N_15526);
xor U16129 (N_16129,N_15308,N_15220);
and U16130 (N_16130,N_15610,N_15167);
or U16131 (N_16131,N_15432,N_15683);
nand U16132 (N_16132,N_15704,N_15832);
xor U16133 (N_16133,N_15656,N_15799);
nor U16134 (N_16134,N_15816,N_15383);
nand U16135 (N_16135,N_15089,N_15253);
and U16136 (N_16136,N_15977,N_15614);
or U16137 (N_16137,N_15002,N_15302);
or U16138 (N_16138,N_15301,N_15427);
xnor U16139 (N_16139,N_15671,N_15256);
or U16140 (N_16140,N_15481,N_15356);
xor U16141 (N_16141,N_15864,N_15747);
nor U16142 (N_16142,N_15322,N_15710);
nand U16143 (N_16143,N_15924,N_15655);
and U16144 (N_16144,N_15126,N_15954);
nand U16145 (N_16145,N_15207,N_15474);
xor U16146 (N_16146,N_15604,N_15130);
xor U16147 (N_16147,N_15409,N_15339);
xor U16148 (N_16148,N_15884,N_15448);
nand U16149 (N_16149,N_15708,N_15331);
or U16150 (N_16150,N_15624,N_15806);
nand U16151 (N_16151,N_15918,N_15401);
and U16152 (N_16152,N_15994,N_15639);
nand U16153 (N_16153,N_15627,N_15344);
xor U16154 (N_16154,N_15605,N_15235);
nor U16155 (N_16155,N_15986,N_15509);
nand U16156 (N_16156,N_15278,N_15348);
nor U16157 (N_16157,N_15521,N_15773);
nor U16158 (N_16158,N_15095,N_15467);
or U16159 (N_16159,N_15752,N_15541);
or U16160 (N_16160,N_15428,N_15254);
xnor U16161 (N_16161,N_15592,N_15693);
nand U16162 (N_16162,N_15326,N_15090);
xor U16163 (N_16163,N_15060,N_15759);
and U16164 (N_16164,N_15613,N_15342);
nand U16165 (N_16165,N_15451,N_15312);
and U16166 (N_16166,N_15158,N_15066);
or U16167 (N_16167,N_15112,N_15384);
nand U16168 (N_16168,N_15965,N_15586);
and U16169 (N_16169,N_15228,N_15291);
nor U16170 (N_16170,N_15597,N_15070);
nor U16171 (N_16171,N_15545,N_15825);
xnor U16172 (N_16172,N_15008,N_15535);
or U16173 (N_16173,N_15949,N_15907);
nand U16174 (N_16174,N_15758,N_15398);
and U16175 (N_16175,N_15041,N_15363);
xor U16176 (N_16176,N_15364,N_15303);
and U16177 (N_16177,N_15574,N_15108);
nand U16178 (N_16178,N_15387,N_15246);
nand U16179 (N_16179,N_15355,N_15860);
or U16180 (N_16180,N_15958,N_15009);
nand U16181 (N_16181,N_15645,N_15776);
nand U16182 (N_16182,N_15067,N_15615);
nor U16183 (N_16183,N_15846,N_15984);
nand U16184 (N_16184,N_15547,N_15566);
nand U16185 (N_16185,N_15910,N_15183);
and U16186 (N_16186,N_15477,N_15082);
nand U16187 (N_16187,N_15836,N_15625);
nor U16188 (N_16188,N_15488,N_15928);
xor U16189 (N_16189,N_15442,N_15793);
and U16190 (N_16190,N_15888,N_15109);
nor U16191 (N_16191,N_15874,N_15245);
nand U16192 (N_16192,N_15857,N_15307);
and U16193 (N_16193,N_15276,N_15916);
or U16194 (N_16194,N_15001,N_15211);
and U16195 (N_16195,N_15735,N_15280);
xor U16196 (N_16196,N_15300,N_15557);
and U16197 (N_16197,N_15007,N_15612);
nor U16198 (N_16198,N_15826,N_15379);
or U16199 (N_16199,N_15110,N_15475);
or U16200 (N_16200,N_15970,N_15635);
nor U16201 (N_16201,N_15804,N_15819);
and U16202 (N_16202,N_15423,N_15328);
or U16203 (N_16203,N_15128,N_15943);
xnor U16204 (N_16204,N_15707,N_15032);
or U16205 (N_16205,N_15603,N_15833);
or U16206 (N_16206,N_15296,N_15159);
nor U16207 (N_16207,N_15282,N_15714);
or U16208 (N_16208,N_15643,N_15071);
and U16209 (N_16209,N_15144,N_15927);
nand U16210 (N_16210,N_15957,N_15016);
xnor U16211 (N_16211,N_15751,N_15879);
and U16212 (N_16212,N_15263,N_15503);
nor U16213 (N_16213,N_15378,N_15673);
or U16214 (N_16214,N_15892,N_15944);
nand U16215 (N_16215,N_15172,N_15425);
nand U16216 (N_16216,N_15261,N_15780);
nor U16217 (N_16217,N_15192,N_15419);
nor U16218 (N_16218,N_15975,N_15084);
or U16219 (N_16219,N_15293,N_15882);
nand U16220 (N_16220,N_15650,N_15470);
nor U16221 (N_16221,N_15632,N_15124);
nor U16222 (N_16222,N_15292,N_15652);
xnor U16223 (N_16223,N_15502,N_15116);
and U16224 (N_16224,N_15807,N_15894);
and U16225 (N_16225,N_15523,N_15148);
or U16226 (N_16226,N_15237,N_15914);
and U16227 (N_16227,N_15657,N_15721);
xor U16228 (N_16228,N_15562,N_15654);
or U16229 (N_16229,N_15559,N_15560);
or U16230 (N_16230,N_15221,N_15299);
nand U16231 (N_16231,N_15289,N_15677);
or U16232 (N_16232,N_15204,N_15305);
xor U16233 (N_16233,N_15354,N_15668);
nor U16234 (N_16234,N_15851,N_15811);
nor U16235 (N_16235,N_15157,N_15168);
and U16236 (N_16236,N_15861,N_15178);
nand U16237 (N_16237,N_15599,N_15913);
xor U16238 (N_16238,N_15528,N_15377);
nand U16239 (N_16239,N_15270,N_15284);
xor U16240 (N_16240,N_15452,N_15319);
xor U16241 (N_16241,N_15877,N_15374);
xnor U16242 (N_16242,N_15930,N_15415);
nor U16243 (N_16243,N_15003,N_15802);
nand U16244 (N_16244,N_15349,N_15794);
nand U16245 (N_16245,N_15317,N_15578);
xor U16246 (N_16246,N_15887,N_15809);
nor U16247 (N_16247,N_15798,N_15695);
nand U16248 (N_16248,N_15487,N_15051);
and U16249 (N_16249,N_15800,N_15154);
or U16250 (N_16250,N_15184,N_15595);
and U16251 (N_16251,N_15744,N_15358);
and U16252 (N_16252,N_15630,N_15103);
nand U16253 (N_16253,N_15337,N_15533);
nor U16254 (N_16254,N_15444,N_15283);
nand U16255 (N_16255,N_15456,N_15602);
nand U16256 (N_16256,N_15830,N_15831);
nor U16257 (N_16257,N_15437,N_15539);
or U16258 (N_16258,N_15623,N_15725);
nand U16259 (N_16259,N_15679,N_15769);
nor U16260 (N_16260,N_15403,N_15083);
nor U16261 (N_16261,N_15329,N_15325);
nor U16262 (N_16262,N_15563,N_15738);
nand U16263 (N_16263,N_15803,N_15929);
or U16264 (N_16264,N_15353,N_15048);
and U16265 (N_16265,N_15956,N_15967);
or U16266 (N_16266,N_15141,N_15113);
nand U16267 (N_16267,N_15194,N_15102);
nor U16268 (N_16268,N_15576,N_15549);
nor U16269 (N_16269,N_15808,N_15405);
nand U16270 (N_16270,N_15005,N_15848);
and U16271 (N_16271,N_15590,N_15086);
nor U16272 (N_16272,N_15689,N_15672);
nand U16273 (N_16273,N_15698,N_15318);
nor U16274 (N_16274,N_15691,N_15591);
nand U16275 (N_16275,N_15734,N_15969);
and U16276 (N_16276,N_15497,N_15870);
nand U16277 (N_16277,N_15472,N_15647);
nor U16278 (N_16278,N_15642,N_15222);
and U16279 (N_16279,N_15197,N_15553);
nand U16280 (N_16280,N_15685,N_15135);
nor U16281 (N_16281,N_15641,N_15760);
xor U16282 (N_16282,N_15837,N_15678);
nor U16283 (N_16283,N_15323,N_15038);
xor U16284 (N_16284,N_15120,N_15266);
nand U16285 (N_16285,N_15506,N_15546);
and U16286 (N_16286,N_15134,N_15840);
xnor U16287 (N_16287,N_15881,N_15013);
or U16288 (N_16288,N_15537,N_15435);
nand U16289 (N_16289,N_15915,N_15885);
nor U16290 (N_16290,N_15249,N_15993);
xnor U16291 (N_16291,N_15859,N_15709);
nor U16292 (N_16292,N_15105,N_15778);
and U16293 (N_16293,N_15675,N_15496);
nor U16294 (N_16294,N_15143,N_15490);
nor U16295 (N_16295,N_15443,N_15680);
nand U16296 (N_16296,N_15863,N_15385);
nand U16297 (N_16297,N_15202,N_15400);
and U16298 (N_16298,N_15436,N_15115);
nor U16299 (N_16299,N_15164,N_15493);
or U16300 (N_16300,N_15171,N_15404);
or U16301 (N_16301,N_15844,N_15988);
and U16302 (N_16302,N_15294,N_15201);
nor U16303 (N_16303,N_15375,N_15438);
xor U16304 (N_16304,N_15408,N_15786);
or U16305 (N_16305,N_15462,N_15466);
nor U16306 (N_16306,N_15324,N_15852);
or U16307 (N_16307,N_15897,N_15440);
or U16308 (N_16308,N_15920,N_15123);
nand U16309 (N_16309,N_15585,N_15351);
and U16310 (N_16310,N_15054,N_15873);
nor U16311 (N_16311,N_15921,N_15023);
and U16312 (N_16312,N_15022,N_15552);
and U16313 (N_16313,N_15111,N_15941);
nand U16314 (N_16314,N_15145,N_15055);
and U16315 (N_16315,N_15163,N_15290);
nor U16316 (N_16316,N_15338,N_15224);
or U16317 (N_16317,N_15434,N_15978);
or U16318 (N_16318,N_15277,N_15429);
nand U16319 (N_16319,N_15565,N_15785);
or U16320 (N_16320,N_15185,N_15227);
xnor U16321 (N_16321,N_15868,N_15607);
or U16322 (N_16322,N_15855,N_15856);
nor U16323 (N_16323,N_15583,N_15996);
or U16324 (N_16324,N_15295,N_15391);
and U16325 (N_16325,N_15935,N_15225);
or U16326 (N_16326,N_15411,N_15188);
nand U16327 (N_16327,N_15987,N_15251);
nand U16328 (N_16328,N_15529,N_15345);
nor U16329 (N_16329,N_15571,N_15511);
nor U16330 (N_16330,N_15454,N_15026);
nor U16331 (N_16331,N_15209,N_15945);
nor U16332 (N_16332,N_15274,N_15596);
and U16333 (N_16333,N_15369,N_15749);
nand U16334 (N_16334,N_15155,N_15681);
xor U16335 (N_16335,N_15039,N_15402);
and U16336 (N_16336,N_15841,N_15771);
nand U16337 (N_16337,N_15754,N_15191);
nor U16338 (N_16338,N_15138,N_15056);
or U16339 (N_16339,N_15099,N_15298);
nor U16340 (N_16340,N_15587,N_15964);
and U16341 (N_16341,N_15350,N_15589);
and U16342 (N_16342,N_15824,N_15046);
xor U16343 (N_16343,N_15577,N_15313);
nand U16344 (N_16344,N_15104,N_15684);
nand U16345 (N_16345,N_15534,N_15370);
nand U16346 (N_16346,N_15457,N_15361);
nor U16347 (N_16347,N_15480,N_15660);
and U16348 (N_16348,N_15330,N_15767);
nor U16349 (N_16349,N_15728,N_15498);
xor U16350 (N_16350,N_15699,N_15979);
nand U16351 (N_16351,N_15584,N_15169);
nand U16352 (N_16352,N_15621,N_15634);
and U16353 (N_16353,N_15426,N_15849);
and U16354 (N_16354,N_15160,N_15933);
nor U16355 (N_16355,N_15079,N_15519);
or U16356 (N_16356,N_15582,N_15761);
and U16357 (N_16357,N_15796,N_15814);
nand U16358 (N_16358,N_15241,N_15702);
xor U16359 (N_16359,N_15004,N_15213);
nand U16360 (N_16360,N_15911,N_15446);
and U16361 (N_16361,N_15564,N_15271);
and U16362 (N_16362,N_15995,N_15062);
nand U16363 (N_16363,N_15542,N_15073);
and U16364 (N_16364,N_15035,N_15600);
and U16365 (N_16365,N_15076,N_15784);
nand U16366 (N_16366,N_15077,N_15114);
nand U16367 (N_16367,N_15686,N_15620);
xor U16368 (N_16368,N_15661,N_15269);
or U16369 (N_16369,N_15031,N_15489);
and U16370 (N_16370,N_15445,N_15146);
and U16371 (N_16371,N_15858,N_15018);
or U16372 (N_16372,N_15606,N_15327);
nand U16373 (N_16373,N_15097,N_15670);
and U16374 (N_16374,N_15206,N_15514);
xor U16375 (N_16375,N_15333,N_15763);
nand U16376 (N_16376,N_15827,N_15359);
or U16377 (N_16377,N_15059,N_15536);
and U16378 (N_16378,N_15854,N_15231);
nand U16379 (N_16379,N_15540,N_15946);
and U16380 (N_16380,N_15193,N_15631);
nand U16381 (N_16381,N_15187,N_15229);
nor U16382 (N_16382,N_15050,N_15649);
and U16383 (N_16383,N_15570,N_15092);
or U16384 (N_16384,N_15766,N_15152);
nor U16385 (N_16385,N_15486,N_15517);
nand U16386 (N_16386,N_15413,N_15061);
or U16387 (N_16387,N_15064,N_15368);
or U16388 (N_16388,N_15119,N_15551);
and U16389 (N_16389,N_15473,N_15394);
nor U16390 (N_16390,N_15835,N_15320);
or U16391 (N_16391,N_15556,N_15453);
and U16392 (N_16392,N_15516,N_15081);
nor U16393 (N_16393,N_15636,N_15588);
xnor U16394 (N_16394,N_15772,N_15925);
nand U16395 (N_16395,N_15019,N_15226);
xnor U16396 (N_16396,N_15199,N_15499);
nand U16397 (N_16397,N_15392,N_15922);
and U16398 (N_16398,N_15257,N_15190);
or U16399 (N_16399,N_15731,N_15561);
and U16400 (N_16400,N_15260,N_15306);
xnor U16401 (N_16401,N_15898,N_15867);
or U16402 (N_16402,N_15815,N_15715);
xor U16403 (N_16403,N_15273,N_15705);
nand U16404 (N_16404,N_15886,N_15373);
or U16405 (N_16405,N_15568,N_15581);
and U16406 (N_16406,N_15281,N_15718);
xor U16407 (N_16407,N_15279,N_15014);
or U16408 (N_16408,N_15173,N_15010);
and U16409 (N_16409,N_15020,N_15658);
and U16410 (N_16410,N_15622,N_15223);
xor U16411 (N_16411,N_15133,N_15156);
nand U16412 (N_16412,N_15593,N_15821);
nand U16413 (N_16413,N_15458,N_15087);
or U16414 (N_16414,N_15459,N_15091);
or U16415 (N_16415,N_15461,N_15341);
or U16416 (N_16416,N_15501,N_15700);
nand U16417 (N_16417,N_15966,N_15029);
and U16418 (N_16418,N_15510,N_15938);
nand U16419 (N_16419,N_15843,N_15983);
and U16420 (N_16420,N_15393,N_15900);
nor U16421 (N_16421,N_15352,N_15998);
xnor U16422 (N_16422,N_15195,N_15981);
nand U16423 (N_16423,N_15768,N_15037);
nand U16424 (N_16424,N_15781,N_15716);
or U16425 (N_16425,N_15455,N_15217);
or U16426 (N_16426,N_15287,N_15687);
xor U16427 (N_16427,N_15972,N_15524);
nor U16428 (N_16428,N_15876,N_15243);
nand U16429 (N_16429,N_15100,N_15006);
nand U16430 (N_16430,N_15748,N_15694);
or U16431 (N_16431,N_15321,N_15640);
xor U16432 (N_16432,N_15117,N_15088);
or U16433 (N_16433,N_15889,N_15770);
nor U16434 (N_16434,N_15788,N_15646);
nor U16435 (N_16435,N_15908,N_15153);
or U16436 (N_16436,N_15464,N_15218);
nand U16437 (N_16437,N_15937,N_15068);
nor U16438 (N_16438,N_15813,N_15450);
xor U16439 (N_16439,N_15386,N_15817);
and U16440 (N_16440,N_15040,N_15181);
and U16441 (N_16441,N_15527,N_15139);
or U16442 (N_16442,N_15629,N_15850);
or U16443 (N_16443,N_15801,N_15476);
xor U16444 (N_16444,N_15810,N_15316);
nor U16445 (N_16445,N_15335,N_15431);
and U16446 (N_16446,N_15940,N_15504);
nand U16447 (N_16447,N_15992,N_15447);
nand U16448 (N_16448,N_15045,N_15791);
nand U16449 (N_16449,N_15787,N_15309);
nand U16450 (N_16450,N_15310,N_15792);
nand U16451 (N_16451,N_15272,N_15601);
nor U16452 (N_16452,N_15422,N_15406);
nand U16453 (N_16453,N_15212,N_15902);
xor U16454 (N_16454,N_15186,N_15774);
or U16455 (N_16455,N_15127,N_15024);
nand U16456 (N_16456,N_15122,N_15982);
nor U16457 (N_16457,N_15057,N_15697);
nor U16458 (N_16458,N_15609,N_15485);
or U16459 (N_16459,N_15343,N_15554);
nor U16460 (N_16460,N_15205,N_15267);
nand U16461 (N_16461,N_15247,N_15275);
nor U16462 (N_16462,N_15548,N_15210);
xnor U16463 (N_16463,N_15449,N_15905);
and U16464 (N_16464,N_15238,N_15034);
nand U16465 (N_16465,N_15931,N_15903);
and U16466 (N_16466,N_15072,N_15465);
nand U16467 (N_16467,N_15616,N_15017);
xor U16468 (N_16468,N_15508,N_15166);
nor U16469 (N_16469,N_15044,N_15366);
nand U16470 (N_16470,N_15463,N_15011);
xor U16471 (N_16471,N_15149,N_15232);
or U16472 (N_16472,N_15471,N_15505);
nand U16473 (N_16473,N_15233,N_15955);
xor U16474 (N_16474,N_15236,N_15742);
nor U16475 (N_16475,N_15332,N_15512);
xnor U16476 (N_16476,N_15912,N_15043);
nor U16477 (N_16477,N_15662,N_15775);
nand U16478 (N_16478,N_15611,N_15847);
or U16479 (N_16479,N_15182,N_15720);
nor U16480 (N_16480,N_15665,N_15822);
nand U16481 (N_16481,N_15371,N_15483);
and U16482 (N_16482,N_15522,N_15567);
xnor U16483 (N_16483,N_15947,N_15525);
nor U16484 (N_16484,N_15936,N_15030);
xor U16485 (N_16485,N_15479,N_15407);
xor U16486 (N_16486,N_15617,N_15314);
xnor U16487 (N_16487,N_15390,N_15797);
nor U16488 (N_16488,N_15142,N_15491);
or U16489 (N_16489,N_15573,N_15736);
nand U16490 (N_16490,N_15682,N_15421);
or U16491 (N_16491,N_15042,N_15380);
xnor U16492 (N_16492,N_15179,N_15845);
and U16493 (N_16493,N_15923,N_15085);
and U16494 (N_16494,N_15520,N_15196);
and U16495 (N_16495,N_15093,N_15106);
or U16496 (N_16496,N_15118,N_15676);
xnor U16497 (N_16497,N_15000,N_15136);
or U16498 (N_16498,N_15065,N_15412);
nand U16499 (N_16499,N_15080,N_15021);
and U16500 (N_16500,N_15930,N_15753);
and U16501 (N_16501,N_15762,N_15310);
and U16502 (N_16502,N_15384,N_15528);
xnor U16503 (N_16503,N_15637,N_15777);
or U16504 (N_16504,N_15531,N_15734);
and U16505 (N_16505,N_15820,N_15448);
nand U16506 (N_16506,N_15312,N_15829);
xnor U16507 (N_16507,N_15033,N_15025);
and U16508 (N_16508,N_15496,N_15599);
nor U16509 (N_16509,N_15433,N_15078);
or U16510 (N_16510,N_15245,N_15189);
xor U16511 (N_16511,N_15688,N_15877);
or U16512 (N_16512,N_15019,N_15423);
nand U16513 (N_16513,N_15851,N_15137);
or U16514 (N_16514,N_15316,N_15970);
or U16515 (N_16515,N_15329,N_15728);
and U16516 (N_16516,N_15836,N_15798);
nor U16517 (N_16517,N_15729,N_15099);
and U16518 (N_16518,N_15636,N_15248);
and U16519 (N_16519,N_15889,N_15314);
nand U16520 (N_16520,N_15476,N_15115);
nand U16521 (N_16521,N_15408,N_15502);
nand U16522 (N_16522,N_15592,N_15582);
xnor U16523 (N_16523,N_15016,N_15979);
nand U16524 (N_16524,N_15173,N_15426);
xnor U16525 (N_16525,N_15020,N_15944);
nor U16526 (N_16526,N_15306,N_15097);
nand U16527 (N_16527,N_15343,N_15053);
xnor U16528 (N_16528,N_15047,N_15294);
and U16529 (N_16529,N_15567,N_15162);
xor U16530 (N_16530,N_15306,N_15477);
and U16531 (N_16531,N_15937,N_15013);
or U16532 (N_16532,N_15751,N_15429);
and U16533 (N_16533,N_15940,N_15356);
xnor U16534 (N_16534,N_15064,N_15142);
or U16535 (N_16535,N_15089,N_15880);
xor U16536 (N_16536,N_15158,N_15088);
nor U16537 (N_16537,N_15559,N_15297);
nand U16538 (N_16538,N_15415,N_15836);
nand U16539 (N_16539,N_15850,N_15291);
or U16540 (N_16540,N_15853,N_15071);
nand U16541 (N_16541,N_15462,N_15599);
xor U16542 (N_16542,N_15017,N_15263);
xnor U16543 (N_16543,N_15886,N_15380);
xor U16544 (N_16544,N_15708,N_15697);
nor U16545 (N_16545,N_15450,N_15216);
and U16546 (N_16546,N_15071,N_15899);
nand U16547 (N_16547,N_15769,N_15962);
nand U16548 (N_16548,N_15768,N_15457);
nor U16549 (N_16549,N_15264,N_15322);
nor U16550 (N_16550,N_15914,N_15279);
or U16551 (N_16551,N_15626,N_15941);
and U16552 (N_16552,N_15012,N_15887);
nor U16553 (N_16553,N_15021,N_15317);
and U16554 (N_16554,N_15635,N_15719);
nand U16555 (N_16555,N_15754,N_15235);
or U16556 (N_16556,N_15334,N_15934);
or U16557 (N_16557,N_15561,N_15554);
xnor U16558 (N_16558,N_15160,N_15647);
and U16559 (N_16559,N_15284,N_15759);
nand U16560 (N_16560,N_15422,N_15171);
xnor U16561 (N_16561,N_15613,N_15703);
nor U16562 (N_16562,N_15050,N_15660);
nor U16563 (N_16563,N_15896,N_15525);
xor U16564 (N_16564,N_15551,N_15245);
nor U16565 (N_16565,N_15747,N_15816);
or U16566 (N_16566,N_15386,N_15927);
nand U16567 (N_16567,N_15366,N_15585);
xor U16568 (N_16568,N_15613,N_15003);
xor U16569 (N_16569,N_15093,N_15038);
or U16570 (N_16570,N_15993,N_15885);
and U16571 (N_16571,N_15494,N_15897);
or U16572 (N_16572,N_15646,N_15679);
xnor U16573 (N_16573,N_15081,N_15304);
nor U16574 (N_16574,N_15667,N_15278);
and U16575 (N_16575,N_15240,N_15826);
nand U16576 (N_16576,N_15110,N_15042);
nor U16577 (N_16577,N_15661,N_15523);
xnor U16578 (N_16578,N_15197,N_15181);
and U16579 (N_16579,N_15605,N_15693);
and U16580 (N_16580,N_15639,N_15910);
xnor U16581 (N_16581,N_15697,N_15328);
and U16582 (N_16582,N_15901,N_15392);
and U16583 (N_16583,N_15995,N_15586);
and U16584 (N_16584,N_15682,N_15134);
nor U16585 (N_16585,N_15646,N_15092);
nor U16586 (N_16586,N_15434,N_15973);
xor U16587 (N_16587,N_15699,N_15354);
nor U16588 (N_16588,N_15840,N_15949);
and U16589 (N_16589,N_15169,N_15382);
xor U16590 (N_16590,N_15385,N_15411);
nor U16591 (N_16591,N_15788,N_15428);
or U16592 (N_16592,N_15683,N_15347);
nor U16593 (N_16593,N_15713,N_15014);
and U16594 (N_16594,N_15357,N_15370);
nand U16595 (N_16595,N_15502,N_15364);
nand U16596 (N_16596,N_15013,N_15085);
nand U16597 (N_16597,N_15866,N_15232);
nor U16598 (N_16598,N_15316,N_15742);
or U16599 (N_16599,N_15720,N_15749);
nand U16600 (N_16600,N_15349,N_15957);
or U16601 (N_16601,N_15449,N_15892);
and U16602 (N_16602,N_15010,N_15181);
or U16603 (N_16603,N_15686,N_15382);
nor U16604 (N_16604,N_15484,N_15501);
xnor U16605 (N_16605,N_15360,N_15895);
xnor U16606 (N_16606,N_15975,N_15867);
and U16607 (N_16607,N_15021,N_15559);
nand U16608 (N_16608,N_15303,N_15025);
nand U16609 (N_16609,N_15796,N_15458);
nand U16610 (N_16610,N_15300,N_15103);
xnor U16611 (N_16611,N_15371,N_15058);
nor U16612 (N_16612,N_15473,N_15172);
nor U16613 (N_16613,N_15688,N_15718);
and U16614 (N_16614,N_15623,N_15952);
and U16615 (N_16615,N_15571,N_15609);
xor U16616 (N_16616,N_15628,N_15764);
xor U16617 (N_16617,N_15338,N_15217);
nand U16618 (N_16618,N_15858,N_15476);
nor U16619 (N_16619,N_15920,N_15943);
xnor U16620 (N_16620,N_15852,N_15658);
xor U16621 (N_16621,N_15293,N_15336);
xor U16622 (N_16622,N_15963,N_15752);
and U16623 (N_16623,N_15690,N_15471);
or U16624 (N_16624,N_15304,N_15880);
or U16625 (N_16625,N_15871,N_15555);
nand U16626 (N_16626,N_15263,N_15096);
nor U16627 (N_16627,N_15646,N_15757);
nand U16628 (N_16628,N_15481,N_15015);
and U16629 (N_16629,N_15250,N_15944);
nand U16630 (N_16630,N_15710,N_15501);
or U16631 (N_16631,N_15136,N_15853);
nor U16632 (N_16632,N_15597,N_15694);
xnor U16633 (N_16633,N_15116,N_15915);
nor U16634 (N_16634,N_15550,N_15418);
or U16635 (N_16635,N_15555,N_15598);
or U16636 (N_16636,N_15147,N_15868);
nand U16637 (N_16637,N_15465,N_15500);
nand U16638 (N_16638,N_15475,N_15662);
nor U16639 (N_16639,N_15021,N_15101);
xnor U16640 (N_16640,N_15869,N_15304);
nor U16641 (N_16641,N_15090,N_15115);
nor U16642 (N_16642,N_15355,N_15584);
nor U16643 (N_16643,N_15691,N_15677);
nor U16644 (N_16644,N_15261,N_15087);
xor U16645 (N_16645,N_15635,N_15069);
nand U16646 (N_16646,N_15201,N_15649);
and U16647 (N_16647,N_15982,N_15495);
nor U16648 (N_16648,N_15548,N_15493);
xnor U16649 (N_16649,N_15408,N_15926);
and U16650 (N_16650,N_15665,N_15975);
and U16651 (N_16651,N_15381,N_15799);
or U16652 (N_16652,N_15831,N_15016);
xnor U16653 (N_16653,N_15259,N_15695);
and U16654 (N_16654,N_15963,N_15530);
nor U16655 (N_16655,N_15219,N_15236);
xor U16656 (N_16656,N_15976,N_15794);
xor U16657 (N_16657,N_15774,N_15558);
xnor U16658 (N_16658,N_15120,N_15654);
and U16659 (N_16659,N_15246,N_15824);
nor U16660 (N_16660,N_15567,N_15149);
nor U16661 (N_16661,N_15062,N_15165);
or U16662 (N_16662,N_15746,N_15512);
and U16663 (N_16663,N_15001,N_15004);
or U16664 (N_16664,N_15220,N_15097);
nor U16665 (N_16665,N_15331,N_15976);
nand U16666 (N_16666,N_15986,N_15264);
nor U16667 (N_16667,N_15946,N_15242);
nand U16668 (N_16668,N_15960,N_15685);
nor U16669 (N_16669,N_15575,N_15016);
nor U16670 (N_16670,N_15874,N_15134);
or U16671 (N_16671,N_15476,N_15171);
and U16672 (N_16672,N_15251,N_15220);
and U16673 (N_16673,N_15249,N_15082);
nor U16674 (N_16674,N_15755,N_15454);
nand U16675 (N_16675,N_15642,N_15605);
and U16676 (N_16676,N_15919,N_15371);
nand U16677 (N_16677,N_15636,N_15552);
and U16678 (N_16678,N_15941,N_15048);
nor U16679 (N_16679,N_15691,N_15623);
nor U16680 (N_16680,N_15084,N_15140);
nand U16681 (N_16681,N_15050,N_15460);
and U16682 (N_16682,N_15362,N_15746);
xor U16683 (N_16683,N_15030,N_15337);
nor U16684 (N_16684,N_15850,N_15842);
nand U16685 (N_16685,N_15545,N_15791);
nor U16686 (N_16686,N_15066,N_15914);
nor U16687 (N_16687,N_15159,N_15187);
xor U16688 (N_16688,N_15020,N_15101);
and U16689 (N_16689,N_15572,N_15433);
or U16690 (N_16690,N_15659,N_15994);
nor U16691 (N_16691,N_15007,N_15316);
and U16692 (N_16692,N_15762,N_15549);
xnor U16693 (N_16693,N_15193,N_15002);
or U16694 (N_16694,N_15354,N_15794);
xor U16695 (N_16695,N_15202,N_15613);
nor U16696 (N_16696,N_15024,N_15104);
or U16697 (N_16697,N_15910,N_15158);
xor U16698 (N_16698,N_15388,N_15438);
nor U16699 (N_16699,N_15443,N_15419);
nor U16700 (N_16700,N_15637,N_15975);
nand U16701 (N_16701,N_15547,N_15368);
nor U16702 (N_16702,N_15776,N_15319);
and U16703 (N_16703,N_15848,N_15695);
nor U16704 (N_16704,N_15709,N_15734);
and U16705 (N_16705,N_15432,N_15372);
nor U16706 (N_16706,N_15831,N_15034);
and U16707 (N_16707,N_15675,N_15948);
or U16708 (N_16708,N_15020,N_15411);
nand U16709 (N_16709,N_15267,N_15865);
xnor U16710 (N_16710,N_15376,N_15732);
and U16711 (N_16711,N_15040,N_15434);
xor U16712 (N_16712,N_15579,N_15652);
and U16713 (N_16713,N_15380,N_15031);
nor U16714 (N_16714,N_15304,N_15549);
nor U16715 (N_16715,N_15750,N_15991);
nand U16716 (N_16716,N_15339,N_15030);
or U16717 (N_16717,N_15088,N_15894);
nand U16718 (N_16718,N_15752,N_15039);
nand U16719 (N_16719,N_15773,N_15870);
nand U16720 (N_16720,N_15401,N_15246);
nand U16721 (N_16721,N_15158,N_15200);
nand U16722 (N_16722,N_15686,N_15781);
nor U16723 (N_16723,N_15670,N_15778);
or U16724 (N_16724,N_15000,N_15367);
and U16725 (N_16725,N_15197,N_15480);
or U16726 (N_16726,N_15962,N_15334);
xnor U16727 (N_16727,N_15708,N_15137);
or U16728 (N_16728,N_15471,N_15899);
nor U16729 (N_16729,N_15184,N_15154);
or U16730 (N_16730,N_15534,N_15742);
or U16731 (N_16731,N_15817,N_15423);
and U16732 (N_16732,N_15409,N_15279);
nor U16733 (N_16733,N_15214,N_15018);
nand U16734 (N_16734,N_15662,N_15367);
and U16735 (N_16735,N_15598,N_15759);
and U16736 (N_16736,N_15427,N_15284);
nor U16737 (N_16737,N_15445,N_15137);
and U16738 (N_16738,N_15472,N_15936);
nor U16739 (N_16739,N_15359,N_15459);
and U16740 (N_16740,N_15423,N_15515);
or U16741 (N_16741,N_15949,N_15413);
or U16742 (N_16742,N_15498,N_15238);
and U16743 (N_16743,N_15173,N_15219);
or U16744 (N_16744,N_15286,N_15891);
and U16745 (N_16745,N_15835,N_15122);
nor U16746 (N_16746,N_15141,N_15154);
nand U16747 (N_16747,N_15296,N_15985);
nor U16748 (N_16748,N_15433,N_15121);
or U16749 (N_16749,N_15799,N_15845);
xnor U16750 (N_16750,N_15054,N_15112);
and U16751 (N_16751,N_15512,N_15377);
and U16752 (N_16752,N_15378,N_15962);
nor U16753 (N_16753,N_15224,N_15815);
xor U16754 (N_16754,N_15239,N_15253);
or U16755 (N_16755,N_15472,N_15242);
nand U16756 (N_16756,N_15928,N_15197);
xor U16757 (N_16757,N_15664,N_15898);
nor U16758 (N_16758,N_15766,N_15344);
xnor U16759 (N_16759,N_15251,N_15300);
nand U16760 (N_16760,N_15539,N_15970);
nor U16761 (N_16761,N_15739,N_15414);
or U16762 (N_16762,N_15313,N_15120);
and U16763 (N_16763,N_15090,N_15353);
xnor U16764 (N_16764,N_15969,N_15537);
nor U16765 (N_16765,N_15692,N_15259);
nor U16766 (N_16766,N_15325,N_15938);
nor U16767 (N_16767,N_15274,N_15696);
and U16768 (N_16768,N_15421,N_15011);
nor U16769 (N_16769,N_15722,N_15190);
and U16770 (N_16770,N_15508,N_15617);
or U16771 (N_16771,N_15865,N_15710);
nor U16772 (N_16772,N_15669,N_15914);
nand U16773 (N_16773,N_15887,N_15135);
and U16774 (N_16774,N_15018,N_15100);
and U16775 (N_16775,N_15735,N_15679);
nor U16776 (N_16776,N_15447,N_15038);
and U16777 (N_16777,N_15782,N_15237);
and U16778 (N_16778,N_15227,N_15730);
xor U16779 (N_16779,N_15093,N_15384);
nor U16780 (N_16780,N_15330,N_15434);
xnor U16781 (N_16781,N_15500,N_15415);
or U16782 (N_16782,N_15403,N_15192);
or U16783 (N_16783,N_15859,N_15100);
and U16784 (N_16784,N_15049,N_15055);
nand U16785 (N_16785,N_15806,N_15659);
nand U16786 (N_16786,N_15857,N_15111);
nand U16787 (N_16787,N_15414,N_15758);
nand U16788 (N_16788,N_15786,N_15134);
xnor U16789 (N_16789,N_15022,N_15316);
xor U16790 (N_16790,N_15492,N_15761);
and U16791 (N_16791,N_15329,N_15759);
or U16792 (N_16792,N_15196,N_15638);
xor U16793 (N_16793,N_15431,N_15741);
nor U16794 (N_16794,N_15245,N_15847);
and U16795 (N_16795,N_15302,N_15238);
nor U16796 (N_16796,N_15850,N_15513);
nand U16797 (N_16797,N_15801,N_15905);
and U16798 (N_16798,N_15339,N_15703);
xnor U16799 (N_16799,N_15285,N_15891);
or U16800 (N_16800,N_15591,N_15301);
nand U16801 (N_16801,N_15772,N_15696);
or U16802 (N_16802,N_15394,N_15116);
and U16803 (N_16803,N_15205,N_15879);
nand U16804 (N_16804,N_15303,N_15196);
and U16805 (N_16805,N_15975,N_15003);
nand U16806 (N_16806,N_15728,N_15451);
nor U16807 (N_16807,N_15570,N_15885);
nand U16808 (N_16808,N_15628,N_15531);
and U16809 (N_16809,N_15187,N_15905);
nand U16810 (N_16810,N_15822,N_15606);
nor U16811 (N_16811,N_15330,N_15260);
and U16812 (N_16812,N_15167,N_15323);
xnor U16813 (N_16813,N_15331,N_15118);
and U16814 (N_16814,N_15161,N_15213);
and U16815 (N_16815,N_15229,N_15722);
and U16816 (N_16816,N_15457,N_15092);
and U16817 (N_16817,N_15302,N_15942);
or U16818 (N_16818,N_15680,N_15968);
nand U16819 (N_16819,N_15567,N_15308);
nand U16820 (N_16820,N_15417,N_15548);
or U16821 (N_16821,N_15397,N_15021);
xor U16822 (N_16822,N_15517,N_15523);
nor U16823 (N_16823,N_15290,N_15808);
and U16824 (N_16824,N_15173,N_15395);
or U16825 (N_16825,N_15946,N_15668);
or U16826 (N_16826,N_15306,N_15664);
nand U16827 (N_16827,N_15815,N_15516);
or U16828 (N_16828,N_15639,N_15847);
and U16829 (N_16829,N_15383,N_15723);
nor U16830 (N_16830,N_15963,N_15106);
nand U16831 (N_16831,N_15557,N_15559);
xnor U16832 (N_16832,N_15041,N_15222);
and U16833 (N_16833,N_15755,N_15914);
and U16834 (N_16834,N_15559,N_15625);
xnor U16835 (N_16835,N_15741,N_15919);
xor U16836 (N_16836,N_15608,N_15970);
nand U16837 (N_16837,N_15030,N_15465);
nand U16838 (N_16838,N_15394,N_15407);
xor U16839 (N_16839,N_15250,N_15612);
or U16840 (N_16840,N_15488,N_15089);
nand U16841 (N_16841,N_15494,N_15535);
nand U16842 (N_16842,N_15196,N_15836);
and U16843 (N_16843,N_15726,N_15271);
or U16844 (N_16844,N_15979,N_15413);
nor U16845 (N_16845,N_15553,N_15263);
nor U16846 (N_16846,N_15248,N_15120);
nand U16847 (N_16847,N_15423,N_15972);
nand U16848 (N_16848,N_15590,N_15909);
nor U16849 (N_16849,N_15298,N_15766);
nor U16850 (N_16850,N_15316,N_15865);
or U16851 (N_16851,N_15232,N_15698);
nor U16852 (N_16852,N_15847,N_15160);
nor U16853 (N_16853,N_15606,N_15995);
nand U16854 (N_16854,N_15621,N_15694);
nand U16855 (N_16855,N_15753,N_15427);
xor U16856 (N_16856,N_15746,N_15520);
xnor U16857 (N_16857,N_15674,N_15498);
and U16858 (N_16858,N_15880,N_15277);
or U16859 (N_16859,N_15209,N_15837);
nor U16860 (N_16860,N_15435,N_15940);
or U16861 (N_16861,N_15834,N_15752);
nor U16862 (N_16862,N_15691,N_15158);
xor U16863 (N_16863,N_15029,N_15376);
nor U16864 (N_16864,N_15209,N_15267);
nor U16865 (N_16865,N_15015,N_15990);
xnor U16866 (N_16866,N_15283,N_15243);
or U16867 (N_16867,N_15537,N_15562);
nor U16868 (N_16868,N_15857,N_15869);
and U16869 (N_16869,N_15838,N_15874);
or U16870 (N_16870,N_15321,N_15008);
nand U16871 (N_16871,N_15548,N_15419);
nor U16872 (N_16872,N_15893,N_15063);
or U16873 (N_16873,N_15365,N_15094);
or U16874 (N_16874,N_15946,N_15925);
nor U16875 (N_16875,N_15957,N_15191);
and U16876 (N_16876,N_15483,N_15687);
xor U16877 (N_16877,N_15611,N_15708);
nor U16878 (N_16878,N_15432,N_15780);
and U16879 (N_16879,N_15780,N_15719);
nand U16880 (N_16880,N_15072,N_15683);
xor U16881 (N_16881,N_15850,N_15532);
nand U16882 (N_16882,N_15943,N_15303);
nand U16883 (N_16883,N_15542,N_15943);
or U16884 (N_16884,N_15850,N_15396);
nand U16885 (N_16885,N_15488,N_15902);
or U16886 (N_16886,N_15274,N_15987);
nand U16887 (N_16887,N_15899,N_15904);
nor U16888 (N_16888,N_15944,N_15698);
nor U16889 (N_16889,N_15967,N_15855);
nor U16890 (N_16890,N_15913,N_15464);
xnor U16891 (N_16891,N_15108,N_15931);
xor U16892 (N_16892,N_15875,N_15782);
and U16893 (N_16893,N_15001,N_15917);
nor U16894 (N_16894,N_15809,N_15637);
nor U16895 (N_16895,N_15501,N_15370);
or U16896 (N_16896,N_15812,N_15193);
xor U16897 (N_16897,N_15663,N_15911);
xnor U16898 (N_16898,N_15672,N_15434);
and U16899 (N_16899,N_15534,N_15597);
and U16900 (N_16900,N_15350,N_15743);
nor U16901 (N_16901,N_15407,N_15030);
and U16902 (N_16902,N_15620,N_15761);
or U16903 (N_16903,N_15141,N_15380);
and U16904 (N_16904,N_15240,N_15856);
nand U16905 (N_16905,N_15513,N_15047);
nand U16906 (N_16906,N_15610,N_15822);
xor U16907 (N_16907,N_15505,N_15854);
nor U16908 (N_16908,N_15397,N_15823);
nor U16909 (N_16909,N_15570,N_15340);
nand U16910 (N_16910,N_15644,N_15325);
xnor U16911 (N_16911,N_15627,N_15811);
nor U16912 (N_16912,N_15791,N_15593);
xnor U16913 (N_16913,N_15496,N_15212);
and U16914 (N_16914,N_15666,N_15374);
nor U16915 (N_16915,N_15304,N_15091);
or U16916 (N_16916,N_15852,N_15794);
and U16917 (N_16917,N_15360,N_15411);
and U16918 (N_16918,N_15426,N_15998);
nor U16919 (N_16919,N_15251,N_15061);
nand U16920 (N_16920,N_15284,N_15472);
xnor U16921 (N_16921,N_15129,N_15105);
xnor U16922 (N_16922,N_15352,N_15448);
xor U16923 (N_16923,N_15929,N_15998);
nor U16924 (N_16924,N_15185,N_15298);
nor U16925 (N_16925,N_15468,N_15361);
xnor U16926 (N_16926,N_15021,N_15807);
nand U16927 (N_16927,N_15045,N_15247);
and U16928 (N_16928,N_15087,N_15859);
nor U16929 (N_16929,N_15870,N_15308);
or U16930 (N_16930,N_15338,N_15326);
nor U16931 (N_16931,N_15235,N_15591);
and U16932 (N_16932,N_15891,N_15067);
nand U16933 (N_16933,N_15347,N_15577);
nand U16934 (N_16934,N_15111,N_15893);
nand U16935 (N_16935,N_15995,N_15566);
and U16936 (N_16936,N_15729,N_15035);
xor U16937 (N_16937,N_15352,N_15761);
or U16938 (N_16938,N_15031,N_15717);
xor U16939 (N_16939,N_15922,N_15167);
and U16940 (N_16940,N_15921,N_15722);
or U16941 (N_16941,N_15075,N_15716);
nor U16942 (N_16942,N_15529,N_15026);
xnor U16943 (N_16943,N_15013,N_15506);
nand U16944 (N_16944,N_15190,N_15360);
nor U16945 (N_16945,N_15222,N_15993);
and U16946 (N_16946,N_15929,N_15574);
xnor U16947 (N_16947,N_15768,N_15352);
and U16948 (N_16948,N_15109,N_15208);
nor U16949 (N_16949,N_15555,N_15241);
xor U16950 (N_16950,N_15236,N_15447);
or U16951 (N_16951,N_15921,N_15254);
xnor U16952 (N_16952,N_15666,N_15581);
and U16953 (N_16953,N_15865,N_15479);
or U16954 (N_16954,N_15773,N_15237);
or U16955 (N_16955,N_15231,N_15018);
xor U16956 (N_16956,N_15104,N_15265);
nand U16957 (N_16957,N_15033,N_15103);
nand U16958 (N_16958,N_15704,N_15794);
nor U16959 (N_16959,N_15805,N_15215);
and U16960 (N_16960,N_15325,N_15800);
xnor U16961 (N_16961,N_15972,N_15617);
nor U16962 (N_16962,N_15877,N_15952);
or U16963 (N_16963,N_15111,N_15679);
nand U16964 (N_16964,N_15822,N_15246);
and U16965 (N_16965,N_15081,N_15351);
nor U16966 (N_16966,N_15906,N_15654);
nand U16967 (N_16967,N_15779,N_15158);
xor U16968 (N_16968,N_15963,N_15375);
or U16969 (N_16969,N_15693,N_15714);
nand U16970 (N_16970,N_15498,N_15882);
xnor U16971 (N_16971,N_15640,N_15707);
and U16972 (N_16972,N_15602,N_15981);
xnor U16973 (N_16973,N_15521,N_15979);
xor U16974 (N_16974,N_15009,N_15185);
nand U16975 (N_16975,N_15380,N_15191);
xor U16976 (N_16976,N_15463,N_15570);
xnor U16977 (N_16977,N_15838,N_15360);
nor U16978 (N_16978,N_15276,N_15968);
and U16979 (N_16979,N_15862,N_15055);
xnor U16980 (N_16980,N_15661,N_15658);
xor U16981 (N_16981,N_15169,N_15220);
and U16982 (N_16982,N_15666,N_15091);
or U16983 (N_16983,N_15005,N_15244);
nand U16984 (N_16984,N_15004,N_15008);
nand U16985 (N_16985,N_15668,N_15147);
nand U16986 (N_16986,N_15482,N_15063);
and U16987 (N_16987,N_15936,N_15444);
or U16988 (N_16988,N_15493,N_15440);
xnor U16989 (N_16989,N_15092,N_15116);
nand U16990 (N_16990,N_15412,N_15369);
or U16991 (N_16991,N_15010,N_15354);
nand U16992 (N_16992,N_15444,N_15312);
xor U16993 (N_16993,N_15485,N_15092);
nand U16994 (N_16994,N_15590,N_15814);
nor U16995 (N_16995,N_15339,N_15461);
nand U16996 (N_16996,N_15226,N_15694);
and U16997 (N_16997,N_15108,N_15573);
and U16998 (N_16998,N_15116,N_15583);
or U16999 (N_16999,N_15304,N_15031);
xor U17000 (N_17000,N_16234,N_16328);
or U17001 (N_17001,N_16284,N_16573);
xnor U17002 (N_17002,N_16504,N_16743);
or U17003 (N_17003,N_16636,N_16276);
and U17004 (N_17004,N_16507,N_16736);
xor U17005 (N_17005,N_16825,N_16875);
nor U17006 (N_17006,N_16505,N_16126);
nor U17007 (N_17007,N_16991,N_16033);
and U17008 (N_17008,N_16125,N_16025);
nor U17009 (N_17009,N_16790,N_16352);
or U17010 (N_17010,N_16915,N_16784);
nor U17011 (N_17011,N_16364,N_16057);
nor U17012 (N_17012,N_16031,N_16828);
and U17013 (N_17013,N_16942,N_16479);
xor U17014 (N_17014,N_16270,N_16837);
xor U17015 (N_17015,N_16229,N_16590);
xor U17016 (N_17016,N_16386,N_16698);
nand U17017 (N_17017,N_16461,N_16560);
nor U17018 (N_17018,N_16946,N_16570);
and U17019 (N_17019,N_16685,N_16975);
nor U17020 (N_17020,N_16863,N_16580);
nand U17021 (N_17021,N_16655,N_16832);
nand U17022 (N_17022,N_16508,N_16645);
or U17023 (N_17023,N_16422,N_16150);
nor U17024 (N_17024,N_16236,N_16435);
or U17025 (N_17025,N_16895,N_16943);
nand U17026 (N_17026,N_16225,N_16614);
and U17027 (N_17027,N_16420,N_16317);
nand U17028 (N_17028,N_16205,N_16273);
and U17029 (N_17029,N_16522,N_16601);
nor U17030 (N_17030,N_16515,N_16903);
and U17031 (N_17031,N_16774,N_16059);
or U17032 (N_17032,N_16390,N_16687);
nand U17033 (N_17033,N_16671,N_16230);
nand U17034 (N_17034,N_16106,N_16546);
or U17035 (N_17035,N_16379,N_16779);
nor U17036 (N_17036,N_16078,N_16908);
nor U17037 (N_17037,N_16968,N_16694);
or U17038 (N_17038,N_16289,N_16921);
nand U17039 (N_17039,N_16410,N_16215);
or U17040 (N_17040,N_16082,N_16911);
nor U17041 (N_17041,N_16416,N_16535);
xor U17042 (N_17042,N_16684,N_16491);
and U17043 (N_17043,N_16476,N_16114);
nand U17044 (N_17044,N_16143,N_16311);
and U17045 (N_17045,N_16353,N_16745);
or U17046 (N_17046,N_16428,N_16979);
nor U17047 (N_17047,N_16224,N_16824);
nand U17048 (N_17048,N_16001,N_16563);
xor U17049 (N_17049,N_16957,N_16287);
or U17050 (N_17050,N_16530,N_16608);
nor U17051 (N_17051,N_16089,N_16301);
xor U17052 (N_17052,N_16906,N_16540);
nand U17053 (N_17053,N_16757,N_16355);
and U17054 (N_17054,N_16233,N_16753);
xnor U17055 (N_17055,N_16146,N_16278);
nand U17056 (N_17056,N_16549,N_16831);
nor U17057 (N_17057,N_16673,N_16241);
xnor U17058 (N_17058,N_16552,N_16962);
xor U17059 (N_17059,N_16760,N_16266);
xnor U17060 (N_17060,N_16814,N_16262);
and U17061 (N_17061,N_16648,N_16376);
xor U17062 (N_17062,N_16396,N_16258);
and U17063 (N_17063,N_16228,N_16852);
nor U17064 (N_17064,N_16080,N_16538);
nor U17065 (N_17065,N_16367,N_16937);
nand U17066 (N_17066,N_16938,N_16475);
and U17067 (N_17067,N_16609,N_16749);
xnor U17068 (N_17068,N_16292,N_16693);
or U17069 (N_17069,N_16716,N_16706);
or U17070 (N_17070,N_16800,N_16669);
xnor U17071 (N_17071,N_16659,N_16347);
and U17072 (N_17072,N_16513,N_16995);
and U17073 (N_17073,N_16081,N_16223);
or U17074 (N_17074,N_16815,N_16724);
or U17075 (N_17075,N_16419,N_16285);
xor U17076 (N_17076,N_16260,N_16633);
and U17077 (N_17077,N_16312,N_16652);
nor U17078 (N_17078,N_16014,N_16849);
and U17079 (N_17079,N_16544,N_16254);
nand U17080 (N_17080,N_16854,N_16060);
nor U17081 (N_17081,N_16209,N_16697);
xor U17082 (N_17082,N_16462,N_16742);
nor U17083 (N_17083,N_16071,N_16850);
xor U17084 (N_17084,N_16555,N_16313);
nand U17085 (N_17085,N_16756,N_16041);
nand U17086 (N_17086,N_16630,N_16651);
nor U17087 (N_17087,N_16926,N_16583);
or U17088 (N_17088,N_16750,N_16067);
nor U17089 (N_17089,N_16965,N_16076);
xor U17090 (N_17090,N_16758,N_16378);
or U17091 (N_17091,N_16449,N_16898);
and U17092 (N_17092,N_16551,N_16454);
nor U17093 (N_17093,N_16877,N_16914);
nor U17094 (N_17094,N_16415,N_16199);
nor U17095 (N_17095,N_16620,N_16565);
xnor U17096 (N_17096,N_16291,N_16783);
or U17097 (N_17097,N_16781,N_16424);
and U17098 (N_17098,N_16807,N_16759);
and U17099 (N_17099,N_16391,N_16872);
and U17100 (N_17100,N_16711,N_16763);
nand U17101 (N_17101,N_16070,N_16989);
or U17102 (N_17102,N_16941,N_16058);
and U17103 (N_17103,N_16145,N_16982);
or U17104 (N_17104,N_16998,N_16970);
and U17105 (N_17105,N_16463,N_16527);
nand U17106 (N_17106,N_16306,N_16383);
xor U17107 (N_17107,N_16747,N_16098);
or U17108 (N_17108,N_16598,N_16471);
nor U17109 (N_17109,N_16751,N_16715);
and U17110 (N_17110,N_16404,N_16548);
or U17111 (N_17111,N_16019,N_16296);
or U17112 (N_17112,N_16242,N_16531);
xor U17113 (N_17113,N_16350,N_16490);
xor U17114 (N_17114,N_16584,N_16916);
and U17115 (N_17115,N_16239,N_16048);
or U17116 (N_17116,N_16533,N_16662);
xor U17117 (N_17117,N_16572,N_16682);
and U17118 (N_17118,N_16618,N_16628);
and U17119 (N_17119,N_16919,N_16622);
xnor U17120 (N_17120,N_16936,N_16950);
xnor U17121 (N_17121,N_16528,N_16894);
or U17122 (N_17122,N_16023,N_16107);
and U17123 (N_17123,N_16331,N_16365);
nand U17124 (N_17124,N_16594,N_16720);
or U17125 (N_17125,N_16450,N_16692);
nor U17126 (N_17126,N_16585,N_16839);
and U17127 (N_17127,N_16882,N_16149);
nor U17128 (N_17128,N_16140,N_16641);
and U17129 (N_17129,N_16297,N_16887);
and U17130 (N_17130,N_16426,N_16413);
and U17131 (N_17131,N_16186,N_16249);
nor U17132 (N_17132,N_16918,N_16142);
and U17133 (N_17133,N_16827,N_16708);
nor U17134 (N_17134,N_16027,N_16073);
xnor U17135 (N_17135,N_16003,N_16137);
nor U17136 (N_17136,N_16309,N_16506);
nor U17137 (N_17137,N_16913,N_16826);
nand U17138 (N_17138,N_16823,N_16087);
or U17139 (N_17139,N_16370,N_16703);
or U17140 (N_17140,N_16524,N_16043);
xor U17141 (N_17141,N_16500,N_16445);
xor U17142 (N_17142,N_16980,N_16302);
xor U17143 (N_17143,N_16765,N_16927);
xor U17144 (N_17144,N_16002,N_16066);
nand U17145 (N_17145,N_16775,N_16681);
or U17146 (N_17146,N_16772,N_16737);
and U17147 (N_17147,N_16016,N_16611);
nand U17148 (N_17148,N_16885,N_16846);
xnor U17149 (N_17149,N_16740,N_16451);
or U17150 (N_17150,N_16647,N_16203);
nand U17151 (N_17151,N_16674,N_16656);
and U17152 (N_17152,N_16503,N_16252);
nand U17153 (N_17153,N_16351,N_16870);
xor U17154 (N_17154,N_16719,N_16575);
or U17155 (N_17155,N_16263,N_16932);
or U17156 (N_17156,N_16766,N_16382);
nor U17157 (N_17157,N_16187,N_16282);
nand U17158 (N_17158,N_16668,N_16822);
xor U17159 (N_17159,N_16362,N_16099);
nor U17160 (N_17160,N_16992,N_16017);
xnor U17161 (N_17161,N_16272,N_16201);
nand U17162 (N_17162,N_16256,N_16539);
nand U17163 (N_17163,N_16712,N_16893);
xnor U17164 (N_17164,N_16956,N_16268);
xor U17165 (N_17165,N_16444,N_16044);
and U17166 (N_17166,N_16933,N_16155);
and U17167 (N_17167,N_16801,N_16520);
nor U17168 (N_17168,N_16342,N_16469);
and U17169 (N_17169,N_16925,N_16380);
nor U17170 (N_17170,N_16477,N_16627);
xnor U17171 (N_17171,N_16954,N_16472);
xor U17172 (N_17172,N_16250,N_16564);
xnor U17173 (N_17173,N_16638,N_16189);
and U17174 (N_17174,N_16497,N_16452);
nor U17175 (N_17175,N_16381,N_16015);
and U17176 (N_17176,N_16153,N_16532);
xnor U17177 (N_17177,N_16458,N_16216);
nand U17178 (N_17178,N_16330,N_16349);
or U17179 (N_17179,N_16212,N_16789);
or U17180 (N_17180,N_16990,N_16022);
nand U17181 (N_17181,N_16884,N_16707);
xor U17182 (N_17182,N_16597,N_16664);
nor U17183 (N_17183,N_16574,N_16221);
nor U17184 (N_17184,N_16857,N_16935);
xnor U17185 (N_17185,N_16389,N_16493);
nor U17186 (N_17186,N_16734,N_16642);
nand U17187 (N_17187,N_16414,N_16295);
or U17188 (N_17188,N_16009,N_16222);
and U17189 (N_17189,N_16495,N_16421);
nand U17190 (N_17190,N_16586,N_16632);
xor U17191 (N_17191,N_16981,N_16514);
nand U17192 (N_17192,N_16136,N_16550);
and U17193 (N_17193,N_16206,N_16762);
nand U17194 (N_17194,N_16977,N_16996);
xor U17195 (N_17195,N_16269,N_16701);
xnor U17196 (N_17196,N_16246,N_16218);
xnor U17197 (N_17197,N_16964,N_16088);
nand U17198 (N_17198,N_16799,N_16714);
or U17199 (N_17199,N_16589,N_16045);
nand U17200 (N_17200,N_16348,N_16448);
xnor U17201 (N_17201,N_16190,N_16314);
and U17202 (N_17202,N_16072,N_16888);
nor U17203 (N_17203,N_16960,N_16804);
nand U17204 (N_17204,N_16244,N_16571);
xor U17205 (N_17205,N_16226,N_16130);
or U17206 (N_17206,N_16417,N_16034);
and U17207 (N_17207,N_16120,N_16326);
nand U17208 (N_17208,N_16184,N_16878);
xor U17209 (N_17209,N_16866,N_16357);
nand U17210 (N_17210,N_16690,N_16439);
nor U17211 (N_17211,N_16117,N_16631);
and U17212 (N_17212,N_16833,N_16780);
xor U17213 (N_17213,N_16786,N_16193);
xnor U17214 (N_17214,N_16769,N_16179);
nand U17215 (N_17215,N_16144,N_16696);
nand U17216 (N_17216,N_16333,N_16257);
xor U17217 (N_17217,N_16961,N_16492);
or U17218 (N_17218,N_16752,N_16024);
and U17219 (N_17219,N_16425,N_16891);
or U17220 (N_17220,N_16634,N_16337);
and U17221 (N_17221,N_16610,N_16124);
or U17222 (N_17222,N_16429,N_16049);
nor U17223 (N_17223,N_16579,N_16489);
and U17224 (N_17224,N_16930,N_16718);
xnor U17225 (N_17225,N_16324,N_16154);
xnor U17226 (N_17226,N_16722,N_16606);
and U17227 (N_17227,N_16578,N_16116);
or U17228 (N_17228,N_16896,N_16812);
nand U17229 (N_17229,N_16486,N_16602);
or U17230 (N_17230,N_16865,N_16660);
and U17231 (N_17231,N_16063,N_16679);
xor U17232 (N_17232,N_16148,N_16018);
nand U17233 (N_17233,N_16141,N_16680);
and U17234 (N_17234,N_16782,N_16286);
or U17235 (N_17235,N_16675,N_16838);
nand U17236 (N_17236,N_16274,N_16065);
nor U17237 (N_17237,N_16346,N_16561);
or U17238 (N_17238,N_16407,N_16227);
and U17239 (N_17239,N_16607,N_16110);
xor U17240 (N_17240,N_16183,N_16686);
or U17241 (N_17241,N_16171,N_16588);
xnor U17242 (N_17242,N_16086,N_16100);
nor U17243 (N_17243,N_16547,N_16678);
and U17244 (N_17244,N_16290,N_16710);
nand U17245 (N_17245,N_16537,N_16543);
nor U17246 (N_17246,N_16591,N_16195);
nor U17247 (N_17247,N_16947,N_16319);
and U17248 (N_17248,N_16835,N_16457);
nand U17249 (N_17249,N_16771,N_16188);
or U17250 (N_17250,N_16966,N_16859);
or U17251 (N_17251,N_16032,N_16177);
xor U17252 (N_17252,N_16643,N_16275);
xor U17253 (N_17253,N_16300,N_16200);
and U17254 (N_17254,N_16411,N_16976);
or U17255 (N_17255,N_16118,N_16358);
nand U17256 (N_17256,N_16851,N_16169);
nand U17257 (N_17257,N_16104,N_16917);
nand U17258 (N_17258,N_16880,N_16243);
xor U17259 (N_17259,N_16322,N_16595);
nor U17260 (N_17260,N_16341,N_16605);
and U17261 (N_17261,N_16501,N_16105);
nand U17262 (N_17262,N_16542,N_16219);
or U17263 (N_17263,N_16037,N_16094);
and U17264 (N_17264,N_16213,N_16480);
xor U17265 (N_17265,N_16581,N_16000);
xnor U17266 (N_17266,N_16972,N_16568);
nand U17267 (N_17267,N_16255,N_16123);
or U17268 (N_17268,N_16897,N_16619);
xor U17269 (N_17269,N_16847,N_16441);
nand U17270 (N_17270,N_16168,N_16375);
nor U17271 (N_17271,N_16802,N_16198);
nor U17272 (N_17272,N_16248,N_16646);
nor U17273 (N_17273,N_16876,N_16446);
nor U17274 (N_17274,N_16251,N_16517);
and U17275 (N_17275,N_16986,N_16470);
and U17276 (N_17276,N_16092,N_16303);
xnor U17277 (N_17277,N_16820,N_16418);
xnor U17278 (N_17278,N_16119,N_16423);
xnor U17279 (N_17279,N_16384,N_16661);
or U17280 (N_17280,N_16436,N_16283);
nor U17281 (N_17281,N_16855,N_16777);
and U17282 (N_17282,N_16402,N_16744);
nand U17283 (N_17283,N_16554,N_16253);
nor U17284 (N_17284,N_16008,N_16385);
nor U17285 (N_17285,N_16558,N_16377);
nor U17286 (N_17286,N_16408,N_16304);
and U17287 (N_17287,N_16810,N_16062);
xnor U17288 (N_17288,N_16929,N_16180);
nand U17289 (N_17289,N_16709,N_16967);
or U17290 (N_17290,N_16856,N_16879);
or U17291 (N_17291,N_16139,N_16842);
nand U17292 (N_17292,N_16085,N_16280);
and U17293 (N_17293,N_16658,N_16288);
and U17294 (N_17294,N_16746,N_16944);
nand U17295 (N_17295,N_16393,N_16987);
and U17296 (N_17296,N_16705,N_16483);
xnor U17297 (N_17297,N_16321,N_16232);
and U17298 (N_17298,N_16738,N_16728);
or U17299 (N_17299,N_16841,N_16629);
and U17300 (N_17300,N_16923,N_16768);
and U17301 (N_17301,N_16848,N_16134);
nor U17302 (N_17302,N_16398,N_16005);
or U17303 (N_17303,N_16173,N_16487);
xnor U17304 (N_17304,N_16663,N_16293);
xnor U17305 (N_17305,N_16264,N_16443);
xnor U17306 (N_17306,N_16792,N_16101);
and U17307 (N_17307,N_16892,N_16277);
xor U17308 (N_17308,N_16093,N_16688);
nand U17309 (N_17309,N_16170,N_16748);
nor U17310 (N_17310,N_16666,N_16600);
nand U17311 (N_17311,N_16108,N_16910);
xnor U17312 (N_17312,N_16021,N_16265);
nand U17313 (N_17313,N_16412,N_16567);
nor U17314 (N_17314,N_16672,N_16447);
or U17315 (N_17315,N_16741,N_16271);
and U17316 (N_17316,N_16160,N_16103);
and U17317 (N_17317,N_16577,N_16077);
or U17318 (N_17318,N_16329,N_16197);
xnor U17319 (N_17319,N_16368,N_16955);
and U17320 (N_17320,N_16334,N_16904);
nor U17321 (N_17321,N_16767,N_16796);
xor U17322 (N_17322,N_16494,N_16521);
or U17323 (N_17323,N_16466,N_16056);
xor U17324 (N_17324,N_16211,N_16909);
nand U17325 (N_17325,N_16730,N_16064);
and U17326 (N_17326,N_16261,N_16862);
nand U17327 (N_17327,N_16433,N_16813);
nor U17328 (N_17328,N_16010,N_16294);
nor U17329 (N_17329,N_16526,N_16090);
and U17330 (N_17330,N_16185,N_16473);
nor U17331 (N_17331,N_16905,N_16963);
and U17332 (N_17332,N_16320,N_16773);
or U17333 (N_17333,N_16613,N_16615);
xor U17334 (N_17334,N_16238,N_16456);
nand U17335 (N_17335,N_16167,N_16042);
nor U17336 (N_17336,N_16361,N_16603);
or U17337 (N_17337,N_16373,N_16949);
and U17338 (N_17338,N_16890,N_16951);
or U17339 (N_17339,N_16158,N_16162);
nand U17340 (N_17340,N_16721,N_16325);
or U17341 (N_17341,N_16702,N_16345);
nand U17342 (N_17342,N_16207,N_16400);
nor U17343 (N_17343,N_16369,N_16068);
nand U17344 (N_17344,N_16478,N_16039);
nor U17345 (N_17345,N_16649,N_16316);
and U17346 (N_17346,N_16793,N_16481);
or U17347 (N_17347,N_16102,N_16845);
or U17348 (N_17348,N_16983,N_16803);
nor U17349 (N_17349,N_16821,N_16061);
or U17350 (N_17350,N_16339,N_16046);
xor U17351 (N_17351,N_16562,N_16650);
or U17352 (N_17352,N_16468,N_16704);
nand U17353 (N_17353,N_16498,N_16791);
nand U17354 (N_17354,N_16079,N_16427);
nand U17355 (N_17355,N_16036,N_16388);
or U17356 (N_17356,N_16113,N_16727);
and U17357 (N_17357,N_16518,N_16245);
or U17358 (N_17358,N_16474,N_16988);
xnor U17359 (N_17359,N_16029,N_16798);
xor U17360 (N_17360,N_16726,N_16829);
nand U17361 (N_17361,N_16174,N_16406);
and U17362 (N_17362,N_16013,N_16165);
nor U17363 (N_17363,N_16509,N_16689);
nor U17364 (N_17364,N_16797,N_16805);
nor U17365 (N_17365,N_16394,N_16735);
and U17366 (N_17366,N_16948,N_16356);
xor U17367 (N_17367,N_16318,N_16359);
and U17368 (N_17368,N_16868,N_16587);
and U17369 (N_17369,N_16132,N_16953);
or U17370 (N_17370,N_16038,N_16576);
xnor U17371 (N_17371,N_16699,N_16844);
and U17372 (N_17372,N_16978,N_16889);
nor U17373 (N_17373,N_16860,N_16074);
and U17374 (N_17374,N_16523,N_16028);
and U17375 (N_17375,N_16157,N_16811);
or U17376 (N_17376,N_16902,N_16442);
xnor U17377 (N_17377,N_16881,N_16545);
xor U17378 (N_17378,N_16653,N_16569);
nor U17379 (N_17379,N_16553,N_16907);
nor U17380 (N_17380,N_16035,N_16091);
nor U17381 (N_17381,N_16795,N_16467);
and U17382 (N_17382,N_16511,N_16592);
nand U17383 (N_17383,N_16175,N_16776);
or U17384 (N_17384,N_16323,N_16050);
or U17385 (N_17385,N_16172,N_16725);
and U17386 (N_17386,N_16464,N_16654);
nor U17387 (N_17387,N_16599,N_16217);
or U17388 (N_17388,N_16194,N_16247);
and U17389 (N_17389,N_16437,N_16861);
or U17390 (N_17390,N_16401,N_16794);
nand U17391 (N_17391,N_16127,N_16399);
nand U17392 (N_17392,N_16308,N_16984);
nand U17393 (N_17393,N_16051,N_16761);
xnor U17394 (N_17394,N_16121,N_16755);
and U17395 (N_17395,N_16971,N_16363);
xor U17396 (N_17396,N_16047,N_16985);
xor U17397 (N_17397,N_16004,N_16785);
nand U17398 (N_17398,N_16624,N_16054);
or U17399 (N_17399,N_16809,N_16639);
nand U17400 (N_17400,N_16431,N_16163);
nand U17401 (N_17401,N_16864,N_16084);
and U17402 (N_17402,N_16525,N_16122);
nor U17403 (N_17403,N_16582,N_16994);
xor U17404 (N_17404,N_16840,N_16883);
nand U17405 (N_17405,N_16940,N_16665);
nand U17406 (N_17406,N_16007,N_16327);
and U17407 (N_17407,N_16181,N_16372);
or U17408 (N_17408,N_16729,N_16488);
nand U17409 (N_17409,N_16635,N_16159);
and U17410 (N_17410,N_16621,N_16997);
and U17411 (N_17411,N_16147,N_16340);
or U17412 (N_17412,N_16700,N_16235);
or U17413 (N_17413,N_16922,N_16465);
and U17414 (N_17414,N_16818,N_16993);
and U17415 (N_17415,N_16109,N_16874);
xor U17416 (N_17416,N_16667,N_16204);
or U17417 (N_17417,N_16438,N_16817);
and U17418 (N_17418,N_16403,N_16529);
nor U17419 (N_17419,N_16405,N_16305);
or U17420 (N_17420,N_16858,N_16516);
nor U17421 (N_17421,N_16011,N_16096);
nand U17422 (N_17422,N_16182,N_16455);
nor U17423 (N_17423,N_16739,N_16536);
and U17424 (N_17424,N_16566,N_16231);
or U17425 (N_17425,N_16901,N_16939);
nand U17426 (N_17426,N_16135,N_16030);
nor U17427 (N_17427,N_16499,N_16626);
nor U17428 (N_17428,N_16220,N_16834);
xor U17429 (N_17429,N_16409,N_16670);
xor U17430 (N_17430,N_16111,N_16723);
or U17431 (N_17431,N_16778,N_16115);
xor U17432 (N_17432,N_16731,N_16453);
nor U17433 (N_17433,N_16208,N_16999);
nor U17434 (N_17434,N_16336,N_16138);
nor U17435 (N_17435,N_16131,N_16151);
nand U17436 (N_17436,N_16617,N_16214);
xor U17437 (N_17437,N_16900,N_16332);
or U17438 (N_17438,N_16460,N_16192);
nand U17439 (N_17439,N_16485,N_16097);
xnor U17440 (N_17440,N_16052,N_16133);
and U17441 (N_17441,N_16166,N_16354);
and U17442 (N_17442,N_16616,N_16315);
xor U17443 (N_17443,N_16637,N_16191);
nand U17444 (N_17444,N_16931,N_16430);
and U17445 (N_17445,N_16557,N_16129);
and U17446 (N_17446,N_16808,N_16816);
and U17447 (N_17447,N_16397,N_16787);
or U17448 (N_17448,N_16974,N_16053);
nor U17449 (N_17449,N_16819,N_16869);
nand U17450 (N_17450,N_16867,N_16434);
and U17451 (N_17451,N_16732,N_16161);
or U17452 (N_17452,N_16676,N_16596);
xnor U17453 (N_17453,N_16806,N_16075);
nor U17454 (N_17454,N_16952,N_16945);
nand U17455 (N_17455,N_16510,N_16459);
nor U17456 (N_17456,N_16788,N_16733);
or U17457 (N_17457,N_16559,N_16912);
and U17458 (N_17458,N_16969,N_16899);
and U17459 (N_17459,N_16069,N_16026);
nand U17460 (N_17460,N_16307,N_16873);
and U17461 (N_17461,N_16623,N_16267);
or U17462 (N_17462,N_16593,N_16344);
or U17463 (N_17463,N_16040,N_16924);
nor U17464 (N_17464,N_16164,N_16112);
nor U17465 (N_17465,N_16387,N_16279);
xnor U17466 (N_17466,N_16625,N_16928);
or U17467 (N_17467,N_16432,N_16482);
nor U17468 (N_17468,N_16830,N_16012);
nor U17469 (N_17469,N_16237,N_16920);
and U17470 (N_17470,N_16502,N_16677);
xor U17471 (N_17471,N_16657,N_16083);
nand U17472 (N_17472,N_16871,N_16371);
nand U17473 (N_17473,N_16343,N_16713);
nand U17474 (N_17474,N_16496,N_16178);
nor U17475 (N_17475,N_16128,N_16695);
nand U17476 (N_17476,N_16176,N_16281);
xnor U17477 (N_17477,N_16210,N_16202);
or U17478 (N_17478,N_16310,N_16196);
nand U17479 (N_17479,N_16843,N_16392);
nor U17480 (N_17480,N_16604,N_16683);
or U17481 (N_17481,N_16374,N_16764);
or U17482 (N_17482,N_16541,N_16259);
and U17483 (N_17483,N_16156,N_16512);
and U17484 (N_17484,N_16754,N_16299);
and U17485 (N_17485,N_16886,N_16534);
and U17486 (N_17486,N_16240,N_16556);
or U17487 (N_17487,N_16335,N_16770);
nor U17488 (N_17488,N_16934,N_16360);
nand U17489 (N_17489,N_16959,N_16973);
and U17490 (N_17490,N_16338,N_16395);
and U17491 (N_17491,N_16055,N_16691);
nor U17492 (N_17492,N_16366,N_16717);
nand U17493 (N_17493,N_16484,N_16095);
nand U17494 (N_17494,N_16640,N_16958);
xor U17495 (N_17495,N_16020,N_16298);
nor U17496 (N_17496,N_16152,N_16440);
and U17497 (N_17497,N_16006,N_16853);
nor U17498 (N_17498,N_16836,N_16519);
nand U17499 (N_17499,N_16644,N_16612);
or U17500 (N_17500,N_16428,N_16341);
nand U17501 (N_17501,N_16755,N_16514);
nand U17502 (N_17502,N_16023,N_16694);
or U17503 (N_17503,N_16075,N_16590);
xnor U17504 (N_17504,N_16647,N_16062);
xnor U17505 (N_17505,N_16992,N_16237);
or U17506 (N_17506,N_16102,N_16175);
nor U17507 (N_17507,N_16057,N_16013);
nand U17508 (N_17508,N_16422,N_16854);
xor U17509 (N_17509,N_16799,N_16492);
or U17510 (N_17510,N_16831,N_16518);
nor U17511 (N_17511,N_16829,N_16595);
xnor U17512 (N_17512,N_16064,N_16243);
nand U17513 (N_17513,N_16023,N_16263);
nand U17514 (N_17514,N_16585,N_16018);
or U17515 (N_17515,N_16920,N_16317);
and U17516 (N_17516,N_16771,N_16124);
nor U17517 (N_17517,N_16767,N_16779);
or U17518 (N_17518,N_16964,N_16580);
and U17519 (N_17519,N_16771,N_16212);
nand U17520 (N_17520,N_16297,N_16359);
xnor U17521 (N_17521,N_16274,N_16233);
and U17522 (N_17522,N_16175,N_16146);
xor U17523 (N_17523,N_16676,N_16114);
or U17524 (N_17524,N_16957,N_16803);
and U17525 (N_17525,N_16439,N_16390);
and U17526 (N_17526,N_16302,N_16976);
xor U17527 (N_17527,N_16715,N_16565);
nor U17528 (N_17528,N_16895,N_16216);
xor U17529 (N_17529,N_16390,N_16000);
nand U17530 (N_17530,N_16076,N_16570);
and U17531 (N_17531,N_16278,N_16471);
or U17532 (N_17532,N_16919,N_16183);
or U17533 (N_17533,N_16021,N_16342);
or U17534 (N_17534,N_16013,N_16467);
xor U17535 (N_17535,N_16616,N_16041);
xor U17536 (N_17536,N_16196,N_16823);
nor U17537 (N_17537,N_16369,N_16485);
or U17538 (N_17538,N_16119,N_16570);
nand U17539 (N_17539,N_16682,N_16872);
nand U17540 (N_17540,N_16512,N_16147);
or U17541 (N_17541,N_16462,N_16888);
or U17542 (N_17542,N_16241,N_16282);
nand U17543 (N_17543,N_16424,N_16174);
xor U17544 (N_17544,N_16598,N_16480);
and U17545 (N_17545,N_16783,N_16916);
xor U17546 (N_17546,N_16443,N_16483);
nand U17547 (N_17547,N_16763,N_16106);
and U17548 (N_17548,N_16614,N_16891);
and U17549 (N_17549,N_16987,N_16894);
xor U17550 (N_17550,N_16759,N_16574);
and U17551 (N_17551,N_16365,N_16347);
nand U17552 (N_17552,N_16539,N_16982);
nor U17553 (N_17553,N_16461,N_16840);
nand U17554 (N_17554,N_16457,N_16487);
xor U17555 (N_17555,N_16035,N_16777);
or U17556 (N_17556,N_16513,N_16394);
or U17557 (N_17557,N_16531,N_16451);
xnor U17558 (N_17558,N_16523,N_16463);
or U17559 (N_17559,N_16210,N_16287);
xnor U17560 (N_17560,N_16649,N_16880);
nor U17561 (N_17561,N_16177,N_16484);
or U17562 (N_17562,N_16061,N_16057);
nand U17563 (N_17563,N_16649,N_16074);
or U17564 (N_17564,N_16441,N_16421);
nor U17565 (N_17565,N_16549,N_16251);
nand U17566 (N_17566,N_16706,N_16294);
nand U17567 (N_17567,N_16153,N_16881);
and U17568 (N_17568,N_16620,N_16829);
and U17569 (N_17569,N_16634,N_16868);
and U17570 (N_17570,N_16091,N_16655);
nor U17571 (N_17571,N_16294,N_16053);
nor U17572 (N_17572,N_16742,N_16173);
and U17573 (N_17573,N_16028,N_16852);
or U17574 (N_17574,N_16158,N_16611);
and U17575 (N_17575,N_16086,N_16409);
or U17576 (N_17576,N_16404,N_16506);
xnor U17577 (N_17577,N_16929,N_16078);
or U17578 (N_17578,N_16166,N_16668);
and U17579 (N_17579,N_16663,N_16491);
xor U17580 (N_17580,N_16926,N_16670);
nor U17581 (N_17581,N_16400,N_16861);
and U17582 (N_17582,N_16796,N_16597);
and U17583 (N_17583,N_16684,N_16911);
and U17584 (N_17584,N_16002,N_16028);
xor U17585 (N_17585,N_16781,N_16187);
and U17586 (N_17586,N_16208,N_16357);
and U17587 (N_17587,N_16971,N_16895);
and U17588 (N_17588,N_16226,N_16551);
xor U17589 (N_17589,N_16695,N_16072);
nand U17590 (N_17590,N_16597,N_16572);
nand U17591 (N_17591,N_16587,N_16531);
xnor U17592 (N_17592,N_16473,N_16595);
nor U17593 (N_17593,N_16686,N_16662);
nand U17594 (N_17594,N_16331,N_16471);
nor U17595 (N_17595,N_16804,N_16319);
xnor U17596 (N_17596,N_16803,N_16900);
xnor U17597 (N_17597,N_16498,N_16229);
or U17598 (N_17598,N_16391,N_16061);
and U17599 (N_17599,N_16913,N_16939);
and U17600 (N_17600,N_16654,N_16829);
or U17601 (N_17601,N_16995,N_16137);
and U17602 (N_17602,N_16483,N_16681);
nand U17603 (N_17603,N_16011,N_16727);
and U17604 (N_17604,N_16784,N_16885);
nand U17605 (N_17605,N_16876,N_16648);
xnor U17606 (N_17606,N_16492,N_16771);
nor U17607 (N_17607,N_16637,N_16615);
and U17608 (N_17608,N_16255,N_16428);
and U17609 (N_17609,N_16021,N_16006);
and U17610 (N_17610,N_16186,N_16146);
or U17611 (N_17611,N_16081,N_16257);
xor U17612 (N_17612,N_16328,N_16649);
nor U17613 (N_17613,N_16351,N_16126);
xor U17614 (N_17614,N_16060,N_16698);
or U17615 (N_17615,N_16276,N_16060);
and U17616 (N_17616,N_16569,N_16217);
nand U17617 (N_17617,N_16071,N_16089);
and U17618 (N_17618,N_16574,N_16842);
xor U17619 (N_17619,N_16391,N_16277);
and U17620 (N_17620,N_16607,N_16358);
nand U17621 (N_17621,N_16517,N_16229);
xor U17622 (N_17622,N_16230,N_16199);
and U17623 (N_17623,N_16201,N_16936);
or U17624 (N_17624,N_16495,N_16170);
nor U17625 (N_17625,N_16578,N_16983);
xnor U17626 (N_17626,N_16158,N_16680);
xor U17627 (N_17627,N_16906,N_16090);
nor U17628 (N_17628,N_16908,N_16471);
and U17629 (N_17629,N_16034,N_16047);
nor U17630 (N_17630,N_16018,N_16462);
xnor U17631 (N_17631,N_16760,N_16403);
nand U17632 (N_17632,N_16257,N_16878);
nand U17633 (N_17633,N_16576,N_16154);
and U17634 (N_17634,N_16811,N_16533);
nand U17635 (N_17635,N_16514,N_16716);
and U17636 (N_17636,N_16399,N_16975);
nor U17637 (N_17637,N_16261,N_16762);
nor U17638 (N_17638,N_16494,N_16074);
nor U17639 (N_17639,N_16547,N_16907);
nor U17640 (N_17640,N_16050,N_16930);
xnor U17641 (N_17641,N_16060,N_16530);
or U17642 (N_17642,N_16375,N_16473);
or U17643 (N_17643,N_16053,N_16345);
or U17644 (N_17644,N_16577,N_16269);
nor U17645 (N_17645,N_16575,N_16541);
nor U17646 (N_17646,N_16426,N_16377);
and U17647 (N_17647,N_16659,N_16784);
or U17648 (N_17648,N_16767,N_16565);
nand U17649 (N_17649,N_16449,N_16941);
xnor U17650 (N_17650,N_16319,N_16953);
or U17651 (N_17651,N_16161,N_16692);
and U17652 (N_17652,N_16509,N_16467);
or U17653 (N_17653,N_16579,N_16303);
xor U17654 (N_17654,N_16841,N_16707);
nand U17655 (N_17655,N_16666,N_16236);
nor U17656 (N_17656,N_16765,N_16925);
nand U17657 (N_17657,N_16626,N_16397);
or U17658 (N_17658,N_16142,N_16998);
and U17659 (N_17659,N_16213,N_16498);
xor U17660 (N_17660,N_16462,N_16905);
nor U17661 (N_17661,N_16604,N_16626);
xnor U17662 (N_17662,N_16957,N_16602);
nor U17663 (N_17663,N_16903,N_16624);
xor U17664 (N_17664,N_16985,N_16613);
and U17665 (N_17665,N_16487,N_16354);
nand U17666 (N_17666,N_16744,N_16036);
or U17667 (N_17667,N_16644,N_16795);
or U17668 (N_17668,N_16764,N_16517);
nor U17669 (N_17669,N_16518,N_16406);
and U17670 (N_17670,N_16205,N_16749);
xnor U17671 (N_17671,N_16770,N_16652);
nor U17672 (N_17672,N_16461,N_16897);
xnor U17673 (N_17673,N_16869,N_16180);
nor U17674 (N_17674,N_16567,N_16310);
nor U17675 (N_17675,N_16348,N_16881);
nand U17676 (N_17676,N_16866,N_16220);
nand U17677 (N_17677,N_16810,N_16919);
nand U17678 (N_17678,N_16683,N_16759);
nor U17679 (N_17679,N_16389,N_16906);
xor U17680 (N_17680,N_16666,N_16886);
or U17681 (N_17681,N_16454,N_16283);
nand U17682 (N_17682,N_16752,N_16394);
and U17683 (N_17683,N_16418,N_16807);
xnor U17684 (N_17684,N_16368,N_16995);
and U17685 (N_17685,N_16069,N_16441);
xnor U17686 (N_17686,N_16386,N_16245);
xnor U17687 (N_17687,N_16047,N_16632);
and U17688 (N_17688,N_16989,N_16786);
and U17689 (N_17689,N_16105,N_16028);
nor U17690 (N_17690,N_16746,N_16977);
nor U17691 (N_17691,N_16839,N_16066);
xor U17692 (N_17692,N_16162,N_16783);
nor U17693 (N_17693,N_16892,N_16646);
nand U17694 (N_17694,N_16726,N_16661);
nand U17695 (N_17695,N_16474,N_16333);
and U17696 (N_17696,N_16692,N_16136);
or U17697 (N_17697,N_16177,N_16941);
nand U17698 (N_17698,N_16878,N_16831);
nand U17699 (N_17699,N_16433,N_16238);
and U17700 (N_17700,N_16425,N_16516);
nor U17701 (N_17701,N_16668,N_16862);
nand U17702 (N_17702,N_16191,N_16616);
and U17703 (N_17703,N_16422,N_16279);
or U17704 (N_17704,N_16533,N_16924);
nor U17705 (N_17705,N_16493,N_16797);
nand U17706 (N_17706,N_16659,N_16113);
nand U17707 (N_17707,N_16619,N_16837);
or U17708 (N_17708,N_16897,N_16135);
nand U17709 (N_17709,N_16938,N_16120);
or U17710 (N_17710,N_16883,N_16533);
nor U17711 (N_17711,N_16077,N_16062);
or U17712 (N_17712,N_16927,N_16297);
xor U17713 (N_17713,N_16022,N_16910);
xor U17714 (N_17714,N_16167,N_16137);
or U17715 (N_17715,N_16633,N_16168);
xor U17716 (N_17716,N_16802,N_16420);
nor U17717 (N_17717,N_16806,N_16780);
or U17718 (N_17718,N_16342,N_16158);
xnor U17719 (N_17719,N_16722,N_16937);
and U17720 (N_17720,N_16143,N_16592);
and U17721 (N_17721,N_16279,N_16893);
and U17722 (N_17722,N_16535,N_16191);
xnor U17723 (N_17723,N_16667,N_16784);
or U17724 (N_17724,N_16057,N_16610);
or U17725 (N_17725,N_16951,N_16872);
nand U17726 (N_17726,N_16271,N_16697);
nand U17727 (N_17727,N_16528,N_16908);
nand U17728 (N_17728,N_16746,N_16164);
nand U17729 (N_17729,N_16075,N_16869);
nand U17730 (N_17730,N_16985,N_16519);
nor U17731 (N_17731,N_16318,N_16125);
nand U17732 (N_17732,N_16721,N_16066);
and U17733 (N_17733,N_16236,N_16080);
nand U17734 (N_17734,N_16075,N_16256);
nor U17735 (N_17735,N_16083,N_16241);
nand U17736 (N_17736,N_16159,N_16417);
or U17737 (N_17737,N_16221,N_16688);
and U17738 (N_17738,N_16529,N_16100);
or U17739 (N_17739,N_16457,N_16361);
nor U17740 (N_17740,N_16128,N_16117);
nor U17741 (N_17741,N_16277,N_16255);
or U17742 (N_17742,N_16284,N_16780);
nand U17743 (N_17743,N_16911,N_16375);
nor U17744 (N_17744,N_16674,N_16397);
xor U17745 (N_17745,N_16407,N_16375);
nand U17746 (N_17746,N_16477,N_16181);
nor U17747 (N_17747,N_16903,N_16345);
nand U17748 (N_17748,N_16600,N_16083);
xnor U17749 (N_17749,N_16424,N_16385);
nor U17750 (N_17750,N_16126,N_16189);
xor U17751 (N_17751,N_16218,N_16773);
nor U17752 (N_17752,N_16821,N_16847);
xor U17753 (N_17753,N_16376,N_16676);
nand U17754 (N_17754,N_16402,N_16938);
and U17755 (N_17755,N_16860,N_16276);
nand U17756 (N_17756,N_16393,N_16831);
nor U17757 (N_17757,N_16252,N_16400);
nand U17758 (N_17758,N_16534,N_16452);
nor U17759 (N_17759,N_16395,N_16842);
nand U17760 (N_17760,N_16094,N_16421);
xor U17761 (N_17761,N_16239,N_16746);
and U17762 (N_17762,N_16742,N_16032);
nand U17763 (N_17763,N_16555,N_16185);
xor U17764 (N_17764,N_16960,N_16381);
xor U17765 (N_17765,N_16195,N_16391);
nor U17766 (N_17766,N_16996,N_16806);
nor U17767 (N_17767,N_16506,N_16346);
xor U17768 (N_17768,N_16926,N_16752);
xor U17769 (N_17769,N_16502,N_16661);
xnor U17770 (N_17770,N_16779,N_16530);
and U17771 (N_17771,N_16156,N_16873);
nand U17772 (N_17772,N_16815,N_16997);
xor U17773 (N_17773,N_16071,N_16974);
nand U17774 (N_17774,N_16429,N_16807);
and U17775 (N_17775,N_16033,N_16520);
xor U17776 (N_17776,N_16932,N_16629);
nand U17777 (N_17777,N_16386,N_16870);
nor U17778 (N_17778,N_16473,N_16502);
xor U17779 (N_17779,N_16681,N_16138);
or U17780 (N_17780,N_16854,N_16416);
or U17781 (N_17781,N_16169,N_16120);
and U17782 (N_17782,N_16921,N_16772);
nand U17783 (N_17783,N_16226,N_16110);
nor U17784 (N_17784,N_16834,N_16405);
nor U17785 (N_17785,N_16527,N_16432);
and U17786 (N_17786,N_16503,N_16148);
xnor U17787 (N_17787,N_16795,N_16085);
and U17788 (N_17788,N_16411,N_16260);
nor U17789 (N_17789,N_16431,N_16208);
nand U17790 (N_17790,N_16583,N_16382);
and U17791 (N_17791,N_16501,N_16343);
nor U17792 (N_17792,N_16994,N_16290);
nor U17793 (N_17793,N_16494,N_16627);
or U17794 (N_17794,N_16678,N_16463);
xnor U17795 (N_17795,N_16001,N_16712);
and U17796 (N_17796,N_16574,N_16472);
nor U17797 (N_17797,N_16303,N_16175);
nand U17798 (N_17798,N_16793,N_16064);
nor U17799 (N_17799,N_16111,N_16285);
xor U17800 (N_17800,N_16653,N_16990);
and U17801 (N_17801,N_16741,N_16013);
nor U17802 (N_17802,N_16501,N_16035);
nand U17803 (N_17803,N_16252,N_16305);
nand U17804 (N_17804,N_16915,N_16461);
and U17805 (N_17805,N_16709,N_16615);
and U17806 (N_17806,N_16747,N_16680);
xnor U17807 (N_17807,N_16111,N_16953);
nor U17808 (N_17808,N_16791,N_16894);
and U17809 (N_17809,N_16024,N_16043);
nor U17810 (N_17810,N_16340,N_16139);
and U17811 (N_17811,N_16720,N_16449);
and U17812 (N_17812,N_16269,N_16674);
and U17813 (N_17813,N_16876,N_16866);
nand U17814 (N_17814,N_16426,N_16280);
nor U17815 (N_17815,N_16482,N_16096);
xnor U17816 (N_17816,N_16004,N_16505);
or U17817 (N_17817,N_16653,N_16794);
nor U17818 (N_17818,N_16729,N_16497);
nand U17819 (N_17819,N_16007,N_16576);
nand U17820 (N_17820,N_16719,N_16387);
xnor U17821 (N_17821,N_16764,N_16285);
xor U17822 (N_17822,N_16107,N_16752);
and U17823 (N_17823,N_16133,N_16159);
and U17824 (N_17824,N_16688,N_16922);
and U17825 (N_17825,N_16409,N_16609);
nand U17826 (N_17826,N_16634,N_16606);
nand U17827 (N_17827,N_16106,N_16755);
and U17828 (N_17828,N_16027,N_16304);
xnor U17829 (N_17829,N_16407,N_16109);
nand U17830 (N_17830,N_16210,N_16007);
or U17831 (N_17831,N_16125,N_16923);
or U17832 (N_17832,N_16378,N_16968);
and U17833 (N_17833,N_16035,N_16008);
nand U17834 (N_17834,N_16833,N_16355);
or U17835 (N_17835,N_16621,N_16771);
nor U17836 (N_17836,N_16594,N_16528);
nand U17837 (N_17837,N_16552,N_16416);
nor U17838 (N_17838,N_16383,N_16940);
nand U17839 (N_17839,N_16157,N_16609);
xor U17840 (N_17840,N_16136,N_16534);
and U17841 (N_17841,N_16649,N_16776);
nand U17842 (N_17842,N_16619,N_16354);
xor U17843 (N_17843,N_16547,N_16552);
xnor U17844 (N_17844,N_16021,N_16272);
xor U17845 (N_17845,N_16089,N_16661);
xor U17846 (N_17846,N_16621,N_16159);
and U17847 (N_17847,N_16142,N_16907);
and U17848 (N_17848,N_16844,N_16632);
nor U17849 (N_17849,N_16558,N_16770);
xnor U17850 (N_17850,N_16432,N_16854);
nor U17851 (N_17851,N_16137,N_16904);
nand U17852 (N_17852,N_16609,N_16830);
nand U17853 (N_17853,N_16070,N_16117);
nand U17854 (N_17854,N_16217,N_16278);
nor U17855 (N_17855,N_16354,N_16879);
nand U17856 (N_17856,N_16601,N_16489);
nor U17857 (N_17857,N_16059,N_16904);
nand U17858 (N_17858,N_16489,N_16568);
and U17859 (N_17859,N_16385,N_16313);
and U17860 (N_17860,N_16383,N_16793);
xnor U17861 (N_17861,N_16209,N_16203);
xor U17862 (N_17862,N_16089,N_16009);
or U17863 (N_17863,N_16029,N_16680);
nand U17864 (N_17864,N_16904,N_16497);
or U17865 (N_17865,N_16453,N_16857);
or U17866 (N_17866,N_16502,N_16015);
nor U17867 (N_17867,N_16528,N_16667);
nand U17868 (N_17868,N_16547,N_16665);
or U17869 (N_17869,N_16915,N_16313);
and U17870 (N_17870,N_16729,N_16457);
or U17871 (N_17871,N_16140,N_16531);
nor U17872 (N_17872,N_16690,N_16492);
and U17873 (N_17873,N_16117,N_16353);
xor U17874 (N_17874,N_16802,N_16479);
nor U17875 (N_17875,N_16258,N_16808);
nor U17876 (N_17876,N_16017,N_16862);
nand U17877 (N_17877,N_16905,N_16127);
nor U17878 (N_17878,N_16871,N_16564);
or U17879 (N_17879,N_16522,N_16560);
or U17880 (N_17880,N_16000,N_16005);
nand U17881 (N_17881,N_16985,N_16661);
and U17882 (N_17882,N_16131,N_16092);
nand U17883 (N_17883,N_16275,N_16497);
nor U17884 (N_17884,N_16333,N_16353);
nand U17885 (N_17885,N_16034,N_16027);
nor U17886 (N_17886,N_16519,N_16049);
nand U17887 (N_17887,N_16749,N_16403);
nand U17888 (N_17888,N_16283,N_16200);
xor U17889 (N_17889,N_16834,N_16223);
xor U17890 (N_17890,N_16519,N_16110);
nand U17891 (N_17891,N_16857,N_16634);
or U17892 (N_17892,N_16047,N_16439);
or U17893 (N_17893,N_16964,N_16997);
and U17894 (N_17894,N_16995,N_16005);
xnor U17895 (N_17895,N_16407,N_16461);
and U17896 (N_17896,N_16753,N_16147);
xor U17897 (N_17897,N_16443,N_16144);
nor U17898 (N_17898,N_16877,N_16726);
or U17899 (N_17899,N_16770,N_16786);
xor U17900 (N_17900,N_16826,N_16102);
and U17901 (N_17901,N_16890,N_16025);
xnor U17902 (N_17902,N_16061,N_16200);
or U17903 (N_17903,N_16735,N_16201);
nand U17904 (N_17904,N_16810,N_16857);
xnor U17905 (N_17905,N_16546,N_16192);
and U17906 (N_17906,N_16354,N_16362);
and U17907 (N_17907,N_16224,N_16329);
xnor U17908 (N_17908,N_16992,N_16818);
or U17909 (N_17909,N_16204,N_16171);
or U17910 (N_17910,N_16763,N_16079);
xnor U17911 (N_17911,N_16824,N_16556);
nand U17912 (N_17912,N_16726,N_16711);
and U17913 (N_17913,N_16708,N_16943);
and U17914 (N_17914,N_16946,N_16807);
and U17915 (N_17915,N_16031,N_16047);
and U17916 (N_17916,N_16193,N_16836);
and U17917 (N_17917,N_16861,N_16058);
and U17918 (N_17918,N_16269,N_16478);
nor U17919 (N_17919,N_16970,N_16363);
or U17920 (N_17920,N_16076,N_16790);
or U17921 (N_17921,N_16861,N_16707);
and U17922 (N_17922,N_16183,N_16466);
xnor U17923 (N_17923,N_16710,N_16118);
nand U17924 (N_17924,N_16068,N_16373);
nand U17925 (N_17925,N_16925,N_16955);
and U17926 (N_17926,N_16003,N_16197);
xor U17927 (N_17927,N_16335,N_16766);
or U17928 (N_17928,N_16498,N_16345);
nor U17929 (N_17929,N_16793,N_16641);
nor U17930 (N_17930,N_16975,N_16443);
nor U17931 (N_17931,N_16686,N_16650);
xor U17932 (N_17932,N_16307,N_16354);
nand U17933 (N_17933,N_16832,N_16470);
nand U17934 (N_17934,N_16561,N_16229);
or U17935 (N_17935,N_16304,N_16907);
and U17936 (N_17936,N_16026,N_16336);
xor U17937 (N_17937,N_16403,N_16813);
or U17938 (N_17938,N_16561,N_16440);
nor U17939 (N_17939,N_16733,N_16654);
and U17940 (N_17940,N_16201,N_16931);
nand U17941 (N_17941,N_16876,N_16242);
xor U17942 (N_17942,N_16581,N_16937);
xnor U17943 (N_17943,N_16760,N_16302);
or U17944 (N_17944,N_16693,N_16192);
nor U17945 (N_17945,N_16486,N_16955);
or U17946 (N_17946,N_16928,N_16122);
and U17947 (N_17947,N_16028,N_16315);
xor U17948 (N_17948,N_16710,N_16948);
xnor U17949 (N_17949,N_16324,N_16866);
nor U17950 (N_17950,N_16745,N_16955);
nand U17951 (N_17951,N_16232,N_16737);
or U17952 (N_17952,N_16870,N_16462);
or U17953 (N_17953,N_16416,N_16261);
nor U17954 (N_17954,N_16378,N_16408);
or U17955 (N_17955,N_16620,N_16821);
xor U17956 (N_17956,N_16633,N_16480);
xor U17957 (N_17957,N_16823,N_16505);
xor U17958 (N_17958,N_16048,N_16287);
nand U17959 (N_17959,N_16854,N_16985);
or U17960 (N_17960,N_16533,N_16808);
xor U17961 (N_17961,N_16246,N_16642);
nand U17962 (N_17962,N_16643,N_16076);
and U17963 (N_17963,N_16051,N_16714);
and U17964 (N_17964,N_16371,N_16533);
or U17965 (N_17965,N_16417,N_16782);
nor U17966 (N_17966,N_16696,N_16425);
nor U17967 (N_17967,N_16937,N_16552);
xor U17968 (N_17968,N_16468,N_16674);
xor U17969 (N_17969,N_16761,N_16415);
or U17970 (N_17970,N_16443,N_16197);
xnor U17971 (N_17971,N_16564,N_16491);
or U17972 (N_17972,N_16302,N_16502);
xor U17973 (N_17973,N_16170,N_16967);
and U17974 (N_17974,N_16740,N_16760);
xor U17975 (N_17975,N_16004,N_16070);
and U17976 (N_17976,N_16172,N_16600);
nand U17977 (N_17977,N_16247,N_16833);
nand U17978 (N_17978,N_16933,N_16729);
nand U17979 (N_17979,N_16956,N_16336);
or U17980 (N_17980,N_16803,N_16643);
xor U17981 (N_17981,N_16526,N_16889);
and U17982 (N_17982,N_16127,N_16559);
nor U17983 (N_17983,N_16252,N_16926);
xnor U17984 (N_17984,N_16714,N_16552);
and U17985 (N_17985,N_16332,N_16852);
and U17986 (N_17986,N_16266,N_16801);
nor U17987 (N_17987,N_16536,N_16838);
xnor U17988 (N_17988,N_16791,N_16708);
or U17989 (N_17989,N_16047,N_16132);
xnor U17990 (N_17990,N_16648,N_16246);
xnor U17991 (N_17991,N_16166,N_16682);
xor U17992 (N_17992,N_16448,N_16995);
nor U17993 (N_17993,N_16687,N_16239);
and U17994 (N_17994,N_16701,N_16012);
nand U17995 (N_17995,N_16206,N_16381);
nand U17996 (N_17996,N_16693,N_16763);
nand U17997 (N_17997,N_16016,N_16675);
or U17998 (N_17998,N_16608,N_16017);
and U17999 (N_17999,N_16554,N_16611);
nand U18000 (N_18000,N_17771,N_17626);
or U18001 (N_18001,N_17438,N_17558);
xor U18002 (N_18002,N_17876,N_17879);
nor U18003 (N_18003,N_17969,N_17726);
and U18004 (N_18004,N_17696,N_17490);
nor U18005 (N_18005,N_17515,N_17158);
nor U18006 (N_18006,N_17561,N_17605);
or U18007 (N_18007,N_17457,N_17367);
and U18008 (N_18008,N_17450,N_17947);
xnor U18009 (N_18009,N_17412,N_17674);
and U18010 (N_18010,N_17730,N_17034);
or U18011 (N_18011,N_17682,N_17645);
and U18012 (N_18012,N_17287,N_17404);
and U18013 (N_18013,N_17036,N_17664);
nand U18014 (N_18014,N_17456,N_17210);
or U18015 (N_18015,N_17591,N_17294);
nand U18016 (N_18016,N_17095,N_17628);
nand U18017 (N_18017,N_17209,N_17550);
xor U18018 (N_18018,N_17604,N_17942);
nand U18019 (N_18019,N_17927,N_17620);
xor U18020 (N_18020,N_17613,N_17756);
nand U18021 (N_18021,N_17476,N_17124);
nand U18022 (N_18022,N_17469,N_17688);
nand U18023 (N_18023,N_17974,N_17486);
and U18024 (N_18024,N_17607,N_17570);
xnor U18025 (N_18025,N_17168,N_17848);
xor U18026 (N_18026,N_17488,N_17527);
or U18027 (N_18027,N_17175,N_17243);
nor U18028 (N_18028,N_17845,N_17082);
nor U18029 (N_18029,N_17010,N_17694);
nand U18030 (N_18030,N_17171,N_17184);
nor U18031 (N_18031,N_17402,N_17325);
xnor U18032 (N_18032,N_17152,N_17827);
xor U18033 (N_18033,N_17295,N_17493);
nor U18034 (N_18034,N_17391,N_17874);
or U18035 (N_18035,N_17277,N_17377);
nand U18036 (N_18036,N_17719,N_17348);
xor U18037 (N_18037,N_17923,N_17500);
nand U18038 (N_18038,N_17100,N_17815);
or U18039 (N_18039,N_17729,N_17042);
nand U18040 (N_18040,N_17776,N_17761);
and U18041 (N_18041,N_17769,N_17569);
xor U18042 (N_18042,N_17275,N_17148);
nand U18043 (N_18043,N_17055,N_17349);
xor U18044 (N_18044,N_17429,N_17700);
and U18045 (N_18045,N_17526,N_17016);
and U18046 (N_18046,N_17079,N_17366);
nor U18047 (N_18047,N_17847,N_17931);
xor U18048 (N_18048,N_17663,N_17985);
xnor U18049 (N_18049,N_17229,N_17618);
or U18050 (N_18050,N_17333,N_17544);
nand U18051 (N_18051,N_17266,N_17763);
nor U18052 (N_18052,N_17522,N_17291);
or U18053 (N_18053,N_17115,N_17997);
and U18054 (N_18054,N_17331,N_17679);
or U18055 (N_18055,N_17789,N_17279);
and U18056 (N_18056,N_17453,N_17482);
and U18057 (N_18057,N_17512,N_17023);
and U18058 (N_18058,N_17015,N_17501);
and U18059 (N_18059,N_17934,N_17314);
nand U18060 (N_18060,N_17956,N_17987);
xnor U18061 (N_18061,N_17669,N_17917);
and U18062 (N_18062,N_17706,N_17345);
nor U18063 (N_18063,N_17661,N_17868);
nor U18064 (N_18064,N_17068,N_17166);
nor U18065 (N_18065,N_17650,N_17720);
nand U18066 (N_18066,N_17810,N_17360);
xnor U18067 (N_18067,N_17610,N_17508);
or U18068 (N_18068,N_17919,N_17714);
or U18069 (N_18069,N_17248,N_17414);
nor U18070 (N_18070,N_17255,N_17154);
nor U18071 (N_18071,N_17315,N_17887);
or U18072 (N_18072,N_17624,N_17652);
and U18073 (N_18073,N_17098,N_17216);
and U18074 (N_18074,N_17920,N_17766);
and U18075 (N_18075,N_17410,N_17841);
and U18076 (N_18076,N_17589,N_17466);
and U18077 (N_18077,N_17894,N_17641);
or U18078 (N_18078,N_17346,N_17639);
or U18079 (N_18079,N_17788,N_17268);
nor U18080 (N_18080,N_17625,N_17926);
and U18081 (N_18081,N_17568,N_17063);
or U18082 (N_18082,N_17698,N_17838);
nor U18083 (N_18083,N_17594,N_17914);
and U18084 (N_18084,N_17566,N_17191);
xnor U18085 (N_18085,N_17257,N_17787);
or U18086 (N_18086,N_17986,N_17276);
and U18087 (N_18087,N_17244,N_17973);
and U18088 (N_18088,N_17783,N_17470);
xor U18089 (N_18089,N_17867,N_17718);
and U18090 (N_18090,N_17830,N_17608);
xnor U18091 (N_18091,N_17144,N_17379);
nand U18092 (N_18092,N_17693,N_17744);
and U18093 (N_18093,N_17891,N_17992);
nor U18094 (N_18094,N_17064,N_17433);
or U18095 (N_18095,N_17617,N_17520);
or U18096 (N_18096,N_17008,N_17965);
and U18097 (N_18097,N_17282,N_17924);
nand U18098 (N_18098,N_17517,N_17001);
nor U18099 (N_18099,N_17196,N_17937);
xnor U18100 (N_18100,N_17150,N_17288);
or U18101 (N_18101,N_17407,N_17996);
xor U18102 (N_18102,N_17472,N_17235);
xor U18103 (N_18103,N_17668,N_17409);
nor U18104 (N_18104,N_17381,N_17609);
and U18105 (N_18105,N_17518,N_17962);
nand U18106 (N_18106,N_17822,N_17577);
nand U18107 (N_18107,N_17363,N_17935);
xnor U18108 (N_18108,N_17084,N_17860);
nand U18109 (N_18109,N_17910,N_17913);
nor U18110 (N_18110,N_17317,N_17305);
xor U18111 (N_18111,N_17840,N_17939);
nand U18112 (N_18112,N_17051,N_17957);
xor U18113 (N_18113,N_17820,N_17012);
xnor U18114 (N_18114,N_17811,N_17353);
nor U18115 (N_18115,N_17795,N_17821);
and U18116 (N_18116,N_17362,N_17826);
and U18117 (N_18117,N_17292,N_17181);
or U18118 (N_18118,N_17227,N_17564);
or U18119 (N_18119,N_17125,N_17989);
xnor U18120 (N_18120,N_17030,N_17339);
nor U18121 (N_18121,N_17651,N_17963);
or U18122 (N_18122,N_17621,N_17280);
nand U18123 (N_18123,N_17185,N_17557);
or U18124 (N_18124,N_17653,N_17751);
xnor U18125 (N_18125,N_17471,N_17683);
nor U18126 (N_18126,N_17473,N_17767);
xnor U18127 (N_18127,N_17107,N_17117);
nand U18128 (N_18128,N_17837,N_17403);
nand U18129 (N_18129,N_17952,N_17932);
xnor U18130 (N_18130,N_17270,N_17858);
xor U18131 (N_18131,N_17418,N_17307);
or U18132 (N_18132,N_17143,N_17780);
xor U18133 (N_18133,N_17662,N_17715);
and U18134 (N_18134,N_17448,N_17734);
nand U18135 (N_18135,N_17073,N_17057);
xor U18136 (N_18136,N_17530,N_17741);
xnor U18137 (N_18137,N_17581,N_17262);
or U18138 (N_18138,N_17510,N_17483);
and U18139 (N_18139,N_17083,N_17463);
nor U18140 (N_18140,N_17648,N_17188);
nor U18141 (N_18141,N_17439,N_17309);
nor U18142 (N_18142,N_17660,N_17053);
or U18143 (N_18143,N_17601,N_17843);
or U18144 (N_18144,N_17772,N_17048);
nand U18145 (N_18145,N_17966,N_17099);
nor U18146 (N_18146,N_17071,N_17330);
or U18147 (N_18147,N_17524,N_17777);
nor U18148 (N_18148,N_17441,N_17793);
xnor U18149 (N_18149,N_17123,N_17673);
nor U18150 (N_18150,N_17708,N_17253);
nor U18151 (N_18151,N_17161,N_17024);
and U18152 (N_18152,N_17237,N_17922);
nor U18153 (N_18153,N_17478,N_17460);
and U18154 (N_18154,N_17695,N_17062);
and U18155 (N_18155,N_17234,N_17654);
nor U18156 (N_18156,N_17261,N_17039);
or U18157 (N_18157,N_17045,N_17643);
or U18158 (N_18158,N_17779,N_17909);
xnor U18159 (N_18159,N_17757,N_17183);
nor U18160 (N_18160,N_17903,N_17802);
or U18161 (N_18161,N_17959,N_17041);
and U18162 (N_18162,N_17028,N_17642);
and U18163 (N_18163,N_17226,N_17753);
or U18164 (N_18164,N_17532,N_17110);
xnor U18165 (N_18165,N_17781,N_17312);
and U18166 (N_18166,N_17893,N_17975);
nand U18167 (N_18167,N_17087,N_17828);
xor U18168 (N_18168,N_17960,N_17467);
nand U18169 (N_18169,N_17611,N_17311);
and U18170 (N_18170,N_17640,N_17598);
or U18171 (N_18171,N_17027,N_17105);
nand U18172 (N_18172,N_17066,N_17218);
nor U18173 (N_18173,N_17022,N_17434);
nand U18174 (N_18174,N_17298,N_17896);
or U18175 (N_18175,N_17101,N_17697);
xnor U18176 (N_18176,N_17529,N_17916);
and U18177 (N_18177,N_17507,N_17880);
or U18178 (N_18178,N_17634,N_17213);
nand U18179 (N_18179,N_17644,N_17908);
xor U18180 (N_18180,N_17387,N_17803);
nor U18181 (N_18181,N_17373,N_17684);
nor U18182 (N_18182,N_17709,N_17356);
nor U18183 (N_18183,N_17449,N_17832);
nand U18184 (N_18184,N_17072,N_17672);
or U18185 (N_18185,N_17316,N_17479);
nor U18186 (N_18186,N_17358,N_17341);
nand U18187 (N_18187,N_17195,N_17186);
nor U18188 (N_18188,N_17225,N_17451);
or U18189 (N_18189,N_17738,N_17852);
nor U18190 (N_18190,N_17372,N_17964);
nor U18191 (N_18191,N_17980,N_17597);
nor U18192 (N_18192,N_17888,N_17406);
and U18193 (N_18193,N_17256,N_17699);
nor U18194 (N_18194,N_17246,N_17020);
nor U18195 (N_18195,N_17770,N_17089);
xnor U18196 (N_18196,N_17205,N_17627);
xor U18197 (N_18197,N_17859,N_17677);
nand U18198 (N_18198,N_17442,N_17572);
xnor U18199 (N_18199,N_17549,N_17681);
nand U18200 (N_18200,N_17386,N_17940);
xor U18201 (N_18201,N_17090,N_17019);
or U18202 (N_18202,N_17798,N_17665);
and U18203 (N_18203,N_17138,N_17602);
nor U18204 (N_18204,N_17806,N_17069);
nand U18205 (N_18205,N_17921,N_17990);
xnor U18206 (N_18206,N_17236,N_17240);
or U18207 (N_18207,N_17915,N_17759);
or U18208 (N_18208,N_17254,N_17269);
nor U18209 (N_18209,N_17374,N_17790);
nand U18210 (N_18210,N_17322,N_17636);
and U18211 (N_18211,N_17263,N_17286);
nor U18212 (N_18212,N_17201,N_17005);
nand U18213 (N_18213,N_17519,N_17422);
nand U18214 (N_18214,N_17174,N_17462);
nand U18215 (N_18215,N_17649,N_17489);
or U18216 (N_18216,N_17513,N_17829);
or U18217 (N_18217,N_17895,N_17369);
xnor U18218 (N_18218,N_17272,N_17856);
and U18219 (N_18219,N_17179,N_17886);
and U18220 (N_18220,N_17578,N_17659);
and U18221 (N_18221,N_17252,N_17637);
or U18222 (N_18222,N_17765,N_17394);
xor U18223 (N_18223,N_17308,N_17250);
xor U18224 (N_18224,N_17862,N_17804);
or U18225 (N_18225,N_17592,N_17492);
nand U18226 (N_18226,N_17542,N_17459);
and U18227 (N_18227,N_17059,N_17354);
or U18228 (N_18228,N_17678,N_17614);
xnor U18229 (N_18229,N_17038,N_17238);
and U18230 (N_18230,N_17742,N_17061);
nand U18231 (N_18231,N_17464,N_17396);
nand U18232 (N_18232,N_17141,N_17052);
nor U18233 (N_18233,N_17713,N_17306);
nor U18234 (N_18234,N_17535,N_17003);
or U18235 (N_18235,N_17575,N_17844);
and U18236 (N_18236,N_17768,N_17378);
nor U18237 (N_18237,N_17259,N_17290);
or U18238 (N_18238,N_17465,N_17521);
or U18239 (N_18239,N_17221,N_17035);
nor U18240 (N_18240,N_17671,N_17554);
and U18241 (N_18241,N_17484,N_17794);
or U18242 (N_18242,N_17206,N_17461);
xnor U18243 (N_18243,N_17562,N_17088);
xnor U18244 (N_18244,N_17251,N_17731);
nor U18245 (N_18245,N_17133,N_17423);
nand U18246 (N_18246,N_17692,N_17274);
and U18247 (N_18247,N_17630,N_17113);
nor U18248 (N_18248,N_17906,N_17687);
and U18249 (N_18249,N_17523,N_17037);
xor U18250 (N_18250,N_17543,N_17408);
or U18251 (N_18251,N_17018,N_17775);
nand U18252 (N_18252,N_17595,N_17116);
and U18253 (N_18253,N_17823,N_17538);
and U18254 (N_18254,N_17157,N_17514);
nor U18255 (N_18255,N_17156,N_17336);
xnor U18256 (N_18256,N_17735,N_17155);
nand U18257 (N_18257,N_17299,N_17623);
or U18258 (N_18258,N_17784,N_17077);
and U18259 (N_18259,N_17043,N_17905);
or U18260 (N_18260,N_17390,N_17297);
or U18261 (N_18261,N_17555,N_17006);
nand U18262 (N_18262,N_17281,N_17056);
nor U18263 (N_18263,N_17146,N_17736);
and U18264 (N_18264,N_17813,N_17176);
or U18265 (N_18265,N_17506,N_17539);
or U18266 (N_18266,N_17106,N_17046);
xor U18267 (N_18267,N_17443,N_17432);
and U18268 (N_18268,N_17496,N_17393);
or U18269 (N_18269,N_17321,N_17785);
nand U18270 (N_18270,N_17603,N_17545);
and U18271 (N_18271,N_17928,N_17782);
nand U18272 (N_18272,N_17481,N_17405);
nor U18273 (N_18273,N_17419,N_17722);
nand U18274 (N_18274,N_17239,N_17212);
xor U18275 (N_18275,N_17170,N_17013);
nand U18276 (N_18276,N_17223,N_17567);
nand U18277 (N_18277,N_17383,N_17067);
or U18278 (N_18278,N_17899,N_17703);
or U18279 (N_18279,N_17375,N_17284);
or U18280 (N_18280,N_17495,N_17491);
xnor U18281 (N_18281,N_17504,N_17967);
xor U18282 (N_18282,N_17998,N_17584);
nor U18283 (N_18283,N_17203,N_17149);
and U18284 (N_18284,N_17565,N_17343);
nand U18285 (N_18285,N_17224,N_17060);
nor U18286 (N_18286,N_17219,N_17727);
xnor U18287 (N_18287,N_17586,N_17850);
nor U18288 (N_18288,N_17885,N_17571);
and U18289 (N_18289,N_17220,N_17177);
and U18290 (N_18290,N_17026,N_17136);
or U18291 (N_18291,N_17892,N_17180);
xnor U18292 (N_18292,N_17118,N_17968);
and U18293 (N_18293,N_17007,N_17395);
xnor U18294 (N_18294,N_17033,N_17951);
nor U18295 (N_18295,N_17548,N_17145);
or U18296 (N_18296,N_17716,N_17428);
nand U18297 (N_18297,N_17445,N_17972);
or U18298 (N_18298,N_17774,N_17392);
or U18299 (N_18299,N_17304,N_17485);
nand U18300 (N_18300,N_17747,N_17446);
or U18301 (N_18301,N_17382,N_17812);
nand U18302 (N_18302,N_17355,N_17400);
and U18303 (N_18303,N_17855,N_17285);
or U18304 (N_18304,N_17108,N_17863);
and U18305 (N_18305,N_17164,N_17198);
nor U18306 (N_18306,N_17208,N_17337);
or U18307 (N_18307,N_17541,N_17137);
nor U18308 (N_18308,N_17163,N_17260);
nand U18309 (N_18309,N_17596,N_17017);
or U18310 (N_18310,N_17458,N_17551);
and U18311 (N_18311,N_17273,N_17616);
nor U18312 (N_18312,N_17323,N_17563);
nor U18313 (N_18313,N_17941,N_17817);
xnor U18314 (N_18314,N_17824,N_17587);
and U18315 (N_18315,N_17352,N_17127);
and U18316 (N_18316,N_17583,N_17502);
xor U18317 (N_18317,N_17897,N_17884);
nor U18318 (N_18318,N_17528,N_17283);
nand U18319 (N_18319,N_17389,N_17749);
or U18320 (N_18320,N_17497,N_17754);
and U18321 (N_18321,N_17870,N_17711);
or U18322 (N_18322,N_17070,N_17267);
or U18323 (N_18323,N_17889,N_17264);
or U18324 (N_18324,N_17875,N_17612);
nor U18325 (N_18325,N_17365,N_17340);
or U18326 (N_18326,N_17086,N_17792);
xor U18327 (N_18327,N_17534,N_17576);
and U18328 (N_18328,N_17417,N_17505);
nor U18329 (N_18329,N_17979,N_17685);
nor U18330 (N_18330,N_17320,N_17574);
nor U18331 (N_18331,N_17376,N_17883);
xnor U18332 (N_18332,N_17955,N_17437);
xnor U18333 (N_18333,N_17958,N_17590);
and U18334 (N_18334,N_17401,N_17540);
and U18335 (N_18335,N_17657,N_17842);
and U18336 (N_18336,N_17200,N_17994);
and U18337 (N_18337,N_17029,N_17691);
nor U18338 (N_18338,N_17839,N_17447);
nand U18339 (N_18339,N_17370,N_17846);
nor U18340 (N_18340,N_17599,N_17525);
or U18341 (N_18341,N_17444,N_17075);
nor U18342 (N_18342,N_17094,N_17516);
or U18343 (N_18343,N_17984,N_17480);
and U18344 (N_18344,N_17878,N_17468);
and U18345 (N_18345,N_17092,N_17153);
or U18346 (N_18346,N_17351,N_17559);
nand U18347 (N_18347,N_17357,N_17078);
nor U18348 (N_18348,N_17494,N_17074);
xor U18349 (N_18349,N_17721,N_17946);
xor U18350 (N_18350,N_17058,N_17385);
nand U18351 (N_18351,N_17364,N_17585);
and U18352 (N_18352,N_17988,N_17904);
or U18353 (N_18353,N_17332,N_17132);
xnor U18354 (N_18354,N_17801,N_17948);
or U18355 (N_18355,N_17420,N_17743);
xnor U18356 (N_18356,N_17799,N_17873);
and U18357 (N_18357,N_17165,N_17936);
and U18358 (N_18358,N_17511,N_17981);
nand U18359 (N_18359,N_17014,N_17139);
nor U18360 (N_18360,N_17953,N_17128);
xor U18361 (N_18361,N_17245,N_17102);
nor U18362 (N_18362,N_17752,N_17553);
or U18363 (N_18363,N_17011,N_17296);
xor U18364 (N_18364,N_17982,N_17580);
and U18365 (N_18365,N_17619,N_17368);
and U18366 (N_18366,N_17631,N_17933);
and U18367 (N_18367,N_17202,N_17430);
nand U18368 (N_18368,N_17725,N_17533);
xor U18369 (N_18369,N_17797,N_17750);
xor U18370 (N_18370,N_17189,N_17537);
xnor U18371 (N_18371,N_17474,N_17871);
or U18372 (N_18372,N_17211,N_17851);
xor U18373 (N_18373,N_17831,N_17938);
xor U18374 (N_18374,N_17204,N_17807);
nand U18375 (N_18375,N_17531,N_17579);
nand U18376 (N_18376,N_17194,N_17380);
or U18377 (N_18377,N_17748,N_17762);
and U18378 (N_18378,N_17593,N_17190);
xnor U18379 (N_18379,N_17600,N_17854);
or U18380 (N_18380,N_17808,N_17324);
and U18381 (N_18381,N_17436,N_17040);
and U18382 (N_18382,N_17977,N_17746);
nand U18383 (N_18383,N_17638,N_17431);
and U18384 (N_18384,N_17278,N_17786);
nor U18385 (N_18385,N_17976,N_17732);
nor U18386 (N_18386,N_17835,N_17398);
and U18387 (N_18387,N_17091,N_17487);
and U18388 (N_18388,N_17773,N_17440);
nand U18389 (N_18389,N_17004,N_17503);
and U18390 (N_18390,N_17907,N_17097);
nor U18391 (N_18391,N_17622,N_17300);
nand U18392 (N_18392,N_17326,N_17676);
and U18393 (N_18393,N_17857,N_17993);
xor U18394 (N_18394,N_17983,N_17103);
xor U18395 (N_18395,N_17944,N_17633);
nor U18396 (N_18396,N_17054,N_17629);
nor U18397 (N_18397,N_17214,N_17778);
or U18398 (N_18398,N_17819,N_17361);
xnor U18399 (N_18399,N_17911,N_17289);
nand U18400 (N_18400,N_17222,N_17995);
nor U18401 (N_18401,N_17950,N_17740);
and U18402 (N_18402,N_17310,N_17758);
nand U18403 (N_18403,N_17151,N_17129);
or U18404 (N_18404,N_17021,N_17881);
or U18405 (N_18405,N_17869,N_17178);
and U18406 (N_18406,N_17547,N_17680);
nand U18407 (N_18407,N_17814,N_17818);
xor U18408 (N_18408,N_17864,N_17536);
xnor U18409 (N_18409,N_17745,N_17302);
nor U18410 (N_18410,N_17546,N_17796);
nand U18411 (N_18411,N_17902,N_17724);
or U18412 (N_18412,N_17388,N_17658);
or U18413 (N_18413,N_17140,N_17560);
nand U18414 (N_18414,N_17615,N_17265);
nor U18415 (N_18415,N_17049,N_17723);
nor U18416 (N_18416,N_17656,N_17647);
nor U18417 (N_18417,N_17872,N_17080);
nor U18418 (N_18418,N_17192,N_17475);
and U18419 (N_18419,N_17241,N_17606);
nand U18420 (N_18420,N_17918,N_17945);
nand U18421 (N_18421,N_17701,N_17159);
nand U18422 (N_18422,N_17833,N_17318);
nor U18423 (N_18423,N_17877,N_17167);
and U18424 (N_18424,N_17109,N_17707);
and U18425 (N_18425,N_17588,N_17454);
nand U18426 (N_18426,N_17834,N_17825);
nor U18427 (N_18427,N_17002,N_17230);
or U18428 (N_18428,N_17415,N_17328);
and U18429 (N_18429,N_17999,N_17791);
or U18430 (N_18430,N_17866,N_17313);
or U18431 (N_18431,N_17717,N_17114);
nor U18432 (N_18432,N_17249,N_17173);
xor U18433 (N_18433,N_17142,N_17667);
nand U18434 (N_18434,N_17978,N_17081);
nand U18435 (N_18435,N_17670,N_17215);
or U18436 (N_18436,N_17131,N_17096);
nand U18437 (N_18437,N_17666,N_17455);
xnor U18438 (N_18438,N_17836,N_17147);
nor U18439 (N_18439,N_17686,N_17632);
xnor U18440 (N_18440,N_17126,N_17705);
or U18441 (N_18441,N_17044,N_17805);
nand U18442 (N_18442,N_17635,N_17217);
or U18443 (N_18443,N_17690,N_17242);
and U18444 (N_18444,N_17231,N_17737);
nor U18445 (N_18445,N_17085,N_17258);
and U18446 (N_18446,N_17093,N_17925);
nor U18447 (N_18447,N_17384,N_17424);
nand U18448 (N_18448,N_17303,N_17853);
xnor U18449 (N_18449,N_17901,N_17344);
and U18450 (N_18450,N_17329,N_17739);
nor U18451 (N_18451,N_17119,N_17452);
and U18452 (N_18452,N_17359,N_17498);
nand U18453 (N_18453,N_17898,N_17882);
nand U18454 (N_18454,N_17232,N_17816);
or U18455 (N_18455,N_17949,N_17961);
nor U18456 (N_18456,N_17025,N_17193);
and U18457 (N_18457,N_17499,N_17065);
and U18458 (N_18458,N_17334,N_17350);
and U18459 (N_18459,N_17970,N_17733);
and U18460 (N_18460,N_17120,N_17032);
nor U18461 (N_18461,N_17122,N_17047);
and U18462 (N_18462,N_17111,N_17197);
and U18463 (N_18463,N_17930,N_17134);
nand U18464 (N_18464,N_17849,N_17427);
xnor U18465 (N_18465,N_17865,N_17076);
nor U18466 (N_18466,N_17509,N_17207);
nand U18467 (N_18467,N_17130,N_17199);
or U18468 (N_18468,N_17421,N_17228);
nand U18469 (N_18469,N_17000,N_17327);
nand U18470 (N_18470,N_17371,N_17675);
nor U18471 (N_18471,N_17031,N_17991);
and U18472 (N_18472,N_17900,N_17556);
and U18473 (N_18473,N_17710,N_17187);
and U18474 (N_18474,N_17172,N_17247);
xnor U18475 (N_18475,N_17943,N_17135);
nand U18476 (N_18476,N_17712,N_17182);
nand U18477 (N_18477,N_17760,N_17890);
and U18478 (N_18478,N_17416,N_17160);
nand U18479 (N_18479,N_17104,N_17347);
nor U18480 (N_18480,N_17335,N_17861);
or U18481 (N_18481,N_17399,N_17552);
and U18482 (N_18482,N_17582,N_17573);
nor U18483 (N_18483,N_17233,N_17397);
xor U18484 (N_18484,N_17271,N_17702);
and U18485 (N_18485,N_17009,N_17169);
nor U18486 (N_18486,N_17646,N_17435);
nor U18487 (N_18487,N_17293,N_17338);
nand U18488 (N_18488,N_17426,N_17477);
and U18489 (N_18489,N_17809,N_17704);
xnor U18490 (N_18490,N_17728,N_17121);
nor U18491 (N_18491,N_17971,N_17112);
xnor U18492 (N_18492,N_17912,N_17689);
or U18493 (N_18493,N_17050,N_17411);
and U18494 (N_18494,N_17954,N_17319);
or U18495 (N_18495,N_17764,N_17929);
xnor U18496 (N_18496,N_17655,N_17413);
nand U18497 (N_18497,N_17800,N_17755);
nor U18498 (N_18498,N_17162,N_17425);
and U18499 (N_18499,N_17342,N_17301);
nand U18500 (N_18500,N_17790,N_17411);
xor U18501 (N_18501,N_17844,N_17991);
nor U18502 (N_18502,N_17633,N_17254);
nand U18503 (N_18503,N_17624,N_17716);
and U18504 (N_18504,N_17247,N_17739);
nand U18505 (N_18505,N_17479,N_17220);
xnor U18506 (N_18506,N_17095,N_17994);
xor U18507 (N_18507,N_17373,N_17204);
nor U18508 (N_18508,N_17124,N_17525);
nor U18509 (N_18509,N_17337,N_17555);
or U18510 (N_18510,N_17109,N_17546);
and U18511 (N_18511,N_17953,N_17544);
nor U18512 (N_18512,N_17611,N_17842);
and U18513 (N_18513,N_17894,N_17690);
xor U18514 (N_18514,N_17862,N_17738);
or U18515 (N_18515,N_17178,N_17845);
or U18516 (N_18516,N_17451,N_17716);
nor U18517 (N_18517,N_17666,N_17952);
xnor U18518 (N_18518,N_17936,N_17610);
or U18519 (N_18519,N_17053,N_17440);
and U18520 (N_18520,N_17398,N_17944);
nor U18521 (N_18521,N_17405,N_17244);
or U18522 (N_18522,N_17066,N_17091);
xor U18523 (N_18523,N_17350,N_17858);
or U18524 (N_18524,N_17075,N_17018);
xor U18525 (N_18525,N_17897,N_17139);
or U18526 (N_18526,N_17270,N_17610);
nand U18527 (N_18527,N_17738,N_17453);
nor U18528 (N_18528,N_17858,N_17848);
nand U18529 (N_18529,N_17014,N_17863);
and U18530 (N_18530,N_17491,N_17115);
or U18531 (N_18531,N_17228,N_17728);
or U18532 (N_18532,N_17492,N_17760);
nand U18533 (N_18533,N_17673,N_17853);
and U18534 (N_18534,N_17456,N_17891);
or U18535 (N_18535,N_17168,N_17478);
nor U18536 (N_18536,N_17819,N_17420);
nand U18537 (N_18537,N_17055,N_17640);
nand U18538 (N_18538,N_17283,N_17060);
or U18539 (N_18539,N_17285,N_17264);
or U18540 (N_18540,N_17470,N_17302);
or U18541 (N_18541,N_17383,N_17539);
and U18542 (N_18542,N_17271,N_17548);
nor U18543 (N_18543,N_17251,N_17239);
and U18544 (N_18544,N_17644,N_17586);
or U18545 (N_18545,N_17388,N_17021);
or U18546 (N_18546,N_17982,N_17820);
or U18547 (N_18547,N_17060,N_17528);
nor U18548 (N_18548,N_17060,N_17114);
and U18549 (N_18549,N_17080,N_17741);
nor U18550 (N_18550,N_17648,N_17905);
nor U18551 (N_18551,N_17251,N_17529);
and U18552 (N_18552,N_17821,N_17511);
xnor U18553 (N_18553,N_17329,N_17255);
nand U18554 (N_18554,N_17051,N_17687);
nor U18555 (N_18555,N_17898,N_17801);
xnor U18556 (N_18556,N_17477,N_17255);
nand U18557 (N_18557,N_17046,N_17574);
or U18558 (N_18558,N_17998,N_17359);
xnor U18559 (N_18559,N_17034,N_17023);
nand U18560 (N_18560,N_17960,N_17711);
nand U18561 (N_18561,N_17589,N_17870);
and U18562 (N_18562,N_17113,N_17612);
nor U18563 (N_18563,N_17485,N_17202);
xor U18564 (N_18564,N_17779,N_17470);
nand U18565 (N_18565,N_17001,N_17095);
nand U18566 (N_18566,N_17475,N_17139);
and U18567 (N_18567,N_17930,N_17607);
nor U18568 (N_18568,N_17284,N_17567);
or U18569 (N_18569,N_17122,N_17747);
xor U18570 (N_18570,N_17223,N_17026);
xnor U18571 (N_18571,N_17880,N_17680);
or U18572 (N_18572,N_17164,N_17369);
and U18573 (N_18573,N_17504,N_17948);
or U18574 (N_18574,N_17385,N_17992);
or U18575 (N_18575,N_17776,N_17174);
nor U18576 (N_18576,N_17608,N_17454);
or U18577 (N_18577,N_17441,N_17360);
or U18578 (N_18578,N_17207,N_17075);
or U18579 (N_18579,N_17173,N_17903);
xor U18580 (N_18580,N_17815,N_17090);
and U18581 (N_18581,N_17599,N_17192);
nor U18582 (N_18582,N_17072,N_17870);
or U18583 (N_18583,N_17813,N_17456);
nor U18584 (N_18584,N_17625,N_17883);
nor U18585 (N_18585,N_17310,N_17463);
xor U18586 (N_18586,N_17303,N_17966);
xor U18587 (N_18587,N_17254,N_17993);
and U18588 (N_18588,N_17794,N_17343);
and U18589 (N_18589,N_17846,N_17067);
or U18590 (N_18590,N_17427,N_17945);
and U18591 (N_18591,N_17337,N_17420);
and U18592 (N_18592,N_17084,N_17806);
xor U18593 (N_18593,N_17001,N_17592);
nand U18594 (N_18594,N_17763,N_17943);
or U18595 (N_18595,N_17975,N_17516);
nand U18596 (N_18596,N_17547,N_17536);
or U18597 (N_18597,N_17885,N_17741);
nor U18598 (N_18598,N_17714,N_17249);
or U18599 (N_18599,N_17231,N_17649);
nand U18600 (N_18600,N_17219,N_17149);
xor U18601 (N_18601,N_17803,N_17077);
nand U18602 (N_18602,N_17849,N_17752);
or U18603 (N_18603,N_17617,N_17137);
xnor U18604 (N_18604,N_17740,N_17492);
and U18605 (N_18605,N_17638,N_17791);
or U18606 (N_18606,N_17872,N_17899);
nand U18607 (N_18607,N_17171,N_17561);
and U18608 (N_18608,N_17217,N_17290);
nor U18609 (N_18609,N_17474,N_17477);
nor U18610 (N_18610,N_17888,N_17325);
and U18611 (N_18611,N_17505,N_17867);
xnor U18612 (N_18612,N_17755,N_17354);
or U18613 (N_18613,N_17327,N_17591);
and U18614 (N_18614,N_17283,N_17305);
and U18615 (N_18615,N_17218,N_17493);
or U18616 (N_18616,N_17477,N_17319);
nor U18617 (N_18617,N_17649,N_17230);
xor U18618 (N_18618,N_17431,N_17763);
xor U18619 (N_18619,N_17851,N_17777);
xnor U18620 (N_18620,N_17302,N_17438);
and U18621 (N_18621,N_17733,N_17553);
or U18622 (N_18622,N_17386,N_17176);
nor U18623 (N_18623,N_17768,N_17553);
xor U18624 (N_18624,N_17693,N_17035);
and U18625 (N_18625,N_17614,N_17626);
nor U18626 (N_18626,N_17276,N_17711);
or U18627 (N_18627,N_17537,N_17014);
nand U18628 (N_18628,N_17613,N_17769);
xor U18629 (N_18629,N_17118,N_17162);
or U18630 (N_18630,N_17868,N_17438);
nand U18631 (N_18631,N_17381,N_17291);
or U18632 (N_18632,N_17378,N_17707);
nand U18633 (N_18633,N_17213,N_17708);
nor U18634 (N_18634,N_17725,N_17376);
xnor U18635 (N_18635,N_17477,N_17214);
xor U18636 (N_18636,N_17877,N_17726);
nor U18637 (N_18637,N_17596,N_17615);
nor U18638 (N_18638,N_17243,N_17745);
xor U18639 (N_18639,N_17738,N_17546);
nor U18640 (N_18640,N_17548,N_17706);
or U18641 (N_18641,N_17426,N_17437);
xnor U18642 (N_18642,N_17173,N_17292);
nand U18643 (N_18643,N_17433,N_17297);
or U18644 (N_18644,N_17115,N_17475);
nand U18645 (N_18645,N_17580,N_17077);
or U18646 (N_18646,N_17583,N_17941);
nor U18647 (N_18647,N_17868,N_17996);
xor U18648 (N_18648,N_17506,N_17655);
nand U18649 (N_18649,N_17102,N_17702);
xor U18650 (N_18650,N_17307,N_17570);
xor U18651 (N_18651,N_17554,N_17096);
or U18652 (N_18652,N_17242,N_17713);
nor U18653 (N_18653,N_17383,N_17251);
or U18654 (N_18654,N_17173,N_17968);
nor U18655 (N_18655,N_17649,N_17178);
and U18656 (N_18656,N_17399,N_17066);
nor U18657 (N_18657,N_17293,N_17472);
xnor U18658 (N_18658,N_17206,N_17873);
nand U18659 (N_18659,N_17021,N_17249);
nand U18660 (N_18660,N_17082,N_17156);
nand U18661 (N_18661,N_17053,N_17600);
and U18662 (N_18662,N_17767,N_17660);
or U18663 (N_18663,N_17558,N_17930);
and U18664 (N_18664,N_17271,N_17823);
nand U18665 (N_18665,N_17898,N_17707);
nor U18666 (N_18666,N_17604,N_17500);
nand U18667 (N_18667,N_17592,N_17468);
xor U18668 (N_18668,N_17135,N_17380);
nand U18669 (N_18669,N_17601,N_17785);
xor U18670 (N_18670,N_17664,N_17120);
or U18671 (N_18671,N_17523,N_17916);
nand U18672 (N_18672,N_17717,N_17119);
nor U18673 (N_18673,N_17698,N_17426);
and U18674 (N_18674,N_17956,N_17951);
nor U18675 (N_18675,N_17560,N_17070);
nand U18676 (N_18676,N_17858,N_17625);
and U18677 (N_18677,N_17729,N_17553);
and U18678 (N_18678,N_17627,N_17733);
xor U18679 (N_18679,N_17197,N_17107);
nor U18680 (N_18680,N_17898,N_17981);
and U18681 (N_18681,N_17889,N_17797);
nand U18682 (N_18682,N_17776,N_17811);
nor U18683 (N_18683,N_17884,N_17134);
xor U18684 (N_18684,N_17534,N_17199);
or U18685 (N_18685,N_17123,N_17574);
or U18686 (N_18686,N_17050,N_17887);
xnor U18687 (N_18687,N_17969,N_17611);
nand U18688 (N_18688,N_17044,N_17174);
xnor U18689 (N_18689,N_17711,N_17900);
xnor U18690 (N_18690,N_17647,N_17770);
nand U18691 (N_18691,N_17481,N_17045);
xor U18692 (N_18692,N_17607,N_17518);
and U18693 (N_18693,N_17253,N_17457);
nor U18694 (N_18694,N_17354,N_17872);
nand U18695 (N_18695,N_17944,N_17667);
xor U18696 (N_18696,N_17234,N_17180);
or U18697 (N_18697,N_17875,N_17273);
xor U18698 (N_18698,N_17142,N_17392);
nor U18699 (N_18699,N_17405,N_17121);
or U18700 (N_18700,N_17028,N_17862);
nor U18701 (N_18701,N_17024,N_17766);
and U18702 (N_18702,N_17628,N_17459);
xnor U18703 (N_18703,N_17346,N_17569);
and U18704 (N_18704,N_17646,N_17721);
nor U18705 (N_18705,N_17608,N_17940);
or U18706 (N_18706,N_17717,N_17253);
and U18707 (N_18707,N_17401,N_17250);
nand U18708 (N_18708,N_17750,N_17438);
nand U18709 (N_18709,N_17765,N_17969);
xor U18710 (N_18710,N_17987,N_17738);
nand U18711 (N_18711,N_17345,N_17259);
and U18712 (N_18712,N_17038,N_17587);
nor U18713 (N_18713,N_17193,N_17365);
nand U18714 (N_18714,N_17995,N_17359);
nor U18715 (N_18715,N_17745,N_17328);
xnor U18716 (N_18716,N_17287,N_17208);
nor U18717 (N_18717,N_17760,N_17759);
and U18718 (N_18718,N_17753,N_17421);
and U18719 (N_18719,N_17692,N_17139);
nand U18720 (N_18720,N_17822,N_17447);
xnor U18721 (N_18721,N_17266,N_17482);
nand U18722 (N_18722,N_17167,N_17002);
or U18723 (N_18723,N_17145,N_17861);
nor U18724 (N_18724,N_17955,N_17930);
and U18725 (N_18725,N_17953,N_17658);
nand U18726 (N_18726,N_17523,N_17471);
or U18727 (N_18727,N_17671,N_17150);
nor U18728 (N_18728,N_17926,N_17401);
nand U18729 (N_18729,N_17688,N_17054);
nor U18730 (N_18730,N_17465,N_17937);
nor U18731 (N_18731,N_17936,N_17750);
xnor U18732 (N_18732,N_17789,N_17259);
and U18733 (N_18733,N_17362,N_17499);
xnor U18734 (N_18734,N_17160,N_17689);
or U18735 (N_18735,N_17492,N_17111);
xnor U18736 (N_18736,N_17463,N_17456);
and U18737 (N_18737,N_17739,N_17799);
nand U18738 (N_18738,N_17853,N_17203);
and U18739 (N_18739,N_17364,N_17052);
nand U18740 (N_18740,N_17121,N_17783);
nand U18741 (N_18741,N_17143,N_17823);
xnor U18742 (N_18742,N_17950,N_17392);
or U18743 (N_18743,N_17928,N_17927);
or U18744 (N_18744,N_17910,N_17897);
nand U18745 (N_18745,N_17453,N_17438);
nor U18746 (N_18746,N_17770,N_17189);
or U18747 (N_18747,N_17368,N_17315);
xor U18748 (N_18748,N_17144,N_17756);
and U18749 (N_18749,N_17795,N_17331);
nor U18750 (N_18750,N_17825,N_17498);
or U18751 (N_18751,N_17727,N_17215);
xnor U18752 (N_18752,N_17485,N_17672);
xor U18753 (N_18753,N_17552,N_17909);
nor U18754 (N_18754,N_17859,N_17525);
nand U18755 (N_18755,N_17007,N_17366);
nor U18756 (N_18756,N_17955,N_17343);
xnor U18757 (N_18757,N_17355,N_17450);
xor U18758 (N_18758,N_17371,N_17644);
xnor U18759 (N_18759,N_17053,N_17930);
nand U18760 (N_18760,N_17261,N_17806);
xnor U18761 (N_18761,N_17084,N_17160);
xor U18762 (N_18762,N_17782,N_17293);
or U18763 (N_18763,N_17580,N_17813);
or U18764 (N_18764,N_17595,N_17991);
nor U18765 (N_18765,N_17127,N_17438);
or U18766 (N_18766,N_17309,N_17358);
or U18767 (N_18767,N_17790,N_17287);
nor U18768 (N_18768,N_17122,N_17050);
nor U18769 (N_18769,N_17843,N_17783);
xnor U18770 (N_18770,N_17734,N_17408);
and U18771 (N_18771,N_17437,N_17872);
xor U18772 (N_18772,N_17833,N_17090);
or U18773 (N_18773,N_17925,N_17269);
nor U18774 (N_18774,N_17968,N_17995);
or U18775 (N_18775,N_17186,N_17274);
nand U18776 (N_18776,N_17403,N_17128);
or U18777 (N_18777,N_17150,N_17841);
nand U18778 (N_18778,N_17617,N_17539);
nand U18779 (N_18779,N_17968,N_17497);
xnor U18780 (N_18780,N_17540,N_17452);
xnor U18781 (N_18781,N_17879,N_17630);
and U18782 (N_18782,N_17039,N_17245);
xor U18783 (N_18783,N_17953,N_17510);
xor U18784 (N_18784,N_17270,N_17455);
nand U18785 (N_18785,N_17848,N_17884);
xor U18786 (N_18786,N_17533,N_17716);
xor U18787 (N_18787,N_17843,N_17038);
xnor U18788 (N_18788,N_17275,N_17245);
nor U18789 (N_18789,N_17729,N_17211);
or U18790 (N_18790,N_17693,N_17337);
nand U18791 (N_18791,N_17368,N_17676);
nand U18792 (N_18792,N_17225,N_17739);
or U18793 (N_18793,N_17022,N_17064);
xnor U18794 (N_18794,N_17921,N_17427);
xor U18795 (N_18795,N_17350,N_17805);
nor U18796 (N_18796,N_17637,N_17477);
nand U18797 (N_18797,N_17558,N_17574);
nor U18798 (N_18798,N_17667,N_17378);
and U18799 (N_18799,N_17752,N_17071);
nand U18800 (N_18800,N_17315,N_17549);
nor U18801 (N_18801,N_17107,N_17271);
nor U18802 (N_18802,N_17778,N_17947);
xnor U18803 (N_18803,N_17964,N_17055);
or U18804 (N_18804,N_17661,N_17054);
nand U18805 (N_18805,N_17778,N_17692);
nand U18806 (N_18806,N_17105,N_17967);
or U18807 (N_18807,N_17788,N_17325);
and U18808 (N_18808,N_17215,N_17366);
nand U18809 (N_18809,N_17678,N_17174);
xor U18810 (N_18810,N_17310,N_17354);
nor U18811 (N_18811,N_17384,N_17348);
or U18812 (N_18812,N_17894,N_17779);
or U18813 (N_18813,N_17942,N_17882);
nor U18814 (N_18814,N_17258,N_17990);
nor U18815 (N_18815,N_17063,N_17651);
xor U18816 (N_18816,N_17832,N_17758);
xnor U18817 (N_18817,N_17304,N_17120);
nor U18818 (N_18818,N_17123,N_17132);
or U18819 (N_18819,N_17774,N_17411);
or U18820 (N_18820,N_17284,N_17674);
nand U18821 (N_18821,N_17544,N_17197);
or U18822 (N_18822,N_17840,N_17627);
nor U18823 (N_18823,N_17438,N_17120);
nor U18824 (N_18824,N_17716,N_17410);
nand U18825 (N_18825,N_17509,N_17565);
and U18826 (N_18826,N_17337,N_17977);
and U18827 (N_18827,N_17038,N_17579);
or U18828 (N_18828,N_17479,N_17917);
and U18829 (N_18829,N_17145,N_17745);
and U18830 (N_18830,N_17622,N_17474);
nor U18831 (N_18831,N_17402,N_17373);
nor U18832 (N_18832,N_17600,N_17495);
xor U18833 (N_18833,N_17473,N_17464);
and U18834 (N_18834,N_17916,N_17245);
xnor U18835 (N_18835,N_17639,N_17408);
xnor U18836 (N_18836,N_17610,N_17493);
nand U18837 (N_18837,N_17575,N_17613);
or U18838 (N_18838,N_17729,N_17518);
nand U18839 (N_18839,N_17146,N_17386);
or U18840 (N_18840,N_17587,N_17263);
xor U18841 (N_18841,N_17992,N_17548);
xnor U18842 (N_18842,N_17433,N_17052);
and U18843 (N_18843,N_17653,N_17437);
nor U18844 (N_18844,N_17738,N_17639);
nand U18845 (N_18845,N_17808,N_17063);
xor U18846 (N_18846,N_17107,N_17571);
nor U18847 (N_18847,N_17957,N_17636);
xnor U18848 (N_18848,N_17622,N_17642);
xor U18849 (N_18849,N_17610,N_17376);
nor U18850 (N_18850,N_17463,N_17770);
nor U18851 (N_18851,N_17367,N_17612);
nand U18852 (N_18852,N_17999,N_17853);
xor U18853 (N_18853,N_17350,N_17645);
nand U18854 (N_18854,N_17509,N_17717);
xor U18855 (N_18855,N_17532,N_17773);
nand U18856 (N_18856,N_17286,N_17986);
nand U18857 (N_18857,N_17683,N_17261);
or U18858 (N_18858,N_17874,N_17055);
and U18859 (N_18859,N_17909,N_17471);
nor U18860 (N_18860,N_17252,N_17685);
and U18861 (N_18861,N_17766,N_17833);
and U18862 (N_18862,N_17705,N_17984);
and U18863 (N_18863,N_17453,N_17114);
or U18864 (N_18864,N_17856,N_17008);
and U18865 (N_18865,N_17291,N_17496);
and U18866 (N_18866,N_17514,N_17449);
nand U18867 (N_18867,N_17618,N_17049);
nand U18868 (N_18868,N_17587,N_17229);
and U18869 (N_18869,N_17407,N_17041);
nand U18870 (N_18870,N_17581,N_17967);
and U18871 (N_18871,N_17270,N_17375);
xor U18872 (N_18872,N_17489,N_17744);
xor U18873 (N_18873,N_17333,N_17782);
and U18874 (N_18874,N_17767,N_17518);
xnor U18875 (N_18875,N_17424,N_17056);
or U18876 (N_18876,N_17942,N_17640);
xnor U18877 (N_18877,N_17438,N_17673);
nor U18878 (N_18878,N_17349,N_17851);
nor U18879 (N_18879,N_17126,N_17921);
nor U18880 (N_18880,N_17401,N_17787);
or U18881 (N_18881,N_17046,N_17602);
xnor U18882 (N_18882,N_17636,N_17282);
xor U18883 (N_18883,N_17249,N_17389);
or U18884 (N_18884,N_17192,N_17578);
xor U18885 (N_18885,N_17838,N_17922);
nand U18886 (N_18886,N_17259,N_17626);
nand U18887 (N_18887,N_17602,N_17343);
xnor U18888 (N_18888,N_17688,N_17265);
and U18889 (N_18889,N_17013,N_17670);
nand U18890 (N_18890,N_17490,N_17908);
nor U18891 (N_18891,N_17068,N_17232);
nor U18892 (N_18892,N_17240,N_17869);
and U18893 (N_18893,N_17151,N_17142);
or U18894 (N_18894,N_17161,N_17127);
nor U18895 (N_18895,N_17680,N_17743);
or U18896 (N_18896,N_17067,N_17045);
and U18897 (N_18897,N_17697,N_17923);
xnor U18898 (N_18898,N_17615,N_17494);
nor U18899 (N_18899,N_17300,N_17815);
nor U18900 (N_18900,N_17082,N_17904);
nand U18901 (N_18901,N_17480,N_17523);
and U18902 (N_18902,N_17541,N_17899);
nand U18903 (N_18903,N_17741,N_17805);
nor U18904 (N_18904,N_17298,N_17569);
nand U18905 (N_18905,N_17410,N_17571);
and U18906 (N_18906,N_17813,N_17060);
nand U18907 (N_18907,N_17705,N_17157);
or U18908 (N_18908,N_17924,N_17551);
xor U18909 (N_18909,N_17609,N_17176);
nor U18910 (N_18910,N_17861,N_17715);
nor U18911 (N_18911,N_17876,N_17655);
xor U18912 (N_18912,N_17448,N_17435);
or U18913 (N_18913,N_17740,N_17932);
or U18914 (N_18914,N_17738,N_17256);
or U18915 (N_18915,N_17295,N_17245);
or U18916 (N_18916,N_17541,N_17874);
or U18917 (N_18917,N_17483,N_17485);
or U18918 (N_18918,N_17824,N_17654);
or U18919 (N_18919,N_17717,N_17608);
and U18920 (N_18920,N_17861,N_17753);
nand U18921 (N_18921,N_17514,N_17727);
nand U18922 (N_18922,N_17381,N_17312);
nand U18923 (N_18923,N_17728,N_17028);
xnor U18924 (N_18924,N_17734,N_17294);
nand U18925 (N_18925,N_17377,N_17757);
and U18926 (N_18926,N_17775,N_17817);
nand U18927 (N_18927,N_17133,N_17062);
xor U18928 (N_18928,N_17174,N_17654);
or U18929 (N_18929,N_17913,N_17920);
nor U18930 (N_18930,N_17708,N_17447);
or U18931 (N_18931,N_17843,N_17513);
or U18932 (N_18932,N_17189,N_17802);
or U18933 (N_18933,N_17096,N_17854);
or U18934 (N_18934,N_17614,N_17232);
and U18935 (N_18935,N_17831,N_17443);
and U18936 (N_18936,N_17279,N_17260);
nor U18937 (N_18937,N_17425,N_17947);
and U18938 (N_18938,N_17784,N_17032);
and U18939 (N_18939,N_17570,N_17182);
and U18940 (N_18940,N_17059,N_17464);
and U18941 (N_18941,N_17946,N_17280);
or U18942 (N_18942,N_17864,N_17977);
xor U18943 (N_18943,N_17458,N_17374);
nand U18944 (N_18944,N_17985,N_17975);
or U18945 (N_18945,N_17450,N_17035);
nor U18946 (N_18946,N_17510,N_17425);
or U18947 (N_18947,N_17470,N_17310);
or U18948 (N_18948,N_17373,N_17440);
or U18949 (N_18949,N_17200,N_17075);
nor U18950 (N_18950,N_17106,N_17296);
nand U18951 (N_18951,N_17684,N_17083);
nor U18952 (N_18952,N_17102,N_17206);
nor U18953 (N_18953,N_17171,N_17478);
nor U18954 (N_18954,N_17833,N_17016);
and U18955 (N_18955,N_17023,N_17688);
or U18956 (N_18956,N_17233,N_17789);
nand U18957 (N_18957,N_17283,N_17606);
or U18958 (N_18958,N_17361,N_17014);
nor U18959 (N_18959,N_17376,N_17249);
nand U18960 (N_18960,N_17736,N_17297);
nor U18961 (N_18961,N_17815,N_17985);
nor U18962 (N_18962,N_17104,N_17981);
nand U18963 (N_18963,N_17568,N_17020);
and U18964 (N_18964,N_17208,N_17251);
or U18965 (N_18965,N_17807,N_17526);
and U18966 (N_18966,N_17812,N_17573);
or U18967 (N_18967,N_17323,N_17264);
nand U18968 (N_18968,N_17156,N_17185);
or U18969 (N_18969,N_17406,N_17394);
xnor U18970 (N_18970,N_17615,N_17951);
and U18971 (N_18971,N_17569,N_17247);
or U18972 (N_18972,N_17044,N_17118);
nand U18973 (N_18973,N_17569,N_17292);
xor U18974 (N_18974,N_17756,N_17795);
nor U18975 (N_18975,N_17000,N_17221);
nand U18976 (N_18976,N_17830,N_17800);
xor U18977 (N_18977,N_17442,N_17133);
and U18978 (N_18978,N_17388,N_17332);
or U18979 (N_18979,N_17089,N_17995);
nand U18980 (N_18980,N_17718,N_17669);
nor U18981 (N_18981,N_17065,N_17943);
or U18982 (N_18982,N_17720,N_17529);
nand U18983 (N_18983,N_17876,N_17187);
nor U18984 (N_18984,N_17645,N_17585);
and U18985 (N_18985,N_17543,N_17339);
nand U18986 (N_18986,N_17491,N_17668);
nand U18987 (N_18987,N_17228,N_17458);
nor U18988 (N_18988,N_17801,N_17463);
nand U18989 (N_18989,N_17684,N_17802);
nor U18990 (N_18990,N_17961,N_17040);
nor U18991 (N_18991,N_17707,N_17055);
or U18992 (N_18992,N_17129,N_17384);
and U18993 (N_18993,N_17007,N_17021);
nor U18994 (N_18994,N_17915,N_17931);
and U18995 (N_18995,N_17724,N_17076);
and U18996 (N_18996,N_17093,N_17700);
and U18997 (N_18997,N_17967,N_17028);
or U18998 (N_18998,N_17655,N_17765);
nand U18999 (N_18999,N_17149,N_17801);
xnor U19000 (N_19000,N_18211,N_18507);
and U19001 (N_19001,N_18321,N_18739);
nand U19002 (N_19002,N_18874,N_18943);
and U19003 (N_19003,N_18264,N_18169);
nor U19004 (N_19004,N_18805,N_18858);
and U19005 (N_19005,N_18661,N_18896);
nand U19006 (N_19006,N_18272,N_18815);
or U19007 (N_19007,N_18377,N_18766);
xor U19008 (N_19008,N_18885,N_18775);
nor U19009 (N_19009,N_18449,N_18487);
xnor U19010 (N_19010,N_18140,N_18654);
or U19011 (N_19011,N_18594,N_18154);
or U19012 (N_19012,N_18286,N_18687);
or U19013 (N_19013,N_18488,N_18907);
or U19014 (N_19014,N_18511,N_18886);
nand U19015 (N_19015,N_18653,N_18655);
nor U19016 (N_19016,N_18365,N_18199);
and U19017 (N_19017,N_18938,N_18109);
xor U19018 (N_19018,N_18521,N_18880);
and U19019 (N_19019,N_18870,N_18191);
or U19020 (N_19020,N_18131,N_18713);
xor U19021 (N_19021,N_18071,N_18577);
nand U19022 (N_19022,N_18470,N_18010);
or U19023 (N_19023,N_18812,N_18080);
and U19024 (N_19024,N_18808,N_18930);
nor U19025 (N_19025,N_18146,N_18659);
and U19026 (N_19026,N_18972,N_18343);
nand U19027 (N_19027,N_18643,N_18961);
xnor U19028 (N_19028,N_18072,N_18899);
nor U19029 (N_19029,N_18416,N_18921);
nor U19030 (N_19030,N_18711,N_18786);
and U19031 (N_19031,N_18218,N_18920);
xor U19032 (N_19032,N_18969,N_18064);
xnor U19033 (N_19033,N_18835,N_18955);
and U19034 (N_19034,N_18161,N_18819);
or U19035 (N_19035,N_18558,N_18166);
nor U19036 (N_19036,N_18438,N_18322);
or U19037 (N_19037,N_18928,N_18867);
nand U19038 (N_19038,N_18872,N_18593);
and U19039 (N_19039,N_18656,N_18219);
xnor U19040 (N_19040,N_18571,N_18890);
xnor U19041 (N_19041,N_18691,N_18601);
or U19042 (N_19042,N_18744,N_18276);
or U19043 (N_19043,N_18228,N_18401);
and U19044 (N_19044,N_18498,N_18101);
or U19045 (N_19045,N_18714,N_18495);
nand U19046 (N_19046,N_18372,N_18663);
nor U19047 (N_19047,N_18927,N_18120);
or U19048 (N_19048,N_18031,N_18328);
or U19049 (N_19049,N_18825,N_18137);
nor U19050 (N_19050,N_18579,N_18528);
nand U19051 (N_19051,N_18142,N_18323);
nand U19052 (N_19052,N_18686,N_18596);
and U19053 (N_19053,N_18809,N_18044);
and U19054 (N_19054,N_18512,N_18701);
or U19055 (N_19055,N_18919,N_18423);
xnor U19056 (N_19056,N_18251,N_18810);
xnor U19057 (N_19057,N_18267,N_18944);
or U19058 (N_19058,N_18113,N_18348);
and U19059 (N_19059,N_18734,N_18982);
nand U19060 (N_19060,N_18906,N_18402);
or U19061 (N_19061,N_18724,N_18300);
xnor U19062 (N_19062,N_18547,N_18623);
and U19063 (N_19063,N_18699,N_18868);
and U19064 (N_19064,N_18570,N_18407);
nand U19065 (N_19065,N_18610,N_18752);
nand U19066 (N_19066,N_18155,N_18774);
nand U19067 (N_19067,N_18616,N_18184);
nor U19068 (N_19068,N_18340,N_18909);
and U19069 (N_19069,N_18222,N_18989);
and U19070 (N_19070,N_18738,N_18213);
nor U19071 (N_19071,N_18134,N_18849);
nand U19072 (N_19072,N_18591,N_18248);
nand U19073 (N_19073,N_18564,N_18991);
or U19074 (N_19074,N_18782,N_18110);
or U19075 (N_19075,N_18959,N_18006);
nand U19076 (N_19076,N_18428,N_18386);
and U19077 (N_19077,N_18204,N_18238);
or U19078 (N_19078,N_18747,N_18794);
xor U19079 (N_19079,N_18865,N_18347);
or U19080 (N_19080,N_18183,N_18116);
nand U19081 (N_19081,N_18135,N_18788);
and U19082 (N_19082,N_18811,N_18274);
and U19083 (N_19083,N_18068,N_18041);
xnor U19084 (N_19084,N_18367,N_18224);
nor U19085 (N_19085,N_18958,N_18692);
nand U19086 (N_19086,N_18668,N_18278);
or U19087 (N_19087,N_18674,N_18524);
or U19088 (N_19088,N_18381,N_18779);
xnor U19089 (N_19089,N_18291,N_18269);
and U19090 (N_19090,N_18995,N_18931);
nor U19091 (N_19091,N_18246,N_18629);
xor U19092 (N_19092,N_18409,N_18063);
xor U19093 (N_19093,N_18985,N_18496);
xnor U19094 (N_19094,N_18467,N_18437);
and U19095 (N_19095,N_18431,N_18342);
and U19096 (N_19096,N_18212,N_18088);
nor U19097 (N_19097,N_18994,N_18285);
xnor U19098 (N_19098,N_18435,N_18133);
or U19099 (N_19099,N_18371,N_18632);
or U19100 (N_19100,N_18060,N_18553);
or U19101 (N_19101,N_18677,N_18647);
xor U19102 (N_19102,N_18589,N_18160);
nand U19103 (N_19103,N_18175,N_18741);
xnor U19104 (N_19104,N_18290,N_18432);
nand U19105 (N_19105,N_18265,N_18688);
nand U19106 (N_19106,N_18270,N_18514);
nand U19107 (N_19107,N_18715,N_18430);
or U19108 (N_19108,N_18020,N_18103);
nor U19109 (N_19109,N_18833,N_18608);
nor U19110 (N_19110,N_18028,N_18427);
xnor U19111 (N_19111,N_18187,N_18007);
or U19112 (N_19112,N_18743,N_18536);
and U19113 (N_19113,N_18149,N_18532);
xnor U19114 (N_19114,N_18882,N_18327);
and U19115 (N_19115,N_18878,N_18025);
xor U19116 (N_19116,N_18009,N_18948);
or U19117 (N_19117,N_18875,N_18311);
or U19118 (N_19118,N_18037,N_18722);
nor U19119 (N_19119,N_18971,N_18112);
xnor U19120 (N_19120,N_18652,N_18602);
or U19121 (N_19121,N_18221,N_18502);
or U19122 (N_19122,N_18551,N_18157);
and U19123 (N_19123,N_18475,N_18406);
nor U19124 (N_19124,N_18719,N_18303);
nand U19125 (N_19125,N_18261,N_18784);
nand U19126 (N_19126,N_18200,N_18911);
xor U19127 (N_19127,N_18313,N_18772);
xor U19128 (N_19128,N_18237,N_18974);
and U19129 (N_19129,N_18820,N_18073);
xnor U19130 (N_19130,N_18873,N_18705);
nand U19131 (N_19131,N_18669,N_18869);
xor U19132 (N_19132,N_18798,N_18888);
nor U19133 (N_19133,N_18454,N_18122);
xor U19134 (N_19134,N_18165,N_18205);
and U19135 (N_19135,N_18754,N_18188);
nand U19136 (N_19136,N_18066,N_18918);
and U19137 (N_19137,N_18693,N_18950);
nor U19138 (N_19138,N_18702,N_18466);
nand U19139 (N_19139,N_18726,N_18453);
xor U19140 (N_19140,N_18823,N_18005);
nand U19141 (N_19141,N_18599,N_18541);
nand U19142 (N_19142,N_18846,N_18544);
xnor U19143 (N_19143,N_18198,N_18736);
or U19144 (N_19144,N_18312,N_18003);
or U19145 (N_19145,N_18986,N_18540);
and U19146 (N_19146,N_18307,N_18642);
nand U19147 (N_19147,N_18095,N_18712);
xnor U19148 (N_19148,N_18843,N_18130);
xor U19149 (N_19149,N_18315,N_18960);
xnor U19150 (N_19150,N_18395,N_18970);
nand U19151 (N_19151,N_18796,N_18979);
xor U19152 (N_19152,N_18929,N_18460);
xnor U19153 (N_19153,N_18508,N_18185);
and U19154 (N_19154,N_18244,N_18389);
nor U19155 (N_19155,N_18145,N_18127);
and U19156 (N_19156,N_18818,N_18203);
xnor U19157 (N_19157,N_18548,N_18412);
nor U19158 (N_19158,N_18740,N_18047);
and U19159 (N_19159,N_18486,N_18152);
or U19160 (N_19160,N_18546,N_18644);
nand U19161 (N_19161,N_18413,N_18525);
or U19162 (N_19162,N_18424,N_18567);
and U19163 (N_19163,N_18163,N_18756);
nand U19164 (N_19164,N_18090,N_18049);
or U19165 (N_19165,N_18055,N_18015);
nand U19166 (N_19166,N_18845,N_18518);
or U19167 (N_19167,N_18338,N_18176);
or U19168 (N_19168,N_18038,N_18337);
xor U19169 (N_19169,N_18639,N_18917);
or U19170 (N_19170,N_18118,N_18761);
nand U19171 (N_19171,N_18834,N_18537);
nand U19172 (N_19172,N_18295,N_18492);
xnor U19173 (N_19173,N_18355,N_18792);
and U19174 (N_19174,N_18026,N_18297);
nor U19175 (N_19175,N_18708,N_18247);
or U19176 (N_19176,N_18399,N_18353);
and U19177 (N_19177,N_18581,N_18832);
and U19178 (N_19178,N_18117,N_18509);
or U19179 (N_19179,N_18036,N_18206);
or U19180 (N_19180,N_18275,N_18617);
or U19181 (N_19181,N_18051,N_18331);
nor U19182 (N_19182,N_18572,N_18704);
nor U19183 (N_19183,N_18790,N_18984);
and U19184 (N_19184,N_18753,N_18364);
and U19185 (N_19185,N_18472,N_18397);
xnor U19186 (N_19186,N_18128,N_18126);
xor U19187 (N_19187,N_18325,N_18650);
or U19188 (N_19188,N_18665,N_18429);
or U19189 (N_19189,N_18672,N_18698);
nand U19190 (N_19190,N_18636,N_18942);
xor U19191 (N_19191,N_18421,N_18294);
xnor U19192 (N_19192,N_18619,N_18083);
xor U19193 (N_19193,N_18844,N_18615);
nand U19194 (N_19194,N_18787,N_18292);
xor U19195 (N_19195,N_18797,N_18012);
nor U19196 (N_19196,N_18027,N_18791);
or U19197 (N_19197,N_18387,N_18143);
nand U19198 (N_19198,N_18543,N_18951);
xnor U19199 (N_19199,N_18515,N_18684);
or U19200 (N_19200,N_18962,N_18123);
or U19201 (N_19201,N_18124,N_18085);
nand U19202 (N_19202,N_18605,N_18763);
nand U19203 (N_19203,N_18059,N_18941);
xor U19204 (N_19204,N_18193,N_18768);
nor U19205 (N_19205,N_18053,N_18657);
nor U19206 (N_19206,N_18630,N_18363);
nor U19207 (N_19207,N_18168,N_18344);
or U19208 (N_19208,N_18745,N_18309);
and U19209 (N_19209,N_18534,N_18923);
or U19210 (N_19210,N_18945,N_18411);
nor U19211 (N_19211,N_18241,N_18717);
nand U19212 (N_19212,N_18132,N_18887);
xnor U19213 (N_19213,N_18861,N_18925);
nand U19214 (N_19214,N_18500,N_18856);
or U19215 (N_19215,N_18765,N_18729);
and U19216 (N_19216,N_18439,N_18946);
xnor U19217 (N_19217,N_18607,N_18280);
nor U19218 (N_19218,N_18370,N_18598);
xor U19219 (N_19219,N_18057,N_18461);
nand U19220 (N_19220,N_18651,N_18405);
and U19221 (N_19221,N_18147,N_18318);
nor U19222 (N_19222,N_18192,N_18326);
xnor U19223 (N_19223,N_18585,N_18474);
and U19224 (N_19224,N_18273,N_18368);
nor U19225 (N_19225,N_18268,N_18759);
nand U19226 (N_19226,N_18664,N_18162);
and U19227 (N_19227,N_18530,N_18554);
xor U19228 (N_19228,N_18732,N_18279);
nor U19229 (N_19229,N_18462,N_18209);
nand U19230 (N_19230,N_18335,N_18125);
or U19231 (N_19231,N_18891,N_18504);
or U19232 (N_19232,N_18358,N_18281);
xnor U19233 (N_19233,N_18750,N_18816);
and U19234 (N_19234,N_18383,N_18838);
and U19235 (N_19235,N_18104,N_18529);
and U19236 (N_19236,N_18803,N_18040);
or U19237 (N_19237,N_18735,N_18023);
nand U19238 (N_19238,N_18054,N_18709);
nand U19239 (N_19239,N_18182,N_18746);
nor U19240 (N_19240,N_18757,N_18662);
or U19241 (N_19241,N_18716,N_18385);
nand U19242 (N_19242,N_18559,N_18822);
or U19243 (N_19243,N_18079,N_18660);
or U19244 (N_19244,N_18513,N_18703);
or U19245 (N_19245,N_18904,N_18912);
nor U19246 (N_19246,N_18349,N_18631);
xor U19247 (N_19247,N_18582,N_18226);
xor U19248 (N_19248,N_18417,N_18254);
and U19249 (N_19249,N_18718,N_18839);
nor U19250 (N_19250,N_18458,N_18233);
nand U19251 (N_19251,N_18785,N_18485);
and U19252 (N_19252,N_18483,N_18978);
or U19253 (N_19253,N_18568,N_18760);
nand U19254 (N_19254,N_18682,N_18077);
nor U19255 (N_19255,N_18635,N_18600);
and U19256 (N_19256,N_18637,N_18356);
and U19257 (N_19257,N_18293,N_18755);
nor U19258 (N_19258,N_18640,N_18499);
and U19259 (N_19259,N_18523,N_18369);
nand U19260 (N_19260,N_18230,N_18024);
xor U19261 (N_19261,N_18783,N_18829);
xnor U19262 (N_19262,N_18841,N_18584);
nor U19263 (N_19263,N_18730,N_18552);
xnor U19264 (N_19264,N_18115,N_18479);
nor U19265 (N_19265,N_18905,N_18093);
xor U19266 (N_19266,N_18403,N_18299);
and U19267 (N_19267,N_18837,N_18645);
and U19268 (N_19268,N_18679,N_18910);
nor U19269 (N_19269,N_18884,N_18813);
nor U19270 (N_19270,N_18098,N_18638);
nand U19271 (N_19271,N_18864,N_18058);
nor U19272 (N_19272,N_18934,N_18778);
xor U19273 (N_19273,N_18310,N_18256);
or U19274 (N_19274,N_18400,N_18334);
xor U19275 (N_19275,N_18604,N_18505);
and U19276 (N_19276,N_18388,N_18721);
nor U19277 (N_19277,N_18129,N_18391);
and U19278 (N_19278,N_18915,N_18266);
and U19279 (N_19279,N_18465,N_18676);
or U19280 (N_19280,N_18916,N_18196);
nor U19281 (N_19281,N_18900,N_18214);
nand U19282 (N_19282,N_18136,N_18180);
or U19283 (N_19283,N_18476,N_18056);
xor U19284 (N_19284,N_18949,N_18179);
xor U19285 (N_19285,N_18450,N_18287);
or U19286 (N_19286,N_18284,N_18243);
and U19287 (N_19287,N_18520,N_18592);
nand U19288 (N_19288,N_18789,N_18578);
nand U19289 (N_19289,N_18586,N_18404);
nor U19290 (N_19290,N_18574,N_18566);
nor U19291 (N_19291,N_18814,N_18913);
nor U19292 (N_19292,N_18232,N_18306);
and U19293 (N_19293,N_18195,N_18621);
nand U19294 (N_19294,N_18097,N_18922);
and U19295 (N_19295,N_18296,N_18376);
nor U19296 (N_19296,N_18469,N_18957);
and U19297 (N_19297,N_18609,N_18625);
nor U19298 (N_19298,N_18542,N_18624);
nand U19299 (N_19299,N_18549,N_18550);
nor U19300 (N_19300,N_18859,N_18382);
nor U19301 (N_19301,N_18392,N_18341);
and U19302 (N_19302,N_18881,N_18197);
and U19303 (N_19303,N_18350,N_18151);
or U19304 (N_19304,N_18332,N_18497);
nand U19305 (N_19305,N_18410,N_18561);
or U19306 (N_19306,N_18419,N_18105);
or U19307 (N_19307,N_18210,N_18422);
or U19308 (N_19308,N_18689,N_18239);
and U19309 (N_19309,N_18262,N_18992);
and U19310 (N_19310,N_18092,N_18277);
or U19311 (N_19311,N_18671,N_18426);
xor U19312 (N_19312,N_18898,N_18622);
nand U19313 (N_19313,N_18614,N_18366);
xor U19314 (N_19314,N_18216,N_18952);
nand U19315 (N_19315,N_18830,N_18987);
or U19316 (N_19316,N_18706,N_18894);
nand U19317 (N_19317,N_18111,N_18648);
xor U19318 (N_19318,N_18854,N_18826);
or U19319 (N_19319,N_18042,N_18414);
or U19320 (N_19320,N_18641,N_18289);
nand U19321 (N_19321,N_18806,N_18091);
or U19322 (N_19322,N_18288,N_18935);
nand U19323 (N_19323,N_18828,N_18250);
nand U19324 (N_19324,N_18490,N_18667);
nor U19325 (N_19325,N_18456,N_18448);
xor U19326 (N_19326,N_18680,N_18597);
xnor U19327 (N_19327,N_18506,N_18876);
xor U19328 (N_19328,N_18078,N_18446);
and U19329 (N_19329,N_18860,N_18831);
and U19330 (N_19330,N_18441,N_18863);
or U19331 (N_19331,N_18357,N_18119);
and U19332 (N_19332,N_18069,N_18626);
or U19333 (N_19333,N_18628,N_18455);
nor U19334 (N_19334,N_18522,N_18777);
or U19335 (N_19335,N_18685,N_18981);
nand U19336 (N_19336,N_18658,N_18897);
nand U19337 (N_19337,N_18780,N_18220);
or U19338 (N_19338,N_18360,N_18560);
or U19339 (N_19339,N_18258,N_18620);
nor U19340 (N_19340,N_18611,N_18045);
xnor U19341 (N_19341,N_18947,N_18144);
and U19342 (N_19342,N_18333,N_18590);
nand U19343 (N_19343,N_18351,N_18425);
nand U19344 (N_19344,N_18562,N_18231);
nor U19345 (N_19345,N_18606,N_18033);
nand U19346 (N_19346,N_18802,N_18603);
nor U19347 (N_19347,N_18800,N_18336);
and U19348 (N_19348,N_18723,N_18393);
and U19349 (N_19349,N_18171,N_18106);
and U19350 (N_19350,N_18993,N_18997);
and U19351 (N_19351,N_18415,N_18016);
xnor U19352 (N_19352,N_18996,N_18362);
and U19353 (N_19353,N_18695,N_18174);
xor U19354 (N_19354,N_18065,N_18048);
nand U19355 (N_19355,N_18418,N_18159);
nor U19356 (N_19356,N_18967,N_18480);
nor U19357 (N_19357,N_18008,N_18074);
xor U19358 (N_19358,N_18234,N_18096);
nand U19359 (N_19359,N_18707,N_18075);
xnor U19360 (N_19360,N_18440,N_18194);
or U19361 (N_19361,N_18473,N_18956);
nor U19362 (N_19362,N_18963,N_18444);
xnor U19363 (N_19363,N_18700,N_18694);
or U19364 (N_19364,N_18965,N_18451);
or U19365 (N_19365,N_18208,N_18725);
nor U19366 (N_19366,N_18742,N_18583);
xor U19367 (N_19367,N_18852,N_18892);
nor U19368 (N_19368,N_18394,N_18793);
nor U19369 (N_19369,N_18298,N_18491);
and U19370 (N_19370,N_18804,N_18673);
or U19371 (N_19371,N_18021,N_18557);
nor U19372 (N_19372,N_18001,N_18002);
nand U19373 (N_19373,N_18764,N_18434);
nand U19374 (N_19374,N_18324,N_18442);
or U19375 (N_19375,N_18384,N_18086);
and U19376 (N_19376,N_18850,N_18516);
and U19377 (N_19377,N_18352,N_18100);
or U19378 (N_19378,N_18148,N_18720);
and U19379 (N_19379,N_18771,N_18980);
and U19380 (N_19380,N_18302,N_18932);
xnor U19381 (N_19381,N_18319,N_18728);
nor U19382 (N_19382,N_18821,N_18201);
or U19383 (N_19383,N_18330,N_18587);
nor U19384 (N_19384,N_18697,N_18178);
and U19385 (N_19385,N_18375,N_18314);
xnor U19386 (N_19386,N_18084,N_18235);
xnor U19387 (N_19387,N_18478,N_18767);
or U19388 (N_19388,N_18308,N_18000);
or U19389 (N_19389,N_18108,N_18908);
xnor U19390 (N_19390,N_18138,N_18769);
xnor U19391 (N_19391,N_18748,N_18373);
or U19392 (N_19392,N_18207,N_18018);
nor U19393 (N_19393,N_18099,N_18052);
and U19394 (N_19394,N_18420,N_18227);
and U19395 (N_19395,N_18801,N_18983);
xnor U19396 (N_19396,N_18731,N_18390);
nand U19397 (N_19397,N_18022,N_18202);
nor U19398 (N_19398,N_18795,N_18445);
xnor U19399 (N_19399,N_18749,N_18489);
and U19400 (N_19400,N_18998,N_18305);
nor U19401 (N_19401,N_18737,N_18436);
or U19402 (N_19402,N_18189,N_18482);
xor U19403 (N_19403,N_18346,N_18217);
and U19404 (N_19404,N_18857,N_18263);
or U19405 (N_19405,N_18902,N_18457);
or U19406 (N_19406,N_18612,N_18646);
xnor U19407 (N_19407,N_18067,N_18862);
nor U19408 (N_19408,N_18866,N_18379);
xor U19409 (N_19409,N_18627,N_18853);
and U19410 (N_19410,N_18339,N_18484);
nor U19411 (N_19411,N_18773,N_18851);
xor U19412 (N_19412,N_18883,N_18519);
xor U19413 (N_19413,N_18172,N_18733);
and U19414 (N_19414,N_18255,N_18538);
or U19415 (N_19415,N_18855,N_18893);
nor U19416 (N_19416,N_18102,N_18249);
and U19417 (N_19417,N_18847,N_18259);
and U19418 (N_19418,N_18988,N_18670);
or U19419 (N_19419,N_18329,N_18153);
nand U19420 (N_19420,N_18190,N_18141);
xor U19421 (N_19421,N_18966,N_18374);
or U19422 (N_19422,N_18493,N_18776);
nor U19423 (N_19423,N_18013,N_18526);
and U19424 (N_19424,N_18173,N_18361);
xnor U19425 (N_19425,N_18588,N_18240);
or U19426 (N_19426,N_18030,N_18799);
and U19427 (N_19427,N_18260,N_18751);
or U19428 (N_19428,N_18903,N_18477);
nand U19429 (N_19429,N_18359,N_18569);
nand U19430 (N_19430,N_18573,N_18150);
and U19431 (N_19431,N_18634,N_18398);
nand U19432 (N_19432,N_18964,N_18345);
xor U19433 (N_19433,N_18253,N_18070);
xor U19434 (N_19434,N_18062,N_18807);
xnor U19435 (N_19435,N_18889,N_18954);
xnor U19436 (N_19436,N_18481,N_18675);
and U19437 (N_19437,N_18936,N_18975);
nand U19438 (N_19438,N_18304,N_18999);
xnor U19439 (N_19439,N_18545,N_18953);
nor U19440 (N_19440,N_18170,N_18976);
xnor U19441 (N_19441,N_18681,N_18004);
and U19442 (N_19442,N_18081,N_18501);
nor U19443 (N_19443,N_18710,N_18937);
nand U19444 (N_19444,N_18181,N_18940);
and U19445 (N_19445,N_18471,N_18575);
xor U19446 (N_19446,N_18046,N_18527);
nand U19447 (N_19447,N_18378,N_18050);
xor U19448 (N_19448,N_18019,N_18613);
and U19449 (N_19449,N_18973,N_18396);
and U19450 (N_19450,N_18082,N_18271);
or U19451 (N_19451,N_18167,N_18895);
or U19452 (N_19452,N_18035,N_18380);
nand U19453 (N_19453,N_18094,N_18158);
nor U19454 (N_19454,N_18690,N_18139);
nor U19455 (N_19455,N_18576,N_18968);
nand U19456 (N_19456,N_18156,N_18186);
and U19457 (N_19457,N_18087,N_18563);
nor U19458 (N_19458,N_18595,N_18463);
xor U19459 (N_19459,N_18565,N_18533);
and U19460 (N_19460,N_18034,N_18245);
and U19461 (N_19461,N_18556,N_18257);
and U19462 (N_19462,N_18555,N_18871);
nand U19463 (N_19463,N_18758,N_18468);
xnor U19464 (N_19464,N_18666,N_18977);
or U19465 (N_19465,N_18252,N_18317);
and U19466 (N_19466,N_18011,N_18452);
nand U19467 (N_19467,N_18114,N_18017);
nand U19468 (N_19468,N_18282,N_18762);
xor U19469 (N_19469,N_18817,N_18089);
nand U19470 (N_19470,N_18539,N_18494);
and U19471 (N_19471,N_18061,N_18618);
and U19472 (N_19472,N_18354,N_18039);
or U19473 (N_19473,N_18827,N_18535);
nand U19474 (N_19474,N_18840,N_18914);
nand U19475 (N_19475,N_18076,N_18229);
nand U19476 (N_19476,N_18770,N_18032);
nand U19477 (N_19477,N_18781,N_18320);
nor U19478 (N_19478,N_18107,N_18447);
xnor U19479 (N_19479,N_18459,N_18649);
nor U19480 (N_19480,N_18242,N_18464);
nor U19481 (N_19481,N_18926,N_18683);
and U19482 (N_19482,N_18879,N_18433);
or U19483 (N_19483,N_18301,N_18678);
nor U19484 (N_19484,N_18236,N_18877);
xor U19485 (N_19485,N_18836,N_18408);
nor U19486 (N_19486,N_18223,N_18933);
or U19487 (N_19487,N_18990,N_18443);
xnor U19488 (N_19488,N_18029,N_18901);
xor U19489 (N_19489,N_18824,N_18164);
xor U19490 (N_19490,N_18848,N_18121);
xor U19491 (N_19491,N_18842,N_18580);
and U19492 (N_19492,N_18316,N_18043);
and U19493 (N_19493,N_18924,N_18727);
xor U19494 (N_19494,N_18531,N_18283);
nand U19495 (N_19495,N_18633,N_18014);
and U19496 (N_19496,N_18517,N_18939);
nor U19497 (N_19497,N_18503,N_18696);
nor U19498 (N_19498,N_18177,N_18225);
nand U19499 (N_19499,N_18215,N_18510);
or U19500 (N_19500,N_18469,N_18317);
xnor U19501 (N_19501,N_18659,N_18058);
nand U19502 (N_19502,N_18756,N_18831);
nor U19503 (N_19503,N_18156,N_18387);
nor U19504 (N_19504,N_18375,N_18786);
nor U19505 (N_19505,N_18014,N_18835);
nor U19506 (N_19506,N_18747,N_18754);
nor U19507 (N_19507,N_18106,N_18134);
nand U19508 (N_19508,N_18132,N_18660);
nor U19509 (N_19509,N_18588,N_18529);
nand U19510 (N_19510,N_18624,N_18636);
or U19511 (N_19511,N_18585,N_18546);
nand U19512 (N_19512,N_18406,N_18089);
or U19513 (N_19513,N_18056,N_18118);
and U19514 (N_19514,N_18431,N_18678);
nand U19515 (N_19515,N_18758,N_18092);
xnor U19516 (N_19516,N_18485,N_18107);
or U19517 (N_19517,N_18332,N_18295);
nor U19518 (N_19518,N_18190,N_18753);
nor U19519 (N_19519,N_18743,N_18346);
or U19520 (N_19520,N_18343,N_18718);
xnor U19521 (N_19521,N_18428,N_18455);
nor U19522 (N_19522,N_18253,N_18210);
nor U19523 (N_19523,N_18051,N_18255);
or U19524 (N_19524,N_18524,N_18041);
or U19525 (N_19525,N_18071,N_18904);
nand U19526 (N_19526,N_18439,N_18773);
and U19527 (N_19527,N_18831,N_18225);
and U19528 (N_19528,N_18094,N_18789);
nor U19529 (N_19529,N_18483,N_18045);
and U19530 (N_19530,N_18014,N_18850);
nand U19531 (N_19531,N_18591,N_18428);
xor U19532 (N_19532,N_18177,N_18344);
nand U19533 (N_19533,N_18387,N_18896);
and U19534 (N_19534,N_18121,N_18174);
xnor U19535 (N_19535,N_18336,N_18121);
and U19536 (N_19536,N_18455,N_18815);
nor U19537 (N_19537,N_18045,N_18222);
nand U19538 (N_19538,N_18570,N_18523);
and U19539 (N_19539,N_18786,N_18129);
and U19540 (N_19540,N_18847,N_18129);
xor U19541 (N_19541,N_18199,N_18489);
nand U19542 (N_19542,N_18750,N_18961);
and U19543 (N_19543,N_18867,N_18720);
nand U19544 (N_19544,N_18263,N_18117);
nor U19545 (N_19545,N_18409,N_18297);
and U19546 (N_19546,N_18149,N_18590);
xor U19547 (N_19547,N_18028,N_18823);
xnor U19548 (N_19548,N_18234,N_18556);
or U19549 (N_19549,N_18462,N_18432);
xor U19550 (N_19550,N_18963,N_18238);
and U19551 (N_19551,N_18887,N_18880);
nand U19552 (N_19552,N_18897,N_18789);
xnor U19553 (N_19553,N_18264,N_18472);
nor U19554 (N_19554,N_18680,N_18539);
or U19555 (N_19555,N_18643,N_18012);
nor U19556 (N_19556,N_18497,N_18205);
nand U19557 (N_19557,N_18742,N_18978);
xnor U19558 (N_19558,N_18517,N_18096);
nor U19559 (N_19559,N_18738,N_18139);
and U19560 (N_19560,N_18031,N_18085);
nand U19561 (N_19561,N_18458,N_18699);
nand U19562 (N_19562,N_18676,N_18887);
xor U19563 (N_19563,N_18031,N_18400);
or U19564 (N_19564,N_18388,N_18806);
nand U19565 (N_19565,N_18319,N_18005);
nand U19566 (N_19566,N_18595,N_18695);
and U19567 (N_19567,N_18561,N_18610);
nand U19568 (N_19568,N_18960,N_18086);
nand U19569 (N_19569,N_18159,N_18091);
and U19570 (N_19570,N_18435,N_18388);
and U19571 (N_19571,N_18957,N_18345);
or U19572 (N_19572,N_18976,N_18897);
xor U19573 (N_19573,N_18853,N_18016);
nand U19574 (N_19574,N_18683,N_18057);
nand U19575 (N_19575,N_18331,N_18261);
or U19576 (N_19576,N_18282,N_18334);
and U19577 (N_19577,N_18056,N_18027);
or U19578 (N_19578,N_18658,N_18372);
nor U19579 (N_19579,N_18554,N_18031);
nand U19580 (N_19580,N_18846,N_18537);
nor U19581 (N_19581,N_18857,N_18838);
and U19582 (N_19582,N_18536,N_18444);
nand U19583 (N_19583,N_18317,N_18107);
nand U19584 (N_19584,N_18170,N_18002);
nor U19585 (N_19585,N_18880,N_18204);
nor U19586 (N_19586,N_18591,N_18021);
or U19587 (N_19587,N_18976,N_18952);
and U19588 (N_19588,N_18033,N_18452);
nand U19589 (N_19589,N_18116,N_18933);
nand U19590 (N_19590,N_18345,N_18491);
nand U19591 (N_19591,N_18380,N_18065);
nand U19592 (N_19592,N_18024,N_18135);
and U19593 (N_19593,N_18644,N_18302);
nand U19594 (N_19594,N_18676,N_18184);
nor U19595 (N_19595,N_18490,N_18101);
nor U19596 (N_19596,N_18686,N_18716);
and U19597 (N_19597,N_18152,N_18327);
and U19598 (N_19598,N_18777,N_18400);
and U19599 (N_19599,N_18324,N_18645);
nor U19600 (N_19600,N_18361,N_18293);
nand U19601 (N_19601,N_18838,N_18812);
or U19602 (N_19602,N_18593,N_18961);
nand U19603 (N_19603,N_18907,N_18454);
and U19604 (N_19604,N_18041,N_18179);
and U19605 (N_19605,N_18809,N_18994);
and U19606 (N_19606,N_18317,N_18225);
nor U19607 (N_19607,N_18280,N_18791);
and U19608 (N_19608,N_18192,N_18459);
nand U19609 (N_19609,N_18306,N_18104);
nand U19610 (N_19610,N_18512,N_18414);
xor U19611 (N_19611,N_18836,N_18076);
or U19612 (N_19612,N_18674,N_18067);
and U19613 (N_19613,N_18547,N_18470);
or U19614 (N_19614,N_18270,N_18306);
nor U19615 (N_19615,N_18615,N_18232);
or U19616 (N_19616,N_18873,N_18341);
xnor U19617 (N_19617,N_18590,N_18888);
xor U19618 (N_19618,N_18974,N_18344);
and U19619 (N_19619,N_18662,N_18205);
nor U19620 (N_19620,N_18961,N_18519);
nor U19621 (N_19621,N_18086,N_18565);
nor U19622 (N_19622,N_18932,N_18900);
nand U19623 (N_19623,N_18634,N_18160);
or U19624 (N_19624,N_18765,N_18202);
xnor U19625 (N_19625,N_18519,N_18612);
or U19626 (N_19626,N_18617,N_18259);
and U19627 (N_19627,N_18794,N_18242);
and U19628 (N_19628,N_18359,N_18278);
xnor U19629 (N_19629,N_18873,N_18477);
xor U19630 (N_19630,N_18751,N_18872);
nand U19631 (N_19631,N_18589,N_18305);
or U19632 (N_19632,N_18554,N_18463);
nand U19633 (N_19633,N_18328,N_18532);
and U19634 (N_19634,N_18020,N_18373);
nand U19635 (N_19635,N_18406,N_18016);
or U19636 (N_19636,N_18331,N_18120);
nor U19637 (N_19637,N_18513,N_18794);
and U19638 (N_19638,N_18543,N_18589);
nor U19639 (N_19639,N_18767,N_18138);
nand U19640 (N_19640,N_18061,N_18066);
nor U19641 (N_19641,N_18941,N_18780);
and U19642 (N_19642,N_18199,N_18028);
and U19643 (N_19643,N_18761,N_18289);
or U19644 (N_19644,N_18336,N_18470);
and U19645 (N_19645,N_18108,N_18797);
or U19646 (N_19646,N_18753,N_18810);
xnor U19647 (N_19647,N_18451,N_18951);
xor U19648 (N_19648,N_18272,N_18714);
nor U19649 (N_19649,N_18855,N_18782);
nand U19650 (N_19650,N_18879,N_18851);
xor U19651 (N_19651,N_18640,N_18510);
xor U19652 (N_19652,N_18848,N_18915);
and U19653 (N_19653,N_18617,N_18944);
and U19654 (N_19654,N_18971,N_18587);
and U19655 (N_19655,N_18506,N_18058);
or U19656 (N_19656,N_18786,N_18854);
nor U19657 (N_19657,N_18408,N_18994);
nand U19658 (N_19658,N_18550,N_18274);
or U19659 (N_19659,N_18422,N_18500);
xor U19660 (N_19660,N_18751,N_18020);
nor U19661 (N_19661,N_18617,N_18274);
xor U19662 (N_19662,N_18136,N_18149);
nor U19663 (N_19663,N_18895,N_18455);
nand U19664 (N_19664,N_18626,N_18255);
nand U19665 (N_19665,N_18962,N_18561);
and U19666 (N_19666,N_18838,N_18394);
or U19667 (N_19667,N_18604,N_18454);
or U19668 (N_19668,N_18592,N_18394);
nor U19669 (N_19669,N_18593,N_18861);
nor U19670 (N_19670,N_18035,N_18145);
nor U19671 (N_19671,N_18788,N_18594);
nor U19672 (N_19672,N_18434,N_18678);
and U19673 (N_19673,N_18078,N_18366);
or U19674 (N_19674,N_18864,N_18701);
nand U19675 (N_19675,N_18274,N_18377);
nor U19676 (N_19676,N_18821,N_18433);
and U19677 (N_19677,N_18118,N_18409);
xnor U19678 (N_19678,N_18027,N_18766);
or U19679 (N_19679,N_18569,N_18036);
or U19680 (N_19680,N_18363,N_18316);
nand U19681 (N_19681,N_18997,N_18731);
nor U19682 (N_19682,N_18414,N_18169);
xor U19683 (N_19683,N_18786,N_18151);
or U19684 (N_19684,N_18952,N_18625);
nand U19685 (N_19685,N_18721,N_18481);
or U19686 (N_19686,N_18161,N_18121);
nor U19687 (N_19687,N_18520,N_18926);
xor U19688 (N_19688,N_18867,N_18594);
or U19689 (N_19689,N_18294,N_18042);
or U19690 (N_19690,N_18181,N_18910);
and U19691 (N_19691,N_18188,N_18116);
nor U19692 (N_19692,N_18782,N_18941);
nor U19693 (N_19693,N_18704,N_18413);
and U19694 (N_19694,N_18582,N_18384);
and U19695 (N_19695,N_18108,N_18075);
or U19696 (N_19696,N_18204,N_18825);
and U19697 (N_19697,N_18080,N_18272);
or U19698 (N_19698,N_18692,N_18984);
and U19699 (N_19699,N_18294,N_18116);
xnor U19700 (N_19700,N_18605,N_18112);
xor U19701 (N_19701,N_18072,N_18589);
nor U19702 (N_19702,N_18168,N_18357);
and U19703 (N_19703,N_18351,N_18538);
xnor U19704 (N_19704,N_18827,N_18430);
xor U19705 (N_19705,N_18857,N_18545);
or U19706 (N_19706,N_18215,N_18028);
and U19707 (N_19707,N_18960,N_18276);
and U19708 (N_19708,N_18239,N_18347);
xnor U19709 (N_19709,N_18603,N_18448);
or U19710 (N_19710,N_18867,N_18553);
nand U19711 (N_19711,N_18396,N_18518);
xor U19712 (N_19712,N_18587,N_18029);
or U19713 (N_19713,N_18476,N_18829);
nand U19714 (N_19714,N_18851,N_18067);
nor U19715 (N_19715,N_18283,N_18060);
or U19716 (N_19716,N_18469,N_18164);
nand U19717 (N_19717,N_18428,N_18852);
or U19718 (N_19718,N_18852,N_18184);
xnor U19719 (N_19719,N_18799,N_18262);
or U19720 (N_19720,N_18766,N_18912);
or U19721 (N_19721,N_18708,N_18689);
and U19722 (N_19722,N_18004,N_18398);
and U19723 (N_19723,N_18377,N_18265);
xnor U19724 (N_19724,N_18271,N_18236);
nand U19725 (N_19725,N_18639,N_18753);
or U19726 (N_19726,N_18497,N_18087);
nand U19727 (N_19727,N_18100,N_18454);
nor U19728 (N_19728,N_18644,N_18980);
nand U19729 (N_19729,N_18268,N_18162);
nand U19730 (N_19730,N_18498,N_18402);
xnor U19731 (N_19731,N_18757,N_18390);
and U19732 (N_19732,N_18870,N_18193);
nor U19733 (N_19733,N_18453,N_18703);
xnor U19734 (N_19734,N_18363,N_18529);
nand U19735 (N_19735,N_18061,N_18702);
nand U19736 (N_19736,N_18068,N_18356);
nor U19737 (N_19737,N_18214,N_18534);
nand U19738 (N_19738,N_18783,N_18465);
xnor U19739 (N_19739,N_18000,N_18250);
nor U19740 (N_19740,N_18954,N_18971);
or U19741 (N_19741,N_18152,N_18792);
xnor U19742 (N_19742,N_18757,N_18642);
nor U19743 (N_19743,N_18711,N_18342);
xnor U19744 (N_19744,N_18574,N_18788);
nor U19745 (N_19745,N_18364,N_18309);
or U19746 (N_19746,N_18751,N_18779);
xor U19747 (N_19747,N_18817,N_18242);
nor U19748 (N_19748,N_18382,N_18874);
nor U19749 (N_19749,N_18571,N_18449);
and U19750 (N_19750,N_18663,N_18622);
nand U19751 (N_19751,N_18028,N_18963);
xor U19752 (N_19752,N_18101,N_18169);
nor U19753 (N_19753,N_18204,N_18026);
nand U19754 (N_19754,N_18783,N_18716);
or U19755 (N_19755,N_18733,N_18437);
xor U19756 (N_19756,N_18879,N_18994);
nor U19757 (N_19757,N_18409,N_18489);
and U19758 (N_19758,N_18372,N_18375);
nor U19759 (N_19759,N_18141,N_18227);
or U19760 (N_19760,N_18674,N_18244);
or U19761 (N_19761,N_18755,N_18647);
and U19762 (N_19762,N_18042,N_18093);
xnor U19763 (N_19763,N_18008,N_18211);
nor U19764 (N_19764,N_18075,N_18142);
or U19765 (N_19765,N_18062,N_18877);
and U19766 (N_19766,N_18222,N_18282);
nand U19767 (N_19767,N_18662,N_18968);
nand U19768 (N_19768,N_18237,N_18813);
and U19769 (N_19769,N_18926,N_18644);
and U19770 (N_19770,N_18689,N_18491);
nand U19771 (N_19771,N_18342,N_18321);
xor U19772 (N_19772,N_18467,N_18523);
nand U19773 (N_19773,N_18246,N_18181);
and U19774 (N_19774,N_18967,N_18569);
xnor U19775 (N_19775,N_18629,N_18637);
xnor U19776 (N_19776,N_18498,N_18698);
nand U19777 (N_19777,N_18582,N_18267);
or U19778 (N_19778,N_18823,N_18510);
xnor U19779 (N_19779,N_18488,N_18670);
xor U19780 (N_19780,N_18763,N_18522);
and U19781 (N_19781,N_18483,N_18347);
xnor U19782 (N_19782,N_18554,N_18791);
nand U19783 (N_19783,N_18487,N_18226);
xnor U19784 (N_19784,N_18941,N_18411);
and U19785 (N_19785,N_18563,N_18905);
or U19786 (N_19786,N_18595,N_18399);
or U19787 (N_19787,N_18083,N_18769);
and U19788 (N_19788,N_18515,N_18484);
and U19789 (N_19789,N_18496,N_18739);
nand U19790 (N_19790,N_18038,N_18974);
or U19791 (N_19791,N_18629,N_18702);
nand U19792 (N_19792,N_18342,N_18030);
nor U19793 (N_19793,N_18946,N_18367);
and U19794 (N_19794,N_18881,N_18994);
nand U19795 (N_19795,N_18791,N_18615);
xor U19796 (N_19796,N_18310,N_18677);
nor U19797 (N_19797,N_18021,N_18560);
nand U19798 (N_19798,N_18026,N_18696);
nor U19799 (N_19799,N_18648,N_18346);
xnor U19800 (N_19800,N_18232,N_18385);
and U19801 (N_19801,N_18869,N_18160);
xnor U19802 (N_19802,N_18940,N_18558);
nor U19803 (N_19803,N_18948,N_18019);
or U19804 (N_19804,N_18583,N_18631);
nor U19805 (N_19805,N_18012,N_18547);
xor U19806 (N_19806,N_18480,N_18839);
nand U19807 (N_19807,N_18167,N_18689);
nor U19808 (N_19808,N_18287,N_18672);
or U19809 (N_19809,N_18518,N_18411);
and U19810 (N_19810,N_18941,N_18207);
and U19811 (N_19811,N_18851,N_18086);
and U19812 (N_19812,N_18538,N_18929);
or U19813 (N_19813,N_18351,N_18757);
and U19814 (N_19814,N_18775,N_18830);
nor U19815 (N_19815,N_18975,N_18163);
nand U19816 (N_19816,N_18678,N_18205);
or U19817 (N_19817,N_18432,N_18324);
nor U19818 (N_19818,N_18598,N_18456);
or U19819 (N_19819,N_18055,N_18120);
and U19820 (N_19820,N_18503,N_18954);
nor U19821 (N_19821,N_18158,N_18176);
nor U19822 (N_19822,N_18309,N_18586);
xnor U19823 (N_19823,N_18572,N_18072);
and U19824 (N_19824,N_18163,N_18780);
nand U19825 (N_19825,N_18978,N_18907);
nor U19826 (N_19826,N_18332,N_18711);
nor U19827 (N_19827,N_18902,N_18575);
or U19828 (N_19828,N_18999,N_18927);
or U19829 (N_19829,N_18378,N_18196);
or U19830 (N_19830,N_18660,N_18011);
xnor U19831 (N_19831,N_18813,N_18390);
nand U19832 (N_19832,N_18067,N_18848);
and U19833 (N_19833,N_18074,N_18025);
and U19834 (N_19834,N_18369,N_18996);
nand U19835 (N_19835,N_18871,N_18107);
xor U19836 (N_19836,N_18890,N_18326);
or U19837 (N_19837,N_18399,N_18123);
nand U19838 (N_19838,N_18201,N_18097);
or U19839 (N_19839,N_18282,N_18927);
xnor U19840 (N_19840,N_18878,N_18200);
nor U19841 (N_19841,N_18966,N_18023);
or U19842 (N_19842,N_18040,N_18655);
or U19843 (N_19843,N_18923,N_18630);
nor U19844 (N_19844,N_18297,N_18267);
xnor U19845 (N_19845,N_18630,N_18108);
nor U19846 (N_19846,N_18565,N_18456);
or U19847 (N_19847,N_18983,N_18255);
nand U19848 (N_19848,N_18081,N_18593);
xnor U19849 (N_19849,N_18983,N_18604);
or U19850 (N_19850,N_18573,N_18590);
and U19851 (N_19851,N_18045,N_18993);
nor U19852 (N_19852,N_18354,N_18615);
nor U19853 (N_19853,N_18163,N_18746);
nand U19854 (N_19854,N_18290,N_18595);
xor U19855 (N_19855,N_18990,N_18079);
nand U19856 (N_19856,N_18575,N_18156);
xor U19857 (N_19857,N_18288,N_18734);
and U19858 (N_19858,N_18370,N_18708);
nand U19859 (N_19859,N_18562,N_18552);
nor U19860 (N_19860,N_18228,N_18719);
nand U19861 (N_19861,N_18396,N_18202);
and U19862 (N_19862,N_18137,N_18586);
and U19863 (N_19863,N_18945,N_18307);
xor U19864 (N_19864,N_18767,N_18852);
nand U19865 (N_19865,N_18889,N_18885);
and U19866 (N_19866,N_18992,N_18113);
or U19867 (N_19867,N_18168,N_18359);
xnor U19868 (N_19868,N_18473,N_18484);
nand U19869 (N_19869,N_18119,N_18507);
or U19870 (N_19870,N_18042,N_18298);
or U19871 (N_19871,N_18425,N_18438);
or U19872 (N_19872,N_18878,N_18976);
nand U19873 (N_19873,N_18814,N_18733);
nor U19874 (N_19874,N_18080,N_18414);
or U19875 (N_19875,N_18422,N_18651);
nor U19876 (N_19876,N_18726,N_18097);
and U19877 (N_19877,N_18093,N_18881);
and U19878 (N_19878,N_18884,N_18181);
nand U19879 (N_19879,N_18344,N_18594);
nor U19880 (N_19880,N_18602,N_18370);
nand U19881 (N_19881,N_18307,N_18014);
nor U19882 (N_19882,N_18560,N_18477);
xnor U19883 (N_19883,N_18229,N_18256);
or U19884 (N_19884,N_18059,N_18777);
nand U19885 (N_19885,N_18309,N_18189);
and U19886 (N_19886,N_18407,N_18677);
and U19887 (N_19887,N_18802,N_18803);
or U19888 (N_19888,N_18551,N_18268);
nand U19889 (N_19889,N_18545,N_18906);
and U19890 (N_19890,N_18437,N_18001);
nand U19891 (N_19891,N_18152,N_18368);
and U19892 (N_19892,N_18804,N_18684);
and U19893 (N_19893,N_18319,N_18626);
nor U19894 (N_19894,N_18446,N_18957);
nand U19895 (N_19895,N_18206,N_18220);
xnor U19896 (N_19896,N_18880,N_18396);
or U19897 (N_19897,N_18012,N_18787);
nand U19898 (N_19898,N_18507,N_18700);
xor U19899 (N_19899,N_18110,N_18591);
xnor U19900 (N_19900,N_18841,N_18448);
nor U19901 (N_19901,N_18242,N_18688);
nor U19902 (N_19902,N_18927,N_18546);
nand U19903 (N_19903,N_18154,N_18727);
and U19904 (N_19904,N_18363,N_18613);
or U19905 (N_19905,N_18291,N_18964);
nor U19906 (N_19906,N_18726,N_18101);
nor U19907 (N_19907,N_18459,N_18455);
nor U19908 (N_19908,N_18643,N_18642);
and U19909 (N_19909,N_18191,N_18691);
and U19910 (N_19910,N_18450,N_18368);
nor U19911 (N_19911,N_18970,N_18310);
or U19912 (N_19912,N_18032,N_18752);
nand U19913 (N_19913,N_18479,N_18837);
or U19914 (N_19914,N_18643,N_18856);
nand U19915 (N_19915,N_18988,N_18190);
nor U19916 (N_19916,N_18262,N_18001);
and U19917 (N_19917,N_18667,N_18525);
nor U19918 (N_19918,N_18992,N_18055);
nor U19919 (N_19919,N_18382,N_18544);
nand U19920 (N_19920,N_18323,N_18804);
nor U19921 (N_19921,N_18779,N_18281);
xnor U19922 (N_19922,N_18642,N_18630);
xnor U19923 (N_19923,N_18846,N_18857);
xor U19924 (N_19924,N_18450,N_18082);
nand U19925 (N_19925,N_18549,N_18682);
nand U19926 (N_19926,N_18541,N_18300);
xor U19927 (N_19927,N_18761,N_18846);
nand U19928 (N_19928,N_18453,N_18622);
and U19929 (N_19929,N_18570,N_18677);
and U19930 (N_19930,N_18220,N_18232);
or U19931 (N_19931,N_18602,N_18390);
and U19932 (N_19932,N_18309,N_18370);
or U19933 (N_19933,N_18357,N_18054);
and U19934 (N_19934,N_18597,N_18050);
nand U19935 (N_19935,N_18485,N_18495);
and U19936 (N_19936,N_18573,N_18605);
nor U19937 (N_19937,N_18373,N_18841);
xnor U19938 (N_19938,N_18661,N_18107);
nor U19939 (N_19939,N_18401,N_18248);
and U19940 (N_19940,N_18754,N_18406);
nor U19941 (N_19941,N_18903,N_18021);
or U19942 (N_19942,N_18511,N_18769);
xor U19943 (N_19943,N_18652,N_18861);
nand U19944 (N_19944,N_18018,N_18638);
or U19945 (N_19945,N_18676,N_18898);
or U19946 (N_19946,N_18457,N_18474);
xor U19947 (N_19947,N_18900,N_18258);
and U19948 (N_19948,N_18215,N_18935);
xor U19949 (N_19949,N_18985,N_18600);
or U19950 (N_19950,N_18377,N_18591);
and U19951 (N_19951,N_18474,N_18149);
nor U19952 (N_19952,N_18690,N_18904);
nand U19953 (N_19953,N_18817,N_18456);
or U19954 (N_19954,N_18700,N_18666);
nand U19955 (N_19955,N_18331,N_18630);
nor U19956 (N_19956,N_18870,N_18298);
nand U19957 (N_19957,N_18660,N_18975);
nor U19958 (N_19958,N_18486,N_18894);
nor U19959 (N_19959,N_18548,N_18612);
nor U19960 (N_19960,N_18901,N_18441);
nand U19961 (N_19961,N_18231,N_18826);
and U19962 (N_19962,N_18026,N_18010);
or U19963 (N_19963,N_18353,N_18169);
nor U19964 (N_19964,N_18588,N_18673);
nor U19965 (N_19965,N_18650,N_18946);
or U19966 (N_19966,N_18089,N_18341);
nand U19967 (N_19967,N_18117,N_18630);
and U19968 (N_19968,N_18674,N_18834);
nor U19969 (N_19969,N_18878,N_18543);
nor U19970 (N_19970,N_18238,N_18617);
xnor U19971 (N_19971,N_18848,N_18563);
xor U19972 (N_19972,N_18131,N_18443);
nor U19973 (N_19973,N_18031,N_18889);
xor U19974 (N_19974,N_18164,N_18623);
xor U19975 (N_19975,N_18552,N_18024);
nor U19976 (N_19976,N_18223,N_18548);
or U19977 (N_19977,N_18278,N_18674);
or U19978 (N_19978,N_18134,N_18498);
nor U19979 (N_19979,N_18183,N_18062);
nand U19980 (N_19980,N_18732,N_18208);
nand U19981 (N_19981,N_18270,N_18050);
nand U19982 (N_19982,N_18114,N_18462);
xnor U19983 (N_19983,N_18081,N_18648);
and U19984 (N_19984,N_18284,N_18872);
and U19985 (N_19985,N_18625,N_18011);
nor U19986 (N_19986,N_18147,N_18353);
nand U19987 (N_19987,N_18649,N_18312);
and U19988 (N_19988,N_18780,N_18829);
or U19989 (N_19989,N_18438,N_18987);
and U19990 (N_19990,N_18392,N_18580);
nand U19991 (N_19991,N_18038,N_18065);
or U19992 (N_19992,N_18795,N_18272);
nor U19993 (N_19993,N_18618,N_18814);
nand U19994 (N_19994,N_18221,N_18007);
and U19995 (N_19995,N_18674,N_18134);
nor U19996 (N_19996,N_18522,N_18252);
nand U19997 (N_19997,N_18973,N_18529);
and U19998 (N_19998,N_18956,N_18874);
nor U19999 (N_19999,N_18030,N_18532);
xor U20000 (N_20000,N_19647,N_19682);
xnor U20001 (N_20001,N_19156,N_19997);
xor U20002 (N_20002,N_19972,N_19629);
nand U20003 (N_20003,N_19628,N_19265);
or U20004 (N_20004,N_19613,N_19644);
and U20005 (N_20005,N_19425,N_19221);
nor U20006 (N_20006,N_19488,N_19732);
xnor U20007 (N_20007,N_19711,N_19392);
and U20008 (N_20008,N_19479,N_19961);
xor U20009 (N_20009,N_19181,N_19755);
nor U20010 (N_20010,N_19578,N_19417);
and U20011 (N_20011,N_19552,N_19528);
and U20012 (N_20012,N_19693,N_19905);
nor U20013 (N_20013,N_19975,N_19505);
nand U20014 (N_20014,N_19098,N_19184);
and U20015 (N_20015,N_19455,N_19390);
xnor U20016 (N_20016,N_19757,N_19564);
nor U20017 (N_20017,N_19470,N_19426);
and U20018 (N_20018,N_19190,N_19193);
nor U20019 (N_20019,N_19700,N_19590);
xor U20020 (N_20020,N_19224,N_19679);
nand U20021 (N_20021,N_19307,N_19282);
or U20022 (N_20022,N_19041,N_19527);
nor U20023 (N_20023,N_19668,N_19883);
nand U20024 (N_20024,N_19441,N_19101);
nand U20025 (N_20025,N_19968,N_19896);
nor U20026 (N_20026,N_19115,N_19235);
or U20027 (N_20027,N_19990,N_19234);
or U20028 (N_20028,N_19168,N_19855);
xor U20029 (N_20029,N_19080,N_19678);
nand U20030 (N_20030,N_19219,N_19302);
xor U20031 (N_20031,N_19976,N_19494);
and U20032 (N_20032,N_19481,N_19349);
or U20033 (N_20033,N_19919,N_19113);
xnor U20034 (N_20034,N_19588,N_19183);
nor U20035 (N_20035,N_19770,N_19971);
or U20036 (N_20036,N_19801,N_19795);
xnor U20037 (N_20037,N_19671,N_19416);
nor U20038 (N_20038,N_19877,N_19172);
or U20039 (N_20039,N_19926,N_19938);
and U20040 (N_20040,N_19012,N_19903);
nand U20041 (N_20041,N_19987,N_19818);
xnor U20042 (N_20042,N_19743,N_19677);
or U20043 (N_20043,N_19728,N_19431);
nand U20044 (N_20044,N_19822,N_19558);
nor U20045 (N_20045,N_19222,N_19240);
nor U20046 (N_20046,N_19639,N_19914);
or U20047 (N_20047,N_19662,N_19969);
xnor U20048 (N_20048,N_19418,N_19446);
xnor U20049 (N_20049,N_19496,N_19097);
nor U20050 (N_20050,N_19011,N_19889);
or U20051 (N_20051,N_19828,N_19544);
and U20052 (N_20052,N_19137,N_19329);
xor U20053 (N_20053,N_19726,N_19569);
and U20054 (N_20054,N_19218,N_19359);
xor U20055 (N_20055,N_19545,N_19956);
and U20056 (N_20056,N_19324,N_19145);
or U20057 (N_20057,N_19264,N_19055);
nor U20058 (N_20058,N_19207,N_19806);
nor U20059 (N_20059,N_19109,N_19713);
nor U20060 (N_20060,N_19745,N_19958);
xnor U20061 (N_20061,N_19461,N_19784);
xnor U20062 (N_20062,N_19837,N_19939);
xor U20063 (N_20063,N_19381,N_19986);
and U20064 (N_20064,N_19999,N_19489);
nand U20065 (N_20065,N_19735,N_19869);
xor U20066 (N_20066,N_19340,N_19909);
nor U20067 (N_20067,N_19402,N_19936);
nor U20068 (N_20068,N_19005,N_19327);
xor U20069 (N_20069,N_19454,N_19541);
xnor U20070 (N_20070,N_19059,N_19686);
and U20071 (N_20071,N_19208,N_19261);
nand U20072 (N_20072,N_19079,N_19603);
nand U20073 (N_20073,N_19439,N_19925);
nand U20074 (N_20074,N_19258,N_19514);
and U20075 (N_20075,N_19309,N_19203);
or U20076 (N_20076,N_19281,N_19069);
or U20077 (N_20077,N_19038,N_19014);
nand U20078 (N_20078,N_19852,N_19305);
or U20079 (N_20079,N_19952,N_19210);
or U20080 (N_20080,N_19449,N_19045);
or U20081 (N_20081,N_19907,N_19859);
xnor U20082 (N_20082,N_19636,N_19260);
nor U20083 (N_20083,N_19949,N_19804);
xnor U20084 (N_20084,N_19727,N_19741);
xor U20085 (N_20085,N_19230,N_19314);
nor U20086 (N_20086,N_19651,N_19681);
xor U20087 (N_20087,N_19597,N_19067);
xor U20088 (N_20088,N_19459,N_19729);
or U20089 (N_20089,N_19540,N_19092);
and U20090 (N_20090,N_19810,N_19974);
nor U20091 (N_20091,N_19391,N_19592);
nor U20092 (N_20092,N_19823,N_19860);
xor U20093 (N_20093,N_19180,N_19328);
nand U20094 (N_20094,N_19771,N_19880);
or U20095 (N_20095,N_19484,N_19007);
nand U20096 (N_20096,N_19389,N_19312);
nand U20097 (N_20097,N_19388,N_19731);
nor U20098 (N_20098,N_19114,N_19386);
and U20099 (N_20099,N_19557,N_19518);
xor U20100 (N_20100,N_19075,N_19460);
and U20101 (N_20101,N_19608,N_19593);
and U20102 (N_20102,N_19847,N_19829);
nand U20103 (N_20103,N_19794,N_19138);
and U20104 (N_20104,N_19524,N_19946);
or U20105 (N_20105,N_19397,N_19793);
nor U20106 (N_20106,N_19815,N_19501);
nand U20107 (N_20107,N_19692,N_19150);
xor U20108 (N_20108,N_19135,N_19212);
nand U20109 (N_20109,N_19303,N_19842);
nand U20110 (N_20110,N_19627,N_19421);
nor U20111 (N_20111,N_19044,N_19228);
and U20112 (N_20112,N_19062,N_19637);
and U20113 (N_20113,N_19875,N_19699);
and U20114 (N_20114,N_19087,N_19957);
or U20115 (N_20115,N_19188,N_19768);
nand U20116 (N_20116,N_19853,N_19435);
xor U20117 (N_20117,N_19635,N_19520);
nand U20118 (N_20118,N_19658,N_19262);
nor U20119 (N_20119,N_19756,N_19963);
nor U20120 (N_20120,N_19721,N_19638);
nor U20121 (N_20121,N_19398,N_19737);
or U20122 (N_20122,N_19531,N_19760);
and U20123 (N_20123,N_19424,N_19444);
and U20124 (N_20124,N_19291,N_19186);
nand U20125 (N_20125,N_19684,N_19707);
nand U20126 (N_20126,N_19015,N_19959);
and U20127 (N_20127,N_19318,N_19201);
or U20128 (N_20128,N_19767,N_19788);
and U20129 (N_20129,N_19802,N_19916);
or U20130 (N_20130,N_19888,N_19551);
nor U20131 (N_20131,N_19370,N_19565);
nor U20132 (N_20132,N_19615,N_19632);
and U20133 (N_20133,N_19123,N_19226);
and U20134 (N_20134,N_19498,N_19348);
nand U20135 (N_20135,N_19690,N_19490);
xnor U20136 (N_20136,N_19994,N_19511);
nand U20137 (N_20137,N_19238,N_19442);
xnor U20138 (N_20138,N_19373,N_19865);
nand U20139 (N_20139,N_19029,N_19427);
xnor U20140 (N_20140,N_19010,N_19472);
nor U20141 (N_20141,N_19004,N_19364);
and U20142 (N_20142,N_19266,N_19019);
nor U20143 (N_20143,N_19550,N_19278);
and U20144 (N_20144,N_19675,N_19652);
xnor U20145 (N_20145,N_19073,N_19716);
or U20146 (N_20146,N_19002,N_19749);
and U20147 (N_20147,N_19081,N_19500);
nor U20148 (N_20148,N_19811,N_19898);
xor U20149 (N_20149,N_19338,N_19153);
xnor U20150 (N_20150,N_19169,N_19339);
nand U20151 (N_20151,N_19509,N_19433);
or U20152 (N_20152,N_19857,N_19131);
nor U20153 (N_20153,N_19213,N_19249);
xnor U20154 (N_20154,N_19485,N_19543);
or U20155 (N_20155,N_19927,N_19600);
xnor U20156 (N_20156,N_19724,N_19667);
or U20157 (N_20157,N_19561,N_19341);
nor U20158 (N_20158,N_19214,N_19110);
nor U20159 (N_20159,N_19812,N_19506);
xnor U20160 (N_20160,N_19033,N_19351);
nand U20161 (N_20161,N_19893,N_19523);
xor U20162 (N_20162,N_19753,N_19962);
nor U20163 (N_20163,N_19432,N_19546);
xnor U20164 (N_20164,N_19268,N_19654);
or U20165 (N_20165,N_19709,N_19199);
nor U20166 (N_20166,N_19864,N_19814);
and U20167 (N_20167,N_19585,N_19083);
xnor U20168 (N_20168,N_19429,N_19923);
nand U20169 (N_20169,N_19185,N_19094);
nor U20170 (N_20170,N_19532,N_19039);
and U20171 (N_20171,N_19293,N_19861);
xnor U20172 (N_20172,N_19453,N_19866);
nor U20173 (N_20173,N_19154,N_19099);
or U20174 (N_20174,N_19664,N_19191);
or U20175 (N_20175,N_19817,N_19910);
xor U20176 (N_20176,N_19360,N_19367);
xor U20177 (N_20177,N_19085,N_19515);
nor U20178 (N_20178,N_19512,N_19572);
or U20179 (N_20179,N_19774,N_19609);
xor U20180 (N_20180,N_19171,N_19142);
xor U20181 (N_20181,N_19161,N_19813);
xnor U20182 (N_20182,N_19537,N_19782);
and U20183 (N_20183,N_19510,N_19881);
and U20184 (N_20184,N_19820,N_19072);
or U20185 (N_20185,N_19844,N_19406);
or U20186 (N_20186,N_19900,N_19495);
xor U20187 (N_20187,N_19042,N_19366);
or U20188 (N_20188,N_19194,N_19430);
nand U20189 (N_20189,N_19502,N_19250);
and U20190 (N_20190,N_19216,N_19619);
and U20191 (N_20191,N_19606,N_19006);
xnor U20192 (N_20192,N_19833,N_19492);
nand U20193 (N_20193,N_19434,N_19333);
xnor U20194 (N_20194,N_19953,N_19577);
or U20195 (N_20195,N_19259,N_19915);
xor U20196 (N_20196,N_19934,N_19263);
and U20197 (N_20197,N_19803,N_19626);
xor U20198 (N_20198,N_19122,N_19955);
nor U20199 (N_20199,N_19000,N_19315);
nor U20200 (N_20200,N_19840,N_19533);
xor U20201 (N_20201,N_19850,N_19854);
and U20202 (N_20202,N_19691,N_19596);
or U20203 (N_20203,N_19331,N_19311);
or U20204 (N_20204,N_19912,N_19808);
or U20205 (N_20205,N_19977,N_19362);
nand U20206 (N_20206,N_19361,N_19908);
or U20207 (N_20207,N_19831,N_19383);
and U20208 (N_20208,N_19008,N_19462);
or U20209 (N_20209,N_19395,N_19027);
nor U20210 (N_20210,N_19750,N_19384);
and U20211 (N_20211,N_19165,N_19605);
nor U20212 (N_20212,N_19878,N_19559);
xor U20213 (N_20213,N_19584,N_19661);
xor U20214 (N_20214,N_19103,N_19330);
or U20215 (N_20215,N_19720,N_19870);
nand U20216 (N_20216,N_19074,N_19299);
xnor U20217 (N_20217,N_19689,N_19112);
or U20218 (N_20218,N_19825,N_19428);
or U20219 (N_20219,N_19068,N_19197);
nand U20220 (N_20220,N_19891,N_19960);
nand U20221 (N_20221,N_19796,N_19215);
or U20222 (N_20222,N_19239,N_19271);
nor U20223 (N_20223,N_19316,N_19294);
xnor U20224 (N_20224,N_19733,N_19924);
nor U20225 (N_20225,N_19344,N_19769);
and U20226 (N_20226,N_19522,N_19136);
and U20227 (N_20227,N_19321,N_19176);
xnor U20228 (N_20228,N_19155,N_19369);
or U20229 (N_20229,N_19827,N_19978);
and U20230 (N_20230,N_19173,N_19824);
nor U20231 (N_20231,N_19941,N_19104);
nor U20232 (N_20232,N_19504,N_19223);
or U20233 (N_20233,N_19775,N_19942);
xor U20234 (N_20234,N_19162,N_19674);
nand U20235 (N_20235,N_19473,N_19935);
nor U20236 (N_20236,N_19621,N_19283);
or U20237 (N_20237,N_19887,N_19149);
nand U20238 (N_20238,N_19687,N_19277);
xnor U20239 (N_20239,N_19175,N_19279);
nor U20240 (N_20240,N_19762,N_19051);
and U20241 (N_20241,N_19730,N_19843);
nor U20242 (N_20242,N_19576,N_19879);
and U20243 (N_20243,N_19868,N_19355);
and U20244 (N_20244,N_19497,N_19319);
or U20245 (N_20245,N_19483,N_19940);
nand U20246 (N_20246,N_19529,N_19419);
nor U20247 (N_20247,N_19121,N_19867);
and U20248 (N_20248,N_19676,N_19673);
nand U20249 (N_20249,N_19983,N_19998);
or U20250 (N_20250,N_19412,N_19013);
xnor U20251 (N_20251,N_19451,N_19407);
nand U20252 (N_20252,N_19284,N_19777);
xnor U20253 (N_20253,N_19920,N_19408);
and U20254 (N_20254,N_19040,N_19158);
and U20255 (N_20255,N_19922,N_19320);
xor U20256 (N_20256,N_19740,N_19107);
nand U20257 (N_20257,N_19555,N_19017);
and U20258 (N_20258,N_19030,N_19243);
and U20259 (N_20259,N_19096,N_19611);
xor U20260 (N_20260,N_19198,N_19549);
nand U20261 (N_20261,N_19140,N_19393);
nor U20262 (N_20262,N_19672,N_19575);
and U20263 (N_20263,N_19163,N_19405);
xor U20264 (N_20264,N_19885,N_19049);
or U20265 (N_20265,N_19325,N_19272);
and U20266 (N_20266,N_19710,N_19274);
and U20267 (N_20267,N_19164,N_19241);
or U20268 (N_20268,N_19290,N_19703);
nand U20269 (N_20269,N_19144,N_19624);
xnor U20270 (N_20270,N_19179,N_19301);
nand U20271 (N_20271,N_19064,N_19300);
or U20272 (N_20272,N_19404,N_19932);
nor U20273 (N_20273,N_19656,N_19884);
nand U20274 (N_20274,N_19317,N_19723);
nor U20275 (N_20275,N_19758,N_19894);
xnor U20276 (N_20276,N_19143,N_19187);
and U20277 (N_20277,N_19102,N_19694);
and U20278 (N_20278,N_19669,N_19204);
xnor U20279 (N_20279,N_19964,N_19789);
nor U20280 (N_20280,N_19902,N_19933);
or U20281 (N_20281,N_19088,N_19126);
nor U20282 (N_20282,N_19587,N_19759);
and U20283 (N_20283,N_19438,N_19437);
and U20284 (N_20284,N_19071,N_19643);
nand U20285 (N_20285,N_19225,N_19851);
xnor U20286 (N_20286,N_19151,N_19568);
or U20287 (N_20287,N_19931,N_19413);
xor U20288 (N_20288,N_19217,N_19354);
or U20289 (N_20289,N_19744,N_19560);
or U20290 (N_20290,N_19090,N_19356);
nand U20291 (N_20291,N_19048,N_19233);
nor U20292 (N_20292,N_19025,N_19474);
or U20293 (N_20293,N_19345,N_19132);
nand U20294 (N_20294,N_19835,N_19979);
xor U20295 (N_20295,N_19120,N_19748);
or U20296 (N_20296,N_19763,N_19834);
and U20297 (N_20297,N_19640,N_19372);
nand U20298 (N_20298,N_19513,N_19872);
or U20299 (N_20299,N_19895,N_19486);
or U20300 (N_20300,N_19819,N_19385);
or U20301 (N_20301,N_19477,N_19981);
and U20302 (N_20302,N_19607,N_19414);
xnor U20303 (N_20303,N_19623,N_19781);
and U20304 (N_20304,N_19751,N_19701);
xnor U20305 (N_20305,N_19858,N_19047);
nor U20306 (N_20306,N_19022,N_19897);
nor U20307 (N_20307,N_19848,N_19196);
and U20308 (N_20308,N_19993,N_19086);
xor U20309 (N_20309,N_19091,N_19947);
xnor U20310 (N_20310,N_19053,N_19747);
or U20311 (N_20311,N_19415,N_19401);
or U20312 (N_20312,N_19009,N_19516);
nor U20313 (N_20313,N_19147,N_19447);
and U20314 (N_20314,N_19660,N_19400);
nor U20315 (N_20315,N_19874,N_19378);
nor U20316 (N_20316,N_19773,N_19478);
and U20317 (N_20317,N_19780,N_19704);
or U20318 (N_20318,N_19705,N_19892);
xor U20319 (N_20319,N_19482,N_19111);
or U20320 (N_20320,N_19467,N_19023);
nor U20321 (N_20321,N_19056,N_19464);
nand U20322 (N_20322,N_19313,N_19698);
nor U20323 (N_20323,N_19616,N_19280);
xnor U20324 (N_20324,N_19521,N_19948);
xnor U20325 (N_20325,N_19070,N_19342);
nor U20326 (N_20326,N_19128,N_19786);
nand U20327 (N_20327,N_19396,N_19166);
or U20328 (N_20328,N_19670,N_19177);
nand U20329 (N_20329,N_19253,N_19346);
nand U20330 (N_20330,N_19211,N_19448);
or U20331 (N_20331,N_19680,N_19178);
nand U20332 (N_20332,N_19754,N_19645);
nand U20333 (N_20333,N_19571,N_19800);
nand U20334 (N_20334,N_19420,N_19967);
nor U20335 (N_20335,N_19141,N_19170);
xnor U20336 (N_20336,N_19220,N_19985);
nor U20337 (N_20337,N_19856,N_19581);
and U20338 (N_20338,N_19547,N_19347);
xor U20339 (N_20339,N_19057,N_19242);
xor U20340 (N_20340,N_19236,N_19129);
nand U20341 (N_20341,N_19245,N_19246);
nor U20342 (N_20342,N_19772,N_19821);
xor U20343 (N_20343,N_19832,N_19655);
nand U20344 (N_20344,N_19950,N_19054);
and U20345 (N_20345,N_19846,N_19805);
and U20346 (N_20346,N_19970,N_19783);
xnor U20347 (N_20347,N_19237,N_19599);
nand U20348 (N_20348,N_19463,N_19625);
xnor U20349 (N_20349,N_19648,N_19422);
and U20350 (N_20350,N_19838,N_19901);
or U20351 (N_20351,N_19229,N_19715);
xnor U20352 (N_20352,N_19989,N_19286);
xnor U20353 (N_20353,N_19016,N_19357);
and U20354 (N_20354,N_19231,N_19612);
or U20355 (N_20355,N_19563,N_19598);
nand U20356 (N_20356,N_19060,N_19882);
nand U20357 (N_20357,N_19666,N_19918);
nand U20358 (N_20358,N_19046,N_19382);
or U20359 (N_20359,N_19148,N_19548);
and U20360 (N_20360,N_19269,N_19984);
and U20361 (N_20361,N_19065,N_19334);
xor U20362 (N_20362,N_19954,N_19873);
nand U20363 (N_20363,N_19790,N_19380);
nor U20364 (N_20364,N_19117,N_19980);
and U20365 (N_20365,N_19586,N_19917);
nor U20366 (N_20366,N_19717,N_19913);
or U20367 (N_20367,N_19475,N_19343);
xnor U20368 (N_20368,N_19517,N_19742);
xnor U20369 (N_20369,N_19020,N_19335);
and U20370 (N_20370,N_19232,N_19403);
xor U20371 (N_20371,N_19061,N_19287);
nand U20372 (N_20372,N_19849,N_19116);
and U20373 (N_20373,N_19244,N_19399);
nand U20374 (N_20374,N_19695,N_19118);
xor U20375 (N_20375,N_19336,N_19580);
nor U20376 (N_20376,N_19778,N_19195);
xnor U20377 (N_20377,N_19379,N_19119);
nor U20378 (N_20378,N_19063,N_19582);
xnor U20379 (N_20379,N_19659,N_19125);
and U20380 (N_20380,N_19440,N_19539);
nor U20381 (N_20381,N_19275,N_19082);
and U20382 (N_20382,N_19052,N_19363);
and U20383 (N_20383,N_19839,N_19298);
xor U20384 (N_20384,N_19722,N_19556);
nand U20385 (N_20385,N_19604,N_19043);
nor U20386 (N_20386,N_19100,N_19465);
or U20387 (N_20387,N_19270,N_19982);
xor U20388 (N_20388,N_19152,N_19944);
nor U20389 (N_20389,N_19276,N_19003);
nor U20390 (N_20390,N_19683,N_19567);
nor U20391 (N_20391,N_19653,N_19937);
nor U20392 (N_20392,N_19921,N_19766);
xor U20393 (N_20393,N_19876,N_19257);
nand U20394 (N_20394,N_19610,N_19579);
nand U20395 (N_20395,N_19322,N_19594);
xnor U20396 (N_20396,N_19765,N_19525);
and U20397 (N_20397,N_19458,N_19353);
nand U20398 (N_20398,N_19738,N_19174);
and U20399 (N_20399,N_19992,N_19066);
nand U20400 (N_20400,N_19863,N_19295);
or U20401 (N_20401,N_19157,N_19256);
xnor U20402 (N_20402,N_19836,N_19306);
xor U20403 (N_20403,N_19566,N_19034);
nand U20404 (N_20404,N_19706,N_19929);
xor U20405 (N_20405,N_19452,N_19206);
or U20406 (N_20406,N_19714,N_19945);
nand U20407 (N_20407,N_19791,N_19906);
nand U20408 (N_20408,N_19991,N_19375);
nand U20409 (N_20409,N_19764,N_19487);
xor U20410 (N_20410,N_19423,N_19205);
nand U20411 (N_20411,N_19718,N_19337);
nor U20412 (N_20412,N_19323,N_19799);
xor U20413 (N_20413,N_19493,N_19622);
xor U20414 (N_20414,N_19614,N_19326);
nand U20415 (N_20415,N_19297,N_19050);
xor U20416 (N_20416,N_19076,N_19292);
xor U20417 (N_20417,N_19503,N_19519);
nor U20418 (N_20418,N_19255,N_19227);
nand U20419 (N_20419,N_19787,N_19641);
or U20420 (N_20420,N_19736,N_19845);
or U20421 (N_20421,N_19209,N_19797);
or U20422 (N_20422,N_19685,N_19352);
nand U20423 (N_20423,N_19037,N_19371);
nand U20424 (N_20424,N_19127,N_19634);
and U20425 (N_20425,N_19776,N_19200);
and U20426 (N_20426,N_19365,N_19089);
nand U20427 (N_20427,N_19332,N_19508);
nand U20428 (N_20428,N_19031,N_19471);
and U20429 (N_20429,N_19024,N_19996);
xor U20430 (N_20430,N_19574,N_19553);
xor U20431 (N_20431,N_19930,N_19308);
xnor U20432 (N_20432,N_19093,N_19965);
or U20433 (N_20433,N_19289,N_19456);
xor U20434 (N_20434,N_19688,N_19871);
or U20435 (N_20435,N_19649,N_19189);
and U20436 (N_20436,N_19443,N_19904);
nor U20437 (N_20437,N_19095,N_19719);
and U20438 (N_20438,N_19663,N_19657);
nand U20439 (N_20439,N_19018,N_19350);
and U20440 (N_20440,N_19591,N_19445);
and U20441 (N_20441,N_19589,N_19146);
nor U20442 (N_20442,N_19450,N_19809);
or U20443 (N_20443,N_19247,N_19077);
nor U20444 (N_20444,N_19358,N_19409);
nand U20445 (N_20445,N_19830,N_19105);
xor U20446 (N_20446,N_19304,N_19001);
nor U20447 (N_20447,N_19374,N_19702);
nand U20448 (N_20448,N_19534,N_19886);
nand U20449 (N_20449,N_19530,N_19583);
and U20450 (N_20450,N_19167,N_19792);
nor U20451 (N_20451,N_19491,N_19890);
and U20452 (N_20452,N_19192,N_19469);
xnor U20453 (N_20453,N_19394,N_19595);
or U20454 (N_20454,N_19841,N_19785);
nor U20455 (N_20455,N_19554,N_19734);
xor U20456 (N_20456,N_19928,N_19028);
and U20457 (N_20457,N_19468,N_19130);
and U20458 (N_20458,N_19480,N_19562);
and U20459 (N_20459,N_19988,N_19032);
nand U20460 (N_20460,N_19570,N_19036);
nand U20461 (N_20461,N_19084,N_19160);
or U20462 (N_20462,N_19712,N_19642);
and U20463 (N_20463,N_19798,N_19725);
or U20464 (N_20464,N_19650,N_19058);
nand U20465 (N_20465,N_19966,N_19526);
nor U20466 (N_20466,N_19746,N_19021);
and U20467 (N_20467,N_19026,N_19368);
and U20468 (N_20468,N_19202,N_19411);
xnor U20469 (N_20469,N_19630,N_19816);
or U20470 (N_20470,N_19752,N_19159);
nand U20471 (N_20471,N_19617,N_19078);
xor U20472 (N_20472,N_19436,N_19133);
xnor U20473 (N_20473,N_19251,N_19285);
xor U20474 (N_20474,N_19807,N_19779);
and U20475 (N_20475,N_19248,N_19862);
nand U20476 (N_20476,N_19601,N_19377);
or U20477 (N_20477,N_19310,N_19108);
nand U20478 (N_20478,N_19254,N_19252);
xor U20479 (N_20479,N_19646,N_19182);
nand U20480 (N_20480,N_19134,N_19457);
or U20481 (N_20481,N_19124,N_19911);
and U20482 (N_20482,N_19633,N_19573);
nand U20483 (N_20483,N_19973,N_19538);
and U20484 (N_20484,N_19995,N_19739);
nand U20485 (N_20485,N_19387,N_19708);
and U20486 (N_20486,N_19620,N_19697);
nand U20487 (N_20487,N_19535,N_19542);
or U20488 (N_20488,N_19631,N_19106);
or U20489 (N_20489,N_19507,N_19296);
nand U20490 (N_20490,N_19665,N_19536);
xnor U20491 (N_20491,N_19602,N_19035);
or U20492 (N_20492,N_19267,N_19951);
nand U20493 (N_20493,N_19139,N_19466);
or U20494 (N_20494,N_19288,N_19618);
or U20495 (N_20495,N_19376,N_19761);
nor U20496 (N_20496,N_19273,N_19826);
nand U20497 (N_20497,N_19410,N_19499);
nor U20498 (N_20498,N_19476,N_19696);
nand U20499 (N_20499,N_19899,N_19943);
xnor U20500 (N_20500,N_19498,N_19844);
xnor U20501 (N_20501,N_19953,N_19089);
xor U20502 (N_20502,N_19643,N_19655);
xnor U20503 (N_20503,N_19872,N_19193);
or U20504 (N_20504,N_19298,N_19790);
nand U20505 (N_20505,N_19439,N_19849);
nand U20506 (N_20506,N_19089,N_19710);
nor U20507 (N_20507,N_19801,N_19490);
nand U20508 (N_20508,N_19031,N_19371);
nor U20509 (N_20509,N_19028,N_19472);
xor U20510 (N_20510,N_19222,N_19723);
and U20511 (N_20511,N_19476,N_19395);
nand U20512 (N_20512,N_19938,N_19324);
nand U20513 (N_20513,N_19353,N_19404);
xnor U20514 (N_20514,N_19817,N_19201);
nand U20515 (N_20515,N_19049,N_19107);
xor U20516 (N_20516,N_19181,N_19891);
and U20517 (N_20517,N_19009,N_19943);
nor U20518 (N_20518,N_19887,N_19187);
nand U20519 (N_20519,N_19324,N_19701);
or U20520 (N_20520,N_19042,N_19390);
nand U20521 (N_20521,N_19387,N_19403);
nor U20522 (N_20522,N_19939,N_19686);
nor U20523 (N_20523,N_19226,N_19573);
nor U20524 (N_20524,N_19913,N_19702);
xor U20525 (N_20525,N_19447,N_19628);
or U20526 (N_20526,N_19095,N_19995);
and U20527 (N_20527,N_19335,N_19235);
nor U20528 (N_20528,N_19765,N_19152);
nor U20529 (N_20529,N_19363,N_19527);
or U20530 (N_20530,N_19621,N_19344);
or U20531 (N_20531,N_19758,N_19070);
nand U20532 (N_20532,N_19361,N_19237);
xor U20533 (N_20533,N_19062,N_19476);
nand U20534 (N_20534,N_19717,N_19768);
or U20535 (N_20535,N_19486,N_19888);
xor U20536 (N_20536,N_19860,N_19585);
xor U20537 (N_20537,N_19507,N_19749);
nor U20538 (N_20538,N_19411,N_19579);
nor U20539 (N_20539,N_19521,N_19250);
or U20540 (N_20540,N_19378,N_19019);
nand U20541 (N_20541,N_19788,N_19104);
xor U20542 (N_20542,N_19427,N_19133);
nor U20543 (N_20543,N_19847,N_19914);
and U20544 (N_20544,N_19662,N_19779);
nand U20545 (N_20545,N_19347,N_19387);
xor U20546 (N_20546,N_19987,N_19455);
and U20547 (N_20547,N_19400,N_19822);
nor U20548 (N_20548,N_19401,N_19823);
nor U20549 (N_20549,N_19811,N_19927);
nor U20550 (N_20550,N_19512,N_19533);
xnor U20551 (N_20551,N_19544,N_19784);
and U20552 (N_20552,N_19950,N_19282);
and U20553 (N_20553,N_19841,N_19771);
nor U20554 (N_20554,N_19607,N_19919);
xor U20555 (N_20555,N_19185,N_19518);
nor U20556 (N_20556,N_19897,N_19995);
and U20557 (N_20557,N_19021,N_19347);
nand U20558 (N_20558,N_19379,N_19538);
or U20559 (N_20559,N_19752,N_19359);
or U20560 (N_20560,N_19151,N_19806);
xor U20561 (N_20561,N_19537,N_19363);
xnor U20562 (N_20562,N_19011,N_19142);
nor U20563 (N_20563,N_19361,N_19021);
or U20564 (N_20564,N_19918,N_19217);
and U20565 (N_20565,N_19978,N_19687);
and U20566 (N_20566,N_19853,N_19590);
nand U20567 (N_20567,N_19160,N_19717);
nand U20568 (N_20568,N_19930,N_19853);
nand U20569 (N_20569,N_19001,N_19428);
nor U20570 (N_20570,N_19651,N_19778);
xor U20571 (N_20571,N_19431,N_19255);
and U20572 (N_20572,N_19785,N_19276);
and U20573 (N_20573,N_19224,N_19241);
nor U20574 (N_20574,N_19259,N_19910);
xnor U20575 (N_20575,N_19467,N_19270);
or U20576 (N_20576,N_19996,N_19145);
xor U20577 (N_20577,N_19685,N_19820);
and U20578 (N_20578,N_19000,N_19186);
nor U20579 (N_20579,N_19368,N_19863);
or U20580 (N_20580,N_19239,N_19228);
nor U20581 (N_20581,N_19056,N_19379);
nor U20582 (N_20582,N_19311,N_19248);
or U20583 (N_20583,N_19925,N_19579);
nand U20584 (N_20584,N_19230,N_19032);
or U20585 (N_20585,N_19205,N_19697);
nand U20586 (N_20586,N_19939,N_19004);
and U20587 (N_20587,N_19171,N_19348);
and U20588 (N_20588,N_19360,N_19571);
xor U20589 (N_20589,N_19906,N_19734);
or U20590 (N_20590,N_19236,N_19738);
and U20591 (N_20591,N_19481,N_19377);
nand U20592 (N_20592,N_19030,N_19242);
nand U20593 (N_20593,N_19152,N_19788);
xnor U20594 (N_20594,N_19503,N_19064);
nand U20595 (N_20595,N_19193,N_19613);
nand U20596 (N_20596,N_19675,N_19097);
nor U20597 (N_20597,N_19321,N_19771);
or U20598 (N_20598,N_19727,N_19859);
nand U20599 (N_20599,N_19842,N_19414);
or U20600 (N_20600,N_19802,N_19427);
nor U20601 (N_20601,N_19692,N_19325);
nor U20602 (N_20602,N_19161,N_19023);
xor U20603 (N_20603,N_19505,N_19297);
and U20604 (N_20604,N_19802,N_19877);
xor U20605 (N_20605,N_19763,N_19096);
nand U20606 (N_20606,N_19039,N_19975);
nor U20607 (N_20607,N_19881,N_19623);
and U20608 (N_20608,N_19451,N_19071);
nor U20609 (N_20609,N_19764,N_19239);
nor U20610 (N_20610,N_19559,N_19182);
nand U20611 (N_20611,N_19739,N_19801);
or U20612 (N_20612,N_19329,N_19126);
xor U20613 (N_20613,N_19754,N_19000);
xor U20614 (N_20614,N_19105,N_19992);
xnor U20615 (N_20615,N_19981,N_19449);
xor U20616 (N_20616,N_19064,N_19919);
xnor U20617 (N_20617,N_19142,N_19445);
xnor U20618 (N_20618,N_19837,N_19980);
or U20619 (N_20619,N_19967,N_19342);
nand U20620 (N_20620,N_19930,N_19914);
xor U20621 (N_20621,N_19465,N_19588);
nor U20622 (N_20622,N_19895,N_19069);
xnor U20623 (N_20623,N_19228,N_19380);
xnor U20624 (N_20624,N_19512,N_19811);
or U20625 (N_20625,N_19528,N_19570);
nor U20626 (N_20626,N_19807,N_19877);
nand U20627 (N_20627,N_19247,N_19842);
nand U20628 (N_20628,N_19955,N_19084);
or U20629 (N_20629,N_19771,N_19764);
and U20630 (N_20630,N_19251,N_19014);
nor U20631 (N_20631,N_19979,N_19475);
nor U20632 (N_20632,N_19426,N_19188);
or U20633 (N_20633,N_19364,N_19750);
nor U20634 (N_20634,N_19815,N_19280);
nand U20635 (N_20635,N_19606,N_19953);
and U20636 (N_20636,N_19646,N_19278);
and U20637 (N_20637,N_19953,N_19910);
or U20638 (N_20638,N_19864,N_19386);
nand U20639 (N_20639,N_19338,N_19330);
nor U20640 (N_20640,N_19808,N_19735);
and U20641 (N_20641,N_19903,N_19401);
or U20642 (N_20642,N_19337,N_19745);
nor U20643 (N_20643,N_19052,N_19535);
nand U20644 (N_20644,N_19306,N_19745);
or U20645 (N_20645,N_19013,N_19572);
xor U20646 (N_20646,N_19799,N_19478);
and U20647 (N_20647,N_19774,N_19210);
nor U20648 (N_20648,N_19977,N_19314);
nand U20649 (N_20649,N_19018,N_19025);
nand U20650 (N_20650,N_19314,N_19491);
xnor U20651 (N_20651,N_19965,N_19450);
nand U20652 (N_20652,N_19537,N_19734);
or U20653 (N_20653,N_19660,N_19437);
nor U20654 (N_20654,N_19757,N_19649);
nand U20655 (N_20655,N_19107,N_19596);
xnor U20656 (N_20656,N_19331,N_19371);
nor U20657 (N_20657,N_19101,N_19633);
nor U20658 (N_20658,N_19310,N_19271);
nor U20659 (N_20659,N_19353,N_19415);
or U20660 (N_20660,N_19080,N_19930);
nor U20661 (N_20661,N_19126,N_19027);
or U20662 (N_20662,N_19548,N_19692);
or U20663 (N_20663,N_19745,N_19555);
nand U20664 (N_20664,N_19210,N_19987);
or U20665 (N_20665,N_19288,N_19743);
nand U20666 (N_20666,N_19643,N_19433);
and U20667 (N_20667,N_19015,N_19407);
or U20668 (N_20668,N_19738,N_19382);
nand U20669 (N_20669,N_19452,N_19909);
xor U20670 (N_20670,N_19992,N_19779);
nand U20671 (N_20671,N_19360,N_19270);
and U20672 (N_20672,N_19737,N_19695);
nor U20673 (N_20673,N_19809,N_19037);
and U20674 (N_20674,N_19284,N_19765);
xor U20675 (N_20675,N_19017,N_19511);
nor U20676 (N_20676,N_19251,N_19576);
or U20677 (N_20677,N_19124,N_19157);
and U20678 (N_20678,N_19664,N_19079);
nor U20679 (N_20679,N_19101,N_19394);
nand U20680 (N_20680,N_19726,N_19148);
nor U20681 (N_20681,N_19216,N_19696);
or U20682 (N_20682,N_19756,N_19370);
and U20683 (N_20683,N_19535,N_19469);
and U20684 (N_20684,N_19476,N_19005);
or U20685 (N_20685,N_19252,N_19684);
nand U20686 (N_20686,N_19989,N_19192);
or U20687 (N_20687,N_19784,N_19536);
and U20688 (N_20688,N_19851,N_19098);
and U20689 (N_20689,N_19028,N_19019);
and U20690 (N_20690,N_19337,N_19184);
and U20691 (N_20691,N_19070,N_19142);
and U20692 (N_20692,N_19331,N_19795);
xnor U20693 (N_20693,N_19079,N_19374);
nor U20694 (N_20694,N_19964,N_19819);
and U20695 (N_20695,N_19730,N_19807);
nor U20696 (N_20696,N_19618,N_19455);
xnor U20697 (N_20697,N_19879,N_19115);
and U20698 (N_20698,N_19471,N_19647);
nand U20699 (N_20699,N_19673,N_19861);
nand U20700 (N_20700,N_19851,N_19215);
nand U20701 (N_20701,N_19506,N_19499);
nor U20702 (N_20702,N_19332,N_19027);
and U20703 (N_20703,N_19099,N_19113);
or U20704 (N_20704,N_19662,N_19915);
nand U20705 (N_20705,N_19816,N_19632);
nor U20706 (N_20706,N_19833,N_19343);
or U20707 (N_20707,N_19100,N_19716);
nand U20708 (N_20708,N_19462,N_19619);
nor U20709 (N_20709,N_19368,N_19859);
or U20710 (N_20710,N_19830,N_19745);
and U20711 (N_20711,N_19639,N_19655);
or U20712 (N_20712,N_19255,N_19828);
and U20713 (N_20713,N_19104,N_19453);
xor U20714 (N_20714,N_19220,N_19111);
and U20715 (N_20715,N_19815,N_19159);
xor U20716 (N_20716,N_19259,N_19295);
nor U20717 (N_20717,N_19076,N_19092);
or U20718 (N_20718,N_19686,N_19135);
and U20719 (N_20719,N_19302,N_19405);
nand U20720 (N_20720,N_19850,N_19759);
and U20721 (N_20721,N_19339,N_19042);
and U20722 (N_20722,N_19052,N_19321);
xnor U20723 (N_20723,N_19862,N_19258);
nor U20724 (N_20724,N_19808,N_19199);
xnor U20725 (N_20725,N_19100,N_19660);
nand U20726 (N_20726,N_19844,N_19843);
or U20727 (N_20727,N_19668,N_19191);
and U20728 (N_20728,N_19111,N_19634);
and U20729 (N_20729,N_19072,N_19661);
and U20730 (N_20730,N_19243,N_19983);
nor U20731 (N_20731,N_19213,N_19606);
or U20732 (N_20732,N_19267,N_19718);
and U20733 (N_20733,N_19215,N_19894);
xnor U20734 (N_20734,N_19144,N_19100);
or U20735 (N_20735,N_19928,N_19585);
and U20736 (N_20736,N_19736,N_19719);
and U20737 (N_20737,N_19752,N_19403);
nor U20738 (N_20738,N_19414,N_19577);
nor U20739 (N_20739,N_19208,N_19031);
or U20740 (N_20740,N_19240,N_19085);
or U20741 (N_20741,N_19260,N_19311);
and U20742 (N_20742,N_19211,N_19775);
nand U20743 (N_20743,N_19928,N_19441);
and U20744 (N_20744,N_19393,N_19351);
nor U20745 (N_20745,N_19177,N_19501);
or U20746 (N_20746,N_19594,N_19161);
nor U20747 (N_20747,N_19247,N_19910);
xor U20748 (N_20748,N_19807,N_19891);
and U20749 (N_20749,N_19542,N_19322);
nor U20750 (N_20750,N_19043,N_19970);
nor U20751 (N_20751,N_19151,N_19720);
nand U20752 (N_20752,N_19501,N_19626);
or U20753 (N_20753,N_19490,N_19464);
and U20754 (N_20754,N_19553,N_19023);
or U20755 (N_20755,N_19881,N_19218);
and U20756 (N_20756,N_19355,N_19953);
nor U20757 (N_20757,N_19594,N_19939);
nand U20758 (N_20758,N_19638,N_19294);
nand U20759 (N_20759,N_19889,N_19239);
nand U20760 (N_20760,N_19909,N_19561);
nand U20761 (N_20761,N_19620,N_19836);
nand U20762 (N_20762,N_19962,N_19983);
nand U20763 (N_20763,N_19644,N_19080);
xor U20764 (N_20764,N_19655,N_19683);
or U20765 (N_20765,N_19789,N_19332);
xnor U20766 (N_20766,N_19216,N_19428);
nand U20767 (N_20767,N_19431,N_19196);
xor U20768 (N_20768,N_19450,N_19997);
xor U20769 (N_20769,N_19072,N_19186);
or U20770 (N_20770,N_19297,N_19888);
or U20771 (N_20771,N_19209,N_19744);
and U20772 (N_20772,N_19738,N_19264);
or U20773 (N_20773,N_19898,N_19212);
or U20774 (N_20774,N_19076,N_19690);
nand U20775 (N_20775,N_19874,N_19170);
nand U20776 (N_20776,N_19081,N_19935);
or U20777 (N_20777,N_19297,N_19452);
nor U20778 (N_20778,N_19642,N_19960);
and U20779 (N_20779,N_19810,N_19190);
or U20780 (N_20780,N_19271,N_19453);
nor U20781 (N_20781,N_19012,N_19111);
nor U20782 (N_20782,N_19543,N_19882);
and U20783 (N_20783,N_19831,N_19772);
nor U20784 (N_20784,N_19668,N_19237);
or U20785 (N_20785,N_19099,N_19744);
nand U20786 (N_20786,N_19633,N_19444);
and U20787 (N_20787,N_19350,N_19269);
nand U20788 (N_20788,N_19607,N_19928);
xor U20789 (N_20789,N_19597,N_19171);
and U20790 (N_20790,N_19970,N_19097);
nand U20791 (N_20791,N_19453,N_19320);
nor U20792 (N_20792,N_19881,N_19317);
xnor U20793 (N_20793,N_19604,N_19310);
and U20794 (N_20794,N_19233,N_19245);
nor U20795 (N_20795,N_19134,N_19262);
xor U20796 (N_20796,N_19597,N_19206);
nand U20797 (N_20797,N_19358,N_19694);
and U20798 (N_20798,N_19840,N_19142);
or U20799 (N_20799,N_19475,N_19110);
nor U20800 (N_20800,N_19555,N_19314);
or U20801 (N_20801,N_19504,N_19399);
or U20802 (N_20802,N_19073,N_19035);
nor U20803 (N_20803,N_19095,N_19127);
nand U20804 (N_20804,N_19386,N_19957);
and U20805 (N_20805,N_19432,N_19425);
nand U20806 (N_20806,N_19002,N_19499);
nand U20807 (N_20807,N_19095,N_19664);
and U20808 (N_20808,N_19242,N_19836);
and U20809 (N_20809,N_19239,N_19836);
and U20810 (N_20810,N_19315,N_19575);
nor U20811 (N_20811,N_19544,N_19628);
nor U20812 (N_20812,N_19997,N_19057);
nand U20813 (N_20813,N_19132,N_19158);
or U20814 (N_20814,N_19848,N_19473);
nor U20815 (N_20815,N_19228,N_19209);
xor U20816 (N_20816,N_19710,N_19461);
xor U20817 (N_20817,N_19111,N_19643);
xnor U20818 (N_20818,N_19991,N_19507);
nand U20819 (N_20819,N_19982,N_19754);
or U20820 (N_20820,N_19610,N_19449);
or U20821 (N_20821,N_19097,N_19250);
or U20822 (N_20822,N_19143,N_19062);
nor U20823 (N_20823,N_19865,N_19329);
nand U20824 (N_20824,N_19639,N_19020);
nand U20825 (N_20825,N_19844,N_19714);
nand U20826 (N_20826,N_19620,N_19925);
nor U20827 (N_20827,N_19288,N_19002);
or U20828 (N_20828,N_19190,N_19189);
xor U20829 (N_20829,N_19494,N_19170);
nand U20830 (N_20830,N_19128,N_19331);
or U20831 (N_20831,N_19080,N_19545);
nor U20832 (N_20832,N_19571,N_19788);
nand U20833 (N_20833,N_19249,N_19085);
nand U20834 (N_20834,N_19903,N_19027);
nor U20835 (N_20835,N_19523,N_19728);
nor U20836 (N_20836,N_19928,N_19025);
nor U20837 (N_20837,N_19232,N_19219);
nand U20838 (N_20838,N_19232,N_19064);
nor U20839 (N_20839,N_19511,N_19558);
nor U20840 (N_20840,N_19210,N_19243);
nand U20841 (N_20841,N_19619,N_19064);
nand U20842 (N_20842,N_19769,N_19628);
or U20843 (N_20843,N_19228,N_19400);
or U20844 (N_20844,N_19654,N_19073);
or U20845 (N_20845,N_19840,N_19740);
or U20846 (N_20846,N_19339,N_19441);
xor U20847 (N_20847,N_19241,N_19158);
xor U20848 (N_20848,N_19378,N_19989);
and U20849 (N_20849,N_19641,N_19252);
nor U20850 (N_20850,N_19858,N_19883);
or U20851 (N_20851,N_19867,N_19151);
or U20852 (N_20852,N_19888,N_19069);
or U20853 (N_20853,N_19715,N_19759);
or U20854 (N_20854,N_19121,N_19214);
nand U20855 (N_20855,N_19396,N_19339);
nand U20856 (N_20856,N_19743,N_19848);
or U20857 (N_20857,N_19550,N_19060);
xor U20858 (N_20858,N_19719,N_19589);
xnor U20859 (N_20859,N_19914,N_19974);
nand U20860 (N_20860,N_19695,N_19546);
and U20861 (N_20861,N_19721,N_19269);
or U20862 (N_20862,N_19270,N_19412);
or U20863 (N_20863,N_19071,N_19477);
and U20864 (N_20864,N_19040,N_19070);
xor U20865 (N_20865,N_19383,N_19575);
nor U20866 (N_20866,N_19548,N_19054);
nand U20867 (N_20867,N_19603,N_19428);
or U20868 (N_20868,N_19168,N_19665);
and U20869 (N_20869,N_19858,N_19238);
xnor U20870 (N_20870,N_19863,N_19406);
nand U20871 (N_20871,N_19705,N_19398);
xor U20872 (N_20872,N_19967,N_19423);
nor U20873 (N_20873,N_19500,N_19451);
nor U20874 (N_20874,N_19484,N_19954);
xnor U20875 (N_20875,N_19098,N_19466);
nor U20876 (N_20876,N_19714,N_19337);
xor U20877 (N_20877,N_19032,N_19670);
nor U20878 (N_20878,N_19095,N_19909);
nand U20879 (N_20879,N_19154,N_19483);
or U20880 (N_20880,N_19435,N_19489);
nor U20881 (N_20881,N_19258,N_19417);
and U20882 (N_20882,N_19351,N_19832);
or U20883 (N_20883,N_19950,N_19961);
or U20884 (N_20884,N_19664,N_19086);
nand U20885 (N_20885,N_19138,N_19125);
nand U20886 (N_20886,N_19474,N_19426);
xor U20887 (N_20887,N_19528,N_19984);
nor U20888 (N_20888,N_19103,N_19669);
and U20889 (N_20889,N_19502,N_19933);
and U20890 (N_20890,N_19417,N_19289);
nand U20891 (N_20891,N_19507,N_19131);
nor U20892 (N_20892,N_19263,N_19100);
or U20893 (N_20893,N_19818,N_19458);
and U20894 (N_20894,N_19072,N_19938);
xnor U20895 (N_20895,N_19129,N_19888);
xnor U20896 (N_20896,N_19818,N_19624);
nor U20897 (N_20897,N_19490,N_19745);
or U20898 (N_20898,N_19555,N_19642);
and U20899 (N_20899,N_19197,N_19366);
and U20900 (N_20900,N_19938,N_19422);
xnor U20901 (N_20901,N_19284,N_19017);
or U20902 (N_20902,N_19126,N_19780);
nor U20903 (N_20903,N_19136,N_19496);
or U20904 (N_20904,N_19897,N_19787);
and U20905 (N_20905,N_19903,N_19773);
xnor U20906 (N_20906,N_19337,N_19246);
and U20907 (N_20907,N_19867,N_19782);
nor U20908 (N_20908,N_19570,N_19115);
or U20909 (N_20909,N_19557,N_19445);
nor U20910 (N_20910,N_19829,N_19775);
xor U20911 (N_20911,N_19298,N_19033);
or U20912 (N_20912,N_19652,N_19636);
or U20913 (N_20913,N_19468,N_19278);
nand U20914 (N_20914,N_19975,N_19191);
or U20915 (N_20915,N_19575,N_19418);
xnor U20916 (N_20916,N_19859,N_19210);
nor U20917 (N_20917,N_19340,N_19870);
or U20918 (N_20918,N_19218,N_19640);
nand U20919 (N_20919,N_19863,N_19349);
xor U20920 (N_20920,N_19963,N_19124);
nor U20921 (N_20921,N_19537,N_19744);
or U20922 (N_20922,N_19640,N_19050);
nand U20923 (N_20923,N_19643,N_19387);
and U20924 (N_20924,N_19734,N_19826);
xor U20925 (N_20925,N_19469,N_19768);
and U20926 (N_20926,N_19954,N_19724);
xnor U20927 (N_20927,N_19076,N_19060);
or U20928 (N_20928,N_19506,N_19296);
nand U20929 (N_20929,N_19413,N_19918);
xor U20930 (N_20930,N_19215,N_19470);
and U20931 (N_20931,N_19094,N_19385);
nor U20932 (N_20932,N_19248,N_19269);
nor U20933 (N_20933,N_19356,N_19899);
nor U20934 (N_20934,N_19111,N_19078);
or U20935 (N_20935,N_19910,N_19884);
and U20936 (N_20936,N_19809,N_19334);
or U20937 (N_20937,N_19978,N_19399);
nand U20938 (N_20938,N_19410,N_19621);
nand U20939 (N_20939,N_19261,N_19568);
or U20940 (N_20940,N_19113,N_19040);
nor U20941 (N_20941,N_19959,N_19030);
xor U20942 (N_20942,N_19211,N_19040);
nand U20943 (N_20943,N_19237,N_19448);
nand U20944 (N_20944,N_19387,N_19150);
or U20945 (N_20945,N_19296,N_19987);
and U20946 (N_20946,N_19195,N_19219);
nor U20947 (N_20947,N_19601,N_19149);
xor U20948 (N_20948,N_19858,N_19904);
and U20949 (N_20949,N_19742,N_19449);
nand U20950 (N_20950,N_19665,N_19939);
nor U20951 (N_20951,N_19099,N_19628);
and U20952 (N_20952,N_19097,N_19734);
or U20953 (N_20953,N_19551,N_19845);
and U20954 (N_20954,N_19205,N_19757);
nand U20955 (N_20955,N_19557,N_19079);
nor U20956 (N_20956,N_19927,N_19464);
or U20957 (N_20957,N_19128,N_19559);
nor U20958 (N_20958,N_19910,N_19236);
and U20959 (N_20959,N_19499,N_19227);
nand U20960 (N_20960,N_19506,N_19099);
xnor U20961 (N_20961,N_19407,N_19789);
xor U20962 (N_20962,N_19690,N_19994);
nor U20963 (N_20963,N_19362,N_19028);
xnor U20964 (N_20964,N_19303,N_19116);
and U20965 (N_20965,N_19934,N_19669);
nor U20966 (N_20966,N_19344,N_19895);
and U20967 (N_20967,N_19830,N_19406);
nand U20968 (N_20968,N_19147,N_19669);
xor U20969 (N_20969,N_19340,N_19826);
xor U20970 (N_20970,N_19220,N_19520);
nand U20971 (N_20971,N_19927,N_19888);
or U20972 (N_20972,N_19344,N_19056);
and U20973 (N_20973,N_19913,N_19530);
or U20974 (N_20974,N_19520,N_19576);
nor U20975 (N_20975,N_19172,N_19930);
nor U20976 (N_20976,N_19242,N_19104);
and U20977 (N_20977,N_19822,N_19608);
nand U20978 (N_20978,N_19140,N_19461);
and U20979 (N_20979,N_19714,N_19763);
xor U20980 (N_20980,N_19449,N_19365);
nand U20981 (N_20981,N_19387,N_19938);
or U20982 (N_20982,N_19540,N_19246);
nand U20983 (N_20983,N_19139,N_19860);
and U20984 (N_20984,N_19140,N_19426);
nor U20985 (N_20985,N_19505,N_19223);
xor U20986 (N_20986,N_19709,N_19425);
and U20987 (N_20987,N_19817,N_19940);
or U20988 (N_20988,N_19610,N_19568);
or U20989 (N_20989,N_19868,N_19395);
nand U20990 (N_20990,N_19057,N_19483);
and U20991 (N_20991,N_19371,N_19373);
nor U20992 (N_20992,N_19124,N_19769);
and U20993 (N_20993,N_19918,N_19743);
nand U20994 (N_20994,N_19920,N_19510);
nand U20995 (N_20995,N_19529,N_19488);
xnor U20996 (N_20996,N_19584,N_19871);
or U20997 (N_20997,N_19624,N_19929);
and U20998 (N_20998,N_19804,N_19217);
xnor U20999 (N_20999,N_19880,N_19993);
nand U21000 (N_21000,N_20143,N_20305);
and U21001 (N_21001,N_20453,N_20053);
nand U21002 (N_21002,N_20370,N_20971);
nor U21003 (N_21003,N_20366,N_20713);
nor U21004 (N_21004,N_20936,N_20446);
nor U21005 (N_21005,N_20645,N_20479);
nand U21006 (N_21006,N_20439,N_20976);
and U21007 (N_21007,N_20888,N_20272);
or U21008 (N_21008,N_20759,N_20559);
and U21009 (N_21009,N_20984,N_20230);
nor U21010 (N_21010,N_20973,N_20749);
and U21011 (N_21011,N_20378,N_20607);
xor U21012 (N_21012,N_20225,N_20140);
or U21013 (N_21013,N_20592,N_20986);
or U21014 (N_21014,N_20867,N_20740);
or U21015 (N_21015,N_20982,N_20322);
nor U21016 (N_21016,N_20285,N_20425);
xnor U21017 (N_21017,N_20518,N_20808);
xor U21018 (N_21018,N_20448,N_20154);
nor U21019 (N_21019,N_20616,N_20841);
nand U21020 (N_21020,N_20754,N_20854);
xnor U21021 (N_21021,N_20006,N_20196);
nand U21022 (N_21022,N_20227,N_20901);
nand U21023 (N_21023,N_20168,N_20344);
xnor U21024 (N_21024,N_20447,N_20144);
or U21025 (N_21025,N_20325,N_20917);
nand U21026 (N_21026,N_20738,N_20727);
and U21027 (N_21027,N_20802,N_20609);
nor U21028 (N_21028,N_20768,N_20711);
or U21029 (N_21029,N_20408,N_20852);
xor U21030 (N_21030,N_20188,N_20342);
nor U21031 (N_21031,N_20517,N_20508);
nand U21032 (N_21032,N_20398,N_20849);
nand U21033 (N_21033,N_20864,N_20847);
xor U21034 (N_21034,N_20523,N_20496);
and U21035 (N_21035,N_20783,N_20379);
xnor U21036 (N_21036,N_20174,N_20644);
nor U21037 (N_21037,N_20511,N_20646);
nor U21038 (N_21038,N_20804,N_20903);
xor U21039 (N_21039,N_20894,N_20811);
xnor U21040 (N_21040,N_20666,N_20674);
nor U21041 (N_21041,N_20928,N_20625);
and U21042 (N_21042,N_20555,N_20362);
nand U21043 (N_21043,N_20582,N_20494);
and U21044 (N_21044,N_20078,N_20293);
xnor U21045 (N_21045,N_20597,N_20529);
or U21046 (N_21046,N_20039,N_20614);
and U21047 (N_21047,N_20076,N_20489);
or U21048 (N_21048,N_20203,N_20070);
or U21049 (N_21049,N_20764,N_20584);
xor U21050 (N_21050,N_20638,N_20710);
nor U21051 (N_21051,N_20530,N_20151);
nor U21052 (N_21052,N_20049,N_20690);
xor U21053 (N_21053,N_20891,N_20139);
nand U21054 (N_21054,N_20406,N_20234);
nand U21055 (N_21055,N_20777,N_20780);
nor U21056 (N_21056,N_20873,N_20624);
nand U21057 (N_21057,N_20637,N_20578);
xor U21058 (N_21058,N_20929,N_20796);
nand U21059 (N_21059,N_20985,N_20748);
nor U21060 (N_21060,N_20267,N_20474);
xnor U21061 (N_21061,N_20488,N_20136);
or U21062 (N_21062,N_20440,N_20159);
and U21063 (N_21063,N_20755,N_20449);
nor U21064 (N_21064,N_20250,N_20031);
nand U21065 (N_21065,N_20392,N_20634);
and U21066 (N_21066,N_20442,N_20138);
or U21067 (N_21067,N_20550,N_20732);
and U21068 (N_21068,N_20246,N_20429);
xor U21069 (N_21069,N_20916,N_20941);
and U21070 (N_21070,N_20712,N_20859);
nand U21071 (N_21071,N_20613,N_20826);
and U21072 (N_21072,N_20918,N_20622);
nor U21073 (N_21073,N_20452,N_20953);
nand U21074 (N_21074,N_20747,N_20235);
nor U21075 (N_21075,N_20153,N_20199);
xor U21076 (N_21076,N_20626,N_20217);
xor U21077 (N_21077,N_20498,N_20456);
nand U21078 (N_21078,N_20851,N_20321);
and U21079 (N_21079,N_20054,N_20506);
or U21080 (N_21080,N_20945,N_20333);
nor U21081 (N_21081,N_20468,N_20532);
nor U21082 (N_21082,N_20141,N_20301);
and U21083 (N_21083,N_20914,N_20944);
and U21084 (N_21084,N_20413,N_20337);
nor U21085 (N_21085,N_20902,N_20156);
nor U21086 (N_21086,N_20739,N_20018);
nand U21087 (N_21087,N_20348,N_20831);
or U21088 (N_21088,N_20603,N_20633);
nor U21089 (N_21089,N_20206,N_20545);
nand U21090 (N_21090,N_20436,N_20784);
or U21091 (N_21091,N_20512,N_20050);
nand U21092 (N_21092,N_20686,N_20654);
nor U21093 (N_21093,N_20191,N_20390);
nor U21094 (N_21094,N_20505,N_20067);
nor U21095 (N_21095,N_20059,N_20270);
and U21096 (N_21096,N_20715,N_20431);
or U21097 (N_21097,N_20595,N_20280);
nor U21098 (N_21098,N_20264,N_20961);
or U21099 (N_21099,N_20781,N_20298);
nand U21100 (N_21100,N_20731,N_20012);
or U21101 (N_21101,N_20495,N_20304);
or U21102 (N_21102,N_20951,N_20040);
nor U21103 (N_21103,N_20351,N_20694);
nor U21104 (N_21104,N_20157,N_20651);
and U21105 (N_21105,N_20382,N_20327);
nand U21106 (N_21106,N_20368,N_20691);
xor U21107 (N_21107,N_20357,N_20315);
and U21108 (N_21108,N_20347,N_20005);
or U21109 (N_21109,N_20499,N_20052);
and U21110 (N_21110,N_20998,N_20687);
nor U21111 (N_21111,N_20164,N_20172);
nand U21112 (N_21112,N_20492,N_20883);
and U21113 (N_21113,N_20701,N_20656);
and U21114 (N_21114,N_20210,N_20407);
xnor U21115 (N_21115,N_20969,N_20311);
nor U21116 (N_21116,N_20466,N_20521);
nor U21117 (N_21117,N_20335,N_20435);
nand U21118 (N_21118,N_20363,N_20332);
or U21119 (N_21119,N_20441,N_20878);
or U21120 (N_21120,N_20548,N_20403);
xor U21121 (N_21121,N_20538,N_20420);
and U21122 (N_21122,N_20433,N_20979);
and U21123 (N_21123,N_20244,N_20612);
nor U21124 (N_21124,N_20471,N_20387);
nand U21125 (N_21125,N_20035,N_20048);
or U21126 (N_21126,N_20991,N_20434);
and U21127 (N_21127,N_20127,N_20528);
nand U21128 (N_21128,N_20079,N_20109);
nor U21129 (N_21129,N_20911,N_20346);
and U21130 (N_21130,N_20650,N_20195);
nand U21131 (N_21131,N_20824,N_20730);
xor U21132 (N_21132,N_20469,N_20047);
nand U21133 (N_21133,N_20800,N_20265);
nand U21134 (N_21134,N_20213,N_20660);
nand U21135 (N_21135,N_20533,N_20340);
nand U21136 (N_21136,N_20177,N_20785);
nand U21137 (N_21137,N_20576,N_20621);
nor U21138 (N_21138,N_20450,N_20775);
nor U21139 (N_21139,N_20323,N_20173);
xor U21140 (N_21140,N_20835,N_20898);
and U21141 (N_21141,N_20557,N_20890);
and U21142 (N_21142,N_20410,N_20519);
nand U21143 (N_21143,N_20776,N_20829);
or U21144 (N_21144,N_20884,N_20258);
nor U21145 (N_21145,N_20721,N_20074);
xor U21146 (N_21146,N_20055,N_20818);
and U21147 (N_21147,N_20013,N_20610);
nor U21148 (N_21148,N_20123,N_20930);
or U21149 (N_21149,N_20572,N_20393);
nand U21150 (N_21150,N_20685,N_20359);
and U21151 (N_21151,N_20683,N_20451);
nor U21152 (N_21152,N_20478,N_20090);
xnor U21153 (N_21153,N_20668,N_20937);
and U21154 (N_21154,N_20960,N_20741);
nor U21155 (N_21155,N_20564,N_20167);
or U21156 (N_21156,N_20030,N_20094);
nand U21157 (N_21157,N_20825,N_20131);
nor U21158 (N_21158,N_20972,N_20038);
or U21159 (N_21159,N_20171,N_20146);
or U21160 (N_21160,N_20099,N_20635);
and U21161 (N_21161,N_20788,N_20628);
or U21162 (N_21162,N_20396,N_20790);
nor U21163 (N_21163,N_20709,N_20120);
nand U21164 (N_21164,N_20667,N_20580);
nor U21165 (N_21165,N_20194,N_20476);
nor U21166 (N_21166,N_20797,N_20111);
xnor U21167 (N_21167,N_20702,N_20827);
xor U21168 (N_21168,N_20515,N_20430);
and U21169 (N_21169,N_20068,N_20661);
nand U21170 (N_21170,N_20920,N_20027);
and U21171 (N_21171,N_20108,N_20490);
nor U21172 (N_21172,N_20836,N_20832);
and U21173 (N_21173,N_20166,N_20229);
or U21174 (N_21174,N_20073,N_20642);
xnor U21175 (N_21175,N_20733,N_20069);
or U21176 (N_21176,N_20716,N_20350);
xor U21177 (N_21177,N_20975,N_20017);
xor U21178 (N_21178,N_20718,N_20641);
nor U21179 (N_21179,N_20988,N_20077);
and U21180 (N_21180,N_20839,N_20266);
nor U21181 (N_21181,N_20724,N_20302);
nor U21182 (N_21182,N_20198,N_20560);
or U21183 (N_21183,N_20245,N_20300);
nand U21184 (N_21184,N_20487,N_20014);
xor U21185 (N_21185,N_20228,N_20662);
and U21186 (N_21186,N_20409,N_20537);
xor U21187 (N_21187,N_20485,N_20980);
nor U21188 (N_21188,N_20653,N_20830);
xnor U21189 (N_21189,N_20799,N_20256);
nand U21190 (N_21190,N_20688,N_20544);
nand U21191 (N_21191,N_20291,N_20855);
nor U21192 (N_21192,N_20161,N_20850);
and U21193 (N_21193,N_20046,N_20795);
or U21194 (N_21194,N_20118,N_20274);
nand U21195 (N_21195,N_20954,N_20218);
and U21196 (N_21196,N_20587,N_20672);
nand U21197 (N_21197,N_20107,N_20925);
nor U21198 (N_21198,N_20947,N_20689);
xnor U21199 (N_21199,N_20414,N_20725);
xnor U21200 (N_21200,N_20756,N_20561);
nand U21201 (N_21201,N_20678,N_20760);
xor U21202 (N_21202,N_20879,N_20583);
nor U21203 (N_21203,N_20990,N_20761);
or U21204 (N_21204,N_20722,N_20513);
nand U21205 (N_21205,N_20170,N_20726);
or U21206 (N_21206,N_20303,N_20290);
xnor U21207 (N_21207,N_20306,N_20381);
nand U21208 (N_21208,N_20862,N_20137);
nor U21209 (N_21209,N_20871,N_20288);
nand U21210 (N_21210,N_20707,N_20509);
nor U21211 (N_21211,N_20966,N_20243);
or U21212 (N_21212,N_20394,N_20126);
and U21213 (N_21213,N_20695,N_20751);
nor U21214 (N_21214,N_20869,N_20639);
or U21215 (N_21215,N_20385,N_20994);
nand U21216 (N_21216,N_20581,N_20135);
and U21217 (N_21217,N_20465,N_20803);
nand U21218 (N_21218,N_20853,N_20910);
nand U21219 (N_21219,N_20921,N_20698);
nand U21220 (N_21220,N_20913,N_20568);
nor U21221 (N_21221,N_20377,N_20556);
xor U21222 (N_21222,N_20791,N_20504);
or U21223 (N_21223,N_20081,N_20673);
xnor U21224 (N_21224,N_20843,N_20432);
or U21225 (N_21225,N_20813,N_20402);
nor U21226 (N_21226,N_20259,N_20062);
nor U21227 (N_21227,N_20838,N_20640);
nand U21228 (N_21228,N_20957,N_20604);
or U21229 (N_21229,N_20185,N_20809);
or U21230 (N_21230,N_20482,N_20636);
nor U21231 (N_21231,N_20949,N_20268);
nand U21232 (N_21232,N_20692,N_20263);
nor U21233 (N_21233,N_20602,N_20223);
nand U21234 (N_21234,N_20993,N_20464);
nand U21235 (N_21235,N_20814,N_20536);
or U21236 (N_21236,N_20475,N_20457);
xor U21237 (N_21237,N_20356,N_20214);
nand U21238 (N_21238,N_20798,N_20992);
and U21239 (N_21239,N_20939,N_20455);
nand U21240 (N_21240,N_20473,N_20297);
xor U21241 (N_21241,N_20887,N_20872);
nor U21242 (N_21242,N_20428,N_20593);
nor U21243 (N_21243,N_20320,N_20282);
nand U21244 (N_21244,N_20423,N_20365);
and U21245 (N_21245,N_20334,N_20591);
xnor U21246 (N_21246,N_20658,N_20411);
nand U21247 (N_21247,N_20178,N_20573);
or U21248 (N_21248,N_20150,N_20345);
xor U21249 (N_21249,N_20906,N_20026);
xnor U21250 (N_21250,N_20620,N_20995);
xnor U21251 (N_21251,N_20208,N_20534);
nand U21252 (N_21252,N_20395,N_20514);
nor U21253 (N_21253,N_20743,N_20909);
nor U21254 (N_21254,N_20096,N_20611);
or U21255 (N_21255,N_20720,N_20866);
or U21256 (N_21256,N_20106,N_20255);
or U21257 (N_21257,N_20946,N_20856);
and U21258 (N_21258,N_20353,N_20343);
or U21259 (N_21259,N_20373,N_20372);
nor U21260 (N_21260,N_20098,N_20480);
xnor U21261 (N_21261,N_20241,N_20585);
and U21262 (N_21262,N_20531,N_20599);
and U21263 (N_21263,N_20842,N_20786);
nor U21264 (N_21264,N_20286,N_20770);
nor U21265 (N_21265,N_20084,N_20287);
nand U21266 (N_21266,N_20367,N_20412);
nand U21267 (N_21267,N_20655,N_20086);
nor U21268 (N_21268,N_20577,N_20181);
xor U21269 (N_21269,N_20184,N_20276);
nand U21270 (N_21270,N_20249,N_20943);
and U21271 (N_21271,N_20773,N_20959);
nor U21272 (N_21272,N_20549,N_20503);
nand U21273 (N_21273,N_20080,N_20215);
or U21274 (N_21274,N_20060,N_20391);
xnor U21275 (N_21275,N_20647,N_20767);
and U21276 (N_21276,N_20977,N_20907);
and U21277 (N_21277,N_20484,N_20175);
and U21278 (N_21278,N_20251,N_20422);
nor U21279 (N_21279,N_20101,N_20817);
and U21280 (N_21280,N_20360,N_20095);
and U21281 (N_21281,N_20438,N_20400);
or U21282 (N_21282,N_20192,N_20664);
or U21283 (N_21283,N_20539,N_20426);
nand U21284 (N_21284,N_20665,N_20324);
or U21285 (N_21285,N_20762,N_20868);
nor U21286 (N_21286,N_20187,N_20397);
nor U21287 (N_21287,N_20216,N_20269);
xor U21288 (N_21288,N_20676,N_20483);
nand U21289 (N_21289,N_20404,N_20844);
nand U21290 (N_21290,N_20331,N_20806);
nand U21291 (N_21291,N_20358,N_20923);
or U21292 (N_21292,N_20354,N_20364);
nand U21293 (N_21293,N_20543,N_20956);
xnor U21294 (N_21294,N_20034,N_20071);
xnor U21295 (N_21295,N_20766,N_20805);
nand U21296 (N_21296,N_20932,N_20222);
nor U21297 (N_21297,N_20043,N_20072);
nor U21298 (N_21298,N_20061,N_20459);
xor U21299 (N_21299,N_20454,N_20097);
nand U21300 (N_21300,N_20815,N_20875);
and U21301 (N_21301,N_20963,N_20083);
nor U21302 (N_21302,N_20242,N_20962);
nor U21303 (N_21303,N_20938,N_20510);
xnor U21304 (N_21304,N_20905,N_20541);
nand U21305 (N_21305,N_20605,N_20057);
or U21306 (N_21306,N_20600,N_20386);
and U21307 (N_21307,N_20794,N_20663);
nor U21308 (N_21308,N_20369,N_20317);
and U21309 (N_21309,N_20204,N_20165);
nor U21310 (N_21310,N_20032,N_20000);
nand U21311 (N_21311,N_20114,N_20970);
and U21312 (N_21312,N_20091,N_20669);
or U21313 (N_21313,N_20629,N_20117);
xnor U21314 (N_21314,N_20190,N_20128);
nand U21315 (N_21315,N_20734,N_20729);
or U21316 (N_21316,N_20024,N_20458);
and U21317 (N_21317,N_20877,N_20893);
nand U21318 (N_21318,N_20289,N_20124);
nand U21319 (N_21319,N_20355,N_20940);
or U21320 (N_21320,N_20586,N_20863);
xnor U21321 (N_21321,N_20374,N_20085);
and U21322 (N_21322,N_20237,N_20226);
nand U21323 (N_21323,N_20328,N_20819);
or U21324 (N_21324,N_20516,N_20443);
and U21325 (N_21325,N_20737,N_20999);
nor U21326 (N_21326,N_20679,N_20326);
nand U21327 (N_21327,N_20179,N_20418);
and U21328 (N_21328,N_20745,N_20082);
or U21329 (N_21329,N_20384,N_20997);
or U21330 (N_21330,N_20981,N_20574);
nand U21331 (N_21331,N_20460,N_20112);
xnor U21332 (N_21332,N_20240,N_20497);
nor U21333 (N_21333,N_20983,N_20820);
nand U21334 (N_21334,N_20763,N_20525);
nor U21335 (N_21335,N_20093,N_20933);
and U21336 (N_21336,N_20389,N_20491);
nor U21337 (N_21337,N_20769,N_20589);
and U21338 (N_21338,N_20472,N_20833);
or U21339 (N_21339,N_20569,N_20105);
nand U21340 (N_21340,N_20704,N_20522);
xnor U21341 (N_21341,N_20121,N_20792);
and U21342 (N_21342,N_20033,N_20912);
or U21343 (N_21343,N_20419,N_20252);
xor U21344 (N_21344,N_20421,N_20044);
nand U21345 (N_21345,N_20020,N_20787);
and U21346 (N_21346,N_20219,N_20857);
nor U21347 (N_21347,N_20296,N_20182);
nor U21348 (N_21348,N_20500,N_20132);
nor U21349 (N_21349,N_20996,N_20899);
or U21350 (N_21350,N_20765,N_20437);
and U21351 (N_21351,N_20160,N_20371);
nand U21352 (N_21352,N_20104,N_20837);
nand U21353 (N_21353,N_20461,N_20526);
and U21354 (N_21354,N_20922,N_20927);
nand U21355 (N_21355,N_20840,N_20858);
nand U21356 (N_21356,N_20313,N_20680);
xnor U21357 (N_21357,N_20757,N_20834);
or U21358 (N_21358,N_20812,N_20520);
nor U21359 (N_21359,N_20008,N_20703);
and U21360 (N_21360,N_20007,N_20036);
or U21361 (N_21361,N_20880,N_20816);
and U21362 (N_21362,N_20260,N_20885);
xnor U21363 (N_21363,N_20895,N_20897);
nor U21364 (N_21364,N_20870,N_20231);
xor U21365 (N_21365,N_20417,N_20349);
nand U21366 (N_21366,N_20952,N_20312);
nand U21367 (N_21367,N_20041,N_20598);
nand U21368 (N_21368,N_20924,N_20562);
or U21369 (N_21369,N_20502,N_20719);
nor U21370 (N_21370,N_20158,N_20958);
xnor U21371 (N_21371,N_20376,N_20019);
xor U21372 (N_21372,N_20279,N_20176);
nor U21373 (N_21373,N_20551,N_20744);
xor U21374 (N_21374,N_20169,N_20009);
xor U21375 (N_21375,N_20205,N_20470);
or U21376 (N_21376,N_20401,N_20643);
nand U21377 (N_21377,N_20463,N_20606);
xnor U21378 (N_21378,N_20115,N_20281);
nand U21379 (N_21379,N_20310,N_20361);
or U21380 (N_21380,N_20671,N_20295);
and U21381 (N_21381,N_20696,N_20129);
nor U21382 (N_21382,N_20527,N_20978);
and U21383 (N_21383,N_20200,N_20066);
and U21384 (N_21384,N_20016,N_20631);
or U21385 (N_21385,N_20771,N_20163);
and U21386 (N_21386,N_20257,N_20180);
or U21387 (N_21387,N_20283,N_20915);
and U21388 (N_21388,N_20388,N_20209);
or U21389 (N_21389,N_20003,N_20728);
xor U21390 (N_21390,N_20567,N_20058);
nand U21391 (N_21391,N_20125,N_20065);
and U21392 (N_21392,N_20779,N_20801);
and U21393 (N_21393,N_20380,N_20247);
nor U21394 (N_21394,N_20197,N_20821);
and U21395 (N_21395,N_20900,N_20162);
nor U21396 (N_21396,N_20659,N_20481);
xnor U21397 (N_21397,N_20271,N_20758);
xnor U21398 (N_21398,N_20789,N_20424);
or U21399 (N_21399,N_20462,N_20233);
nor U21400 (N_21400,N_20029,N_20964);
xnor U21401 (N_21401,N_20028,N_20845);
xor U21402 (N_21402,N_20861,N_20236);
xor U21403 (N_21403,N_20684,N_20699);
nand U21404 (N_21404,N_20700,N_20261);
nor U21405 (N_21405,N_20588,N_20735);
xor U21406 (N_21406,N_20697,N_20056);
and U21407 (N_21407,N_20113,N_20089);
nor U21408 (N_21408,N_20717,N_20427);
nor U21409 (N_21409,N_20254,N_20753);
xnor U21410 (N_21410,N_20063,N_20299);
or U21411 (N_21411,N_20778,N_20565);
nor U21412 (N_21412,N_20087,N_20212);
xnor U21413 (N_21413,N_20336,N_20193);
xor U21414 (N_21414,N_20535,N_20022);
nor U21415 (N_21415,N_20860,N_20186);
nand U21416 (N_21416,N_20823,N_20262);
and U21417 (N_21417,N_20563,N_20399);
nor U21418 (N_21418,N_20445,N_20493);
and U21419 (N_21419,N_20968,N_20284);
xnor U21420 (N_21420,N_20736,N_20554);
xor U21421 (N_21421,N_20706,N_20675);
nor U21422 (N_21422,N_20375,N_20708);
and U21423 (N_21423,N_20571,N_20810);
nor U21424 (N_21424,N_20618,N_20277);
xor U21425 (N_21425,N_20596,N_20075);
and U21426 (N_21426,N_20546,N_20248);
or U21427 (N_21427,N_20989,N_20133);
nand U21428 (N_21428,N_20318,N_20896);
xor U21429 (N_21429,N_20705,N_20103);
and U21430 (N_21430,N_20221,N_20207);
nand U21431 (N_21431,N_20025,N_20822);
or U21432 (N_21432,N_20148,N_20339);
or U21433 (N_21433,N_20967,N_20122);
and U21434 (N_21434,N_20881,N_20308);
and U21435 (N_21435,N_20416,N_20552);
and U21436 (N_21436,N_20950,N_20590);
and U21437 (N_21437,N_20130,N_20627);
xnor U21438 (N_21438,N_20201,N_20100);
nor U21439 (N_21439,N_20874,N_20886);
nor U21440 (N_21440,N_20615,N_20682);
nor U21441 (N_21441,N_20149,N_20575);
nand U21442 (N_21442,N_20045,N_20278);
nand U21443 (N_21443,N_20330,N_20892);
and U21444 (N_21444,N_20579,N_20011);
and U21445 (N_21445,N_20558,N_20594);
nand U21446 (N_21446,N_20782,N_20623);
and U21447 (N_21447,N_20486,N_20352);
nand U21448 (N_21448,N_20329,N_20467);
and U21449 (N_21449,N_20919,N_20183);
or U21450 (N_21450,N_20142,N_20064);
nand U21451 (N_21451,N_20649,N_20772);
xor U21452 (N_21452,N_20232,N_20652);
or U21453 (N_21453,N_20846,N_20002);
and U21454 (N_21454,N_20010,N_20238);
nor U21455 (N_21455,N_20848,N_20542);
and U21456 (N_21456,N_20934,N_20092);
nand U21457 (N_21457,N_20601,N_20015);
xor U21458 (N_21458,N_20608,N_20714);
and U21459 (N_21459,N_20224,N_20974);
or U21460 (N_21460,N_20189,N_20220);
and U21461 (N_21461,N_20147,N_20774);
or U21462 (N_21462,N_20405,N_20630);
xnor U21463 (N_21463,N_20524,N_20904);
nor U21464 (N_21464,N_20501,N_20338);
and U21465 (N_21465,N_20617,N_20145);
and U21466 (N_21466,N_20273,N_20965);
nand U21467 (N_21467,N_20004,N_20648);
and U21468 (N_21468,N_20632,N_20987);
or U21469 (N_21469,N_20807,N_20001);
or U21470 (N_21470,N_20110,N_20152);
and U21471 (N_21471,N_20507,N_20926);
or U21472 (N_21472,N_20314,N_20307);
or U21473 (N_21473,N_20828,N_20211);
or U21474 (N_21474,N_20677,N_20116);
xor U21475 (N_21475,N_20746,N_20742);
xnor U21476 (N_21476,N_20253,N_20309);
nor U21477 (N_21477,N_20239,N_20444);
nand U21478 (N_21478,N_20134,N_20119);
nor U21479 (N_21479,N_20876,N_20292);
nor U21480 (N_21480,N_20570,N_20316);
nor U21481 (N_21481,N_20383,N_20882);
nor U21482 (N_21482,N_20553,N_20415);
or U21483 (N_21483,N_20657,N_20793);
xor U21484 (N_21484,N_20931,N_20202);
nand U21485 (N_21485,N_20681,N_20540);
and U21486 (N_21486,N_20723,N_20942);
or U21487 (N_21487,N_20319,N_20037);
or U21488 (N_21488,N_20935,N_20341);
nor U21489 (N_21489,N_20619,N_20566);
nor U21490 (N_21490,N_20088,N_20948);
xnor U21491 (N_21491,N_20750,N_20023);
or U21492 (N_21492,N_20865,N_20155);
and U21493 (N_21493,N_20294,N_20275);
nand U21494 (N_21494,N_20477,N_20889);
and U21495 (N_21495,N_20547,N_20752);
nor U21496 (N_21496,N_20051,N_20670);
or U21497 (N_21497,N_20693,N_20102);
xor U21498 (N_21498,N_20908,N_20042);
nor U21499 (N_21499,N_20955,N_20021);
nand U21500 (N_21500,N_20097,N_20989);
and U21501 (N_21501,N_20477,N_20468);
xor U21502 (N_21502,N_20092,N_20821);
nand U21503 (N_21503,N_20297,N_20081);
or U21504 (N_21504,N_20499,N_20890);
nor U21505 (N_21505,N_20940,N_20854);
nand U21506 (N_21506,N_20522,N_20762);
or U21507 (N_21507,N_20475,N_20538);
and U21508 (N_21508,N_20996,N_20184);
or U21509 (N_21509,N_20666,N_20137);
xnor U21510 (N_21510,N_20696,N_20783);
and U21511 (N_21511,N_20942,N_20568);
and U21512 (N_21512,N_20783,N_20012);
or U21513 (N_21513,N_20767,N_20886);
nor U21514 (N_21514,N_20628,N_20816);
nand U21515 (N_21515,N_20553,N_20348);
nand U21516 (N_21516,N_20414,N_20598);
and U21517 (N_21517,N_20693,N_20588);
nor U21518 (N_21518,N_20721,N_20583);
and U21519 (N_21519,N_20445,N_20574);
and U21520 (N_21520,N_20840,N_20259);
or U21521 (N_21521,N_20778,N_20701);
xnor U21522 (N_21522,N_20932,N_20542);
or U21523 (N_21523,N_20393,N_20364);
and U21524 (N_21524,N_20220,N_20393);
nor U21525 (N_21525,N_20975,N_20495);
nor U21526 (N_21526,N_20547,N_20263);
nor U21527 (N_21527,N_20342,N_20072);
or U21528 (N_21528,N_20929,N_20217);
xnor U21529 (N_21529,N_20081,N_20204);
and U21530 (N_21530,N_20728,N_20779);
and U21531 (N_21531,N_20622,N_20471);
and U21532 (N_21532,N_20456,N_20085);
or U21533 (N_21533,N_20988,N_20473);
nand U21534 (N_21534,N_20988,N_20846);
nand U21535 (N_21535,N_20390,N_20244);
nand U21536 (N_21536,N_20531,N_20613);
nand U21537 (N_21537,N_20839,N_20982);
and U21538 (N_21538,N_20604,N_20356);
and U21539 (N_21539,N_20296,N_20400);
or U21540 (N_21540,N_20333,N_20319);
xor U21541 (N_21541,N_20913,N_20215);
and U21542 (N_21542,N_20849,N_20333);
xor U21543 (N_21543,N_20799,N_20890);
or U21544 (N_21544,N_20892,N_20672);
and U21545 (N_21545,N_20687,N_20848);
nand U21546 (N_21546,N_20797,N_20529);
and U21547 (N_21547,N_20392,N_20941);
or U21548 (N_21548,N_20795,N_20115);
and U21549 (N_21549,N_20936,N_20310);
and U21550 (N_21550,N_20612,N_20621);
xor U21551 (N_21551,N_20363,N_20508);
nor U21552 (N_21552,N_20197,N_20486);
nand U21553 (N_21553,N_20310,N_20133);
or U21554 (N_21554,N_20567,N_20568);
nor U21555 (N_21555,N_20006,N_20756);
nor U21556 (N_21556,N_20992,N_20660);
or U21557 (N_21557,N_20772,N_20089);
nand U21558 (N_21558,N_20439,N_20023);
nand U21559 (N_21559,N_20191,N_20209);
nor U21560 (N_21560,N_20310,N_20450);
or U21561 (N_21561,N_20443,N_20271);
xnor U21562 (N_21562,N_20257,N_20813);
or U21563 (N_21563,N_20564,N_20957);
nor U21564 (N_21564,N_20623,N_20892);
nand U21565 (N_21565,N_20289,N_20971);
or U21566 (N_21566,N_20464,N_20188);
or U21567 (N_21567,N_20844,N_20992);
xnor U21568 (N_21568,N_20758,N_20335);
nand U21569 (N_21569,N_20017,N_20920);
xnor U21570 (N_21570,N_20314,N_20842);
and U21571 (N_21571,N_20419,N_20255);
or U21572 (N_21572,N_20634,N_20631);
or U21573 (N_21573,N_20856,N_20640);
nand U21574 (N_21574,N_20570,N_20129);
xor U21575 (N_21575,N_20995,N_20904);
and U21576 (N_21576,N_20144,N_20974);
xnor U21577 (N_21577,N_20985,N_20991);
nor U21578 (N_21578,N_20245,N_20790);
xnor U21579 (N_21579,N_20313,N_20489);
nand U21580 (N_21580,N_20705,N_20861);
and U21581 (N_21581,N_20637,N_20034);
nand U21582 (N_21582,N_20261,N_20668);
xnor U21583 (N_21583,N_20074,N_20126);
and U21584 (N_21584,N_20393,N_20489);
or U21585 (N_21585,N_20611,N_20805);
and U21586 (N_21586,N_20395,N_20680);
xnor U21587 (N_21587,N_20228,N_20726);
and U21588 (N_21588,N_20704,N_20854);
or U21589 (N_21589,N_20197,N_20156);
nor U21590 (N_21590,N_20271,N_20214);
or U21591 (N_21591,N_20945,N_20034);
and U21592 (N_21592,N_20156,N_20417);
xor U21593 (N_21593,N_20842,N_20977);
nor U21594 (N_21594,N_20035,N_20566);
nor U21595 (N_21595,N_20562,N_20887);
xor U21596 (N_21596,N_20211,N_20075);
and U21597 (N_21597,N_20006,N_20340);
and U21598 (N_21598,N_20162,N_20460);
nand U21599 (N_21599,N_20021,N_20202);
or U21600 (N_21600,N_20810,N_20683);
xnor U21601 (N_21601,N_20343,N_20495);
or U21602 (N_21602,N_20243,N_20457);
nor U21603 (N_21603,N_20524,N_20607);
nand U21604 (N_21604,N_20281,N_20807);
or U21605 (N_21605,N_20352,N_20328);
nor U21606 (N_21606,N_20572,N_20040);
nor U21607 (N_21607,N_20879,N_20435);
xnor U21608 (N_21608,N_20493,N_20031);
or U21609 (N_21609,N_20760,N_20894);
nor U21610 (N_21610,N_20655,N_20259);
xnor U21611 (N_21611,N_20963,N_20881);
nor U21612 (N_21612,N_20787,N_20103);
or U21613 (N_21613,N_20780,N_20466);
or U21614 (N_21614,N_20743,N_20346);
and U21615 (N_21615,N_20317,N_20150);
xnor U21616 (N_21616,N_20782,N_20592);
xnor U21617 (N_21617,N_20425,N_20815);
xnor U21618 (N_21618,N_20940,N_20199);
nor U21619 (N_21619,N_20303,N_20472);
nand U21620 (N_21620,N_20885,N_20962);
or U21621 (N_21621,N_20357,N_20820);
nand U21622 (N_21622,N_20005,N_20436);
nand U21623 (N_21623,N_20589,N_20634);
xnor U21624 (N_21624,N_20758,N_20464);
or U21625 (N_21625,N_20203,N_20330);
nor U21626 (N_21626,N_20917,N_20304);
nand U21627 (N_21627,N_20422,N_20303);
nand U21628 (N_21628,N_20126,N_20906);
and U21629 (N_21629,N_20000,N_20994);
or U21630 (N_21630,N_20868,N_20890);
xnor U21631 (N_21631,N_20447,N_20927);
or U21632 (N_21632,N_20944,N_20635);
or U21633 (N_21633,N_20671,N_20335);
nand U21634 (N_21634,N_20195,N_20133);
and U21635 (N_21635,N_20217,N_20407);
and U21636 (N_21636,N_20038,N_20886);
and U21637 (N_21637,N_20097,N_20581);
and U21638 (N_21638,N_20437,N_20033);
nand U21639 (N_21639,N_20202,N_20158);
xnor U21640 (N_21640,N_20667,N_20759);
nand U21641 (N_21641,N_20007,N_20487);
nor U21642 (N_21642,N_20139,N_20903);
nor U21643 (N_21643,N_20498,N_20003);
or U21644 (N_21644,N_20545,N_20761);
xor U21645 (N_21645,N_20440,N_20592);
and U21646 (N_21646,N_20502,N_20893);
xnor U21647 (N_21647,N_20746,N_20498);
and U21648 (N_21648,N_20366,N_20103);
nor U21649 (N_21649,N_20343,N_20554);
nor U21650 (N_21650,N_20304,N_20272);
nor U21651 (N_21651,N_20378,N_20079);
or U21652 (N_21652,N_20592,N_20690);
or U21653 (N_21653,N_20685,N_20204);
nand U21654 (N_21654,N_20597,N_20306);
nor U21655 (N_21655,N_20374,N_20494);
xnor U21656 (N_21656,N_20638,N_20946);
nand U21657 (N_21657,N_20081,N_20174);
xnor U21658 (N_21658,N_20880,N_20960);
nand U21659 (N_21659,N_20906,N_20394);
nand U21660 (N_21660,N_20123,N_20745);
and U21661 (N_21661,N_20629,N_20850);
nor U21662 (N_21662,N_20781,N_20665);
nor U21663 (N_21663,N_20345,N_20725);
nor U21664 (N_21664,N_20295,N_20519);
or U21665 (N_21665,N_20826,N_20898);
nor U21666 (N_21666,N_20685,N_20620);
nand U21667 (N_21667,N_20733,N_20008);
nand U21668 (N_21668,N_20449,N_20304);
and U21669 (N_21669,N_20612,N_20413);
xor U21670 (N_21670,N_20458,N_20422);
or U21671 (N_21671,N_20327,N_20793);
and U21672 (N_21672,N_20281,N_20931);
nand U21673 (N_21673,N_20328,N_20524);
or U21674 (N_21674,N_20928,N_20530);
nand U21675 (N_21675,N_20086,N_20576);
xor U21676 (N_21676,N_20867,N_20542);
or U21677 (N_21677,N_20902,N_20945);
or U21678 (N_21678,N_20834,N_20591);
or U21679 (N_21679,N_20967,N_20715);
nand U21680 (N_21680,N_20039,N_20564);
nand U21681 (N_21681,N_20750,N_20145);
nor U21682 (N_21682,N_20087,N_20717);
nor U21683 (N_21683,N_20866,N_20479);
and U21684 (N_21684,N_20576,N_20036);
nor U21685 (N_21685,N_20408,N_20659);
xnor U21686 (N_21686,N_20344,N_20235);
or U21687 (N_21687,N_20896,N_20953);
xor U21688 (N_21688,N_20534,N_20658);
nand U21689 (N_21689,N_20793,N_20557);
or U21690 (N_21690,N_20050,N_20668);
xnor U21691 (N_21691,N_20138,N_20811);
or U21692 (N_21692,N_20876,N_20114);
nor U21693 (N_21693,N_20815,N_20634);
nand U21694 (N_21694,N_20310,N_20806);
or U21695 (N_21695,N_20994,N_20584);
nor U21696 (N_21696,N_20487,N_20216);
nor U21697 (N_21697,N_20716,N_20170);
nor U21698 (N_21698,N_20882,N_20314);
or U21699 (N_21699,N_20773,N_20531);
nor U21700 (N_21700,N_20201,N_20192);
xnor U21701 (N_21701,N_20247,N_20653);
and U21702 (N_21702,N_20182,N_20523);
nor U21703 (N_21703,N_20507,N_20963);
and U21704 (N_21704,N_20084,N_20948);
or U21705 (N_21705,N_20968,N_20356);
and U21706 (N_21706,N_20093,N_20214);
nor U21707 (N_21707,N_20352,N_20565);
xnor U21708 (N_21708,N_20954,N_20729);
or U21709 (N_21709,N_20347,N_20244);
or U21710 (N_21710,N_20290,N_20167);
nor U21711 (N_21711,N_20285,N_20884);
nor U21712 (N_21712,N_20457,N_20014);
or U21713 (N_21713,N_20559,N_20062);
xor U21714 (N_21714,N_20357,N_20171);
nor U21715 (N_21715,N_20724,N_20896);
nand U21716 (N_21716,N_20280,N_20952);
nand U21717 (N_21717,N_20575,N_20897);
or U21718 (N_21718,N_20892,N_20298);
xor U21719 (N_21719,N_20285,N_20321);
or U21720 (N_21720,N_20654,N_20388);
and U21721 (N_21721,N_20081,N_20086);
and U21722 (N_21722,N_20034,N_20143);
xnor U21723 (N_21723,N_20309,N_20519);
and U21724 (N_21724,N_20400,N_20613);
nand U21725 (N_21725,N_20720,N_20242);
or U21726 (N_21726,N_20668,N_20648);
nor U21727 (N_21727,N_20668,N_20044);
or U21728 (N_21728,N_20585,N_20259);
or U21729 (N_21729,N_20886,N_20756);
xor U21730 (N_21730,N_20719,N_20826);
nand U21731 (N_21731,N_20618,N_20003);
nor U21732 (N_21732,N_20162,N_20596);
and U21733 (N_21733,N_20450,N_20839);
nand U21734 (N_21734,N_20178,N_20419);
or U21735 (N_21735,N_20187,N_20488);
nand U21736 (N_21736,N_20055,N_20073);
xnor U21737 (N_21737,N_20632,N_20921);
nor U21738 (N_21738,N_20062,N_20965);
and U21739 (N_21739,N_20543,N_20752);
and U21740 (N_21740,N_20874,N_20527);
and U21741 (N_21741,N_20712,N_20484);
and U21742 (N_21742,N_20017,N_20749);
or U21743 (N_21743,N_20973,N_20927);
and U21744 (N_21744,N_20782,N_20382);
xnor U21745 (N_21745,N_20067,N_20902);
and U21746 (N_21746,N_20623,N_20887);
nand U21747 (N_21747,N_20461,N_20131);
xnor U21748 (N_21748,N_20448,N_20043);
nand U21749 (N_21749,N_20317,N_20447);
and U21750 (N_21750,N_20920,N_20708);
or U21751 (N_21751,N_20991,N_20964);
nand U21752 (N_21752,N_20051,N_20896);
xnor U21753 (N_21753,N_20565,N_20732);
nor U21754 (N_21754,N_20519,N_20369);
nand U21755 (N_21755,N_20502,N_20096);
nor U21756 (N_21756,N_20836,N_20921);
xnor U21757 (N_21757,N_20611,N_20397);
xnor U21758 (N_21758,N_20269,N_20376);
and U21759 (N_21759,N_20063,N_20992);
xnor U21760 (N_21760,N_20451,N_20480);
or U21761 (N_21761,N_20684,N_20047);
nor U21762 (N_21762,N_20754,N_20936);
nor U21763 (N_21763,N_20587,N_20017);
and U21764 (N_21764,N_20513,N_20965);
or U21765 (N_21765,N_20289,N_20172);
or U21766 (N_21766,N_20372,N_20120);
or U21767 (N_21767,N_20460,N_20847);
xor U21768 (N_21768,N_20366,N_20083);
nor U21769 (N_21769,N_20451,N_20875);
xor U21770 (N_21770,N_20965,N_20073);
or U21771 (N_21771,N_20855,N_20936);
nor U21772 (N_21772,N_20207,N_20367);
or U21773 (N_21773,N_20945,N_20955);
or U21774 (N_21774,N_20552,N_20130);
nand U21775 (N_21775,N_20521,N_20535);
xor U21776 (N_21776,N_20867,N_20198);
and U21777 (N_21777,N_20877,N_20322);
nor U21778 (N_21778,N_20201,N_20723);
and U21779 (N_21779,N_20977,N_20994);
xnor U21780 (N_21780,N_20689,N_20057);
or U21781 (N_21781,N_20794,N_20023);
xnor U21782 (N_21782,N_20163,N_20445);
or U21783 (N_21783,N_20997,N_20425);
or U21784 (N_21784,N_20496,N_20055);
or U21785 (N_21785,N_20518,N_20363);
nor U21786 (N_21786,N_20433,N_20092);
nand U21787 (N_21787,N_20027,N_20522);
and U21788 (N_21788,N_20560,N_20262);
or U21789 (N_21789,N_20051,N_20305);
and U21790 (N_21790,N_20579,N_20739);
nor U21791 (N_21791,N_20802,N_20560);
or U21792 (N_21792,N_20917,N_20094);
or U21793 (N_21793,N_20054,N_20452);
or U21794 (N_21794,N_20482,N_20040);
or U21795 (N_21795,N_20601,N_20512);
and U21796 (N_21796,N_20736,N_20130);
nor U21797 (N_21797,N_20764,N_20215);
xnor U21798 (N_21798,N_20885,N_20156);
nor U21799 (N_21799,N_20462,N_20377);
nor U21800 (N_21800,N_20914,N_20066);
and U21801 (N_21801,N_20591,N_20498);
and U21802 (N_21802,N_20642,N_20048);
nor U21803 (N_21803,N_20983,N_20362);
nor U21804 (N_21804,N_20944,N_20637);
nand U21805 (N_21805,N_20547,N_20809);
nor U21806 (N_21806,N_20657,N_20981);
and U21807 (N_21807,N_20545,N_20742);
xnor U21808 (N_21808,N_20544,N_20158);
xnor U21809 (N_21809,N_20217,N_20953);
xnor U21810 (N_21810,N_20054,N_20218);
nor U21811 (N_21811,N_20175,N_20971);
nand U21812 (N_21812,N_20430,N_20171);
and U21813 (N_21813,N_20754,N_20962);
nand U21814 (N_21814,N_20568,N_20014);
nand U21815 (N_21815,N_20851,N_20124);
or U21816 (N_21816,N_20068,N_20594);
and U21817 (N_21817,N_20010,N_20786);
and U21818 (N_21818,N_20700,N_20231);
xor U21819 (N_21819,N_20845,N_20766);
xnor U21820 (N_21820,N_20276,N_20503);
and U21821 (N_21821,N_20644,N_20805);
and U21822 (N_21822,N_20896,N_20602);
or U21823 (N_21823,N_20223,N_20144);
nor U21824 (N_21824,N_20168,N_20719);
and U21825 (N_21825,N_20919,N_20793);
and U21826 (N_21826,N_20515,N_20019);
and U21827 (N_21827,N_20329,N_20861);
or U21828 (N_21828,N_20040,N_20212);
or U21829 (N_21829,N_20514,N_20912);
and U21830 (N_21830,N_20026,N_20810);
nand U21831 (N_21831,N_20846,N_20695);
and U21832 (N_21832,N_20953,N_20353);
xnor U21833 (N_21833,N_20335,N_20318);
and U21834 (N_21834,N_20512,N_20966);
and U21835 (N_21835,N_20990,N_20227);
xnor U21836 (N_21836,N_20344,N_20874);
xnor U21837 (N_21837,N_20770,N_20634);
nand U21838 (N_21838,N_20177,N_20472);
nand U21839 (N_21839,N_20954,N_20000);
xnor U21840 (N_21840,N_20391,N_20519);
and U21841 (N_21841,N_20541,N_20718);
xor U21842 (N_21842,N_20592,N_20051);
or U21843 (N_21843,N_20962,N_20667);
nor U21844 (N_21844,N_20517,N_20393);
and U21845 (N_21845,N_20261,N_20342);
nor U21846 (N_21846,N_20713,N_20394);
nand U21847 (N_21847,N_20942,N_20396);
xnor U21848 (N_21848,N_20439,N_20269);
and U21849 (N_21849,N_20528,N_20558);
nand U21850 (N_21850,N_20084,N_20748);
or U21851 (N_21851,N_20009,N_20260);
and U21852 (N_21852,N_20865,N_20696);
nor U21853 (N_21853,N_20236,N_20314);
nand U21854 (N_21854,N_20318,N_20342);
xnor U21855 (N_21855,N_20566,N_20791);
nor U21856 (N_21856,N_20946,N_20435);
or U21857 (N_21857,N_20939,N_20605);
or U21858 (N_21858,N_20538,N_20697);
nor U21859 (N_21859,N_20367,N_20817);
nand U21860 (N_21860,N_20429,N_20883);
or U21861 (N_21861,N_20080,N_20715);
nor U21862 (N_21862,N_20748,N_20248);
or U21863 (N_21863,N_20750,N_20286);
and U21864 (N_21864,N_20066,N_20373);
xnor U21865 (N_21865,N_20058,N_20275);
xnor U21866 (N_21866,N_20813,N_20900);
nor U21867 (N_21867,N_20075,N_20015);
or U21868 (N_21868,N_20108,N_20596);
nor U21869 (N_21869,N_20827,N_20533);
nand U21870 (N_21870,N_20005,N_20096);
xor U21871 (N_21871,N_20967,N_20237);
and U21872 (N_21872,N_20987,N_20580);
and U21873 (N_21873,N_20456,N_20352);
and U21874 (N_21874,N_20470,N_20579);
or U21875 (N_21875,N_20006,N_20900);
or U21876 (N_21876,N_20907,N_20054);
nor U21877 (N_21877,N_20835,N_20323);
and U21878 (N_21878,N_20610,N_20611);
and U21879 (N_21879,N_20295,N_20408);
nor U21880 (N_21880,N_20601,N_20388);
nor U21881 (N_21881,N_20805,N_20383);
and U21882 (N_21882,N_20420,N_20682);
and U21883 (N_21883,N_20186,N_20110);
and U21884 (N_21884,N_20118,N_20984);
nor U21885 (N_21885,N_20289,N_20220);
nor U21886 (N_21886,N_20833,N_20526);
and U21887 (N_21887,N_20075,N_20470);
xor U21888 (N_21888,N_20430,N_20330);
nand U21889 (N_21889,N_20885,N_20879);
nor U21890 (N_21890,N_20063,N_20610);
nand U21891 (N_21891,N_20735,N_20420);
xnor U21892 (N_21892,N_20130,N_20775);
and U21893 (N_21893,N_20102,N_20471);
or U21894 (N_21894,N_20883,N_20896);
nor U21895 (N_21895,N_20219,N_20150);
and U21896 (N_21896,N_20989,N_20173);
or U21897 (N_21897,N_20861,N_20800);
or U21898 (N_21898,N_20940,N_20841);
and U21899 (N_21899,N_20052,N_20003);
or U21900 (N_21900,N_20498,N_20634);
nor U21901 (N_21901,N_20922,N_20598);
nand U21902 (N_21902,N_20710,N_20577);
and U21903 (N_21903,N_20716,N_20646);
nor U21904 (N_21904,N_20999,N_20505);
nor U21905 (N_21905,N_20555,N_20410);
or U21906 (N_21906,N_20283,N_20900);
xor U21907 (N_21907,N_20240,N_20999);
and U21908 (N_21908,N_20797,N_20433);
nand U21909 (N_21909,N_20470,N_20929);
or U21910 (N_21910,N_20681,N_20298);
xor U21911 (N_21911,N_20213,N_20425);
nand U21912 (N_21912,N_20959,N_20623);
and U21913 (N_21913,N_20219,N_20264);
or U21914 (N_21914,N_20759,N_20758);
nor U21915 (N_21915,N_20228,N_20907);
and U21916 (N_21916,N_20939,N_20023);
or U21917 (N_21917,N_20271,N_20735);
and U21918 (N_21918,N_20156,N_20442);
nand U21919 (N_21919,N_20611,N_20244);
and U21920 (N_21920,N_20351,N_20726);
and U21921 (N_21921,N_20894,N_20566);
and U21922 (N_21922,N_20876,N_20773);
nor U21923 (N_21923,N_20941,N_20351);
and U21924 (N_21924,N_20964,N_20151);
and U21925 (N_21925,N_20530,N_20001);
nor U21926 (N_21926,N_20344,N_20132);
nor U21927 (N_21927,N_20694,N_20463);
or U21928 (N_21928,N_20133,N_20614);
xor U21929 (N_21929,N_20463,N_20590);
nand U21930 (N_21930,N_20498,N_20078);
nor U21931 (N_21931,N_20887,N_20776);
and U21932 (N_21932,N_20638,N_20839);
or U21933 (N_21933,N_20600,N_20243);
nor U21934 (N_21934,N_20806,N_20140);
nor U21935 (N_21935,N_20322,N_20291);
and U21936 (N_21936,N_20091,N_20027);
or U21937 (N_21937,N_20528,N_20458);
or U21938 (N_21938,N_20570,N_20597);
xnor U21939 (N_21939,N_20352,N_20415);
nor U21940 (N_21940,N_20289,N_20070);
and U21941 (N_21941,N_20799,N_20655);
nor U21942 (N_21942,N_20950,N_20586);
and U21943 (N_21943,N_20476,N_20311);
or U21944 (N_21944,N_20925,N_20930);
xnor U21945 (N_21945,N_20476,N_20833);
nand U21946 (N_21946,N_20281,N_20722);
xor U21947 (N_21947,N_20562,N_20556);
xnor U21948 (N_21948,N_20253,N_20528);
nand U21949 (N_21949,N_20618,N_20221);
nand U21950 (N_21950,N_20406,N_20135);
or U21951 (N_21951,N_20423,N_20322);
or U21952 (N_21952,N_20829,N_20653);
or U21953 (N_21953,N_20509,N_20347);
nor U21954 (N_21954,N_20937,N_20132);
xor U21955 (N_21955,N_20583,N_20802);
and U21956 (N_21956,N_20899,N_20540);
and U21957 (N_21957,N_20822,N_20557);
or U21958 (N_21958,N_20651,N_20981);
xnor U21959 (N_21959,N_20692,N_20667);
nand U21960 (N_21960,N_20012,N_20648);
or U21961 (N_21961,N_20857,N_20416);
nand U21962 (N_21962,N_20107,N_20303);
nor U21963 (N_21963,N_20859,N_20974);
nand U21964 (N_21964,N_20494,N_20280);
and U21965 (N_21965,N_20653,N_20630);
and U21966 (N_21966,N_20618,N_20875);
and U21967 (N_21967,N_20536,N_20487);
nand U21968 (N_21968,N_20351,N_20673);
and U21969 (N_21969,N_20430,N_20143);
xor U21970 (N_21970,N_20383,N_20077);
xor U21971 (N_21971,N_20155,N_20919);
nand U21972 (N_21972,N_20073,N_20048);
or U21973 (N_21973,N_20171,N_20691);
and U21974 (N_21974,N_20066,N_20288);
nor U21975 (N_21975,N_20527,N_20578);
and U21976 (N_21976,N_20425,N_20341);
xor U21977 (N_21977,N_20647,N_20000);
nand U21978 (N_21978,N_20519,N_20556);
or U21979 (N_21979,N_20714,N_20126);
xnor U21980 (N_21980,N_20303,N_20046);
nand U21981 (N_21981,N_20797,N_20836);
xor U21982 (N_21982,N_20075,N_20149);
nor U21983 (N_21983,N_20978,N_20610);
xor U21984 (N_21984,N_20944,N_20503);
xnor U21985 (N_21985,N_20509,N_20480);
or U21986 (N_21986,N_20752,N_20313);
nor U21987 (N_21987,N_20451,N_20290);
or U21988 (N_21988,N_20074,N_20865);
or U21989 (N_21989,N_20308,N_20001);
and U21990 (N_21990,N_20202,N_20255);
and U21991 (N_21991,N_20799,N_20462);
or U21992 (N_21992,N_20520,N_20710);
and U21993 (N_21993,N_20229,N_20368);
or U21994 (N_21994,N_20459,N_20919);
xor U21995 (N_21995,N_20989,N_20700);
and U21996 (N_21996,N_20179,N_20940);
nor U21997 (N_21997,N_20954,N_20870);
nor U21998 (N_21998,N_20592,N_20667);
xnor U21999 (N_21999,N_20283,N_20783);
xnor U22000 (N_22000,N_21769,N_21980);
or U22001 (N_22001,N_21312,N_21317);
nand U22002 (N_22002,N_21437,N_21793);
and U22003 (N_22003,N_21589,N_21081);
and U22004 (N_22004,N_21920,N_21994);
nand U22005 (N_22005,N_21204,N_21785);
or U22006 (N_22006,N_21502,N_21251);
xnor U22007 (N_22007,N_21211,N_21135);
xnor U22008 (N_22008,N_21602,N_21756);
nand U22009 (N_22009,N_21051,N_21588);
and U22010 (N_22010,N_21667,N_21885);
xnor U22011 (N_22011,N_21604,N_21388);
nand U22012 (N_22012,N_21201,N_21596);
nand U22013 (N_22013,N_21150,N_21877);
nand U22014 (N_22014,N_21361,N_21291);
and U22015 (N_22015,N_21083,N_21727);
and U22016 (N_22016,N_21503,N_21273);
and U22017 (N_22017,N_21746,N_21630);
nor U22018 (N_22018,N_21780,N_21940);
nand U22019 (N_22019,N_21024,N_21278);
nand U22020 (N_22020,N_21640,N_21322);
nand U22021 (N_22021,N_21360,N_21028);
nor U22022 (N_22022,N_21035,N_21993);
nand U22023 (N_22023,N_21040,N_21709);
xnor U22024 (N_22024,N_21260,N_21538);
nor U22025 (N_22025,N_21900,N_21315);
or U22026 (N_22026,N_21745,N_21944);
nand U22027 (N_22027,N_21334,N_21364);
and U22028 (N_22028,N_21883,N_21753);
nand U22029 (N_22029,N_21698,N_21832);
nand U22030 (N_22030,N_21782,N_21678);
nor U22031 (N_22031,N_21850,N_21449);
nor U22032 (N_22032,N_21916,N_21326);
or U22033 (N_22033,N_21122,N_21776);
nor U22034 (N_22034,N_21608,N_21348);
and U22035 (N_22035,N_21929,N_21359);
xor U22036 (N_22036,N_21739,N_21510);
nor U22037 (N_22037,N_21959,N_21610);
or U22038 (N_22038,N_21127,N_21844);
and U22039 (N_22039,N_21455,N_21418);
or U22040 (N_22040,N_21297,N_21012);
nor U22041 (N_22041,N_21060,N_21209);
nand U22042 (N_22042,N_21728,N_21740);
nor U22043 (N_22043,N_21521,N_21501);
xor U22044 (N_22044,N_21622,N_21332);
nor U22045 (N_22045,N_21186,N_21705);
and U22046 (N_22046,N_21659,N_21718);
nand U22047 (N_22047,N_21500,N_21970);
nor U22048 (N_22048,N_21385,N_21473);
xnor U22049 (N_22049,N_21077,N_21446);
nor U22050 (N_22050,N_21025,N_21898);
nand U22051 (N_22051,N_21719,N_21380);
or U22052 (N_22052,N_21232,N_21631);
nor U22053 (N_22053,N_21813,N_21258);
nor U22054 (N_22054,N_21091,N_21629);
nand U22055 (N_22055,N_21062,N_21262);
nor U22056 (N_22056,N_21654,N_21400);
nand U22057 (N_22057,N_21316,N_21816);
nand U22058 (N_22058,N_21600,N_21003);
xor U22059 (N_22059,N_21442,N_21810);
and U22060 (N_22060,N_21223,N_21457);
xor U22061 (N_22061,N_21242,N_21568);
or U22062 (N_22062,N_21427,N_21528);
or U22063 (N_22063,N_21218,N_21264);
nand U22064 (N_22064,N_21915,N_21021);
or U22065 (N_22065,N_21178,N_21912);
nand U22066 (N_22066,N_21147,N_21982);
nor U22067 (N_22067,N_21206,N_21445);
and U22068 (N_22068,N_21107,N_21389);
or U22069 (N_22069,N_21814,N_21358);
or U22070 (N_22070,N_21742,N_21914);
or U22071 (N_22071,N_21013,N_21737);
nor U22072 (N_22072,N_21639,N_21027);
or U22073 (N_22073,N_21493,N_21414);
or U22074 (N_22074,N_21807,N_21868);
nor U22075 (N_22075,N_21398,N_21078);
xor U22076 (N_22076,N_21646,N_21839);
nand U22077 (N_22077,N_21975,N_21430);
and U22078 (N_22078,N_21717,N_21625);
or U22079 (N_22079,N_21517,N_21570);
xor U22080 (N_22080,N_21365,N_21979);
or U22081 (N_22081,N_21489,N_21046);
or U22082 (N_22082,N_21231,N_21461);
nor U22083 (N_22083,N_21536,N_21840);
nand U22084 (N_22084,N_21886,N_21221);
nand U22085 (N_22085,N_21137,N_21843);
nand U22086 (N_22086,N_21955,N_21567);
xnor U22087 (N_22087,N_21601,N_21337);
nor U22088 (N_22088,N_21302,N_21309);
nand U22089 (N_22089,N_21664,N_21349);
nand U22090 (N_22090,N_21061,N_21274);
and U22091 (N_22091,N_21887,N_21675);
or U22092 (N_22092,N_21762,N_21324);
nor U22093 (N_22093,N_21464,N_21587);
and U22094 (N_22094,N_21577,N_21965);
nor U22095 (N_22095,N_21269,N_21421);
and U22096 (N_22096,N_21874,N_21121);
or U22097 (N_22097,N_21339,N_21833);
or U22098 (N_22098,N_21645,N_21954);
nor U22099 (N_22099,N_21633,N_21956);
or U22100 (N_22100,N_21634,N_21628);
and U22101 (N_22101,N_21522,N_21275);
xnor U22102 (N_22102,N_21548,N_21961);
and U22103 (N_22103,N_21544,N_21376);
or U22104 (N_22104,N_21058,N_21243);
or U22105 (N_22105,N_21110,N_21809);
nand U22106 (N_22106,N_21808,N_21722);
nand U22107 (N_22107,N_21561,N_21716);
or U22108 (N_22108,N_21171,N_21197);
or U22109 (N_22109,N_21476,N_21902);
or U22110 (N_22110,N_21619,N_21736);
or U22111 (N_22111,N_21084,N_21069);
nand U22112 (N_22112,N_21882,N_21781);
and U22113 (N_22113,N_21116,N_21155);
nor U22114 (N_22114,N_21656,N_21199);
and U22115 (N_22115,N_21163,N_21164);
nand U22116 (N_22116,N_21165,N_21922);
and U22117 (N_22117,N_21448,N_21525);
and U22118 (N_22118,N_21347,N_21276);
nor U22119 (N_22119,N_21946,N_21866);
or U22120 (N_22120,N_21724,N_21194);
or U22121 (N_22121,N_21233,N_21033);
nand U22122 (N_22122,N_21255,N_21837);
nor U22123 (N_22123,N_21114,N_21344);
or U22124 (N_22124,N_21237,N_21647);
nor U22125 (N_22125,N_21524,N_21225);
or U22126 (N_22126,N_21481,N_21370);
or U22127 (N_22127,N_21512,N_21001);
and U22128 (N_22128,N_21498,N_21362);
or U22129 (N_22129,N_21168,N_21467);
xor U22130 (N_22130,N_21950,N_21649);
nand U22131 (N_22131,N_21182,N_21087);
nor U22132 (N_22132,N_21433,N_21265);
xor U22133 (N_22133,N_21226,N_21465);
xor U22134 (N_22134,N_21353,N_21227);
nand U22135 (N_22135,N_21638,N_21969);
or U22136 (N_22136,N_21185,N_21937);
and U22137 (N_22137,N_21609,N_21008);
nand U22138 (N_22138,N_21469,N_21945);
or U22139 (N_22139,N_21824,N_21540);
or U22140 (N_22140,N_21917,N_21890);
nand U22141 (N_22141,N_21410,N_21170);
or U22142 (N_22142,N_21997,N_21801);
or U22143 (N_22143,N_21686,N_21118);
and U22144 (N_22144,N_21098,N_21637);
nand U22145 (N_22145,N_21141,N_21848);
nor U22146 (N_22146,N_21819,N_21751);
and U22147 (N_22147,N_21603,N_21558);
or U22148 (N_22148,N_21838,N_21531);
nand U22149 (N_22149,N_21779,N_21803);
and U22150 (N_22150,N_21962,N_21597);
nor U22151 (N_22151,N_21599,N_21173);
and U22152 (N_22152,N_21766,N_21342);
and U22153 (N_22153,N_21372,N_21188);
nor U22154 (N_22154,N_21142,N_21787);
or U22155 (N_22155,N_21552,N_21918);
or U22156 (N_22156,N_21723,N_21483);
nor U22157 (N_22157,N_21303,N_21933);
nand U22158 (N_22158,N_21384,N_21484);
xnor U22159 (N_22159,N_21480,N_21909);
nand U22160 (N_22160,N_21331,N_21492);
xor U22161 (N_22161,N_21574,N_21055);
and U22162 (N_22162,N_21156,N_21229);
xnor U22163 (N_22163,N_21714,N_21180);
or U22164 (N_22164,N_21829,N_21554);
nor U22165 (N_22165,N_21191,N_21123);
xnor U22166 (N_22166,N_21113,N_21845);
nor U22167 (N_22167,N_21236,N_21126);
or U22168 (N_22168,N_21093,N_21771);
and U22169 (N_22169,N_21879,N_21875);
nor U22170 (N_22170,N_21439,N_21487);
nor U22171 (N_22171,N_21624,N_21715);
or U22172 (N_22172,N_21470,N_21863);
nor U22173 (N_22173,N_21054,N_21261);
nor U22174 (N_22174,N_21131,N_21249);
xor U22175 (N_22175,N_21905,N_21726);
and U22176 (N_22176,N_21246,N_21973);
and U22177 (N_22177,N_21452,N_21202);
nor U22178 (N_22178,N_21862,N_21856);
xnor U22179 (N_22179,N_21660,N_21284);
nor U22180 (N_22180,N_21669,N_21217);
nor U22181 (N_22181,N_21230,N_21496);
and U22182 (N_22182,N_21674,N_21108);
nand U22183 (N_22183,N_21125,N_21318);
and U22184 (N_22184,N_21533,N_21541);
and U22185 (N_22185,N_21795,N_21402);
xnor U22186 (N_22186,N_21696,N_21611);
or U22187 (N_22187,N_21958,N_21689);
xor U22188 (N_22188,N_21263,N_21311);
or U22189 (N_22189,N_21403,N_21778);
nand U22190 (N_22190,N_21507,N_21774);
xor U22191 (N_22191,N_21636,N_21187);
or U22192 (N_22192,N_21578,N_21450);
nand U22193 (N_22193,N_21352,N_21042);
or U22194 (N_22194,N_21468,N_21132);
nor U22195 (N_22195,N_21495,N_21010);
nand U22196 (N_22196,N_21394,N_21749);
xor U22197 (N_22197,N_21878,N_21466);
nand U22198 (N_22198,N_21009,N_21295);
nand U22199 (N_22199,N_21148,N_21555);
xnor U22200 (N_22200,N_21157,N_21546);
nand U22201 (N_22201,N_21030,N_21786);
nor U22202 (N_22202,N_21831,N_21151);
nand U22203 (N_22203,N_21576,N_21934);
xnor U22204 (N_22204,N_21189,N_21300);
nor U22205 (N_22205,N_21992,N_21072);
xor U22206 (N_22206,N_21444,N_21880);
and U22207 (N_22207,N_21330,N_21989);
nor U22208 (N_22208,N_21901,N_21612);
nand U22209 (N_22209,N_21579,N_21802);
and U22210 (N_22210,N_21953,N_21712);
nor U22211 (N_22211,N_21938,N_21685);
and U22212 (N_22212,N_21732,N_21981);
nand U22213 (N_22213,N_21591,N_21161);
or U22214 (N_22214,N_21984,N_21543);
nor U22215 (N_22215,N_21535,N_21420);
or U22216 (N_22216,N_21090,N_21289);
or U22217 (N_22217,N_21998,N_21671);
xor U22218 (N_22218,N_21143,N_21569);
or U22219 (N_22219,N_21635,N_21064);
nor U22220 (N_22220,N_21508,N_21662);
nand U22221 (N_22221,N_21144,N_21595);
xor U22222 (N_22222,N_21505,N_21089);
xnor U22223 (N_22223,N_21436,N_21852);
nand U22224 (N_22224,N_21710,N_21499);
nor U22225 (N_22225,N_21690,N_21767);
xor U22226 (N_22226,N_21488,N_21799);
or U22227 (N_22227,N_21212,N_21294);
and U22228 (N_22228,N_21458,N_21811);
nand U22229 (N_22229,N_21818,N_21516);
nand U22230 (N_22230,N_21826,N_21205);
nand U22231 (N_22231,N_21725,N_21057);
and U22232 (N_22232,N_21351,N_21566);
nand U22233 (N_22233,N_21438,N_21704);
nor U22234 (N_22234,N_21872,N_21523);
nand U22235 (N_22235,N_21575,N_21415);
nor U22236 (N_22236,N_21124,N_21584);
nor U22237 (N_22237,N_21419,N_21085);
or U22238 (N_22238,N_21680,N_21004);
and U22239 (N_22239,N_21082,N_21834);
and U22240 (N_22240,N_21999,N_21477);
nand U22241 (N_22241,N_21293,N_21235);
nor U22242 (N_22242,N_21748,N_21247);
and U22243 (N_22243,N_21412,N_21471);
nand U22244 (N_22244,N_21643,N_21172);
or U22245 (N_22245,N_21429,N_21744);
or U22246 (N_22246,N_21299,N_21853);
nand U22247 (N_22247,N_21830,N_21677);
and U22248 (N_22248,N_21043,N_21514);
xnor U22249 (N_22249,N_21277,N_21286);
or U22250 (N_22250,N_21272,N_21198);
xnor U22251 (N_22251,N_21397,N_21153);
or U22252 (N_22252,N_21960,N_21195);
xor U22253 (N_22253,N_21386,N_21063);
and U22254 (N_22254,N_21932,N_21908);
and U22255 (N_22255,N_21310,N_21582);
and U22256 (N_22256,N_21821,N_21738);
and U22257 (N_22257,N_21335,N_21149);
xor U22258 (N_22258,N_21478,N_21761);
nand U22259 (N_22259,N_21513,N_21943);
nor U22260 (N_22260,N_21177,N_21250);
and U22261 (N_22261,N_21426,N_21134);
nor U22262 (N_22262,N_21621,N_21383);
xnor U22263 (N_22263,N_21256,N_21836);
nand U22264 (N_22264,N_21045,N_21655);
or U22265 (N_22265,N_21102,N_21099);
nand U22266 (N_22266,N_21129,N_21325);
xor U22267 (N_22267,N_21020,N_21976);
nor U22268 (N_22268,N_21941,N_21354);
xor U22269 (N_22269,N_21765,N_21565);
nor U22270 (N_22270,N_21861,N_21720);
and U22271 (N_22271,N_21835,N_21571);
or U22272 (N_22272,N_21416,N_21530);
nor U22273 (N_22273,N_21443,N_21699);
or U22274 (N_22274,N_21983,N_21292);
nand U22275 (N_22275,N_21367,N_21340);
nor U22276 (N_22276,N_21592,N_21889);
nor U22277 (N_22277,N_21788,N_21755);
xnor U22278 (N_22278,N_21563,N_21296);
and U22279 (N_22279,N_21447,N_21606);
xnor U22280 (N_22280,N_21697,N_21796);
or U22281 (N_22281,N_21894,N_21891);
or U22282 (N_22282,N_21893,N_21036);
nor U22283 (N_22283,N_21871,N_21949);
or U22284 (N_22284,N_21648,N_21130);
nand U22285 (N_22285,N_21580,N_21391);
xnor U22286 (N_22286,N_21138,N_21849);
nor U22287 (N_22287,N_21708,N_21381);
xnor U22288 (N_22288,N_21100,N_21537);
nor U22289 (N_22289,N_21996,N_21103);
and U22290 (N_22290,N_21074,N_21752);
nor U22291 (N_22291,N_21822,N_21076);
or U22292 (N_22292,N_21392,N_21721);
nor U22293 (N_22293,N_21313,N_21551);
nand U22294 (N_22294,N_21355,N_21080);
xnor U22295 (N_22295,N_21966,N_21038);
xnor U22296 (N_22296,N_21870,N_21145);
nand U22297 (N_22297,N_21271,N_21120);
and U22298 (N_22298,N_21701,N_21482);
xor U22299 (N_22299,N_21390,N_21401);
nor U22300 (N_22300,N_21991,N_21166);
or U22301 (N_22301,N_21518,N_21146);
nand U22302 (N_22302,N_21456,N_21181);
and U22303 (N_22303,N_21693,N_21928);
xor U22304 (N_22304,N_21015,N_21096);
nor U22305 (N_22305,N_21428,N_21176);
nand U22306 (N_22306,N_21216,N_21101);
or U22307 (N_22307,N_21935,N_21616);
xor U22308 (N_22308,N_21346,N_21865);
and U22309 (N_22309,N_21474,N_21179);
xnor U22310 (N_22310,N_21930,N_21435);
or U22311 (N_22311,N_21222,N_21684);
or U22312 (N_22312,N_21618,N_21408);
and U22313 (N_22313,N_21692,N_21486);
or U22314 (N_22314,N_21159,N_21773);
nand U22315 (N_22315,N_21881,N_21792);
xor U22316 (N_22316,N_21343,N_21174);
and U22317 (N_22317,N_21208,N_21073);
xor U22318 (N_22318,N_21658,N_21549);
and U22319 (N_22319,N_21282,N_21425);
or U22320 (N_22320,N_21651,N_21632);
and U22321 (N_22321,N_21963,N_21356);
nor U22322 (N_22322,N_21193,N_21985);
nor U22323 (N_22323,N_21519,N_21133);
and U22324 (N_22324,N_21037,N_21244);
or U22325 (N_22325,N_21441,N_21534);
xnor U22326 (N_22326,N_21047,N_21504);
xnor U22327 (N_22327,N_21192,N_21184);
xnor U22328 (N_22328,N_21884,N_21497);
nand U22329 (N_22329,N_21097,N_21210);
or U22330 (N_22330,N_21283,N_21104);
nand U22331 (N_22331,N_21931,N_21775);
nor U22332 (N_22332,N_21019,N_21014);
nor U22333 (N_22333,N_21238,N_21615);
or U22334 (N_22334,N_21321,N_21770);
and U22335 (N_22335,N_21735,N_21105);
nor U22336 (N_22336,N_21140,N_21215);
xor U22337 (N_22337,N_21371,N_21424);
nand U22338 (N_22338,N_21128,N_21759);
xnor U22339 (N_22339,N_21196,N_21338);
xnor U22340 (N_22340,N_21368,N_21016);
or U22341 (N_22341,N_21911,N_21828);
and U22342 (N_22342,N_21617,N_21784);
and U22343 (N_22343,N_21031,N_21079);
and U22344 (N_22344,N_21298,N_21373);
nand U22345 (N_22345,N_21657,N_21017);
xnor U22346 (N_22346,N_21026,N_21494);
and U22347 (N_22347,N_21220,N_21942);
nand U22348 (N_22348,N_21422,N_21254);
and U22349 (N_22349,N_21924,N_21453);
or U22350 (N_22350,N_21075,N_21094);
or U22351 (N_22351,N_21794,N_21048);
nand U22352 (N_22352,N_21404,N_21268);
nand U22353 (N_22353,N_21764,N_21320);
xnor U22354 (N_22354,N_21305,N_21864);
and U22355 (N_22355,N_21903,N_21772);
nand U22356 (N_22356,N_21406,N_21234);
nor U22357 (N_22357,N_21252,N_21539);
xnor U22358 (N_22358,N_21066,N_21224);
nand U22359 (N_22359,N_21323,N_21253);
nor U22360 (N_22360,N_21357,N_21855);
nand U22361 (N_22361,N_21377,N_21023);
and U22362 (N_22362,N_21396,N_21627);
nand U22363 (N_22363,N_21594,N_21741);
nor U22364 (N_22364,N_21266,N_21672);
xor U22365 (N_22365,N_21641,N_21183);
or U22366 (N_22366,N_21379,N_21395);
nor U22367 (N_22367,N_21964,N_21053);
nor U22368 (N_22368,N_21842,N_21411);
xnor U22369 (N_22369,N_21827,N_21586);
nor U22370 (N_22370,N_21939,N_21977);
and U22371 (N_22371,N_21666,N_21022);
xor U22372 (N_22372,N_21713,N_21515);
or U22373 (N_22373,N_21650,N_21859);
or U22374 (N_22374,N_21434,N_21694);
or U22375 (N_22375,N_21460,N_21175);
nand U22376 (N_22376,N_21306,N_21095);
xnor U22377 (N_22377,N_21613,N_21162);
nor U22378 (N_22378,N_21729,N_21440);
nand U22379 (N_22379,N_21511,N_21590);
or U22380 (N_22380,N_21585,N_21791);
xnor U22381 (N_22381,N_21583,N_21919);
and U22382 (N_22382,N_21169,N_21869);
and U22383 (N_22383,N_21923,N_21070);
and U22384 (N_22384,N_21988,N_21413);
nand U22385 (N_22385,N_21860,N_21279);
nand U22386 (N_22386,N_21490,N_21896);
nor U22387 (N_22387,N_21858,N_21851);
or U22388 (N_22388,N_21327,N_21547);
or U22389 (N_22389,N_21812,N_21730);
and U22390 (N_22390,N_21971,N_21280);
or U22391 (N_22391,N_21270,N_21581);
or U22392 (N_22392,N_21550,N_21319);
nor U22393 (N_22393,N_21947,N_21329);
xnor U22394 (N_22394,N_21387,N_21707);
xor U22395 (N_22395,N_21951,N_21910);
nand U22396 (N_22396,N_21783,N_21068);
and U22397 (N_22397,N_21806,N_21032);
or U22398 (N_22398,N_21207,N_21065);
nand U22399 (N_22399,N_21854,N_21995);
nor U22400 (N_22400,N_21542,N_21560);
and U22401 (N_22401,N_21899,N_21366);
nand U22402 (N_22402,N_21620,N_21248);
and U22403 (N_22403,N_21768,N_21451);
or U22404 (N_22404,N_21825,N_21239);
and U22405 (N_22405,N_21459,N_21614);
xnor U22406 (N_22406,N_21086,N_21763);
nand U22407 (N_22407,N_21341,N_21990);
and U22408 (N_22408,N_21805,N_21847);
and U22409 (N_22409,N_21369,N_21287);
nand U22410 (N_22410,N_21158,N_21846);
xnor U22411 (N_22411,N_21423,N_21154);
nand U22412 (N_22412,N_21691,N_21485);
xnor U22413 (N_22413,N_21049,N_21041);
or U22414 (N_22414,N_21472,N_21733);
nor U22415 (N_22415,N_21867,N_21000);
xor U22416 (N_22416,N_21245,N_21703);
and U22417 (N_22417,N_21475,N_21029);
nand U22418 (N_22418,N_21559,N_21820);
and U22419 (N_22419,N_21407,N_21463);
nor U22420 (N_22420,N_21006,N_21823);
nand U22421 (N_22421,N_21350,N_21405);
nor U22422 (N_22422,N_21986,N_21607);
or U22423 (N_22423,N_21797,N_21545);
nor U22424 (N_22424,N_21112,N_21160);
nand U22425 (N_22425,N_21683,N_21532);
or U22426 (N_22426,N_21240,N_21375);
xnor U22427 (N_22427,N_21479,N_21876);
xor U22428 (N_22428,N_21167,N_21743);
nand U22429 (N_22429,N_21007,N_21681);
and U22430 (N_22430,N_21092,N_21071);
xor U22431 (N_22431,N_21241,N_21301);
xnor U22432 (N_22432,N_21978,N_21790);
nand U22433 (N_22433,N_21682,N_21213);
nor U22434 (N_22434,N_21598,N_21815);
or U22435 (N_22435,N_21925,N_21661);
xor U22436 (N_22436,N_21011,N_21152);
or U22437 (N_22437,N_21926,N_21052);
or U22438 (N_22438,N_21409,N_21564);
or U22439 (N_22439,N_21431,N_21777);
nand U22440 (N_22440,N_21139,N_21281);
or U22441 (N_22441,N_21626,N_21623);
nand U22442 (N_22442,N_21257,N_21314);
and U22443 (N_22443,N_21804,N_21593);
or U22444 (N_22444,N_21904,N_21927);
and U22445 (N_22445,N_21288,N_21670);
or U22446 (N_22446,N_21018,N_21382);
nand U22447 (N_22447,N_21800,N_21760);
nor U22448 (N_22448,N_21203,N_21688);
or U22449 (N_22449,N_21747,N_21734);
and U22450 (N_22450,N_21378,N_21228);
or U22451 (N_22451,N_21115,N_21967);
nand U22452 (N_22452,N_21034,N_21817);
xnor U22453 (N_22453,N_21557,N_21957);
nand U22454 (N_22454,N_21679,N_21374);
nor U22455 (N_22455,N_21921,N_21285);
nand U22456 (N_22456,N_21948,N_21111);
and U22457 (N_22457,N_21892,N_21527);
or U22458 (N_22458,N_21039,N_21290);
or U22459 (N_22459,N_21758,N_21754);
xnor U22460 (N_22460,N_21706,N_21336);
nor U22461 (N_22461,N_21987,N_21750);
or U22462 (N_22462,N_21259,N_21642);
nor U22463 (N_22463,N_21906,N_21462);
or U22464 (N_22464,N_21731,N_21067);
nor U22465 (N_22465,N_21328,N_21572);
nor U22466 (N_22466,N_21700,N_21644);
nor U22467 (N_22467,N_21873,N_21002);
nor U22468 (N_22468,N_21219,N_21562);
xnor U22469 (N_22469,N_21556,N_21044);
xor U22470 (N_22470,N_21454,N_21702);
or U22471 (N_22471,N_21695,N_21895);
nand U22472 (N_22472,N_21972,N_21897);
xor U22473 (N_22473,N_21857,N_21757);
nor U22474 (N_22474,N_21665,N_21907);
nor U22475 (N_22475,N_21307,N_21050);
or U22476 (N_22476,N_21117,N_21399);
nand U22477 (N_22477,N_21393,N_21304);
and U22478 (N_22478,N_21553,N_21789);
or U22479 (N_22479,N_21520,N_21432);
or U22480 (N_22480,N_21652,N_21056);
and U22481 (N_22481,N_21509,N_21059);
nand U22482 (N_22482,N_21363,N_21200);
nand U22483 (N_22483,N_21136,N_21668);
xnor U22484 (N_22484,N_21109,N_21267);
nand U22485 (N_22485,N_21190,N_21663);
nand U22486 (N_22486,N_21506,N_21529);
and U22487 (N_22487,N_21308,N_21974);
nand U22488 (N_22488,N_21106,N_21888);
and U22489 (N_22489,N_21653,N_21005);
or U22490 (N_22490,N_21605,N_21345);
nand U22491 (N_22491,N_21968,N_21913);
and U22492 (N_22492,N_21676,N_21526);
xnor U22493 (N_22493,N_21088,N_21491);
and U22494 (N_22494,N_21333,N_21936);
nand U22495 (N_22495,N_21417,N_21214);
or U22496 (N_22496,N_21673,N_21841);
and U22497 (N_22497,N_21119,N_21573);
nand U22498 (N_22498,N_21711,N_21798);
nand U22499 (N_22499,N_21687,N_21952);
xor U22500 (N_22500,N_21554,N_21934);
nand U22501 (N_22501,N_21531,N_21877);
and U22502 (N_22502,N_21267,N_21245);
nor U22503 (N_22503,N_21604,N_21509);
and U22504 (N_22504,N_21266,N_21696);
or U22505 (N_22505,N_21286,N_21723);
or U22506 (N_22506,N_21274,N_21604);
or U22507 (N_22507,N_21043,N_21126);
and U22508 (N_22508,N_21884,N_21459);
and U22509 (N_22509,N_21412,N_21936);
or U22510 (N_22510,N_21266,N_21311);
and U22511 (N_22511,N_21275,N_21878);
nand U22512 (N_22512,N_21826,N_21990);
nor U22513 (N_22513,N_21761,N_21556);
nand U22514 (N_22514,N_21842,N_21646);
xor U22515 (N_22515,N_21394,N_21946);
or U22516 (N_22516,N_21851,N_21586);
and U22517 (N_22517,N_21496,N_21844);
or U22518 (N_22518,N_21238,N_21626);
nor U22519 (N_22519,N_21686,N_21707);
and U22520 (N_22520,N_21657,N_21049);
or U22521 (N_22521,N_21514,N_21802);
xnor U22522 (N_22522,N_21488,N_21558);
nand U22523 (N_22523,N_21754,N_21423);
or U22524 (N_22524,N_21941,N_21614);
nand U22525 (N_22525,N_21607,N_21857);
nor U22526 (N_22526,N_21445,N_21915);
nand U22527 (N_22527,N_21020,N_21195);
nand U22528 (N_22528,N_21897,N_21847);
nor U22529 (N_22529,N_21216,N_21384);
nand U22530 (N_22530,N_21850,N_21058);
nand U22531 (N_22531,N_21107,N_21367);
or U22532 (N_22532,N_21502,N_21051);
nor U22533 (N_22533,N_21613,N_21389);
or U22534 (N_22534,N_21994,N_21237);
nand U22535 (N_22535,N_21196,N_21200);
xnor U22536 (N_22536,N_21217,N_21095);
xnor U22537 (N_22537,N_21406,N_21730);
and U22538 (N_22538,N_21504,N_21182);
nand U22539 (N_22539,N_21861,N_21780);
xnor U22540 (N_22540,N_21587,N_21282);
nor U22541 (N_22541,N_21009,N_21139);
and U22542 (N_22542,N_21457,N_21845);
or U22543 (N_22543,N_21786,N_21763);
or U22544 (N_22544,N_21058,N_21900);
and U22545 (N_22545,N_21410,N_21304);
and U22546 (N_22546,N_21993,N_21934);
nor U22547 (N_22547,N_21608,N_21359);
and U22548 (N_22548,N_21522,N_21556);
nor U22549 (N_22549,N_21305,N_21454);
xor U22550 (N_22550,N_21237,N_21078);
xor U22551 (N_22551,N_21654,N_21700);
nor U22552 (N_22552,N_21939,N_21110);
and U22553 (N_22553,N_21322,N_21889);
or U22554 (N_22554,N_21257,N_21794);
or U22555 (N_22555,N_21885,N_21060);
nor U22556 (N_22556,N_21001,N_21143);
nor U22557 (N_22557,N_21937,N_21033);
nor U22558 (N_22558,N_21955,N_21160);
nor U22559 (N_22559,N_21819,N_21737);
nand U22560 (N_22560,N_21467,N_21941);
xnor U22561 (N_22561,N_21628,N_21857);
xnor U22562 (N_22562,N_21125,N_21208);
xnor U22563 (N_22563,N_21061,N_21044);
or U22564 (N_22564,N_21469,N_21216);
nand U22565 (N_22565,N_21703,N_21752);
or U22566 (N_22566,N_21215,N_21038);
or U22567 (N_22567,N_21762,N_21011);
and U22568 (N_22568,N_21567,N_21848);
or U22569 (N_22569,N_21586,N_21910);
and U22570 (N_22570,N_21469,N_21948);
and U22571 (N_22571,N_21722,N_21063);
or U22572 (N_22572,N_21323,N_21445);
nor U22573 (N_22573,N_21211,N_21519);
or U22574 (N_22574,N_21656,N_21546);
xnor U22575 (N_22575,N_21402,N_21471);
or U22576 (N_22576,N_21852,N_21012);
or U22577 (N_22577,N_21178,N_21270);
nor U22578 (N_22578,N_21055,N_21297);
or U22579 (N_22579,N_21276,N_21536);
nor U22580 (N_22580,N_21578,N_21637);
nor U22581 (N_22581,N_21114,N_21976);
nand U22582 (N_22582,N_21145,N_21819);
nand U22583 (N_22583,N_21263,N_21347);
and U22584 (N_22584,N_21571,N_21438);
or U22585 (N_22585,N_21701,N_21113);
nor U22586 (N_22586,N_21781,N_21656);
xnor U22587 (N_22587,N_21754,N_21587);
and U22588 (N_22588,N_21140,N_21153);
or U22589 (N_22589,N_21304,N_21384);
nor U22590 (N_22590,N_21855,N_21950);
or U22591 (N_22591,N_21777,N_21512);
nor U22592 (N_22592,N_21715,N_21465);
or U22593 (N_22593,N_21960,N_21222);
or U22594 (N_22594,N_21525,N_21185);
nor U22595 (N_22595,N_21834,N_21464);
nand U22596 (N_22596,N_21959,N_21919);
nor U22597 (N_22597,N_21747,N_21217);
and U22598 (N_22598,N_21512,N_21423);
or U22599 (N_22599,N_21511,N_21095);
or U22600 (N_22600,N_21187,N_21816);
nor U22601 (N_22601,N_21298,N_21233);
or U22602 (N_22602,N_21673,N_21472);
or U22603 (N_22603,N_21721,N_21436);
nand U22604 (N_22604,N_21398,N_21596);
xnor U22605 (N_22605,N_21239,N_21344);
xor U22606 (N_22606,N_21830,N_21904);
xnor U22607 (N_22607,N_21694,N_21289);
nand U22608 (N_22608,N_21237,N_21931);
nand U22609 (N_22609,N_21959,N_21864);
and U22610 (N_22610,N_21733,N_21600);
and U22611 (N_22611,N_21419,N_21641);
nand U22612 (N_22612,N_21490,N_21562);
xor U22613 (N_22613,N_21754,N_21229);
nor U22614 (N_22614,N_21957,N_21789);
xor U22615 (N_22615,N_21135,N_21471);
nor U22616 (N_22616,N_21554,N_21872);
or U22617 (N_22617,N_21137,N_21773);
or U22618 (N_22618,N_21818,N_21292);
nand U22619 (N_22619,N_21273,N_21420);
xnor U22620 (N_22620,N_21419,N_21925);
nand U22621 (N_22621,N_21083,N_21612);
and U22622 (N_22622,N_21651,N_21560);
and U22623 (N_22623,N_21491,N_21950);
nor U22624 (N_22624,N_21554,N_21931);
and U22625 (N_22625,N_21611,N_21850);
nand U22626 (N_22626,N_21955,N_21355);
xnor U22627 (N_22627,N_21393,N_21685);
and U22628 (N_22628,N_21473,N_21144);
or U22629 (N_22629,N_21145,N_21212);
or U22630 (N_22630,N_21332,N_21815);
and U22631 (N_22631,N_21313,N_21229);
xor U22632 (N_22632,N_21618,N_21821);
xor U22633 (N_22633,N_21836,N_21457);
nand U22634 (N_22634,N_21769,N_21793);
xnor U22635 (N_22635,N_21737,N_21139);
or U22636 (N_22636,N_21055,N_21843);
nand U22637 (N_22637,N_21964,N_21703);
xor U22638 (N_22638,N_21268,N_21667);
xnor U22639 (N_22639,N_21880,N_21003);
nand U22640 (N_22640,N_21363,N_21507);
xnor U22641 (N_22641,N_21364,N_21826);
or U22642 (N_22642,N_21307,N_21591);
nand U22643 (N_22643,N_21285,N_21403);
nor U22644 (N_22644,N_21068,N_21388);
and U22645 (N_22645,N_21580,N_21304);
nor U22646 (N_22646,N_21474,N_21132);
and U22647 (N_22647,N_21342,N_21871);
and U22648 (N_22648,N_21915,N_21184);
or U22649 (N_22649,N_21528,N_21016);
nor U22650 (N_22650,N_21025,N_21113);
or U22651 (N_22651,N_21564,N_21244);
nand U22652 (N_22652,N_21321,N_21773);
and U22653 (N_22653,N_21188,N_21197);
or U22654 (N_22654,N_21614,N_21139);
nand U22655 (N_22655,N_21578,N_21849);
or U22656 (N_22656,N_21989,N_21456);
nand U22657 (N_22657,N_21453,N_21019);
or U22658 (N_22658,N_21559,N_21937);
or U22659 (N_22659,N_21566,N_21515);
xor U22660 (N_22660,N_21804,N_21869);
or U22661 (N_22661,N_21903,N_21479);
or U22662 (N_22662,N_21788,N_21055);
nand U22663 (N_22663,N_21447,N_21917);
nand U22664 (N_22664,N_21617,N_21389);
or U22665 (N_22665,N_21007,N_21650);
and U22666 (N_22666,N_21773,N_21394);
nor U22667 (N_22667,N_21872,N_21379);
xnor U22668 (N_22668,N_21563,N_21782);
xnor U22669 (N_22669,N_21893,N_21466);
and U22670 (N_22670,N_21323,N_21681);
xnor U22671 (N_22671,N_21013,N_21271);
and U22672 (N_22672,N_21986,N_21360);
nand U22673 (N_22673,N_21589,N_21652);
and U22674 (N_22674,N_21244,N_21182);
nand U22675 (N_22675,N_21057,N_21488);
nand U22676 (N_22676,N_21427,N_21989);
nor U22677 (N_22677,N_21839,N_21270);
nor U22678 (N_22678,N_21821,N_21159);
xnor U22679 (N_22679,N_21111,N_21059);
or U22680 (N_22680,N_21805,N_21014);
nand U22681 (N_22681,N_21528,N_21780);
nor U22682 (N_22682,N_21280,N_21578);
and U22683 (N_22683,N_21154,N_21109);
and U22684 (N_22684,N_21801,N_21526);
or U22685 (N_22685,N_21668,N_21184);
and U22686 (N_22686,N_21822,N_21751);
and U22687 (N_22687,N_21292,N_21791);
nor U22688 (N_22688,N_21255,N_21358);
and U22689 (N_22689,N_21376,N_21815);
nor U22690 (N_22690,N_21400,N_21348);
and U22691 (N_22691,N_21147,N_21534);
xnor U22692 (N_22692,N_21358,N_21791);
nor U22693 (N_22693,N_21091,N_21550);
xnor U22694 (N_22694,N_21910,N_21236);
nand U22695 (N_22695,N_21569,N_21743);
xnor U22696 (N_22696,N_21801,N_21316);
or U22697 (N_22697,N_21588,N_21206);
nand U22698 (N_22698,N_21187,N_21098);
xor U22699 (N_22699,N_21201,N_21045);
xor U22700 (N_22700,N_21522,N_21187);
xor U22701 (N_22701,N_21103,N_21762);
nor U22702 (N_22702,N_21338,N_21044);
nand U22703 (N_22703,N_21029,N_21189);
nand U22704 (N_22704,N_21424,N_21164);
xnor U22705 (N_22705,N_21603,N_21485);
and U22706 (N_22706,N_21497,N_21505);
nand U22707 (N_22707,N_21369,N_21179);
and U22708 (N_22708,N_21046,N_21637);
nor U22709 (N_22709,N_21308,N_21313);
or U22710 (N_22710,N_21150,N_21975);
nand U22711 (N_22711,N_21354,N_21168);
or U22712 (N_22712,N_21887,N_21721);
nand U22713 (N_22713,N_21155,N_21187);
nor U22714 (N_22714,N_21823,N_21301);
xor U22715 (N_22715,N_21748,N_21479);
nand U22716 (N_22716,N_21143,N_21204);
nand U22717 (N_22717,N_21727,N_21467);
xnor U22718 (N_22718,N_21382,N_21698);
or U22719 (N_22719,N_21463,N_21861);
or U22720 (N_22720,N_21797,N_21942);
or U22721 (N_22721,N_21186,N_21501);
nand U22722 (N_22722,N_21516,N_21531);
or U22723 (N_22723,N_21538,N_21912);
and U22724 (N_22724,N_21097,N_21565);
and U22725 (N_22725,N_21847,N_21948);
or U22726 (N_22726,N_21878,N_21308);
xor U22727 (N_22727,N_21893,N_21929);
and U22728 (N_22728,N_21825,N_21381);
nor U22729 (N_22729,N_21765,N_21888);
nand U22730 (N_22730,N_21769,N_21021);
xnor U22731 (N_22731,N_21156,N_21245);
nor U22732 (N_22732,N_21225,N_21059);
xnor U22733 (N_22733,N_21860,N_21014);
or U22734 (N_22734,N_21847,N_21024);
xor U22735 (N_22735,N_21704,N_21096);
nor U22736 (N_22736,N_21877,N_21071);
or U22737 (N_22737,N_21132,N_21956);
or U22738 (N_22738,N_21926,N_21333);
nor U22739 (N_22739,N_21987,N_21994);
xor U22740 (N_22740,N_21654,N_21186);
nand U22741 (N_22741,N_21071,N_21846);
nor U22742 (N_22742,N_21860,N_21495);
and U22743 (N_22743,N_21075,N_21079);
nor U22744 (N_22744,N_21748,N_21510);
and U22745 (N_22745,N_21847,N_21540);
xnor U22746 (N_22746,N_21822,N_21759);
and U22747 (N_22747,N_21508,N_21716);
nand U22748 (N_22748,N_21155,N_21282);
nand U22749 (N_22749,N_21482,N_21727);
or U22750 (N_22750,N_21989,N_21638);
or U22751 (N_22751,N_21107,N_21375);
nor U22752 (N_22752,N_21537,N_21312);
or U22753 (N_22753,N_21298,N_21108);
xor U22754 (N_22754,N_21365,N_21039);
nand U22755 (N_22755,N_21787,N_21010);
or U22756 (N_22756,N_21692,N_21571);
xnor U22757 (N_22757,N_21348,N_21362);
xor U22758 (N_22758,N_21261,N_21666);
xor U22759 (N_22759,N_21308,N_21873);
xnor U22760 (N_22760,N_21460,N_21932);
nor U22761 (N_22761,N_21261,N_21671);
or U22762 (N_22762,N_21281,N_21220);
and U22763 (N_22763,N_21737,N_21396);
nor U22764 (N_22764,N_21805,N_21799);
or U22765 (N_22765,N_21318,N_21315);
nand U22766 (N_22766,N_21773,N_21741);
or U22767 (N_22767,N_21355,N_21120);
or U22768 (N_22768,N_21344,N_21211);
nor U22769 (N_22769,N_21413,N_21168);
or U22770 (N_22770,N_21913,N_21580);
xnor U22771 (N_22771,N_21265,N_21727);
nor U22772 (N_22772,N_21161,N_21499);
and U22773 (N_22773,N_21539,N_21585);
and U22774 (N_22774,N_21459,N_21112);
nor U22775 (N_22775,N_21331,N_21154);
and U22776 (N_22776,N_21197,N_21515);
and U22777 (N_22777,N_21270,N_21899);
xor U22778 (N_22778,N_21469,N_21084);
nand U22779 (N_22779,N_21752,N_21631);
and U22780 (N_22780,N_21441,N_21403);
and U22781 (N_22781,N_21210,N_21245);
nand U22782 (N_22782,N_21020,N_21779);
nand U22783 (N_22783,N_21169,N_21786);
nand U22784 (N_22784,N_21170,N_21024);
or U22785 (N_22785,N_21639,N_21764);
nand U22786 (N_22786,N_21875,N_21644);
or U22787 (N_22787,N_21183,N_21572);
nor U22788 (N_22788,N_21794,N_21351);
xor U22789 (N_22789,N_21854,N_21479);
or U22790 (N_22790,N_21134,N_21252);
and U22791 (N_22791,N_21770,N_21624);
nand U22792 (N_22792,N_21750,N_21986);
and U22793 (N_22793,N_21076,N_21268);
nand U22794 (N_22794,N_21947,N_21824);
or U22795 (N_22795,N_21564,N_21917);
and U22796 (N_22796,N_21702,N_21521);
nor U22797 (N_22797,N_21847,N_21562);
nand U22798 (N_22798,N_21848,N_21908);
nand U22799 (N_22799,N_21894,N_21779);
nor U22800 (N_22800,N_21154,N_21351);
xnor U22801 (N_22801,N_21508,N_21371);
xor U22802 (N_22802,N_21733,N_21643);
xor U22803 (N_22803,N_21303,N_21156);
or U22804 (N_22804,N_21104,N_21049);
and U22805 (N_22805,N_21023,N_21776);
xor U22806 (N_22806,N_21350,N_21790);
nor U22807 (N_22807,N_21185,N_21409);
nand U22808 (N_22808,N_21576,N_21895);
xor U22809 (N_22809,N_21572,N_21874);
nand U22810 (N_22810,N_21405,N_21193);
nand U22811 (N_22811,N_21439,N_21129);
nand U22812 (N_22812,N_21867,N_21151);
nand U22813 (N_22813,N_21935,N_21879);
nor U22814 (N_22814,N_21609,N_21384);
and U22815 (N_22815,N_21746,N_21582);
nand U22816 (N_22816,N_21246,N_21176);
nor U22817 (N_22817,N_21206,N_21828);
xnor U22818 (N_22818,N_21771,N_21211);
nor U22819 (N_22819,N_21332,N_21506);
nor U22820 (N_22820,N_21895,N_21547);
xnor U22821 (N_22821,N_21974,N_21944);
and U22822 (N_22822,N_21345,N_21633);
nor U22823 (N_22823,N_21168,N_21332);
and U22824 (N_22824,N_21283,N_21479);
xor U22825 (N_22825,N_21098,N_21369);
and U22826 (N_22826,N_21392,N_21053);
or U22827 (N_22827,N_21085,N_21793);
and U22828 (N_22828,N_21736,N_21626);
xnor U22829 (N_22829,N_21735,N_21484);
xnor U22830 (N_22830,N_21650,N_21827);
xnor U22831 (N_22831,N_21563,N_21710);
nor U22832 (N_22832,N_21367,N_21835);
and U22833 (N_22833,N_21750,N_21663);
and U22834 (N_22834,N_21180,N_21692);
xor U22835 (N_22835,N_21318,N_21449);
xnor U22836 (N_22836,N_21121,N_21789);
and U22837 (N_22837,N_21320,N_21947);
or U22838 (N_22838,N_21923,N_21393);
xor U22839 (N_22839,N_21036,N_21400);
or U22840 (N_22840,N_21637,N_21210);
and U22841 (N_22841,N_21146,N_21873);
or U22842 (N_22842,N_21751,N_21108);
nor U22843 (N_22843,N_21058,N_21247);
nor U22844 (N_22844,N_21069,N_21407);
xor U22845 (N_22845,N_21833,N_21531);
xor U22846 (N_22846,N_21796,N_21322);
or U22847 (N_22847,N_21393,N_21367);
or U22848 (N_22848,N_21944,N_21529);
and U22849 (N_22849,N_21031,N_21744);
or U22850 (N_22850,N_21786,N_21447);
nand U22851 (N_22851,N_21671,N_21835);
or U22852 (N_22852,N_21516,N_21671);
nand U22853 (N_22853,N_21377,N_21524);
and U22854 (N_22854,N_21144,N_21725);
nand U22855 (N_22855,N_21433,N_21063);
and U22856 (N_22856,N_21332,N_21423);
and U22857 (N_22857,N_21517,N_21795);
nand U22858 (N_22858,N_21661,N_21967);
and U22859 (N_22859,N_21700,N_21659);
nand U22860 (N_22860,N_21796,N_21407);
or U22861 (N_22861,N_21096,N_21887);
xnor U22862 (N_22862,N_21313,N_21736);
nand U22863 (N_22863,N_21663,N_21817);
nand U22864 (N_22864,N_21619,N_21549);
and U22865 (N_22865,N_21332,N_21667);
and U22866 (N_22866,N_21693,N_21582);
nand U22867 (N_22867,N_21191,N_21809);
and U22868 (N_22868,N_21850,N_21196);
nand U22869 (N_22869,N_21851,N_21991);
nor U22870 (N_22870,N_21122,N_21340);
nor U22871 (N_22871,N_21726,N_21006);
xnor U22872 (N_22872,N_21481,N_21237);
nor U22873 (N_22873,N_21658,N_21230);
nor U22874 (N_22874,N_21863,N_21081);
nand U22875 (N_22875,N_21466,N_21205);
or U22876 (N_22876,N_21567,N_21434);
and U22877 (N_22877,N_21069,N_21479);
nand U22878 (N_22878,N_21364,N_21059);
and U22879 (N_22879,N_21528,N_21690);
nand U22880 (N_22880,N_21987,N_21981);
xor U22881 (N_22881,N_21521,N_21805);
nor U22882 (N_22882,N_21144,N_21254);
or U22883 (N_22883,N_21205,N_21967);
nor U22884 (N_22884,N_21636,N_21609);
or U22885 (N_22885,N_21739,N_21059);
xnor U22886 (N_22886,N_21706,N_21831);
or U22887 (N_22887,N_21741,N_21645);
nand U22888 (N_22888,N_21282,N_21512);
xor U22889 (N_22889,N_21171,N_21029);
and U22890 (N_22890,N_21154,N_21681);
nand U22891 (N_22891,N_21676,N_21110);
or U22892 (N_22892,N_21694,N_21542);
and U22893 (N_22893,N_21084,N_21654);
nand U22894 (N_22894,N_21298,N_21571);
nand U22895 (N_22895,N_21127,N_21631);
or U22896 (N_22896,N_21812,N_21877);
xor U22897 (N_22897,N_21764,N_21294);
or U22898 (N_22898,N_21441,N_21706);
nor U22899 (N_22899,N_21507,N_21247);
nand U22900 (N_22900,N_21532,N_21102);
nand U22901 (N_22901,N_21490,N_21939);
xnor U22902 (N_22902,N_21608,N_21456);
nor U22903 (N_22903,N_21770,N_21360);
nand U22904 (N_22904,N_21699,N_21282);
nand U22905 (N_22905,N_21795,N_21854);
or U22906 (N_22906,N_21063,N_21673);
xor U22907 (N_22907,N_21498,N_21341);
and U22908 (N_22908,N_21618,N_21381);
or U22909 (N_22909,N_21789,N_21052);
and U22910 (N_22910,N_21714,N_21879);
and U22911 (N_22911,N_21500,N_21704);
or U22912 (N_22912,N_21180,N_21005);
nor U22913 (N_22913,N_21740,N_21528);
or U22914 (N_22914,N_21006,N_21348);
or U22915 (N_22915,N_21247,N_21818);
and U22916 (N_22916,N_21128,N_21570);
and U22917 (N_22917,N_21212,N_21857);
or U22918 (N_22918,N_21001,N_21778);
or U22919 (N_22919,N_21811,N_21683);
and U22920 (N_22920,N_21195,N_21924);
xor U22921 (N_22921,N_21902,N_21686);
nor U22922 (N_22922,N_21969,N_21547);
xnor U22923 (N_22923,N_21834,N_21846);
xor U22924 (N_22924,N_21159,N_21459);
and U22925 (N_22925,N_21073,N_21686);
nor U22926 (N_22926,N_21434,N_21017);
nor U22927 (N_22927,N_21976,N_21290);
or U22928 (N_22928,N_21758,N_21173);
xnor U22929 (N_22929,N_21473,N_21903);
xor U22930 (N_22930,N_21669,N_21472);
nand U22931 (N_22931,N_21733,N_21818);
nor U22932 (N_22932,N_21525,N_21987);
nand U22933 (N_22933,N_21443,N_21726);
nand U22934 (N_22934,N_21254,N_21404);
nand U22935 (N_22935,N_21307,N_21360);
or U22936 (N_22936,N_21189,N_21578);
nor U22937 (N_22937,N_21591,N_21779);
xnor U22938 (N_22938,N_21594,N_21428);
nor U22939 (N_22939,N_21713,N_21144);
nor U22940 (N_22940,N_21879,N_21473);
nand U22941 (N_22941,N_21083,N_21486);
and U22942 (N_22942,N_21525,N_21271);
or U22943 (N_22943,N_21806,N_21375);
or U22944 (N_22944,N_21339,N_21635);
nand U22945 (N_22945,N_21346,N_21569);
nor U22946 (N_22946,N_21126,N_21317);
and U22947 (N_22947,N_21836,N_21887);
nand U22948 (N_22948,N_21064,N_21638);
xnor U22949 (N_22949,N_21006,N_21301);
nand U22950 (N_22950,N_21686,N_21599);
or U22951 (N_22951,N_21182,N_21755);
nand U22952 (N_22952,N_21103,N_21298);
and U22953 (N_22953,N_21659,N_21744);
nor U22954 (N_22954,N_21931,N_21484);
nor U22955 (N_22955,N_21756,N_21859);
and U22956 (N_22956,N_21906,N_21569);
xnor U22957 (N_22957,N_21418,N_21192);
nor U22958 (N_22958,N_21069,N_21730);
and U22959 (N_22959,N_21208,N_21357);
xnor U22960 (N_22960,N_21987,N_21486);
and U22961 (N_22961,N_21206,N_21567);
or U22962 (N_22962,N_21561,N_21009);
or U22963 (N_22963,N_21224,N_21476);
xor U22964 (N_22964,N_21011,N_21239);
nor U22965 (N_22965,N_21491,N_21640);
xor U22966 (N_22966,N_21914,N_21075);
xnor U22967 (N_22967,N_21485,N_21915);
or U22968 (N_22968,N_21765,N_21649);
and U22969 (N_22969,N_21229,N_21940);
nor U22970 (N_22970,N_21122,N_21667);
and U22971 (N_22971,N_21712,N_21620);
or U22972 (N_22972,N_21661,N_21994);
nand U22973 (N_22973,N_21111,N_21985);
and U22974 (N_22974,N_21165,N_21992);
xor U22975 (N_22975,N_21391,N_21643);
nand U22976 (N_22976,N_21013,N_21180);
xnor U22977 (N_22977,N_21622,N_21550);
or U22978 (N_22978,N_21160,N_21267);
nor U22979 (N_22979,N_21377,N_21749);
and U22980 (N_22980,N_21218,N_21930);
or U22981 (N_22981,N_21103,N_21125);
nor U22982 (N_22982,N_21480,N_21504);
nor U22983 (N_22983,N_21998,N_21754);
nand U22984 (N_22984,N_21959,N_21978);
nand U22985 (N_22985,N_21191,N_21044);
and U22986 (N_22986,N_21588,N_21339);
xor U22987 (N_22987,N_21930,N_21413);
xnor U22988 (N_22988,N_21530,N_21517);
or U22989 (N_22989,N_21203,N_21604);
xor U22990 (N_22990,N_21473,N_21755);
nor U22991 (N_22991,N_21506,N_21505);
nor U22992 (N_22992,N_21256,N_21639);
nor U22993 (N_22993,N_21260,N_21210);
xor U22994 (N_22994,N_21535,N_21818);
and U22995 (N_22995,N_21679,N_21304);
or U22996 (N_22996,N_21809,N_21268);
xor U22997 (N_22997,N_21706,N_21684);
or U22998 (N_22998,N_21713,N_21908);
or U22999 (N_22999,N_21682,N_21202);
nor U23000 (N_23000,N_22948,N_22135);
and U23001 (N_23001,N_22678,N_22764);
nor U23002 (N_23002,N_22860,N_22241);
xnor U23003 (N_23003,N_22535,N_22268);
and U23004 (N_23004,N_22592,N_22902);
or U23005 (N_23005,N_22240,N_22757);
or U23006 (N_23006,N_22547,N_22417);
nor U23007 (N_23007,N_22248,N_22273);
nor U23008 (N_23008,N_22529,N_22447);
nand U23009 (N_23009,N_22053,N_22664);
xnor U23010 (N_23010,N_22340,N_22020);
or U23011 (N_23011,N_22416,N_22243);
xnor U23012 (N_23012,N_22088,N_22175);
nand U23013 (N_23013,N_22207,N_22393);
xor U23014 (N_23014,N_22496,N_22706);
and U23015 (N_23015,N_22328,N_22477);
nor U23016 (N_23016,N_22455,N_22443);
nor U23017 (N_23017,N_22519,N_22392);
xor U23018 (N_23018,N_22675,N_22472);
or U23019 (N_23019,N_22450,N_22296);
or U23020 (N_23020,N_22224,N_22137);
and U23021 (N_23021,N_22863,N_22532);
or U23022 (N_23022,N_22636,N_22069);
nor U23023 (N_23023,N_22728,N_22196);
nor U23024 (N_23024,N_22335,N_22935);
nor U23025 (N_23025,N_22537,N_22278);
xnor U23026 (N_23026,N_22688,N_22559);
nand U23027 (N_23027,N_22884,N_22620);
or U23028 (N_23028,N_22879,N_22584);
and U23029 (N_23029,N_22050,N_22075);
or U23030 (N_23030,N_22616,N_22955);
and U23031 (N_23031,N_22815,N_22512);
nand U23032 (N_23032,N_22352,N_22025);
xor U23033 (N_23033,N_22520,N_22787);
and U23034 (N_23034,N_22601,N_22263);
xnor U23035 (N_23035,N_22441,N_22101);
nand U23036 (N_23036,N_22148,N_22431);
xnor U23037 (N_23037,N_22065,N_22323);
nand U23038 (N_23038,N_22700,N_22799);
xnor U23039 (N_23039,N_22722,N_22538);
nor U23040 (N_23040,N_22324,N_22821);
nor U23041 (N_23041,N_22168,N_22357);
and U23042 (N_23042,N_22848,N_22056);
nand U23043 (N_23043,N_22531,N_22912);
and U23044 (N_23044,N_22483,N_22172);
xor U23045 (N_23045,N_22910,N_22800);
or U23046 (N_23046,N_22375,N_22112);
nand U23047 (N_23047,N_22167,N_22811);
or U23048 (N_23048,N_22680,N_22322);
xnor U23049 (N_23049,N_22140,N_22694);
and U23050 (N_23050,N_22151,N_22609);
or U23051 (N_23051,N_22561,N_22841);
and U23052 (N_23052,N_22981,N_22638);
nand U23053 (N_23053,N_22824,N_22959);
or U23054 (N_23054,N_22937,N_22313);
or U23055 (N_23055,N_22369,N_22656);
nand U23056 (N_23056,N_22994,N_22999);
xor U23057 (N_23057,N_22578,N_22777);
xnor U23058 (N_23058,N_22671,N_22725);
xor U23059 (N_23059,N_22621,N_22349);
and U23060 (N_23060,N_22696,N_22499);
nand U23061 (N_23061,N_22522,N_22767);
or U23062 (N_23062,N_22100,N_22061);
nor U23063 (N_23063,N_22095,N_22729);
and U23064 (N_23064,N_22844,N_22864);
nand U23065 (N_23065,N_22640,N_22002);
xor U23066 (N_23066,N_22201,N_22708);
and U23067 (N_23067,N_22752,N_22735);
nor U23068 (N_23068,N_22284,N_22422);
xor U23069 (N_23069,N_22571,N_22145);
and U23070 (N_23070,N_22200,N_22896);
nand U23071 (N_23071,N_22992,N_22227);
nand U23072 (N_23072,N_22486,N_22070);
xor U23073 (N_23073,N_22454,N_22551);
nand U23074 (N_23074,N_22698,N_22338);
xnor U23075 (N_23075,N_22469,N_22911);
or U23076 (N_23076,N_22288,N_22781);
nor U23077 (N_23077,N_22693,N_22627);
and U23078 (N_23078,N_22615,N_22297);
or U23079 (N_23079,N_22083,N_22921);
or U23080 (N_23080,N_22104,N_22952);
nor U23081 (N_23081,N_22134,N_22331);
nor U23082 (N_23082,N_22947,N_22042);
xor U23083 (N_23083,N_22479,N_22176);
or U23084 (N_23084,N_22403,N_22822);
nor U23085 (N_23085,N_22110,N_22527);
and U23086 (N_23086,N_22978,N_22272);
nand U23087 (N_23087,N_22464,N_22173);
or U23088 (N_23088,N_22114,N_22541);
xnor U23089 (N_23089,N_22673,N_22548);
nor U23090 (N_23090,N_22440,N_22304);
nor U23091 (N_23091,N_22745,N_22690);
or U23092 (N_23092,N_22966,N_22583);
nand U23093 (N_23093,N_22186,N_22309);
or U23094 (N_23094,N_22399,N_22652);
nand U23095 (N_23095,N_22368,N_22345);
nor U23096 (N_23096,N_22610,N_22869);
nand U23097 (N_23097,N_22497,N_22475);
nor U23098 (N_23098,N_22995,N_22596);
nand U23099 (N_23099,N_22813,N_22790);
xnor U23100 (N_23100,N_22556,N_22149);
or U23101 (N_23101,N_22852,N_22803);
and U23102 (N_23102,N_22925,N_22669);
and U23103 (N_23103,N_22190,N_22147);
and U23104 (N_23104,N_22348,N_22819);
nand U23105 (N_23105,N_22015,N_22302);
xor U23106 (N_23106,N_22810,N_22940);
xnor U23107 (N_23107,N_22846,N_22883);
and U23108 (N_23108,N_22740,N_22458);
and U23109 (N_23109,N_22318,N_22234);
nor U23110 (N_23110,N_22866,N_22446);
nor U23111 (N_23111,N_22985,N_22677);
nand U23112 (N_23112,N_22377,N_22518);
nor U23113 (N_23113,N_22398,N_22188);
xnor U23114 (N_23114,N_22644,N_22271);
and U23115 (N_23115,N_22950,N_22954);
and U23116 (N_23116,N_22320,N_22132);
xor U23117 (N_23117,N_22526,N_22027);
and U23118 (N_23118,N_22256,N_22709);
nand U23119 (N_23119,N_22506,N_22951);
nand U23120 (N_23120,N_22975,N_22424);
and U23121 (N_23121,N_22834,N_22292);
and U23122 (N_23122,N_22639,N_22407);
and U23123 (N_23123,N_22624,N_22946);
nand U23124 (N_23124,N_22276,N_22521);
nor U23125 (N_23125,N_22942,N_22908);
and U23126 (N_23126,N_22542,N_22774);
and U23127 (N_23127,N_22130,N_22931);
nand U23128 (N_23128,N_22353,N_22468);
xor U23129 (N_23129,N_22182,N_22222);
or U23130 (N_23130,N_22979,N_22895);
xnor U23131 (N_23131,N_22901,N_22588);
or U23132 (N_23132,N_22713,N_22419);
nor U23133 (N_23133,N_22058,N_22829);
or U23134 (N_23134,N_22124,N_22524);
or U23135 (N_23135,N_22603,N_22772);
or U23136 (N_23136,N_22004,N_22258);
nor U23137 (N_23137,N_22120,N_22433);
nand U23138 (N_23138,N_22067,N_22612);
xnor U23139 (N_23139,N_22456,N_22528);
nand U23140 (N_23140,N_22406,N_22637);
xnor U23141 (N_23141,N_22213,N_22789);
or U23142 (N_23142,N_22501,N_22193);
nand U23143 (N_23143,N_22043,N_22899);
and U23144 (N_23144,N_22650,N_22174);
and U23145 (N_23145,N_22969,N_22773);
or U23146 (N_23146,N_22593,N_22429);
or U23147 (N_23147,N_22641,N_22461);
and U23148 (N_23148,N_22044,N_22298);
nor U23149 (N_23149,N_22041,N_22106);
and U23150 (N_23150,N_22129,N_22093);
nand U23151 (N_23151,N_22651,N_22888);
or U23152 (N_23152,N_22554,N_22462);
and U23153 (N_23153,N_22388,N_22972);
xnor U23154 (N_23154,N_22923,N_22037);
nand U23155 (N_23155,N_22039,N_22536);
xnor U23156 (N_23156,N_22974,N_22870);
and U23157 (N_23157,N_22460,N_22223);
or U23158 (N_23158,N_22607,N_22802);
and U23159 (N_23159,N_22160,N_22481);
nand U23160 (N_23160,N_22293,N_22687);
nand U23161 (N_23161,N_22126,N_22714);
xor U23162 (N_23162,N_22394,N_22395);
or U23163 (N_23163,N_22289,N_22927);
xor U23164 (N_23164,N_22382,N_22307);
nor U23165 (N_23165,N_22915,N_22146);
nor U23166 (N_23166,N_22847,N_22859);
and U23167 (N_23167,N_22500,N_22003);
nor U23168 (N_23168,N_22991,N_22558);
nand U23169 (N_23169,N_22262,N_22152);
nand U23170 (N_23170,N_22105,N_22676);
nor U23171 (N_23171,N_22574,N_22759);
nand U23172 (N_23172,N_22643,N_22435);
or U23173 (N_23173,N_22316,N_22026);
xor U23174 (N_23174,N_22202,N_22198);
xor U23175 (N_23175,N_22311,N_22195);
or U23176 (N_23176,N_22898,N_22466);
and U23177 (N_23177,N_22618,N_22473);
nor U23178 (N_23178,N_22366,N_22376);
or U23179 (N_23179,N_22763,N_22438);
and U23180 (N_23180,N_22566,N_22900);
nor U23181 (N_23181,N_22683,N_22448);
and U23182 (N_23182,N_22890,N_22667);
xor U23183 (N_23183,N_22237,N_22494);
and U23184 (N_23184,N_22049,N_22098);
and U23185 (N_23185,N_22963,N_22017);
nand U23186 (N_23186,N_22699,N_22875);
xnor U23187 (N_23187,N_22502,N_22582);
or U23188 (N_23188,N_22107,N_22205);
nor U23189 (N_23189,N_22540,N_22389);
and U23190 (N_23190,N_22054,N_22250);
nand U23191 (N_23191,N_22219,N_22747);
nor U23192 (N_23192,N_22600,N_22555);
nor U23193 (N_23193,N_22177,N_22823);
xor U23194 (N_23194,N_22836,N_22893);
nand U23195 (N_23195,N_22346,N_22267);
nor U23196 (N_23196,N_22515,N_22046);
nor U23197 (N_23197,N_22034,N_22367);
and U23198 (N_23198,N_22679,N_22619);
xor U23199 (N_23199,N_22136,N_22756);
xor U23200 (N_23200,N_22956,N_22031);
and U23201 (N_23201,N_22573,N_22997);
xnor U23202 (N_23202,N_22712,N_22692);
xor U23203 (N_23203,N_22760,N_22445);
and U23204 (N_23204,N_22336,N_22442);
and U23205 (N_23205,N_22845,N_22854);
nor U23206 (N_23206,N_22837,N_22185);
and U23207 (N_23207,N_22478,N_22791);
or U23208 (N_23208,N_22741,N_22206);
nand U23209 (N_23209,N_22192,N_22986);
and U23210 (N_23210,N_22505,N_22119);
nor U23211 (N_23211,N_22337,N_22021);
and U23212 (N_23212,N_22342,N_22255);
and U23213 (N_23213,N_22743,N_22907);
nand U23214 (N_23214,N_22371,N_22567);
nand U23215 (N_23215,N_22586,N_22560);
and U23216 (N_23216,N_22798,N_22507);
nand U23217 (N_23217,N_22611,N_22572);
and U23218 (N_23218,N_22654,N_22855);
and U23219 (N_23219,N_22066,N_22405);
or U23220 (N_23220,N_22047,N_22727);
and U23221 (N_23221,N_22629,N_22029);
nand U23222 (N_23222,N_22154,N_22139);
nor U23223 (N_23223,N_22370,N_22666);
nand U23224 (N_23224,N_22749,N_22511);
nand U23225 (N_23225,N_22242,N_22339);
nor U23226 (N_23226,N_22958,N_22885);
or U23227 (N_23227,N_22363,N_22606);
and U23228 (N_23228,N_22783,N_22330);
and U23229 (N_23229,N_22674,N_22019);
or U23230 (N_23230,N_22504,N_22295);
xor U23231 (N_23231,N_22544,N_22608);
or U23232 (N_23232,N_22327,N_22045);
nor U23233 (N_23233,N_22482,N_22878);
nand U23234 (N_23234,N_22932,N_22938);
nand U23235 (N_23235,N_22082,N_22816);
xor U23236 (N_23236,N_22232,N_22568);
xnor U23237 (N_23237,N_22007,N_22962);
nor U23238 (N_23238,N_22736,N_22385);
and U23239 (N_23239,N_22489,N_22916);
nand U23240 (N_23240,N_22917,N_22287);
and U23241 (N_23241,N_22751,N_22081);
nor U23242 (N_23242,N_22808,N_22886);
xnor U23243 (N_23243,N_22432,N_22633);
or U23244 (N_23244,N_22270,N_22539);
nor U23245 (N_23245,N_22861,N_22071);
nor U23246 (N_23246,N_22453,N_22077);
nor U23247 (N_23247,N_22068,N_22707);
or U23248 (N_23248,N_22239,N_22372);
and U23249 (N_23249,N_22150,N_22018);
nor U23250 (N_23250,N_22035,N_22228);
nand U23251 (N_23251,N_22118,N_22929);
nand U23252 (N_23252,N_22503,N_22575);
nor U23253 (N_23253,N_22839,N_22257);
or U23254 (N_23254,N_22514,N_22159);
nor U23255 (N_23255,N_22761,N_22853);
and U23256 (N_23256,N_22299,N_22812);
xnor U23257 (N_23257,N_22161,N_22973);
xnor U23258 (N_23258,N_22244,N_22856);
or U23259 (N_23259,N_22079,N_22589);
or U23260 (N_23260,N_22006,N_22795);
nor U23261 (N_23261,N_22825,N_22216);
nor U23262 (N_23262,N_22701,N_22344);
and U23263 (N_23263,N_22252,N_22413);
or U23264 (N_23264,N_22133,N_22628);
nand U23265 (N_23265,N_22748,N_22960);
and U23266 (N_23266,N_22657,N_22212);
xor U23267 (N_23267,N_22880,N_22164);
nor U23268 (N_23268,N_22581,N_22378);
xnor U23269 (N_23269,N_22534,N_22076);
or U23270 (N_23270,N_22251,N_22265);
xor U23271 (N_23271,N_22961,N_22982);
or U23272 (N_23272,N_22365,N_22163);
or U23273 (N_23273,N_22922,N_22421);
or U23274 (N_23274,N_22968,N_22204);
or U23275 (N_23275,N_22980,N_22341);
xor U23276 (N_23276,N_22488,N_22742);
xnor U23277 (N_23277,N_22439,N_22509);
nand U23278 (N_23278,N_22919,N_22495);
nor U23279 (N_23279,N_22734,N_22487);
nor U23280 (N_23280,N_22631,N_22569);
and U23281 (N_23281,N_22402,N_22380);
or U23282 (N_23282,N_22724,N_22356);
or U23283 (N_23283,N_22412,N_22142);
nor U23284 (N_23284,N_22051,N_22930);
or U23285 (N_23285,N_22842,N_22702);
nand U23286 (N_23286,N_22807,N_22218);
and U23287 (N_23287,N_22545,N_22310);
nor U23288 (N_23288,N_22233,N_22953);
or U23289 (N_23289,N_22964,N_22939);
nand U23290 (N_23290,N_22806,N_22943);
nor U23291 (N_23291,N_22788,N_22993);
nand U23292 (N_23292,N_22024,N_22291);
or U23293 (N_23293,N_22715,N_22203);
or U23294 (N_23294,N_22474,N_22274);
xnor U23295 (N_23295,N_22321,N_22125);
nor U23296 (N_23296,N_22220,N_22074);
or U23297 (N_23297,N_22697,N_22165);
nor U23298 (N_23298,N_22226,N_22040);
or U23299 (N_23299,N_22197,N_22622);
nor U23300 (N_23300,N_22379,N_22723);
and U23301 (N_23301,N_22123,N_22452);
nor U23302 (N_23302,N_22894,N_22072);
nand U23303 (N_23303,N_22648,N_22794);
xnor U23304 (N_23304,N_22704,N_22786);
nand U23305 (N_23305,N_22092,N_22306);
nand U23306 (N_23306,N_22796,N_22977);
xnor U23307 (N_23307,N_22094,N_22036);
nand U23308 (N_23308,N_22209,N_22384);
or U23309 (N_23309,N_22818,N_22418);
xor U23310 (N_23310,N_22513,N_22334);
or U23311 (N_23311,N_22891,N_22383);
nand U23312 (N_23312,N_22828,N_22108);
xnor U23313 (N_23313,N_22765,N_22457);
and U23314 (N_23314,N_22102,N_22766);
and U23315 (N_23315,N_22523,N_22549);
nand U23316 (N_23316,N_22934,N_22158);
nor U23317 (N_23317,N_22936,N_22604);
nor U23318 (N_23318,N_22871,N_22892);
nand U23319 (N_23319,N_22199,N_22180);
nand U23320 (N_23320,N_22281,N_22113);
and U23321 (N_23321,N_22266,N_22630);
xor U23322 (N_23322,N_22645,N_22290);
nand U23323 (N_23323,N_22685,N_22703);
and U23324 (N_23324,N_22231,N_22033);
nor U23325 (N_23325,N_22762,N_22913);
nor U23326 (N_23326,N_22022,N_22359);
nor U23327 (N_23327,N_22711,N_22672);
and U23328 (N_23328,N_22738,N_22613);
nand U23329 (N_23329,N_22183,N_22705);
and U23330 (N_23330,N_22401,N_22391);
nand U23331 (N_23331,N_22928,N_22470);
nand U23332 (N_23332,N_22013,N_22784);
and U23333 (N_23333,N_22510,N_22873);
xor U23334 (N_23334,N_22990,N_22373);
xor U23335 (N_23335,N_22691,N_22351);
xor U23336 (N_23336,N_22062,N_22286);
and U23337 (N_23337,N_22400,N_22909);
nand U23338 (N_23338,N_22642,N_22492);
nand U23339 (N_23339,N_22277,N_22625);
nand U23340 (N_23340,N_22597,N_22089);
or U23341 (N_23341,N_22109,N_22484);
nand U23342 (N_23342,N_22670,N_22996);
and U23343 (N_23343,N_22355,N_22755);
or U23344 (N_23344,N_22782,N_22647);
xnor U23345 (N_23345,N_22830,N_22721);
nand U23346 (N_23346,N_22655,N_22000);
nor U23347 (N_23347,N_22360,N_22116);
and U23348 (N_23348,N_22849,N_22169);
xor U23349 (N_23349,N_22976,N_22087);
nand U23350 (N_23350,N_22319,N_22598);
nor U23351 (N_23351,N_22591,N_22579);
nand U23352 (N_23352,N_22801,N_22662);
and U23353 (N_23353,N_22533,N_22970);
nor U23354 (N_23354,N_22785,N_22594);
xnor U23355 (N_23355,N_22386,N_22471);
and U23356 (N_23356,N_22858,N_22754);
or U23357 (N_23357,N_22967,N_22153);
nor U23358 (N_23358,N_22737,N_22236);
xor U23359 (N_23359,N_22122,N_22280);
and U23360 (N_23360,N_22476,N_22155);
and U23361 (N_23361,N_22595,N_22221);
nand U23362 (N_23362,N_22817,N_22364);
nand U23363 (N_23363,N_22868,N_22649);
xnor U23364 (N_23364,N_22557,N_22746);
or U23365 (N_23365,N_22301,N_22465);
nor U23366 (N_23366,N_22410,N_22874);
nand U23367 (N_23367,N_22001,N_22732);
xor U23368 (N_23368,N_22792,N_22838);
or U23369 (N_23369,N_22390,N_22904);
nor U23370 (N_23370,N_22260,N_22623);
nor U23371 (N_23371,N_22553,N_22332);
xor U23372 (N_23372,N_22127,N_22944);
nand U23373 (N_23373,N_22329,N_22420);
nand U23374 (N_23374,N_22686,N_22753);
xor U23375 (N_23375,N_22181,N_22779);
and U23376 (N_23376,N_22872,N_22739);
nor U23377 (N_23377,N_22189,N_22682);
or U23378 (N_23378,N_22905,N_22317);
or U23379 (N_23379,N_22771,N_22121);
xor U23380 (N_23380,N_22211,N_22315);
nor U23381 (N_23381,N_22987,N_22245);
or U23382 (N_23382,N_22249,N_22217);
xor U23383 (N_23383,N_22264,N_22343);
and U23384 (N_23384,N_22178,N_22411);
nor U23385 (N_23385,N_22646,N_22354);
and U23386 (N_23386,N_22776,N_22063);
nand U23387 (N_23387,N_22850,N_22867);
nor U23388 (N_23388,N_22726,N_22451);
xnor U23389 (N_23389,N_22490,N_22425);
and U23390 (N_23390,N_22924,N_22926);
and U23391 (N_23391,N_22187,N_22428);
or U23392 (N_23392,N_22530,N_22414);
or U23393 (N_23393,N_22660,N_22409);
xor U23394 (N_23394,N_22617,N_22009);
or U23395 (N_23395,N_22971,N_22312);
xor U23396 (N_23396,N_22793,N_22259);
nor U23397 (N_23397,N_22358,N_22308);
xor U23398 (N_23398,N_22933,N_22170);
and U23399 (N_23399,N_22897,N_22750);
and U23400 (N_23400,N_22920,N_22733);
or U23401 (N_23401,N_22073,N_22498);
nand U23402 (N_23402,N_22246,N_22294);
xor U23403 (N_23403,N_22731,N_22957);
or U23404 (N_23404,N_22508,N_22230);
xor U23405 (N_23405,N_22626,N_22326);
and U23406 (N_23406,N_22179,N_22546);
xnor U23407 (N_23407,N_22570,N_22350);
nand U23408 (N_23408,N_22303,N_22023);
nor U23409 (N_23409,N_22718,N_22166);
nand U23410 (N_23410,N_22064,N_22614);
nand U23411 (N_23411,N_22084,N_22491);
xnor U23412 (N_23412,N_22577,N_22668);
or U23413 (N_23413,N_22827,N_22275);
or U23414 (N_23414,N_22998,N_22983);
or U23415 (N_23415,N_22843,N_22404);
and U23416 (N_23416,N_22214,N_22215);
and U23417 (N_23417,N_22730,N_22208);
and U23418 (N_23418,N_22325,N_22634);
and U23419 (N_23419,N_22171,N_22988);
nor U23420 (N_23420,N_22184,N_22397);
nand U23421 (N_23421,N_22374,N_22032);
or U23422 (N_23422,N_22914,N_22467);
nor U23423 (N_23423,N_22157,N_22744);
and U23424 (N_23424,N_22805,N_22225);
and U23425 (N_23425,N_22918,N_22543);
or U23426 (N_23426,N_22085,N_22525);
nor U23427 (N_23427,N_22989,N_22261);
and U23428 (N_23428,N_22396,N_22096);
xnor U23429 (N_23429,N_22661,N_22632);
or U23430 (N_23430,N_22059,N_22057);
and U23431 (N_23431,N_22768,N_22117);
or U23432 (N_23432,N_22434,N_22048);
or U23433 (N_23433,N_22717,N_22635);
nand U23434 (N_23434,N_22493,N_22889);
xnor U23435 (N_23435,N_22882,N_22887);
or U23436 (N_23436,N_22949,N_22014);
xor U23437 (N_23437,N_22832,N_22463);
nor U23438 (N_23438,N_22078,N_22695);
nor U23439 (N_23439,N_22103,N_22945);
nand U23440 (N_23440,N_22086,N_22162);
nor U23441 (N_23441,N_22903,N_22758);
xnor U23442 (N_23442,N_22144,N_22052);
and U23443 (N_23443,N_22143,N_22194);
xor U23444 (N_23444,N_22444,N_22279);
and U23445 (N_23445,N_22247,N_22480);
xor U23446 (N_23446,N_22285,N_22599);
or U23447 (N_23447,N_22235,N_22851);
nand U23448 (N_23448,N_22585,N_22877);
or U23449 (N_23449,N_22770,N_22865);
nor U23450 (N_23450,N_22826,N_22115);
nand U23451 (N_23451,N_22333,N_22381);
nor U23452 (N_23452,N_22128,N_22253);
nor U23453 (N_23453,N_22016,N_22833);
or U23454 (N_23454,N_22011,N_22430);
nor U23455 (N_23455,N_22716,N_22881);
and U23456 (N_23456,N_22387,N_22038);
nand U23457 (N_23457,N_22191,N_22459);
nand U23458 (N_23458,N_22131,N_22965);
nand U23459 (N_23459,N_22562,N_22552);
xor U23460 (N_23460,N_22550,N_22080);
nand U23461 (N_23461,N_22769,N_22138);
nand U23462 (N_23462,N_22111,N_22254);
nand U23463 (N_23463,N_22099,N_22269);
nor U23464 (N_23464,N_22775,N_22097);
xor U23465 (N_23465,N_22415,N_22005);
and U23466 (N_23466,N_22587,N_22576);
or U23467 (N_23467,N_22426,N_22229);
nor U23468 (N_23468,N_22408,N_22485);
nor U23469 (N_23469,N_22564,N_22804);
nand U23470 (N_23470,N_22156,N_22030);
nor U23471 (N_23471,N_22659,N_22090);
and U23472 (N_23472,N_22862,N_22427);
and U23473 (N_23473,N_22362,N_22300);
or U23474 (N_23474,N_22437,N_22565);
xor U23475 (N_23475,N_22602,N_22580);
or U23476 (N_23476,N_22941,N_22684);
nand U23477 (N_23477,N_22141,N_22517);
xor U23478 (N_23478,N_22347,N_22361);
nor U23479 (N_23479,N_22835,N_22857);
nand U23480 (N_23480,N_22010,N_22663);
nor U23481 (N_23481,N_22665,N_22436);
and U23482 (N_23482,N_22563,N_22778);
nand U23483 (N_23483,N_22605,N_22658);
or U23484 (N_23484,N_22720,N_22423);
xnor U23485 (N_23485,N_22814,N_22305);
xor U23486 (N_23486,N_22055,N_22210);
or U23487 (N_23487,N_22028,N_22653);
and U23488 (N_23488,N_22516,N_22710);
xnor U23489 (N_23489,N_22283,N_22282);
nor U23490 (N_23490,N_22840,N_22906);
nor U23491 (N_23491,N_22689,N_22797);
nand U23492 (N_23492,N_22809,N_22012);
xor U23493 (N_23493,N_22780,N_22449);
nand U23494 (N_23494,N_22820,N_22719);
xor U23495 (N_23495,N_22876,N_22590);
xor U23496 (N_23496,N_22314,N_22238);
xor U23497 (N_23497,N_22091,N_22008);
nand U23498 (N_23498,N_22060,N_22831);
nand U23499 (N_23499,N_22681,N_22984);
and U23500 (N_23500,N_22441,N_22764);
nand U23501 (N_23501,N_22248,N_22953);
nand U23502 (N_23502,N_22034,N_22515);
nor U23503 (N_23503,N_22393,N_22924);
nor U23504 (N_23504,N_22860,N_22944);
or U23505 (N_23505,N_22023,N_22489);
nand U23506 (N_23506,N_22630,N_22645);
or U23507 (N_23507,N_22633,N_22329);
nand U23508 (N_23508,N_22587,N_22003);
xor U23509 (N_23509,N_22058,N_22543);
nand U23510 (N_23510,N_22156,N_22580);
and U23511 (N_23511,N_22774,N_22607);
nor U23512 (N_23512,N_22292,N_22527);
or U23513 (N_23513,N_22964,N_22994);
xnor U23514 (N_23514,N_22258,N_22625);
or U23515 (N_23515,N_22303,N_22687);
or U23516 (N_23516,N_22733,N_22224);
and U23517 (N_23517,N_22725,N_22308);
and U23518 (N_23518,N_22535,N_22294);
nand U23519 (N_23519,N_22301,N_22080);
or U23520 (N_23520,N_22803,N_22624);
nand U23521 (N_23521,N_22909,N_22851);
xor U23522 (N_23522,N_22832,N_22599);
nor U23523 (N_23523,N_22575,N_22070);
and U23524 (N_23524,N_22183,N_22846);
nand U23525 (N_23525,N_22946,N_22426);
xor U23526 (N_23526,N_22523,N_22952);
nand U23527 (N_23527,N_22233,N_22493);
and U23528 (N_23528,N_22417,N_22695);
xnor U23529 (N_23529,N_22950,N_22009);
xor U23530 (N_23530,N_22844,N_22723);
nor U23531 (N_23531,N_22077,N_22957);
nor U23532 (N_23532,N_22757,N_22207);
or U23533 (N_23533,N_22317,N_22164);
or U23534 (N_23534,N_22351,N_22125);
xor U23535 (N_23535,N_22936,N_22162);
nor U23536 (N_23536,N_22213,N_22624);
nand U23537 (N_23537,N_22958,N_22303);
nor U23538 (N_23538,N_22786,N_22858);
or U23539 (N_23539,N_22901,N_22832);
nand U23540 (N_23540,N_22288,N_22148);
or U23541 (N_23541,N_22625,N_22731);
xnor U23542 (N_23542,N_22248,N_22478);
nand U23543 (N_23543,N_22797,N_22075);
or U23544 (N_23544,N_22271,N_22740);
nand U23545 (N_23545,N_22993,N_22072);
xor U23546 (N_23546,N_22282,N_22863);
nor U23547 (N_23547,N_22060,N_22801);
nand U23548 (N_23548,N_22559,N_22642);
nand U23549 (N_23549,N_22871,N_22115);
xor U23550 (N_23550,N_22856,N_22798);
or U23551 (N_23551,N_22984,N_22678);
or U23552 (N_23552,N_22485,N_22971);
xor U23553 (N_23553,N_22586,N_22671);
and U23554 (N_23554,N_22734,N_22346);
xor U23555 (N_23555,N_22501,N_22024);
nand U23556 (N_23556,N_22674,N_22882);
nor U23557 (N_23557,N_22322,N_22624);
nor U23558 (N_23558,N_22898,N_22463);
and U23559 (N_23559,N_22421,N_22364);
and U23560 (N_23560,N_22518,N_22674);
nand U23561 (N_23561,N_22429,N_22813);
and U23562 (N_23562,N_22547,N_22589);
nand U23563 (N_23563,N_22289,N_22850);
xnor U23564 (N_23564,N_22681,N_22258);
xor U23565 (N_23565,N_22122,N_22463);
xor U23566 (N_23566,N_22291,N_22111);
nand U23567 (N_23567,N_22139,N_22838);
nor U23568 (N_23568,N_22067,N_22943);
nand U23569 (N_23569,N_22778,N_22992);
nor U23570 (N_23570,N_22315,N_22923);
nand U23571 (N_23571,N_22559,N_22305);
xor U23572 (N_23572,N_22506,N_22821);
and U23573 (N_23573,N_22352,N_22441);
nor U23574 (N_23574,N_22113,N_22920);
or U23575 (N_23575,N_22738,N_22222);
xor U23576 (N_23576,N_22122,N_22903);
nand U23577 (N_23577,N_22577,N_22782);
xnor U23578 (N_23578,N_22052,N_22562);
xor U23579 (N_23579,N_22159,N_22343);
nor U23580 (N_23580,N_22390,N_22046);
nand U23581 (N_23581,N_22114,N_22291);
xnor U23582 (N_23582,N_22707,N_22470);
xor U23583 (N_23583,N_22086,N_22391);
or U23584 (N_23584,N_22535,N_22266);
xor U23585 (N_23585,N_22695,N_22014);
nand U23586 (N_23586,N_22113,N_22060);
nand U23587 (N_23587,N_22563,N_22819);
xor U23588 (N_23588,N_22092,N_22257);
nand U23589 (N_23589,N_22001,N_22338);
or U23590 (N_23590,N_22151,N_22473);
nand U23591 (N_23591,N_22894,N_22524);
xnor U23592 (N_23592,N_22402,N_22840);
and U23593 (N_23593,N_22096,N_22285);
or U23594 (N_23594,N_22199,N_22889);
xor U23595 (N_23595,N_22816,N_22174);
nand U23596 (N_23596,N_22781,N_22798);
nand U23597 (N_23597,N_22349,N_22963);
xor U23598 (N_23598,N_22177,N_22022);
xor U23599 (N_23599,N_22939,N_22830);
nand U23600 (N_23600,N_22961,N_22551);
nand U23601 (N_23601,N_22617,N_22065);
nor U23602 (N_23602,N_22658,N_22645);
nand U23603 (N_23603,N_22770,N_22723);
and U23604 (N_23604,N_22003,N_22529);
or U23605 (N_23605,N_22641,N_22292);
or U23606 (N_23606,N_22040,N_22605);
and U23607 (N_23607,N_22596,N_22555);
and U23608 (N_23608,N_22918,N_22786);
or U23609 (N_23609,N_22922,N_22814);
nor U23610 (N_23610,N_22636,N_22834);
nand U23611 (N_23611,N_22614,N_22457);
nand U23612 (N_23612,N_22276,N_22623);
and U23613 (N_23613,N_22036,N_22425);
nand U23614 (N_23614,N_22171,N_22006);
or U23615 (N_23615,N_22972,N_22009);
xnor U23616 (N_23616,N_22097,N_22384);
and U23617 (N_23617,N_22429,N_22666);
nor U23618 (N_23618,N_22939,N_22063);
nor U23619 (N_23619,N_22674,N_22253);
xnor U23620 (N_23620,N_22031,N_22252);
xnor U23621 (N_23621,N_22904,N_22855);
nand U23622 (N_23622,N_22881,N_22966);
nor U23623 (N_23623,N_22722,N_22945);
and U23624 (N_23624,N_22644,N_22636);
or U23625 (N_23625,N_22930,N_22874);
or U23626 (N_23626,N_22056,N_22490);
or U23627 (N_23627,N_22727,N_22152);
nor U23628 (N_23628,N_22519,N_22931);
and U23629 (N_23629,N_22945,N_22962);
or U23630 (N_23630,N_22552,N_22771);
xnor U23631 (N_23631,N_22035,N_22492);
nand U23632 (N_23632,N_22735,N_22854);
and U23633 (N_23633,N_22937,N_22319);
nor U23634 (N_23634,N_22392,N_22868);
nand U23635 (N_23635,N_22499,N_22120);
and U23636 (N_23636,N_22752,N_22959);
nor U23637 (N_23637,N_22419,N_22387);
xor U23638 (N_23638,N_22348,N_22812);
nor U23639 (N_23639,N_22282,N_22331);
xor U23640 (N_23640,N_22169,N_22081);
nand U23641 (N_23641,N_22189,N_22907);
or U23642 (N_23642,N_22436,N_22698);
or U23643 (N_23643,N_22502,N_22079);
nor U23644 (N_23644,N_22578,N_22038);
xor U23645 (N_23645,N_22932,N_22283);
or U23646 (N_23646,N_22897,N_22779);
nor U23647 (N_23647,N_22422,N_22304);
or U23648 (N_23648,N_22293,N_22760);
and U23649 (N_23649,N_22535,N_22473);
xnor U23650 (N_23650,N_22021,N_22084);
and U23651 (N_23651,N_22870,N_22088);
nand U23652 (N_23652,N_22561,N_22973);
nand U23653 (N_23653,N_22099,N_22428);
nand U23654 (N_23654,N_22909,N_22311);
nor U23655 (N_23655,N_22898,N_22468);
or U23656 (N_23656,N_22834,N_22442);
nor U23657 (N_23657,N_22202,N_22415);
nor U23658 (N_23658,N_22551,N_22806);
nand U23659 (N_23659,N_22627,N_22282);
or U23660 (N_23660,N_22656,N_22212);
nand U23661 (N_23661,N_22409,N_22303);
nor U23662 (N_23662,N_22427,N_22044);
or U23663 (N_23663,N_22343,N_22988);
nand U23664 (N_23664,N_22337,N_22009);
and U23665 (N_23665,N_22149,N_22143);
or U23666 (N_23666,N_22274,N_22857);
nor U23667 (N_23667,N_22049,N_22073);
xnor U23668 (N_23668,N_22463,N_22115);
and U23669 (N_23669,N_22503,N_22113);
nand U23670 (N_23670,N_22344,N_22372);
nor U23671 (N_23671,N_22890,N_22784);
or U23672 (N_23672,N_22667,N_22083);
nand U23673 (N_23673,N_22686,N_22009);
or U23674 (N_23674,N_22639,N_22267);
nor U23675 (N_23675,N_22745,N_22801);
xnor U23676 (N_23676,N_22081,N_22757);
nand U23677 (N_23677,N_22220,N_22403);
xor U23678 (N_23678,N_22785,N_22211);
xnor U23679 (N_23679,N_22687,N_22311);
xnor U23680 (N_23680,N_22447,N_22686);
and U23681 (N_23681,N_22930,N_22081);
nor U23682 (N_23682,N_22149,N_22233);
nor U23683 (N_23683,N_22263,N_22194);
and U23684 (N_23684,N_22549,N_22536);
or U23685 (N_23685,N_22109,N_22960);
nor U23686 (N_23686,N_22427,N_22382);
and U23687 (N_23687,N_22921,N_22524);
nand U23688 (N_23688,N_22301,N_22894);
and U23689 (N_23689,N_22930,N_22014);
xnor U23690 (N_23690,N_22333,N_22152);
nand U23691 (N_23691,N_22794,N_22350);
nor U23692 (N_23692,N_22968,N_22152);
nor U23693 (N_23693,N_22271,N_22790);
or U23694 (N_23694,N_22743,N_22627);
and U23695 (N_23695,N_22166,N_22029);
nor U23696 (N_23696,N_22387,N_22471);
or U23697 (N_23697,N_22384,N_22835);
nand U23698 (N_23698,N_22954,N_22933);
or U23699 (N_23699,N_22418,N_22036);
and U23700 (N_23700,N_22735,N_22706);
xnor U23701 (N_23701,N_22709,N_22708);
nand U23702 (N_23702,N_22090,N_22730);
nor U23703 (N_23703,N_22713,N_22056);
or U23704 (N_23704,N_22884,N_22742);
nor U23705 (N_23705,N_22643,N_22473);
nor U23706 (N_23706,N_22663,N_22090);
and U23707 (N_23707,N_22641,N_22383);
or U23708 (N_23708,N_22217,N_22944);
xnor U23709 (N_23709,N_22789,N_22075);
or U23710 (N_23710,N_22397,N_22122);
nor U23711 (N_23711,N_22409,N_22333);
xnor U23712 (N_23712,N_22243,N_22418);
nand U23713 (N_23713,N_22580,N_22600);
xor U23714 (N_23714,N_22327,N_22395);
xor U23715 (N_23715,N_22644,N_22702);
nand U23716 (N_23716,N_22047,N_22039);
xnor U23717 (N_23717,N_22126,N_22544);
xnor U23718 (N_23718,N_22639,N_22396);
and U23719 (N_23719,N_22266,N_22186);
and U23720 (N_23720,N_22757,N_22363);
xor U23721 (N_23721,N_22273,N_22285);
nand U23722 (N_23722,N_22942,N_22162);
xnor U23723 (N_23723,N_22727,N_22212);
xor U23724 (N_23724,N_22342,N_22171);
or U23725 (N_23725,N_22672,N_22442);
or U23726 (N_23726,N_22848,N_22805);
nand U23727 (N_23727,N_22709,N_22953);
xor U23728 (N_23728,N_22235,N_22400);
nor U23729 (N_23729,N_22312,N_22175);
nor U23730 (N_23730,N_22925,N_22149);
xnor U23731 (N_23731,N_22414,N_22682);
xnor U23732 (N_23732,N_22514,N_22509);
nand U23733 (N_23733,N_22398,N_22263);
xor U23734 (N_23734,N_22716,N_22110);
nand U23735 (N_23735,N_22666,N_22396);
or U23736 (N_23736,N_22207,N_22157);
xnor U23737 (N_23737,N_22303,N_22317);
or U23738 (N_23738,N_22002,N_22854);
nor U23739 (N_23739,N_22799,N_22749);
or U23740 (N_23740,N_22262,N_22837);
nor U23741 (N_23741,N_22856,N_22759);
nand U23742 (N_23742,N_22998,N_22913);
nand U23743 (N_23743,N_22375,N_22401);
nand U23744 (N_23744,N_22812,N_22566);
nor U23745 (N_23745,N_22126,N_22465);
nor U23746 (N_23746,N_22826,N_22267);
or U23747 (N_23747,N_22109,N_22348);
nand U23748 (N_23748,N_22038,N_22186);
or U23749 (N_23749,N_22147,N_22824);
xor U23750 (N_23750,N_22934,N_22657);
and U23751 (N_23751,N_22237,N_22512);
and U23752 (N_23752,N_22041,N_22074);
nor U23753 (N_23753,N_22708,N_22452);
xnor U23754 (N_23754,N_22780,N_22166);
nand U23755 (N_23755,N_22277,N_22828);
or U23756 (N_23756,N_22330,N_22687);
nand U23757 (N_23757,N_22904,N_22580);
and U23758 (N_23758,N_22258,N_22313);
nand U23759 (N_23759,N_22203,N_22620);
nor U23760 (N_23760,N_22462,N_22079);
nor U23761 (N_23761,N_22427,N_22617);
or U23762 (N_23762,N_22631,N_22316);
and U23763 (N_23763,N_22317,N_22063);
xnor U23764 (N_23764,N_22183,N_22427);
or U23765 (N_23765,N_22279,N_22960);
xnor U23766 (N_23766,N_22181,N_22288);
and U23767 (N_23767,N_22064,N_22768);
nand U23768 (N_23768,N_22093,N_22025);
xor U23769 (N_23769,N_22625,N_22847);
and U23770 (N_23770,N_22841,N_22066);
nor U23771 (N_23771,N_22400,N_22620);
xor U23772 (N_23772,N_22439,N_22557);
nor U23773 (N_23773,N_22389,N_22221);
or U23774 (N_23774,N_22636,N_22232);
xnor U23775 (N_23775,N_22181,N_22317);
and U23776 (N_23776,N_22566,N_22661);
nor U23777 (N_23777,N_22011,N_22032);
nand U23778 (N_23778,N_22412,N_22681);
nand U23779 (N_23779,N_22119,N_22517);
xnor U23780 (N_23780,N_22940,N_22159);
nor U23781 (N_23781,N_22122,N_22577);
nor U23782 (N_23782,N_22096,N_22893);
or U23783 (N_23783,N_22161,N_22846);
or U23784 (N_23784,N_22782,N_22495);
and U23785 (N_23785,N_22245,N_22674);
xnor U23786 (N_23786,N_22290,N_22781);
xnor U23787 (N_23787,N_22675,N_22209);
nor U23788 (N_23788,N_22794,N_22448);
xor U23789 (N_23789,N_22160,N_22385);
nor U23790 (N_23790,N_22440,N_22709);
or U23791 (N_23791,N_22567,N_22241);
nor U23792 (N_23792,N_22623,N_22175);
or U23793 (N_23793,N_22850,N_22701);
nand U23794 (N_23794,N_22020,N_22069);
nand U23795 (N_23795,N_22323,N_22648);
or U23796 (N_23796,N_22328,N_22003);
nand U23797 (N_23797,N_22215,N_22293);
and U23798 (N_23798,N_22497,N_22621);
and U23799 (N_23799,N_22437,N_22354);
nor U23800 (N_23800,N_22655,N_22317);
xnor U23801 (N_23801,N_22992,N_22328);
and U23802 (N_23802,N_22926,N_22257);
xor U23803 (N_23803,N_22581,N_22046);
or U23804 (N_23804,N_22107,N_22308);
xor U23805 (N_23805,N_22424,N_22694);
and U23806 (N_23806,N_22798,N_22875);
nor U23807 (N_23807,N_22326,N_22239);
and U23808 (N_23808,N_22800,N_22783);
xnor U23809 (N_23809,N_22568,N_22308);
nand U23810 (N_23810,N_22394,N_22129);
nor U23811 (N_23811,N_22110,N_22617);
xor U23812 (N_23812,N_22168,N_22051);
and U23813 (N_23813,N_22227,N_22540);
and U23814 (N_23814,N_22959,N_22397);
nor U23815 (N_23815,N_22595,N_22000);
nand U23816 (N_23816,N_22008,N_22075);
or U23817 (N_23817,N_22418,N_22584);
nand U23818 (N_23818,N_22499,N_22519);
and U23819 (N_23819,N_22649,N_22921);
nand U23820 (N_23820,N_22058,N_22919);
nor U23821 (N_23821,N_22825,N_22403);
or U23822 (N_23822,N_22317,N_22152);
and U23823 (N_23823,N_22147,N_22104);
nand U23824 (N_23824,N_22419,N_22165);
xor U23825 (N_23825,N_22979,N_22623);
nor U23826 (N_23826,N_22137,N_22000);
and U23827 (N_23827,N_22810,N_22628);
nand U23828 (N_23828,N_22818,N_22825);
or U23829 (N_23829,N_22886,N_22518);
and U23830 (N_23830,N_22610,N_22063);
nand U23831 (N_23831,N_22213,N_22133);
and U23832 (N_23832,N_22697,N_22150);
or U23833 (N_23833,N_22463,N_22118);
and U23834 (N_23834,N_22584,N_22562);
nor U23835 (N_23835,N_22764,N_22689);
or U23836 (N_23836,N_22501,N_22359);
nand U23837 (N_23837,N_22746,N_22878);
nor U23838 (N_23838,N_22455,N_22137);
and U23839 (N_23839,N_22763,N_22248);
xor U23840 (N_23840,N_22800,N_22451);
or U23841 (N_23841,N_22929,N_22797);
xnor U23842 (N_23842,N_22278,N_22319);
nor U23843 (N_23843,N_22302,N_22407);
nor U23844 (N_23844,N_22602,N_22419);
or U23845 (N_23845,N_22674,N_22158);
nor U23846 (N_23846,N_22054,N_22033);
and U23847 (N_23847,N_22485,N_22593);
nand U23848 (N_23848,N_22098,N_22470);
or U23849 (N_23849,N_22194,N_22118);
or U23850 (N_23850,N_22414,N_22541);
xor U23851 (N_23851,N_22942,N_22763);
nand U23852 (N_23852,N_22791,N_22556);
nand U23853 (N_23853,N_22404,N_22745);
nor U23854 (N_23854,N_22690,N_22607);
or U23855 (N_23855,N_22079,N_22103);
or U23856 (N_23856,N_22964,N_22109);
nand U23857 (N_23857,N_22754,N_22133);
or U23858 (N_23858,N_22103,N_22798);
xor U23859 (N_23859,N_22689,N_22735);
nor U23860 (N_23860,N_22290,N_22005);
nor U23861 (N_23861,N_22350,N_22520);
and U23862 (N_23862,N_22583,N_22616);
xor U23863 (N_23863,N_22493,N_22641);
nor U23864 (N_23864,N_22675,N_22855);
nor U23865 (N_23865,N_22523,N_22210);
nor U23866 (N_23866,N_22156,N_22589);
and U23867 (N_23867,N_22864,N_22035);
nor U23868 (N_23868,N_22593,N_22430);
xnor U23869 (N_23869,N_22192,N_22795);
xor U23870 (N_23870,N_22229,N_22706);
nor U23871 (N_23871,N_22758,N_22882);
and U23872 (N_23872,N_22667,N_22810);
nand U23873 (N_23873,N_22648,N_22053);
and U23874 (N_23874,N_22837,N_22298);
xor U23875 (N_23875,N_22441,N_22202);
xnor U23876 (N_23876,N_22158,N_22714);
nand U23877 (N_23877,N_22436,N_22246);
nand U23878 (N_23878,N_22251,N_22939);
and U23879 (N_23879,N_22781,N_22379);
xor U23880 (N_23880,N_22698,N_22157);
nor U23881 (N_23881,N_22129,N_22085);
nor U23882 (N_23882,N_22963,N_22344);
or U23883 (N_23883,N_22942,N_22002);
and U23884 (N_23884,N_22946,N_22987);
nand U23885 (N_23885,N_22393,N_22330);
or U23886 (N_23886,N_22971,N_22713);
and U23887 (N_23887,N_22431,N_22282);
and U23888 (N_23888,N_22382,N_22508);
xnor U23889 (N_23889,N_22026,N_22857);
xnor U23890 (N_23890,N_22841,N_22961);
or U23891 (N_23891,N_22059,N_22287);
or U23892 (N_23892,N_22090,N_22888);
nand U23893 (N_23893,N_22245,N_22965);
or U23894 (N_23894,N_22162,N_22527);
nor U23895 (N_23895,N_22205,N_22161);
and U23896 (N_23896,N_22489,N_22543);
or U23897 (N_23897,N_22214,N_22983);
xor U23898 (N_23898,N_22700,N_22410);
and U23899 (N_23899,N_22426,N_22901);
and U23900 (N_23900,N_22714,N_22458);
or U23901 (N_23901,N_22909,N_22566);
xor U23902 (N_23902,N_22605,N_22811);
nor U23903 (N_23903,N_22863,N_22041);
nand U23904 (N_23904,N_22898,N_22614);
xnor U23905 (N_23905,N_22722,N_22706);
and U23906 (N_23906,N_22615,N_22579);
or U23907 (N_23907,N_22021,N_22279);
or U23908 (N_23908,N_22887,N_22012);
nand U23909 (N_23909,N_22943,N_22791);
and U23910 (N_23910,N_22874,N_22077);
and U23911 (N_23911,N_22698,N_22310);
and U23912 (N_23912,N_22756,N_22515);
nand U23913 (N_23913,N_22217,N_22557);
nor U23914 (N_23914,N_22956,N_22759);
or U23915 (N_23915,N_22815,N_22656);
or U23916 (N_23916,N_22800,N_22641);
and U23917 (N_23917,N_22019,N_22929);
nor U23918 (N_23918,N_22633,N_22115);
and U23919 (N_23919,N_22391,N_22209);
nand U23920 (N_23920,N_22657,N_22023);
nand U23921 (N_23921,N_22841,N_22436);
and U23922 (N_23922,N_22945,N_22969);
nor U23923 (N_23923,N_22431,N_22856);
and U23924 (N_23924,N_22713,N_22292);
nand U23925 (N_23925,N_22307,N_22095);
xor U23926 (N_23926,N_22861,N_22547);
nor U23927 (N_23927,N_22860,N_22305);
xor U23928 (N_23928,N_22471,N_22559);
nand U23929 (N_23929,N_22983,N_22111);
nand U23930 (N_23930,N_22113,N_22065);
nor U23931 (N_23931,N_22401,N_22154);
or U23932 (N_23932,N_22995,N_22893);
or U23933 (N_23933,N_22391,N_22640);
and U23934 (N_23934,N_22493,N_22328);
or U23935 (N_23935,N_22721,N_22560);
or U23936 (N_23936,N_22547,N_22867);
or U23937 (N_23937,N_22868,N_22748);
nand U23938 (N_23938,N_22066,N_22691);
and U23939 (N_23939,N_22939,N_22692);
xor U23940 (N_23940,N_22078,N_22126);
nor U23941 (N_23941,N_22981,N_22837);
nor U23942 (N_23942,N_22008,N_22432);
nor U23943 (N_23943,N_22853,N_22891);
nor U23944 (N_23944,N_22370,N_22054);
and U23945 (N_23945,N_22231,N_22856);
or U23946 (N_23946,N_22698,N_22260);
and U23947 (N_23947,N_22218,N_22568);
and U23948 (N_23948,N_22643,N_22496);
or U23949 (N_23949,N_22512,N_22390);
and U23950 (N_23950,N_22812,N_22514);
nor U23951 (N_23951,N_22987,N_22566);
xor U23952 (N_23952,N_22686,N_22833);
nor U23953 (N_23953,N_22587,N_22881);
xnor U23954 (N_23954,N_22149,N_22471);
nor U23955 (N_23955,N_22692,N_22679);
nand U23956 (N_23956,N_22908,N_22458);
or U23957 (N_23957,N_22140,N_22980);
xor U23958 (N_23958,N_22344,N_22680);
nor U23959 (N_23959,N_22208,N_22198);
xnor U23960 (N_23960,N_22997,N_22251);
nand U23961 (N_23961,N_22094,N_22190);
xnor U23962 (N_23962,N_22857,N_22471);
or U23963 (N_23963,N_22028,N_22250);
xnor U23964 (N_23964,N_22251,N_22257);
and U23965 (N_23965,N_22155,N_22964);
nor U23966 (N_23966,N_22163,N_22754);
xor U23967 (N_23967,N_22428,N_22811);
or U23968 (N_23968,N_22649,N_22321);
xor U23969 (N_23969,N_22157,N_22522);
nor U23970 (N_23970,N_22495,N_22976);
and U23971 (N_23971,N_22017,N_22646);
or U23972 (N_23972,N_22116,N_22563);
nor U23973 (N_23973,N_22025,N_22250);
nand U23974 (N_23974,N_22909,N_22130);
nor U23975 (N_23975,N_22218,N_22821);
and U23976 (N_23976,N_22774,N_22998);
and U23977 (N_23977,N_22981,N_22449);
nor U23978 (N_23978,N_22252,N_22436);
or U23979 (N_23979,N_22518,N_22918);
or U23980 (N_23980,N_22953,N_22315);
nor U23981 (N_23981,N_22756,N_22526);
nor U23982 (N_23982,N_22119,N_22391);
and U23983 (N_23983,N_22683,N_22347);
nand U23984 (N_23984,N_22914,N_22013);
or U23985 (N_23985,N_22175,N_22591);
and U23986 (N_23986,N_22768,N_22150);
nand U23987 (N_23987,N_22518,N_22287);
xnor U23988 (N_23988,N_22192,N_22847);
xor U23989 (N_23989,N_22231,N_22433);
nor U23990 (N_23990,N_22617,N_22495);
or U23991 (N_23991,N_22182,N_22102);
or U23992 (N_23992,N_22837,N_22843);
nor U23993 (N_23993,N_22474,N_22428);
or U23994 (N_23994,N_22160,N_22797);
or U23995 (N_23995,N_22860,N_22470);
nor U23996 (N_23996,N_22920,N_22953);
xnor U23997 (N_23997,N_22350,N_22623);
nor U23998 (N_23998,N_22785,N_22768);
nand U23999 (N_23999,N_22781,N_22277);
xor U24000 (N_24000,N_23748,N_23638);
nand U24001 (N_24001,N_23344,N_23622);
and U24002 (N_24002,N_23330,N_23438);
nand U24003 (N_24003,N_23113,N_23349);
nor U24004 (N_24004,N_23908,N_23375);
and U24005 (N_24005,N_23241,N_23271);
xnor U24006 (N_24006,N_23810,N_23140);
or U24007 (N_24007,N_23822,N_23726);
nor U24008 (N_24008,N_23343,N_23619);
nor U24009 (N_24009,N_23813,N_23503);
nand U24010 (N_24010,N_23450,N_23099);
nor U24011 (N_24011,N_23197,N_23529);
or U24012 (N_24012,N_23571,N_23307);
nor U24013 (N_24013,N_23646,N_23969);
or U24014 (N_24014,N_23968,N_23776);
or U24015 (N_24015,N_23561,N_23306);
nand U24016 (N_24016,N_23878,N_23530);
nor U24017 (N_24017,N_23870,N_23556);
xnor U24018 (N_24018,N_23889,N_23335);
and U24019 (N_24019,N_23996,N_23441);
and U24020 (N_24020,N_23742,N_23225);
xor U24021 (N_24021,N_23366,N_23336);
xor U24022 (N_24022,N_23210,N_23934);
nor U24023 (N_24023,N_23141,N_23370);
nand U24024 (N_24024,N_23784,N_23679);
or U24025 (N_24025,N_23924,N_23753);
nor U24026 (N_24026,N_23567,N_23433);
xor U24027 (N_24027,N_23300,N_23605);
nor U24028 (N_24028,N_23329,N_23513);
nor U24029 (N_24029,N_23305,N_23904);
nand U24030 (N_24030,N_23475,N_23712);
xor U24031 (N_24031,N_23175,N_23490);
or U24032 (N_24032,N_23518,N_23055);
nand U24033 (N_24033,N_23695,N_23459);
xnor U24034 (N_24034,N_23224,N_23069);
or U24035 (N_24035,N_23642,N_23521);
or U24036 (N_24036,N_23121,N_23227);
nand U24037 (N_24037,N_23458,N_23684);
nand U24038 (N_24038,N_23002,N_23570);
and U24039 (N_24039,N_23692,N_23274);
nand U24040 (N_24040,N_23579,N_23858);
or U24041 (N_24041,N_23593,N_23451);
and U24042 (N_24042,N_23833,N_23364);
nand U24043 (N_24043,N_23671,N_23043);
xnor U24044 (N_24044,N_23010,N_23954);
nor U24045 (N_24045,N_23909,N_23818);
and U24046 (N_24046,N_23406,N_23417);
xnor U24047 (N_24047,N_23469,N_23738);
xnor U24048 (N_24048,N_23412,N_23708);
or U24049 (N_24049,N_23755,N_23232);
nand U24050 (N_24050,N_23609,N_23396);
and U24051 (N_24051,N_23394,N_23104);
nor U24052 (N_24052,N_23269,N_23114);
and U24053 (N_24053,N_23920,N_23297);
nor U24054 (N_24054,N_23144,N_23186);
nand U24055 (N_24055,N_23097,N_23844);
or U24056 (N_24056,N_23369,N_23656);
xor U24057 (N_24057,N_23301,N_23201);
nor U24058 (N_24058,N_23273,N_23725);
nor U24059 (N_24059,N_23624,N_23047);
xnor U24060 (N_24060,N_23156,N_23773);
and U24061 (N_24061,N_23495,N_23082);
and U24062 (N_24062,N_23506,N_23351);
xor U24063 (N_24063,N_23399,N_23194);
nor U24064 (N_24064,N_23426,N_23942);
and U24065 (N_24065,N_23100,N_23633);
nand U24066 (N_24066,N_23196,N_23480);
or U24067 (N_24067,N_23652,N_23309);
xnor U24068 (N_24068,N_23294,N_23084);
nand U24069 (N_24069,N_23740,N_23377);
or U24070 (N_24070,N_23255,N_23544);
nand U24071 (N_24071,N_23569,N_23325);
nor U24072 (N_24072,N_23699,N_23973);
xor U24073 (N_24073,N_23400,N_23950);
nand U24074 (N_24074,N_23859,N_23541);
nor U24075 (N_24075,N_23006,N_23487);
and U24076 (N_24076,N_23632,N_23922);
nor U24077 (N_24077,N_23660,N_23425);
xor U24078 (N_24078,N_23392,N_23110);
or U24079 (N_24079,N_23543,N_23875);
and U24080 (N_24080,N_23508,N_23342);
nor U24081 (N_24081,N_23857,N_23333);
nor U24082 (N_24082,N_23731,N_23431);
and U24083 (N_24083,N_23191,N_23730);
or U24084 (N_24084,N_23783,N_23957);
or U24085 (N_24085,N_23038,N_23226);
nor U24086 (N_24086,N_23239,N_23222);
nor U24087 (N_24087,N_23621,N_23162);
nor U24088 (N_24088,N_23310,N_23161);
and U24089 (N_24089,N_23296,N_23603);
xor U24090 (N_24090,N_23018,N_23492);
nand U24091 (N_24091,N_23563,N_23163);
and U24092 (N_24092,N_23644,N_23456);
nand U24093 (N_24093,N_23353,N_23963);
or U24094 (N_24094,N_23248,N_23661);
nor U24095 (N_24095,N_23802,N_23068);
nand U24096 (N_24096,N_23277,N_23929);
and U24097 (N_24097,N_23065,N_23581);
nor U24098 (N_24098,N_23295,N_23494);
and U24099 (N_24099,N_23597,N_23443);
and U24100 (N_24100,N_23537,N_23378);
xor U24101 (N_24101,N_23686,N_23205);
and U24102 (N_24102,N_23463,N_23976);
nor U24103 (N_24103,N_23631,N_23505);
and U24104 (N_24104,N_23359,N_23989);
xnor U24105 (N_24105,N_23702,N_23614);
or U24106 (N_24106,N_23860,N_23123);
nand U24107 (N_24107,N_23618,N_23538);
xnor U24108 (N_24108,N_23265,N_23474);
nor U24109 (N_24109,N_23437,N_23217);
and U24110 (N_24110,N_23171,N_23466);
nand U24111 (N_24111,N_23982,N_23944);
nor U24112 (N_24112,N_23135,N_23629);
or U24113 (N_24113,N_23497,N_23083);
nand U24114 (N_24114,N_23781,N_23917);
or U24115 (N_24115,N_23796,N_23423);
nor U24116 (N_24116,N_23283,N_23160);
and U24117 (N_24117,N_23173,N_23254);
and U24118 (N_24118,N_23133,N_23914);
or U24119 (N_24119,N_23007,N_23230);
nor U24120 (N_24120,N_23106,N_23941);
or U24121 (N_24121,N_23384,N_23233);
xnor U24122 (N_24122,N_23293,N_23899);
nand U24123 (N_24123,N_23720,N_23798);
xor U24124 (N_24124,N_23876,N_23620);
nand U24125 (N_24125,N_23872,N_23312);
xnor U24126 (N_24126,N_23498,N_23547);
nor U24127 (N_24127,N_23211,N_23303);
nand U24128 (N_24128,N_23484,N_23677);
and U24129 (N_24129,N_23235,N_23522);
nor U24130 (N_24130,N_23088,N_23081);
and U24131 (N_24131,N_23535,N_23984);
xnor U24132 (N_24132,N_23752,N_23031);
nand U24133 (N_24133,N_23252,N_23473);
nor U24134 (N_24134,N_23797,N_23409);
or U24135 (N_24135,N_23866,N_23835);
nand U24136 (N_24136,N_23940,N_23648);
xor U24137 (N_24137,N_23395,N_23855);
nor U24138 (N_24138,N_23849,N_23769);
or U24139 (N_24139,N_23789,N_23843);
and U24140 (N_24140,N_23383,N_23869);
xnor U24141 (N_24141,N_23767,N_23771);
xnor U24142 (N_24142,N_23542,N_23777);
and U24143 (N_24143,N_23072,N_23562);
or U24144 (N_24144,N_23019,N_23694);
and U24145 (N_24145,N_23650,N_23288);
and U24146 (N_24146,N_23026,N_23788);
xor U24147 (N_24147,N_23009,N_23625);
nand U24148 (N_24148,N_23604,N_23534);
xnor U24149 (N_24149,N_23095,N_23645);
and U24150 (N_24150,N_23687,N_23812);
xor U24151 (N_24151,N_23402,N_23896);
nand U24152 (N_24152,N_23707,N_23246);
and U24153 (N_24153,N_23683,N_23137);
nand U24154 (N_24154,N_23017,N_23829);
and U24155 (N_24155,N_23555,N_23219);
xor U24156 (N_24156,N_23820,N_23884);
or U24157 (N_24157,N_23256,N_23129);
nand U24158 (N_24158,N_23127,N_23637);
or U24159 (N_24159,N_23803,N_23643);
and U24160 (N_24160,N_23496,N_23594);
xnor U24161 (N_24161,N_23167,N_23061);
xnor U24162 (N_24162,N_23454,N_23046);
nand U24163 (N_24163,N_23733,N_23356);
xnor U24164 (N_24164,N_23589,N_23240);
or U24165 (N_24165,N_23745,N_23736);
xnor U24166 (N_24166,N_23856,N_23413);
xor U24167 (N_24167,N_23471,N_23037);
nand U24168 (N_24168,N_23952,N_23805);
nor U24169 (N_24169,N_23049,N_23410);
and U24170 (N_24170,N_23094,N_23415);
nor U24171 (N_24171,N_23758,N_23582);
or U24172 (N_24172,N_23299,N_23887);
xnor U24173 (N_24173,N_23890,N_23981);
nand U24174 (N_24174,N_23724,N_23659);
and U24175 (N_24175,N_23615,N_23690);
nor U24176 (N_24176,N_23174,N_23602);
nand U24177 (N_24177,N_23931,N_23445);
xor U24178 (N_24178,N_23845,N_23338);
and U24179 (N_24179,N_23770,N_23735);
nor U24180 (N_24180,N_23024,N_23236);
nor U24181 (N_24181,N_23190,N_23568);
and U24182 (N_24182,N_23001,N_23444);
and U24183 (N_24183,N_23220,N_23536);
and U24184 (N_24184,N_23765,N_23979);
xor U24185 (N_24185,N_23022,N_23251);
xor U24186 (N_24186,N_23257,N_23838);
xnor U24187 (N_24187,N_23937,N_23640);
xor U24188 (N_24188,N_23754,N_23716);
and U24189 (N_24189,N_23959,N_23282);
nor U24190 (N_24190,N_23169,N_23290);
xor U24191 (N_24191,N_23033,N_23528);
xnor U24192 (N_24192,N_23961,N_23780);
xnor U24193 (N_24193,N_23397,N_23587);
or U24194 (N_24194,N_23675,N_23158);
or U24195 (N_24195,N_23322,N_23907);
nand U24196 (N_24196,N_23964,N_23749);
nor U24197 (N_24197,N_23595,N_23653);
nand U24198 (N_24198,N_23831,N_23418);
nor U24199 (N_24199,N_23063,N_23086);
or U24200 (N_24200,N_23268,N_23548);
and U24201 (N_24201,N_23560,N_23928);
xnor U24202 (N_24202,N_23314,N_23811);
and U24203 (N_24203,N_23793,N_23678);
and U24204 (N_24204,N_23885,N_23125);
or U24205 (N_24205,N_23434,N_23967);
or U24206 (N_24206,N_23546,N_23539);
nor U24207 (N_24207,N_23786,N_23662);
and U24208 (N_24208,N_23421,N_23554);
and U24209 (N_24209,N_23170,N_23216);
nor U24210 (N_24210,N_23936,N_23391);
nand U24211 (N_24211,N_23477,N_23586);
nor U24212 (N_24212,N_23817,N_23382);
nand U24213 (N_24213,N_23292,N_23746);
nor U24214 (N_24214,N_23639,N_23946);
nand U24215 (N_24215,N_23237,N_23590);
or U24216 (N_24216,N_23898,N_23098);
and U24217 (N_24217,N_23926,N_23634);
or U24218 (N_24218,N_23516,N_23883);
xor U24219 (N_24219,N_23368,N_23130);
xnor U24220 (N_24220,N_23500,N_23118);
and U24221 (N_24221,N_23575,N_23092);
nand U24222 (N_24222,N_23672,N_23668);
nor U24223 (N_24223,N_23109,N_23892);
xnor U24224 (N_24224,N_23150,N_23628);
and U24225 (N_24225,N_23682,N_23839);
or U24226 (N_24226,N_23131,N_23461);
nor U24227 (N_24227,N_23930,N_23401);
xnor U24228 (N_24228,N_23040,N_23956);
nor U24229 (N_24229,N_23440,N_23693);
and U24230 (N_24230,N_23717,N_23550);
and U24231 (N_24231,N_23916,N_23840);
nand U24232 (N_24232,N_23111,N_23278);
and U24233 (N_24233,N_23572,N_23116);
nor U24234 (N_24234,N_23734,N_23374);
and U24235 (N_24235,N_23371,N_23923);
xor U24236 (N_24236,N_23919,N_23862);
or U24237 (N_24237,N_23393,N_23341);
nor U24238 (N_24238,N_23520,N_23050);
xnor U24239 (N_24239,N_23103,N_23332);
and U24240 (N_24240,N_23654,N_23585);
xnor U24241 (N_24241,N_23258,N_23795);
nand U24242 (N_24242,N_23517,N_23779);
xnor U24243 (N_24243,N_23148,N_23549);
nand U24244 (N_24244,N_23302,N_23483);
nand U24245 (N_24245,N_23361,N_23760);
xor U24246 (N_24246,N_23172,N_23138);
xor U24247 (N_24247,N_23367,N_23387);
and U24248 (N_24248,N_23218,N_23380);
xnor U24249 (N_24249,N_23943,N_23179);
and U24250 (N_24250,N_23253,N_23819);
nor U24251 (N_24251,N_23326,N_23407);
nand U24252 (N_24252,N_23918,N_23067);
xor U24253 (N_24253,N_23446,N_23180);
nor U24254 (N_24254,N_23192,N_23991);
xnor U24255 (N_24255,N_23214,N_23193);
or U24256 (N_24256,N_23939,N_23023);
nand U24257 (N_24257,N_23790,N_23317);
or U24258 (N_24258,N_23807,N_23348);
or U24259 (N_24259,N_23510,N_23910);
nor U24260 (N_24260,N_23763,N_23977);
and U24261 (N_24261,N_23373,N_23455);
nor U24262 (N_24262,N_23076,N_23729);
nor U24263 (N_24263,N_23608,N_23264);
nor U24264 (N_24264,N_23090,N_23559);
or U24265 (N_24265,N_23379,N_23958);
xor U24266 (N_24266,N_23524,N_23705);
xnor U24267 (N_24267,N_23424,N_23995);
or U24268 (N_24268,N_23003,N_23911);
xor U24269 (N_24269,N_23584,N_23809);
nand U24270 (N_24270,N_23250,N_23921);
and U24271 (N_24271,N_23328,N_23867);
or U24272 (N_24272,N_23276,N_23155);
nand U24273 (N_24273,N_23741,N_23863);
or U24274 (N_24274,N_23664,N_23029);
or U24275 (N_24275,N_23323,N_23347);
or U24276 (N_24276,N_23073,N_23154);
and U24277 (N_24277,N_23994,N_23157);
nor U24278 (N_24278,N_23533,N_23365);
xor U24279 (N_24279,N_23757,N_23165);
nor U24280 (N_24280,N_23189,N_23178);
and U24281 (N_24281,N_23853,N_23281);
nor U24282 (N_24282,N_23071,N_23102);
xor U24283 (N_24283,N_23501,N_23962);
nor U24284 (N_24284,N_23949,N_23657);
nor U24285 (N_24285,N_23107,N_23478);
and U24286 (N_24286,N_23526,N_23195);
xnor U24287 (N_24287,N_23039,N_23551);
xor U24288 (N_24288,N_23901,N_23245);
nor U24289 (N_24289,N_23053,N_23821);
or U24290 (N_24290,N_23275,N_23999);
and U24291 (N_24291,N_23126,N_23626);
or U24292 (N_24292,N_23851,N_23703);
or U24293 (N_24293,N_23270,N_23184);
and U24294 (N_24294,N_23512,N_23128);
xnor U24295 (N_24295,N_23457,N_23641);
nor U24296 (N_24296,N_23945,N_23915);
and U24297 (N_24297,N_23698,N_23052);
and U24298 (N_24298,N_23404,N_23827);
nor U24299 (N_24299,N_23011,N_23249);
nand U24300 (N_24300,N_23489,N_23826);
or U24301 (N_24301,N_23188,N_23578);
nand U24302 (N_24302,N_23491,N_23966);
nand U24303 (N_24303,N_23636,N_23079);
xor U24304 (N_24304,N_23481,N_23948);
or U24305 (N_24305,N_23873,N_23286);
or U24306 (N_24306,N_23493,N_23714);
and U24307 (N_24307,N_23509,N_23223);
or U24308 (N_24308,N_23352,N_23381);
or U24309 (N_24309,N_23244,N_23566);
nor U24310 (N_24310,N_23564,N_23647);
xnor U24311 (N_24311,N_23327,N_23975);
nand U24312 (N_24312,N_23136,N_23231);
nand U24313 (N_24313,N_23965,N_23261);
or U24314 (N_24314,N_23722,N_23048);
or U24315 (N_24315,N_23337,N_23091);
nand U24316 (N_24316,N_23432,N_23600);
xor U24317 (N_24317,N_23468,N_23987);
nand U24318 (N_24318,N_23439,N_23861);
nor U24319 (N_24319,N_23577,N_23247);
and U24320 (N_24320,N_23649,N_23658);
xnor U24321 (N_24321,N_23674,N_23616);
or U24322 (N_24322,N_23280,N_23764);
or U24323 (N_24323,N_23842,N_23778);
or U24324 (N_24324,N_23350,N_23830);
or U24325 (N_24325,N_23666,N_23263);
xor U24326 (N_24326,N_23713,N_23519);
and U24327 (N_24327,N_23854,N_23895);
nor U24328 (N_24328,N_23836,N_23685);
nor U24329 (N_24329,N_23514,N_23891);
xnor U24330 (N_24330,N_23960,N_23787);
nor U24331 (N_24331,N_23164,N_23215);
nand U24332 (N_24332,N_23146,N_23362);
and U24333 (N_24333,N_23837,N_23354);
and U24334 (N_24334,N_23176,N_23689);
nand U24335 (N_24335,N_23363,N_23502);
xor U24336 (N_24336,N_23428,N_23208);
nor U24337 (N_24337,N_23670,N_23202);
nor U24338 (N_24338,N_23183,N_23613);
or U24339 (N_24339,N_23667,N_23004);
nand U24340 (N_24340,N_23750,N_23598);
or U24341 (N_24341,N_23447,N_23070);
or U24342 (N_24342,N_23846,N_23986);
nor U24343 (N_24343,N_23591,N_23185);
nor U24344 (N_24344,N_23800,N_23893);
and U24345 (N_24345,N_23558,N_23515);
or U24346 (N_24346,N_23711,N_23243);
or U24347 (N_24347,N_23997,N_23864);
and U24348 (N_24348,N_23630,N_23436);
nand U24349 (N_24349,N_23229,N_23078);
xor U24350 (N_24350,N_23772,N_23452);
nand U24351 (N_24351,N_23988,N_23700);
nand U24352 (N_24352,N_23877,N_23990);
or U24353 (N_24353,N_23576,N_23774);
nand U24354 (N_24354,N_23422,N_23152);
xor U24355 (N_24355,N_23723,N_23304);
or U24356 (N_24356,N_23120,N_23311);
nor U24357 (N_24357,N_23834,N_23782);
and U24358 (N_24358,N_23499,N_23291);
xor U24359 (N_24359,N_23766,N_23540);
nor U24360 (N_24360,N_23978,N_23971);
nand U24361 (N_24361,N_23992,N_23467);
or U24362 (N_24362,N_23358,N_23177);
nor U24363 (N_24363,N_23228,N_23955);
or U24364 (N_24364,N_23785,N_23709);
nand U24365 (N_24365,N_23112,N_23565);
nor U24366 (N_24366,N_23035,N_23187);
and U24367 (N_24367,N_23611,N_23881);
nand U24368 (N_24368,N_23238,N_23768);
nand U24369 (N_24369,N_23420,N_23847);
or U24370 (N_24370,N_23479,N_23612);
or U24371 (N_24371,N_23430,N_23021);
and U24372 (N_24372,N_23080,N_23599);
and U24373 (N_24373,N_23761,N_23824);
nand U24374 (N_24374,N_23912,N_23606);
or U24375 (N_24375,N_23744,N_23020);
nor U24376 (N_24376,N_23886,N_23815);
or U24377 (N_24377,N_23028,N_23013);
xnor U24378 (N_24378,N_23719,N_23429);
nor U24379 (N_24379,N_23879,N_23791);
and U24380 (N_24380,N_23848,N_23357);
nor U24381 (N_24381,N_23718,N_23315);
xnor U24382 (N_24382,N_23775,N_23209);
nand U24383 (N_24383,N_23408,N_23124);
and U24384 (N_24384,N_23925,N_23673);
and U24385 (N_24385,N_23034,N_23823);
nor U24386 (N_24386,N_23262,N_23903);
or U24387 (N_24387,N_23865,N_23372);
and U24388 (N_24388,N_23610,N_23108);
nor U24389 (N_24389,N_23287,N_23284);
xor U24390 (N_24390,N_23448,N_23727);
or U24391 (N_24391,N_23181,N_23308);
nor U24392 (N_24392,N_23117,N_23405);
xnor U24393 (N_24393,N_23340,N_23145);
and U24394 (N_24394,N_23828,N_23472);
or U24395 (N_24395,N_23132,N_23388);
and U24396 (N_24396,N_23663,N_23168);
xor U24397 (N_24397,N_23974,N_23607);
nor U24398 (N_24398,N_23665,N_23696);
nor U24399 (N_24399,N_23453,N_23042);
nor U24400 (N_24400,N_23360,N_23557);
nor U24401 (N_24401,N_23932,N_23321);
and U24402 (N_24402,N_23045,N_23355);
nor U24403 (N_24403,N_23669,N_23583);
and U24404 (N_24404,N_23651,N_23016);
nand U24405 (N_24405,N_23882,N_23427);
nor U24406 (N_24406,N_23710,N_23119);
nor U24407 (N_24407,N_23200,N_23320);
or U24408 (N_24408,N_23897,N_23743);
nand U24409 (N_24409,N_23464,N_23051);
nor U24410 (N_24410,N_23234,N_23204);
or U24411 (N_24411,N_23390,N_23850);
xnor U24412 (N_24412,N_23139,N_23462);
nor U24413 (N_24413,N_23087,N_23970);
xnor U24414 (N_24414,N_23093,N_23025);
and U24415 (N_24415,N_23953,N_23319);
and U24416 (N_24416,N_23331,N_23266);
or U24417 (N_24417,N_23935,N_23085);
nor U24418 (N_24418,N_23313,N_23816);
xnor U24419 (N_24419,N_23627,N_23801);
and U24420 (N_24420,N_23721,N_23596);
nor U24421 (N_24421,N_23066,N_23507);
or U24422 (N_24422,N_23058,N_23096);
nand U24423 (N_24423,N_23985,N_23077);
and U24424 (N_24424,N_23635,N_23905);
or U24425 (N_24425,N_23617,N_23166);
xnor U24426 (N_24426,N_23318,N_23676);
nor U24427 (N_24427,N_23900,N_23880);
or U24428 (N_24428,N_23792,N_23386);
and U24429 (N_24429,N_23825,N_23101);
and U24430 (N_24430,N_23206,N_23588);
or U24431 (N_24431,N_23523,N_23060);
or U24432 (N_24432,N_23913,N_23623);
and U24433 (N_24433,N_23142,N_23005);
and U24434 (N_24434,N_23115,N_23527);
nor U24435 (N_24435,N_23159,N_23075);
and U24436 (N_24436,N_23376,N_23655);
nand U24437 (N_24437,N_23041,N_23927);
nor U24438 (N_24438,N_23756,N_23704);
xor U24439 (N_24439,N_23691,N_23601);
xnor U24440 (N_24440,N_23852,N_23947);
and U24441 (N_24441,N_23794,N_23014);
or U24442 (N_24442,N_23751,N_23339);
and U24443 (N_24443,N_23983,N_23762);
nor U24444 (N_24444,N_23532,N_23681);
xor U24445 (N_24445,N_23151,N_23574);
nand U24446 (N_24446,N_23054,N_23874);
or U24447 (N_24447,N_23182,N_23398);
nor U24448 (N_24448,N_23147,N_23411);
nand U24449 (N_24449,N_23346,N_23064);
and U24450 (N_24450,N_23012,N_23841);
and U24451 (N_24451,N_23153,N_23998);
nand U24452 (N_24452,N_23938,N_23199);
nand U24453 (N_24453,N_23089,N_23486);
nand U24454 (N_24454,N_23573,N_23272);
or U24455 (N_24455,N_23799,N_23808);
xor U24456 (N_24456,N_23894,N_23706);
xnor U24457 (N_24457,N_23580,N_23980);
or U24458 (N_24458,N_23134,N_23385);
nand U24459 (N_24459,N_23902,N_23008);
or U24460 (N_24460,N_23122,N_23525);
nand U24461 (N_24461,N_23056,N_23149);
xnor U24462 (N_24462,N_23485,N_23747);
or U24463 (N_24463,N_23972,N_23511);
xnor U24464 (N_24464,N_23260,N_23553);
and U24465 (N_24465,N_23465,N_23488);
and U24466 (N_24466,N_23015,N_23531);
nand U24467 (N_24467,N_23739,N_23298);
or U24468 (N_24468,N_23221,N_23806);
or U24469 (N_24469,N_23203,N_23267);
nand U24470 (N_24470,N_23403,N_23832);
or U24471 (N_24471,N_23552,N_23993);
and U24472 (N_24472,N_23285,N_23728);
xor U24473 (N_24473,N_23814,N_23030);
xnor U24474 (N_24474,N_23105,N_23759);
and U24475 (N_24475,N_23482,N_23435);
xnor U24476 (N_24476,N_23074,N_23414);
xor U24477 (N_24477,N_23476,N_23868);
xnor U24478 (N_24478,N_23198,N_23460);
or U24479 (N_24479,N_23242,N_23213);
and U24480 (N_24480,N_23334,N_23057);
nor U24481 (N_24481,N_23688,N_23888);
nand U24482 (N_24482,N_23737,N_23279);
nand U24483 (N_24483,N_23951,N_23804);
xor U24484 (N_24484,N_23449,N_23545);
and U24485 (N_24485,N_23207,N_23143);
or U24486 (N_24486,N_23715,N_23871);
or U24487 (N_24487,N_23062,N_23697);
nor U24488 (N_24488,N_23389,N_23592);
nor U24489 (N_24489,N_23470,N_23036);
and U24490 (N_24490,N_23316,N_23442);
or U24491 (N_24491,N_23212,N_23059);
xor U24492 (N_24492,N_23259,N_23732);
and U24493 (N_24493,N_23000,N_23324);
nand U24494 (N_24494,N_23419,N_23680);
xnor U24495 (N_24495,N_23701,N_23416);
xnor U24496 (N_24496,N_23933,N_23032);
or U24497 (N_24497,N_23345,N_23289);
xnor U24498 (N_24498,N_23044,N_23027);
and U24499 (N_24499,N_23504,N_23906);
nand U24500 (N_24500,N_23313,N_23035);
nor U24501 (N_24501,N_23387,N_23246);
nand U24502 (N_24502,N_23288,N_23817);
or U24503 (N_24503,N_23398,N_23024);
or U24504 (N_24504,N_23069,N_23774);
or U24505 (N_24505,N_23352,N_23511);
and U24506 (N_24506,N_23162,N_23396);
nor U24507 (N_24507,N_23206,N_23890);
nand U24508 (N_24508,N_23315,N_23241);
xor U24509 (N_24509,N_23199,N_23245);
or U24510 (N_24510,N_23967,N_23597);
nand U24511 (N_24511,N_23292,N_23867);
nor U24512 (N_24512,N_23211,N_23301);
and U24513 (N_24513,N_23387,N_23547);
xor U24514 (N_24514,N_23401,N_23104);
or U24515 (N_24515,N_23298,N_23770);
nand U24516 (N_24516,N_23754,N_23023);
xnor U24517 (N_24517,N_23671,N_23331);
nand U24518 (N_24518,N_23307,N_23736);
or U24519 (N_24519,N_23520,N_23570);
nand U24520 (N_24520,N_23258,N_23893);
xor U24521 (N_24521,N_23357,N_23672);
nand U24522 (N_24522,N_23119,N_23127);
and U24523 (N_24523,N_23167,N_23678);
nor U24524 (N_24524,N_23297,N_23697);
or U24525 (N_24525,N_23569,N_23508);
and U24526 (N_24526,N_23851,N_23407);
nand U24527 (N_24527,N_23266,N_23296);
nand U24528 (N_24528,N_23924,N_23045);
nand U24529 (N_24529,N_23928,N_23143);
and U24530 (N_24530,N_23330,N_23147);
or U24531 (N_24531,N_23249,N_23893);
and U24532 (N_24532,N_23276,N_23410);
xor U24533 (N_24533,N_23694,N_23338);
and U24534 (N_24534,N_23567,N_23830);
nand U24535 (N_24535,N_23597,N_23115);
xor U24536 (N_24536,N_23068,N_23940);
and U24537 (N_24537,N_23599,N_23415);
nor U24538 (N_24538,N_23598,N_23327);
or U24539 (N_24539,N_23582,N_23157);
or U24540 (N_24540,N_23277,N_23265);
nor U24541 (N_24541,N_23937,N_23265);
nand U24542 (N_24542,N_23923,N_23329);
xnor U24543 (N_24543,N_23171,N_23168);
or U24544 (N_24544,N_23586,N_23345);
and U24545 (N_24545,N_23458,N_23632);
nor U24546 (N_24546,N_23604,N_23337);
xnor U24547 (N_24547,N_23628,N_23690);
xor U24548 (N_24548,N_23325,N_23823);
xnor U24549 (N_24549,N_23391,N_23618);
or U24550 (N_24550,N_23087,N_23373);
xor U24551 (N_24551,N_23255,N_23402);
and U24552 (N_24552,N_23767,N_23636);
xnor U24553 (N_24553,N_23898,N_23002);
and U24554 (N_24554,N_23337,N_23777);
nor U24555 (N_24555,N_23719,N_23397);
or U24556 (N_24556,N_23561,N_23793);
and U24557 (N_24557,N_23235,N_23810);
nor U24558 (N_24558,N_23936,N_23063);
nand U24559 (N_24559,N_23020,N_23441);
and U24560 (N_24560,N_23920,N_23929);
nand U24561 (N_24561,N_23603,N_23530);
nand U24562 (N_24562,N_23027,N_23810);
or U24563 (N_24563,N_23754,N_23445);
nor U24564 (N_24564,N_23697,N_23328);
or U24565 (N_24565,N_23332,N_23792);
and U24566 (N_24566,N_23315,N_23489);
xor U24567 (N_24567,N_23984,N_23812);
nor U24568 (N_24568,N_23946,N_23836);
and U24569 (N_24569,N_23001,N_23632);
nand U24570 (N_24570,N_23539,N_23741);
xnor U24571 (N_24571,N_23636,N_23934);
or U24572 (N_24572,N_23648,N_23634);
or U24573 (N_24573,N_23393,N_23099);
nand U24574 (N_24574,N_23692,N_23882);
nand U24575 (N_24575,N_23289,N_23849);
or U24576 (N_24576,N_23206,N_23949);
xor U24577 (N_24577,N_23564,N_23164);
and U24578 (N_24578,N_23099,N_23816);
or U24579 (N_24579,N_23747,N_23175);
or U24580 (N_24580,N_23892,N_23252);
nor U24581 (N_24581,N_23630,N_23729);
xnor U24582 (N_24582,N_23578,N_23918);
or U24583 (N_24583,N_23929,N_23412);
xnor U24584 (N_24584,N_23955,N_23509);
or U24585 (N_24585,N_23674,N_23630);
xor U24586 (N_24586,N_23175,N_23793);
xor U24587 (N_24587,N_23581,N_23763);
nand U24588 (N_24588,N_23236,N_23279);
nor U24589 (N_24589,N_23271,N_23102);
xor U24590 (N_24590,N_23113,N_23456);
and U24591 (N_24591,N_23567,N_23310);
or U24592 (N_24592,N_23309,N_23690);
nand U24593 (N_24593,N_23067,N_23155);
and U24594 (N_24594,N_23131,N_23769);
or U24595 (N_24595,N_23018,N_23710);
nand U24596 (N_24596,N_23996,N_23563);
nand U24597 (N_24597,N_23701,N_23328);
xnor U24598 (N_24598,N_23022,N_23331);
and U24599 (N_24599,N_23623,N_23240);
xor U24600 (N_24600,N_23407,N_23727);
nor U24601 (N_24601,N_23363,N_23315);
xor U24602 (N_24602,N_23009,N_23821);
nor U24603 (N_24603,N_23410,N_23655);
nor U24604 (N_24604,N_23740,N_23824);
nor U24605 (N_24605,N_23113,N_23879);
or U24606 (N_24606,N_23960,N_23535);
nand U24607 (N_24607,N_23418,N_23825);
nand U24608 (N_24608,N_23515,N_23137);
nand U24609 (N_24609,N_23302,N_23227);
xnor U24610 (N_24610,N_23603,N_23487);
nor U24611 (N_24611,N_23897,N_23518);
or U24612 (N_24612,N_23873,N_23262);
nand U24613 (N_24613,N_23566,N_23719);
and U24614 (N_24614,N_23654,N_23160);
or U24615 (N_24615,N_23075,N_23560);
nor U24616 (N_24616,N_23524,N_23966);
or U24617 (N_24617,N_23095,N_23167);
or U24618 (N_24618,N_23209,N_23848);
nor U24619 (N_24619,N_23133,N_23205);
or U24620 (N_24620,N_23486,N_23848);
and U24621 (N_24621,N_23058,N_23060);
nor U24622 (N_24622,N_23487,N_23126);
nand U24623 (N_24623,N_23404,N_23071);
or U24624 (N_24624,N_23190,N_23140);
nand U24625 (N_24625,N_23797,N_23266);
nand U24626 (N_24626,N_23051,N_23375);
or U24627 (N_24627,N_23903,N_23589);
and U24628 (N_24628,N_23756,N_23533);
or U24629 (N_24629,N_23863,N_23320);
xnor U24630 (N_24630,N_23788,N_23820);
xor U24631 (N_24631,N_23962,N_23947);
nand U24632 (N_24632,N_23545,N_23588);
nor U24633 (N_24633,N_23886,N_23687);
and U24634 (N_24634,N_23782,N_23886);
or U24635 (N_24635,N_23866,N_23273);
nor U24636 (N_24636,N_23732,N_23213);
and U24637 (N_24637,N_23045,N_23966);
or U24638 (N_24638,N_23552,N_23825);
nand U24639 (N_24639,N_23000,N_23958);
and U24640 (N_24640,N_23011,N_23239);
or U24641 (N_24641,N_23571,N_23330);
xnor U24642 (N_24642,N_23322,N_23471);
or U24643 (N_24643,N_23088,N_23865);
xnor U24644 (N_24644,N_23714,N_23146);
and U24645 (N_24645,N_23495,N_23923);
xnor U24646 (N_24646,N_23881,N_23029);
nand U24647 (N_24647,N_23207,N_23168);
and U24648 (N_24648,N_23989,N_23138);
and U24649 (N_24649,N_23586,N_23305);
nor U24650 (N_24650,N_23230,N_23622);
nor U24651 (N_24651,N_23452,N_23765);
nand U24652 (N_24652,N_23777,N_23229);
nor U24653 (N_24653,N_23785,N_23299);
nand U24654 (N_24654,N_23680,N_23298);
nor U24655 (N_24655,N_23180,N_23105);
or U24656 (N_24656,N_23772,N_23733);
and U24657 (N_24657,N_23836,N_23603);
and U24658 (N_24658,N_23318,N_23276);
or U24659 (N_24659,N_23723,N_23411);
or U24660 (N_24660,N_23962,N_23770);
or U24661 (N_24661,N_23480,N_23831);
xor U24662 (N_24662,N_23684,N_23291);
nor U24663 (N_24663,N_23721,N_23885);
nand U24664 (N_24664,N_23158,N_23502);
and U24665 (N_24665,N_23277,N_23715);
and U24666 (N_24666,N_23223,N_23319);
nand U24667 (N_24667,N_23796,N_23951);
or U24668 (N_24668,N_23020,N_23555);
xnor U24669 (N_24669,N_23152,N_23079);
or U24670 (N_24670,N_23451,N_23939);
nand U24671 (N_24671,N_23300,N_23329);
nor U24672 (N_24672,N_23753,N_23953);
and U24673 (N_24673,N_23926,N_23295);
or U24674 (N_24674,N_23148,N_23441);
or U24675 (N_24675,N_23293,N_23066);
nand U24676 (N_24676,N_23667,N_23465);
and U24677 (N_24677,N_23901,N_23751);
xnor U24678 (N_24678,N_23488,N_23338);
nand U24679 (N_24679,N_23566,N_23578);
xor U24680 (N_24680,N_23085,N_23125);
or U24681 (N_24681,N_23156,N_23132);
nand U24682 (N_24682,N_23241,N_23927);
nand U24683 (N_24683,N_23062,N_23573);
or U24684 (N_24684,N_23064,N_23315);
and U24685 (N_24685,N_23319,N_23913);
nand U24686 (N_24686,N_23777,N_23608);
xnor U24687 (N_24687,N_23646,N_23982);
and U24688 (N_24688,N_23132,N_23036);
xor U24689 (N_24689,N_23067,N_23376);
nand U24690 (N_24690,N_23221,N_23583);
xnor U24691 (N_24691,N_23771,N_23164);
nor U24692 (N_24692,N_23782,N_23483);
and U24693 (N_24693,N_23942,N_23177);
xor U24694 (N_24694,N_23431,N_23960);
and U24695 (N_24695,N_23990,N_23263);
or U24696 (N_24696,N_23324,N_23147);
nor U24697 (N_24697,N_23336,N_23193);
xnor U24698 (N_24698,N_23291,N_23213);
or U24699 (N_24699,N_23509,N_23638);
xnor U24700 (N_24700,N_23449,N_23973);
nor U24701 (N_24701,N_23847,N_23073);
xor U24702 (N_24702,N_23729,N_23725);
xnor U24703 (N_24703,N_23670,N_23206);
and U24704 (N_24704,N_23806,N_23514);
or U24705 (N_24705,N_23332,N_23568);
xor U24706 (N_24706,N_23934,N_23207);
and U24707 (N_24707,N_23260,N_23557);
nand U24708 (N_24708,N_23003,N_23334);
or U24709 (N_24709,N_23127,N_23787);
or U24710 (N_24710,N_23907,N_23665);
nor U24711 (N_24711,N_23378,N_23855);
nor U24712 (N_24712,N_23997,N_23824);
nand U24713 (N_24713,N_23543,N_23045);
and U24714 (N_24714,N_23761,N_23068);
xor U24715 (N_24715,N_23467,N_23436);
xnor U24716 (N_24716,N_23013,N_23913);
nor U24717 (N_24717,N_23401,N_23688);
and U24718 (N_24718,N_23452,N_23136);
xor U24719 (N_24719,N_23086,N_23562);
xor U24720 (N_24720,N_23178,N_23947);
and U24721 (N_24721,N_23026,N_23395);
or U24722 (N_24722,N_23808,N_23964);
and U24723 (N_24723,N_23109,N_23773);
or U24724 (N_24724,N_23410,N_23827);
xnor U24725 (N_24725,N_23330,N_23893);
or U24726 (N_24726,N_23142,N_23911);
nor U24727 (N_24727,N_23104,N_23167);
or U24728 (N_24728,N_23368,N_23447);
xor U24729 (N_24729,N_23787,N_23719);
and U24730 (N_24730,N_23361,N_23671);
nand U24731 (N_24731,N_23960,N_23258);
and U24732 (N_24732,N_23228,N_23382);
nand U24733 (N_24733,N_23527,N_23072);
and U24734 (N_24734,N_23791,N_23679);
or U24735 (N_24735,N_23816,N_23681);
and U24736 (N_24736,N_23914,N_23046);
and U24737 (N_24737,N_23941,N_23134);
or U24738 (N_24738,N_23419,N_23929);
xnor U24739 (N_24739,N_23400,N_23071);
xor U24740 (N_24740,N_23372,N_23935);
and U24741 (N_24741,N_23431,N_23581);
or U24742 (N_24742,N_23659,N_23278);
nor U24743 (N_24743,N_23373,N_23431);
nand U24744 (N_24744,N_23726,N_23206);
nand U24745 (N_24745,N_23314,N_23559);
xor U24746 (N_24746,N_23728,N_23764);
xnor U24747 (N_24747,N_23267,N_23131);
xnor U24748 (N_24748,N_23020,N_23495);
nand U24749 (N_24749,N_23859,N_23820);
xor U24750 (N_24750,N_23110,N_23268);
nor U24751 (N_24751,N_23846,N_23254);
nor U24752 (N_24752,N_23319,N_23153);
or U24753 (N_24753,N_23033,N_23434);
nand U24754 (N_24754,N_23480,N_23093);
or U24755 (N_24755,N_23908,N_23706);
nor U24756 (N_24756,N_23490,N_23131);
or U24757 (N_24757,N_23455,N_23454);
nand U24758 (N_24758,N_23248,N_23074);
nor U24759 (N_24759,N_23794,N_23977);
and U24760 (N_24760,N_23532,N_23535);
or U24761 (N_24761,N_23738,N_23071);
or U24762 (N_24762,N_23597,N_23044);
and U24763 (N_24763,N_23525,N_23899);
and U24764 (N_24764,N_23982,N_23541);
and U24765 (N_24765,N_23293,N_23616);
or U24766 (N_24766,N_23898,N_23773);
nand U24767 (N_24767,N_23882,N_23864);
nor U24768 (N_24768,N_23486,N_23339);
nand U24769 (N_24769,N_23643,N_23891);
and U24770 (N_24770,N_23540,N_23543);
or U24771 (N_24771,N_23940,N_23742);
or U24772 (N_24772,N_23220,N_23888);
or U24773 (N_24773,N_23859,N_23959);
or U24774 (N_24774,N_23190,N_23971);
and U24775 (N_24775,N_23279,N_23072);
nand U24776 (N_24776,N_23854,N_23457);
xor U24777 (N_24777,N_23976,N_23880);
and U24778 (N_24778,N_23656,N_23074);
and U24779 (N_24779,N_23117,N_23159);
and U24780 (N_24780,N_23335,N_23924);
xnor U24781 (N_24781,N_23423,N_23757);
and U24782 (N_24782,N_23936,N_23881);
nand U24783 (N_24783,N_23418,N_23814);
or U24784 (N_24784,N_23389,N_23745);
and U24785 (N_24785,N_23579,N_23358);
nor U24786 (N_24786,N_23786,N_23951);
and U24787 (N_24787,N_23539,N_23973);
or U24788 (N_24788,N_23022,N_23753);
and U24789 (N_24789,N_23758,N_23475);
nor U24790 (N_24790,N_23908,N_23112);
xor U24791 (N_24791,N_23277,N_23383);
nand U24792 (N_24792,N_23440,N_23182);
or U24793 (N_24793,N_23891,N_23942);
nor U24794 (N_24794,N_23796,N_23996);
nor U24795 (N_24795,N_23591,N_23213);
xnor U24796 (N_24796,N_23747,N_23037);
xor U24797 (N_24797,N_23873,N_23040);
nor U24798 (N_24798,N_23988,N_23912);
nand U24799 (N_24799,N_23832,N_23097);
xnor U24800 (N_24800,N_23895,N_23257);
nor U24801 (N_24801,N_23313,N_23302);
xor U24802 (N_24802,N_23298,N_23069);
nand U24803 (N_24803,N_23379,N_23538);
xor U24804 (N_24804,N_23794,N_23169);
xnor U24805 (N_24805,N_23846,N_23722);
xnor U24806 (N_24806,N_23735,N_23057);
xor U24807 (N_24807,N_23905,N_23545);
xor U24808 (N_24808,N_23335,N_23879);
xnor U24809 (N_24809,N_23887,N_23219);
and U24810 (N_24810,N_23185,N_23404);
or U24811 (N_24811,N_23979,N_23806);
nand U24812 (N_24812,N_23544,N_23356);
nor U24813 (N_24813,N_23215,N_23385);
or U24814 (N_24814,N_23387,N_23103);
xor U24815 (N_24815,N_23392,N_23993);
nand U24816 (N_24816,N_23693,N_23530);
nor U24817 (N_24817,N_23502,N_23461);
nand U24818 (N_24818,N_23908,N_23341);
and U24819 (N_24819,N_23918,N_23540);
and U24820 (N_24820,N_23085,N_23953);
and U24821 (N_24821,N_23566,N_23322);
or U24822 (N_24822,N_23943,N_23247);
nand U24823 (N_24823,N_23091,N_23017);
nand U24824 (N_24824,N_23732,N_23508);
xnor U24825 (N_24825,N_23604,N_23676);
nor U24826 (N_24826,N_23129,N_23959);
xnor U24827 (N_24827,N_23913,N_23802);
and U24828 (N_24828,N_23411,N_23364);
nor U24829 (N_24829,N_23796,N_23922);
xnor U24830 (N_24830,N_23724,N_23839);
xor U24831 (N_24831,N_23509,N_23866);
and U24832 (N_24832,N_23588,N_23818);
nor U24833 (N_24833,N_23669,N_23681);
nor U24834 (N_24834,N_23841,N_23209);
nor U24835 (N_24835,N_23384,N_23078);
and U24836 (N_24836,N_23020,N_23189);
nand U24837 (N_24837,N_23851,N_23776);
xnor U24838 (N_24838,N_23779,N_23923);
or U24839 (N_24839,N_23625,N_23605);
nor U24840 (N_24840,N_23257,N_23161);
nor U24841 (N_24841,N_23706,N_23498);
nand U24842 (N_24842,N_23971,N_23735);
nand U24843 (N_24843,N_23278,N_23686);
nand U24844 (N_24844,N_23168,N_23724);
or U24845 (N_24845,N_23330,N_23795);
or U24846 (N_24846,N_23808,N_23973);
nand U24847 (N_24847,N_23408,N_23600);
nand U24848 (N_24848,N_23952,N_23037);
and U24849 (N_24849,N_23270,N_23422);
and U24850 (N_24850,N_23892,N_23654);
nor U24851 (N_24851,N_23930,N_23432);
and U24852 (N_24852,N_23373,N_23976);
nand U24853 (N_24853,N_23477,N_23280);
or U24854 (N_24854,N_23811,N_23968);
nand U24855 (N_24855,N_23439,N_23386);
and U24856 (N_24856,N_23850,N_23703);
nand U24857 (N_24857,N_23609,N_23181);
xor U24858 (N_24858,N_23537,N_23068);
and U24859 (N_24859,N_23749,N_23327);
xor U24860 (N_24860,N_23813,N_23605);
or U24861 (N_24861,N_23855,N_23390);
nor U24862 (N_24862,N_23752,N_23441);
or U24863 (N_24863,N_23095,N_23582);
nand U24864 (N_24864,N_23713,N_23046);
nand U24865 (N_24865,N_23603,N_23896);
xor U24866 (N_24866,N_23322,N_23692);
and U24867 (N_24867,N_23305,N_23966);
xor U24868 (N_24868,N_23547,N_23728);
or U24869 (N_24869,N_23624,N_23481);
nand U24870 (N_24870,N_23749,N_23635);
nand U24871 (N_24871,N_23598,N_23808);
nor U24872 (N_24872,N_23271,N_23606);
nor U24873 (N_24873,N_23006,N_23081);
xnor U24874 (N_24874,N_23951,N_23603);
and U24875 (N_24875,N_23282,N_23947);
nand U24876 (N_24876,N_23587,N_23979);
or U24877 (N_24877,N_23633,N_23129);
nor U24878 (N_24878,N_23632,N_23534);
xor U24879 (N_24879,N_23046,N_23737);
xor U24880 (N_24880,N_23940,N_23841);
nor U24881 (N_24881,N_23125,N_23166);
and U24882 (N_24882,N_23919,N_23239);
or U24883 (N_24883,N_23016,N_23598);
and U24884 (N_24884,N_23143,N_23163);
or U24885 (N_24885,N_23547,N_23981);
nor U24886 (N_24886,N_23116,N_23006);
nand U24887 (N_24887,N_23942,N_23605);
xor U24888 (N_24888,N_23189,N_23651);
or U24889 (N_24889,N_23568,N_23272);
and U24890 (N_24890,N_23047,N_23053);
nor U24891 (N_24891,N_23330,N_23537);
nand U24892 (N_24892,N_23156,N_23075);
xor U24893 (N_24893,N_23810,N_23510);
and U24894 (N_24894,N_23055,N_23257);
nor U24895 (N_24895,N_23176,N_23027);
nor U24896 (N_24896,N_23347,N_23053);
nand U24897 (N_24897,N_23101,N_23666);
xor U24898 (N_24898,N_23738,N_23101);
and U24899 (N_24899,N_23835,N_23886);
or U24900 (N_24900,N_23193,N_23222);
nor U24901 (N_24901,N_23850,N_23278);
nand U24902 (N_24902,N_23403,N_23314);
xor U24903 (N_24903,N_23241,N_23558);
nor U24904 (N_24904,N_23034,N_23347);
nand U24905 (N_24905,N_23584,N_23668);
or U24906 (N_24906,N_23281,N_23945);
or U24907 (N_24907,N_23498,N_23662);
nand U24908 (N_24908,N_23895,N_23153);
nor U24909 (N_24909,N_23655,N_23082);
xor U24910 (N_24910,N_23878,N_23663);
nand U24911 (N_24911,N_23608,N_23446);
nor U24912 (N_24912,N_23506,N_23786);
xnor U24913 (N_24913,N_23966,N_23265);
nand U24914 (N_24914,N_23398,N_23295);
and U24915 (N_24915,N_23804,N_23522);
and U24916 (N_24916,N_23291,N_23606);
and U24917 (N_24917,N_23045,N_23263);
xor U24918 (N_24918,N_23534,N_23598);
nand U24919 (N_24919,N_23182,N_23441);
and U24920 (N_24920,N_23373,N_23657);
and U24921 (N_24921,N_23591,N_23210);
nand U24922 (N_24922,N_23194,N_23227);
and U24923 (N_24923,N_23362,N_23368);
xnor U24924 (N_24924,N_23507,N_23961);
and U24925 (N_24925,N_23973,N_23454);
or U24926 (N_24926,N_23915,N_23709);
or U24927 (N_24927,N_23312,N_23112);
xnor U24928 (N_24928,N_23296,N_23754);
and U24929 (N_24929,N_23494,N_23320);
xnor U24930 (N_24930,N_23819,N_23653);
xor U24931 (N_24931,N_23169,N_23569);
nand U24932 (N_24932,N_23935,N_23272);
or U24933 (N_24933,N_23089,N_23861);
nand U24934 (N_24934,N_23033,N_23899);
nor U24935 (N_24935,N_23385,N_23597);
nand U24936 (N_24936,N_23438,N_23220);
nor U24937 (N_24937,N_23645,N_23083);
xor U24938 (N_24938,N_23243,N_23385);
nor U24939 (N_24939,N_23727,N_23966);
nor U24940 (N_24940,N_23603,N_23235);
nand U24941 (N_24941,N_23263,N_23156);
nor U24942 (N_24942,N_23663,N_23332);
and U24943 (N_24943,N_23151,N_23858);
nand U24944 (N_24944,N_23981,N_23576);
and U24945 (N_24945,N_23966,N_23956);
xor U24946 (N_24946,N_23421,N_23332);
and U24947 (N_24947,N_23200,N_23979);
xnor U24948 (N_24948,N_23779,N_23300);
nand U24949 (N_24949,N_23678,N_23448);
xnor U24950 (N_24950,N_23034,N_23568);
nand U24951 (N_24951,N_23771,N_23631);
nor U24952 (N_24952,N_23034,N_23848);
and U24953 (N_24953,N_23386,N_23628);
or U24954 (N_24954,N_23694,N_23586);
nand U24955 (N_24955,N_23710,N_23756);
nor U24956 (N_24956,N_23643,N_23310);
xor U24957 (N_24957,N_23225,N_23717);
nand U24958 (N_24958,N_23756,N_23085);
nand U24959 (N_24959,N_23513,N_23064);
and U24960 (N_24960,N_23866,N_23382);
xor U24961 (N_24961,N_23812,N_23493);
nor U24962 (N_24962,N_23308,N_23405);
nor U24963 (N_24963,N_23653,N_23502);
xor U24964 (N_24964,N_23357,N_23293);
nand U24965 (N_24965,N_23090,N_23757);
xor U24966 (N_24966,N_23050,N_23344);
and U24967 (N_24967,N_23791,N_23460);
xor U24968 (N_24968,N_23672,N_23175);
xor U24969 (N_24969,N_23434,N_23972);
or U24970 (N_24970,N_23786,N_23503);
xor U24971 (N_24971,N_23978,N_23349);
and U24972 (N_24972,N_23955,N_23843);
nand U24973 (N_24973,N_23983,N_23006);
and U24974 (N_24974,N_23901,N_23678);
nand U24975 (N_24975,N_23905,N_23504);
and U24976 (N_24976,N_23056,N_23428);
and U24977 (N_24977,N_23554,N_23219);
nand U24978 (N_24978,N_23797,N_23093);
and U24979 (N_24979,N_23474,N_23903);
nand U24980 (N_24980,N_23488,N_23317);
nand U24981 (N_24981,N_23906,N_23872);
xnor U24982 (N_24982,N_23491,N_23642);
nand U24983 (N_24983,N_23369,N_23256);
nor U24984 (N_24984,N_23143,N_23000);
or U24985 (N_24985,N_23256,N_23426);
nor U24986 (N_24986,N_23351,N_23975);
and U24987 (N_24987,N_23359,N_23218);
and U24988 (N_24988,N_23798,N_23245);
nor U24989 (N_24989,N_23620,N_23796);
xnor U24990 (N_24990,N_23950,N_23866);
and U24991 (N_24991,N_23187,N_23977);
nor U24992 (N_24992,N_23164,N_23623);
nor U24993 (N_24993,N_23388,N_23197);
nand U24994 (N_24994,N_23921,N_23207);
nand U24995 (N_24995,N_23611,N_23667);
nand U24996 (N_24996,N_23875,N_23956);
nor U24997 (N_24997,N_23250,N_23790);
nor U24998 (N_24998,N_23104,N_23291);
xor U24999 (N_24999,N_23953,N_23321);
and U25000 (N_25000,N_24540,N_24257);
xor U25001 (N_25001,N_24104,N_24439);
and U25002 (N_25002,N_24773,N_24967);
or U25003 (N_25003,N_24782,N_24736);
or U25004 (N_25004,N_24120,N_24381);
or U25005 (N_25005,N_24735,N_24207);
and U25006 (N_25006,N_24327,N_24486);
nand U25007 (N_25007,N_24793,N_24291);
or U25008 (N_25008,N_24930,N_24810);
nor U25009 (N_25009,N_24124,N_24901);
and U25010 (N_25010,N_24390,N_24923);
xnor U25011 (N_25011,N_24700,N_24081);
or U25012 (N_25012,N_24477,N_24572);
nor U25013 (N_25013,N_24666,N_24959);
nand U25014 (N_25014,N_24693,N_24647);
xor U25015 (N_25015,N_24558,N_24749);
nor U25016 (N_25016,N_24905,N_24117);
or U25017 (N_25017,N_24323,N_24788);
xor U25018 (N_25018,N_24529,N_24834);
or U25019 (N_25019,N_24660,N_24935);
and U25020 (N_25020,N_24239,N_24550);
nor U25021 (N_25021,N_24182,N_24944);
nor U25022 (N_25022,N_24803,N_24171);
and U25023 (N_25023,N_24546,N_24979);
and U25024 (N_25024,N_24850,N_24586);
and U25025 (N_25025,N_24204,N_24135);
and U25026 (N_25026,N_24873,N_24051);
and U25027 (N_25027,N_24436,N_24538);
or U25028 (N_25028,N_24630,N_24494);
nor U25029 (N_25029,N_24380,N_24136);
and U25030 (N_25030,N_24756,N_24157);
nor U25031 (N_25031,N_24802,N_24075);
or U25032 (N_25032,N_24837,N_24779);
and U25033 (N_25033,N_24328,N_24535);
nor U25034 (N_25034,N_24044,N_24234);
nand U25035 (N_25035,N_24928,N_24311);
nor U25036 (N_25036,N_24106,N_24615);
xnor U25037 (N_25037,N_24305,N_24791);
nor U25038 (N_25038,N_24007,N_24842);
or U25039 (N_25039,N_24116,N_24325);
nand U25040 (N_25040,N_24753,N_24441);
and U25041 (N_25041,N_24459,N_24038);
nor U25042 (N_25042,N_24225,N_24744);
nand U25043 (N_25043,N_24306,N_24512);
xnor U25044 (N_25044,N_24806,N_24021);
nand U25045 (N_25045,N_24835,N_24358);
nand U25046 (N_25046,N_24611,N_24169);
nand U25047 (N_25047,N_24228,N_24315);
xor U25048 (N_25048,N_24298,N_24409);
and U25049 (N_25049,N_24657,N_24478);
xor U25050 (N_25050,N_24539,N_24829);
nand U25051 (N_25051,N_24401,N_24078);
or U25052 (N_25052,N_24142,N_24922);
nor U25053 (N_25053,N_24556,N_24440);
xnor U25054 (N_25054,N_24527,N_24153);
nand U25055 (N_25055,N_24451,N_24145);
or U25056 (N_25056,N_24368,N_24200);
or U25057 (N_25057,N_24552,N_24988);
and U25058 (N_25058,N_24896,N_24815);
and U25059 (N_25059,N_24524,N_24033);
nand U25060 (N_25060,N_24448,N_24350);
xor U25061 (N_25061,N_24346,N_24956);
xnor U25062 (N_25062,N_24085,N_24613);
nand U25063 (N_25063,N_24721,N_24268);
nand U25064 (N_25064,N_24969,N_24816);
nor U25065 (N_25065,N_24692,N_24212);
nand U25066 (N_25066,N_24553,N_24671);
or U25067 (N_25067,N_24746,N_24367);
nor U25068 (N_25068,N_24783,N_24186);
or U25069 (N_25069,N_24121,N_24688);
xor U25070 (N_25070,N_24277,N_24899);
nand U25071 (N_25071,N_24673,N_24370);
xor U25072 (N_25072,N_24296,N_24581);
nor U25073 (N_25073,N_24464,N_24465);
xnor U25074 (N_25074,N_24644,N_24310);
xor U25075 (N_25075,N_24684,N_24826);
nor U25076 (N_25076,N_24592,N_24591);
and U25077 (N_25077,N_24545,N_24003);
nand U25078 (N_25078,N_24821,N_24322);
nand U25079 (N_25079,N_24397,N_24326);
nor U25080 (N_25080,N_24544,N_24187);
and U25081 (N_25081,N_24845,N_24993);
xor U25082 (N_25082,N_24992,N_24455);
nor U25083 (N_25083,N_24488,N_24208);
xor U25084 (N_25084,N_24415,N_24866);
xnor U25085 (N_25085,N_24391,N_24050);
nand U25086 (N_25086,N_24867,N_24340);
nor U25087 (N_25087,N_24167,N_24561);
nor U25088 (N_25088,N_24017,N_24522);
and U25089 (N_25089,N_24934,N_24795);
nand U25090 (N_25090,N_24881,N_24412);
xnor U25091 (N_25091,N_24520,N_24012);
nand U25092 (N_25092,N_24908,N_24787);
xor U25093 (N_25093,N_24047,N_24203);
and U25094 (N_25094,N_24205,N_24898);
nor U25095 (N_25095,N_24589,N_24070);
or U25096 (N_25096,N_24357,N_24991);
and U25097 (N_25097,N_24468,N_24600);
nor U25098 (N_25098,N_24906,N_24197);
and U25099 (N_25099,N_24710,N_24961);
and U25100 (N_25100,N_24472,N_24062);
or U25101 (N_25101,N_24109,N_24708);
xnor U25102 (N_25102,N_24879,N_24634);
nand U25103 (N_25103,N_24086,N_24606);
nor U25104 (N_25104,N_24264,N_24649);
and U25105 (N_25105,N_24139,N_24083);
xnor U25106 (N_25106,N_24292,N_24836);
nor U25107 (N_25107,N_24875,N_24759);
nand U25108 (N_25108,N_24669,N_24309);
and U25109 (N_25109,N_24609,N_24694);
xor U25110 (N_25110,N_24832,N_24536);
nand U25111 (N_25111,N_24662,N_24838);
nand U25112 (N_25112,N_24531,N_24450);
nor U25113 (N_25113,N_24579,N_24925);
nand U25114 (N_25114,N_24030,N_24608);
nand U25115 (N_25115,N_24717,N_24330);
xnor U25116 (N_25116,N_24607,N_24285);
nand U25117 (N_25117,N_24172,N_24011);
nand U25118 (N_25118,N_24105,N_24699);
or U25119 (N_25119,N_24764,N_24162);
or U25120 (N_25120,N_24218,N_24166);
and U25121 (N_25121,N_24254,N_24195);
nor U25122 (N_25122,N_24363,N_24823);
or U25123 (N_25123,N_24951,N_24920);
xnor U25124 (N_25124,N_24126,N_24943);
nor U25125 (N_25125,N_24261,N_24729);
or U25126 (N_25126,N_24960,N_24064);
nor U25127 (N_25127,N_24903,N_24314);
xor U25128 (N_25128,N_24937,N_24789);
and U25129 (N_25129,N_24331,N_24076);
and U25130 (N_25130,N_24774,N_24854);
nor U25131 (N_25131,N_24971,N_24256);
nor U25132 (N_25132,N_24022,N_24709);
or U25133 (N_25133,N_24933,N_24792);
or U25134 (N_25134,N_24929,N_24860);
nand U25135 (N_25135,N_24616,N_24469);
xor U25136 (N_25136,N_24491,N_24910);
xor U25137 (N_25137,N_24319,N_24580);
nand U25138 (N_25138,N_24237,N_24730);
and U25139 (N_25139,N_24131,N_24884);
or U25140 (N_25140,N_24278,N_24707);
xnor U25141 (N_25141,N_24683,N_24599);
and U25142 (N_25142,N_24054,N_24094);
nor U25143 (N_25143,N_24113,N_24772);
nor U25144 (N_25144,N_24247,N_24534);
nor U25145 (N_25145,N_24273,N_24295);
xor U25146 (N_25146,N_24794,N_24696);
nor U25147 (N_25147,N_24411,N_24290);
xor U25148 (N_25148,N_24159,N_24019);
or U25149 (N_25149,N_24165,N_24621);
nor U25150 (N_25150,N_24432,N_24697);
or U25151 (N_25151,N_24542,N_24986);
xor U25152 (N_25152,N_24214,N_24267);
and U25153 (N_25153,N_24084,N_24500);
and U25154 (N_25154,N_24185,N_24138);
nand U25155 (N_25155,N_24049,N_24229);
nand U25156 (N_25156,N_24698,N_24476);
nor U25157 (N_25157,N_24931,N_24423);
nor U25158 (N_25158,N_24701,N_24042);
and U25159 (N_25159,N_24874,N_24963);
or U25160 (N_25160,N_24945,N_24637);
and U25161 (N_25161,N_24110,N_24775);
or U25162 (N_25162,N_24897,N_24997);
nor U25163 (N_25163,N_24020,N_24828);
xnor U25164 (N_25164,N_24955,N_24382);
or U25165 (N_25165,N_24416,N_24217);
xor U25166 (N_25166,N_24888,N_24509);
nand U25167 (N_25167,N_24386,N_24479);
nand U25168 (N_25168,N_24577,N_24994);
nand U25169 (N_25169,N_24378,N_24324);
xnor U25170 (N_25170,N_24069,N_24886);
nor U25171 (N_25171,N_24525,N_24372);
xnor U25172 (N_25172,N_24046,N_24584);
xor U25173 (N_25173,N_24130,N_24058);
nand U25174 (N_25174,N_24023,N_24668);
or U25175 (N_25175,N_24487,N_24461);
xnor U25176 (N_25176,N_24495,N_24972);
xor U25177 (N_25177,N_24734,N_24576);
xnor U25178 (N_25178,N_24442,N_24804);
xnor U25179 (N_25179,N_24626,N_24618);
or U25180 (N_25180,N_24027,N_24807);
or U25181 (N_25181,N_24318,N_24950);
nand U25182 (N_25182,N_24780,N_24633);
or U25183 (N_25183,N_24303,N_24354);
nand U25184 (N_25184,N_24154,N_24199);
xor U25185 (N_25185,N_24489,N_24163);
nand U25186 (N_25186,N_24446,N_24080);
nand U25187 (N_25187,N_24031,N_24808);
and U25188 (N_25188,N_24739,N_24505);
xor U25189 (N_25189,N_24151,N_24192);
xor U25190 (N_25190,N_24987,N_24258);
nor U25191 (N_25191,N_24176,N_24393);
or U25192 (N_25192,N_24429,N_24691);
or U25193 (N_25193,N_24682,N_24024);
xor U25194 (N_25194,N_24443,N_24371);
and U25195 (N_25195,N_24438,N_24048);
nor U25196 (N_25196,N_24175,N_24034);
or U25197 (N_25197,N_24851,N_24376);
nand U25198 (N_25198,N_24082,N_24052);
nand U25199 (N_25199,N_24067,N_24173);
nand U25200 (N_25200,N_24039,N_24653);
xor U25201 (N_25201,N_24307,N_24032);
nor U25202 (N_25202,N_24010,N_24876);
nor U25203 (N_25203,N_24210,N_24118);
and U25204 (N_25204,N_24623,N_24015);
nor U25205 (N_25205,N_24585,N_24918);
and U25206 (N_25206,N_24975,N_24818);
nand U25207 (N_25207,N_24720,N_24578);
nor U25208 (N_25208,N_24868,N_24410);
nor U25209 (N_25209,N_24639,N_24865);
nand U25210 (N_25210,N_24748,N_24335);
and U25211 (N_25211,N_24344,N_24652);
or U25212 (N_25212,N_24885,N_24504);
or U25213 (N_25213,N_24170,N_24341);
xor U25214 (N_25214,N_24638,N_24762);
xnor U25215 (N_25215,N_24902,N_24374);
or U25216 (N_25216,N_24356,N_24732);
xor U25217 (N_25217,N_24066,N_24947);
nand U25218 (N_25218,N_24800,N_24702);
or U25219 (N_25219,N_24388,N_24541);
nand U25220 (N_25220,N_24687,N_24796);
or U25221 (N_25221,N_24308,N_24904);
or U25222 (N_25222,N_24279,N_24202);
and U25223 (N_25223,N_24213,N_24907);
nor U25224 (N_25224,N_24765,N_24651);
or U25225 (N_25225,N_24663,N_24559);
or U25226 (N_25226,N_24492,N_24911);
and U25227 (N_25227,N_24364,N_24394);
and U25228 (N_25228,N_24565,N_24650);
nor U25229 (N_25229,N_24516,N_24568);
nand U25230 (N_25230,N_24063,N_24714);
or U25231 (N_25231,N_24098,N_24751);
xor U25232 (N_25232,N_24127,N_24026);
and U25233 (N_25233,N_24685,N_24777);
nand U25234 (N_25234,N_24570,N_24016);
nand U25235 (N_25235,N_24575,N_24601);
nand U25236 (N_25236,N_24705,N_24270);
and U25237 (N_25237,N_24824,N_24255);
nor U25238 (N_25238,N_24071,N_24724);
xor U25239 (N_25239,N_24675,N_24402);
nand U25240 (N_25240,N_24119,N_24799);
and U25241 (N_25241,N_24502,N_24990);
nor U25242 (N_25242,N_24594,N_24260);
xnor U25243 (N_25243,N_24619,N_24089);
xnor U25244 (N_25244,N_24862,N_24164);
xor U25245 (N_25245,N_24593,N_24434);
xnor U25246 (N_25246,N_24574,N_24345);
xor U25247 (N_25247,N_24392,N_24786);
nand U25248 (N_25248,N_24526,N_24598);
nor U25249 (N_25249,N_24863,N_24820);
xnor U25250 (N_25250,N_24661,N_24413);
xnor U25251 (N_25251,N_24848,N_24280);
or U25252 (N_25252,N_24916,N_24706);
nand U25253 (N_25253,N_24877,N_24968);
or U25254 (N_25254,N_24554,N_24758);
nand U25255 (N_25255,N_24755,N_24395);
xnor U25256 (N_25256,N_24266,N_24014);
nor U25257 (N_25257,N_24499,N_24373);
and U25258 (N_25258,N_24506,N_24833);
xnor U25259 (N_25259,N_24814,N_24895);
or U25260 (N_25260,N_24425,N_24747);
nor U25261 (N_25261,N_24405,N_24056);
xor U25262 (N_25262,N_24533,N_24900);
nand U25263 (N_25263,N_24317,N_24114);
xnor U25264 (N_25264,N_24767,N_24811);
and U25265 (N_25265,N_24343,N_24595);
and U25266 (N_25266,N_24471,N_24548);
and U25267 (N_25267,N_24407,N_24603);
or U25268 (N_25268,N_24635,N_24355);
xor U25269 (N_25269,N_24913,N_24801);
nor U25270 (N_25270,N_24713,N_24271);
xnor U25271 (N_25271,N_24060,N_24417);
and U25272 (N_25272,N_24179,N_24099);
and U25273 (N_25273,N_24422,N_24115);
xor U25274 (N_25274,N_24158,N_24909);
and U25275 (N_25275,N_24057,N_24236);
xnor U25276 (N_25276,N_24846,N_24617);
xnor U25277 (N_25277,N_24244,N_24333);
nand U25278 (N_25278,N_24511,N_24293);
xnor U25279 (N_25279,N_24133,N_24191);
and U25280 (N_25280,N_24625,N_24629);
or U25281 (N_25281,N_24738,N_24072);
or U25282 (N_25282,N_24286,N_24265);
nand U25283 (N_25283,N_24396,N_24223);
or U25284 (N_25284,N_24695,N_24513);
xor U25285 (N_25285,N_24242,N_24462);
nor U25286 (N_25286,N_24948,N_24564);
and U25287 (N_25287,N_24596,N_24435);
xor U25288 (N_25288,N_24125,N_24137);
xnor U25289 (N_25289,N_24112,N_24641);
nor U25290 (N_25290,N_24320,N_24065);
and U25291 (N_25291,N_24983,N_24831);
xor U25292 (N_25292,N_24359,N_24250);
and U25293 (N_25293,N_24674,N_24861);
nor U25294 (N_25294,N_24883,N_24129);
and U25295 (N_25295,N_24398,N_24002);
or U25296 (N_25296,N_24924,N_24146);
or U25297 (N_25297,N_24628,N_24059);
xnor U25298 (N_25298,N_24768,N_24272);
nor U25299 (N_25299,N_24299,N_24349);
nand U25300 (N_25300,N_24149,N_24103);
or U25301 (N_25301,N_24101,N_24369);
nand U25302 (N_25302,N_24013,N_24073);
and U25303 (N_25303,N_24893,N_24406);
nand U25304 (N_25304,N_24915,N_24233);
and U25305 (N_25305,N_24177,N_24111);
and U25306 (N_25306,N_24754,N_24160);
nand U25307 (N_25307,N_24532,N_24074);
and U25308 (N_25308,N_24090,N_24745);
and U25309 (N_25309,N_24521,N_24573);
and U25310 (N_25310,N_24858,N_24238);
nand U25311 (N_25311,N_24679,N_24812);
nor U25312 (N_25312,N_24178,N_24703);
nor U25313 (N_25313,N_24232,N_24152);
and U25314 (N_25314,N_24981,N_24283);
or U25315 (N_25315,N_24362,N_24055);
xor U25316 (N_25316,N_24087,N_24555);
and U25317 (N_25317,N_24891,N_24966);
and U25318 (N_25318,N_24453,N_24181);
nor U25319 (N_25319,N_24813,N_24817);
xor U25320 (N_25320,N_24672,N_24560);
xor U25321 (N_25321,N_24156,N_24953);
nand U25322 (N_25322,N_24632,N_24365);
xnor U25323 (N_25323,N_24235,N_24590);
and U25324 (N_25324,N_24543,N_24107);
xor U25325 (N_25325,N_24664,N_24843);
nor U25326 (N_25326,N_24704,N_24518);
and U25327 (N_25327,N_24686,N_24562);
nor U25328 (N_25328,N_24061,N_24092);
and U25329 (N_25329,N_24750,N_24760);
nand U25330 (N_25330,N_24778,N_24088);
or U25331 (N_25331,N_24294,N_24211);
or U25332 (N_25332,N_24939,N_24917);
and U25333 (N_25333,N_24096,N_24690);
or U25334 (N_25334,N_24769,N_24827);
nand U25335 (N_25335,N_24996,N_24977);
and U25336 (N_25336,N_24419,N_24612);
nor U25337 (N_25337,N_24770,N_24482);
nand U25338 (N_25338,N_24313,N_24077);
or U25339 (N_25339,N_24712,N_24849);
nor U25340 (N_25340,N_24856,N_24781);
and U25341 (N_25341,N_24245,N_24643);
nand U25342 (N_25342,N_24517,N_24045);
or U25343 (N_25343,N_24936,N_24946);
or U25344 (N_25344,N_24467,N_24337);
and U25345 (N_25345,N_24602,N_24711);
nand U25346 (N_25346,N_24029,N_24740);
or U25347 (N_25347,N_24426,N_24507);
nand U25348 (N_25348,N_24825,N_24196);
nor U25349 (N_25349,N_24230,N_24215);
nor U25350 (N_25350,N_24722,N_24454);
xor U25351 (N_25351,N_24147,N_24183);
nand U25352 (N_25352,N_24882,N_24338);
or U25353 (N_25353,N_24670,N_24274);
nor U25354 (N_25354,N_24557,N_24890);
xor U25355 (N_25355,N_24190,N_24880);
xor U25356 (N_25356,N_24927,N_24384);
nand U25357 (N_25357,N_24352,N_24892);
and U25358 (N_25358,N_24474,N_24155);
xnor U25359 (N_25359,N_24610,N_24537);
or U25360 (N_25360,N_24004,N_24300);
nand U25361 (N_25361,N_24725,N_24716);
nand U25362 (N_25362,N_24231,N_24853);
nand U25363 (N_25363,N_24731,N_24418);
and U25364 (N_25364,N_24025,N_24473);
nor U25365 (N_25365,N_24414,N_24962);
or U25366 (N_25366,N_24188,N_24408);
xnor U25367 (N_25367,N_24456,N_24132);
xnor U25368 (N_25368,N_24001,N_24859);
or U25369 (N_25369,N_24091,N_24437);
nor U25370 (N_25370,N_24457,N_24246);
and U25371 (N_25371,N_24949,N_24912);
or U25372 (N_25372,N_24387,N_24588);
xor U25373 (N_25373,N_24503,N_24184);
or U25374 (N_25374,N_24941,N_24470);
xor U25375 (N_25375,N_24515,N_24134);
and U25376 (N_25376,N_24965,N_24297);
and U25377 (N_25377,N_24715,N_24389);
xor U25378 (N_25378,N_24102,N_24351);
or U25379 (N_25379,N_24312,N_24678);
or U25380 (N_25380,N_24219,N_24144);
nand U25381 (N_25381,N_24932,N_24805);
nor U25382 (N_25382,N_24424,N_24743);
or U25383 (N_25383,N_24719,N_24222);
or U25384 (N_25384,N_24510,N_24493);
nor U25385 (N_25385,N_24128,N_24742);
or U25386 (N_25386,N_24347,N_24490);
nand U25387 (N_25387,N_24501,N_24940);
nand U25388 (N_25388,N_24321,N_24206);
xnor U25389 (N_25389,N_24276,N_24403);
or U25390 (N_25390,N_24844,N_24035);
xnor U25391 (N_25391,N_24248,N_24399);
or U25392 (N_25392,N_24645,N_24984);
xnor U25393 (N_25393,N_24658,N_24037);
and U25394 (N_25394,N_24444,N_24226);
and U25395 (N_25395,N_24974,N_24938);
or U25396 (N_25396,N_24872,N_24995);
nor U25397 (N_25397,N_24809,N_24161);
and U25398 (N_25398,N_24921,N_24243);
and U25399 (N_25399,N_24269,N_24108);
or U25400 (N_25400,N_24819,N_24659);
nor U25401 (N_25401,N_24018,N_24334);
nor U25402 (N_25402,N_24463,N_24665);
or U25403 (N_25403,N_24342,N_24361);
nor U25404 (N_25404,N_24209,N_24053);
and U25405 (N_25405,N_24894,N_24180);
nand U25406 (N_25406,N_24980,N_24201);
xnor U25407 (N_25407,N_24360,N_24332);
or U25408 (N_25408,N_24733,N_24249);
nor U25409 (N_25409,N_24919,N_24251);
and U25410 (N_25410,N_24514,N_24123);
nor U25411 (N_25411,N_24563,N_24449);
nand U25412 (N_25412,N_24785,N_24302);
or U25413 (N_25413,N_24718,N_24431);
xnor U25414 (N_25414,N_24379,N_24336);
nand U25415 (N_25415,N_24329,N_24766);
nand U25416 (N_25416,N_24587,N_24957);
nor U25417 (N_25417,N_24648,N_24433);
nor U25418 (N_25418,N_24847,N_24627);
or U25419 (N_25419,N_24677,N_24954);
xnor U25420 (N_25420,N_24631,N_24241);
nor U25421 (N_25421,N_24339,N_24040);
xnor U25422 (N_25422,N_24227,N_24871);
or U25423 (N_25423,N_24976,N_24989);
nor U25424 (N_25424,N_24452,N_24041);
and U25425 (N_25425,N_24275,N_24008);
and U25426 (N_25426,N_24485,N_24043);
nor U25427 (N_25427,N_24150,N_24840);
and U25428 (N_25428,N_24421,N_24519);
nand U25429 (N_25429,N_24569,N_24097);
and U25430 (N_25430,N_24189,N_24723);
nand U25431 (N_25431,N_24385,N_24353);
and U25432 (N_25432,N_24009,N_24667);
and U25433 (N_25433,N_24252,N_24839);
nor U25434 (N_25434,N_24727,N_24240);
or U25435 (N_25435,N_24737,N_24262);
nand U25436 (N_25436,N_24484,N_24728);
nand U25437 (N_25437,N_24301,N_24752);
or U25438 (N_25438,N_24926,N_24497);
or U25439 (N_25439,N_24460,N_24857);
xnor U25440 (N_25440,N_24224,N_24889);
and U25441 (N_25441,N_24642,N_24428);
and U25442 (N_25442,N_24680,N_24289);
nand U25443 (N_25443,N_24466,N_24597);
nor U25444 (N_25444,N_24348,N_24583);
xnor U25445 (N_25445,N_24761,N_24952);
and U25446 (N_25446,N_24654,N_24475);
or U25447 (N_25447,N_24726,N_24614);
nand U25448 (N_25448,N_24168,N_24776);
nand U25449 (N_25449,N_24604,N_24304);
or U25450 (N_25450,N_24194,N_24458);
nor U25451 (N_25451,N_24140,N_24481);
nor U25452 (N_25452,N_24483,N_24771);
and U25453 (N_25453,N_24624,N_24143);
nand U25454 (N_25454,N_24622,N_24068);
nor U25455 (N_25455,N_24790,N_24741);
or U25456 (N_25456,N_24571,N_24079);
and U25457 (N_25457,N_24420,N_24445);
xnor U25458 (N_25458,N_24122,N_24549);
nand U25459 (N_25459,N_24582,N_24377);
nand U25460 (N_25460,N_24383,N_24528);
and U25461 (N_25461,N_24498,N_24028);
nand U25462 (N_25462,N_24427,N_24978);
nand U25463 (N_25463,N_24964,N_24655);
nor U25464 (N_25464,N_24852,N_24404);
and U25465 (N_25465,N_24447,N_24830);
xnor U25466 (N_25466,N_24193,N_24620);
and U25467 (N_25467,N_24982,N_24366);
or U25468 (N_25468,N_24640,N_24095);
nor U25469 (N_25469,N_24676,N_24006);
nand U25470 (N_25470,N_24797,N_24220);
or U25471 (N_25471,N_24822,N_24855);
nor U25472 (N_25472,N_24887,N_24656);
and U25473 (N_25473,N_24681,N_24281);
nor U25474 (N_25474,N_24985,N_24970);
xor U25475 (N_25475,N_24174,N_24496);
nand U25476 (N_25476,N_24005,N_24869);
nor U25477 (N_25477,N_24998,N_24316);
and U25478 (N_25478,N_24757,N_24689);
xor U25479 (N_25479,N_24284,N_24198);
nor U25480 (N_25480,N_24841,N_24636);
or U25481 (N_25481,N_24942,N_24973);
and U25482 (N_25482,N_24878,N_24263);
nand U25483 (N_25483,N_24282,N_24000);
nor U25484 (N_25484,N_24508,N_24523);
and U25485 (N_25485,N_24551,N_24288);
nand U25486 (N_25486,N_24914,N_24530);
xnor U25487 (N_25487,N_24605,N_24547);
nor U25488 (N_25488,N_24141,N_24566);
and U25489 (N_25489,N_24430,N_24100);
and U25490 (N_25490,N_24036,N_24216);
or U25491 (N_25491,N_24480,N_24646);
xnor U25492 (N_25492,N_24400,N_24221);
or U25493 (N_25493,N_24784,N_24567);
and U25494 (N_25494,N_24864,N_24798);
or U25495 (N_25495,N_24763,N_24870);
or U25496 (N_25496,N_24999,N_24375);
or U25497 (N_25497,N_24148,N_24287);
or U25498 (N_25498,N_24253,N_24093);
nand U25499 (N_25499,N_24259,N_24958);
or U25500 (N_25500,N_24821,N_24939);
or U25501 (N_25501,N_24631,N_24617);
nor U25502 (N_25502,N_24553,N_24403);
xor U25503 (N_25503,N_24754,N_24335);
nor U25504 (N_25504,N_24357,N_24691);
nand U25505 (N_25505,N_24790,N_24570);
nor U25506 (N_25506,N_24400,N_24701);
or U25507 (N_25507,N_24502,N_24935);
nand U25508 (N_25508,N_24503,N_24449);
or U25509 (N_25509,N_24425,N_24769);
xnor U25510 (N_25510,N_24803,N_24174);
nand U25511 (N_25511,N_24600,N_24700);
nand U25512 (N_25512,N_24808,N_24587);
and U25513 (N_25513,N_24390,N_24479);
or U25514 (N_25514,N_24603,N_24606);
or U25515 (N_25515,N_24245,N_24779);
nor U25516 (N_25516,N_24497,N_24554);
nand U25517 (N_25517,N_24929,N_24752);
nor U25518 (N_25518,N_24284,N_24329);
nand U25519 (N_25519,N_24119,N_24514);
and U25520 (N_25520,N_24328,N_24989);
or U25521 (N_25521,N_24801,N_24677);
nand U25522 (N_25522,N_24745,N_24270);
nor U25523 (N_25523,N_24904,N_24187);
or U25524 (N_25524,N_24925,N_24948);
or U25525 (N_25525,N_24345,N_24484);
nor U25526 (N_25526,N_24251,N_24323);
nand U25527 (N_25527,N_24703,N_24066);
xnor U25528 (N_25528,N_24314,N_24797);
nor U25529 (N_25529,N_24300,N_24339);
xor U25530 (N_25530,N_24744,N_24596);
nor U25531 (N_25531,N_24553,N_24857);
or U25532 (N_25532,N_24275,N_24215);
or U25533 (N_25533,N_24573,N_24086);
nor U25534 (N_25534,N_24208,N_24708);
or U25535 (N_25535,N_24369,N_24284);
and U25536 (N_25536,N_24647,N_24464);
nand U25537 (N_25537,N_24636,N_24237);
or U25538 (N_25538,N_24134,N_24341);
nor U25539 (N_25539,N_24092,N_24362);
nand U25540 (N_25540,N_24190,N_24652);
nand U25541 (N_25541,N_24649,N_24816);
and U25542 (N_25542,N_24410,N_24673);
and U25543 (N_25543,N_24497,N_24930);
nor U25544 (N_25544,N_24833,N_24805);
and U25545 (N_25545,N_24009,N_24989);
nor U25546 (N_25546,N_24226,N_24150);
xnor U25547 (N_25547,N_24598,N_24646);
or U25548 (N_25548,N_24748,N_24732);
nor U25549 (N_25549,N_24663,N_24050);
nand U25550 (N_25550,N_24350,N_24177);
nor U25551 (N_25551,N_24896,N_24860);
or U25552 (N_25552,N_24629,N_24566);
or U25553 (N_25553,N_24039,N_24975);
nor U25554 (N_25554,N_24771,N_24590);
nand U25555 (N_25555,N_24868,N_24186);
xor U25556 (N_25556,N_24287,N_24789);
nand U25557 (N_25557,N_24553,N_24386);
xnor U25558 (N_25558,N_24213,N_24817);
or U25559 (N_25559,N_24899,N_24357);
and U25560 (N_25560,N_24524,N_24496);
nor U25561 (N_25561,N_24297,N_24726);
and U25562 (N_25562,N_24006,N_24219);
or U25563 (N_25563,N_24349,N_24033);
and U25564 (N_25564,N_24450,N_24497);
xnor U25565 (N_25565,N_24277,N_24688);
nand U25566 (N_25566,N_24868,N_24510);
and U25567 (N_25567,N_24345,N_24314);
nand U25568 (N_25568,N_24991,N_24554);
and U25569 (N_25569,N_24171,N_24614);
xnor U25570 (N_25570,N_24240,N_24229);
nand U25571 (N_25571,N_24691,N_24976);
or U25572 (N_25572,N_24778,N_24196);
nor U25573 (N_25573,N_24618,N_24004);
and U25574 (N_25574,N_24089,N_24691);
xor U25575 (N_25575,N_24028,N_24221);
and U25576 (N_25576,N_24802,N_24549);
and U25577 (N_25577,N_24563,N_24015);
and U25578 (N_25578,N_24292,N_24879);
nand U25579 (N_25579,N_24506,N_24181);
nor U25580 (N_25580,N_24280,N_24943);
or U25581 (N_25581,N_24648,N_24153);
and U25582 (N_25582,N_24061,N_24010);
nand U25583 (N_25583,N_24495,N_24935);
xor U25584 (N_25584,N_24425,N_24202);
nand U25585 (N_25585,N_24191,N_24079);
or U25586 (N_25586,N_24098,N_24070);
or U25587 (N_25587,N_24372,N_24423);
xnor U25588 (N_25588,N_24239,N_24606);
nand U25589 (N_25589,N_24919,N_24785);
or U25590 (N_25590,N_24968,N_24564);
nand U25591 (N_25591,N_24722,N_24422);
xor U25592 (N_25592,N_24499,N_24076);
or U25593 (N_25593,N_24800,N_24301);
nor U25594 (N_25594,N_24763,N_24630);
nor U25595 (N_25595,N_24359,N_24227);
and U25596 (N_25596,N_24648,N_24476);
nand U25597 (N_25597,N_24505,N_24878);
or U25598 (N_25598,N_24062,N_24486);
and U25599 (N_25599,N_24174,N_24316);
nand U25600 (N_25600,N_24224,N_24308);
or U25601 (N_25601,N_24195,N_24141);
nor U25602 (N_25602,N_24881,N_24345);
or U25603 (N_25603,N_24533,N_24604);
or U25604 (N_25604,N_24458,N_24218);
and U25605 (N_25605,N_24017,N_24657);
or U25606 (N_25606,N_24727,N_24572);
nor U25607 (N_25607,N_24240,N_24246);
nor U25608 (N_25608,N_24621,N_24672);
nand U25609 (N_25609,N_24681,N_24860);
or U25610 (N_25610,N_24514,N_24380);
nor U25611 (N_25611,N_24468,N_24745);
and U25612 (N_25612,N_24931,N_24863);
and U25613 (N_25613,N_24415,N_24875);
xnor U25614 (N_25614,N_24018,N_24172);
xor U25615 (N_25615,N_24574,N_24177);
and U25616 (N_25616,N_24863,N_24043);
and U25617 (N_25617,N_24594,N_24024);
nor U25618 (N_25618,N_24961,N_24117);
and U25619 (N_25619,N_24452,N_24000);
nor U25620 (N_25620,N_24054,N_24460);
nor U25621 (N_25621,N_24958,N_24922);
nor U25622 (N_25622,N_24392,N_24483);
xor U25623 (N_25623,N_24482,N_24693);
and U25624 (N_25624,N_24638,N_24753);
nor U25625 (N_25625,N_24951,N_24761);
xnor U25626 (N_25626,N_24176,N_24792);
and U25627 (N_25627,N_24338,N_24012);
nor U25628 (N_25628,N_24624,N_24376);
and U25629 (N_25629,N_24402,N_24624);
nor U25630 (N_25630,N_24077,N_24163);
nor U25631 (N_25631,N_24195,N_24202);
nand U25632 (N_25632,N_24789,N_24912);
or U25633 (N_25633,N_24405,N_24857);
and U25634 (N_25634,N_24380,N_24693);
nor U25635 (N_25635,N_24521,N_24930);
nor U25636 (N_25636,N_24273,N_24588);
and U25637 (N_25637,N_24696,N_24564);
and U25638 (N_25638,N_24318,N_24396);
and U25639 (N_25639,N_24738,N_24180);
xor U25640 (N_25640,N_24757,N_24439);
xor U25641 (N_25641,N_24190,N_24031);
nor U25642 (N_25642,N_24697,N_24796);
or U25643 (N_25643,N_24856,N_24545);
and U25644 (N_25644,N_24414,N_24247);
or U25645 (N_25645,N_24387,N_24927);
nor U25646 (N_25646,N_24912,N_24155);
nand U25647 (N_25647,N_24137,N_24080);
or U25648 (N_25648,N_24175,N_24255);
nor U25649 (N_25649,N_24286,N_24346);
xnor U25650 (N_25650,N_24392,N_24578);
nor U25651 (N_25651,N_24960,N_24331);
nand U25652 (N_25652,N_24044,N_24616);
nor U25653 (N_25653,N_24766,N_24690);
nor U25654 (N_25654,N_24982,N_24760);
nor U25655 (N_25655,N_24563,N_24623);
nor U25656 (N_25656,N_24860,N_24288);
or U25657 (N_25657,N_24692,N_24898);
xnor U25658 (N_25658,N_24856,N_24454);
xnor U25659 (N_25659,N_24766,N_24217);
or U25660 (N_25660,N_24272,N_24560);
nand U25661 (N_25661,N_24882,N_24217);
xnor U25662 (N_25662,N_24231,N_24263);
nand U25663 (N_25663,N_24538,N_24349);
nor U25664 (N_25664,N_24131,N_24427);
and U25665 (N_25665,N_24008,N_24070);
xnor U25666 (N_25666,N_24495,N_24985);
or U25667 (N_25667,N_24668,N_24993);
or U25668 (N_25668,N_24254,N_24489);
and U25669 (N_25669,N_24389,N_24544);
nand U25670 (N_25670,N_24580,N_24290);
nor U25671 (N_25671,N_24126,N_24340);
and U25672 (N_25672,N_24207,N_24077);
or U25673 (N_25673,N_24396,N_24872);
and U25674 (N_25674,N_24367,N_24323);
and U25675 (N_25675,N_24201,N_24296);
nand U25676 (N_25676,N_24029,N_24463);
nand U25677 (N_25677,N_24140,N_24499);
and U25678 (N_25678,N_24893,N_24508);
or U25679 (N_25679,N_24723,N_24345);
or U25680 (N_25680,N_24951,N_24420);
xnor U25681 (N_25681,N_24429,N_24572);
or U25682 (N_25682,N_24958,N_24280);
and U25683 (N_25683,N_24165,N_24779);
or U25684 (N_25684,N_24737,N_24980);
nand U25685 (N_25685,N_24923,N_24222);
or U25686 (N_25686,N_24350,N_24757);
nor U25687 (N_25687,N_24097,N_24021);
nor U25688 (N_25688,N_24467,N_24351);
nand U25689 (N_25689,N_24150,N_24582);
xor U25690 (N_25690,N_24689,N_24075);
nor U25691 (N_25691,N_24171,N_24834);
or U25692 (N_25692,N_24441,N_24344);
and U25693 (N_25693,N_24171,N_24814);
nand U25694 (N_25694,N_24927,N_24684);
nand U25695 (N_25695,N_24696,N_24362);
or U25696 (N_25696,N_24570,N_24030);
and U25697 (N_25697,N_24472,N_24605);
or U25698 (N_25698,N_24535,N_24069);
or U25699 (N_25699,N_24951,N_24727);
and U25700 (N_25700,N_24411,N_24862);
xor U25701 (N_25701,N_24401,N_24654);
nor U25702 (N_25702,N_24147,N_24273);
nand U25703 (N_25703,N_24477,N_24472);
or U25704 (N_25704,N_24602,N_24687);
and U25705 (N_25705,N_24551,N_24100);
and U25706 (N_25706,N_24567,N_24014);
or U25707 (N_25707,N_24980,N_24702);
or U25708 (N_25708,N_24771,N_24835);
nor U25709 (N_25709,N_24703,N_24333);
nand U25710 (N_25710,N_24383,N_24391);
nor U25711 (N_25711,N_24508,N_24211);
and U25712 (N_25712,N_24708,N_24879);
nand U25713 (N_25713,N_24140,N_24227);
or U25714 (N_25714,N_24553,N_24865);
nor U25715 (N_25715,N_24652,N_24297);
nand U25716 (N_25716,N_24736,N_24988);
xor U25717 (N_25717,N_24390,N_24223);
nor U25718 (N_25718,N_24931,N_24606);
or U25719 (N_25719,N_24477,N_24895);
or U25720 (N_25720,N_24925,N_24331);
nand U25721 (N_25721,N_24915,N_24949);
nor U25722 (N_25722,N_24306,N_24076);
nor U25723 (N_25723,N_24739,N_24257);
and U25724 (N_25724,N_24337,N_24763);
and U25725 (N_25725,N_24635,N_24653);
nor U25726 (N_25726,N_24466,N_24464);
nand U25727 (N_25727,N_24738,N_24759);
and U25728 (N_25728,N_24388,N_24180);
xnor U25729 (N_25729,N_24826,N_24490);
nand U25730 (N_25730,N_24508,N_24888);
nor U25731 (N_25731,N_24616,N_24617);
xor U25732 (N_25732,N_24901,N_24973);
xor U25733 (N_25733,N_24182,N_24090);
nand U25734 (N_25734,N_24600,N_24147);
and U25735 (N_25735,N_24479,N_24275);
nor U25736 (N_25736,N_24026,N_24083);
or U25737 (N_25737,N_24709,N_24145);
nor U25738 (N_25738,N_24210,N_24649);
nand U25739 (N_25739,N_24400,N_24795);
or U25740 (N_25740,N_24887,N_24250);
nor U25741 (N_25741,N_24224,N_24946);
or U25742 (N_25742,N_24959,N_24800);
xor U25743 (N_25743,N_24855,N_24427);
or U25744 (N_25744,N_24467,N_24842);
nand U25745 (N_25745,N_24367,N_24392);
xor U25746 (N_25746,N_24296,N_24978);
xnor U25747 (N_25747,N_24302,N_24900);
nor U25748 (N_25748,N_24731,N_24533);
xnor U25749 (N_25749,N_24643,N_24134);
nand U25750 (N_25750,N_24475,N_24916);
xnor U25751 (N_25751,N_24656,N_24547);
xor U25752 (N_25752,N_24026,N_24221);
xnor U25753 (N_25753,N_24801,N_24016);
and U25754 (N_25754,N_24624,N_24719);
nand U25755 (N_25755,N_24399,N_24241);
nor U25756 (N_25756,N_24110,N_24162);
and U25757 (N_25757,N_24414,N_24753);
nor U25758 (N_25758,N_24532,N_24658);
and U25759 (N_25759,N_24196,N_24892);
and U25760 (N_25760,N_24482,N_24200);
and U25761 (N_25761,N_24955,N_24381);
nand U25762 (N_25762,N_24663,N_24624);
or U25763 (N_25763,N_24288,N_24548);
nand U25764 (N_25764,N_24543,N_24814);
nand U25765 (N_25765,N_24146,N_24764);
or U25766 (N_25766,N_24516,N_24838);
and U25767 (N_25767,N_24427,N_24607);
and U25768 (N_25768,N_24374,N_24611);
or U25769 (N_25769,N_24154,N_24585);
nand U25770 (N_25770,N_24817,N_24005);
nand U25771 (N_25771,N_24096,N_24330);
nor U25772 (N_25772,N_24879,N_24695);
and U25773 (N_25773,N_24634,N_24838);
xor U25774 (N_25774,N_24488,N_24663);
xnor U25775 (N_25775,N_24893,N_24368);
or U25776 (N_25776,N_24991,N_24403);
nor U25777 (N_25777,N_24313,N_24662);
nor U25778 (N_25778,N_24934,N_24680);
or U25779 (N_25779,N_24275,N_24504);
nand U25780 (N_25780,N_24328,N_24814);
xor U25781 (N_25781,N_24971,N_24699);
xnor U25782 (N_25782,N_24839,N_24773);
nor U25783 (N_25783,N_24011,N_24410);
nor U25784 (N_25784,N_24107,N_24748);
and U25785 (N_25785,N_24535,N_24013);
and U25786 (N_25786,N_24232,N_24136);
or U25787 (N_25787,N_24688,N_24232);
or U25788 (N_25788,N_24266,N_24581);
xnor U25789 (N_25789,N_24055,N_24196);
nand U25790 (N_25790,N_24199,N_24621);
or U25791 (N_25791,N_24622,N_24934);
xnor U25792 (N_25792,N_24978,N_24238);
nor U25793 (N_25793,N_24617,N_24869);
xnor U25794 (N_25794,N_24837,N_24208);
nand U25795 (N_25795,N_24703,N_24855);
or U25796 (N_25796,N_24148,N_24476);
or U25797 (N_25797,N_24533,N_24763);
nand U25798 (N_25798,N_24483,N_24385);
xor U25799 (N_25799,N_24424,N_24850);
nand U25800 (N_25800,N_24789,N_24860);
nand U25801 (N_25801,N_24213,N_24244);
nor U25802 (N_25802,N_24405,N_24527);
nor U25803 (N_25803,N_24721,N_24026);
and U25804 (N_25804,N_24116,N_24967);
xnor U25805 (N_25805,N_24384,N_24432);
or U25806 (N_25806,N_24174,N_24972);
xnor U25807 (N_25807,N_24252,N_24561);
and U25808 (N_25808,N_24758,N_24190);
nor U25809 (N_25809,N_24891,N_24558);
and U25810 (N_25810,N_24655,N_24480);
nand U25811 (N_25811,N_24084,N_24586);
nor U25812 (N_25812,N_24816,N_24535);
or U25813 (N_25813,N_24211,N_24300);
or U25814 (N_25814,N_24386,N_24346);
nand U25815 (N_25815,N_24153,N_24888);
nor U25816 (N_25816,N_24651,N_24064);
nor U25817 (N_25817,N_24745,N_24478);
nand U25818 (N_25818,N_24236,N_24091);
xnor U25819 (N_25819,N_24349,N_24618);
or U25820 (N_25820,N_24322,N_24408);
and U25821 (N_25821,N_24256,N_24506);
and U25822 (N_25822,N_24074,N_24627);
nand U25823 (N_25823,N_24925,N_24381);
nor U25824 (N_25824,N_24060,N_24487);
and U25825 (N_25825,N_24123,N_24897);
or U25826 (N_25826,N_24476,N_24650);
or U25827 (N_25827,N_24826,N_24966);
or U25828 (N_25828,N_24859,N_24976);
nand U25829 (N_25829,N_24764,N_24241);
or U25830 (N_25830,N_24908,N_24666);
nor U25831 (N_25831,N_24236,N_24440);
nor U25832 (N_25832,N_24829,N_24351);
nor U25833 (N_25833,N_24741,N_24955);
nand U25834 (N_25834,N_24737,N_24816);
nor U25835 (N_25835,N_24098,N_24515);
or U25836 (N_25836,N_24972,N_24328);
xnor U25837 (N_25837,N_24976,N_24868);
xor U25838 (N_25838,N_24632,N_24211);
nand U25839 (N_25839,N_24839,N_24457);
nor U25840 (N_25840,N_24414,N_24601);
nand U25841 (N_25841,N_24241,N_24242);
or U25842 (N_25842,N_24961,N_24782);
nand U25843 (N_25843,N_24228,N_24185);
and U25844 (N_25844,N_24199,N_24561);
and U25845 (N_25845,N_24839,N_24851);
nand U25846 (N_25846,N_24831,N_24523);
or U25847 (N_25847,N_24425,N_24891);
and U25848 (N_25848,N_24748,N_24642);
nor U25849 (N_25849,N_24050,N_24348);
and U25850 (N_25850,N_24856,N_24144);
xor U25851 (N_25851,N_24947,N_24757);
and U25852 (N_25852,N_24096,N_24371);
xnor U25853 (N_25853,N_24934,N_24342);
and U25854 (N_25854,N_24071,N_24925);
or U25855 (N_25855,N_24780,N_24561);
or U25856 (N_25856,N_24383,N_24293);
nor U25857 (N_25857,N_24178,N_24144);
xor U25858 (N_25858,N_24520,N_24002);
nor U25859 (N_25859,N_24387,N_24188);
or U25860 (N_25860,N_24046,N_24930);
nor U25861 (N_25861,N_24945,N_24513);
or U25862 (N_25862,N_24484,N_24734);
xnor U25863 (N_25863,N_24247,N_24188);
and U25864 (N_25864,N_24229,N_24257);
or U25865 (N_25865,N_24764,N_24914);
or U25866 (N_25866,N_24504,N_24969);
nand U25867 (N_25867,N_24577,N_24492);
or U25868 (N_25868,N_24668,N_24940);
and U25869 (N_25869,N_24392,N_24146);
xor U25870 (N_25870,N_24828,N_24437);
xnor U25871 (N_25871,N_24541,N_24393);
xor U25872 (N_25872,N_24403,N_24566);
nor U25873 (N_25873,N_24072,N_24395);
nor U25874 (N_25874,N_24983,N_24969);
or U25875 (N_25875,N_24513,N_24691);
xnor U25876 (N_25876,N_24327,N_24979);
nand U25877 (N_25877,N_24366,N_24680);
xnor U25878 (N_25878,N_24931,N_24016);
nor U25879 (N_25879,N_24278,N_24423);
nand U25880 (N_25880,N_24195,N_24773);
xnor U25881 (N_25881,N_24357,N_24825);
nor U25882 (N_25882,N_24638,N_24504);
nor U25883 (N_25883,N_24378,N_24706);
or U25884 (N_25884,N_24618,N_24005);
nor U25885 (N_25885,N_24627,N_24676);
nand U25886 (N_25886,N_24790,N_24990);
xnor U25887 (N_25887,N_24145,N_24644);
or U25888 (N_25888,N_24282,N_24883);
or U25889 (N_25889,N_24869,N_24789);
xnor U25890 (N_25890,N_24013,N_24864);
or U25891 (N_25891,N_24715,N_24846);
nand U25892 (N_25892,N_24130,N_24551);
and U25893 (N_25893,N_24545,N_24630);
or U25894 (N_25894,N_24136,N_24298);
nor U25895 (N_25895,N_24307,N_24348);
xnor U25896 (N_25896,N_24301,N_24264);
xor U25897 (N_25897,N_24362,N_24662);
nand U25898 (N_25898,N_24760,N_24607);
xnor U25899 (N_25899,N_24715,N_24325);
xor U25900 (N_25900,N_24888,N_24271);
nor U25901 (N_25901,N_24464,N_24564);
and U25902 (N_25902,N_24351,N_24187);
nand U25903 (N_25903,N_24098,N_24856);
nor U25904 (N_25904,N_24871,N_24611);
xor U25905 (N_25905,N_24998,N_24213);
xor U25906 (N_25906,N_24089,N_24947);
nor U25907 (N_25907,N_24934,N_24088);
nand U25908 (N_25908,N_24434,N_24459);
or U25909 (N_25909,N_24464,N_24480);
or U25910 (N_25910,N_24579,N_24399);
nand U25911 (N_25911,N_24246,N_24943);
and U25912 (N_25912,N_24398,N_24408);
xnor U25913 (N_25913,N_24780,N_24119);
nand U25914 (N_25914,N_24081,N_24324);
xnor U25915 (N_25915,N_24854,N_24226);
or U25916 (N_25916,N_24480,N_24038);
and U25917 (N_25917,N_24870,N_24775);
nor U25918 (N_25918,N_24472,N_24869);
nor U25919 (N_25919,N_24702,N_24856);
and U25920 (N_25920,N_24648,N_24148);
nand U25921 (N_25921,N_24237,N_24434);
nand U25922 (N_25922,N_24406,N_24818);
nand U25923 (N_25923,N_24051,N_24491);
and U25924 (N_25924,N_24476,N_24303);
nor U25925 (N_25925,N_24931,N_24207);
xor U25926 (N_25926,N_24014,N_24742);
or U25927 (N_25927,N_24966,N_24368);
nor U25928 (N_25928,N_24816,N_24531);
and U25929 (N_25929,N_24207,N_24289);
or U25930 (N_25930,N_24591,N_24789);
xor U25931 (N_25931,N_24678,N_24035);
nand U25932 (N_25932,N_24430,N_24127);
xor U25933 (N_25933,N_24341,N_24708);
nor U25934 (N_25934,N_24380,N_24628);
nand U25935 (N_25935,N_24916,N_24669);
nand U25936 (N_25936,N_24828,N_24070);
nand U25937 (N_25937,N_24972,N_24324);
or U25938 (N_25938,N_24536,N_24230);
and U25939 (N_25939,N_24146,N_24955);
and U25940 (N_25940,N_24479,N_24477);
and U25941 (N_25941,N_24585,N_24622);
xor U25942 (N_25942,N_24069,N_24048);
xnor U25943 (N_25943,N_24658,N_24242);
nand U25944 (N_25944,N_24552,N_24748);
nand U25945 (N_25945,N_24866,N_24831);
nand U25946 (N_25946,N_24487,N_24684);
or U25947 (N_25947,N_24629,N_24972);
nor U25948 (N_25948,N_24974,N_24065);
nand U25949 (N_25949,N_24844,N_24813);
nor U25950 (N_25950,N_24235,N_24714);
or U25951 (N_25951,N_24238,N_24332);
xnor U25952 (N_25952,N_24795,N_24782);
or U25953 (N_25953,N_24823,N_24730);
or U25954 (N_25954,N_24083,N_24475);
xor U25955 (N_25955,N_24960,N_24661);
xnor U25956 (N_25956,N_24940,N_24966);
nor U25957 (N_25957,N_24208,N_24337);
and U25958 (N_25958,N_24366,N_24145);
nand U25959 (N_25959,N_24684,N_24786);
nand U25960 (N_25960,N_24693,N_24799);
or U25961 (N_25961,N_24156,N_24902);
nor U25962 (N_25962,N_24624,N_24277);
nor U25963 (N_25963,N_24141,N_24637);
or U25964 (N_25964,N_24909,N_24557);
nor U25965 (N_25965,N_24539,N_24289);
nand U25966 (N_25966,N_24961,N_24550);
and U25967 (N_25967,N_24600,N_24028);
nand U25968 (N_25968,N_24187,N_24919);
nand U25969 (N_25969,N_24629,N_24022);
and U25970 (N_25970,N_24986,N_24605);
nand U25971 (N_25971,N_24159,N_24767);
xnor U25972 (N_25972,N_24196,N_24294);
or U25973 (N_25973,N_24411,N_24692);
and U25974 (N_25974,N_24483,N_24148);
xnor U25975 (N_25975,N_24601,N_24740);
xor U25976 (N_25976,N_24894,N_24617);
nor U25977 (N_25977,N_24581,N_24776);
nor U25978 (N_25978,N_24754,N_24354);
xor U25979 (N_25979,N_24005,N_24635);
nor U25980 (N_25980,N_24051,N_24919);
nor U25981 (N_25981,N_24133,N_24759);
or U25982 (N_25982,N_24490,N_24473);
and U25983 (N_25983,N_24412,N_24287);
and U25984 (N_25984,N_24433,N_24601);
or U25985 (N_25985,N_24512,N_24397);
and U25986 (N_25986,N_24628,N_24202);
nand U25987 (N_25987,N_24896,N_24025);
xnor U25988 (N_25988,N_24933,N_24665);
nand U25989 (N_25989,N_24596,N_24437);
nor U25990 (N_25990,N_24754,N_24903);
nand U25991 (N_25991,N_24630,N_24570);
nand U25992 (N_25992,N_24767,N_24674);
nor U25993 (N_25993,N_24444,N_24150);
or U25994 (N_25994,N_24302,N_24606);
or U25995 (N_25995,N_24005,N_24577);
xnor U25996 (N_25996,N_24541,N_24791);
xnor U25997 (N_25997,N_24531,N_24227);
nand U25998 (N_25998,N_24900,N_24733);
nand U25999 (N_25999,N_24995,N_24533);
and U26000 (N_26000,N_25181,N_25304);
nor U26001 (N_26001,N_25872,N_25258);
and U26002 (N_26002,N_25243,N_25906);
nand U26003 (N_26003,N_25740,N_25577);
or U26004 (N_26004,N_25589,N_25285);
nor U26005 (N_26005,N_25964,N_25163);
nor U26006 (N_26006,N_25913,N_25961);
xor U26007 (N_26007,N_25466,N_25045);
or U26008 (N_26008,N_25886,N_25346);
xnor U26009 (N_26009,N_25752,N_25804);
nor U26010 (N_26010,N_25713,N_25338);
nor U26011 (N_26011,N_25691,N_25493);
xor U26012 (N_26012,N_25729,N_25788);
nor U26013 (N_26013,N_25647,N_25301);
nor U26014 (N_26014,N_25296,N_25094);
or U26015 (N_26015,N_25649,N_25267);
and U26016 (N_26016,N_25079,N_25499);
nor U26017 (N_26017,N_25411,N_25785);
nand U26018 (N_26018,N_25707,N_25238);
and U26019 (N_26019,N_25613,N_25453);
or U26020 (N_26020,N_25309,N_25474);
nor U26021 (N_26021,N_25391,N_25443);
or U26022 (N_26022,N_25814,N_25731);
nor U26023 (N_26023,N_25706,N_25699);
or U26024 (N_26024,N_25171,N_25746);
nand U26025 (N_26025,N_25637,N_25152);
and U26026 (N_26026,N_25695,N_25794);
nor U26027 (N_26027,N_25584,N_25147);
and U26028 (N_26028,N_25719,N_25869);
xnor U26029 (N_26029,N_25290,N_25970);
xnor U26030 (N_26030,N_25641,N_25182);
and U26031 (N_26031,N_25583,N_25481);
nand U26032 (N_26032,N_25862,N_25011);
or U26033 (N_26033,N_25421,N_25907);
or U26034 (N_26034,N_25401,N_25784);
nand U26035 (N_26035,N_25573,N_25984);
or U26036 (N_26036,N_25703,N_25217);
xnor U26037 (N_26037,N_25292,N_25263);
nor U26038 (N_26038,N_25146,N_25418);
xnor U26039 (N_26039,N_25787,N_25980);
and U26040 (N_26040,N_25435,N_25708);
or U26041 (N_26041,N_25333,N_25128);
and U26042 (N_26042,N_25259,N_25680);
and U26043 (N_26043,N_25926,N_25008);
nor U26044 (N_26044,N_25324,N_25640);
nor U26045 (N_26045,N_25711,N_25581);
nor U26046 (N_26046,N_25039,N_25818);
xnor U26047 (N_26047,N_25714,N_25214);
nor U26048 (N_26048,N_25870,N_25656);
xnor U26049 (N_26049,N_25168,N_25652);
nor U26050 (N_26050,N_25227,N_25810);
xnor U26051 (N_26051,N_25132,N_25200);
or U26052 (N_26052,N_25251,N_25479);
nand U26053 (N_26053,N_25544,N_25464);
nand U26054 (N_26054,N_25115,N_25622);
nand U26055 (N_26055,N_25275,N_25545);
or U26056 (N_26056,N_25276,N_25305);
or U26057 (N_26057,N_25611,N_25898);
xor U26058 (N_26058,N_25193,N_25023);
xor U26059 (N_26059,N_25032,N_25547);
nand U26060 (N_26060,N_25187,N_25004);
or U26061 (N_26061,N_25874,N_25058);
nand U26062 (N_26062,N_25475,N_25674);
nand U26063 (N_26063,N_25815,N_25018);
xor U26064 (N_26064,N_25138,N_25060);
and U26065 (N_26065,N_25384,N_25437);
nor U26066 (N_26066,N_25976,N_25949);
or U26067 (N_26067,N_25635,N_25295);
xor U26068 (N_26068,N_25073,N_25014);
xnor U26069 (N_26069,N_25722,N_25001);
and U26070 (N_26070,N_25151,N_25609);
and U26071 (N_26071,N_25947,N_25038);
or U26072 (N_26072,N_25113,N_25955);
xnor U26073 (N_26073,N_25123,N_25610);
or U26074 (N_26074,N_25894,N_25929);
and U26075 (N_26075,N_25413,N_25364);
and U26076 (N_26076,N_25447,N_25972);
or U26077 (N_26077,N_25239,N_25742);
or U26078 (N_26078,N_25412,N_25716);
nor U26079 (N_26079,N_25944,N_25678);
or U26080 (N_26080,N_25865,N_25877);
nand U26081 (N_26081,N_25724,N_25519);
or U26082 (N_26082,N_25288,N_25308);
xor U26083 (N_26083,N_25672,N_25013);
nand U26084 (N_26084,N_25530,N_25236);
nand U26085 (N_26085,N_25310,N_25910);
nand U26086 (N_26086,N_25670,N_25378);
nor U26087 (N_26087,N_25504,N_25988);
nand U26088 (N_26088,N_25556,N_25423);
xnor U26089 (N_26089,N_25667,N_25974);
nor U26090 (N_26090,N_25527,N_25415);
and U26091 (N_26091,N_25650,N_25173);
or U26092 (N_26092,N_25780,N_25921);
nand U26093 (N_26093,N_25912,N_25766);
or U26094 (N_26094,N_25330,N_25127);
or U26095 (N_26095,N_25511,N_25157);
and U26096 (N_26096,N_25449,N_25800);
nor U26097 (N_26097,N_25122,N_25430);
and U26098 (N_26098,N_25931,N_25560);
or U26099 (N_26099,N_25158,N_25407);
nor U26100 (N_26100,N_25653,N_25823);
nor U26101 (N_26101,N_25260,N_25646);
or U26102 (N_26102,N_25344,N_25059);
or U26103 (N_26103,N_25489,N_25782);
or U26104 (N_26104,N_25508,N_25044);
nor U26105 (N_26105,N_25375,N_25194);
or U26106 (N_26106,N_25935,N_25126);
and U26107 (N_26107,N_25328,N_25743);
nor U26108 (N_26108,N_25473,N_25916);
or U26109 (N_26109,N_25091,N_25728);
nor U26110 (N_26110,N_25311,N_25734);
xnor U26111 (N_26111,N_25410,N_25468);
or U26112 (N_26112,N_25130,N_25586);
nor U26113 (N_26113,N_25027,N_25639);
xnor U26114 (N_26114,N_25454,N_25587);
xor U26115 (N_26115,N_25566,N_25306);
and U26116 (N_26116,N_25958,N_25179);
xnor U26117 (N_26117,N_25188,N_25186);
xnor U26118 (N_26118,N_25209,N_25141);
nand U26119 (N_26119,N_25593,N_25078);
and U26120 (N_26120,N_25503,N_25167);
and U26121 (N_26121,N_25007,N_25245);
nor U26122 (N_26122,N_25117,N_25143);
xor U26123 (N_26123,N_25485,N_25879);
nand U26124 (N_26124,N_25568,N_25360);
nor U26125 (N_26125,N_25222,N_25244);
nor U26126 (N_26126,N_25325,N_25085);
nand U26127 (N_26127,N_25923,N_25993);
xor U26128 (N_26128,N_25054,N_25737);
nand U26129 (N_26129,N_25274,N_25416);
and U26130 (N_26130,N_25831,N_25162);
and U26131 (N_26131,N_25010,N_25514);
nor U26132 (N_26132,N_25405,N_25658);
or U26133 (N_26133,N_25465,N_25192);
nor U26134 (N_26134,N_25500,N_25121);
xnor U26135 (N_26135,N_25074,N_25442);
or U26136 (N_26136,N_25172,N_25751);
and U26137 (N_26137,N_25666,N_25139);
and U26138 (N_26138,N_25878,N_25889);
nand U26139 (N_26139,N_25155,N_25567);
and U26140 (N_26140,N_25299,N_25377);
or U26141 (N_26141,N_25273,N_25843);
nor U26142 (N_26142,N_25215,N_25882);
nor U26143 (N_26143,N_25166,N_25165);
nor U26144 (N_26144,N_25506,N_25943);
or U26145 (N_26145,N_25914,N_25374);
nor U26146 (N_26146,N_25924,N_25414);
and U26147 (N_26147,N_25019,N_25402);
xnor U26148 (N_26148,N_25739,N_25960);
xnor U26149 (N_26149,N_25406,N_25394);
or U26150 (N_26150,N_25681,N_25210);
and U26151 (N_26151,N_25314,N_25232);
or U26152 (N_26152,N_25517,N_25749);
nor U26153 (N_26153,N_25125,N_25833);
nand U26154 (N_26154,N_25067,N_25247);
or U26155 (N_26155,N_25747,N_25745);
xnor U26156 (N_26156,N_25837,N_25438);
and U26157 (N_26157,N_25962,N_25642);
or U26158 (N_26158,N_25389,N_25266);
or U26159 (N_26159,N_25012,N_25286);
and U26160 (N_26160,N_25118,N_25614);
and U26161 (N_26161,N_25081,N_25180);
or U26162 (N_26162,N_25189,N_25633);
and U26163 (N_26163,N_25645,N_25093);
nor U26164 (N_26164,N_25852,N_25026);
nand U26165 (N_26165,N_25665,N_25873);
and U26166 (N_26166,N_25417,N_25813);
or U26167 (N_26167,N_25994,N_25548);
xnor U26168 (N_26168,N_25488,N_25730);
nand U26169 (N_26169,N_25327,N_25805);
xor U26170 (N_26170,N_25520,N_25677);
or U26171 (N_26171,N_25630,N_25591);
or U26172 (N_26172,N_25682,N_25967);
and U26173 (N_26173,N_25846,N_25709);
nor U26174 (N_26174,N_25601,N_25732);
or U26175 (N_26175,N_25144,N_25900);
nor U26176 (N_26176,N_25190,N_25684);
or U26177 (N_26177,N_25829,N_25408);
xor U26178 (N_26178,N_25204,N_25765);
xnor U26179 (N_26179,N_25340,N_25509);
xor U26180 (N_26180,N_25973,N_25808);
nor U26181 (N_26181,N_25398,N_25097);
and U26182 (N_26182,N_25277,N_25062);
or U26183 (N_26183,N_25319,N_25977);
nor U26184 (N_26184,N_25524,N_25817);
or U26185 (N_26185,N_25542,N_25801);
or U26186 (N_26186,N_25753,N_25133);
or U26187 (N_26187,N_25875,N_25033);
and U26188 (N_26188,N_25480,N_25693);
or U26189 (N_26189,N_25009,N_25469);
nor U26190 (N_26190,N_25307,N_25925);
xnor U26191 (N_26191,N_25380,N_25868);
and U26192 (N_26192,N_25890,N_25712);
nor U26193 (N_26193,N_25688,N_25441);
and U26194 (N_26194,N_25331,N_25848);
xnor U26195 (N_26195,N_25066,N_25888);
xor U26196 (N_26196,N_25024,N_25904);
and U26197 (N_26197,N_25250,N_25426);
nand U26198 (N_26198,N_25390,N_25359);
xnor U26199 (N_26199,N_25679,N_25803);
nor U26200 (N_26200,N_25648,N_25068);
and U26201 (N_26201,N_25574,N_25521);
or U26202 (N_26202,N_25917,N_25588);
xor U26203 (N_26203,N_25150,N_25940);
and U26204 (N_26204,N_25554,N_25347);
nand U26205 (N_26205,N_25439,N_25183);
xor U26206 (N_26206,N_25300,N_25725);
or U26207 (N_26207,N_25042,N_25109);
nor U26208 (N_26208,N_25756,N_25733);
or U26209 (N_26209,N_25120,N_25358);
nor U26210 (N_26210,N_25992,N_25897);
xor U26211 (N_26211,N_25356,N_25534);
or U26212 (N_26212,N_25885,N_25616);
and U26213 (N_26213,N_25603,N_25891);
nand U26214 (N_26214,N_25065,N_25839);
or U26215 (N_26215,N_25116,N_25371);
xor U26216 (N_26216,N_25908,N_25536);
nand U26217 (N_26217,N_25860,N_25219);
and U26218 (N_26218,N_25284,N_25088);
and U26219 (N_26219,N_25516,N_25883);
and U26220 (N_26220,N_25821,N_25856);
xor U26221 (N_26221,N_25540,N_25563);
or U26222 (N_26222,N_25963,N_25137);
nor U26223 (N_26223,N_25156,N_25332);
or U26224 (N_26224,N_25802,N_25807);
xnor U26225 (N_26225,N_25927,N_25768);
xor U26226 (N_26226,N_25754,N_25741);
or U26227 (N_26227,N_25507,N_25099);
or U26228 (N_26228,N_25792,N_25220);
or U26229 (N_26229,N_25990,N_25965);
xnor U26230 (N_26230,N_25142,N_25847);
nand U26231 (N_26231,N_25386,N_25979);
xor U26232 (N_26232,N_25098,N_25261);
nand U26233 (N_26233,N_25558,N_25483);
or U26234 (N_26234,N_25694,N_25953);
nand U26235 (N_26235,N_25427,N_25580);
xor U26236 (N_26236,N_25450,N_25590);
nand U26237 (N_26237,N_25820,N_25363);
nor U26238 (N_26238,N_25498,N_25177);
nor U26239 (N_26239,N_25382,N_25549);
nor U26240 (N_26240,N_25030,N_25854);
and U26241 (N_26241,N_25592,N_25842);
and U26242 (N_26242,N_25050,N_25760);
xor U26243 (N_26243,N_25899,N_25859);
nand U26244 (N_26244,N_25697,N_25218);
and U26245 (N_26245,N_25928,N_25880);
nand U26246 (N_26246,N_25954,N_25775);
or U26247 (N_26247,N_25777,N_25996);
or U26248 (N_26248,N_25104,N_25750);
or U26249 (N_26249,N_25089,N_25334);
or U26250 (N_26250,N_25832,N_25323);
nor U26251 (N_26251,N_25281,N_25084);
nor U26252 (N_26252,N_25564,N_25106);
nor U26253 (N_26253,N_25216,N_25235);
and U26254 (N_26254,N_25983,N_25770);
nor U26255 (N_26255,N_25518,N_25298);
or U26256 (N_26256,N_25830,N_25255);
nor U26257 (N_26257,N_25531,N_25772);
xor U26258 (N_26258,N_25134,N_25294);
nand U26259 (N_26259,N_25687,N_25903);
xor U26260 (N_26260,N_25096,N_25896);
nor U26261 (N_26261,N_25392,N_25029);
and U26262 (N_26262,N_25322,N_25625);
nor U26263 (N_26263,N_25257,N_25835);
nand U26264 (N_26264,N_25605,N_25948);
or U26265 (N_26265,N_25495,N_25755);
nor U26266 (N_26266,N_25595,N_25505);
or U26267 (N_26267,N_25981,N_25178);
and U26268 (N_26268,N_25971,N_25486);
and U26269 (N_26269,N_25072,N_25361);
nand U26270 (N_26270,N_25381,N_25002);
nand U26271 (N_26271,N_25783,N_25000);
or U26272 (N_26272,N_25069,N_25812);
nor U26273 (N_26273,N_25892,N_25048);
or U26274 (N_26274,N_25434,N_25119);
nor U26275 (N_26275,N_25339,N_25234);
nand U26276 (N_26276,N_25689,N_25102);
nor U26277 (N_26277,N_25368,N_25020);
xnor U26278 (N_26278,N_25211,N_25612);
and U26279 (N_26279,N_25440,N_25692);
xor U26280 (N_26280,N_25901,N_25834);
xnor U26281 (N_26281,N_25477,N_25607);
xor U26282 (N_26282,N_25422,N_25491);
nand U26283 (N_26283,N_25715,N_25055);
and U26284 (N_26284,N_25893,N_25525);
nor U26285 (N_26285,N_25052,N_25930);
nand U26286 (N_26286,N_25387,N_25199);
xor U26287 (N_26287,N_25826,N_25271);
nand U26288 (N_26288,N_25723,N_25664);
and U26289 (N_26289,N_25950,N_25510);
nand U26290 (N_26290,N_25087,N_25773);
or U26291 (N_26291,N_25424,N_25279);
xnor U26292 (N_26292,N_25425,N_25638);
xnor U26293 (N_26293,N_25982,N_25482);
and U26294 (N_26294,N_25532,N_25655);
or U26295 (N_26295,N_25017,N_25539);
and U26296 (N_26296,N_25562,N_25629);
xor U26297 (N_26297,N_25341,N_25861);
xnor U26298 (N_26298,N_25683,N_25129);
or U26299 (N_26299,N_25397,N_25557);
and U26300 (N_26300,N_25372,N_25103);
or U26301 (N_26301,N_25432,N_25938);
nand U26302 (N_26302,N_25105,N_25720);
or U26303 (N_26303,N_25207,N_25080);
xnor U26304 (N_26304,N_25999,N_25932);
and U26305 (N_26305,N_25618,N_25623);
nor U26306 (N_26306,N_25902,N_25634);
xnor U26307 (N_26307,N_25201,N_25543);
xor U26308 (N_26308,N_25660,N_25791);
nor U26309 (N_26309,N_25855,N_25918);
xnor U26310 (N_26310,N_25185,N_25701);
or U26311 (N_26311,N_25806,N_25668);
xnor U26312 (N_26312,N_25778,N_25654);
or U26313 (N_26313,N_25352,N_25051);
nand U26314 (N_26314,N_25169,N_25090);
or U26315 (N_26315,N_25253,N_25241);
nor U26316 (N_26316,N_25035,N_25986);
nand U26317 (N_26317,N_25569,N_25597);
nor U26318 (N_26318,N_25721,N_25797);
or U26319 (N_26319,N_25462,N_25537);
and U26320 (N_26320,N_25124,N_25991);
or U26321 (N_26321,N_25501,N_25620);
nor U26322 (N_26322,N_25249,N_25686);
nor U26323 (N_26323,N_25700,N_25799);
xnor U26324 (N_26324,N_25451,N_25049);
or U26325 (N_26325,N_25436,N_25936);
nor U26326 (N_26326,N_25946,N_25196);
nor U26327 (N_26327,N_25448,N_25184);
nor U26328 (N_26328,N_25403,N_25095);
xnor U26329 (N_26329,N_25457,N_25578);
nand U26330 (N_26330,N_25366,N_25937);
and U26331 (N_26331,N_25348,N_25321);
nand U26332 (N_26332,N_25718,N_25283);
and U26333 (N_26333,N_25552,N_25576);
nand U26334 (N_26334,N_25675,N_25853);
or U26335 (N_26335,N_25248,N_25396);
nor U26336 (N_26336,N_25798,N_25452);
and U26337 (N_26337,N_25351,N_25786);
and U26338 (N_26338,N_25819,N_25496);
xor U26339 (N_26339,N_25355,N_25082);
or U26340 (N_26340,N_25343,N_25037);
nor U26341 (N_26341,N_25758,N_25114);
nor U26342 (N_26342,N_25353,N_25269);
and U26343 (N_26343,N_25342,N_25529);
and U26344 (N_26344,N_25278,N_25467);
nor U26345 (N_26345,N_25769,N_25998);
xnor U26346 (N_26346,N_25841,N_25598);
xnor U26347 (N_26347,N_25456,N_25828);
or U26348 (N_26348,N_25206,N_25570);
and U26349 (N_26349,N_25604,N_25825);
xnor U26350 (N_26350,N_25282,N_25100);
nand U26351 (N_26351,N_25594,N_25208);
or U26352 (N_26352,N_25111,N_25659);
and U26353 (N_26353,N_25148,N_25617);
xor U26354 (N_26354,N_25523,N_25636);
nor U26355 (N_26355,N_25256,N_25393);
nand U26356 (N_26356,N_25911,N_25112);
or U26357 (N_26357,N_25779,N_25136);
or U26358 (N_26358,N_25565,N_25851);
nand U26359 (N_26359,N_25264,N_25350);
nor U26360 (N_26360,N_25316,N_25538);
or U26361 (N_26361,N_25388,N_25280);
xnor U26362 (N_26362,N_25909,N_25744);
and U26363 (N_26363,N_25761,N_25661);
xor U26364 (N_26364,N_25915,N_25034);
nand U26365 (N_26365,N_25795,N_25108);
xnor U26366 (N_26366,N_25223,N_25313);
and U26367 (N_26367,N_25064,N_25240);
nor U26368 (N_26368,N_25864,N_25345);
xnor U26369 (N_26369,N_25838,N_25989);
nor U26370 (N_26370,N_25513,N_25561);
nand U26371 (N_26371,N_25671,N_25231);
xor U26372 (N_26372,N_25246,N_25336);
nor U26373 (N_26373,N_25252,N_25289);
nor U26374 (N_26374,N_25458,N_25337);
nand U26375 (N_26375,N_25871,N_25317);
and U26376 (N_26376,N_25383,N_25349);
xor U26377 (N_26377,N_25365,N_25022);
xnor U26378 (N_26378,N_25478,N_25226);
and U26379 (N_26379,N_25431,N_25400);
nand U26380 (N_26380,N_25161,N_25229);
xnor U26381 (N_26381,N_25484,N_25367);
and U26382 (N_26382,N_25164,N_25939);
or U26383 (N_26383,N_25702,N_25762);
xnor U26384 (N_26384,N_25016,N_25522);
nand U26385 (N_26385,N_25789,N_25228);
nor U26386 (N_26386,N_25541,N_25419);
nand U26387 (N_26387,N_25320,N_25941);
nand U26388 (N_26388,N_25003,N_25881);
nand U26389 (N_26389,N_25420,N_25985);
nor U26390 (N_26390,N_25959,N_25767);
nor U26391 (N_26391,N_25738,N_25781);
nand U26392 (N_26392,N_25905,N_25370);
nand U26393 (N_26393,N_25487,N_25302);
nand U26394 (N_26394,N_25698,N_25312);
and U26395 (N_26395,N_25174,N_25175);
nor U26396 (N_26396,N_25673,N_25476);
or U26397 (N_26397,N_25705,N_25662);
nand U26398 (N_26398,N_25101,N_25056);
and U26399 (N_26399,N_25533,N_25585);
nand U26400 (N_26400,N_25727,N_25836);
or U26401 (N_26401,N_25497,N_25197);
xnor U26402 (N_26402,N_25224,N_25041);
and U26403 (N_26403,N_25287,N_25445);
nand U26404 (N_26404,N_25061,N_25070);
nor U26405 (N_26405,N_25472,N_25212);
or U26406 (N_26406,N_25512,N_25811);
and U26407 (N_26407,N_25053,N_25006);
and U26408 (N_26408,N_25028,N_25376);
and U26409 (N_26409,N_25043,N_25460);
nor U26410 (N_26410,N_25131,N_25771);
xnor U26411 (N_26411,N_25546,N_25774);
nand U26412 (N_26412,N_25357,N_25515);
xnor U26413 (N_26413,N_25876,N_25047);
nand U26414 (N_26414,N_25233,N_25599);
or U26415 (N_26415,N_25303,N_25942);
or U26416 (N_26416,N_25202,N_25968);
xor U26417 (N_26417,N_25957,N_25373);
nand U26418 (N_26418,N_25490,N_25225);
or U26419 (N_26419,N_25385,N_25444);
and U26420 (N_26420,N_25628,N_25262);
nor U26421 (N_26421,N_25643,N_25575);
nand U26422 (N_26422,N_25685,N_25757);
nor U26423 (N_26423,N_25987,N_25297);
xor U26424 (N_26424,N_25572,N_25461);
and U26425 (N_26425,N_25696,N_25615);
nor U26426 (N_26426,N_25135,N_25031);
xor U26427 (N_26427,N_25046,N_25887);
xnor U26428 (N_26428,N_25149,N_25471);
or U26429 (N_26429,N_25827,N_25040);
or U26430 (N_26430,N_25850,N_25763);
nor U26431 (N_26431,N_25369,N_25748);
nand U26432 (N_26432,N_25221,N_25845);
nor U26433 (N_26433,N_25145,N_25822);
xor U26434 (N_26434,N_25550,N_25951);
nor U26435 (N_26435,N_25626,N_25857);
and U26436 (N_26436,N_25934,N_25717);
and U26437 (N_26437,N_25764,N_25619);
or U26438 (N_26438,N_25559,N_25866);
and U26439 (N_26439,N_25291,N_25463);
nor U26440 (N_26440,N_25057,N_25867);
nand U26441 (N_26441,N_25608,N_25395);
and U26442 (N_26442,N_25690,N_25657);
xnor U26443 (N_26443,N_25600,N_25796);
nor U26444 (N_26444,N_25315,N_25083);
nand U26445 (N_26445,N_25154,N_25021);
nor U26446 (N_26446,N_25956,N_25176);
or U26447 (N_26447,N_25759,N_25663);
or U26448 (N_26448,N_25621,N_25318);
xnor U26449 (N_26449,N_25110,N_25997);
or U26450 (N_26450,N_25840,N_25596);
nor U26451 (N_26451,N_25726,N_25428);
and U26452 (N_26452,N_25704,N_25293);
nand U26453 (N_26453,N_25254,N_25502);
xor U26454 (N_26454,N_25409,N_25242);
nor U26455 (N_26455,N_25553,N_25230);
nor U26456 (N_26456,N_25526,N_25107);
nor U26457 (N_26457,N_25459,N_25092);
and U26458 (N_26458,N_25535,N_25582);
xor U26459 (N_26459,N_25790,N_25995);
nand U26460 (N_26460,N_25579,N_25237);
and U26461 (N_26461,N_25071,N_25433);
xnor U26462 (N_26462,N_25153,N_25268);
or U26463 (N_26463,N_25858,N_25933);
and U26464 (N_26464,N_25606,N_25159);
and U26465 (N_26465,N_25969,N_25270);
nor U26466 (N_26466,N_25492,N_25555);
xor U26467 (N_26467,N_25494,N_25329);
and U26468 (N_26468,N_25076,N_25624);
and U26469 (N_26469,N_25326,N_25170);
xnor U26470 (N_26470,N_25335,N_25404);
nand U26471 (N_26471,N_25651,N_25455);
nor U26472 (N_26472,N_25191,N_25140);
nor U26473 (N_26473,N_25005,N_25816);
or U26474 (N_26474,N_25922,N_25863);
nor U26475 (N_26475,N_25205,N_25015);
nor U26476 (N_26476,N_25776,N_25978);
nor U26477 (N_26477,N_25793,N_25919);
nand U26478 (N_26478,N_25362,N_25824);
nand U26479 (N_26479,N_25470,N_25429);
nand U26480 (N_26480,N_25920,N_25945);
or U26481 (N_26481,N_25195,N_25446);
xnor U26482 (N_26482,N_25075,N_25086);
nand U26483 (N_26483,N_25602,N_25036);
nor U26484 (N_26484,N_25399,N_25631);
xor U26485 (N_26485,N_25077,N_25644);
xnor U26486 (N_26486,N_25952,N_25735);
nand U26487 (N_26487,N_25632,N_25966);
nor U26488 (N_26488,N_25975,N_25379);
nor U26489 (N_26489,N_25272,N_25895);
nor U26490 (N_26490,N_25213,N_25809);
nand U26491 (N_26491,N_25884,N_25669);
or U26492 (N_26492,N_25203,N_25627);
nor U26493 (N_26493,N_25849,N_25571);
nand U26494 (N_26494,N_25063,N_25198);
xor U26495 (N_26495,N_25160,N_25265);
or U26496 (N_26496,N_25710,N_25736);
or U26497 (N_26497,N_25528,N_25025);
xnor U26498 (N_26498,N_25354,N_25551);
nand U26499 (N_26499,N_25676,N_25844);
and U26500 (N_26500,N_25073,N_25142);
xnor U26501 (N_26501,N_25840,N_25212);
nor U26502 (N_26502,N_25246,N_25230);
nand U26503 (N_26503,N_25938,N_25672);
nand U26504 (N_26504,N_25553,N_25697);
and U26505 (N_26505,N_25302,N_25062);
nand U26506 (N_26506,N_25933,N_25633);
nor U26507 (N_26507,N_25941,N_25767);
nor U26508 (N_26508,N_25393,N_25803);
nor U26509 (N_26509,N_25015,N_25283);
xor U26510 (N_26510,N_25263,N_25169);
nor U26511 (N_26511,N_25057,N_25395);
nor U26512 (N_26512,N_25181,N_25509);
xor U26513 (N_26513,N_25060,N_25687);
and U26514 (N_26514,N_25578,N_25454);
and U26515 (N_26515,N_25315,N_25880);
xor U26516 (N_26516,N_25566,N_25371);
or U26517 (N_26517,N_25049,N_25956);
nand U26518 (N_26518,N_25820,N_25271);
and U26519 (N_26519,N_25711,N_25396);
xor U26520 (N_26520,N_25532,N_25615);
and U26521 (N_26521,N_25071,N_25202);
or U26522 (N_26522,N_25998,N_25197);
xnor U26523 (N_26523,N_25045,N_25343);
and U26524 (N_26524,N_25334,N_25196);
nor U26525 (N_26525,N_25777,N_25170);
xnor U26526 (N_26526,N_25163,N_25503);
and U26527 (N_26527,N_25280,N_25917);
and U26528 (N_26528,N_25729,N_25156);
nor U26529 (N_26529,N_25816,N_25160);
and U26530 (N_26530,N_25527,N_25479);
and U26531 (N_26531,N_25077,N_25711);
nor U26532 (N_26532,N_25448,N_25511);
and U26533 (N_26533,N_25070,N_25623);
nand U26534 (N_26534,N_25248,N_25432);
nand U26535 (N_26535,N_25060,N_25805);
and U26536 (N_26536,N_25644,N_25700);
nor U26537 (N_26537,N_25699,N_25325);
or U26538 (N_26538,N_25847,N_25632);
nor U26539 (N_26539,N_25815,N_25918);
nor U26540 (N_26540,N_25728,N_25042);
nand U26541 (N_26541,N_25972,N_25001);
nand U26542 (N_26542,N_25761,N_25689);
xnor U26543 (N_26543,N_25191,N_25968);
nand U26544 (N_26544,N_25407,N_25417);
xnor U26545 (N_26545,N_25885,N_25272);
xnor U26546 (N_26546,N_25644,N_25044);
and U26547 (N_26547,N_25923,N_25700);
xnor U26548 (N_26548,N_25556,N_25668);
nor U26549 (N_26549,N_25775,N_25766);
and U26550 (N_26550,N_25513,N_25627);
or U26551 (N_26551,N_25790,N_25042);
xor U26552 (N_26552,N_25528,N_25576);
or U26553 (N_26553,N_25727,N_25096);
nor U26554 (N_26554,N_25487,N_25418);
nand U26555 (N_26555,N_25352,N_25261);
xnor U26556 (N_26556,N_25205,N_25615);
and U26557 (N_26557,N_25982,N_25439);
and U26558 (N_26558,N_25307,N_25630);
and U26559 (N_26559,N_25767,N_25578);
nor U26560 (N_26560,N_25286,N_25402);
xor U26561 (N_26561,N_25674,N_25794);
nand U26562 (N_26562,N_25000,N_25722);
or U26563 (N_26563,N_25565,N_25770);
or U26564 (N_26564,N_25808,N_25719);
and U26565 (N_26565,N_25835,N_25612);
or U26566 (N_26566,N_25087,N_25342);
and U26567 (N_26567,N_25604,N_25023);
xnor U26568 (N_26568,N_25387,N_25538);
xnor U26569 (N_26569,N_25181,N_25614);
and U26570 (N_26570,N_25842,N_25738);
xor U26571 (N_26571,N_25634,N_25673);
or U26572 (N_26572,N_25809,N_25990);
xnor U26573 (N_26573,N_25383,N_25309);
or U26574 (N_26574,N_25009,N_25927);
nand U26575 (N_26575,N_25785,N_25045);
nor U26576 (N_26576,N_25034,N_25141);
nand U26577 (N_26577,N_25344,N_25417);
nor U26578 (N_26578,N_25155,N_25244);
or U26579 (N_26579,N_25383,N_25641);
and U26580 (N_26580,N_25487,N_25887);
and U26581 (N_26581,N_25595,N_25164);
and U26582 (N_26582,N_25881,N_25057);
and U26583 (N_26583,N_25654,N_25503);
nand U26584 (N_26584,N_25124,N_25690);
and U26585 (N_26585,N_25391,N_25093);
xnor U26586 (N_26586,N_25094,N_25031);
nor U26587 (N_26587,N_25244,N_25274);
and U26588 (N_26588,N_25479,N_25923);
and U26589 (N_26589,N_25583,N_25623);
xor U26590 (N_26590,N_25168,N_25251);
nor U26591 (N_26591,N_25641,N_25761);
xor U26592 (N_26592,N_25672,N_25727);
nand U26593 (N_26593,N_25747,N_25808);
xnor U26594 (N_26594,N_25758,N_25693);
or U26595 (N_26595,N_25171,N_25205);
xnor U26596 (N_26596,N_25281,N_25324);
or U26597 (N_26597,N_25501,N_25164);
and U26598 (N_26598,N_25851,N_25077);
nor U26599 (N_26599,N_25265,N_25429);
and U26600 (N_26600,N_25489,N_25461);
xnor U26601 (N_26601,N_25638,N_25709);
nand U26602 (N_26602,N_25309,N_25001);
nand U26603 (N_26603,N_25739,N_25962);
nand U26604 (N_26604,N_25663,N_25550);
nor U26605 (N_26605,N_25789,N_25721);
xor U26606 (N_26606,N_25470,N_25358);
nor U26607 (N_26607,N_25498,N_25125);
and U26608 (N_26608,N_25760,N_25598);
nor U26609 (N_26609,N_25686,N_25741);
xnor U26610 (N_26610,N_25623,N_25513);
nor U26611 (N_26611,N_25143,N_25249);
nor U26612 (N_26612,N_25407,N_25133);
xnor U26613 (N_26613,N_25617,N_25561);
xnor U26614 (N_26614,N_25519,N_25226);
nand U26615 (N_26615,N_25146,N_25179);
or U26616 (N_26616,N_25863,N_25168);
or U26617 (N_26617,N_25568,N_25907);
nor U26618 (N_26618,N_25617,N_25269);
and U26619 (N_26619,N_25594,N_25967);
nand U26620 (N_26620,N_25376,N_25706);
nand U26621 (N_26621,N_25701,N_25258);
and U26622 (N_26622,N_25872,N_25109);
or U26623 (N_26623,N_25658,N_25153);
nor U26624 (N_26624,N_25389,N_25324);
or U26625 (N_26625,N_25821,N_25639);
and U26626 (N_26626,N_25506,N_25439);
nor U26627 (N_26627,N_25265,N_25872);
nand U26628 (N_26628,N_25777,N_25269);
xnor U26629 (N_26629,N_25329,N_25252);
or U26630 (N_26630,N_25906,N_25500);
nor U26631 (N_26631,N_25589,N_25498);
or U26632 (N_26632,N_25991,N_25977);
and U26633 (N_26633,N_25289,N_25766);
nand U26634 (N_26634,N_25336,N_25756);
xor U26635 (N_26635,N_25129,N_25632);
nor U26636 (N_26636,N_25799,N_25053);
and U26637 (N_26637,N_25781,N_25197);
or U26638 (N_26638,N_25755,N_25140);
nor U26639 (N_26639,N_25662,N_25152);
nand U26640 (N_26640,N_25829,N_25620);
nor U26641 (N_26641,N_25287,N_25152);
nor U26642 (N_26642,N_25063,N_25315);
and U26643 (N_26643,N_25319,N_25378);
nand U26644 (N_26644,N_25880,N_25327);
nor U26645 (N_26645,N_25867,N_25846);
xnor U26646 (N_26646,N_25313,N_25290);
or U26647 (N_26647,N_25814,N_25902);
and U26648 (N_26648,N_25340,N_25117);
xor U26649 (N_26649,N_25557,N_25205);
nand U26650 (N_26650,N_25747,N_25555);
nand U26651 (N_26651,N_25031,N_25911);
nand U26652 (N_26652,N_25045,N_25403);
xor U26653 (N_26653,N_25282,N_25693);
nand U26654 (N_26654,N_25597,N_25070);
or U26655 (N_26655,N_25013,N_25573);
nor U26656 (N_26656,N_25174,N_25504);
and U26657 (N_26657,N_25791,N_25729);
xnor U26658 (N_26658,N_25042,N_25205);
nand U26659 (N_26659,N_25393,N_25921);
and U26660 (N_26660,N_25124,N_25513);
nand U26661 (N_26661,N_25865,N_25153);
or U26662 (N_26662,N_25219,N_25787);
nand U26663 (N_26663,N_25637,N_25339);
xor U26664 (N_26664,N_25903,N_25256);
nor U26665 (N_26665,N_25608,N_25788);
nor U26666 (N_26666,N_25581,N_25878);
nor U26667 (N_26667,N_25401,N_25150);
and U26668 (N_26668,N_25554,N_25071);
or U26669 (N_26669,N_25079,N_25322);
or U26670 (N_26670,N_25664,N_25073);
nand U26671 (N_26671,N_25956,N_25303);
nor U26672 (N_26672,N_25269,N_25789);
and U26673 (N_26673,N_25443,N_25601);
and U26674 (N_26674,N_25597,N_25544);
nand U26675 (N_26675,N_25242,N_25563);
and U26676 (N_26676,N_25184,N_25217);
and U26677 (N_26677,N_25030,N_25682);
nor U26678 (N_26678,N_25083,N_25817);
and U26679 (N_26679,N_25241,N_25354);
nand U26680 (N_26680,N_25821,N_25137);
nor U26681 (N_26681,N_25962,N_25258);
nand U26682 (N_26682,N_25286,N_25078);
nor U26683 (N_26683,N_25546,N_25290);
and U26684 (N_26684,N_25925,N_25728);
and U26685 (N_26685,N_25438,N_25619);
and U26686 (N_26686,N_25650,N_25340);
or U26687 (N_26687,N_25160,N_25176);
or U26688 (N_26688,N_25936,N_25543);
nor U26689 (N_26689,N_25570,N_25710);
nor U26690 (N_26690,N_25514,N_25518);
xnor U26691 (N_26691,N_25595,N_25387);
and U26692 (N_26692,N_25019,N_25487);
nor U26693 (N_26693,N_25708,N_25084);
and U26694 (N_26694,N_25544,N_25166);
nand U26695 (N_26695,N_25166,N_25167);
nand U26696 (N_26696,N_25619,N_25061);
or U26697 (N_26697,N_25172,N_25679);
and U26698 (N_26698,N_25258,N_25097);
nor U26699 (N_26699,N_25624,N_25321);
or U26700 (N_26700,N_25956,N_25094);
and U26701 (N_26701,N_25890,N_25810);
nand U26702 (N_26702,N_25759,N_25557);
nor U26703 (N_26703,N_25656,N_25102);
and U26704 (N_26704,N_25083,N_25815);
or U26705 (N_26705,N_25223,N_25834);
nor U26706 (N_26706,N_25186,N_25076);
or U26707 (N_26707,N_25115,N_25432);
nand U26708 (N_26708,N_25668,N_25899);
and U26709 (N_26709,N_25609,N_25463);
nand U26710 (N_26710,N_25456,N_25461);
nand U26711 (N_26711,N_25335,N_25814);
xnor U26712 (N_26712,N_25019,N_25721);
nand U26713 (N_26713,N_25003,N_25949);
and U26714 (N_26714,N_25437,N_25648);
nand U26715 (N_26715,N_25701,N_25327);
and U26716 (N_26716,N_25836,N_25417);
xor U26717 (N_26717,N_25009,N_25467);
or U26718 (N_26718,N_25085,N_25947);
xor U26719 (N_26719,N_25821,N_25185);
or U26720 (N_26720,N_25743,N_25750);
xnor U26721 (N_26721,N_25035,N_25969);
or U26722 (N_26722,N_25518,N_25094);
xor U26723 (N_26723,N_25680,N_25668);
and U26724 (N_26724,N_25031,N_25068);
xnor U26725 (N_26725,N_25890,N_25649);
or U26726 (N_26726,N_25267,N_25918);
xor U26727 (N_26727,N_25864,N_25423);
or U26728 (N_26728,N_25347,N_25575);
or U26729 (N_26729,N_25912,N_25293);
and U26730 (N_26730,N_25983,N_25648);
nand U26731 (N_26731,N_25390,N_25059);
and U26732 (N_26732,N_25855,N_25866);
and U26733 (N_26733,N_25374,N_25411);
nand U26734 (N_26734,N_25882,N_25241);
or U26735 (N_26735,N_25162,N_25264);
nand U26736 (N_26736,N_25100,N_25575);
nor U26737 (N_26737,N_25535,N_25863);
nand U26738 (N_26738,N_25714,N_25946);
or U26739 (N_26739,N_25676,N_25236);
or U26740 (N_26740,N_25032,N_25221);
nor U26741 (N_26741,N_25794,N_25995);
or U26742 (N_26742,N_25913,N_25940);
nor U26743 (N_26743,N_25149,N_25341);
and U26744 (N_26744,N_25334,N_25689);
xnor U26745 (N_26745,N_25914,N_25252);
and U26746 (N_26746,N_25860,N_25636);
nand U26747 (N_26747,N_25461,N_25125);
nor U26748 (N_26748,N_25242,N_25182);
and U26749 (N_26749,N_25955,N_25671);
or U26750 (N_26750,N_25172,N_25382);
and U26751 (N_26751,N_25101,N_25256);
nand U26752 (N_26752,N_25539,N_25525);
nor U26753 (N_26753,N_25603,N_25215);
nand U26754 (N_26754,N_25783,N_25790);
nor U26755 (N_26755,N_25593,N_25693);
or U26756 (N_26756,N_25513,N_25949);
or U26757 (N_26757,N_25938,N_25167);
xor U26758 (N_26758,N_25971,N_25758);
nand U26759 (N_26759,N_25343,N_25321);
nand U26760 (N_26760,N_25341,N_25955);
and U26761 (N_26761,N_25240,N_25312);
nor U26762 (N_26762,N_25643,N_25007);
nand U26763 (N_26763,N_25191,N_25272);
xor U26764 (N_26764,N_25703,N_25244);
and U26765 (N_26765,N_25550,N_25377);
nor U26766 (N_26766,N_25132,N_25741);
or U26767 (N_26767,N_25808,N_25070);
or U26768 (N_26768,N_25102,N_25163);
or U26769 (N_26769,N_25976,N_25977);
nand U26770 (N_26770,N_25796,N_25087);
nor U26771 (N_26771,N_25204,N_25034);
and U26772 (N_26772,N_25076,N_25956);
nand U26773 (N_26773,N_25028,N_25868);
and U26774 (N_26774,N_25817,N_25102);
nand U26775 (N_26775,N_25362,N_25841);
xor U26776 (N_26776,N_25612,N_25426);
nand U26777 (N_26777,N_25834,N_25950);
nand U26778 (N_26778,N_25025,N_25399);
nor U26779 (N_26779,N_25905,N_25178);
or U26780 (N_26780,N_25987,N_25018);
xor U26781 (N_26781,N_25033,N_25405);
xnor U26782 (N_26782,N_25590,N_25054);
or U26783 (N_26783,N_25325,N_25493);
nor U26784 (N_26784,N_25734,N_25356);
and U26785 (N_26785,N_25931,N_25641);
or U26786 (N_26786,N_25524,N_25420);
or U26787 (N_26787,N_25647,N_25079);
nor U26788 (N_26788,N_25643,N_25271);
or U26789 (N_26789,N_25306,N_25019);
or U26790 (N_26790,N_25458,N_25482);
nand U26791 (N_26791,N_25084,N_25590);
xnor U26792 (N_26792,N_25605,N_25491);
xnor U26793 (N_26793,N_25222,N_25556);
nor U26794 (N_26794,N_25452,N_25846);
nor U26795 (N_26795,N_25030,N_25572);
nand U26796 (N_26796,N_25481,N_25450);
nand U26797 (N_26797,N_25548,N_25920);
xor U26798 (N_26798,N_25255,N_25525);
xor U26799 (N_26799,N_25192,N_25274);
xor U26800 (N_26800,N_25718,N_25919);
nor U26801 (N_26801,N_25967,N_25509);
nand U26802 (N_26802,N_25457,N_25127);
nor U26803 (N_26803,N_25883,N_25978);
nor U26804 (N_26804,N_25060,N_25927);
xnor U26805 (N_26805,N_25396,N_25282);
nor U26806 (N_26806,N_25588,N_25855);
nor U26807 (N_26807,N_25184,N_25883);
xnor U26808 (N_26808,N_25630,N_25119);
and U26809 (N_26809,N_25193,N_25851);
nor U26810 (N_26810,N_25394,N_25585);
xnor U26811 (N_26811,N_25163,N_25123);
or U26812 (N_26812,N_25249,N_25446);
nor U26813 (N_26813,N_25740,N_25485);
nor U26814 (N_26814,N_25479,N_25672);
nor U26815 (N_26815,N_25673,N_25701);
nor U26816 (N_26816,N_25573,N_25025);
xor U26817 (N_26817,N_25102,N_25678);
and U26818 (N_26818,N_25949,N_25102);
xor U26819 (N_26819,N_25848,N_25484);
nor U26820 (N_26820,N_25452,N_25992);
nor U26821 (N_26821,N_25593,N_25955);
and U26822 (N_26822,N_25171,N_25206);
nand U26823 (N_26823,N_25413,N_25634);
or U26824 (N_26824,N_25767,N_25958);
or U26825 (N_26825,N_25585,N_25471);
nor U26826 (N_26826,N_25729,N_25990);
and U26827 (N_26827,N_25545,N_25334);
nor U26828 (N_26828,N_25758,N_25773);
and U26829 (N_26829,N_25340,N_25995);
nor U26830 (N_26830,N_25626,N_25062);
nand U26831 (N_26831,N_25895,N_25348);
and U26832 (N_26832,N_25710,N_25056);
xor U26833 (N_26833,N_25446,N_25040);
xnor U26834 (N_26834,N_25427,N_25809);
nand U26835 (N_26835,N_25328,N_25832);
xnor U26836 (N_26836,N_25529,N_25330);
nor U26837 (N_26837,N_25011,N_25904);
xor U26838 (N_26838,N_25121,N_25462);
nor U26839 (N_26839,N_25585,N_25774);
and U26840 (N_26840,N_25885,N_25226);
and U26841 (N_26841,N_25907,N_25492);
nand U26842 (N_26842,N_25542,N_25767);
nor U26843 (N_26843,N_25045,N_25971);
nand U26844 (N_26844,N_25084,N_25476);
xnor U26845 (N_26845,N_25807,N_25927);
nor U26846 (N_26846,N_25720,N_25605);
nand U26847 (N_26847,N_25501,N_25974);
or U26848 (N_26848,N_25210,N_25798);
nand U26849 (N_26849,N_25578,N_25036);
nand U26850 (N_26850,N_25362,N_25785);
or U26851 (N_26851,N_25162,N_25573);
or U26852 (N_26852,N_25686,N_25082);
xnor U26853 (N_26853,N_25186,N_25374);
and U26854 (N_26854,N_25951,N_25015);
or U26855 (N_26855,N_25289,N_25500);
xor U26856 (N_26856,N_25188,N_25147);
and U26857 (N_26857,N_25522,N_25623);
nor U26858 (N_26858,N_25804,N_25254);
nor U26859 (N_26859,N_25315,N_25074);
nor U26860 (N_26860,N_25934,N_25123);
and U26861 (N_26861,N_25568,N_25658);
nor U26862 (N_26862,N_25116,N_25045);
xor U26863 (N_26863,N_25740,N_25784);
nor U26864 (N_26864,N_25841,N_25825);
nand U26865 (N_26865,N_25927,N_25554);
nand U26866 (N_26866,N_25119,N_25290);
xor U26867 (N_26867,N_25115,N_25687);
nor U26868 (N_26868,N_25754,N_25170);
nand U26869 (N_26869,N_25536,N_25754);
xnor U26870 (N_26870,N_25468,N_25208);
or U26871 (N_26871,N_25191,N_25149);
nand U26872 (N_26872,N_25993,N_25327);
xnor U26873 (N_26873,N_25127,N_25311);
xnor U26874 (N_26874,N_25394,N_25225);
nor U26875 (N_26875,N_25470,N_25810);
nor U26876 (N_26876,N_25523,N_25138);
nor U26877 (N_26877,N_25758,N_25300);
or U26878 (N_26878,N_25874,N_25615);
nand U26879 (N_26879,N_25495,N_25686);
or U26880 (N_26880,N_25610,N_25906);
nand U26881 (N_26881,N_25750,N_25056);
xnor U26882 (N_26882,N_25041,N_25833);
nand U26883 (N_26883,N_25852,N_25209);
nor U26884 (N_26884,N_25541,N_25467);
nand U26885 (N_26885,N_25367,N_25390);
xor U26886 (N_26886,N_25525,N_25724);
nand U26887 (N_26887,N_25513,N_25111);
nand U26888 (N_26888,N_25110,N_25831);
nor U26889 (N_26889,N_25481,N_25134);
or U26890 (N_26890,N_25881,N_25419);
and U26891 (N_26891,N_25205,N_25565);
nor U26892 (N_26892,N_25890,N_25372);
xor U26893 (N_26893,N_25356,N_25553);
xnor U26894 (N_26894,N_25806,N_25858);
xor U26895 (N_26895,N_25539,N_25306);
xor U26896 (N_26896,N_25643,N_25955);
or U26897 (N_26897,N_25208,N_25637);
xor U26898 (N_26898,N_25824,N_25205);
and U26899 (N_26899,N_25705,N_25533);
nor U26900 (N_26900,N_25371,N_25190);
and U26901 (N_26901,N_25172,N_25961);
xor U26902 (N_26902,N_25161,N_25381);
nand U26903 (N_26903,N_25272,N_25045);
and U26904 (N_26904,N_25622,N_25150);
xnor U26905 (N_26905,N_25274,N_25892);
or U26906 (N_26906,N_25245,N_25931);
or U26907 (N_26907,N_25377,N_25674);
nor U26908 (N_26908,N_25277,N_25167);
and U26909 (N_26909,N_25503,N_25668);
nand U26910 (N_26910,N_25974,N_25235);
xnor U26911 (N_26911,N_25855,N_25365);
xnor U26912 (N_26912,N_25676,N_25636);
or U26913 (N_26913,N_25930,N_25625);
or U26914 (N_26914,N_25642,N_25964);
and U26915 (N_26915,N_25921,N_25564);
nor U26916 (N_26916,N_25229,N_25822);
xnor U26917 (N_26917,N_25836,N_25005);
and U26918 (N_26918,N_25776,N_25112);
or U26919 (N_26919,N_25744,N_25370);
xor U26920 (N_26920,N_25976,N_25172);
and U26921 (N_26921,N_25415,N_25602);
nand U26922 (N_26922,N_25638,N_25671);
nor U26923 (N_26923,N_25955,N_25818);
xnor U26924 (N_26924,N_25392,N_25724);
and U26925 (N_26925,N_25253,N_25387);
and U26926 (N_26926,N_25660,N_25975);
xor U26927 (N_26927,N_25732,N_25971);
nand U26928 (N_26928,N_25817,N_25609);
nand U26929 (N_26929,N_25075,N_25627);
nand U26930 (N_26930,N_25458,N_25411);
xnor U26931 (N_26931,N_25963,N_25887);
or U26932 (N_26932,N_25552,N_25405);
nor U26933 (N_26933,N_25098,N_25616);
xnor U26934 (N_26934,N_25534,N_25175);
or U26935 (N_26935,N_25400,N_25884);
nand U26936 (N_26936,N_25865,N_25550);
nor U26937 (N_26937,N_25884,N_25055);
nand U26938 (N_26938,N_25781,N_25664);
nand U26939 (N_26939,N_25079,N_25403);
and U26940 (N_26940,N_25479,N_25382);
xor U26941 (N_26941,N_25652,N_25759);
and U26942 (N_26942,N_25021,N_25719);
and U26943 (N_26943,N_25952,N_25681);
xnor U26944 (N_26944,N_25806,N_25908);
nor U26945 (N_26945,N_25347,N_25921);
or U26946 (N_26946,N_25891,N_25757);
and U26947 (N_26947,N_25378,N_25728);
nor U26948 (N_26948,N_25875,N_25428);
nand U26949 (N_26949,N_25741,N_25260);
and U26950 (N_26950,N_25942,N_25423);
nand U26951 (N_26951,N_25268,N_25736);
nor U26952 (N_26952,N_25102,N_25838);
and U26953 (N_26953,N_25691,N_25975);
nor U26954 (N_26954,N_25365,N_25746);
or U26955 (N_26955,N_25110,N_25542);
and U26956 (N_26956,N_25589,N_25583);
and U26957 (N_26957,N_25084,N_25491);
nand U26958 (N_26958,N_25691,N_25891);
and U26959 (N_26959,N_25055,N_25079);
or U26960 (N_26960,N_25991,N_25338);
or U26961 (N_26961,N_25568,N_25931);
nand U26962 (N_26962,N_25274,N_25632);
nor U26963 (N_26963,N_25589,N_25369);
or U26964 (N_26964,N_25235,N_25211);
nand U26965 (N_26965,N_25950,N_25302);
nand U26966 (N_26966,N_25466,N_25418);
or U26967 (N_26967,N_25209,N_25721);
xor U26968 (N_26968,N_25952,N_25130);
or U26969 (N_26969,N_25176,N_25110);
xor U26970 (N_26970,N_25164,N_25984);
nand U26971 (N_26971,N_25971,N_25322);
nand U26972 (N_26972,N_25379,N_25201);
and U26973 (N_26973,N_25049,N_25669);
xor U26974 (N_26974,N_25666,N_25044);
nor U26975 (N_26975,N_25976,N_25287);
nand U26976 (N_26976,N_25059,N_25381);
nand U26977 (N_26977,N_25507,N_25522);
nor U26978 (N_26978,N_25225,N_25263);
or U26979 (N_26979,N_25314,N_25567);
nor U26980 (N_26980,N_25512,N_25309);
nor U26981 (N_26981,N_25205,N_25089);
nor U26982 (N_26982,N_25637,N_25994);
nor U26983 (N_26983,N_25571,N_25934);
xnor U26984 (N_26984,N_25939,N_25141);
or U26985 (N_26985,N_25809,N_25504);
or U26986 (N_26986,N_25234,N_25726);
and U26987 (N_26987,N_25789,N_25676);
nand U26988 (N_26988,N_25172,N_25124);
nand U26989 (N_26989,N_25637,N_25615);
nor U26990 (N_26990,N_25937,N_25854);
and U26991 (N_26991,N_25079,N_25344);
nand U26992 (N_26992,N_25282,N_25313);
nor U26993 (N_26993,N_25016,N_25544);
nand U26994 (N_26994,N_25896,N_25521);
nor U26995 (N_26995,N_25434,N_25552);
nand U26996 (N_26996,N_25444,N_25431);
or U26997 (N_26997,N_25488,N_25550);
or U26998 (N_26998,N_25087,N_25620);
nor U26999 (N_26999,N_25447,N_25207);
nor U27000 (N_27000,N_26468,N_26105);
or U27001 (N_27001,N_26632,N_26529);
nor U27002 (N_27002,N_26354,N_26482);
and U27003 (N_27003,N_26780,N_26146);
or U27004 (N_27004,N_26211,N_26360);
or U27005 (N_27005,N_26807,N_26194);
or U27006 (N_27006,N_26478,N_26302);
nor U27007 (N_27007,N_26594,N_26068);
and U27008 (N_27008,N_26984,N_26810);
or U27009 (N_27009,N_26580,N_26481);
nor U27010 (N_27010,N_26473,N_26367);
xor U27011 (N_27011,N_26329,N_26259);
nor U27012 (N_27012,N_26326,N_26791);
nor U27013 (N_27013,N_26823,N_26287);
nand U27014 (N_27014,N_26042,N_26066);
or U27015 (N_27015,N_26979,N_26218);
xnor U27016 (N_27016,N_26988,N_26583);
xor U27017 (N_27017,N_26688,N_26362);
nor U27018 (N_27018,N_26390,N_26880);
nor U27019 (N_27019,N_26512,N_26395);
and U27020 (N_27020,N_26852,N_26694);
nand U27021 (N_27021,N_26322,N_26845);
and U27022 (N_27022,N_26489,N_26802);
xor U27023 (N_27023,N_26531,N_26461);
xnor U27024 (N_27024,N_26051,N_26808);
and U27025 (N_27025,N_26806,N_26956);
and U27026 (N_27026,N_26117,N_26497);
or U27027 (N_27027,N_26408,N_26556);
nand U27028 (N_27028,N_26385,N_26515);
xnor U27029 (N_27029,N_26865,N_26714);
nor U27030 (N_27030,N_26924,N_26667);
nor U27031 (N_27031,N_26587,N_26566);
nand U27032 (N_27032,N_26371,N_26022);
nor U27033 (N_27033,N_26909,N_26342);
xnor U27034 (N_27034,N_26450,N_26937);
nand U27035 (N_27035,N_26129,N_26162);
nand U27036 (N_27036,N_26666,N_26401);
xor U27037 (N_27037,N_26402,N_26631);
nand U27038 (N_27038,N_26809,N_26319);
or U27039 (N_27039,N_26745,N_26555);
nor U27040 (N_27040,N_26538,N_26734);
or U27041 (N_27041,N_26870,N_26544);
or U27042 (N_27042,N_26707,N_26421);
nand U27043 (N_27043,N_26436,N_26103);
and U27044 (N_27044,N_26973,N_26641);
or U27045 (N_27045,N_26801,N_26673);
xnor U27046 (N_27046,N_26081,N_26908);
nor U27047 (N_27047,N_26837,N_26996);
xnor U27048 (N_27048,N_26149,N_26676);
or U27049 (N_27049,N_26586,N_26494);
xor U27050 (N_27050,N_26256,N_26364);
and U27051 (N_27051,N_26039,N_26994);
nor U27052 (N_27052,N_26127,N_26411);
or U27053 (N_27053,N_26835,N_26934);
xnor U27054 (N_27054,N_26295,N_26179);
nand U27055 (N_27055,N_26240,N_26314);
or U27056 (N_27056,N_26917,N_26422);
or U27057 (N_27057,N_26704,N_26552);
xor U27058 (N_27058,N_26783,N_26310);
or U27059 (N_27059,N_26141,N_26742);
or U27060 (N_27060,N_26782,N_26236);
nor U27061 (N_27061,N_26569,N_26217);
nand U27062 (N_27062,N_26004,N_26346);
xnor U27063 (N_27063,N_26132,N_26751);
and U27064 (N_27064,N_26718,N_26486);
nor U27065 (N_27065,N_26216,N_26678);
or U27066 (N_27066,N_26978,N_26206);
nor U27067 (N_27067,N_26001,N_26100);
or U27068 (N_27068,N_26311,N_26359);
and U27069 (N_27069,N_26156,N_26998);
xor U27070 (N_27070,N_26054,N_26763);
nand U27071 (N_27071,N_26611,N_26230);
or U27072 (N_27072,N_26774,N_26093);
nand U27073 (N_27073,N_26237,N_26091);
or U27074 (N_27074,N_26281,N_26242);
nand U27075 (N_27075,N_26062,N_26625);
xor U27076 (N_27076,N_26510,N_26831);
and U27077 (N_27077,N_26970,N_26733);
or U27078 (N_27078,N_26374,N_26854);
or U27079 (N_27079,N_26285,N_26916);
nand U27080 (N_27080,N_26710,N_26928);
nand U27081 (N_27081,N_26317,N_26316);
nand U27082 (N_27082,N_26511,N_26993);
and U27083 (N_27083,N_26543,N_26500);
nand U27084 (N_27084,N_26768,N_26833);
or U27085 (N_27085,N_26366,N_26198);
nor U27086 (N_27086,N_26106,N_26098);
and U27087 (N_27087,N_26679,N_26223);
and U27088 (N_27088,N_26723,N_26219);
nor U27089 (N_27089,N_26116,N_26212);
nor U27090 (N_27090,N_26257,N_26244);
xor U27091 (N_27091,N_26448,N_26907);
nand U27092 (N_27092,N_26588,N_26112);
nand U27093 (N_27093,N_26377,N_26392);
xor U27094 (N_27094,N_26172,N_26487);
xnor U27095 (N_27095,N_26744,N_26614);
and U27096 (N_27096,N_26672,N_26071);
or U27097 (N_27097,N_26128,N_26232);
and U27098 (N_27098,N_26581,N_26405);
xnor U27099 (N_27099,N_26070,N_26031);
nor U27100 (N_27100,N_26797,N_26905);
nor U27101 (N_27101,N_26592,N_26509);
or U27102 (N_27102,N_26739,N_26847);
or U27103 (N_27103,N_26125,N_26102);
and U27104 (N_27104,N_26189,N_26557);
nor U27105 (N_27105,N_26372,N_26624);
nand U27106 (N_27106,N_26365,N_26947);
xor U27107 (N_27107,N_26861,N_26019);
or U27108 (N_27108,N_26079,N_26178);
or U27109 (N_27109,N_26024,N_26113);
nand U27110 (N_27110,N_26550,N_26938);
or U27111 (N_27111,N_26469,N_26668);
nor U27112 (N_27112,N_26502,N_26275);
xnor U27113 (N_27113,N_26191,N_26406);
nand U27114 (N_27114,N_26139,N_26018);
xnor U27115 (N_27115,N_26029,N_26058);
and U27116 (N_27116,N_26685,N_26902);
nand U27117 (N_27117,N_26415,N_26787);
nand U27118 (N_27118,N_26437,N_26789);
xor U27119 (N_27119,N_26349,N_26276);
and U27120 (N_27120,N_26130,N_26589);
nor U27121 (N_27121,N_26653,N_26353);
nand U27122 (N_27122,N_26052,N_26386);
xor U27123 (N_27123,N_26951,N_26866);
nor U27124 (N_27124,N_26944,N_26331);
or U27125 (N_27125,N_26239,N_26897);
nor U27126 (N_27126,N_26063,N_26452);
nor U27127 (N_27127,N_26060,N_26713);
nor U27128 (N_27128,N_26300,N_26357);
or U27129 (N_27129,N_26496,N_26968);
nor U27130 (N_27130,N_26137,N_26930);
or U27131 (N_27131,N_26634,N_26110);
xnor U27132 (N_27132,N_26380,N_26278);
or U27133 (N_27133,N_26161,N_26757);
xor U27134 (N_27134,N_26165,N_26090);
and U27135 (N_27135,N_26343,N_26306);
and U27136 (N_27136,N_26006,N_26335);
and U27137 (N_27137,N_26350,N_26023);
xor U27138 (N_27138,N_26047,N_26115);
nor U27139 (N_27139,N_26148,N_26345);
and U27140 (N_27140,N_26684,N_26182);
or U27141 (N_27141,N_26279,N_26712);
nor U27142 (N_27142,N_26779,N_26107);
and U27143 (N_27143,N_26792,N_26554);
xor U27144 (N_27144,N_26197,N_26072);
nor U27145 (N_27145,N_26417,N_26088);
nand U27146 (N_27146,N_26546,N_26518);
nor U27147 (N_27147,N_26010,N_26294);
and U27148 (N_27148,N_26728,N_26860);
xnor U27149 (N_27149,N_26681,N_26598);
nor U27150 (N_27150,N_26635,N_26123);
or U27151 (N_27151,N_26633,N_26076);
and U27152 (N_27152,N_26756,N_26457);
and U27153 (N_27153,N_26073,N_26725);
and U27154 (N_27154,N_26389,N_26126);
or U27155 (N_27155,N_26827,N_26654);
nand U27156 (N_27156,N_26629,N_26307);
nor U27157 (N_27157,N_26894,N_26766);
and U27158 (N_27158,N_26596,N_26521);
nor U27159 (N_27159,N_26409,N_26608);
nand U27160 (N_27160,N_26025,N_26134);
and U27161 (N_27161,N_26332,N_26991);
nor U27162 (N_27162,N_26449,N_26637);
xor U27163 (N_27163,N_26009,N_26454);
nand U27164 (N_27164,N_26948,N_26315);
nand U27165 (N_27165,N_26539,N_26412);
nand U27166 (N_27166,N_26690,N_26325);
and U27167 (N_27167,N_26950,N_26677);
nand U27168 (N_27168,N_26087,N_26826);
xor U27169 (N_27169,N_26579,N_26922);
xor U27170 (N_27170,N_26561,N_26876);
or U27171 (N_27171,N_26292,N_26208);
nor U27172 (N_27172,N_26460,N_26818);
nand U27173 (N_27173,N_26328,N_26157);
and U27174 (N_27174,N_26413,N_26083);
nand U27175 (N_27175,N_26699,N_26923);
and U27176 (N_27176,N_26946,N_26485);
and U27177 (N_27177,N_26470,N_26442);
or U27178 (N_27178,N_26693,N_26272);
and U27179 (N_27179,N_26958,N_26656);
or U27180 (N_27180,N_26160,N_26504);
nor U27181 (N_27181,N_26935,N_26565);
or U27182 (N_27182,N_26921,N_26659);
nor U27183 (N_27183,N_26007,N_26778);
and U27184 (N_27184,N_26501,N_26361);
or U27185 (N_27185,N_26424,N_26868);
and U27186 (N_27186,N_26691,N_26857);
xor U27187 (N_27187,N_26444,N_26636);
xor U27188 (N_27188,N_26145,N_26288);
xor U27189 (N_27189,N_26892,N_26174);
xor U27190 (N_27190,N_26247,N_26974);
and U27191 (N_27191,N_26597,N_26534);
nor U27192 (N_27192,N_26709,N_26265);
nor U27193 (N_27193,N_26798,N_26432);
nor U27194 (N_27194,N_26604,N_26225);
nor U27195 (N_27195,N_26983,N_26812);
or U27196 (N_27196,N_26525,N_26570);
nor U27197 (N_27197,N_26911,N_26784);
and U27198 (N_27198,N_26114,N_26925);
nor U27199 (N_27199,N_26159,N_26945);
nand U27200 (N_27200,N_26730,N_26906);
nand U27201 (N_27201,N_26686,N_26423);
nand U27202 (N_27202,N_26879,N_26765);
xor U27203 (N_27203,N_26755,N_26615);
nor U27204 (N_27204,N_26607,N_26255);
nand U27205 (N_27205,N_26170,N_26560);
xnor U27206 (N_27206,N_26788,N_26612);
nor U27207 (N_27207,N_26736,N_26193);
nor U27208 (N_27208,N_26492,N_26877);
or U27209 (N_27209,N_26942,N_26726);
nor U27210 (N_27210,N_26936,N_26832);
nor U27211 (N_27211,N_26375,N_26391);
xnor U27212 (N_27212,N_26456,N_26324);
or U27213 (N_27213,N_26548,N_26347);
or U27214 (N_27214,N_26972,N_26853);
nand U27215 (N_27215,N_26841,N_26542);
nand U27216 (N_27216,N_26344,N_26234);
or U27217 (N_27217,N_26507,N_26228);
xor U27218 (N_27218,N_26644,N_26601);
nand U27219 (N_27219,N_26387,N_26416);
and U27220 (N_27220,N_26277,N_26049);
or U27221 (N_27221,N_26772,N_26889);
xnor U27222 (N_27222,N_26817,N_26533);
nand U27223 (N_27223,N_26671,N_26382);
or U27224 (N_27224,N_26439,N_26011);
nand U27225 (N_27225,N_26800,N_26167);
or U27226 (N_27226,N_26138,N_26397);
or U27227 (N_27227,N_26793,N_26171);
and U27228 (N_27228,N_26702,N_26005);
and U27229 (N_27229,N_26927,N_26410);
xor U27230 (N_27230,N_26796,N_26855);
and U27231 (N_27231,N_26235,N_26899);
nand U27232 (N_27232,N_26075,N_26394);
nor U27233 (N_27233,N_26041,N_26836);
or U27234 (N_27234,N_26535,N_26252);
nor U27235 (N_27235,N_26708,N_26697);
nand U27236 (N_27236,N_26250,N_26333);
xnor U27237 (N_27237,N_26192,N_26645);
or U27238 (N_27238,N_26484,N_26888);
xor U27239 (N_27239,N_26213,N_26195);
xnor U27240 (N_27240,N_26616,N_26163);
and U27241 (N_27241,N_26229,N_26519);
nor U27242 (N_27242,N_26269,N_26603);
xor U27243 (N_27243,N_26600,N_26465);
nor U27244 (N_27244,N_26312,N_26867);
nand U27245 (N_27245,N_26263,N_26819);
nand U27246 (N_27246,N_26053,N_26627);
and U27247 (N_27247,N_26573,N_26186);
xnor U27248 (N_27248,N_26069,N_26433);
and U27249 (N_27249,N_26981,N_26050);
nor U27250 (N_27250,N_26602,N_26610);
and U27251 (N_27251,N_26582,N_26746);
xor U27252 (N_27252,N_26918,N_26190);
xor U27253 (N_27253,N_26843,N_26786);
xor U27254 (N_27254,N_26522,N_26963);
nor U27255 (N_27255,N_26418,N_26683);
or U27256 (N_27256,N_26932,N_26910);
and U27257 (N_27257,N_26527,N_26403);
and U27258 (N_27258,N_26297,N_26856);
xnor U27259 (N_27259,N_26447,N_26222);
xnor U27260 (N_27260,N_26077,N_26620);
nor U27261 (N_27261,N_26874,N_26274);
nand U27262 (N_27262,N_26997,N_26578);
nor U27263 (N_27263,N_26859,N_26204);
xnor U27264 (N_27264,N_26400,N_26987);
nor U27265 (N_27265,N_26962,N_26655);
nand U27266 (N_27266,N_26096,N_26455);
xnor U27267 (N_27267,N_26133,N_26722);
xnor U27268 (N_27268,N_26036,N_26663);
xnor U27269 (N_27269,N_26441,N_26308);
nor U27270 (N_27270,N_26358,N_26131);
and U27271 (N_27271,N_26176,N_26082);
xor U27272 (N_27272,N_26313,N_26305);
xor U27273 (N_27273,N_26609,N_26551);
or U27274 (N_27274,N_26327,N_26743);
nand U27275 (N_27275,N_26642,N_26187);
or U27276 (N_27276,N_26919,N_26532);
nand U27277 (N_27277,N_26985,N_26270);
and U27278 (N_27278,N_26399,N_26640);
nor U27279 (N_27279,N_26330,N_26245);
xnor U27280 (N_27280,N_26903,N_26593);
xor U27281 (N_27281,N_26296,N_26762);
xor U27282 (N_27282,N_26619,N_26982);
xnor U27283 (N_27283,N_26828,N_26754);
xnor U27284 (N_27284,N_26700,N_26846);
xnor U27285 (N_27285,N_26687,N_26526);
and U27286 (N_27286,N_26658,N_26420);
nand U27287 (N_27287,N_26341,N_26630);
and U27288 (N_27288,N_26046,N_26271);
nor U27289 (N_27289,N_26508,N_26283);
and U27290 (N_27290,N_26967,N_26776);
or U27291 (N_27291,N_26089,N_26435);
or U27292 (N_27292,N_26184,N_26724);
or U27293 (N_27293,N_26811,N_26748);
nor U27294 (N_27294,N_26825,N_26196);
nor U27295 (N_27295,N_26266,N_26258);
nor U27296 (N_27296,N_26995,N_26241);
nand U27297 (N_27297,N_26621,N_26506);
nand U27298 (N_27298,N_26430,N_26251);
xnor U27299 (N_27299,N_26384,N_26398);
nand U27300 (N_27300,N_26605,N_26839);
nor U27301 (N_27301,N_26498,N_26085);
and U27302 (N_27302,N_26689,N_26254);
nor U27303 (N_27303,N_26849,N_26056);
nand U27304 (N_27304,N_26564,N_26503);
and U27305 (N_27305,N_26805,N_26002);
nor U27306 (N_27306,N_26393,N_26021);
and U27307 (N_27307,N_26568,N_26261);
nand U27308 (N_27308,N_26080,N_26540);
and U27309 (N_27309,N_26092,N_26822);
xor U27310 (N_27310,N_26177,N_26639);
xnor U27311 (N_27311,N_26992,N_26871);
and U27312 (N_27312,N_26559,N_26940);
nand U27313 (N_27313,N_26523,N_26061);
and U27314 (N_27314,N_26169,N_26652);
nand U27315 (N_27315,N_26553,N_26142);
or U27316 (N_27316,N_26869,N_26154);
nor U27317 (N_27317,N_26858,N_26851);
or U27318 (N_27318,N_26576,N_26719);
xor U27319 (N_27319,N_26872,N_26363);
nand U27320 (N_27320,N_26571,N_26680);
xor U27321 (N_27321,N_26013,N_26370);
nor U27322 (N_27322,N_26661,N_26558);
xor U27323 (N_27323,N_26721,N_26814);
and U27324 (N_27324,N_26065,N_26595);
nand U27325 (N_27325,N_26717,N_26108);
nand U27326 (N_27326,N_26959,N_26971);
nand U27327 (N_27327,N_26122,N_26221);
or U27328 (N_27328,N_26750,N_26084);
nor U27329 (N_27329,N_26696,N_26731);
and U27330 (N_27330,N_26882,N_26181);
nor U27331 (N_27331,N_26824,N_26650);
and U27332 (N_27332,N_26379,N_26900);
nand U27333 (N_27333,N_26121,N_26505);
or U27334 (N_27334,N_26862,N_26233);
or U27335 (N_27335,N_26647,N_26622);
or U27336 (N_27336,N_26451,N_26960);
nor U27337 (N_27337,N_26381,N_26623);
nor U27338 (N_27338,N_26887,N_26585);
nand U27339 (N_27339,N_26976,N_26286);
or U27340 (N_27340,N_26590,N_26760);
xor U27341 (N_27341,N_26040,N_26443);
and U27342 (N_27342,N_26574,N_26957);
xor U27343 (N_27343,N_26803,N_26155);
xor U27344 (N_27344,N_26617,N_26705);
nor U27345 (N_27345,N_26057,N_26878);
or U27346 (N_27346,N_26434,N_26769);
and U27347 (N_27347,N_26419,N_26537);
nor U27348 (N_27348,N_26729,N_26210);
and U27349 (N_27349,N_26273,N_26291);
and U27350 (N_27350,N_26698,N_26429);
nor U27351 (N_27351,N_26764,N_26203);
nand U27352 (N_27352,N_26290,N_26584);
nor U27353 (N_27353,N_26830,N_26716);
nor U27354 (N_27354,N_26476,N_26144);
nand U27355 (N_27355,N_26220,N_26323);
and U27356 (N_27356,N_26920,N_26893);
xor U27357 (N_27357,N_26966,N_26701);
or U27358 (N_27358,N_26577,N_26513);
or U27359 (N_27359,N_26012,N_26111);
and U27360 (N_27360,N_26753,N_26901);
and U27361 (N_27361,N_26376,N_26086);
nor U27362 (N_27362,N_26912,N_26064);
nor U27363 (N_27363,N_26545,N_26915);
and U27364 (N_27364,N_26795,N_26665);
nand U27365 (N_27365,N_26166,N_26045);
xor U27366 (N_27366,N_26109,N_26599);
nand U27367 (N_27367,N_26474,N_26264);
nand U27368 (N_27368,N_26188,N_26767);
or U27369 (N_27369,N_26720,N_26775);
and U27370 (N_27370,N_26520,N_26575);
nand U27371 (N_27371,N_26741,N_26885);
nand U27372 (N_27372,N_26475,N_26883);
and U27373 (N_27373,N_26838,N_26675);
xor U27374 (N_27374,N_26334,N_26952);
and U27375 (N_27375,N_26933,N_26202);
or U27376 (N_27376,N_26850,N_26483);
nor U27377 (N_27377,N_26816,N_26896);
or U27378 (N_27378,N_26453,N_26758);
and U27379 (N_27379,N_26471,N_26977);
nor U27380 (N_27380,N_26227,N_26514);
xor U27381 (N_27381,N_26516,N_26340);
nor U27382 (N_27382,N_26821,N_26043);
or U27383 (N_27383,N_26248,N_26299);
xor U27384 (N_27384,N_26462,N_26136);
nor U27385 (N_27385,N_26549,N_26657);
and U27386 (N_27386,N_26185,N_26094);
nand U27387 (N_27387,N_26628,N_26955);
nand U27388 (N_27388,N_26695,N_26246);
nor U27389 (N_27389,N_26231,N_26711);
and U27390 (N_27390,N_26638,N_26014);
xor U27391 (N_27391,N_26033,N_26280);
and U27392 (N_27392,N_26355,N_26304);
and U27393 (N_27393,N_26648,N_26790);
xor U27394 (N_27394,N_26651,N_26268);
xor U27395 (N_27395,N_26794,N_26530);
nor U27396 (N_27396,N_26785,N_26613);
nand U27397 (N_27397,N_26941,N_26759);
nand U27398 (N_27398,N_26458,N_26238);
nor U27399 (N_27399,N_26591,N_26761);
or U27400 (N_27400,N_26426,N_26048);
xor U27401 (N_27401,N_26368,N_26017);
xnor U27402 (N_27402,N_26662,N_26243);
or U27403 (N_27403,N_26820,N_26175);
or U27404 (N_27404,N_26961,N_26727);
xnor U27405 (N_27405,N_26618,N_26173);
or U27406 (N_27406,N_26226,N_26431);
and U27407 (N_27407,N_26352,N_26044);
and U27408 (N_27408,N_26528,N_26369);
and U27409 (N_27409,N_26118,N_26032);
xnor U27410 (N_27410,N_26253,N_26493);
or U27411 (N_27411,N_26035,N_26477);
xnor U27412 (N_27412,N_26781,N_26151);
nor U27413 (N_27413,N_26964,N_26517);
xor U27414 (N_27414,N_26003,N_26873);
and U27415 (N_27415,N_26480,N_26337);
nand U27416 (N_27416,N_26224,N_26038);
nor U27417 (N_27417,N_26008,N_26124);
xnor U27418 (N_27418,N_26931,N_26703);
nor U27419 (N_27419,N_26886,N_26840);
nand U27420 (N_27420,N_26829,N_26104);
xnor U27421 (N_27421,N_26943,N_26881);
nand U27422 (N_27422,N_26267,N_26965);
xnor U27423 (N_27423,N_26459,N_26771);
nand U27424 (N_27424,N_26670,N_26309);
and U27425 (N_27425,N_26864,N_26143);
nand U27426 (N_27426,N_26562,N_26904);
nand U27427 (N_27427,N_26863,N_26135);
xor U27428 (N_27428,N_26318,N_26205);
xor U27429 (N_27429,N_26986,N_26301);
or U27430 (N_27430,N_26164,N_26438);
nor U27431 (N_27431,N_26692,N_26954);
xnor U27432 (N_27432,N_26740,N_26183);
or U27433 (N_27433,N_26078,N_26660);
or U27434 (N_27434,N_26463,N_26215);
and U27435 (N_27435,N_26715,N_26643);
or U27436 (N_27436,N_26491,N_26467);
xnor U27437 (N_27437,N_26199,N_26488);
xor U27438 (N_27438,N_26338,N_26207);
xnor U27439 (N_27439,N_26284,N_26844);
nand U27440 (N_27440,N_26773,N_26388);
nor U27441 (N_27441,N_26875,N_26034);
or U27442 (N_27442,N_26201,N_26348);
nand U27443 (N_27443,N_26152,N_26020);
or U27444 (N_27444,N_26752,N_26834);
nor U27445 (N_27445,N_26282,N_26214);
nand U27446 (N_27446,N_26848,N_26396);
or U27447 (N_27447,N_26799,N_26815);
or U27448 (N_27448,N_26262,N_26336);
xnor U27449 (N_27449,N_26339,N_26440);
nand U27450 (N_27450,N_26646,N_26898);
and U27451 (N_27451,N_26926,N_26298);
nand U27452 (N_27452,N_26466,N_26158);
or U27453 (N_27453,N_26674,N_26028);
and U27454 (N_27454,N_26737,N_26260);
nor U27455 (N_27455,N_26140,N_26321);
xnor U27456 (N_27456,N_26929,N_26682);
and U27457 (N_27457,N_26884,N_26074);
nand U27458 (N_27458,N_26027,N_26249);
xor U27459 (N_27459,N_26563,N_26969);
xnor U27460 (N_27460,N_26059,N_26425);
nand U27461 (N_27461,N_26567,N_26030);
xnor U27462 (N_27462,N_26572,N_26407);
and U27463 (N_27463,N_26464,N_26738);
xor U27464 (N_27464,N_26541,N_26939);
and U27465 (N_27465,N_26606,N_26891);
and U27466 (N_27466,N_26351,N_26289);
xor U27467 (N_27467,N_26320,N_26383);
nand U27468 (N_27468,N_26097,N_26949);
xor U27469 (N_27469,N_26747,N_26209);
xor U27470 (N_27470,N_26895,N_26649);
nor U27471 (N_27471,N_26414,N_26168);
and U27472 (N_27472,N_26180,N_26914);
nand U27473 (N_27473,N_26446,N_26055);
nand U27474 (N_27474,N_26524,N_26777);
nand U27475 (N_27475,N_26813,N_26953);
and U27476 (N_27476,N_26842,N_26999);
and U27477 (N_27477,N_26293,N_26479);
and U27478 (N_27478,N_26147,N_26373);
or U27479 (N_27479,N_26445,N_26095);
nor U27480 (N_27480,N_26153,N_26015);
nand U27481 (N_27481,N_26356,N_26890);
xnor U27482 (N_27482,N_26472,N_26990);
nor U27483 (N_27483,N_26101,N_26975);
nand U27484 (N_27484,N_26200,N_26989);
or U27485 (N_27485,N_26404,N_26016);
xnor U27486 (N_27486,N_26120,N_26303);
or U27487 (N_27487,N_26732,N_26000);
or U27488 (N_27488,N_26026,N_26378);
nor U27489 (N_27489,N_26547,N_26150);
and U27490 (N_27490,N_26626,N_26428);
or U27491 (N_27491,N_26119,N_26495);
xnor U27492 (N_27492,N_26913,N_26664);
and U27493 (N_27493,N_26536,N_26980);
nor U27494 (N_27494,N_26804,N_26749);
xnor U27495 (N_27495,N_26490,N_26067);
nand U27496 (N_27496,N_26770,N_26099);
and U27497 (N_27497,N_26499,N_26735);
xnor U27498 (N_27498,N_26427,N_26669);
nand U27499 (N_27499,N_26706,N_26037);
or U27500 (N_27500,N_26209,N_26694);
and U27501 (N_27501,N_26196,N_26256);
or U27502 (N_27502,N_26671,N_26933);
xnor U27503 (N_27503,N_26389,N_26199);
nor U27504 (N_27504,N_26865,N_26032);
nand U27505 (N_27505,N_26426,N_26661);
and U27506 (N_27506,N_26290,N_26561);
or U27507 (N_27507,N_26145,N_26066);
nand U27508 (N_27508,N_26727,N_26735);
or U27509 (N_27509,N_26288,N_26961);
or U27510 (N_27510,N_26219,N_26589);
and U27511 (N_27511,N_26505,N_26562);
xor U27512 (N_27512,N_26611,N_26071);
and U27513 (N_27513,N_26712,N_26016);
nor U27514 (N_27514,N_26339,N_26193);
nand U27515 (N_27515,N_26498,N_26339);
xnor U27516 (N_27516,N_26745,N_26039);
nand U27517 (N_27517,N_26432,N_26573);
xnor U27518 (N_27518,N_26001,N_26745);
and U27519 (N_27519,N_26062,N_26140);
nand U27520 (N_27520,N_26970,N_26434);
xnor U27521 (N_27521,N_26995,N_26538);
xor U27522 (N_27522,N_26982,N_26100);
or U27523 (N_27523,N_26014,N_26844);
nand U27524 (N_27524,N_26852,N_26323);
nand U27525 (N_27525,N_26859,N_26863);
nand U27526 (N_27526,N_26050,N_26293);
nor U27527 (N_27527,N_26425,N_26676);
nand U27528 (N_27528,N_26748,N_26062);
nor U27529 (N_27529,N_26387,N_26886);
and U27530 (N_27530,N_26380,N_26582);
or U27531 (N_27531,N_26707,N_26664);
and U27532 (N_27532,N_26926,N_26714);
nand U27533 (N_27533,N_26822,N_26428);
xor U27534 (N_27534,N_26242,N_26802);
xor U27535 (N_27535,N_26458,N_26560);
nand U27536 (N_27536,N_26858,N_26618);
and U27537 (N_27537,N_26696,N_26931);
and U27538 (N_27538,N_26187,N_26529);
xnor U27539 (N_27539,N_26055,N_26337);
xnor U27540 (N_27540,N_26896,N_26474);
and U27541 (N_27541,N_26417,N_26374);
nor U27542 (N_27542,N_26675,N_26070);
or U27543 (N_27543,N_26506,N_26937);
nor U27544 (N_27544,N_26633,N_26797);
nand U27545 (N_27545,N_26256,N_26347);
or U27546 (N_27546,N_26400,N_26346);
xor U27547 (N_27547,N_26745,N_26202);
xor U27548 (N_27548,N_26724,N_26650);
and U27549 (N_27549,N_26178,N_26978);
and U27550 (N_27550,N_26586,N_26195);
and U27551 (N_27551,N_26388,N_26739);
or U27552 (N_27552,N_26056,N_26391);
and U27553 (N_27553,N_26852,N_26977);
or U27554 (N_27554,N_26398,N_26276);
nand U27555 (N_27555,N_26530,N_26373);
xnor U27556 (N_27556,N_26995,N_26420);
and U27557 (N_27557,N_26925,N_26173);
nor U27558 (N_27558,N_26006,N_26849);
xnor U27559 (N_27559,N_26020,N_26051);
or U27560 (N_27560,N_26265,N_26832);
or U27561 (N_27561,N_26492,N_26332);
nand U27562 (N_27562,N_26183,N_26538);
or U27563 (N_27563,N_26575,N_26128);
nor U27564 (N_27564,N_26566,N_26025);
or U27565 (N_27565,N_26286,N_26015);
or U27566 (N_27566,N_26321,N_26474);
xor U27567 (N_27567,N_26249,N_26724);
nand U27568 (N_27568,N_26356,N_26729);
or U27569 (N_27569,N_26361,N_26042);
or U27570 (N_27570,N_26528,N_26374);
xnor U27571 (N_27571,N_26745,N_26809);
xnor U27572 (N_27572,N_26646,N_26608);
or U27573 (N_27573,N_26209,N_26318);
xnor U27574 (N_27574,N_26833,N_26877);
nand U27575 (N_27575,N_26419,N_26773);
or U27576 (N_27576,N_26108,N_26179);
xor U27577 (N_27577,N_26534,N_26056);
or U27578 (N_27578,N_26097,N_26244);
or U27579 (N_27579,N_26751,N_26675);
nor U27580 (N_27580,N_26968,N_26449);
or U27581 (N_27581,N_26636,N_26269);
or U27582 (N_27582,N_26696,N_26323);
xnor U27583 (N_27583,N_26587,N_26665);
nor U27584 (N_27584,N_26956,N_26606);
xor U27585 (N_27585,N_26526,N_26730);
or U27586 (N_27586,N_26316,N_26403);
or U27587 (N_27587,N_26359,N_26480);
and U27588 (N_27588,N_26662,N_26768);
xor U27589 (N_27589,N_26997,N_26989);
nor U27590 (N_27590,N_26147,N_26473);
nor U27591 (N_27591,N_26221,N_26126);
or U27592 (N_27592,N_26774,N_26262);
nor U27593 (N_27593,N_26233,N_26723);
and U27594 (N_27594,N_26987,N_26809);
or U27595 (N_27595,N_26994,N_26189);
nand U27596 (N_27596,N_26420,N_26044);
and U27597 (N_27597,N_26135,N_26817);
nor U27598 (N_27598,N_26019,N_26430);
or U27599 (N_27599,N_26269,N_26322);
nor U27600 (N_27600,N_26782,N_26621);
nor U27601 (N_27601,N_26251,N_26263);
and U27602 (N_27602,N_26130,N_26612);
and U27603 (N_27603,N_26751,N_26013);
nor U27604 (N_27604,N_26492,N_26128);
nand U27605 (N_27605,N_26318,N_26816);
xor U27606 (N_27606,N_26378,N_26551);
xor U27607 (N_27607,N_26325,N_26429);
or U27608 (N_27608,N_26174,N_26889);
xnor U27609 (N_27609,N_26367,N_26237);
nand U27610 (N_27610,N_26703,N_26125);
nand U27611 (N_27611,N_26540,N_26881);
nand U27612 (N_27612,N_26001,N_26737);
or U27613 (N_27613,N_26933,N_26737);
xor U27614 (N_27614,N_26359,N_26294);
and U27615 (N_27615,N_26125,N_26936);
xor U27616 (N_27616,N_26731,N_26290);
and U27617 (N_27617,N_26561,N_26452);
and U27618 (N_27618,N_26943,N_26949);
nor U27619 (N_27619,N_26860,N_26558);
or U27620 (N_27620,N_26241,N_26684);
or U27621 (N_27621,N_26690,N_26121);
nand U27622 (N_27622,N_26747,N_26056);
nand U27623 (N_27623,N_26054,N_26171);
and U27624 (N_27624,N_26149,N_26137);
and U27625 (N_27625,N_26524,N_26922);
and U27626 (N_27626,N_26314,N_26808);
nor U27627 (N_27627,N_26524,N_26785);
or U27628 (N_27628,N_26894,N_26558);
or U27629 (N_27629,N_26691,N_26607);
and U27630 (N_27630,N_26365,N_26803);
or U27631 (N_27631,N_26017,N_26553);
nor U27632 (N_27632,N_26103,N_26227);
nor U27633 (N_27633,N_26830,N_26101);
and U27634 (N_27634,N_26330,N_26576);
xor U27635 (N_27635,N_26742,N_26211);
or U27636 (N_27636,N_26256,N_26613);
and U27637 (N_27637,N_26467,N_26166);
nor U27638 (N_27638,N_26377,N_26308);
nand U27639 (N_27639,N_26890,N_26677);
or U27640 (N_27640,N_26399,N_26852);
xnor U27641 (N_27641,N_26964,N_26163);
and U27642 (N_27642,N_26085,N_26043);
or U27643 (N_27643,N_26236,N_26680);
and U27644 (N_27644,N_26572,N_26899);
nor U27645 (N_27645,N_26801,N_26233);
or U27646 (N_27646,N_26915,N_26638);
xor U27647 (N_27647,N_26383,N_26203);
nand U27648 (N_27648,N_26743,N_26118);
nor U27649 (N_27649,N_26555,N_26515);
nand U27650 (N_27650,N_26910,N_26393);
or U27651 (N_27651,N_26168,N_26079);
and U27652 (N_27652,N_26311,N_26173);
and U27653 (N_27653,N_26176,N_26341);
xnor U27654 (N_27654,N_26358,N_26175);
nor U27655 (N_27655,N_26806,N_26862);
nor U27656 (N_27656,N_26991,N_26344);
nand U27657 (N_27657,N_26247,N_26588);
xor U27658 (N_27658,N_26068,N_26643);
nor U27659 (N_27659,N_26638,N_26010);
and U27660 (N_27660,N_26267,N_26002);
and U27661 (N_27661,N_26535,N_26295);
or U27662 (N_27662,N_26181,N_26088);
nor U27663 (N_27663,N_26723,N_26472);
xor U27664 (N_27664,N_26022,N_26435);
xnor U27665 (N_27665,N_26630,N_26917);
or U27666 (N_27666,N_26071,N_26581);
nor U27667 (N_27667,N_26592,N_26348);
nor U27668 (N_27668,N_26468,N_26380);
xnor U27669 (N_27669,N_26867,N_26857);
nor U27670 (N_27670,N_26728,N_26096);
nand U27671 (N_27671,N_26899,N_26019);
nor U27672 (N_27672,N_26313,N_26414);
and U27673 (N_27673,N_26683,N_26879);
xnor U27674 (N_27674,N_26369,N_26049);
nor U27675 (N_27675,N_26653,N_26879);
nor U27676 (N_27676,N_26959,N_26407);
or U27677 (N_27677,N_26306,N_26761);
or U27678 (N_27678,N_26485,N_26182);
xnor U27679 (N_27679,N_26664,N_26922);
xnor U27680 (N_27680,N_26876,N_26539);
nor U27681 (N_27681,N_26147,N_26203);
xnor U27682 (N_27682,N_26369,N_26425);
and U27683 (N_27683,N_26712,N_26370);
nor U27684 (N_27684,N_26176,N_26516);
and U27685 (N_27685,N_26465,N_26739);
nor U27686 (N_27686,N_26262,N_26813);
nor U27687 (N_27687,N_26968,N_26391);
or U27688 (N_27688,N_26397,N_26654);
or U27689 (N_27689,N_26059,N_26632);
xor U27690 (N_27690,N_26176,N_26037);
nand U27691 (N_27691,N_26105,N_26844);
nor U27692 (N_27692,N_26825,N_26131);
or U27693 (N_27693,N_26326,N_26666);
or U27694 (N_27694,N_26958,N_26333);
nand U27695 (N_27695,N_26539,N_26384);
nor U27696 (N_27696,N_26661,N_26567);
xor U27697 (N_27697,N_26355,N_26480);
nor U27698 (N_27698,N_26247,N_26611);
xnor U27699 (N_27699,N_26142,N_26689);
nor U27700 (N_27700,N_26076,N_26038);
nand U27701 (N_27701,N_26806,N_26538);
xnor U27702 (N_27702,N_26174,N_26015);
or U27703 (N_27703,N_26489,N_26840);
nor U27704 (N_27704,N_26934,N_26234);
nor U27705 (N_27705,N_26174,N_26209);
xor U27706 (N_27706,N_26338,N_26149);
nand U27707 (N_27707,N_26461,N_26394);
xor U27708 (N_27708,N_26193,N_26803);
nand U27709 (N_27709,N_26214,N_26364);
nand U27710 (N_27710,N_26892,N_26472);
nor U27711 (N_27711,N_26482,N_26200);
or U27712 (N_27712,N_26813,N_26567);
xnor U27713 (N_27713,N_26464,N_26192);
nor U27714 (N_27714,N_26753,N_26683);
or U27715 (N_27715,N_26087,N_26297);
and U27716 (N_27716,N_26483,N_26268);
xnor U27717 (N_27717,N_26627,N_26594);
nand U27718 (N_27718,N_26984,N_26816);
xnor U27719 (N_27719,N_26324,N_26775);
or U27720 (N_27720,N_26541,N_26270);
and U27721 (N_27721,N_26052,N_26241);
and U27722 (N_27722,N_26111,N_26148);
or U27723 (N_27723,N_26504,N_26183);
nand U27724 (N_27724,N_26436,N_26746);
xor U27725 (N_27725,N_26197,N_26382);
nor U27726 (N_27726,N_26690,N_26736);
xnor U27727 (N_27727,N_26915,N_26246);
nand U27728 (N_27728,N_26960,N_26217);
or U27729 (N_27729,N_26132,N_26115);
nand U27730 (N_27730,N_26543,N_26353);
nand U27731 (N_27731,N_26051,N_26648);
nand U27732 (N_27732,N_26077,N_26085);
or U27733 (N_27733,N_26959,N_26485);
and U27734 (N_27734,N_26460,N_26122);
nand U27735 (N_27735,N_26112,N_26472);
and U27736 (N_27736,N_26556,N_26149);
xnor U27737 (N_27737,N_26160,N_26233);
nor U27738 (N_27738,N_26857,N_26825);
and U27739 (N_27739,N_26720,N_26034);
nor U27740 (N_27740,N_26762,N_26481);
xnor U27741 (N_27741,N_26844,N_26082);
xnor U27742 (N_27742,N_26085,N_26922);
xor U27743 (N_27743,N_26705,N_26210);
nand U27744 (N_27744,N_26629,N_26433);
xnor U27745 (N_27745,N_26978,N_26867);
xor U27746 (N_27746,N_26502,N_26599);
nand U27747 (N_27747,N_26823,N_26749);
and U27748 (N_27748,N_26094,N_26951);
nor U27749 (N_27749,N_26306,N_26232);
and U27750 (N_27750,N_26440,N_26679);
nor U27751 (N_27751,N_26989,N_26986);
nand U27752 (N_27752,N_26324,N_26839);
and U27753 (N_27753,N_26806,N_26931);
nor U27754 (N_27754,N_26054,N_26870);
nor U27755 (N_27755,N_26120,N_26560);
xnor U27756 (N_27756,N_26242,N_26150);
nand U27757 (N_27757,N_26379,N_26302);
nand U27758 (N_27758,N_26335,N_26298);
xor U27759 (N_27759,N_26055,N_26880);
nand U27760 (N_27760,N_26553,N_26443);
xor U27761 (N_27761,N_26957,N_26467);
nor U27762 (N_27762,N_26885,N_26388);
xnor U27763 (N_27763,N_26104,N_26999);
or U27764 (N_27764,N_26717,N_26295);
and U27765 (N_27765,N_26294,N_26289);
nand U27766 (N_27766,N_26904,N_26293);
xnor U27767 (N_27767,N_26730,N_26318);
or U27768 (N_27768,N_26469,N_26096);
and U27769 (N_27769,N_26659,N_26439);
and U27770 (N_27770,N_26484,N_26147);
nand U27771 (N_27771,N_26126,N_26866);
xnor U27772 (N_27772,N_26511,N_26728);
and U27773 (N_27773,N_26186,N_26368);
nand U27774 (N_27774,N_26976,N_26245);
xor U27775 (N_27775,N_26802,N_26572);
and U27776 (N_27776,N_26841,N_26496);
or U27777 (N_27777,N_26183,N_26071);
nand U27778 (N_27778,N_26191,N_26868);
nand U27779 (N_27779,N_26876,N_26849);
nor U27780 (N_27780,N_26417,N_26908);
nor U27781 (N_27781,N_26443,N_26284);
and U27782 (N_27782,N_26377,N_26130);
or U27783 (N_27783,N_26086,N_26213);
nor U27784 (N_27784,N_26157,N_26696);
xnor U27785 (N_27785,N_26658,N_26690);
and U27786 (N_27786,N_26010,N_26787);
nor U27787 (N_27787,N_26613,N_26567);
nor U27788 (N_27788,N_26948,N_26280);
and U27789 (N_27789,N_26098,N_26277);
nor U27790 (N_27790,N_26927,N_26517);
or U27791 (N_27791,N_26028,N_26432);
nand U27792 (N_27792,N_26353,N_26779);
nand U27793 (N_27793,N_26545,N_26393);
or U27794 (N_27794,N_26286,N_26437);
xnor U27795 (N_27795,N_26226,N_26625);
nand U27796 (N_27796,N_26824,N_26462);
nor U27797 (N_27797,N_26904,N_26017);
nand U27798 (N_27798,N_26187,N_26439);
nor U27799 (N_27799,N_26662,N_26719);
or U27800 (N_27800,N_26429,N_26362);
xnor U27801 (N_27801,N_26053,N_26969);
nand U27802 (N_27802,N_26761,N_26290);
xor U27803 (N_27803,N_26191,N_26913);
nand U27804 (N_27804,N_26978,N_26202);
xor U27805 (N_27805,N_26469,N_26490);
nand U27806 (N_27806,N_26467,N_26743);
xnor U27807 (N_27807,N_26945,N_26238);
nor U27808 (N_27808,N_26024,N_26879);
nor U27809 (N_27809,N_26882,N_26751);
nor U27810 (N_27810,N_26598,N_26233);
or U27811 (N_27811,N_26686,N_26216);
nand U27812 (N_27812,N_26337,N_26120);
xnor U27813 (N_27813,N_26273,N_26903);
or U27814 (N_27814,N_26121,N_26399);
nand U27815 (N_27815,N_26906,N_26365);
and U27816 (N_27816,N_26789,N_26634);
nor U27817 (N_27817,N_26255,N_26495);
and U27818 (N_27818,N_26053,N_26523);
nor U27819 (N_27819,N_26478,N_26406);
and U27820 (N_27820,N_26588,N_26467);
nor U27821 (N_27821,N_26552,N_26480);
xor U27822 (N_27822,N_26900,N_26753);
or U27823 (N_27823,N_26009,N_26127);
and U27824 (N_27824,N_26376,N_26395);
nand U27825 (N_27825,N_26120,N_26428);
xnor U27826 (N_27826,N_26499,N_26722);
nor U27827 (N_27827,N_26294,N_26648);
xnor U27828 (N_27828,N_26735,N_26012);
xor U27829 (N_27829,N_26937,N_26335);
or U27830 (N_27830,N_26381,N_26449);
nor U27831 (N_27831,N_26712,N_26689);
or U27832 (N_27832,N_26264,N_26038);
nor U27833 (N_27833,N_26182,N_26403);
xor U27834 (N_27834,N_26845,N_26209);
and U27835 (N_27835,N_26261,N_26786);
xnor U27836 (N_27836,N_26766,N_26775);
nand U27837 (N_27837,N_26344,N_26608);
nand U27838 (N_27838,N_26881,N_26558);
nor U27839 (N_27839,N_26339,N_26748);
nand U27840 (N_27840,N_26535,N_26987);
and U27841 (N_27841,N_26948,N_26673);
nand U27842 (N_27842,N_26661,N_26357);
xnor U27843 (N_27843,N_26895,N_26848);
nand U27844 (N_27844,N_26963,N_26957);
and U27845 (N_27845,N_26132,N_26522);
xnor U27846 (N_27846,N_26508,N_26441);
and U27847 (N_27847,N_26843,N_26980);
and U27848 (N_27848,N_26785,N_26516);
xnor U27849 (N_27849,N_26641,N_26989);
and U27850 (N_27850,N_26676,N_26472);
and U27851 (N_27851,N_26779,N_26961);
nor U27852 (N_27852,N_26721,N_26850);
xor U27853 (N_27853,N_26339,N_26658);
nor U27854 (N_27854,N_26222,N_26145);
nor U27855 (N_27855,N_26034,N_26384);
or U27856 (N_27856,N_26491,N_26770);
xnor U27857 (N_27857,N_26325,N_26107);
nor U27858 (N_27858,N_26603,N_26595);
or U27859 (N_27859,N_26085,N_26248);
nor U27860 (N_27860,N_26615,N_26061);
xnor U27861 (N_27861,N_26534,N_26334);
nor U27862 (N_27862,N_26439,N_26995);
xor U27863 (N_27863,N_26472,N_26237);
and U27864 (N_27864,N_26134,N_26123);
nor U27865 (N_27865,N_26379,N_26033);
or U27866 (N_27866,N_26053,N_26683);
xnor U27867 (N_27867,N_26249,N_26092);
or U27868 (N_27868,N_26276,N_26114);
or U27869 (N_27869,N_26942,N_26757);
and U27870 (N_27870,N_26376,N_26829);
nand U27871 (N_27871,N_26977,N_26839);
nand U27872 (N_27872,N_26301,N_26077);
and U27873 (N_27873,N_26465,N_26985);
xor U27874 (N_27874,N_26392,N_26150);
xor U27875 (N_27875,N_26417,N_26229);
or U27876 (N_27876,N_26728,N_26304);
nand U27877 (N_27877,N_26191,N_26404);
nor U27878 (N_27878,N_26782,N_26394);
xor U27879 (N_27879,N_26441,N_26974);
or U27880 (N_27880,N_26330,N_26687);
or U27881 (N_27881,N_26668,N_26372);
or U27882 (N_27882,N_26953,N_26008);
nand U27883 (N_27883,N_26864,N_26345);
and U27884 (N_27884,N_26911,N_26016);
xnor U27885 (N_27885,N_26702,N_26756);
nor U27886 (N_27886,N_26428,N_26918);
or U27887 (N_27887,N_26788,N_26324);
or U27888 (N_27888,N_26134,N_26291);
and U27889 (N_27889,N_26940,N_26049);
nor U27890 (N_27890,N_26670,N_26462);
and U27891 (N_27891,N_26685,N_26610);
nand U27892 (N_27892,N_26763,N_26019);
and U27893 (N_27893,N_26912,N_26755);
or U27894 (N_27894,N_26976,N_26918);
and U27895 (N_27895,N_26309,N_26273);
or U27896 (N_27896,N_26760,N_26666);
or U27897 (N_27897,N_26703,N_26477);
xnor U27898 (N_27898,N_26853,N_26774);
nor U27899 (N_27899,N_26234,N_26130);
nor U27900 (N_27900,N_26651,N_26563);
nor U27901 (N_27901,N_26063,N_26703);
and U27902 (N_27902,N_26097,N_26904);
or U27903 (N_27903,N_26726,N_26953);
nor U27904 (N_27904,N_26548,N_26410);
nor U27905 (N_27905,N_26787,N_26947);
nand U27906 (N_27906,N_26219,N_26664);
and U27907 (N_27907,N_26363,N_26050);
xnor U27908 (N_27908,N_26870,N_26505);
or U27909 (N_27909,N_26142,N_26103);
and U27910 (N_27910,N_26114,N_26325);
or U27911 (N_27911,N_26007,N_26945);
nand U27912 (N_27912,N_26894,N_26978);
or U27913 (N_27913,N_26667,N_26392);
xor U27914 (N_27914,N_26291,N_26014);
nor U27915 (N_27915,N_26364,N_26102);
xor U27916 (N_27916,N_26411,N_26736);
or U27917 (N_27917,N_26309,N_26068);
or U27918 (N_27918,N_26411,N_26327);
nand U27919 (N_27919,N_26351,N_26377);
nand U27920 (N_27920,N_26338,N_26573);
xor U27921 (N_27921,N_26807,N_26734);
or U27922 (N_27922,N_26833,N_26711);
nor U27923 (N_27923,N_26127,N_26597);
nor U27924 (N_27924,N_26033,N_26885);
nor U27925 (N_27925,N_26037,N_26013);
and U27926 (N_27926,N_26062,N_26693);
and U27927 (N_27927,N_26688,N_26205);
and U27928 (N_27928,N_26011,N_26364);
nand U27929 (N_27929,N_26927,N_26923);
nand U27930 (N_27930,N_26590,N_26505);
nor U27931 (N_27931,N_26336,N_26066);
xor U27932 (N_27932,N_26885,N_26951);
nand U27933 (N_27933,N_26787,N_26625);
and U27934 (N_27934,N_26040,N_26630);
xor U27935 (N_27935,N_26991,N_26755);
nand U27936 (N_27936,N_26423,N_26756);
xor U27937 (N_27937,N_26568,N_26701);
nand U27938 (N_27938,N_26752,N_26366);
nor U27939 (N_27939,N_26422,N_26435);
or U27940 (N_27940,N_26247,N_26060);
nor U27941 (N_27941,N_26778,N_26512);
and U27942 (N_27942,N_26052,N_26504);
nand U27943 (N_27943,N_26247,N_26267);
nor U27944 (N_27944,N_26934,N_26946);
or U27945 (N_27945,N_26694,N_26829);
and U27946 (N_27946,N_26182,N_26177);
and U27947 (N_27947,N_26768,N_26101);
and U27948 (N_27948,N_26227,N_26119);
nor U27949 (N_27949,N_26004,N_26879);
xnor U27950 (N_27950,N_26018,N_26457);
or U27951 (N_27951,N_26462,N_26616);
or U27952 (N_27952,N_26372,N_26856);
xor U27953 (N_27953,N_26162,N_26164);
or U27954 (N_27954,N_26564,N_26420);
nor U27955 (N_27955,N_26194,N_26037);
and U27956 (N_27956,N_26163,N_26227);
and U27957 (N_27957,N_26489,N_26796);
and U27958 (N_27958,N_26883,N_26928);
xnor U27959 (N_27959,N_26219,N_26495);
nand U27960 (N_27960,N_26850,N_26195);
xor U27961 (N_27961,N_26410,N_26485);
or U27962 (N_27962,N_26300,N_26431);
or U27963 (N_27963,N_26755,N_26500);
xnor U27964 (N_27964,N_26211,N_26992);
nor U27965 (N_27965,N_26459,N_26661);
xnor U27966 (N_27966,N_26017,N_26123);
or U27967 (N_27967,N_26217,N_26645);
xnor U27968 (N_27968,N_26867,N_26969);
xnor U27969 (N_27969,N_26593,N_26717);
nor U27970 (N_27970,N_26805,N_26108);
xnor U27971 (N_27971,N_26079,N_26917);
xnor U27972 (N_27972,N_26458,N_26214);
nor U27973 (N_27973,N_26152,N_26467);
and U27974 (N_27974,N_26226,N_26079);
nor U27975 (N_27975,N_26407,N_26601);
nand U27976 (N_27976,N_26833,N_26319);
xnor U27977 (N_27977,N_26685,N_26047);
xor U27978 (N_27978,N_26394,N_26079);
or U27979 (N_27979,N_26050,N_26284);
xor U27980 (N_27980,N_26059,N_26053);
xor U27981 (N_27981,N_26673,N_26942);
nand U27982 (N_27982,N_26252,N_26827);
or U27983 (N_27983,N_26840,N_26730);
nor U27984 (N_27984,N_26951,N_26423);
and U27985 (N_27985,N_26425,N_26682);
and U27986 (N_27986,N_26266,N_26607);
nand U27987 (N_27987,N_26971,N_26043);
and U27988 (N_27988,N_26626,N_26951);
nor U27989 (N_27989,N_26098,N_26555);
nand U27990 (N_27990,N_26060,N_26347);
xor U27991 (N_27991,N_26645,N_26023);
xnor U27992 (N_27992,N_26624,N_26183);
xnor U27993 (N_27993,N_26014,N_26246);
nand U27994 (N_27994,N_26336,N_26101);
or U27995 (N_27995,N_26646,N_26648);
nand U27996 (N_27996,N_26545,N_26755);
and U27997 (N_27997,N_26191,N_26516);
nand U27998 (N_27998,N_26441,N_26185);
nand U27999 (N_27999,N_26168,N_26812);
xnor U28000 (N_28000,N_27357,N_27933);
or U28001 (N_28001,N_27219,N_27495);
nor U28002 (N_28002,N_27665,N_27330);
xor U28003 (N_28003,N_27459,N_27356);
nor U28004 (N_28004,N_27764,N_27501);
and U28005 (N_28005,N_27490,N_27398);
nor U28006 (N_28006,N_27925,N_27691);
nand U28007 (N_28007,N_27508,N_27715);
nor U28008 (N_28008,N_27127,N_27405);
nand U28009 (N_28009,N_27023,N_27808);
nand U28010 (N_28010,N_27589,N_27008);
nor U28011 (N_28011,N_27460,N_27977);
nor U28012 (N_28012,N_27523,N_27548);
nand U28013 (N_28013,N_27367,N_27617);
or U28014 (N_28014,N_27497,N_27165);
nand U28015 (N_28015,N_27536,N_27346);
and U28016 (N_28016,N_27325,N_27269);
and U28017 (N_28017,N_27760,N_27472);
or U28018 (N_28018,N_27615,N_27794);
and U28019 (N_28019,N_27602,N_27897);
xor U28020 (N_28020,N_27362,N_27716);
nand U28021 (N_28021,N_27452,N_27049);
and U28022 (N_28022,N_27669,N_27254);
xnor U28023 (N_28023,N_27743,N_27124);
nor U28024 (N_28024,N_27146,N_27877);
nor U28025 (N_28025,N_27597,N_27579);
nand U28026 (N_28026,N_27853,N_27500);
nor U28027 (N_28027,N_27327,N_27004);
nor U28028 (N_28028,N_27899,N_27159);
nor U28029 (N_28029,N_27521,N_27735);
xor U28030 (N_28030,N_27571,N_27749);
xor U28031 (N_28031,N_27667,N_27510);
xnor U28032 (N_28032,N_27390,N_27946);
or U28033 (N_28033,N_27134,N_27728);
or U28034 (N_28034,N_27678,N_27085);
and U28035 (N_28035,N_27135,N_27038);
and U28036 (N_28036,N_27368,N_27120);
xor U28037 (N_28037,N_27941,N_27377);
nand U28038 (N_28038,N_27827,N_27240);
nand U28039 (N_28039,N_27378,N_27092);
nor U28040 (N_28040,N_27221,N_27410);
nand U28041 (N_28041,N_27328,N_27932);
nor U28042 (N_28042,N_27507,N_27117);
and U28043 (N_28043,N_27496,N_27971);
nand U28044 (N_28044,N_27005,N_27304);
or U28045 (N_28045,N_27839,N_27097);
or U28046 (N_28046,N_27995,N_27567);
and U28047 (N_28047,N_27639,N_27379);
nor U28048 (N_28048,N_27297,N_27973);
nand U28049 (N_28049,N_27953,N_27638);
nand U28050 (N_28050,N_27040,N_27236);
nor U28051 (N_28051,N_27207,N_27684);
nand U28052 (N_28052,N_27782,N_27891);
nor U28053 (N_28053,N_27758,N_27317);
or U28054 (N_28054,N_27551,N_27320);
xor U28055 (N_28055,N_27746,N_27876);
and U28056 (N_28056,N_27401,N_27302);
and U28057 (N_28057,N_27599,N_27710);
xor U28058 (N_28058,N_27337,N_27614);
nand U28059 (N_28059,N_27871,N_27563);
and U28060 (N_28060,N_27612,N_27613);
xnor U28061 (N_28061,N_27588,N_27966);
nand U28062 (N_28062,N_27059,N_27074);
xnor U28063 (N_28063,N_27306,N_27314);
nor U28064 (N_28064,N_27300,N_27545);
xnor U28065 (N_28065,N_27142,N_27313);
or U28066 (N_28066,N_27064,N_27343);
xor U28067 (N_28067,N_27132,N_27391);
and U28068 (N_28068,N_27642,N_27817);
and U28069 (N_28069,N_27882,N_27262);
xor U28070 (N_28070,N_27018,N_27998);
nor U28071 (N_28071,N_27821,N_27984);
nor U28072 (N_28072,N_27136,N_27596);
nor U28073 (N_28073,N_27488,N_27073);
xor U28074 (N_28074,N_27887,N_27261);
or U28075 (N_28075,N_27895,N_27920);
and U28076 (N_28076,N_27316,N_27771);
xor U28077 (N_28077,N_27232,N_27532);
nor U28078 (N_28078,N_27978,N_27147);
nor U28079 (N_28079,N_27637,N_27937);
xor U28080 (N_28080,N_27110,N_27543);
nor U28081 (N_28081,N_27033,N_27699);
nor U28082 (N_28082,N_27283,N_27475);
nor U28083 (N_28083,N_27241,N_27079);
or U28084 (N_28084,N_27450,N_27983);
and U28085 (N_28085,N_27656,N_27264);
or U28086 (N_28086,N_27089,N_27326);
and U28087 (N_28087,N_27019,N_27039);
or U28088 (N_28088,N_27260,N_27807);
xor U28089 (N_28089,N_27845,N_27526);
xnor U28090 (N_28090,N_27756,N_27359);
nand U28091 (N_28091,N_27867,N_27347);
and U28092 (N_28092,N_27619,N_27572);
or U28093 (N_28093,N_27291,N_27651);
nand U28094 (N_28094,N_27530,N_27943);
nand U28095 (N_28095,N_27773,N_27395);
xor U28096 (N_28096,N_27417,N_27892);
and U28097 (N_28097,N_27139,N_27029);
and U28098 (N_28098,N_27099,N_27842);
xnor U28099 (N_28099,N_27030,N_27901);
and U28100 (N_28100,N_27277,N_27797);
nor U28101 (N_28101,N_27854,N_27374);
nand U28102 (N_28102,N_27516,N_27265);
nor U28103 (N_28103,N_27954,N_27633);
nor U28104 (N_28104,N_27091,N_27032);
nor U28105 (N_28105,N_27829,N_27657);
xnor U28106 (N_28106,N_27394,N_27921);
and U28107 (N_28107,N_27409,N_27974);
nor U28108 (N_28108,N_27245,N_27365);
xnor U28109 (N_28109,N_27286,N_27484);
nor U28110 (N_28110,N_27779,N_27744);
or U28111 (N_28111,N_27708,N_27012);
nor U28112 (N_28112,N_27389,N_27754);
nand U28113 (N_28113,N_27476,N_27422);
nand U28114 (N_28114,N_27875,N_27042);
nand U28115 (N_28115,N_27352,N_27942);
and U28116 (N_28116,N_27202,N_27908);
nor U28117 (N_28117,N_27385,N_27466);
nand U28118 (N_28118,N_27082,N_27905);
nor U28119 (N_28119,N_27664,N_27911);
and U28120 (N_28120,N_27148,N_27483);
nor U28121 (N_28121,N_27800,N_27424);
nor U28122 (N_28122,N_27991,N_27319);
nor U28123 (N_28123,N_27094,N_27885);
xnor U28124 (N_28124,N_27980,N_27230);
or U28125 (N_28125,N_27690,N_27421);
and U28126 (N_28126,N_27119,N_27441);
nand U28127 (N_28127,N_27611,N_27701);
and U28128 (N_28128,N_27267,N_27775);
or U28129 (N_28129,N_27786,N_27680);
xor U28130 (N_28130,N_27272,N_27924);
and U28131 (N_28131,N_27169,N_27175);
xnor U28132 (N_28132,N_27338,N_27949);
nor U28133 (N_28133,N_27962,N_27520);
and U28134 (N_28134,N_27115,N_27540);
nand U28135 (N_28135,N_27366,N_27737);
xnor U28136 (N_28136,N_27558,N_27770);
nor U28137 (N_28137,N_27522,N_27204);
nand U28138 (N_28138,N_27434,N_27098);
nand U28139 (N_28139,N_27080,N_27060);
or U28140 (N_28140,N_27268,N_27806);
nor U28141 (N_28141,N_27907,N_27519);
nor U28142 (N_28142,N_27125,N_27732);
xnor U28143 (N_28143,N_27810,N_27185);
nand U28144 (N_28144,N_27799,N_27178);
or U28145 (N_28145,N_27312,N_27601);
and U28146 (N_28146,N_27252,N_27214);
nand U28147 (N_28147,N_27288,N_27833);
xor U28148 (N_28148,N_27632,N_27965);
or U28149 (N_28149,N_27658,N_27741);
and U28150 (N_28150,N_27284,N_27156);
nand U28151 (N_28151,N_27518,N_27725);
and U28152 (N_28152,N_27149,N_27045);
and U28153 (N_28153,N_27796,N_27071);
xnor U28154 (N_28154,N_27028,N_27618);
nor U28155 (N_28155,N_27511,N_27890);
nand U28156 (N_28156,N_27076,N_27246);
nand U28157 (N_28157,N_27950,N_27660);
and U28158 (N_28158,N_27208,N_27711);
and U28159 (N_28159,N_27333,N_27512);
and U28160 (N_28160,N_27605,N_27626);
and U28161 (N_28161,N_27439,N_27504);
and U28162 (N_28162,N_27593,N_27928);
nor U28163 (N_28163,N_27467,N_27227);
xnor U28164 (N_28164,N_27836,N_27580);
xnor U28165 (N_28165,N_27873,N_27830);
or U28166 (N_28166,N_27964,N_27449);
or U28167 (N_28167,N_27988,N_27888);
xor U28168 (N_28168,N_27783,N_27247);
xnor U28169 (N_28169,N_27989,N_27406);
xnor U28170 (N_28170,N_27948,N_27544);
xor U28171 (N_28171,N_27557,N_27233);
and U28172 (N_28172,N_27868,N_27024);
and U28173 (N_28173,N_27751,N_27457);
and U28174 (N_28174,N_27322,N_27055);
xor U28175 (N_28175,N_27858,N_27163);
nand U28176 (N_28176,N_27184,N_27713);
xor U28177 (N_28177,N_27704,N_27380);
xor U28178 (N_28178,N_27348,N_27620);
or U28179 (N_28179,N_27863,N_27113);
nor U28180 (N_28180,N_27056,N_27213);
nand U28181 (N_28181,N_27963,N_27813);
nand U28182 (N_28182,N_27279,N_27766);
nand U28183 (N_28183,N_27041,N_27193);
nor U28184 (N_28184,N_27654,N_27755);
nand U28185 (N_28185,N_27884,N_27682);
or U28186 (N_28186,N_27253,N_27600);
nand U28187 (N_28187,N_27479,N_27739);
nor U28188 (N_28188,N_27959,N_27538);
and U28189 (N_28189,N_27592,N_27492);
or U28190 (N_28190,N_27513,N_27485);
xnor U28191 (N_28191,N_27017,N_27332);
xnor U28192 (N_28192,N_27688,N_27429);
xnor U28193 (N_28193,N_27609,N_27740);
nor U28194 (N_28194,N_27116,N_27956);
xor U28195 (N_28195,N_27199,N_27590);
and U28196 (N_28196,N_27634,N_27331);
or U28197 (N_28197,N_27862,N_27900);
or U28198 (N_28198,N_27418,N_27805);
nor U28199 (N_28199,N_27586,N_27936);
nor U28200 (N_28200,N_27090,N_27561);
xor U28201 (N_28201,N_27748,N_27225);
nor U28202 (N_28202,N_27624,N_27224);
or U28203 (N_28203,N_27237,N_27341);
xor U28204 (N_28204,N_27172,N_27180);
xnor U28205 (N_28205,N_27370,N_27730);
nor U28206 (N_28206,N_27934,N_27420);
xor U28207 (N_28207,N_27187,N_27635);
nand U28208 (N_28208,N_27058,N_27249);
or U28209 (N_28209,N_27493,N_27077);
nand U28210 (N_28210,N_27273,N_27909);
nand U28211 (N_28211,N_27547,N_27803);
nor U28212 (N_28212,N_27879,N_27448);
and U28213 (N_28213,N_27161,N_27471);
or U28214 (N_28214,N_27869,N_27062);
nand U28215 (N_28215,N_27549,N_27130);
or U28216 (N_28216,N_27747,N_27198);
or U28217 (N_28217,N_27044,N_27242);
xor U28218 (N_28218,N_27404,N_27128);
xnor U28219 (N_28219,N_27792,N_27043);
nor U28220 (N_28220,N_27458,N_27509);
nor U28221 (N_28221,N_27757,N_27673);
nor U28222 (N_28222,N_27902,N_27969);
nand U28223 (N_28223,N_27220,N_27923);
nand U28224 (N_28224,N_27036,N_27164);
and U28225 (N_28225,N_27777,N_27358);
and U28226 (N_28226,N_27203,N_27290);
xor U28227 (N_28227,N_27675,N_27848);
or U28228 (N_28228,N_27481,N_27468);
or U28229 (N_28229,N_27195,N_27918);
xnor U28230 (N_28230,N_27311,N_27408);
xnor U28231 (N_28231,N_27057,N_27436);
or U28232 (N_28232,N_27020,N_27705);
nand U28233 (N_28233,N_27298,N_27835);
and U28234 (N_28234,N_27650,N_27702);
and U28235 (N_28235,N_27299,N_27679);
or U28236 (N_28236,N_27722,N_27065);
or U28237 (N_28237,N_27210,N_27816);
nor U28238 (N_28238,N_27625,N_27307);
and U28239 (N_28239,N_27698,N_27010);
xor U28240 (N_28240,N_27640,N_27898);
xnor U28241 (N_28241,N_27251,N_27647);
nor U28242 (N_28242,N_27832,N_27369);
nor U28243 (N_28243,N_27910,N_27912);
and U28244 (N_28244,N_27896,N_27455);
xnor U28245 (N_28245,N_27721,N_27353);
and U28246 (N_28246,N_27565,N_27981);
and U28247 (N_28247,N_27411,N_27067);
xnor U28248 (N_28248,N_27430,N_27529);
xnor U28249 (N_28249,N_27840,N_27072);
xor U28250 (N_28250,N_27917,N_27822);
or U28251 (N_28251,N_27222,N_27712);
nor U28252 (N_28252,N_27677,N_27778);
xnor U28253 (N_28253,N_27216,N_27000);
nand U28254 (N_28254,N_27636,N_27972);
or U28255 (N_28255,N_27407,N_27886);
and U28256 (N_28256,N_27960,N_27088);
or U28257 (N_28257,N_27445,N_27916);
xnor U28258 (N_28258,N_27021,N_27206);
nor U28259 (N_28259,N_27997,N_27753);
nand U28260 (N_28260,N_27958,N_27537);
and U28261 (N_28261,N_27011,N_27026);
nand U28262 (N_28262,N_27123,N_27692);
xor U28263 (N_28263,N_27013,N_27608);
nor U28264 (N_28264,N_27843,N_27825);
and U28265 (N_28265,N_27776,N_27865);
nor U28266 (N_28266,N_27718,N_27461);
or U28267 (N_28267,N_27939,N_27733);
and U28268 (N_28268,N_27745,N_27812);
nand U28269 (N_28269,N_27938,N_27629);
or U28270 (N_28270,N_27102,N_27447);
xnor U28271 (N_28271,N_27838,N_27014);
xor U28272 (N_28272,N_27282,N_27594);
nor U28273 (N_28273,N_27546,N_27456);
nand U28274 (N_28274,N_27940,N_27433);
nor U28275 (N_28275,N_27604,N_27388);
nor U28276 (N_28276,N_27955,N_27787);
and U28277 (N_28277,N_27087,N_27336);
or U28278 (N_28278,N_27524,N_27138);
xor U28279 (N_28279,N_27315,N_27505);
xnor U28280 (N_28280,N_27437,N_27454);
and U28281 (N_28281,N_27414,N_27935);
and U28282 (N_28282,N_27155,N_27952);
and U28283 (N_28283,N_27703,N_27212);
or U28284 (N_28284,N_27627,N_27861);
nand U28285 (N_28285,N_27681,N_27293);
and U28286 (N_28286,N_27689,N_27630);
xnor U28287 (N_28287,N_27785,N_27235);
or U28288 (N_28288,N_27375,N_27982);
and U28289 (N_28289,N_27815,N_27086);
nand U28290 (N_28290,N_27576,N_27303);
nor U28291 (N_28291,N_27478,N_27761);
or U28292 (N_28292,N_27399,N_27724);
nand U28293 (N_28293,N_27050,N_27736);
nor U28294 (N_28294,N_27685,N_27841);
nand U28295 (N_28295,N_27223,N_27157);
and U28296 (N_28296,N_27616,N_27001);
nor U28297 (N_28297,N_27976,N_27687);
nand U28298 (N_28298,N_27371,N_27443);
nor U28299 (N_28299,N_27824,N_27874);
nor U28300 (N_28300,N_27181,N_27750);
or U28301 (N_28301,N_27256,N_27999);
nand U28302 (N_28302,N_27258,N_27037);
nor U28303 (N_28303,N_27350,N_27427);
nor U28304 (N_28304,N_27052,N_27031);
xnor U28305 (N_28305,N_27788,N_27309);
or U28306 (N_28306,N_27670,N_27162);
nor U28307 (N_28307,N_27061,N_27103);
xnor U28308 (N_28308,N_27859,N_27100);
or U28309 (N_28309,N_27553,N_27402);
or U28310 (N_28310,N_27384,N_27849);
and U28311 (N_28311,N_27083,N_27591);
nor U28312 (N_28312,N_27662,N_27345);
nand U28313 (N_28313,N_27914,N_27700);
and U28314 (N_28314,N_27387,N_27819);
nand U28315 (N_28315,N_27883,N_27944);
or U28316 (N_28316,N_27349,N_27270);
nor U28317 (N_28317,N_27494,N_27506);
and U28318 (N_28318,N_27392,N_27412);
nor U28319 (N_28319,N_27706,N_27428);
nor U28320 (N_28320,N_27166,N_27578);
nand U28321 (N_28321,N_27930,N_27373);
nand U28322 (N_28322,N_27560,N_27595);
nor U28323 (N_28323,N_27351,N_27329);
nor U28324 (N_28324,N_27763,N_27465);
or U28325 (N_28325,N_27781,N_27503);
nor U28326 (N_28326,N_27967,N_27355);
or U28327 (N_28327,N_27133,N_27575);
nor U28328 (N_28328,N_27525,N_27025);
nor U28329 (N_28329,N_27729,N_27364);
xnor U28330 (N_28330,N_27719,N_27393);
nor U28331 (N_28331,N_27108,N_27573);
or U28332 (N_28332,N_27961,N_27112);
nand U28333 (N_28333,N_27182,N_27582);
nor U28334 (N_28334,N_27975,N_27823);
nand U28335 (N_28335,N_27188,N_27354);
xor U28336 (N_28336,N_27340,N_27574);
nor U28337 (N_28337,N_27416,N_27531);
xnor U28338 (N_28338,N_27655,N_27697);
nor U28339 (N_28339,N_27742,N_27913);
nor U28340 (N_28340,N_27360,N_27915);
and U28341 (N_28341,N_27860,N_27141);
nand U28342 (N_28342,N_27793,N_27970);
nand U28343 (N_28343,N_27628,N_27372);
nand U28344 (N_28344,N_27047,N_27238);
or U28345 (N_28345,N_27432,N_27323);
nand U28346 (N_28346,N_27022,N_27790);
nor U28347 (N_28347,N_27415,N_27562);
or U28348 (N_28348,N_27696,N_27568);
and U28349 (N_28349,N_27857,N_27603);
xor U28350 (N_28350,N_27271,N_27979);
or U28351 (N_28351,N_27774,N_27668);
and U28352 (N_28352,N_27831,N_27186);
nand U28353 (N_28353,N_27535,N_27643);
nand U28354 (N_28354,N_27851,N_27446);
nor U28355 (N_28355,N_27791,N_27714);
xnor U28356 (N_28356,N_27435,N_27906);
nor U28357 (N_28357,N_27581,N_27903);
xor U28358 (N_28358,N_27266,N_27487);
xnor U28359 (N_28359,N_27016,N_27275);
or U28360 (N_28360,N_27880,N_27310);
nor U28361 (N_28361,N_27872,N_27334);
and U28362 (N_28362,N_27992,N_27243);
and U28363 (N_28363,N_27814,N_27381);
or U28364 (N_28364,N_27344,N_27095);
nand U28365 (N_28365,N_27878,N_27734);
or U28366 (N_28366,N_27864,N_27287);
or U28367 (N_28367,N_27190,N_27649);
or U28368 (N_28368,N_27197,N_27144);
or U28369 (N_28369,N_27259,N_27027);
and U28370 (N_28370,N_27189,N_27015);
nor U28371 (N_28371,N_27587,N_27321);
and U28372 (N_28372,N_27659,N_27767);
xnor U28373 (N_28373,N_27564,N_27081);
or U28374 (N_28374,N_27818,N_27462);
nand U28375 (N_28375,N_27541,N_27683);
xnor U28376 (N_28376,N_27376,N_27051);
or U28377 (N_28377,N_27795,N_27723);
or U28378 (N_28378,N_27569,N_27693);
nand U28379 (N_28379,N_27996,N_27515);
nand U28380 (N_28380,N_27167,N_27866);
nand U28381 (N_28381,N_27985,N_27550);
and U28382 (N_28382,N_27285,N_27661);
nor U28383 (N_28383,N_27176,N_27470);
or U28384 (N_28384,N_27486,N_27585);
or U28385 (N_28385,N_27844,N_27947);
and U28386 (N_28386,N_27606,N_27295);
xnor U28387 (N_28387,N_27396,N_27179);
nor U28388 (N_28388,N_27281,N_27834);
nor U28389 (N_28389,N_27440,N_27759);
xnor U28390 (N_28390,N_27663,N_27644);
or U28391 (N_28391,N_27382,N_27438);
or U28392 (N_28392,N_27610,N_27068);
or U28393 (N_28393,N_27598,N_27168);
nand U28394 (N_28394,N_27464,N_27765);
xor U28395 (N_28395,N_27276,N_27482);
and U28396 (N_28396,N_27046,N_27200);
or U28397 (N_28397,N_27122,N_27583);
or U28398 (N_28398,N_27318,N_27106);
nand U28399 (N_28399,N_27114,N_27686);
and U28400 (N_28400,N_27768,N_27226);
or U28401 (N_28401,N_27986,N_27847);
nor U28402 (N_28402,N_27666,N_27096);
nor U28403 (N_28403,N_27403,N_27442);
xnor U28404 (N_28404,N_27217,N_27170);
or U28405 (N_28405,N_27623,N_27801);
nand U28406 (N_28406,N_27652,N_27250);
xnor U28407 (N_28407,N_27720,N_27489);
or U28408 (N_28408,N_27889,N_27078);
and U28409 (N_28409,N_27707,N_27231);
and U28410 (N_28410,N_27158,N_27263);
or U28411 (N_28411,N_27552,N_27257);
xor U28412 (N_28412,N_27305,N_27856);
nor U28413 (N_28413,N_27646,N_27607);
nor U28414 (N_28414,N_27363,N_27957);
and U28415 (N_28415,N_27993,N_27361);
nor U28416 (N_28416,N_27278,N_27527);
nand U28417 (N_28417,N_27931,N_27676);
nor U28418 (N_28418,N_27499,N_27534);
xor U28419 (N_28419,N_27093,N_27160);
xor U28420 (N_28420,N_27577,N_27426);
or U28421 (N_28421,N_27566,N_27002);
nor U28422 (N_28422,N_27870,N_27280);
nand U28423 (N_28423,N_27927,N_27131);
xor U28424 (N_28424,N_27811,N_27274);
or U28425 (N_28425,N_27852,N_27945);
xnor U28426 (N_28426,N_27211,N_27752);
nor U28427 (N_28427,N_27453,N_27215);
or U28428 (N_28428,N_27622,N_27709);
nor U28429 (N_28429,N_27694,N_27383);
nor U28430 (N_28430,N_27951,N_27126);
and U28431 (N_28431,N_27335,N_27990);
and U28432 (N_28432,N_27926,N_27121);
nand U28433 (N_28433,N_27035,N_27150);
nand U28434 (N_28434,N_27296,N_27006);
and U28435 (N_28435,N_27053,N_27339);
xnor U28436 (N_28436,N_27554,N_27192);
nor U28437 (N_28437,N_27784,N_27145);
or U28438 (N_28438,N_27772,N_27301);
and U28439 (N_28439,N_27674,N_27539);
xor U28440 (N_28440,N_27431,N_27101);
and U28441 (N_28441,N_27469,N_27894);
nor U28442 (N_28442,N_27229,N_27828);
or U28443 (N_28443,N_27183,N_27555);
nor U28444 (N_28444,N_27292,N_27473);
and U28445 (N_28445,N_27480,N_27502);
and U28446 (N_28446,N_27528,N_27419);
and U28447 (N_28447,N_27413,N_27152);
or U28448 (N_28448,N_27228,N_27463);
xnor U28449 (N_28449,N_27671,N_27118);
or U28450 (N_28450,N_27919,N_27007);
or U28451 (N_28451,N_27798,N_27584);
nor U28452 (N_28452,N_27570,N_27342);
and U28453 (N_28453,N_27922,N_27929);
nor U28454 (N_28454,N_27234,N_27727);
or U28455 (N_28455,N_27542,N_27653);
and U28456 (N_28456,N_27645,N_27672);
nand U28457 (N_28457,N_27474,N_27621);
nand U28458 (N_28458,N_27324,N_27174);
nand U28459 (N_28459,N_27717,N_27194);
nor U28460 (N_28460,N_27173,N_27809);
xnor U28461 (N_28461,N_27738,N_27731);
nand U28462 (N_28462,N_27850,N_27804);
nor U28463 (N_28463,N_27151,N_27987);
and U28464 (N_28464,N_27196,N_27386);
nor U28465 (N_28465,N_27137,N_27968);
xnor U28466 (N_28466,N_27075,N_27255);
xor U28467 (N_28467,N_27239,N_27111);
and U28468 (N_28468,N_27054,N_27153);
nor U28469 (N_28469,N_27425,N_27105);
or U28470 (N_28470,N_27726,N_27009);
nor U28471 (N_28471,N_27129,N_27904);
and U28472 (N_28472,N_27034,N_27994);
nor U28473 (N_28473,N_27191,N_27209);
and U28474 (N_28474,N_27451,N_27881);
and U28475 (N_28475,N_27171,N_27109);
nor U28476 (N_28476,N_27769,N_27143);
nor U28477 (N_28477,N_27248,N_27063);
nand U28478 (N_28478,N_27066,N_27444);
xnor U28479 (N_28479,N_27289,N_27517);
xnor U28480 (N_28480,N_27559,N_27294);
xnor U28481 (N_28481,N_27177,N_27244);
nand U28482 (N_28482,N_27789,N_27048);
nor U28483 (N_28483,N_27069,N_27140);
xnor U28484 (N_28484,N_27397,N_27154);
nor U28485 (N_28485,N_27498,N_27893);
nand U28486 (N_28486,N_27802,N_27205);
xnor U28487 (N_28487,N_27648,N_27400);
nor U28488 (N_28488,N_27695,N_27201);
xor U28489 (N_28489,N_27423,N_27491);
or U28490 (N_28490,N_27820,N_27780);
nand U28491 (N_28491,N_27846,N_27084);
nor U28492 (N_28492,N_27837,N_27641);
or U28493 (N_28493,N_27514,N_27762);
nand U28494 (N_28494,N_27533,N_27556);
nand U28495 (N_28495,N_27003,N_27107);
and U28496 (N_28496,N_27855,N_27826);
xor U28497 (N_28497,N_27104,N_27477);
or U28498 (N_28498,N_27308,N_27070);
and U28499 (N_28499,N_27218,N_27631);
nor U28500 (N_28500,N_27379,N_27306);
nand U28501 (N_28501,N_27203,N_27128);
xor U28502 (N_28502,N_27261,N_27526);
nand U28503 (N_28503,N_27469,N_27513);
or U28504 (N_28504,N_27297,N_27734);
and U28505 (N_28505,N_27993,N_27456);
nor U28506 (N_28506,N_27375,N_27436);
xnor U28507 (N_28507,N_27076,N_27775);
and U28508 (N_28508,N_27699,N_27802);
nand U28509 (N_28509,N_27845,N_27978);
and U28510 (N_28510,N_27217,N_27556);
nor U28511 (N_28511,N_27846,N_27473);
and U28512 (N_28512,N_27424,N_27177);
xor U28513 (N_28513,N_27966,N_27679);
and U28514 (N_28514,N_27014,N_27683);
nand U28515 (N_28515,N_27012,N_27815);
and U28516 (N_28516,N_27672,N_27602);
and U28517 (N_28517,N_27411,N_27499);
and U28518 (N_28518,N_27844,N_27948);
or U28519 (N_28519,N_27049,N_27981);
and U28520 (N_28520,N_27554,N_27544);
nor U28521 (N_28521,N_27484,N_27006);
nor U28522 (N_28522,N_27388,N_27996);
and U28523 (N_28523,N_27211,N_27310);
nand U28524 (N_28524,N_27044,N_27107);
nand U28525 (N_28525,N_27129,N_27404);
nor U28526 (N_28526,N_27057,N_27209);
nor U28527 (N_28527,N_27481,N_27340);
and U28528 (N_28528,N_27953,N_27416);
or U28529 (N_28529,N_27956,N_27150);
nand U28530 (N_28530,N_27379,N_27848);
or U28531 (N_28531,N_27798,N_27220);
and U28532 (N_28532,N_27985,N_27911);
xor U28533 (N_28533,N_27112,N_27122);
and U28534 (N_28534,N_27982,N_27546);
or U28535 (N_28535,N_27695,N_27013);
nand U28536 (N_28536,N_27017,N_27756);
nor U28537 (N_28537,N_27982,N_27435);
and U28538 (N_28538,N_27648,N_27031);
and U28539 (N_28539,N_27228,N_27772);
nor U28540 (N_28540,N_27381,N_27577);
or U28541 (N_28541,N_27415,N_27249);
nand U28542 (N_28542,N_27099,N_27044);
nand U28543 (N_28543,N_27944,N_27223);
and U28544 (N_28544,N_27266,N_27445);
and U28545 (N_28545,N_27713,N_27517);
nand U28546 (N_28546,N_27814,N_27869);
or U28547 (N_28547,N_27826,N_27003);
and U28548 (N_28548,N_27825,N_27186);
nor U28549 (N_28549,N_27791,N_27559);
and U28550 (N_28550,N_27975,N_27219);
and U28551 (N_28551,N_27009,N_27579);
nand U28552 (N_28552,N_27696,N_27570);
or U28553 (N_28553,N_27847,N_27525);
nand U28554 (N_28554,N_27218,N_27248);
or U28555 (N_28555,N_27096,N_27059);
nor U28556 (N_28556,N_27913,N_27240);
xor U28557 (N_28557,N_27972,N_27878);
or U28558 (N_28558,N_27727,N_27179);
nor U28559 (N_28559,N_27155,N_27481);
xor U28560 (N_28560,N_27116,N_27961);
nand U28561 (N_28561,N_27938,N_27162);
or U28562 (N_28562,N_27155,N_27548);
nor U28563 (N_28563,N_27275,N_27348);
nand U28564 (N_28564,N_27033,N_27230);
xnor U28565 (N_28565,N_27825,N_27810);
xor U28566 (N_28566,N_27407,N_27012);
xnor U28567 (N_28567,N_27601,N_27619);
xor U28568 (N_28568,N_27824,N_27025);
nand U28569 (N_28569,N_27953,N_27300);
xor U28570 (N_28570,N_27233,N_27744);
and U28571 (N_28571,N_27001,N_27776);
nor U28572 (N_28572,N_27943,N_27998);
nor U28573 (N_28573,N_27979,N_27387);
nor U28574 (N_28574,N_27459,N_27329);
nand U28575 (N_28575,N_27438,N_27460);
nand U28576 (N_28576,N_27336,N_27797);
xnor U28577 (N_28577,N_27084,N_27609);
xor U28578 (N_28578,N_27302,N_27866);
nor U28579 (N_28579,N_27130,N_27471);
xnor U28580 (N_28580,N_27993,N_27031);
nand U28581 (N_28581,N_27526,N_27164);
nand U28582 (N_28582,N_27539,N_27248);
xor U28583 (N_28583,N_27427,N_27353);
nor U28584 (N_28584,N_27390,N_27736);
and U28585 (N_28585,N_27829,N_27472);
and U28586 (N_28586,N_27689,N_27382);
xor U28587 (N_28587,N_27676,N_27451);
nor U28588 (N_28588,N_27538,N_27560);
and U28589 (N_28589,N_27003,N_27322);
nand U28590 (N_28590,N_27108,N_27442);
and U28591 (N_28591,N_27805,N_27937);
or U28592 (N_28592,N_27640,N_27743);
nand U28593 (N_28593,N_27652,N_27479);
nand U28594 (N_28594,N_27207,N_27572);
nand U28595 (N_28595,N_27025,N_27698);
xnor U28596 (N_28596,N_27081,N_27190);
nor U28597 (N_28597,N_27440,N_27225);
or U28598 (N_28598,N_27272,N_27255);
nand U28599 (N_28599,N_27577,N_27114);
nor U28600 (N_28600,N_27057,N_27721);
and U28601 (N_28601,N_27416,N_27145);
nand U28602 (N_28602,N_27785,N_27439);
xor U28603 (N_28603,N_27269,N_27758);
and U28604 (N_28604,N_27073,N_27459);
or U28605 (N_28605,N_27337,N_27546);
and U28606 (N_28606,N_27226,N_27442);
and U28607 (N_28607,N_27189,N_27659);
nand U28608 (N_28608,N_27041,N_27975);
nand U28609 (N_28609,N_27996,N_27637);
and U28610 (N_28610,N_27093,N_27166);
or U28611 (N_28611,N_27520,N_27265);
nand U28612 (N_28612,N_27337,N_27568);
and U28613 (N_28613,N_27770,N_27375);
or U28614 (N_28614,N_27533,N_27417);
nand U28615 (N_28615,N_27292,N_27253);
or U28616 (N_28616,N_27319,N_27378);
and U28617 (N_28617,N_27664,N_27390);
or U28618 (N_28618,N_27361,N_27489);
nor U28619 (N_28619,N_27415,N_27131);
xnor U28620 (N_28620,N_27163,N_27481);
nor U28621 (N_28621,N_27969,N_27683);
or U28622 (N_28622,N_27366,N_27419);
or U28623 (N_28623,N_27132,N_27013);
or U28624 (N_28624,N_27935,N_27356);
or U28625 (N_28625,N_27170,N_27824);
or U28626 (N_28626,N_27862,N_27102);
or U28627 (N_28627,N_27050,N_27806);
or U28628 (N_28628,N_27120,N_27162);
xnor U28629 (N_28629,N_27930,N_27394);
nor U28630 (N_28630,N_27436,N_27295);
nor U28631 (N_28631,N_27401,N_27856);
nand U28632 (N_28632,N_27384,N_27647);
or U28633 (N_28633,N_27563,N_27179);
nand U28634 (N_28634,N_27987,N_27989);
nor U28635 (N_28635,N_27453,N_27820);
xor U28636 (N_28636,N_27057,N_27941);
nor U28637 (N_28637,N_27754,N_27903);
xor U28638 (N_28638,N_27122,N_27828);
nor U28639 (N_28639,N_27484,N_27934);
and U28640 (N_28640,N_27554,N_27785);
nor U28641 (N_28641,N_27231,N_27365);
nand U28642 (N_28642,N_27155,N_27124);
nand U28643 (N_28643,N_27619,N_27521);
nand U28644 (N_28644,N_27811,N_27319);
xor U28645 (N_28645,N_27796,N_27932);
xnor U28646 (N_28646,N_27048,N_27991);
xor U28647 (N_28647,N_27223,N_27498);
nand U28648 (N_28648,N_27099,N_27752);
nand U28649 (N_28649,N_27698,N_27753);
and U28650 (N_28650,N_27257,N_27950);
nor U28651 (N_28651,N_27810,N_27655);
and U28652 (N_28652,N_27144,N_27896);
xnor U28653 (N_28653,N_27169,N_27654);
nor U28654 (N_28654,N_27445,N_27464);
nor U28655 (N_28655,N_27185,N_27555);
or U28656 (N_28656,N_27262,N_27524);
nor U28657 (N_28657,N_27846,N_27484);
and U28658 (N_28658,N_27936,N_27432);
nand U28659 (N_28659,N_27743,N_27923);
or U28660 (N_28660,N_27269,N_27498);
nor U28661 (N_28661,N_27415,N_27827);
xnor U28662 (N_28662,N_27428,N_27632);
xnor U28663 (N_28663,N_27685,N_27064);
xor U28664 (N_28664,N_27935,N_27474);
or U28665 (N_28665,N_27103,N_27194);
nand U28666 (N_28666,N_27874,N_27307);
nor U28667 (N_28667,N_27178,N_27650);
or U28668 (N_28668,N_27461,N_27086);
or U28669 (N_28669,N_27434,N_27610);
nand U28670 (N_28670,N_27876,N_27963);
nand U28671 (N_28671,N_27952,N_27000);
or U28672 (N_28672,N_27854,N_27119);
nand U28673 (N_28673,N_27315,N_27798);
and U28674 (N_28674,N_27575,N_27935);
nor U28675 (N_28675,N_27320,N_27362);
or U28676 (N_28676,N_27941,N_27592);
nor U28677 (N_28677,N_27825,N_27051);
xor U28678 (N_28678,N_27032,N_27432);
xor U28679 (N_28679,N_27464,N_27812);
xnor U28680 (N_28680,N_27728,N_27300);
nand U28681 (N_28681,N_27125,N_27629);
nand U28682 (N_28682,N_27641,N_27233);
or U28683 (N_28683,N_27095,N_27335);
nand U28684 (N_28684,N_27928,N_27728);
and U28685 (N_28685,N_27880,N_27463);
nand U28686 (N_28686,N_27242,N_27400);
or U28687 (N_28687,N_27692,N_27686);
nor U28688 (N_28688,N_27645,N_27904);
nor U28689 (N_28689,N_27874,N_27180);
nor U28690 (N_28690,N_27138,N_27631);
or U28691 (N_28691,N_27119,N_27431);
and U28692 (N_28692,N_27426,N_27470);
nand U28693 (N_28693,N_27664,N_27073);
xor U28694 (N_28694,N_27977,N_27123);
xor U28695 (N_28695,N_27635,N_27387);
xnor U28696 (N_28696,N_27357,N_27026);
xor U28697 (N_28697,N_27639,N_27448);
nor U28698 (N_28698,N_27401,N_27454);
nand U28699 (N_28699,N_27768,N_27460);
nor U28700 (N_28700,N_27796,N_27066);
nor U28701 (N_28701,N_27045,N_27788);
nand U28702 (N_28702,N_27943,N_27260);
xnor U28703 (N_28703,N_27321,N_27383);
nand U28704 (N_28704,N_27420,N_27427);
and U28705 (N_28705,N_27651,N_27780);
xnor U28706 (N_28706,N_27658,N_27014);
or U28707 (N_28707,N_27541,N_27748);
nor U28708 (N_28708,N_27219,N_27986);
nor U28709 (N_28709,N_27947,N_27854);
or U28710 (N_28710,N_27007,N_27933);
and U28711 (N_28711,N_27860,N_27052);
and U28712 (N_28712,N_27547,N_27512);
nand U28713 (N_28713,N_27722,N_27485);
nor U28714 (N_28714,N_27538,N_27998);
nor U28715 (N_28715,N_27319,N_27372);
nand U28716 (N_28716,N_27313,N_27901);
nor U28717 (N_28717,N_27155,N_27189);
or U28718 (N_28718,N_27155,N_27890);
nand U28719 (N_28719,N_27607,N_27485);
xor U28720 (N_28720,N_27605,N_27151);
xor U28721 (N_28721,N_27642,N_27057);
or U28722 (N_28722,N_27756,N_27295);
nand U28723 (N_28723,N_27243,N_27939);
nor U28724 (N_28724,N_27917,N_27876);
xnor U28725 (N_28725,N_27570,N_27969);
nor U28726 (N_28726,N_27237,N_27782);
or U28727 (N_28727,N_27909,N_27801);
or U28728 (N_28728,N_27643,N_27350);
xnor U28729 (N_28729,N_27675,N_27092);
nand U28730 (N_28730,N_27862,N_27849);
or U28731 (N_28731,N_27681,N_27424);
nor U28732 (N_28732,N_27925,N_27158);
and U28733 (N_28733,N_27047,N_27175);
and U28734 (N_28734,N_27973,N_27733);
or U28735 (N_28735,N_27094,N_27980);
xor U28736 (N_28736,N_27331,N_27186);
and U28737 (N_28737,N_27415,N_27875);
and U28738 (N_28738,N_27876,N_27301);
nor U28739 (N_28739,N_27468,N_27227);
and U28740 (N_28740,N_27211,N_27416);
or U28741 (N_28741,N_27728,N_27109);
and U28742 (N_28742,N_27525,N_27502);
nand U28743 (N_28743,N_27592,N_27607);
xor U28744 (N_28744,N_27317,N_27709);
nor U28745 (N_28745,N_27038,N_27287);
nand U28746 (N_28746,N_27941,N_27189);
and U28747 (N_28747,N_27701,N_27342);
nor U28748 (N_28748,N_27580,N_27465);
nand U28749 (N_28749,N_27431,N_27173);
xor U28750 (N_28750,N_27680,N_27230);
and U28751 (N_28751,N_27772,N_27928);
or U28752 (N_28752,N_27893,N_27071);
or U28753 (N_28753,N_27655,N_27803);
or U28754 (N_28754,N_27112,N_27187);
nand U28755 (N_28755,N_27645,N_27231);
nor U28756 (N_28756,N_27380,N_27493);
and U28757 (N_28757,N_27074,N_27980);
or U28758 (N_28758,N_27285,N_27337);
nand U28759 (N_28759,N_27159,N_27283);
nor U28760 (N_28760,N_27953,N_27527);
or U28761 (N_28761,N_27763,N_27194);
xnor U28762 (N_28762,N_27085,N_27210);
nor U28763 (N_28763,N_27798,N_27639);
xnor U28764 (N_28764,N_27765,N_27924);
xnor U28765 (N_28765,N_27410,N_27996);
nor U28766 (N_28766,N_27545,N_27171);
nand U28767 (N_28767,N_27466,N_27102);
nor U28768 (N_28768,N_27070,N_27606);
nand U28769 (N_28769,N_27836,N_27233);
xor U28770 (N_28770,N_27046,N_27638);
nand U28771 (N_28771,N_27882,N_27730);
xor U28772 (N_28772,N_27839,N_27060);
xnor U28773 (N_28773,N_27564,N_27563);
or U28774 (N_28774,N_27752,N_27083);
or U28775 (N_28775,N_27142,N_27386);
and U28776 (N_28776,N_27111,N_27188);
and U28777 (N_28777,N_27290,N_27047);
nor U28778 (N_28778,N_27113,N_27286);
and U28779 (N_28779,N_27599,N_27204);
nor U28780 (N_28780,N_27774,N_27968);
nor U28781 (N_28781,N_27629,N_27682);
nand U28782 (N_28782,N_27449,N_27171);
nand U28783 (N_28783,N_27092,N_27399);
or U28784 (N_28784,N_27240,N_27246);
nand U28785 (N_28785,N_27039,N_27515);
or U28786 (N_28786,N_27277,N_27704);
nand U28787 (N_28787,N_27698,N_27465);
or U28788 (N_28788,N_27168,N_27864);
or U28789 (N_28789,N_27116,N_27051);
nor U28790 (N_28790,N_27892,N_27745);
nand U28791 (N_28791,N_27283,N_27595);
or U28792 (N_28792,N_27102,N_27506);
or U28793 (N_28793,N_27271,N_27392);
nand U28794 (N_28794,N_27860,N_27011);
and U28795 (N_28795,N_27375,N_27993);
nor U28796 (N_28796,N_27056,N_27440);
or U28797 (N_28797,N_27986,N_27087);
xnor U28798 (N_28798,N_27834,N_27878);
nand U28799 (N_28799,N_27562,N_27053);
nor U28800 (N_28800,N_27792,N_27129);
nor U28801 (N_28801,N_27600,N_27165);
nor U28802 (N_28802,N_27114,N_27235);
and U28803 (N_28803,N_27366,N_27572);
nor U28804 (N_28804,N_27161,N_27212);
nor U28805 (N_28805,N_27410,N_27292);
nor U28806 (N_28806,N_27479,N_27335);
nand U28807 (N_28807,N_27133,N_27750);
or U28808 (N_28808,N_27848,N_27879);
xor U28809 (N_28809,N_27675,N_27871);
xnor U28810 (N_28810,N_27360,N_27407);
and U28811 (N_28811,N_27967,N_27158);
nor U28812 (N_28812,N_27819,N_27887);
and U28813 (N_28813,N_27336,N_27287);
nand U28814 (N_28814,N_27035,N_27831);
nor U28815 (N_28815,N_27394,N_27734);
xor U28816 (N_28816,N_27976,N_27751);
nand U28817 (N_28817,N_27644,N_27634);
nand U28818 (N_28818,N_27589,N_27893);
and U28819 (N_28819,N_27980,N_27313);
nand U28820 (N_28820,N_27605,N_27477);
nand U28821 (N_28821,N_27552,N_27547);
nor U28822 (N_28822,N_27708,N_27194);
nand U28823 (N_28823,N_27454,N_27013);
and U28824 (N_28824,N_27288,N_27113);
nand U28825 (N_28825,N_27327,N_27143);
nand U28826 (N_28826,N_27610,N_27939);
or U28827 (N_28827,N_27692,N_27833);
or U28828 (N_28828,N_27034,N_27035);
and U28829 (N_28829,N_27393,N_27385);
and U28830 (N_28830,N_27244,N_27597);
xnor U28831 (N_28831,N_27011,N_27672);
xnor U28832 (N_28832,N_27880,N_27080);
or U28833 (N_28833,N_27673,N_27393);
and U28834 (N_28834,N_27278,N_27039);
or U28835 (N_28835,N_27952,N_27145);
or U28836 (N_28836,N_27931,N_27726);
nand U28837 (N_28837,N_27195,N_27052);
nand U28838 (N_28838,N_27414,N_27757);
xor U28839 (N_28839,N_27758,N_27669);
or U28840 (N_28840,N_27435,N_27653);
and U28841 (N_28841,N_27980,N_27867);
nor U28842 (N_28842,N_27122,N_27220);
nor U28843 (N_28843,N_27589,N_27320);
and U28844 (N_28844,N_27563,N_27480);
or U28845 (N_28845,N_27517,N_27673);
nand U28846 (N_28846,N_27717,N_27699);
xnor U28847 (N_28847,N_27093,N_27540);
or U28848 (N_28848,N_27173,N_27450);
nor U28849 (N_28849,N_27275,N_27478);
nor U28850 (N_28850,N_27213,N_27579);
nand U28851 (N_28851,N_27822,N_27124);
xor U28852 (N_28852,N_27837,N_27275);
nand U28853 (N_28853,N_27673,N_27257);
nor U28854 (N_28854,N_27687,N_27842);
nand U28855 (N_28855,N_27455,N_27196);
nand U28856 (N_28856,N_27260,N_27322);
xnor U28857 (N_28857,N_27394,N_27526);
xnor U28858 (N_28858,N_27927,N_27210);
nand U28859 (N_28859,N_27590,N_27077);
or U28860 (N_28860,N_27976,N_27288);
nand U28861 (N_28861,N_27868,N_27323);
or U28862 (N_28862,N_27061,N_27401);
and U28863 (N_28863,N_27454,N_27726);
nor U28864 (N_28864,N_27684,N_27644);
xor U28865 (N_28865,N_27275,N_27978);
or U28866 (N_28866,N_27053,N_27887);
nand U28867 (N_28867,N_27784,N_27665);
and U28868 (N_28868,N_27681,N_27590);
xnor U28869 (N_28869,N_27784,N_27948);
nor U28870 (N_28870,N_27596,N_27870);
xnor U28871 (N_28871,N_27623,N_27708);
nor U28872 (N_28872,N_27672,N_27465);
or U28873 (N_28873,N_27812,N_27148);
or U28874 (N_28874,N_27933,N_27112);
and U28875 (N_28875,N_27379,N_27084);
and U28876 (N_28876,N_27747,N_27286);
xor U28877 (N_28877,N_27010,N_27518);
nand U28878 (N_28878,N_27149,N_27300);
and U28879 (N_28879,N_27855,N_27416);
nand U28880 (N_28880,N_27779,N_27348);
nor U28881 (N_28881,N_27008,N_27182);
nor U28882 (N_28882,N_27715,N_27459);
nor U28883 (N_28883,N_27960,N_27819);
xor U28884 (N_28884,N_27162,N_27808);
xnor U28885 (N_28885,N_27947,N_27769);
nor U28886 (N_28886,N_27775,N_27372);
and U28887 (N_28887,N_27396,N_27524);
or U28888 (N_28888,N_27537,N_27123);
and U28889 (N_28889,N_27527,N_27866);
nand U28890 (N_28890,N_27460,N_27852);
nor U28891 (N_28891,N_27078,N_27024);
or U28892 (N_28892,N_27314,N_27284);
nand U28893 (N_28893,N_27853,N_27293);
nand U28894 (N_28894,N_27647,N_27094);
nor U28895 (N_28895,N_27427,N_27813);
xor U28896 (N_28896,N_27832,N_27958);
nand U28897 (N_28897,N_27614,N_27861);
and U28898 (N_28898,N_27419,N_27363);
nand U28899 (N_28899,N_27513,N_27311);
or U28900 (N_28900,N_27634,N_27913);
xor U28901 (N_28901,N_27880,N_27404);
or U28902 (N_28902,N_27466,N_27715);
xnor U28903 (N_28903,N_27935,N_27452);
or U28904 (N_28904,N_27986,N_27524);
and U28905 (N_28905,N_27518,N_27089);
nor U28906 (N_28906,N_27637,N_27968);
and U28907 (N_28907,N_27418,N_27915);
or U28908 (N_28908,N_27369,N_27605);
and U28909 (N_28909,N_27756,N_27018);
nand U28910 (N_28910,N_27744,N_27291);
and U28911 (N_28911,N_27315,N_27342);
nor U28912 (N_28912,N_27871,N_27558);
nor U28913 (N_28913,N_27284,N_27687);
or U28914 (N_28914,N_27995,N_27801);
nand U28915 (N_28915,N_27437,N_27578);
nor U28916 (N_28916,N_27564,N_27609);
xor U28917 (N_28917,N_27949,N_27158);
and U28918 (N_28918,N_27923,N_27928);
nand U28919 (N_28919,N_27084,N_27482);
nor U28920 (N_28920,N_27152,N_27250);
nor U28921 (N_28921,N_27892,N_27507);
nor U28922 (N_28922,N_27221,N_27273);
nor U28923 (N_28923,N_27737,N_27692);
xor U28924 (N_28924,N_27734,N_27891);
or U28925 (N_28925,N_27686,N_27531);
nand U28926 (N_28926,N_27568,N_27559);
nand U28927 (N_28927,N_27746,N_27776);
nand U28928 (N_28928,N_27214,N_27876);
and U28929 (N_28929,N_27988,N_27225);
and U28930 (N_28930,N_27713,N_27276);
xnor U28931 (N_28931,N_27328,N_27272);
xor U28932 (N_28932,N_27145,N_27481);
nand U28933 (N_28933,N_27003,N_27876);
nor U28934 (N_28934,N_27275,N_27934);
nor U28935 (N_28935,N_27081,N_27804);
xnor U28936 (N_28936,N_27439,N_27806);
xor U28937 (N_28937,N_27791,N_27189);
nand U28938 (N_28938,N_27983,N_27430);
nand U28939 (N_28939,N_27061,N_27118);
and U28940 (N_28940,N_27495,N_27419);
xnor U28941 (N_28941,N_27869,N_27825);
nand U28942 (N_28942,N_27814,N_27391);
nor U28943 (N_28943,N_27350,N_27165);
and U28944 (N_28944,N_27881,N_27190);
or U28945 (N_28945,N_27665,N_27560);
and U28946 (N_28946,N_27853,N_27411);
nand U28947 (N_28947,N_27938,N_27878);
xnor U28948 (N_28948,N_27640,N_27985);
or U28949 (N_28949,N_27617,N_27508);
xnor U28950 (N_28950,N_27717,N_27822);
and U28951 (N_28951,N_27658,N_27003);
nor U28952 (N_28952,N_27939,N_27161);
nand U28953 (N_28953,N_27411,N_27611);
xnor U28954 (N_28954,N_27806,N_27193);
nor U28955 (N_28955,N_27459,N_27638);
and U28956 (N_28956,N_27356,N_27623);
or U28957 (N_28957,N_27549,N_27678);
nand U28958 (N_28958,N_27663,N_27682);
and U28959 (N_28959,N_27791,N_27709);
nand U28960 (N_28960,N_27317,N_27634);
and U28961 (N_28961,N_27437,N_27599);
and U28962 (N_28962,N_27888,N_27698);
nand U28963 (N_28963,N_27222,N_27340);
xnor U28964 (N_28964,N_27686,N_27474);
or U28965 (N_28965,N_27906,N_27742);
and U28966 (N_28966,N_27344,N_27670);
or U28967 (N_28967,N_27733,N_27223);
xor U28968 (N_28968,N_27454,N_27552);
nor U28969 (N_28969,N_27912,N_27329);
nor U28970 (N_28970,N_27342,N_27434);
xor U28971 (N_28971,N_27999,N_27068);
nor U28972 (N_28972,N_27753,N_27689);
xnor U28973 (N_28973,N_27857,N_27108);
nor U28974 (N_28974,N_27745,N_27148);
nor U28975 (N_28975,N_27407,N_27721);
nor U28976 (N_28976,N_27831,N_27247);
nor U28977 (N_28977,N_27046,N_27344);
and U28978 (N_28978,N_27289,N_27367);
or U28979 (N_28979,N_27285,N_27274);
nand U28980 (N_28980,N_27698,N_27161);
or U28981 (N_28981,N_27628,N_27283);
or U28982 (N_28982,N_27089,N_27017);
nor U28983 (N_28983,N_27317,N_27874);
nand U28984 (N_28984,N_27048,N_27579);
nand U28985 (N_28985,N_27188,N_27896);
and U28986 (N_28986,N_27021,N_27134);
nor U28987 (N_28987,N_27523,N_27297);
xnor U28988 (N_28988,N_27399,N_27811);
nor U28989 (N_28989,N_27904,N_27054);
nand U28990 (N_28990,N_27243,N_27452);
nor U28991 (N_28991,N_27559,N_27963);
nor U28992 (N_28992,N_27026,N_27101);
xor U28993 (N_28993,N_27658,N_27376);
and U28994 (N_28994,N_27619,N_27183);
xnor U28995 (N_28995,N_27029,N_27571);
xor U28996 (N_28996,N_27673,N_27202);
or U28997 (N_28997,N_27527,N_27174);
nand U28998 (N_28998,N_27927,N_27764);
nor U28999 (N_28999,N_27169,N_27187);
xor U29000 (N_29000,N_28246,N_28680);
nand U29001 (N_29001,N_28217,N_28556);
xnor U29002 (N_29002,N_28096,N_28451);
nand U29003 (N_29003,N_28097,N_28040);
xnor U29004 (N_29004,N_28961,N_28903);
nand U29005 (N_29005,N_28768,N_28271);
or U29006 (N_29006,N_28298,N_28391);
xnor U29007 (N_29007,N_28606,N_28491);
and U29008 (N_29008,N_28579,N_28781);
nor U29009 (N_29009,N_28538,N_28321);
nand U29010 (N_29010,N_28790,N_28181);
or U29011 (N_29011,N_28733,N_28034);
or U29012 (N_29012,N_28964,N_28726);
xor U29013 (N_29013,N_28693,N_28369);
xor U29014 (N_29014,N_28707,N_28174);
xnor U29015 (N_29015,N_28967,N_28895);
and U29016 (N_29016,N_28980,N_28350);
and U29017 (N_29017,N_28496,N_28249);
and U29018 (N_29018,N_28682,N_28081);
nor U29019 (N_29019,N_28786,N_28544);
and U29020 (N_29020,N_28639,N_28337);
nor U29021 (N_29021,N_28603,N_28276);
xor U29022 (N_29022,N_28340,N_28219);
or U29023 (N_29023,N_28974,N_28555);
nand U29024 (N_29024,N_28193,N_28258);
or U29025 (N_29025,N_28857,N_28828);
or U29026 (N_29026,N_28890,N_28493);
or U29027 (N_29027,N_28564,N_28410);
or U29028 (N_29028,N_28216,N_28776);
nand U29029 (N_29029,N_28207,N_28586);
and U29030 (N_29030,N_28613,N_28952);
nand U29031 (N_29031,N_28844,N_28362);
nand U29032 (N_29032,N_28747,N_28566);
or U29033 (N_29033,N_28284,N_28968);
nor U29034 (N_29034,N_28438,N_28226);
xor U29035 (N_29035,N_28529,N_28721);
or U29036 (N_29036,N_28699,N_28705);
nand U29037 (N_29037,N_28200,N_28696);
or U29038 (N_29038,N_28942,N_28933);
xor U29039 (N_29039,N_28342,N_28615);
and U29040 (N_29040,N_28486,N_28110);
xnor U29041 (N_29041,N_28503,N_28013);
nand U29042 (N_29042,N_28701,N_28750);
and U29043 (N_29043,N_28734,N_28637);
or U29044 (N_29044,N_28794,N_28822);
nand U29045 (N_29045,N_28035,N_28230);
xnor U29046 (N_29046,N_28457,N_28435);
nand U29047 (N_29047,N_28584,N_28977);
nand U29048 (N_29048,N_28854,N_28415);
or U29049 (N_29049,N_28558,N_28979);
nor U29050 (N_29050,N_28038,N_28542);
nor U29051 (N_29051,N_28091,N_28837);
nor U29052 (N_29052,N_28899,N_28047);
nor U29053 (N_29053,N_28384,N_28178);
and U29054 (N_29054,N_28946,N_28100);
or U29055 (N_29055,N_28652,N_28166);
nor U29056 (N_29056,N_28028,N_28567);
nor U29057 (N_29057,N_28459,N_28136);
and U29058 (N_29058,N_28473,N_28239);
nand U29059 (N_29059,N_28052,N_28996);
and U29060 (N_29060,N_28803,N_28312);
or U29061 (N_29061,N_28888,N_28860);
and U29062 (N_29062,N_28763,N_28474);
xor U29063 (N_29063,N_28441,N_28562);
nor U29064 (N_29064,N_28196,N_28908);
xor U29065 (N_29065,N_28154,N_28611);
nor U29066 (N_29066,N_28653,N_28422);
nor U29067 (N_29067,N_28029,N_28001);
or U29068 (N_29068,N_28630,N_28525);
and U29069 (N_29069,N_28450,N_28158);
or U29070 (N_29070,N_28983,N_28121);
nor U29071 (N_29071,N_28501,N_28328);
nor U29072 (N_29072,N_28924,N_28736);
or U29073 (N_29073,N_28155,N_28290);
xnor U29074 (N_29074,N_28066,N_28043);
or U29075 (N_29075,N_28805,N_28931);
or U29076 (N_29076,N_28840,N_28278);
or U29077 (N_29077,N_28190,N_28229);
nor U29078 (N_29078,N_28801,N_28521);
nand U29079 (N_29079,N_28004,N_28850);
xnor U29080 (N_29080,N_28070,N_28541);
nand U29081 (N_29081,N_28411,N_28080);
xor U29082 (N_29082,N_28398,N_28170);
nor U29083 (N_29083,N_28728,N_28685);
or U29084 (N_29084,N_28011,N_28918);
nand U29085 (N_29085,N_28616,N_28359);
nor U29086 (N_29086,N_28690,N_28151);
xnor U29087 (N_29087,N_28462,N_28966);
and U29088 (N_29088,N_28746,N_28718);
nand U29089 (N_29089,N_28116,N_28530);
xnor U29090 (N_29090,N_28570,N_28167);
xor U29091 (N_29091,N_28655,N_28823);
and U29092 (N_29092,N_28316,N_28995);
and U29093 (N_29093,N_28565,N_28259);
nand U29094 (N_29094,N_28470,N_28389);
xor U29095 (N_29095,N_28508,N_28999);
or U29096 (N_29096,N_28304,N_28399);
and U29097 (N_29097,N_28793,N_28623);
nor U29098 (N_29098,N_28779,N_28785);
xor U29099 (N_29099,N_28099,N_28471);
or U29100 (N_29100,N_28631,N_28578);
and U29101 (N_29101,N_28550,N_28626);
and U29102 (N_29102,N_28852,N_28078);
and U29103 (N_29103,N_28585,N_28408);
xnor U29104 (N_29104,N_28303,N_28695);
nor U29105 (N_29105,N_28020,N_28195);
nor U29106 (N_29106,N_28686,N_28617);
and U29107 (N_29107,N_28014,N_28346);
or U29108 (N_29108,N_28629,N_28310);
or U29109 (N_29109,N_28376,N_28758);
nor U29110 (N_29110,N_28559,N_28935);
nor U29111 (N_29111,N_28065,N_28939);
and U29112 (N_29112,N_28605,N_28694);
nand U29113 (N_29113,N_28660,N_28609);
or U29114 (N_29114,N_28390,N_28403);
and U29115 (N_29115,N_28622,N_28291);
nand U29116 (N_29116,N_28628,N_28039);
xnor U29117 (N_29117,N_28753,N_28663);
xor U29118 (N_29118,N_28744,N_28460);
xnor U29119 (N_29119,N_28743,N_28560);
nand U29120 (N_29120,N_28168,N_28197);
and U29121 (N_29121,N_28073,N_28830);
xor U29122 (N_29122,N_28642,N_28444);
nand U29123 (N_29123,N_28351,N_28377);
nor U29124 (N_29124,N_28745,N_28475);
or U29125 (N_29125,N_28452,N_28874);
nor U29126 (N_29126,N_28702,N_28127);
nor U29127 (N_29127,N_28727,N_28107);
nor U29128 (N_29128,N_28997,N_28152);
or U29129 (N_29129,N_28101,N_28401);
xor U29130 (N_29130,N_28150,N_28773);
or U29131 (N_29131,N_28597,N_28302);
xnor U29132 (N_29132,N_28943,N_28042);
and U29133 (N_29133,N_28787,N_28932);
nand U29134 (N_29134,N_28719,N_28976);
or U29135 (N_29135,N_28945,N_28331);
xnor U29136 (N_29136,N_28810,N_28296);
or U29137 (N_29137,N_28311,N_28654);
nand U29138 (N_29138,N_28214,N_28905);
nor U29139 (N_29139,N_28133,N_28792);
nand U29140 (N_29140,N_28128,N_28700);
or U29141 (N_29141,N_28956,N_28650);
nor U29142 (N_29142,N_28082,N_28199);
nor U29143 (N_29143,N_28295,N_28349);
or U29144 (N_29144,N_28755,N_28769);
nand U29145 (N_29145,N_28594,N_28009);
nand U29146 (N_29146,N_28656,N_28068);
or U29147 (N_29147,N_28417,N_28426);
or U29148 (N_29148,N_28649,N_28292);
and U29149 (N_29149,N_28533,N_28254);
or U29150 (N_29150,N_28641,N_28927);
nand U29151 (N_29151,N_28665,N_28250);
nor U29152 (N_29152,N_28049,N_28969);
and U29153 (N_29153,N_28075,N_28490);
or U29154 (N_29154,N_28126,N_28892);
and U29155 (N_29155,N_28179,N_28524);
and U29156 (N_29156,N_28545,N_28056);
nor U29157 (N_29157,N_28139,N_28855);
nand U29158 (N_29158,N_28534,N_28002);
nor U29159 (N_29159,N_28306,N_28808);
xnor U29160 (N_29160,N_28574,N_28954);
xor U29161 (N_29161,N_28413,N_28762);
xor U29162 (N_29162,N_28730,N_28251);
and U29163 (N_29163,N_28703,N_28428);
nand U29164 (N_29164,N_28064,N_28016);
and U29165 (N_29165,N_28458,N_28802);
nor U29166 (N_29166,N_28988,N_28737);
and U29167 (N_29167,N_28683,N_28554);
xor U29168 (N_29168,N_28887,N_28963);
xnor U29169 (N_29169,N_28248,N_28050);
nand U29170 (N_29170,N_28947,N_28386);
xor U29171 (N_29171,N_28374,N_28354);
xnor U29172 (N_29172,N_28352,N_28124);
and U29173 (N_29173,N_28183,N_28972);
xor U29174 (N_29174,N_28835,N_28433);
nand U29175 (N_29175,N_28661,N_28848);
and U29176 (N_29176,N_28880,N_28468);
or U29177 (N_29177,N_28711,N_28114);
nor U29178 (N_29178,N_28396,N_28575);
xor U29179 (N_29179,N_28878,N_28227);
xnor U29180 (N_29180,N_28893,N_28506);
or U29181 (N_29181,N_28201,N_28313);
or U29182 (N_29182,N_28838,N_28083);
or U29183 (N_29183,N_28060,N_28361);
and U29184 (N_29184,N_28958,N_28007);
and U29185 (N_29185,N_28112,N_28537);
nand U29186 (N_29186,N_28244,N_28818);
nand U29187 (N_29187,N_28599,N_28089);
xor U29188 (N_29188,N_28169,N_28072);
xnor U29189 (N_29189,N_28164,N_28740);
nor U29190 (N_29190,N_28797,N_28940);
xor U29191 (N_29191,N_28382,N_28233);
nand U29192 (N_29192,N_28627,N_28406);
nand U29193 (N_29193,N_28449,N_28900);
xnor U29194 (N_29194,N_28681,N_28345);
and U29195 (N_29195,N_28867,N_28125);
and U29196 (N_29196,N_28981,N_28273);
and U29197 (N_29197,N_28795,N_28540);
or U29198 (N_29198,N_28677,N_28286);
and U29199 (N_29199,N_28962,N_28548);
or U29200 (N_29200,N_28592,N_28657);
xnor U29201 (N_29201,N_28380,N_28531);
nand U29202 (N_29202,N_28242,N_28647);
xnor U29203 (N_29203,N_28180,N_28388);
nand U29204 (N_29204,N_28536,N_28373);
or U29205 (N_29205,N_28488,N_28061);
and U29206 (N_29206,N_28353,N_28079);
nor U29207 (N_29207,N_28829,N_28057);
or U29208 (N_29208,N_28172,N_28577);
nand U29209 (N_29209,N_28679,N_28381);
nand U29210 (N_29210,N_28055,N_28825);
xor U29211 (N_29211,N_28324,N_28025);
nand U29212 (N_29212,N_28668,N_28601);
or U29213 (N_29213,N_28751,N_28713);
or U29214 (N_29214,N_28416,N_28804);
and U29215 (N_29215,N_28409,N_28670);
and U29216 (N_29216,N_28884,N_28156);
nor U29217 (N_29217,N_28404,N_28317);
and U29218 (N_29218,N_28712,N_28600);
and U29219 (N_29219,N_28624,N_28272);
nand U29220 (N_29220,N_28059,N_28607);
and U29221 (N_29221,N_28191,N_28799);
and U29222 (N_29222,N_28209,N_28383);
nand U29223 (N_29223,N_28175,N_28970);
xnor U29224 (N_29224,N_28319,N_28062);
and U29225 (N_29225,N_28861,N_28847);
xor U29226 (N_29226,N_28722,N_28687);
or U29227 (N_29227,N_28485,N_28777);
and U29228 (N_29228,N_28618,N_28614);
nor U29229 (N_29229,N_28134,N_28315);
nand U29230 (N_29230,N_28561,N_28378);
nand U29231 (N_29231,N_28395,N_28407);
and U29232 (N_29232,N_28784,N_28348);
xor U29233 (N_29233,N_28904,N_28551);
nand U29234 (N_29234,N_28929,N_28138);
nand U29235 (N_29235,N_28765,N_28046);
nor U29236 (N_29236,N_28153,N_28301);
nor U29237 (N_29237,N_28405,N_28975);
xnor U29238 (N_29238,N_28252,N_28775);
nor U29239 (N_29239,N_28005,N_28343);
nand U29240 (N_29240,N_28697,N_28902);
nand U29241 (N_29241,N_28876,N_28309);
nand U29242 (N_29242,N_28044,N_28806);
nor U29243 (N_29243,N_28111,N_28645);
nand U29244 (N_29244,N_28090,N_28421);
or U29245 (N_29245,N_28232,N_28741);
and U29246 (N_29246,N_28820,N_28833);
nor U29247 (N_29247,N_28873,N_28300);
or U29248 (N_29248,N_28184,N_28135);
or U29249 (N_29249,N_28141,N_28287);
xnor U29250 (N_29250,N_28826,N_28698);
nor U29251 (N_29251,N_28516,N_28335);
and U29252 (N_29252,N_28928,N_28739);
xnor U29253 (N_29253,N_28824,N_28221);
or U29254 (N_29254,N_28280,N_28048);
nor U29255 (N_29255,N_28102,N_28595);
nand U29256 (N_29256,N_28394,N_28243);
nand U29257 (N_29257,N_28591,N_28402);
xor U29258 (N_29258,N_28322,N_28400);
nor U29259 (N_29259,N_28710,N_28742);
xnor U29260 (N_29260,N_28211,N_28717);
xnor U29261 (N_29261,N_28092,N_28633);
and U29262 (N_29262,N_28881,N_28288);
or U29263 (N_29263,N_28669,N_28467);
xor U29264 (N_29264,N_28953,N_28103);
xnor U29265 (N_29265,N_28915,N_28610);
and U29266 (N_29266,N_28858,N_28379);
nor U29267 (N_29267,N_28883,N_28187);
xor U29268 (N_29268,N_28263,N_28220);
nor U29269 (N_29269,N_28487,N_28708);
and U29270 (N_29270,N_28326,N_28749);
and U29271 (N_29271,N_28563,N_28285);
or U29272 (N_29272,N_28957,N_28998);
or U29273 (N_29273,N_28236,N_28118);
or U29274 (N_29274,N_28891,N_28788);
nand U29275 (N_29275,N_28791,N_28224);
or U29276 (N_29276,N_28913,N_28872);
nand U29277 (N_29277,N_28638,N_28003);
nor U29278 (N_29278,N_28397,N_28203);
xor U29279 (N_29279,N_28519,N_28885);
nor U29280 (N_29280,N_28356,N_28619);
nand U29281 (N_29281,N_28465,N_28063);
nor U29282 (N_29282,N_28948,N_28691);
nor U29283 (N_29283,N_28176,N_28817);
nand U29284 (N_29284,N_28909,N_28173);
xnor U29285 (N_29285,N_28307,N_28770);
xor U29286 (N_29286,N_28439,N_28257);
nand U29287 (N_29287,N_28420,N_28573);
nor U29288 (N_29288,N_28965,N_28000);
or U29289 (N_29289,N_28704,N_28552);
and U29290 (N_29290,N_28914,N_28440);
nand U29291 (N_29291,N_28274,N_28989);
xor U29292 (N_29292,N_28643,N_28032);
nand U29293 (N_29293,N_28210,N_28582);
nand U29294 (N_29294,N_28821,N_28067);
nor U29295 (N_29295,N_28523,N_28960);
nand U29296 (N_29296,N_28058,N_28546);
nand U29297 (N_29297,N_28780,N_28332);
xnor U29298 (N_29298,N_28188,N_28146);
or U29299 (N_29299,N_28510,N_28093);
nor U29300 (N_29300,N_28204,N_28198);
nor U29301 (N_29301,N_28569,N_28576);
or U29302 (N_29302,N_28715,N_28901);
or U29303 (N_29303,N_28425,N_28938);
nor U29304 (N_29304,N_28430,N_28666);
nand U29305 (N_29305,N_28483,N_28984);
xnor U29306 (N_29306,N_28434,N_28978);
or U29307 (N_29307,N_28723,N_28725);
xor U29308 (N_29308,N_28033,N_28074);
nand U29309 (N_29309,N_28419,N_28667);
nor U29310 (N_29310,N_28509,N_28453);
or U29311 (N_29311,N_28502,N_28228);
nor U29312 (N_29312,N_28796,N_28030);
and U29313 (N_29313,N_28492,N_28235);
or U29314 (N_29314,N_28461,N_28937);
xor U29315 (N_29315,N_28476,N_28906);
nor U29316 (N_29316,N_28256,N_28265);
nand U29317 (N_29317,N_28478,N_28774);
or U29318 (N_29318,N_28323,N_28495);
and U29319 (N_29319,N_28163,N_28270);
xnor U29320 (N_29320,N_28836,N_28879);
xor U29321 (N_29321,N_28731,N_28392);
and U29322 (N_29322,N_28841,N_28941);
xor U29323 (N_29323,N_28076,N_28431);
nor U29324 (N_29324,N_28129,N_28936);
nand U29325 (N_29325,N_28771,N_28675);
nand U29326 (N_29326,N_28706,N_28161);
and U29327 (N_29327,N_28950,N_28087);
nor U29328 (N_29328,N_28442,N_28177);
or U29329 (N_29329,N_28789,N_28489);
nand U29330 (N_29330,N_28593,N_28208);
nand U29331 (N_29331,N_28289,N_28297);
or U29332 (N_29332,N_28539,N_28299);
nor U29333 (N_29333,N_28934,N_28517);
and U29334 (N_29334,N_28782,N_28333);
or U29335 (N_29335,N_28571,N_28859);
nand U29336 (N_29336,N_28532,N_28807);
nor U29337 (N_29337,N_28281,N_28819);
xnor U29338 (N_29338,N_28839,N_28527);
and U29339 (N_29339,N_28264,N_28674);
and U29340 (N_29340,N_28222,N_28990);
nor U29341 (N_29341,N_28477,N_28115);
xor U29342 (N_29342,N_28992,N_28522);
and U29343 (N_29343,N_28088,N_28865);
nand U29344 (N_29344,N_28543,N_28526);
xor U29345 (N_29345,N_28620,N_28305);
nor U29346 (N_29346,N_28756,N_28590);
or U29347 (N_29347,N_28621,N_28646);
and U29348 (N_29348,N_28371,N_28636);
nor U29349 (N_29349,N_28015,N_28507);
and U29350 (N_29350,N_28393,N_28499);
nor U29351 (N_29351,N_28266,N_28366);
or U29352 (N_29352,N_28863,N_28535);
xor U29353 (N_29353,N_28689,N_28240);
or U29354 (N_29354,N_28864,N_28596);
xor U29355 (N_29355,N_28358,N_28283);
nor U29356 (N_29356,N_28238,N_28910);
or U29357 (N_29357,N_28418,N_28385);
and U29358 (N_29358,N_28500,N_28446);
and U29359 (N_29359,N_28484,N_28277);
and U29360 (N_29360,N_28511,N_28759);
nand U29361 (N_29361,N_28955,N_28549);
nor U29362 (N_29362,N_28800,N_28767);
or U29363 (N_29363,N_28123,N_28186);
and U29364 (N_29364,N_28761,N_28024);
xor U29365 (N_29365,N_28144,N_28189);
or U29366 (N_29366,N_28279,N_28951);
nand U29367 (N_29367,N_28424,N_28816);
and U29368 (N_29368,N_28925,N_28206);
nand U29369 (N_29369,N_28031,N_28497);
and U29370 (N_29370,N_28583,N_28520);
nor U29371 (N_29371,N_28512,N_28482);
and U29372 (N_29372,N_28026,N_28877);
nand U29373 (N_29373,N_28991,N_28454);
nor U29374 (N_29374,N_28017,N_28132);
nor U29375 (N_29375,N_28023,N_28772);
nand U29376 (N_29376,N_28131,N_28959);
nor U29377 (N_29377,N_28130,N_28944);
or U29378 (N_29378,N_28095,N_28672);
xor U29379 (N_29379,N_28729,N_28845);
xor U29380 (N_29380,N_28515,N_28357);
or U29381 (N_29381,N_28973,N_28084);
and U29382 (N_29382,N_28308,N_28363);
nand U29383 (N_29383,N_28145,N_28664);
nand U29384 (N_29384,N_28320,N_28027);
or U29385 (N_29385,N_28432,N_28387);
or U29386 (N_29386,N_28119,N_28513);
and U29387 (N_29387,N_28827,N_28994);
nor U29388 (N_29388,N_28160,N_28853);
or U29389 (N_29389,N_28194,N_28368);
nor U29390 (N_29390,N_28692,N_28037);
xor U29391 (N_29391,N_28157,N_28815);
nor U29392 (N_29392,N_28455,N_28949);
nor U29393 (N_29393,N_28241,N_28602);
xnor U29394 (N_29394,N_28720,N_28783);
and U29395 (N_29395,N_28447,N_28262);
nand U29396 (N_29396,N_28896,N_28247);
or U29397 (N_29397,N_28113,N_28868);
nand U29398 (N_29398,N_28588,N_28856);
nand U29399 (N_29399,N_28448,N_28137);
nand U29400 (N_29400,N_28370,N_28923);
nor U29401 (N_29401,N_28735,N_28445);
nor U29402 (N_29402,N_28494,N_28143);
or U29403 (N_29403,N_28843,N_28469);
and U29404 (N_29404,N_28754,N_28897);
nand U29405 (N_29405,N_28504,N_28098);
or U29406 (N_29406,N_28917,N_28269);
nand U29407 (N_29407,N_28580,N_28464);
and U29408 (N_29408,N_28165,N_28648);
or U29409 (N_29409,N_28481,N_28054);
nand U29410 (N_29410,N_28336,N_28245);
and U29411 (N_29411,N_28053,N_28659);
nand U29412 (N_29412,N_28261,N_28866);
nand U29413 (N_29413,N_28218,N_28021);
xor U29414 (N_29414,N_28748,N_28738);
nand U29415 (N_29415,N_28987,N_28640);
or U29416 (N_29416,N_28105,N_28347);
nor U29417 (N_29417,N_28231,N_28926);
nor U29418 (N_29418,N_28022,N_28634);
nor U29419 (N_29419,N_28557,N_28104);
and U29420 (N_29420,N_28724,N_28255);
xnor U29421 (N_29421,N_28849,N_28671);
nor U29422 (N_29422,N_28916,N_28598);
xor U29423 (N_29423,N_28466,N_28752);
nor U29424 (N_29424,N_28365,N_28911);
or U29425 (N_29425,N_28182,N_28282);
and U29426 (N_29426,N_28612,N_28071);
or U29427 (N_29427,N_28684,N_28069);
or U29428 (N_29428,N_28882,N_28012);
and U29429 (N_29429,N_28045,N_28871);
xnor U29430 (N_29430,N_28572,N_28812);
nand U29431 (N_29431,N_28809,N_28443);
nor U29432 (N_29432,N_28919,N_28437);
and U29433 (N_29433,N_28875,N_28212);
xor U29434 (N_29434,N_28094,N_28798);
nand U29435 (N_29435,N_28842,N_28479);
nand U29436 (N_29436,N_28036,N_28514);
nor U29437 (N_29437,N_28709,N_28851);
nor U29438 (N_29438,N_28528,N_28355);
and U29439 (N_29439,N_28676,N_28846);
or U29440 (N_29440,N_28688,N_28215);
or U29441 (N_29441,N_28472,N_28547);
nor U29442 (N_29442,N_28314,N_28427);
xor U29443 (N_29443,N_28498,N_28921);
xnor U29444 (N_29444,N_28898,N_28294);
and U29445 (N_29445,N_28162,N_28912);
nor U29446 (N_29446,N_28225,N_28714);
nor U29447 (N_29447,N_28429,N_28553);
and U29448 (N_29448,N_28051,N_28006);
and U29449 (N_29449,N_28364,N_28732);
nand U29450 (N_29450,N_28625,N_28814);
or U29451 (N_29451,N_28202,N_28367);
nor U29452 (N_29452,N_28922,N_28159);
and U29453 (N_29453,N_28993,N_28318);
nor U29454 (N_29454,N_28673,N_28985);
or U29455 (N_29455,N_28907,N_28632);
nor U29456 (N_29456,N_28658,N_28608);
xor U29457 (N_29457,N_28436,N_28260);
nor U29458 (N_29458,N_28171,N_28117);
xnor U29459 (N_29459,N_28360,N_28223);
nor U29460 (N_29460,N_28518,N_28760);
nand U29461 (N_29461,N_28108,N_28832);
xnor U29462 (N_29462,N_28334,N_28275);
or U29463 (N_29463,N_28267,N_28192);
nor U29464 (N_29464,N_28678,N_28644);
xor U29465 (N_29465,N_28041,N_28010);
nand U29466 (N_29466,N_28920,N_28831);
nor U29467 (N_29467,N_28834,N_28106);
nor U29468 (N_29468,N_28412,N_28930);
or U29469 (N_29469,N_28982,N_28237);
nand U29470 (N_29470,N_28463,N_28587);
and U29471 (N_29471,N_28766,N_28505);
nor U29472 (N_29472,N_28869,N_28019);
nand U29473 (N_29473,N_28568,N_28148);
nor U29474 (N_29474,N_28344,N_28662);
and U29475 (N_29475,N_28339,N_28140);
nand U29476 (N_29476,N_28778,N_28341);
or U29477 (N_29477,N_28716,N_28372);
nor U29478 (N_29478,N_28338,N_28077);
and U29479 (N_29479,N_28651,N_28120);
xor U29480 (N_29480,N_28894,N_28862);
xor U29481 (N_29481,N_28889,N_28764);
or U29482 (N_29482,N_28122,N_28604);
and U29483 (N_29483,N_28147,N_28635);
and U29484 (N_29484,N_28142,N_28329);
xor U29485 (N_29485,N_28293,N_28986);
nand U29486 (N_29486,N_28480,N_28589);
or U29487 (N_29487,N_28456,N_28018);
nand U29488 (N_29488,N_28213,N_28375);
and U29489 (N_29489,N_28813,N_28185);
or U29490 (N_29490,N_28886,N_28234);
nand U29491 (N_29491,N_28086,N_28205);
nor U29492 (N_29492,N_28008,N_28109);
and U29493 (N_29493,N_28325,N_28581);
nand U29494 (N_29494,N_28423,N_28971);
or U29495 (N_29495,N_28414,N_28757);
xnor U29496 (N_29496,N_28253,N_28870);
or U29497 (N_29497,N_28811,N_28085);
or U29498 (N_29498,N_28268,N_28149);
xnor U29499 (N_29499,N_28330,N_28327);
nor U29500 (N_29500,N_28926,N_28714);
xnor U29501 (N_29501,N_28988,N_28326);
nor U29502 (N_29502,N_28582,N_28092);
or U29503 (N_29503,N_28889,N_28501);
xnor U29504 (N_29504,N_28411,N_28329);
nor U29505 (N_29505,N_28741,N_28788);
nand U29506 (N_29506,N_28225,N_28660);
nand U29507 (N_29507,N_28118,N_28052);
and U29508 (N_29508,N_28899,N_28524);
or U29509 (N_29509,N_28311,N_28914);
or U29510 (N_29510,N_28016,N_28354);
xor U29511 (N_29511,N_28382,N_28895);
nor U29512 (N_29512,N_28175,N_28559);
nor U29513 (N_29513,N_28207,N_28089);
xor U29514 (N_29514,N_28867,N_28640);
nand U29515 (N_29515,N_28830,N_28726);
xor U29516 (N_29516,N_28510,N_28244);
nand U29517 (N_29517,N_28812,N_28983);
and U29518 (N_29518,N_28343,N_28945);
or U29519 (N_29519,N_28713,N_28280);
or U29520 (N_29520,N_28008,N_28207);
nand U29521 (N_29521,N_28249,N_28603);
nor U29522 (N_29522,N_28050,N_28657);
and U29523 (N_29523,N_28616,N_28245);
or U29524 (N_29524,N_28986,N_28378);
nand U29525 (N_29525,N_28360,N_28726);
and U29526 (N_29526,N_28228,N_28335);
and U29527 (N_29527,N_28622,N_28552);
and U29528 (N_29528,N_28053,N_28432);
or U29529 (N_29529,N_28557,N_28065);
and U29530 (N_29530,N_28905,N_28522);
or U29531 (N_29531,N_28438,N_28531);
or U29532 (N_29532,N_28757,N_28129);
xnor U29533 (N_29533,N_28711,N_28512);
xnor U29534 (N_29534,N_28266,N_28614);
or U29535 (N_29535,N_28150,N_28607);
nor U29536 (N_29536,N_28324,N_28948);
nor U29537 (N_29537,N_28583,N_28709);
nor U29538 (N_29538,N_28452,N_28997);
nand U29539 (N_29539,N_28421,N_28317);
nor U29540 (N_29540,N_28743,N_28540);
nand U29541 (N_29541,N_28058,N_28463);
or U29542 (N_29542,N_28502,N_28942);
or U29543 (N_29543,N_28239,N_28996);
or U29544 (N_29544,N_28214,N_28064);
xnor U29545 (N_29545,N_28883,N_28102);
xnor U29546 (N_29546,N_28110,N_28263);
or U29547 (N_29547,N_28543,N_28709);
nand U29548 (N_29548,N_28403,N_28646);
or U29549 (N_29549,N_28964,N_28817);
xor U29550 (N_29550,N_28915,N_28237);
and U29551 (N_29551,N_28904,N_28760);
nand U29552 (N_29552,N_28010,N_28937);
xnor U29553 (N_29553,N_28958,N_28532);
or U29554 (N_29554,N_28561,N_28689);
xnor U29555 (N_29555,N_28589,N_28043);
nand U29556 (N_29556,N_28282,N_28899);
nor U29557 (N_29557,N_28913,N_28498);
nand U29558 (N_29558,N_28708,N_28130);
and U29559 (N_29559,N_28510,N_28898);
and U29560 (N_29560,N_28579,N_28882);
nand U29561 (N_29561,N_28692,N_28522);
xnor U29562 (N_29562,N_28065,N_28052);
or U29563 (N_29563,N_28930,N_28946);
or U29564 (N_29564,N_28609,N_28256);
and U29565 (N_29565,N_28015,N_28525);
nand U29566 (N_29566,N_28585,N_28844);
xor U29567 (N_29567,N_28893,N_28654);
nor U29568 (N_29568,N_28723,N_28996);
xnor U29569 (N_29569,N_28873,N_28472);
nor U29570 (N_29570,N_28282,N_28895);
and U29571 (N_29571,N_28547,N_28436);
and U29572 (N_29572,N_28485,N_28186);
xnor U29573 (N_29573,N_28853,N_28399);
nand U29574 (N_29574,N_28060,N_28005);
xnor U29575 (N_29575,N_28558,N_28883);
xor U29576 (N_29576,N_28920,N_28134);
nor U29577 (N_29577,N_28859,N_28580);
xnor U29578 (N_29578,N_28388,N_28951);
xor U29579 (N_29579,N_28908,N_28337);
and U29580 (N_29580,N_28766,N_28148);
nand U29581 (N_29581,N_28298,N_28853);
xnor U29582 (N_29582,N_28695,N_28076);
nor U29583 (N_29583,N_28411,N_28870);
or U29584 (N_29584,N_28525,N_28442);
xor U29585 (N_29585,N_28492,N_28327);
nand U29586 (N_29586,N_28596,N_28656);
nor U29587 (N_29587,N_28345,N_28218);
nand U29588 (N_29588,N_28521,N_28675);
and U29589 (N_29589,N_28759,N_28226);
or U29590 (N_29590,N_28807,N_28567);
or U29591 (N_29591,N_28610,N_28586);
nand U29592 (N_29592,N_28962,N_28970);
or U29593 (N_29593,N_28539,N_28781);
xor U29594 (N_29594,N_28242,N_28069);
nand U29595 (N_29595,N_28326,N_28416);
or U29596 (N_29596,N_28520,N_28958);
and U29597 (N_29597,N_28992,N_28057);
xnor U29598 (N_29598,N_28106,N_28509);
nand U29599 (N_29599,N_28697,N_28156);
and U29600 (N_29600,N_28296,N_28531);
nand U29601 (N_29601,N_28656,N_28065);
nor U29602 (N_29602,N_28429,N_28086);
or U29603 (N_29603,N_28073,N_28510);
xor U29604 (N_29604,N_28373,N_28680);
nor U29605 (N_29605,N_28913,N_28203);
and U29606 (N_29606,N_28194,N_28462);
nand U29607 (N_29607,N_28866,N_28541);
or U29608 (N_29608,N_28877,N_28668);
nor U29609 (N_29609,N_28159,N_28528);
and U29610 (N_29610,N_28439,N_28997);
or U29611 (N_29611,N_28705,N_28118);
nand U29612 (N_29612,N_28810,N_28906);
and U29613 (N_29613,N_28428,N_28440);
xor U29614 (N_29614,N_28522,N_28824);
or U29615 (N_29615,N_28348,N_28891);
nor U29616 (N_29616,N_28675,N_28754);
nor U29617 (N_29617,N_28479,N_28772);
nand U29618 (N_29618,N_28028,N_28122);
xnor U29619 (N_29619,N_28973,N_28278);
or U29620 (N_29620,N_28393,N_28336);
or U29621 (N_29621,N_28315,N_28359);
nor U29622 (N_29622,N_28442,N_28220);
xor U29623 (N_29623,N_28388,N_28249);
nor U29624 (N_29624,N_28099,N_28451);
xnor U29625 (N_29625,N_28097,N_28541);
nor U29626 (N_29626,N_28183,N_28165);
xnor U29627 (N_29627,N_28364,N_28217);
nand U29628 (N_29628,N_28724,N_28216);
nand U29629 (N_29629,N_28655,N_28700);
xnor U29630 (N_29630,N_28526,N_28130);
nand U29631 (N_29631,N_28756,N_28362);
nor U29632 (N_29632,N_28492,N_28084);
or U29633 (N_29633,N_28743,N_28539);
xor U29634 (N_29634,N_28107,N_28495);
and U29635 (N_29635,N_28699,N_28317);
xnor U29636 (N_29636,N_28673,N_28709);
and U29637 (N_29637,N_28274,N_28795);
xnor U29638 (N_29638,N_28912,N_28588);
or U29639 (N_29639,N_28535,N_28649);
xor U29640 (N_29640,N_28370,N_28520);
or U29641 (N_29641,N_28113,N_28809);
or U29642 (N_29642,N_28144,N_28722);
nor U29643 (N_29643,N_28231,N_28042);
and U29644 (N_29644,N_28419,N_28757);
nor U29645 (N_29645,N_28900,N_28680);
nand U29646 (N_29646,N_28553,N_28401);
or U29647 (N_29647,N_28433,N_28607);
or U29648 (N_29648,N_28595,N_28040);
or U29649 (N_29649,N_28902,N_28359);
nand U29650 (N_29650,N_28054,N_28335);
nand U29651 (N_29651,N_28517,N_28658);
and U29652 (N_29652,N_28456,N_28356);
nor U29653 (N_29653,N_28316,N_28300);
or U29654 (N_29654,N_28310,N_28684);
xor U29655 (N_29655,N_28608,N_28838);
and U29656 (N_29656,N_28814,N_28985);
nand U29657 (N_29657,N_28798,N_28044);
or U29658 (N_29658,N_28108,N_28147);
or U29659 (N_29659,N_28838,N_28109);
nor U29660 (N_29660,N_28203,N_28299);
nand U29661 (N_29661,N_28525,N_28666);
or U29662 (N_29662,N_28989,N_28552);
xnor U29663 (N_29663,N_28864,N_28687);
xnor U29664 (N_29664,N_28611,N_28087);
xor U29665 (N_29665,N_28779,N_28433);
or U29666 (N_29666,N_28213,N_28688);
or U29667 (N_29667,N_28971,N_28656);
and U29668 (N_29668,N_28090,N_28629);
or U29669 (N_29669,N_28327,N_28507);
or U29670 (N_29670,N_28891,N_28376);
xnor U29671 (N_29671,N_28628,N_28993);
xnor U29672 (N_29672,N_28253,N_28984);
or U29673 (N_29673,N_28527,N_28854);
and U29674 (N_29674,N_28584,N_28140);
nor U29675 (N_29675,N_28408,N_28638);
or U29676 (N_29676,N_28140,N_28758);
xor U29677 (N_29677,N_28122,N_28660);
or U29678 (N_29678,N_28421,N_28469);
nor U29679 (N_29679,N_28491,N_28673);
xnor U29680 (N_29680,N_28189,N_28545);
or U29681 (N_29681,N_28032,N_28743);
nor U29682 (N_29682,N_28164,N_28383);
or U29683 (N_29683,N_28847,N_28282);
or U29684 (N_29684,N_28098,N_28449);
xnor U29685 (N_29685,N_28415,N_28687);
nor U29686 (N_29686,N_28647,N_28411);
nor U29687 (N_29687,N_28098,N_28873);
nor U29688 (N_29688,N_28963,N_28709);
nand U29689 (N_29689,N_28537,N_28987);
and U29690 (N_29690,N_28156,N_28422);
or U29691 (N_29691,N_28976,N_28702);
nand U29692 (N_29692,N_28921,N_28068);
nand U29693 (N_29693,N_28699,N_28422);
xor U29694 (N_29694,N_28801,N_28800);
and U29695 (N_29695,N_28094,N_28989);
nor U29696 (N_29696,N_28223,N_28261);
nor U29697 (N_29697,N_28514,N_28430);
nor U29698 (N_29698,N_28721,N_28413);
nand U29699 (N_29699,N_28086,N_28191);
nand U29700 (N_29700,N_28780,N_28739);
or U29701 (N_29701,N_28313,N_28572);
nand U29702 (N_29702,N_28172,N_28439);
or U29703 (N_29703,N_28860,N_28303);
or U29704 (N_29704,N_28085,N_28298);
and U29705 (N_29705,N_28939,N_28692);
and U29706 (N_29706,N_28472,N_28860);
or U29707 (N_29707,N_28489,N_28059);
xor U29708 (N_29708,N_28561,N_28709);
nand U29709 (N_29709,N_28885,N_28419);
and U29710 (N_29710,N_28742,N_28739);
or U29711 (N_29711,N_28293,N_28772);
and U29712 (N_29712,N_28761,N_28931);
xnor U29713 (N_29713,N_28667,N_28144);
or U29714 (N_29714,N_28257,N_28015);
xnor U29715 (N_29715,N_28447,N_28156);
and U29716 (N_29716,N_28696,N_28396);
nor U29717 (N_29717,N_28000,N_28728);
xnor U29718 (N_29718,N_28005,N_28954);
nand U29719 (N_29719,N_28594,N_28130);
and U29720 (N_29720,N_28042,N_28606);
nor U29721 (N_29721,N_28664,N_28209);
or U29722 (N_29722,N_28826,N_28270);
and U29723 (N_29723,N_28835,N_28872);
or U29724 (N_29724,N_28345,N_28119);
and U29725 (N_29725,N_28969,N_28229);
xor U29726 (N_29726,N_28918,N_28185);
and U29727 (N_29727,N_28322,N_28560);
nand U29728 (N_29728,N_28090,N_28988);
nor U29729 (N_29729,N_28247,N_28130);
xor U29730 (N_29730,N_28740,N_28242);
xor U29731 (N_29731,N_28503,N_28115);
and U29732 (N_29732,N_28007,N_28806);
and U29733 (N_29733,N_28351,N_28614);
and U29734 (N_29734,N_28280,N_28474);
and U29735 (N_29735,N_28063,N_28499);
nor U29736 (N_29736,N_28417,N_28396);
xnor U29737 (N_29737,N_28950,N_28915);
or U29738 (N_29738,N_28713,N_28100);
or U29739 (N_29739,N_28644,N_28608);
nand U29740 (N_29740,N_28779,N_28491);
nand U29741 (N_29741,N_28231,N_28248);
nor U29742 (N_29742,N_28195,N_28946);
or U29743 (N_29743,N_28485,N_28133);
xnor U29744 (N_29744,N_28453,N_28214);
and U29745 (N_29745,N_28152,N_28851);
xor U29746 (N_29746,N_28986,N_28405);
and U29747 (N_29747,N_28416,N_28767);
nor U29748 (N_29748,N_28427,N_28872);
xor U29749 (N_29749,N_28946,N_28274);
xor U29750 (N_29750,N_28626,N_28622);
xnor U29751 (N_29751,N_28909,N_28245);
and U29752 (N_29752,N_28259,N_28622);
xor U29753 (N_29753,N_28070,N_28488);
nand U29754 (N_29754,N_28415,N_28890);
nor U29755 (N_29755,N_28507,N_28304);
or U29756 (N_29756,N_28760,N_28307);
or U29757 (N_29757,N_28678,N_28534);
or U29758 (N_29758,N_28456,N_28726);
nand U29759 (N_29759,N_28005,N_28971);
xor U29760 (N_29760,N_28377,N_28208);
or U29761 (N_29761,N_28006,N_28654);
or U29762 (N_29762,N_28851,N_28577);
or U29763 (N_29763,N_28936,N_28848);
nor U29764 (N_29764,N_28668,N_28177);
and U29765 (N_29765,N_28954,N_28100);
nand U29766 (N_29766,N_28536,N_28140);
xor U29767 (N_29767,N_28635,N_28222);
xor U29768 (N_29768,N_28265,N_28368);
and U29769 (N_29769,N_28513,N_28948);
nand U29770 (N_29770,N_28068,N_28073);
nand U29771 (N_29771,N_28703,N_28101);
or U29772 (N_29772,N_28850,N_28672);
and U29773 (N_29773,N_28316,N_28241);
and U29774 (N_29774,N_28425,N_28784);
and U29775 (N_29775,N_28125,N_28869);
or U29776 (N_29776,N_28147,N_28068);
xnor U29777 (N_29777,N_28590,N_28406);
xor U29778 (N_29778,N_28440,N_28457);
xnor U29779 (N_29779,N_28675,N_28213);
xor U29780 (N_29780,N_28068,N_28162);
xor U29781 (N_29781,N_28823,N_28765);
xnor U29782 (N_29782,N_28215,N_28661);
nor U29783 (N_29783,N_28486,N_28270);
and U29784 (N_29784,N_28468,N_28454);
or U29785 (N_29785,N_28382,N_28528);
nor U29786 (N_29786,N_28570,N_28430);
xor U29787 (N_29787,N_28260,N_28669);
nand U29788 (N_29788,N_28833,N_28642);
nand U29789 (N_29789,N_28671,N_28357);
nand U29790 (N_29790,N_28231,N_28992);
nor U29791 (N_29791,N_28882,N_28896);
nor U29792 (N_29792,N_28072,N_28623);
nor U29793 (N_29793,N_28447,N_28142);
or U29794 (N_29794,N_28531,N_28818);
or U29795 (N_29795,N_28835,N_28815);
xor U29796 (N_29796,N_28859,N_28834);
and U29797 (N_29797,N_28960,N_28332);
or U29798 (N_29798,N_28534,N_28786);
and U29799 (N_29799,N_28012,N_28916);
xnor U29800 (N_29800,N_28605,N_28995);
nor U29801 (N_29801,N_28730,N_28708);
or U29802 (N_29802,N_28113,N_28499);
nand U29803 (N_29803,N_28874,N_28416);
nand U29804 (N_29804,N_28292,N_28862);
nand U29805 (N_29805,N_28178,N_28834);
nor U29806 (N_29806,N_28868,N_28082);
and U29807 (N_29807,N_28298,N_28195);
xor U29808 (N_29808,N_28541,N_28902);
or U29809 (N_29809,N_28495,N_28688);
nand U29810 (N_29810,N_28396,N_28391);
and U29811 (N_29811,N_28942,N_28864);
or U29812 (N_29812,N_28895,N_28208);
or U29813 (N_29813,N_28855,N_28026);
nand U29814 (N_29814,N_28641,N_28134);
and U29815 (N_29815,N_28013,N_28695);
and U29816 (N_29816,N_28756,N_28625);
nor U29817 (N_29817,N_28083,N_28044);
nor U29818 (N_29818,N_28280,N_28886);
nor U29819 (N_29819,N_28030,N_28539);
and U29820 (N_29820,N_28445,N_28461);
and U29821 (N_29821,N_28672,N_28373);
nor U29822 (N_29822,N_28418,N_28886);
xnor U29823 (N_29823,N_28635,N_28965);
nor U29824 (N_29824,N_28706,N_28097);
nor U29825 (N_29825,N_28019,N_28717);
nand U29826 (N_29826,N_28443,N_28551);
and U29827 (N_29827,N_28392,N_28126);
xor U29828 (N_29828,N_28774,N_28218);
nand U29829 (N_29829,N_28455,N_28733);
and U29830 (N_29830,N_28429,N_28624);
xnor U29831 (N_29831,N_28804,N_28285);
nor U29832 (N_29832,N_28166,N_28918);
nand U29833 (N_29833,N_28520,N_28366);
xnor U29834 (N_29834,N_28922,N_28705);
nor U29835 (N_29835,N_28282,N_28805);
nor U29836 (N_29836,N_28371,N_28848);
xor U29837 (N_29837,N_28647,N_28366);
nor U29838 (N_29838,N_28898,N_28446);
nand U29839 (N_29839,N_28598,N_28124);
and U29840 (N_29840,N_28604,N_28096);
nand U29841 (N_29841,N_28332,N_28171);
xor U29842 (N_29842,N_28576,N_28990);
and U29843 (N_29843,N_28581,N_28497);
or U29844 (N_29844,N_28213,N_28117);
nor U29845 (N_29845,N_28476,N_28388);
nor U29846 (N_29846,N_28505,N_28037);
and U29847 (N_29847,N_28404,N_28374);
nor U29848 (N_29848,N_28901,N_28313);
nor U29849 (N_29849,N_28316,N_28057);
xor U29850 (N_29850,N_28080,N_28524);
nor U29851 (N_29851,N_28881,N_28236);
or U29852 (N_29852,N_28852,N_28103);
nor U29853 (N_29853,N_28391,N_28056);
nand U29854 (N_29854,N_28104,N_28291);
and U29855 (N_29855,N_28497,N_28015);
nand U29856 (N_29856,N_28104,N_28012);
nand U29857 (N_29857,N_28028,N_28079);
xnor U29858 (N_29858,N_28914,N_28714);
and U29859 (N_29859,N_28743,N_28053);
and U29860 (N_29860,N_28703,N_28035);
xor U29861 (N_29861,N_28509,N_28443);
xnor U29862 (N_29862,N_28921,N_28412);
nand U29863 (N_29863,N_28998,N_28712);
nor U29864 (N_29864,N_28324,N_28173);
xor U29865 (N_29865,N_28882,N_28954);
or U29866 (N_29866,N_28673,N_28213);
xor U29867 (N_29867,N_28897,N_28451);
or U29868 (N_29868,N_28306,N_28234);
xnor U29869 (N_29869,N_28248,N_28115);
xnor U29870 (N_29870,N_28379,N_28689);
and U29871 (N_29871,N_28885,N_28438);
xor U29872 (N_29872,N_28302,N_28288);
and U29873 (N_29873,N_28626,N_28311);
nand U29874 (N_29874,N_28793,N_28857);
and U29875 (N_29875,N_28463,N_28688);
nand U29876 (N_29876,N_28216,N_28413);
xnor U29877 (N_29877,N_28381,N_28468);
or U29878 (N_29878,N_28634,N_28470);
or U29879 (N_29879,N_28257,N_28422);
nand U29880 (N_29880,N_28948,N_28416);
nand U29881 (N_29881,N_28108,N_28275);
xor U29882 (N_29882,N_28253,N_28786);
nand U29883 (N_29883,N_28960,N_28138);
and U29884 (N_29884,N_28348,N_28904);
or U29885 (N_29885,N_28936,N_28667);
nand U29886 (N_29886,N_28306,N_28561);
xor U29887 (N_29887,N_28765,N_28432);
nand U29888 (N_29888,N_28541,N_28229);
or U29889 (N_29889,N_28587,N_28414);
nor U29890 (N_29890,N_28332,N_28916);
xnor U29891 (N_29891,N_28168,N_28745);
nor U29892 (N_29892,N_28365,N_28953);
nor U29893 (N_29893,N_28353,N_28022);
xor U29894 (N_29894,N_28137,N_28502);
nor U29895 (N_29895,N_28171,N_28932);
xor U29896 (N_29896,N_28054,N_28020);
nor U29897 (N_29897,N_28992,N_28128);
nand U29898 (N_29898,N_28411,N_28997);
or U29899 (N_29899,N_28006,N_28047);
nor U29900 (N_29900,N_28219,N_28132);
nor U29901 (N_29901,N_28469,N_28826);
nor U29902 (N_29902,N_28821,N_28887);
or U29903 (N_29903,N_28489,N_28047);
and U29904 (N_29904,N_28613,N_28023);
xor U29905 (N_29905,N_28036,N_28563);
or U29906 (N_29906,N_28124,N_28022);
nand U29907 (N_29907,N_28360,N_28155);
nand U29908 (N_29908,N_28329,N_28697);
xor U29909 (N_29909,N_28947,N_28124);
xnor U29910 (N_29910,N_28395,N_28491);
and U29911 (N_29911,N_28462,N_28366);
or U29912 (N_29912,N_28479,N_28960);
xor U29913 (N_29913,N_28168,N_28279);
nor U29914 (N_29914,N_28337,N_28769);
nor U29915 (N_29915,N_28728,N_28018);
xor U29916 (N_29916,N_28874,N_28661);
xor U29917 (N_29917,N_28916,N_28565);
and U29918 (N_29918,N_28235,N_28048);
nand U29919 (N_29919,N_28685,N_28329);
or U29920 (N_29920,N_28110,N_28196);
and U29921 (N_29921,N_28283,N_28905);
and U29922 (N_29922,N_28198,N_28999);
and U29923 (N_29923,N_28223,N_28156);
xnor U29924 (N_29924,N_28939,N_28843);
nor U29925 (N_29925,N_28536,N_28416);
xor U29926 (N_29926,N_28903,N_28204);
nand U29927 (N_29927,N_28516,N_28284);
nand U29928 (N_29928,N_28800,N_28017);
xnor U29929 (N_29929,N_28100,N_28995);
nand U29930 (N_29930,N_28293,N_28183);
nor U29931 (N_29931,N_28410,N_28590);
nor U29932 (N_29932,N_28136,N_28627);
nor U29933 (N_29933,N_28487,N_28990);
or U29934 (N_29934,N_28412,N_28812);
nand U29935 (N_29935,N_28248,N_28326);
and U29936 (N_29936,N_28701,N_28854);
xnor U29937 (N_29937,N_28080,N_28780);
and U29938 (N_29938,N_28096,N_28391);
xnor U29939 (N_29939,N_28332,N_28092);
xor U29940 (N_29940,N_28296,N_28820);
or U29941 (N_29941,N_28791,N_28496);
or U29942 (N_29942,N_28047,N_28800);
nor U29943 (N_29943,N_28914,N_28629);
and U29944 (N_29944,N_28285,N_28196);
xor U29945 (N_29945,N_28179,N_28974);
and U29946 (N_29946,N_28293,N_28787);
nand U29947 (N_29947,N_28297,N_28582);
nor U29948 (N_29948,N_28266,N_28844);
nor U29949 (N_29949,N_28739,N_28921);
xnor U29950 (N_29950,N_28938,N_28681);
nor U29951 (N_29951,N_28799,N_28083);
nor U29952 (N_29952,N_28524,N_28871);
or U29953 (N_29953,N_28556,N_28416);
xor U29954 (N_29954,N_28174,N_28779);
or U29955 (N_29955,N_28892,N_28987);
nor U29956 (N_29956,N_28351,N_28602);
nor U29957 (N_29957,N_28658,N_28285);
xnor U29958 (N_29958,N_28358,N_28400);
and U29959 (N_29959,N_28412,N_28624);
xnor U29960 (N_29960,N_28415,N_28323);
or U29961 (N_29961,N_28972,N_28765);
nand U29962 (N_29962,N_28235,N_28798);
nor U29963 (N_29963,N_28713,N_28048);
nor U29964 (N_29964,N_28841,N_28363);
nand U29965 (N_29965,N_28569,N_28066);
xor U29966 (N_29966,N_28235,N_28599);
or U29967 (N_29967,N_28246,N_28403);
nand U29968 (N_29968,N_28087,N_28024);
nor U29969 (N_29969,N_28084,N_28593);
nand U29970 (N_29970,N_28316,N_28881);
nand U29971 (N_29971,N_28213,N_28538);
xnor U29972 (N_29972,N_28574,N_28049);
nand U29973 (N_29973,N_28592,N_28161);
and U29974 (N_29974,N_28639,N_28671);
xnor U29975 (N_29975,N_28321,N_28669);
and U29976 (N_29976,N_28425,N_28819);
or U29977 (N_29977,N_28025,N_28576);
xor U29978 (N_29978,N_28679,N_28235);
and U29979 (N_29979,N_28682,N_28979);
and U29980 (N_29980,N_28477,N_28697);
nor U29981 (N_29981,N_28524,N_28795);
xnor U29982 (N_29982,N_28633,N_28261);
or U29983 (N_29983,N_28732,N_28380);
nand U29984 (N_29984,N_28922,N_28130);
nor U29985 (N_29985,N_28259,N_28490);
and U29986 (N_29986,N_28304,N_28604);
nand U29987 (N_29987,N_28597,N_28887);
nor U29988 (N_29988,N_28334,N_28144);
and U29989 (N_29989,N_28355,N_28488);
nand U29990 (N_29990,N_28339,N_28754);
nor U29991 (N_29991,N_28183,N_28580);
xor U29992 (N_29992,N_28092,N_28416);
nand U29993 (N_29993,N_28153,N_28292);
and U29994 (N_29994,N_28600,N_28094);
xor U29995 (N_29995,N_28061,N_28437);
nor U29996 (N_29996,N_28894,N_28551);
nor U29997 (N_29997,N_28438,N_28142);
or U29998 (N_29998,N_28912,N_28848);
xnor U29999 (N_29999,N_28619,N_28582);
xor UO_0 (O_0,N_29695,N_29256);
nand UO_1 (O_1,N_29290,N_29633);
or UO_2 (O_2,N_29306,N_29229);
xor UO_3 (O_3,N_29706,N_29001);
nor UO_4 (O_4,N_29884,N_29462);
nor UO_5 (O_5,N_29682,N_29025);
nand UO_6 (O_6,N_29796,N_29645);
and UO_7 (O_7,N_29248,N_29745);
xnor UO_8 (O_8,N_29322,N_29039);
and UO_9 (O_9,N_29947,N_29576);
or UO_10 (O_10,N_29874,N_29662);
nor UO_11 (O_11,N_29658,N_29530);
or UO_12 (O_12,N_29062,N_29605);
and UO_13 (O_13,N_29054,N_29644);
and UO_14 (O_14,N_29035,N_29066);
and UO_15 (O_15,N_29582,N_29601);
xnor UO_16 (O_16,N_29751,N_29596);
or UO_17 (O_17,N_29474,N_29413);
and UO_18 (O_18,N_29034,N_29466);
nor UO_19 (O_19,N_29610,N_29259);
nor UO_20 (O_20,N_29908,N_29973);
or UO_21 (O_21,N_29059,N_29245);
nor UO_22 (O_22,N_29449,N_29443);
or UO_23 (O_23,N_29079,N_29611);
and UO_24 (O_24,N_29409,N_29758);
or UO_25 (O_25,N_29505,N_29102);
nand UO_26 (O_26,N_29371,N_29381);
nor UO_27 (O_27,N_29113,N_29261);
or UO_28 (O_28,N_29703,N_29196);
nand UO_29 (O_29,N_29497,N_29157);
xnor UO_30 (O_30,N_29429,N_29217);
or UO_31 (O_31,N_29845,N_29965);
nor UO_32 (O_32,N_29383,N_29628);
or UO_33 (O_33,N_29425,N_29395);
nand UO_34 (O_34,N_29327,N_29856);
nand UO_35 (O_35,N_29094,N_29617);
or UO_36 (O_36,N_29026,N_29643);
and UO_37 (O_37,N_29942,N_29360);
nand UO_38 (O_38,N_29233,N_29219);
or UO_39 (O_39,N_29971,N_29587);
xor UO_40 (O_40,N_29387,N_29069);
and UO_41 (O_41,N_29733,N_29927);
nand UO_42 (O_42,N_29201,N_29969);
xor UO_43 (O_43,N_29269,N_29777);
nand UO_44 (O_44,N_29657,N_29281);
nor UO_45 (O_45,N_29762,N_29549);
nor UO_46 (O_46,N_29406,N_29373);
xnor UO_47 (O_47,N_29844,N_29779);
and UO_48 (O_48,N_29095,N_29498);
and UO_49 (O_49,N_29347,N_29323);
xnor UO_50 (O_50,N_29535,N_29980);
nand UO_51 (O_51,N_29393,N_29366);
nor UO_52 (O_52,N_29647,N_29590);
or UO_53 (O_53,N_29895,N_29005);
xor UO_54 (O_54,N_29129,N_29548);
or UO_55 (O_55,N_29053,N_29822);
xnor UO_56 (O_56,N_29485,N_29194);
xnor UO_57 (O_57,N_29080,N_29048);
nand UO_58 (O_58,N_29835,N_29468);
nand UO_59 (O_59,N_29921,N_29382);
and UO_60 (O_60,N_29769,N_29679);
and UO_61 (O_61,N_29190,N_29709);
or UO_62 (O_62,N_29283,N_29834);
or UO_63 (O_63,N_29532,N_29772);
xor UO_64 (O_64,N_29586,N_29782);
nor UO_65 (O_65,N_29197,N_29631);
nand UO_66 (O_66,N_29184,N_29896);
nor UO_67 (O_67,N_29447,N_29802);
nand UO_68 (O_68,N_29038,N_29188);
or UO_69 (O_69,N_29791,N_29220);
nor UO_70 (O_70,N_29700,N_29664);
nand UO_71 (O_71,N_29369,N_29930);
nand UO_72 (O_72,N_29433,N_29206);
or UO_73 (O_73,N_29148,N_29444);
xnor UO_74 (O_74,N_29212,N_29492);
and UO_75 (O_75,N_29952,N_29132);
or UO_76 (O_76,N_29082,N_29254);
or UO_77 (O_77,N_29356,N_29391);
nor UO_78 (O_78,N_29008,N_29678);
xnor UO_79 (O_79,N_29746,N_29002);
nor UO_80 (O_80,N_29508,N_29367);
or UO_81 (O_81,N_29031,N_29959);
or UO_82 (O_82,N_29340,N_29686);
nor UO_83 (O_83,N_29307,N_29108);
nand UO_84 (O_84,N_29117,N_29096);
nand UO_85 (O_85,N_29236,N_29422);
nor UO_86 (O_86,N_29512,N_29516);
and UO_87 (O_87,N_29408,N_29978);
nor UO_88 (O_88,N_29774,N_29636);
xor UO_89 (O_89,N_29618,N_29321);
xor UO_90 (O_90,N_29208,N_29260);
xor UO_91 (O_91,N_29264,N_29150);
nand UO_92 (O_92,N_29226,N_29007);
xor UO_93 (O_93,N_29024,N_29640);
xnor UO_94 (O_94,N_29670,N_29228);
or UO_95 (O_95,N_29421,N_29883);
xor UO_96 (O_96,N_29339,N_29882);
nand UO_97 (O_97,N_29297,N_29519);
xor UO_98 (O_98,N_29893,N_29126);
nor UO_99 (O_99,N_29503,N_29881);
nor UO_100 (O_100,N_29575,N_29250);
and UO_101 (O_101,N_29140,N_29593);
nor UO_102 (O_102,N_29534,N_29727);
or UO_103 (O_103,N_29273,N_29302);
xor UO_104 (O_104,N_29017,N_29651);
or UO_105 (O_105,N_29903,N_29546);
nor UO_106 (O_106,N_29225,N_29081);
nor UO_107 (O_107,N_29583,N_29011);
and UO_108 (O_108,N_29814,N_29098);
nand UO_109 (O_109,N_29487,N_29389);
nor UO_110 (O_110,N_29115,N_29699);
and UO_111 (O_111,N_29850,N_29671);
nand UO_112 (O_112,N_29456,N_29704);
or UO_113 (O_113,N_29757,N_29010);
and UO_114 (O_114,N_29213,N_29013);
nand UO_115 (O_115,N_29486,N_29730);
nor UO_116 (O_116,N_29402,N_29571);
and UO_117 (O_117,N_29763,N_29146);
nor UO_118 (O_118,N_29130,N_29860);
and UO_119 (O_119,N_29142,N_29904);
nand UO_120 (O_120,N_29055,N_29825);
or UO_121 (O_121,N_29067,N_29049);
nand UO_122 (O_122,N_29337,N_29171);
nor UO_123 (O_123,N_29813,N_29780);
nand UO_124 (O_124,N_29613,N_29314);
and UO_125 (O_125,N_29285,N_29328);
nand UO_126 (O_126,N_29318,N_29705);
nand UO_127 (O_127,N_29278,N_29405);
nor UO_128 (O_128,N_29642,N_29623);
and UO_129 (O_129,N_29070,N_29615);
xor UO_130 (O_130,N_29204,N_29713);
nor UO_131 (O_131,N_29205,N_29821);
nand UO_132 (O_132,N_29114,N_29165);
nand UO_133 (O_133,N_29607,N_29974);
nor UO_134 (O_134,N_29877,N_29654);
and UO_135 (O_135,N_29159,N_29370);
and UO_136 (O_136,N_29787,N_29394);
nand UO_137 (O_137,N_29385,N_29364);
and UO_138 (O_138,N_29805,N_29175);
or UO_139 (O_139,N_29710,N_29771);
and UO_140 (O_140,N_29475,N_29119);
or UO_141 (O_141,N_29224,N_29725);
or UO_142 (O_142,N_29920,N_29831);
nand UO_143 (O_143,N_29798,N_29101);
and UO_144 (O_144,N_29040,N_29263);
nor UO_145 (O_145,N_29870,N_29392);
and UO_146 (O_146,N_29180,N_29346);
xor UO_147 (O_147,N_29917,N_29543);
or UO_148 (O_148,N_29690,N_29953);
nand UO_149 (O_149,N_29694,N_29450);
nand UO_150 (O_150,N_29818,N_29766);
nand UO_151 (O_151,N_29234,N_29741);
or UO_152 (O_152,N_29423,N_29153);
and UO_153 (O_153,N_29279,N_29215);
and UO_154 (O_154,N_29961,N_29437);
and UO_155 (O_155,N_29313,N_29811);
and UO_156 (O_156,N_29262,N_29178);
and UO_157 (O_157,N_29134,N_29830);
or UO_158 (O_158,N_29889,N_29941);
nor UO_159 (O_159,N_29970,N_29430);
nand UO_160 (O_160,N_29529,N_29734);
nand UO_161 (O_161,N_29252,N_29324);
and UO_162 (O_162,N_29399,N_29111);
nand UO_163 (O_163,N_29300,N_29442);
xnor UO_164 (O_164,N_29926,N_29990);
or UO_165 (O_165,N_29265,N_29750);
xnor UO_166 (O_166,N_29648,N_29698);
and UO_167 (O_167,N_29832,N_29077);
nand UO_168 (O_168,N_29723,N_29398);
nor UO_169 (O_169,N_29085,N_29925);
or UO_170 (O_170,N_29992,N_29354);
and UO_171 (O_171,N_29143,N_29988);
and UO_172 (O_172,N_29918,N_29783);
nand UO_173 (O_173,N_29088,N_29464);
or UO_174 (O_174,N_29149,N_29849);
or UO_175 (O_175,N_29985,N_29557);
or UO_176 (O_176,N_29473,N_29414);
or UO_177 (O_177,N_29268,N_29815);
xor UO_178 (O_178,N_29072,N_29790);
nand UO_179 (O_179,N_29600,N_29445);
and UO_180 (O_180,N_29014,N_29739);
and UO_181 (O_181,N_29438,N_29674);
or UO_182 (O_182,N_29198,N_29871);
or UO_183 (O_183,N_29491,N_29786);
or UO_184 (O_184,N_29998,N_29736);
nand UO_185 (O_185,N_29460,N_29416);
and UO_186 (O_186,N_29968,N_29781);
nor UO_187 (O_187,N_29488,N_29312);
or UO_188 (O_188,N_29355,N_29192);
xnor UO_189 (O_189,N_29606,N_29552);
or UO_190 (O_190,N_29501,N_29493);
xnor UO_191 (O_191,N_29520,N_29632);
xnor UO_192 (O_192,N_29076,N_29037);
or UO_193 (O_193,N_29086,N_29218);
nor UO_194 (O_194,N_29045,N_29061);
xor UO_195 (O_195,N_29894,N_29139);
xnor UO_196 (O_196,N_29060,N_29227);
or UO_197 (O_197,N_29960,N_29826);
nor UO_198 (O_198,N_29851,N_29022);
or UO_199 (O_199,N_29480,N_29897);
xor UO_200 (O_200,N_29484,N_29465);
and UO_201 (O_201,N_29839,N_29743);
xor UO_202 (O_202,N_29057,N_29342);
xor UO_203 (O_203,N_29122,N_29044);
nor UO_204 (O_204,N_29999,N_29905);
xor UO_205 (O_205,N_29513,N_29428);
xor UO_206 (O_206,N_29431,N_29345);
or UO_207 (O_207,N_29418,N_29351);
or UO_208 (O_208,N_29625,N_29363);
or UO_209 (O_209,N_29829,N_29544);
xor UO_210 (O_210,N_29560,N_29740);
or UO_211 (O_211,N_29052,N_29434);
or UO_212 (O_212,N_29556,N_29804);
or UO_213 (O_213,N_29847,N_29004);
nand UO_214 (O_214,N_29716,N_29246);
xor UO_215 (O_215,N_29809,N_29685);
nor UO_216 (O_216,N_29099,N_29158);
xor UO_217 (O_217,N_29656,N_29731);
or UO_218 (O_218,N_29420,N_29435);
xnor UO_219 (O_219,N_29838,N_29187);
nor UO_220 (O_220,N_29693,N_29331);
xor UO_221 (O_221,N_29352,N_29732);
or UO_222 (O_222,N_29304,N_29275);
or UO_223 (O_223,N_29711,N_29580);
or UO_224 (O_224,N_29914,N_29368);
xor UO_225 (O_225,N_29778,N_29043);
xor UO_226 (O_226,N_29471,N_29030);
xor UO_227 (O_227,N_29928,N_29608);
and UO_228 (O_228,N_29888,N_29987);
nor UO_229 (O_229,N_29193,N_29511);
nor UO_230 (O_230,N_29329,N_29948);
nor UO_231 (O_231,N_29050,N_29979);
nor UO_232 (O_232,N_29000,N_29274);
and UO_233 (O_233,N_29993,N_29752);
and UO_234 (O_234,N_29164,N_29154);
nand UO_235 (O_235,N_29595,N_29846);
nand UO_236 (O_236,N_29841,N_29317);
nor UO_237 (O_237,N_29292,N_29189);
xnor UO_238 (O_238,N_29046,N_29715);
xnor UO_239 (O_239,N_29842,N_29490);
nand UO_240 (O_240,N_29110,N_29604);
nor UO_241 (O_241,N_29966,N_29997);
nand UO_242 (O_242,N_29909,N_29879);
nor UO_243 (O_243,N_29962,N_29564);
nor UO_244 (O_244,N_29287,N_29946);
or UO_245 (O_245,N_29559,N_29121);
or UO_246 (O_246,N_29691,N_29852);
nor UO_247 (O_247,N_29963,N_29932);
or UO_248 (O_248,N_29477,N_29019);
nor UO_249 (O_249,N_29986,N_29714);
and UO_250 (O_250,N_29463,N_29074);
nor UO_251 (O_251,N_29799,N_29202);
nor UO_252 (O_252,N_29326,N_29308);
and UO_253 (O_253,N_29956,N_29989);
xnor UO_254 (O_254,N_29334,N_29854);
and UO_255 (O_255,N_29768,N_29358);
nor UO_256 (O_256,N_29561,N_29181);
nor UO_257 (O_257,N_29996,N_29721);
and UO_258 (O_258,N_29012,N_29380);
nand UO_259 (O_259,N_29761,N_29824);
nor UO_260 (O_260,N_29770,N_29609);
xor UO_261 (O_261,N_29124,N_29892);
nand UO_262 (O_262,N_29350,N_29539);
nand UO_263 (O_263,N_29319,N_29288);
nand UO_264 (O_264,N_29955,N_29286);
or UO_265 (O_265,N_29021,N_29820);
xnor UO_266 (O_266,N_29837,N_29667);
and UO_267 (O_267,N_29843,N_29396);
or UO_268 (O_268,N_29665,N_29807);
nor UO_269 (O_269,N_29898,N_29502);
xnor UO_270 (O_270,N_29507,N_29784);
and UO_271 (O_271,N_29934,N_29776);
and UO_272 (O_272,N_29470,N_29362);
or UO_273 (O_273,N_29147,N_29090);
xnor UO_274 (O_274,N_29467,N_29775);
xor UO_275 (O_275,N_29424,N_29239);
or UO_276 (O_276,N_29943,N_29554);
xnor UO_277 (O_277,N_29537,N_29602);
and UO_278 (O_278,N_29170,N_29689);
xnor UO_279 (O_279,N_29562,N_29816);
xor UO_280 (O_280,N_29296,N_29375);
or UO_281 (O_281,N_29104,N_29855);
or UO_282 (O_282,N_29598,N_29106);
and UO_283 (O_283,N_29680,N_29812);
or UO_284 (O_284,N_29128,N_29747);
nor UO_285 (O_285,N_29630,N_29504);
nand UO_286 (O_286,N_29759,N_29634);
nand UO_287 (O_287,N_29167,N_29144);
nor UO_288 (O_288,N_29627,N_29808);
and UO_289 (O_289,N_29517,N_29541);
nor UO_290 (O_290,N_29301,N_29748);
nor UO_291 (O_291,N_29828,N_29801);
and UO_292 (O_292,N_29717,N_29599);
xor UO_293 (O_293,N_29635,N_29091);
or UO_294 (O_294,N_29793,N_29168);
nand UO_295 (O_295,N_29570,N_29173);
xor UO_296 (O_296,N_29100,N_29440);
and UO_297 (O_297,N_29071,N_29016);
nor UO_298 (O_298,N_29675,N_29078);
or UO_299 (O_299,N_29489,N_29255);
nor UO_300 (O_300,N_29047,N_29325);
or UO_301 (O_301,N_29857,N_29869);
nor UO_302 (O_302,N_29868,N_29116);
nand UO_303 (O_303,N_29075,N_29199);
nor UO_304 (O_304,N_29872,N_29336);
and UO_305 (O_305,N_29472,N_29744);
xnor UO_306 (O_306,N_29311,N_29027);
and UO_307 (O_307,N_29668,N_29683);
and UO_308 (O_308,N_29298,N_29861);
or UO_309 (O_309,N_29994,N_29103);
nand UO_310 (O_310,N_29885,N_29840);
xnor UO_311 (O_311,N_29588,N_29257);
nor UO_312 (O_312,N_29803,N_29912);
nor UO_313 (O_313,N_29753,N_29064);
xnor UO_314 (O_314,N_29901,N_29120);
nand UO_315 (O_315,N_29379,N_29145);
and UO_316 (O_316,N_29616,N_29289);
xnor UO_317 (O_317,N_29481,N_29692);
or UO_318 (O_318,N_29003,N_29891);
and UO_319 (O_319,N_29403,N_29890);
nand UO_320 (O_320,N_29374,N_29887);
or UO_321 (O_321,N_29669,N_29823);
xor UO_322 (O_322,N_29163,N_29911);
or UO_323 (O_323,N_29722,N_29267);
nor UO_324 (O_324,N_29320,N_29310);
or UO_325 (O_325,N_29899,N_29247);
nor UO_326 (O_326,N_29578,N_29315);
and UO_327 (O_327,N_29726,N_29388);
nand UO_328 (O_328,N_29641,N_29957);
nand UO_329 (O_329,N_29365,N_29191);
or UO_330 (O_330,N_29230,N_29677);
nand UO_331 (O_331,N_29975,N_29929);
and UO_332 (O_332,N_29496,N_29333);
or UO_333 (O_333,N_29087,N_29410);
nand UO_334 (O_334,N_29574,N_29185);
or UO_335 (O_335,N_29880,N_29451);
xor UO_336 (O_336,N_29266,N_29036);
or UO_337 (O_337,N_29672,N_29933);
nand UO_338 (O_338,N_29951,N_29810);
nand UO_339 (O_339,N_29687,N_29935);
or UO_340 (O_340,N_29531,N_29702);
and UO_341 (O_341,N_29785,N_29419);
or UO_342 (O_342,N_29284,N_29125);
nand UO_343 (O_343,N_29506,N_29166);
nand UO_344 (O_344,N_29457,N_29299);
and UO_345 (O_345,N_29755,N_29523);
xor UO_346 (O_346,N_29084,N_29765);
nor UO_347 (O_347,N_29789,N_29461);
nand UO_348 (O_348,N_29684,N_29991);
or UO_349 (O_349,N_29728,N_29591);
and UO_350 (O_350,N_29660,N_29169);
nand UO_351 (O_351,N_29436,N_29231);
nor UO_352 (O_352,N_29967,N_29253);
or UO_353 (O_353,N_29981,N_29009);
and UO_354 (O_354,N_29131,N_29386);
or UO_355 (O_355,N_29524,N_29303);
nand UO_356 (O_356,N_29718,N_29873);
xor UO_357 (O_357,N_29162,N_29558);
xor UO_358 (O_358,N_29827,N_29833);
nand UO_359 (O_359,N_29384,N_29361);
nand UO_360 (O_360,N_29332,N_29650);
or UO_361 (O_361,N_29316,N_29545);
and UO_362 (O_362,N_29666,N_29209);
or UO_363 (O_363,N_29020,N_29764);
xor UO_364 (O_364,N_29910,N_29915);
and UO_365 (O_365,N_29754,N_29688);
and UO_366 (O_366,N_29742,N_29518);
and UO_367 (O_367,N_29063,N_29936);
nor UO_368 (O_368,N_29923,N_29540);
and UO_369 (O_369,N_29707,N_29448);
xor UO_370 (O_370,N_29652,N_29439);
xor UO_371 (O_371,N_29353,N_29309);
or UO_372 (O_372,N_29950,N_29377);
nor UO_373 (O_373,N_29417,N_29900);
and UO_374 (O_374,N_29876,N_29982);
nor UO_375 (O_375,N_29359,N_29089);
nand UO_376 (O_376,N_29214,N_29525);
xnor UO_377 (O_377,N_29294,N_29865);
xor UO_378 (O_378,N_29945,N_29673);
nand UO_379 (O_379,N_29696,N_29614);
or UO_380 (O_380,N_29156,N_29183);
and UO_381 (O_381,N_29788,N_29152);
nor UO_382 (O_382,N_29984,N_29579);
and UO_383 (O_383,N_29412,N_29092);
or UO_384 (O_384,N_29922,N_29767);
nor UO_385 (O_385,N_29724,N_29330);
nor UO_386 (O_386,N_29649,N_29565);
or UO_387 (O_387,N_29712,N_29051);
nor UO_388 (O_388,N_29944,N_29015);
nand UO_389 (O_389,N_29585,N_29795);
or UO_390 (O_390,N_29924,N_29182);
nor UO_391 (O_391,N_29568,N_29127);
nand UO_392 (O_392,N_29797,N_29172);
nor UO_393 (O_393,N_29338,N_29135);
nand UO_394 (O_394,N_29028,N_29240);
and UO_395 (O_395,N_29836,N_29573);
xnor UO_396 (O_396,N_29581,N_29863);
nor UO_397 (O_397,N_29729,N_29223);
xnor UO_398 (O_398,N_29629,N_29138);
xor UO_399 (O_399,N_29272,N_29577);
xnor UO_400 (O_400,N_29033,N_29536);
and UO_401 (O_401,N_29939,N_29109);
nor UO_402 (O_402,N_29211,N_29792);
and UO_403 (O_403,N_29136,N_29906);
xor UO_404 (O_404,N_29105,N_29902);
nand UO_405 (O_405,N_29749,N_29701);
xnor UO_406 (O_406,N_29348,N_29404);
nor UO_407 (O_407,N_29295,N_29452);
or UO_408 (O_408,N_29249,N_29042);
or UO_409 (O_409,N_29864,N_29232);
xnor UO_410 (O_410,N_29118,N_29859);
and UO_411 (O_411,N_29241,N_29235);
xnor UO_412 (O_412,N_29954,N_29773);
or UO_413 (O_413,N_29760,N_29141);
or UO_414 (O_414,N_29446,N_29553);
nand UO_415 (O_415,N_29862,N_29216);
or UO_416 (O_416,N_29478,N_29867);
nor UO_417 (O_417,N_29972,N_29238);
nor UO_418 (O_418,N_29006,N_29938);
and UO_419 (O_419,N_29343,N_29569);
and UO_420 (O_420,N_29174,N_29058);
and UO_421 (O_421,N_29794,N_29919);
nor UO_422 (O_422,N_29258,N_29555);
nor UO_423 (O_423,N_29547,N_29495);
nor UO_424 (O_424,N_29427,N_29029);
and UO_425 (O_425,N_29594,N_29756);
and UO_426 (O_426,N_29415,N_29200);
nor UO_427 (O_427,N_29976,N_29958);
xor UO_428 (O_428,N_29023,N_29293);
nand UO_429 (O_429,N_29372,N_29107);
and UO_430 (O_430,N_29179,N_29655);
xnor UO_431 (O_431,N_29376,N_29646);
xnor UO_432 (O_432,N_29663,N_29661);
and UO_433 (O_433,N_29597,N_29619);
and UO_434 (O_434,N_29277,N_29866);
nor UO_435 (O_435,N_29638,N_29551);
nor UO_436 (O_436,N_29515,N_29177);
nor UO_437 (O_437,N_29276,N_29800);
nor UO_438 (O_438,N_29572,N_29056);
and UO_439 (O_439,N_29068,N_29550);
nand UO_440 (O_440,N_29341,N_29995);
nor UO_441 (O_441,N_29563,N_29280);
and UO_442 (O_442,N_29291,N_29407);
nor UO_443 (O_443,N_29203,N_29401);
or UO_444 (O_444,N_29697,N_29708);
or UO_445 (O_445,N_29738,N_29542);
nor UO_446 (O_446,N_29032,N_29983);
nor UO_447 (O_447,N_29397,N_29411);
nand UO_448 (O_448,N_29521,N_29848);
nand UO_449 (O_449,N_29137,N_29858);
and UO_450 (O_450,N_29242,N_29526);
nor UO_451 (O_451,N_29509,N_29806);
nand UO_452 (O_452,N_29907,N_29186);
nand UO_453 (O_453,N_29612,N_29349);
nor UO_454 (O_454,N_29681,N_29949);
nand UO_455 (O_455,N_29237,N_29271);
xnor UO_456 (O_456,N_29018,N_29123);
nand UO_457 (O_457,N_29913,N_29878);
or UO_458 (O_458,N_29931,N_29305);
or UO_459 (O_459,N_29522,N_29916);
and UO_460 (O_460,N_29455,N_29528);
nor UO_461 (O_461,N_29426,N_29432);
nor UO_462 (O_462,N_29161,N_29160);
xor UO_463 (O_463,N_29817,N_29195);
and UO_464 (O_464,N_29494,N_29243);
or UO_465 (O_465,N_29222,N_29476);
and UO_466 (O_466,N_29112,N_29886);
nand UO_467 (O_467,N_29357,N_29735);
nand UO_468 (O_468,N_29875,N_29282);
nand UO_469 (O_469,N_29479,N_29603);
nor UO_470 (O_470,N_29176,N_29483);
or UO_471 (O_471,N_29400,N_29500);
xor UO_472 (O_472,N_29566,N_29533);
or UO_473 (O_473,N_29454,N_29653);
and UO_474 (O_474,N_29073,N_29207);
or UO_475 (O_475,N_29589,N_29527);
and UO_476 (O_476,N_29719,N_29083);
or UO_477 (O_477,N_29937,N_29221);
xor UO_478 (O_478,N_29621,N_29626);
and UO_479 (O_479,N_29065,N_29469);
nand UO_480 (O_480,N_29819,N_29499);
or UO_481 (O_481,N_29538,N_29335);
and UO_482 (O_482,N_29390,N_29097);
nand UO_483 (O_483,N_29964,N_29041);
nor UO_484 (O_484,N_29344,N_29720);
nor UO_485 (O_485,N_29639,N_29210);
nand UO_486 (O_486,N_29093,N_29482);
nand UO_487 (O_487,N_29155,N_29453);
or UO_488 (O_488,N_29151,N_29378);
nand UO_489 (O_489,N_29940,N_29676);
nor UO_490 (O_490,N_29244,N_29637);
nor UO_491 (O_491,N_29567,N_29622);
nor UO_492 (O_492,N_29270,N_29510);
nand UO_493 (O_493,N_29592,N_29737);
and UO_494 (O_494,N_29624,N_29659);
nand UO_495 (O_495,N_29620,N_29441);
nand UO_496 (O_496,N_29853,N_29584);
or UO_497 (O_497,N_29458,N_29459);
nand UO_498 (O_498,N_29514,N_29133);
nor UO_499 (O_499,N_29977,N_29251);
and UO_500 (O_500,N_29209,N_29759);
or UO_501 (O_501,N_29372,N_29955);
nor UO_502 (O_502,N_29249,N_29885);
nor UO_503 (O_503,N_29350,N_29229);
or UO_504 (O_504,N_29836,N_29727);
xnor UO_505 (O_505,N_29484,N_29970);
nor UO_506 (O_506,N_29976,N_29962);
nor UO_507 (O_507,N_29277,N_29149);
or UO_508 (O_508,N_29284,N_29900);
nand UO_509 (O_509,N_29472,N_29878);
and UO_510 (O_510,N_29575,N_29545);
or UO_511 (O_511,N_29258,N_29043);
xor UO_512 (O_512,N_29814,N_29594);
and UO_513 (O_513,N_29188,N_29800);
nand UO_514 (O_514,N_29550,N_29846);
or UO_515 (O_515,N_29721,N_29885);
or UO_516 (O_516,N_29658,N_29986);
and UO_517 (O_517,N_29095,N_29393);
and UO_518 (O_518,N_29982,N_29977);
nand UO_519 (O_519,N_29978,N_29839);
and UO_520 (O_520,N_29321,N_29546);
xor UO_521 (O_521,N_29477,N_29065);
or UO_522 (O_522,N_29676,N_29777);
xnor UO_523 (O_523,N_29943,N_29622);
xnor UO_524 (O_524,N_29524,N_29951);
nor UO_525 (O_525,N_29425,N_29840);
or UO_526 (O_526,N_29707,N_29294);
nor UO_527 (O_527,N_29362,N_29455);
nand UO_528 (O_528,N_29640,N_29888);
nand UO_529 (O_529,N_29218,N_29068);
nor UO_530 (O_530,N_29427,N_29409);
nand UO_531 (O_531,N_29828,N_29152);
xor UO_532 (O_532,N_29975,N_29536);
and UO_533 (O_533,N_29832,N_29058);
nor UO_534 (O_534,N_29150,N_29604);
or UO_535 (O_535,N_29478,N_29814);
nor UO_536 (O_536,N_29051,N_29176);
and UO_537 (O_537,N_29199,N_29287);
xor UO_538 (O_538,N_29908,N_29925);
nor UO_539 (O_539,N_29780,N_29803);
nand UO_540 (O_540,N_29769,N_29812);
nand UO_541 (O_541,N_29452,N_29606);
or UO_542 (O_542,N_29113,N_29856);
nor UO_543 (O_543,N_29589,N_29324);
nor UO_544 (O_544,N_29183,N_29378);
xnor UO_545 (O_545,N_29528,N_29729);
or UO_546 (O_546,N_29279,N_29663);
xnor UO_547 (O_547,N_29243,N_29067);
or UO_548 (O_548,N_29104,N_29785);
or UO_549 (O_549,N_29282,N_29477);
nand UO_550 (O_550,N_29204,N_29718);
xor UO_551 (O_551,N_29334,N_29183);
nor UO_552 (O_552,N_29071,N_29720);
or UO_553 (O_553,N_29340,N_29440);
xor UO_554 (O_554,N_29319,N_29714);
xnor UO_555 (O_555,N_29370,N_29448);
xor UO_556 (O_556,N_29440,N_29831);
and UO_557 (O_557,N_29261,N_29864);
or UO_558 (O_558,N_29143,N_29992);
nor UO_559 (O_559,N_29123,N_29735);
nand UO_560 (O_560,N_29768,N_29268);
nor UO_561 (O_561,N_29784,N_29061);
or UO_562 (O_562,N_29257,N_29340);
nor UO_563 (O_563,N_29437,N_29559);
xnor UO_564 (O_564,N_29683,N_29472);
or UO_565 (O_565,N_29726,N_29729);
and UO_566 (O_566,N_29861,N_29637);
nor UO_567 (O_567,N_29565,N_29940);
xor UO_568 (O_568,N_29989,N_29262);
or UO_569 (O_569,N_29135,N_29624);
nor UO_570 (O_570,N_29304,N_29165);
and UO_571 (O_571,N_29981,N_29722);
nand UO_572 (O_572,N_29770,N_29585);
nor UO_573 (O_573,N_29819,N_29082);
nor UO_574 (O_574,N_29400,N_29652);
nand UO_575 (O_575,N_29287,N_29892);
nand UO_576 (O_576,N_29129,N_29641);
nand UO_577 (O_577,N_29282,N_29869);
and UO_578 (O_578,N_29385,N_29887);
xor UO_579 (O_579,N_29053,N_29781);
nand UO_580 (O_580,N_29162,N_29475);
nand UO_581 (O_581,N_29156,N_29841);
xor UO_582 (O_582,N_29970,N_29203);
and UO_583 (O_583,N_29139,N_29847);
or UO_584 (O_584,N_29329,N_29910);
and UO_585 (O_585,N_29038,N_29247);
nand UO_586 (O_586,N_29601,N_29727);
nor UO_587 (O_587,N_29729,N_29920);
and UO_588 (O_588,N_29231,N_29166);
nor UO_589 (O_589,N_29499,N_29239);
and UO_590 (O_590,N_29812,N_29029);
or UO_591 (O_591,N_29890,N_29805);
and UO_592 (O_592,N_29230,N_29586);
nor UO_593 (O_593,N_29946,N_29298);
or UO_594 (O_594,N_29751,N_29867);
nor UO_595 (O_595,N_29186,N_29004);
xor UO_596 (O_596,N_29834,N_29224);
and UO_597 (O_597,N_29082,N_29258);
xor UO_598 (O_598,N_29280,N_29777);
nor UO_599 (O_599,N_29236,N_29309);
nor UO_600 (O_600,N_29118,N_29188);
or UO_601 (O_601,N_29971,N_29781);
nor UO_602 (O_602,N_29575,N_29193);
nand UO_603 (O_603,N_29273,N_29268);
or UO_604 (O_604,N_29309,N_29347);
xor UO_605 (O_605,N_29092,N_29231);
or UO_606 (O_606,N_29769,N_29088);
or UO_607 (O_607,N_29536,N_29501);
and UO_608 (O_608,N_29848,N_29397);
nand UO_609 (O_609,N_29330,N_29380);
nand UO_610 (O_610,N_29222,N_29032);
nor UO_611 (O_611,N_29307,N_29838);
xnor UO_612 (O_612,N_29710,N_29294);
and UO_613 (O_613,N_29645,N_29667);
nand UO_614 (O_614,N_29307,N_29336);
nor UO_615 (O_615,N_29471,N_29614);
nor UO_616 (O_616,N_29945,N_29786);
or UO_617 (O_617,N_29426,N_29610);
xor UO_618 (O_618,N_29129,N_29807);
nand UO_619 (O_619,N_29124,N_29725);
and UO_620 (O_620,N_29506,N_29363);
and UO_621 (O_621,N_29727,N_29029);
and UO_622 (O_622,N_29771,N_29459);
xor UO_623 (O_623,N_29145,N_29611);
nand UO_624 (O_624,N_29172,N_29175);
or UO_625 (O_625,N_29007,N_29572);
xor UO_626 (O_626,N_29972,N_29148);
or UO_627 (O_627,N_29236,N_29560);
xnor UO_628 (O_628,N_29464,N_29389);
xor UO_629 (O_629,N_29489,N_29355);
nor UO_630 (O_630,N_29985,N_29054);
or UO_631 (O_631,N_29021,N_29992);
or UO_632 (O_632,N_29638,N_29565);
nor UO_633 (O_633,N_29448,N_29556);
and UO_634 (O_634,N_29481,N_29071);
nand UO_635 (O_635,N_29657,N_29969);
or UO_636 (O_636,N_29446,N_29691);
nand UO_637 (O_637,N_29103,N_29367);
or UO_638 (O_638,N_29192,N_29271);
xor UO_639 (O_639,N_29290,N_29150);
nor UO_640 (O_640,N_29057,N_29217);
xor UO_641 (O_641,N_29617,N_29654);
nand UO_642 (O_642,N_29127,N_29359);
and UO_643 (O_643,N_29122,N_29780);
or UO_644 (O_644,N_29050,N_29051);
or UO_645 (O_645,N_29963,N_29612);
nor UO_646 (O_646,N_29069,N_29216);
and UO_647 (O_647,N_29531,N_29259);
xnor UO_648 (O_648,N_29421,N_29332);
nand UO_649 (O_649,N_29184,N_29419);
xor UO_650 (O_650,N_29126,N_29212);
or UO_651 (O_651,N_29112,N_29557);
or UO_652 (O_652,N_29285,N_29781);
nor UO_653 (O_653,N_29821,N_29596);
xor UO_654 (O_654,N_29746,N_29969);
nand UO_655 (O_655,N_29332,N_29187);
xor UO_656 (O_656,N_29837,N_29411);
or UO_657 (O_657,N_29708,N_29489);
nand UO_658 (O_658,N_29427,N_29608);
xnor UO_659 (O_659,N_29933,N_29276);
xor UO_660 (O_660,N_29892,N_29109);
or UO_661 (O_661,N_29877,N_29010);
or UO_662 (O_662,N_29726,N_29761);
xor UO_663 (O_663,N_29403,N_29533);
nor UO_664 (O_664,N_29148,N_29950);
nand UO_665 (O_665,N_29635,N_29580);
nand UO_666 (O_666,N_29020,N_29905);
nor UO_667 (O_667,N_29228,N_29426);
nand UO_668 (O_668,N_29875,N_29664);
xnor UO_669 (O_669,N_29934,N_29520);
nand UO_670 (O_670,N_29347,N_29993);
or UO_671 (O_671,N_29903,N_29008);
or UO_672 (O_672,N_29960,N_29644);
nand UO_673 (O_673,N_29290,N_29688);
nand UO_674 (O_674,N_29693,N_29502);
and UO_675 (O_675,N_29408,N_29156);
xnor UO_676 (O_676,N_29761,N_29882);
nand UO_677 (O_677,N_29855,N_29846);
or UO_678 (O_678,N_29168,N_29039);
and UO_679 (O_679,N_29702,N_29170);
nand UO_680 (O_680,N_29708,N_29446);
nor UO_681 (O_681,N_29807,N_29716);
and UO_682 (O_682,N_29988,N_29549);
nor UO_683 (O_683,N_29390,N_29468);
and UO_684 (O_684,N_29637,N_29590);
nor UO_685 (O_685,N_29372,N_29189);
nor UO_686 (O_686,N_29205,N_29359);
nand UO_687 (O_687,N_29301,N_29832);
or UO_688 (O_688,N_29595,N_29203);
and UO_689 (O_689,N_29547,N_29191);
and UO_690 (O_690,N_29446,N_29088);
xor UO_691 (O_691,N_29394,N_29371);
or UO_692 (O_692,N_29410,N_29047);
and UO_693 (O_693,N_29037,N_29787);
nor UO_694 (O_694,N_29419,N_29991);
nor UO_695 (O_695,N_29042,N_29946);
nand UO_696 (O_696,N_29725,N_29444);
or UO_697 (O_697,N_29103,N_29997);
and UO_698 (O_698,N_29312,N_29229);
and UO_699 (O_699,N_29866,N_29392);
xnor UO_700 (O_700,N_29025,N_29388);
nor UO_701 (O_701,N_29910,N_29693);
and UO_702 (O_702,N_29364,N_29462);
xnor UO_703 (O_703,N_29889,N_29667);
or UO_704 (O_704,N_29698,N_29602);
nor UO_705 (O_705,N_29655,N_29027);
nand UO_706 (O_706,N_29822,N_29710);
or UO_707 (O_707,N_29064,N_29863);
or UO_708 (O_708,N_29295,N_29803);
xor UO_709 (O_709,N_29551,N_29469);
nor UO_710 (O_710,N_29759,N_29860);
xnor UO_711 (O_711,N_29410,N_29853);
or UO_712 (O_712,N_29746,N_29156);
or UO_713 (O_713,N_29575,N_29936);
or UO_714 (O_714,N_29625,N_29376);
xnor UO_715 (O_715,N_29589,N_29377);
nand UO_716 (O_716,N_29272,N_29562);
xnor UO_717 (O_717,N_29530,N_29182);
xnor UO_718 (O_718,N_29248,N_29287);
nand UO_719 (O_719,N_29294,N_29980);
and UO_720 (O_720,N_29261,N_29850);
or UO_721 (O_721,N_29259,N_29854);
and UO_722 (O_722,N_29292,N_29196);
nand UO_723 (O_723,N_29925,N_29478);
and UO_724 (O_724,N_29222,N_29503);
xor UO_725 (O_725,N_29948,N_29724);
nand UO_726 (O_726,N_29537,N_29786);
or UO_727 (O_727,N_29070,N_29227);
xor UO_728 (O_728,N_29412,N_29202);
or UO_729 (O_729,N_29276,N_29590);
and UO_730 (O_730,N_29036,N_29899);
xnor UO_731 (O_731,N_29915,N_29824);
and UO_732 (O_732,N_29732,N_29608);
xnor UO_733 (O_733,N_29728,N_29664);
and UO_734 (O_734,N_29903,N_29635);
nor UO_735 (O_735,N_29532,N_29866);
xnor UO_736 (O_736,N_29749,N_29452);
or UO_737 (O_737,N_29679,N_29671);
or UO_738 (O_738,N_29035,N_29824);
and UO_739 (O_739,N_29660,N_29062);
nand UO_740 (O_740,N_29844,N_29494);
or UO_741 (O_741,N_29243,N_29849);
nor UO_742 (O_742,N_29272,N_29063);
or UO_743 (O_743,N_29656,N_29473);
xnor UO_744 (O_744,N_29557,N_29114);
nor UO_745 (O_745,N_29086,N_29592);
nand UO_746 (O_746,N_29817,N_29794);
nand UO_747 (O_747,N_29268,N_29448);
xnor UO_748 (O_748,N_29828,N_29573);
or UO_749 (O_749,N_29690,N_29074);
xnor UO_750 (O_750,N_29283,N_29188);
nor UO_751 (O_751,N_29077,N_29169);
xnor UO_752 (O_752,N_29769,N_29772);
nand UO_753 (O_753,N_29087,N_29908);
nand UO_754 (O_754,N_29820,N_29794);
xnor UO_755 (O_755,N_29860,N_29178);
and UO_756 (O_756,N_29621,N_29756);
nor UO_757 (O_757,N_29362,N_29508);
nand UO_758 (O_758,N_29926,N_29573);
xor UO_759 (O_759,N_29595,N_29660);
xor UO_760 (O_760,N_29262,N_29260);
and UO_761 (O_761,N_29137,N_29772);
and UO_762 (O_762,N_29062,N_29478);
and UO_763 (O_763,N_29095,N_29199);
xnor UO_764 (O_764,N_29464,N_29240);
and UO_765 (O_765,N_29396,N_29685);
nand UO_766 (O_766,N_29447,N_29894);
nor UO_767 (O_767,N_29662,N_29438);
and UO_768 (O_768,N_29323,N_29199);
xnor UO_769 (O_769,N_29440,N_29981);
or UO_770 (O_770,N_29302,N_29018);
nand UO_771 (O_771,N_29386,N_29976);
nand UO_772 (O_772,N_29327,N_29299);
xnor UO_773 (O_773,N_29788,N_29015);
or UO_774 (O_774,N_29790,N_29989);
nor UO_775 (O_775,N_29523,N_29049);
nand UO_776 (O_776,N_29596,N_29261);
or UO_777 (O_777,N_29860,N_29686);
or UO_778 (O_778,N_29557,N_29973);
and UO_779 (O_779,N_29714,N_29789);
nor UO_780 (O_780,N_29854,N_29458);
or UO_781 (O_781,N_29576,N_29535);
xor UO_782 (O_782,N_29172,N_29642);
xnor UO_783 (O_783,N_29536,N_29649);
nand UO_784 (O_784,N_29977,N_29044);
nand UO_785 (O_785,N_29820,N_29779);
nand UO_786 (O_786,N_29844,N_29714);
or UO_787 (O_787,N_29971,N_29009);
xor UO_788 (O_788,N_29843,N_29641);
xnor UO_789 (O_789,N_29654,N_29861);
and UO_790 (O_790,N_29304,N_29200);
or UO_791 (O_791,N_29924,N_29684);
or UO_792 (O_792,N_29164,N_29147);
or UO_793 (O_793,N_29223,N_29024);
nor UO_794 (O_794,N_29907,N_29139);
and UO_795 (O_795,N_29765,N_29008);
xnor UO_796 (O_796,N_29151,N_29802);
nand UO_797 (O_797,N_29924,N_29694);
nand UO_798 (O_798,N_29563,N_29063);
and UO_799 (O_799,N_29379,N_29712);
nor UO_800 (O_800,N_29866,N_29758);
nand UO_801 (O_801,N_29169,N_29197);
or UO_802 (O_802,N_29797,N_29538);
nor UO_803 (O_803,N_29843,N_29689);
nor UO_804 (O_804,N_29185,N_29092);
nand UO_805 (O_805,N_29944,N_29143);
or UO_806 (O_806,N_29844,N_29833);
or UO_807 (O_807,N_29762,N_29764);
and UO_808 (O_808,N_29842,N_29457);
nand UO_809 (O_809,N_29980,N_29945);
nand UO_810 (O_810,N_29820,N_29851);
nor UO_811 (O_811,N_29397,N_29268);
or UO_812 (O_812,N_29411,N_29774);
xor UO_813 (O_813,N_29771,N_29920);
nor UO_814 (O_814,N_29594,N_29060);
xor UO_815 (O_815,N_29611,N_29065);
xnor UO_816 (O_816,N_29578,N_29027);
xnor UO_817 (O_817,N_29322,N_29709);
and UO_818 (O_818,N_29291,N_29885);
and UO_819 (O_819,N_29230,N_29657);
nor UO_820 (O_820,N_29961,N_29470);
or UO_821 (O_821,N_29619,N_29813);
and UO_822 (O_822,N_29360,N_29707);
nand UO_823 (O_823,N_29868,N_29896);
nand UO_824 (O_824,N_29981,N_29668);
nor UO_825 (O_825,N_29719,N_29169);
or UO_826 (O_826,N_29269,N_29055);
xor UO_827 (O_827,N_29005,N_29231);
and UO_828 (O_828,N_29997,N_29357);
nor UO_829 (O_829,N_29752,N_29466);
and UO_830 (O_830,N_29646,N_29627);
nand UO_831 (O_831,N_29798,N_29147);
and UO_832 (O_832,N_29898,N_29837);
or UO_833 (O_833,N_29845,N_29440);
nand UO_834 (O_834,N_29167,N_29579);
or UO_835 (O_835,N_29691,N_29504);
or UO_836 (O_836,N_29197,N_29618);
or UO_837 (O_837,N_29504,N_29566);
or UO_838 (O_838,N_29578,N_29256);
xor UO_839 (O_839,N_29914,N_29867);
xnor UO_840 (O_840,N_29445,N_29647);
xor UO_841 (O_841,N_29211,N_29724);
or UO_842 (O_842,N_29323,N_29050);
and UO_843 (O_843,N_29671,N_29673);
or UO_844 (O_844,N_29595,N_29775);
and UO_845 (O_845,N_29104,N_29121);
nor UO_846 (O_846,N_29707,N_29700);
nand UO_847 (O_847,N_29589,N_29288);
xor UO_848 (O_848,N_29563,N_29149);
xnor UO_849 (O_849,N_29804,N_29501);
xor UO_850 (O_850,N_29131,N_29521);
nand UO_851 (O_851,N_29772,N_29199);
or UO_852 (O_852,N_29155,N_29582);
nor UO_853 (O_853,N_29025,N_29407);
and UO_854 (O_854,N_29841,N_29383);
nor UO_855 (O_855,N_29255,N_29024);
xnor UO_856 (O_856,N_29917,N_29293);
xnor UO_857 (O_857,N_29926,N_29867);
and UO_858 (O_858,N_29033,N_29742);
xor UO_859 (O_859,N_29256,N_29328);
xnor UO_860 (O_860,N_29300,N_29772);
nor UO_861 (O_861,N_29199,N_29266);
xor UO_862 (O_862,N_29307,N_29994);
xor UO_863 (O_863,N_29797,N_29133);
and UO_864 (O_864,N_29058,N_29231);
nand UO_865 (O_865,N_29872,N_29923);
and UO_866 (O_866,N_29153,N_29506);
nand UO_867 (O_867,N_29956,N_29643);
nor UO_868 (O_868,N_29637,N_29666);
nor UO_869 (O_869,N_29529,N_29237);
xor UO_870 (O_870,N_29620,N_29315);
nand UO_871 (O_871,N_29733,N_29161);
nand UO_872 (O_872,N_29165,N_29803);
or UO_873 (O_873,N_29475,N_29472);
nand UO_874 (O_874,N_29439,N_29175);
or UO_875 (O_875,N_29280,N_29377);
xnor UO_876 (O_876,N_29780,N_29241);
nor UO_877 (O_877,N_29183,N_29209);
nand UO_878 (O_878,N_29320,N_29712);
nor UO_879 (O_879,N_29063,N_29137);
xor UO_880 (O_880,N_29912,N_29191);
xnor UO_881 (O_881,N_29338,N_29239);
and UO_882 (O_882,N_29203,N_29603);
or UO_883 (O_883,N_29795,N_29173);
or UO_884 (O_884,N_29110,N_29483);
nor UO_885 (O_885,N_29771,N_29128);
and UO_886 (O_886,N_29864,N_29407);
xor UO_887 (O_887,N_29521,N_29786);
and UO_888 (O_888,N_29799,N_29116);
or UO_889 (O_889,N_29015,N_29459);
xnor UO_890 (O_890,N_29135,N_29647);
xnor UO_891 (O_891,N_29441,N_29761);
and UO_892 (O_892,N_29425,N_29909);
nor UO_893 (O_893,N_29290,N_29746);
nand UO_894 (O_894,N_29968,N_29228);
or UO_895 (O_895,N_29552,N_29105);
and UO_896 (O_896,N_29590,N_29667);
nor UO_897 (O_897,N_29736,N_29945);
and UO_898 (O_898,N_29698,N_29424);
nor UO_899 (O_899,N_29449,N_29540);
or UO_900 (O_900,N_29630,N_29750);
and UO_901 (O_901,N_29307,N_29573);
and UO_902 (O_902,N_29498,N_29511);
nand UO_903 (O_903,N_29983,N_29481);
xnor UO_904 (O_904,N_29243,N_29544);
and UO_905 (O_905,N_29051,N_29239);
or UO_906 (O_906,N_29596,N_29585);
nand UO_907 (O_907,N_29985,N_29085);
or UO_908 (O_908,N_29932,N_29625);
and UO_909 (O_909,N_29840,N_29138);
or UO_910 (O_910,N_29773,N_29475);
xnor UO_911 (O_911,N_29528,N_29453);
and UO_912 (O_912,N_29569,N_29106);
nand UO_913 (O_913,N_29014,N_29548);
nand UO_914 (O_914,N_29596,N_29449);
nor UO_915 (O_915,N_29157,N_29117);
nor UO_916 (O_916,N_29338,N_29119);
nor UO_917 (O_917,N_29114,N_29863);
xor UO_918 (O_918,N_29383,N_29648);
nand UO_919 (O_919,N_29316,N_29566);
and UO_920 (O_920,N_29370,N_29898);
or UO_921 (O_921,N_29961,N_29504);
or UO_922 (O_922,N_29553,N_29462);
and UO_923 (O_923,N_29523,N_29240);
and UO_924 (O_924,N_29886,N_29260);
nand UO_925 (O_925,N_29126,N_29749);
nor UO_926 (O_926,N_29719,N_29933);
nand UO_927 (O_927,N_29947,N_29957);
xor UO_928 (O_928,N_29747,N_29851);
xnor UO_929 (O_929,N_29776,N_29699);
or UO_930 (O_930,N_29055,N_29963);
or UO_931 (O_931,N_29465,N_29623);
nand UO_932 (O_932,N_29043,N_29881);
and UO_933 (O_933,N_29154,N_29954);
xnor UO_934 (O_934,N_29293,N_29106);
nor UO_935 (O_935,N_29808,N_29671);
or UO_936 (O_936,N_29350,N_29650);
and UO_937 (O_937,N_29115,N_29526);
xor UO_938 (O_938,N_29400,N_29787);
or UO_939 (O_939,N_29515,N_29167);
or UO_940 (O_940,N_29030,N_29806);
and UO_941 (O_941,N_29564,N_29446);
nand UO_942 (O_942,N_29707,N_29074);
nand UO_943 (O_943,N_29901,N_29085);
or UO_944 (O_944,N_29052,N_29214);
xnor UO_945 (O_945,N_29997,N_29352);
or UO_946 (O_946,N_29634,N_29957);
and UO_947 (O_947,N_29237,N_29632);
xnor UO_948 (O_948,N_29654,N_29445);
nor UO_949 (O_949,N_29431,N_29054);
and UO_950 (O_950,N_29528,N_29586);
and UO_951 (O_951,N_29858,N_29555);
and UO_952 (O_952,N_29060,N_29437);
and UO_953 (O_953,N_29033,N_29570);
or UO_954 (O_954,N_29700,N_29742);
or UO_955 (O_955,N_29228,N_29832);
or UO_956 (O_956,N_29934,N_29007);
xnor UO_957 (O_957,N_29503,N_29298);
nor UO_958 (O_958,N_29334,N_29828);
nand UO_959 (O_959,N_29182,N_29724);
nand UO_960 (O_960,N_29687,N_29303);
and UO_961 (O_961,N_29457,N_29582);
xor UO_962 (O_962,N_29459,N_29465);
xnor UO_963 (O_963,N_29816,N_29036);
nand UO_964 (O_964,N_29935,N_29162);
xnor UO_965 (O_965,N_29087,N_29406);
or UO_966 (O_966,N_29724,N_29844);
and UO_967 (O_967,N_29527,N_29763);
or UO_968 (O_968,N_29325,N_29304);
nor UO_969 (O_969,N_29049,N_29895);
or UO_970 (O_970,N_29022,N_29606);
xnor UO_971 (O_971,N_29697,N_29352);
nand UO_972 (O_972,N_29926,N_29595);
nand UO_973 (O_973,N_29340,N_29205);
nand UO_974 (O_974,N_29598,N_29125);
nor UO_975 (O_975,N_29618,N_29672);
nor UO_976 (O_976,N_29448,N_29966);
or UO_977 (O_977,N_29260,N_29882);
xor UO_978 (O_978,N_29750,N_29405);
nor UO_979 (O_979,N_29177,N_29418);
xor UO_980 (O_980,N_29408,N_29370);
nand UO_981 (O_981,N_29978,N_29970);
or UO_982 (O_982,N_29187,N_29120);
nand UO_983 (O_983,N_29088,N_29856);
nor UO_984 (O_984,N_29620,N_29600);
or UO_985 (O_985,N_29483,N_29689);
or UO_986 (O_986,N_29870,N_29111);
and UO_987 (O_987,N_29811,N_29496);
xor UO_988 (O_988,N_29917,N_29612);
or UO_989 (O_989,N_29612,N_29368);
nand UO_990 (O_990,N_29225,N_29170);
xor UO_991 (O_991,N_29657,N_29319);
nor UO_992 (O_992,N_29919,N_29185);
or UO_993 (O_993,N_29400,N_29421);
and UO_994 (O_994,N_29836,N_29060);
or UO_995 (O_995,N_29339,N_29818);
or UO_996 (O_996,N_29133,N_29297);
xnor UO_997 (O_997,N_29890,N_29371);
and UO_998 (O_998,N_29905,N_29874);
nand UO_999 (O_999,N_29829,N_29988);
nor UO_1000 (O_1000,N_29592,N_29113);
nor UO_1001 (O_1001,N_29545,N_29362);
nor UO_1002 (O_1002,N_29244,N_29457);
or UO_1003 (O_1003,N_29083,N_29171);
and UO_1004 (O_1004,N_29908,N_29569);
nor UO_1005 (O_1005,N_29923,N_29595);
nor UO_1006 (O_1006,N_29572,N_29475);
xor UO_1007 (O_1007,N_29710,N_29796);
and UO_1008 (O_1008,N_29053,N_29802);
nand UO_1009 (O_1009,N_29214,N_29051);
nor UO_1010 (O_1010,N_29068,N_29451);
nand UO_1011 (O_1011,N_29739,N_29082);
and UO_1012 (O_1012,N_29650,N_29363);
nand UO_1013 (O_1013,N_29068,N_29095);
nand UO_1014 (O_1014,N_29304,N_29906);
nor UO_1015 (O_1015,N_29228,N_29613);
nor UO_1016 (O_1016,N_29572,N_29232);
and UO_1017 (O_1017,N_29998,N_29704);
xor UO_1018 (O_1018,N_29444,N_29886);
nor UO_1019 (O_1019,N_29926,N_29654);
nand UO_1020 (O_1020,N_29487,N_29542);
xor UO_1021 (O_1021,N_29505,N_29253);
xnor UO_1022 (O_1022,N_29935,N_29507);
and UO_1023 (O_1023,N_29883,N_29247);
xor UO_1024 (O_1024,N_29746,N_29112);
nand UO_1025 (O_1025,N_29200,N_29113);
nand UO_1026 (O_1026,N_29480,N_29826);
nand UO_1027 (O_1027,N_29689,N_29941);
nand UO_1028 (O_1028,N_29987,N_29994);
xor UO_1029 (O_1029,N_29923,N_29635);
xnor UO_1030 (O_1030,N_29986,N_29209);
or UO_1031 (O_1031,N_29232,N_29731);
xor UO_1032 (O_1032,N_29225,N_29685);
xnor UO_1033 (O_1033,N_29714,N_29270);
or UO_1034 (O_1034,N_29240,N_29493);
nor UO_1035 (O_1035,N_29230,N_29307);
nor UO_1036 (O_1036,N_29503,N_29679);
xnor UO_1037 (O_1037,N_29684,N_29090);
nand UO_1038 (O_1038,N_29774,N_29764);
and UO_1039 (O_1039,N_29431,N_29052);
nand UO_1040 (O_1040,N_29016,N_29751);
or UO_1041 (O_1041,N_29930,N_29674);
nor UO_1042 (O_1042,N_29181,N_29274);
and UO_1043 (O_1043,N_29128,N_29500);
or UO_1044 (O_1044,N_29884,N_29943);
xor UO_1045 (O_1045,N_29566,N_29263);
and UO_1046 (O_1046,N_29860,N_29300);
nor UO_1047 (O_1047,N_29069,N_29329);
or UO_1048 (O_1048,N_29424,N_29204);
and UO_1049 (O_1049,N_29693,N_29408);
nor UO_1050 (O_1050,N_29294,N_29206);
nand UO_1051 (O_1051,N_29045,N_29312);
and UO_1052 (O_1052,N_29412,N_29814);
nand UO_1053 (O_1053,N_29468,N_29700);
and UO_1054 (O_1054,N_29735,N_29504);
xor UO_1055 (O_1055,N_29307,N_29171);
nand UO_1056 (O_1056,N_29224,N_29985);
and UO_1057 (O_1057,N_29947,N_29898);
xnor UO_1058 (O_1058,N_29553,N_29045);
and UO_1059 (O_1059,N_29171,N_29286);
or UO_1060 (O_1060,N_29714,N_29191);
or UO_1061 (O_1061,N_29728,N_29628);
nand UO_1062 (O_1062,N_29704,N_29494);
and UO_1063 (O_1063,N_29499,N_29770);
or UO_1064 (O_1064,N_29309,N_29924);
and UO_1065 (O_1065,N_29606,N_29758);
and UO_1066 (O_1066,N_29232,N_29435);
xor UO_1067 (O_1067,N_29431,N_29095);
and UO_1068 (O_1068,N_29510,N_29341);
nor UO_1069 (O_1069,N_29745,N_29672);
or UO_1070 (O_1070,N_29127,N_29927);
xor UO_1071 (O_1071,N_29942,N_29249);
nor UO_1072 (O_1072,N_29951,N_29844);
xor UO_1073 (O_1073,N_29287,N_29242);
or UO_1074 (O_1074,N_29146,N_29759);
nand UO_1075 (O_1075,N_29985,N_29786);
nand UO_1076 (O_1076,N_29298,N_29476);
nand UO_1077 (O_1077,N_29407,N_29623);
nor UO_1078 (O_1078,N_29658,N_29951);
nor UO_1079 (O_1079,N_29249,N_29855);
and UO_1080 (O_1080,N_29482,N_29927);
nor UO_1081 (O_1081,N_29530,N_29934);
nor UO_1082 (O_1082,N_29694,N_29751);
and UO_1083 (O_1083,N_29920,N_29306);
xnor UO_1084 (O_1084,N_29821,N_29193);
and UO_1085 (O_1085,N_29988,N_29630);
or UO_1086 (O_1086,N_29323,N_29125);
nand UO_1087 (O_1087,N_29187,N_29179);
xor UO_1088 (O_1088,N_29143,N_29685);
nor UO_1089 (O_1089,N_29116,N_29075);
nand UO_1090 (O_1090,N_29277,N_29293);
nor UO_1091 (O_1091,N_29895,N_29477);
xnor UO_1092 (O_1092,N_29730,N_29268);
nand UO_1093 (O_1093,N_29491,N_29647);
nand UO_1094 (O_1094,N_29683,N_29117);
xnor UO_1095 (O_1095,N_29850,N_29435);
nor UO_1096 (O_1096,N_29307,N_29347);
nand UO_1097 (O_1097,N_29300,N_29399);
and UO_1098 (O_1098,N_29032,N_29486);
nand UO_1099 (O_1099,N_29567,N_29250);
xnor UO_1100 (O_1100,N_29109,N_29819);
or UO_1101 (O_1101,N_29341,N_29009);
or UO_1102 (O_1102,N_29778,N_29510);
or UO_1103 (O_1103,N_29735,N_29136);
and UO_1104 (O_1104,N_29849,N_29069);
nand UO_1105 (O_1105,N_29128,N_29733);
xnor UO_1106 (O_1106,N_29128,N_29930);
nand UO_1107 (O_1107,N_29939,N_29912);
or UO_1108 (O_1108,N_29850,N_29395);
or UO_1109 (O_1109,N_29500,N_29088);
nor UO_1110 (O_1110,N_29876,N_29344);
and UO_1111 (O_1111,N_29354,N_29467);
nor UO_1112 (O_1112,N_29307,N_29204);
nand UO_1113 (O_1113,N_29692,N_29076);
nor UO_1114 (O_1114,N_29740,N_29918);
nor UO_1115 (O_1115,N_29600,N_29883);
nand UO_1116 (O_1116,N_29124,N_29912);
nor UO_1117 (O_1117,N_29470,N_29965);
and UO_1118 (O_1118,N_29454,N_29947);
or UO_1119 (O_1119,N_29368,N_29475);
xnor UO_1120 (O_1120,N_29618,N_29653);
or UO_1121 (O_1121,N_29950,N_29535);
or UO_1122 (O_1122,N_29038,N_29243);
or UO_1123 (O_1123,N_29157,N_29986);
or UO_1124 (O_1124,N_29112,N_29593);
nor UO_1125 (O_1125,N_29228,N_29709);
nor UO_1126 (O_1126,N_29770,N_29790);
or UO_1127 (O_1127,N_29733,N_29665);
nor UO_1128 (O_1128,N_29563,N_29438);
xor UO_1129 (O_1129,N_29757,N_29014);
xor UO_1130 (O_1130,N_29410,N_29080);
and UO_1131 (O_1131,N_29448,N_29434);
xor UO_1132 (O_1132,N_29331,N_29178);
nand UO_1133 (O_1133,N_29987,N_29261);
nand UO_1134 (O_1134,N_29598,N_29093);
or UO_1135 (O_1135,N_29284,N_29306);
nor UO_1136 (O_1136,N_29974,N_29938);
xnor UO_1137 (O_1137,N_29219,N_29453);
or UO_1138 (O_1138,N_29398,N_29588);
xnor UO_1139 (O_1139,N_29275,N_29532);
nor UO_1140 (O_1140,N_29555,N_29429);
or UO_1141 (O_1141,N_29482,N_29999);
nor UO_1142 (O_1142,N_29725,N_29757);
nor UO_1143 (O_1143,N_29204,N_29732);
nand UO_1144 (O_1144,N_29472,N_29802);
nand UO_1145 (O_1145,N_29963,N_29931);
and UO_1146 (O_1146,N_29561,N_29555);
or UO_1147 (O_1147,N_29268,N_29539);
xnor UO_1148 (O_1148,N_29026,N_29956);
or UO_1149 (O_1149,N_29991,N_29839);
or UO_1150 (O_1150,N_29567,N_29547);
or UO_1151 (O_1151,N_29820,N_29691);
xor UO_1152 (O_1152,N_29874,N_29152);
nand UO_1153 (O_1153,N_29183,N_29751);
or UO_1154 (O_1154,N_29992,N_29608);
xor UO_1155 (O_1155,N_29529,N_29714);
and UO_1156 (O_1156,N_29132,N_29229);
or UO_1157 (O_1157,N_29216,N_29540);
nor UO_1158 (O_1158,N_29797,N_29825);
nand UO_1159 (O_1159,N_29398,N_29165);
and UO_1160 (O_1160,N_29113,N_29460);
xor UO_1161 (O_1161,N_29457,N_29579);
xor UO_1162 (O_1162,N_29000,N_29408);
nor UO_1163 (O_1163,N_29688,N_29304);
nand UO_1164 (O_1164,N_29675,N_29516);
and UO_1165 (O_1165,N_29181,N_29535);
and UO_1166 (O_1166,N_29609,N_29588);
and UO_1167 (O_1167,N_29391,N_29221);
nand UO_1168 (O_1168,N_29746,N_29854);
xor UO_1169 (O_1169,N_29281,N_29325);
xor UO_1170 (O_1170,N_29365,N_29379);
nand UO_1171 (O_1171,N_29332,N_29135);
or UO_1172 (O_1172,N_29340,N_29714);
nor UO_1173 (O_1173,N_29241,N_29628);
nor UO_1174 (O_1174,N_29720,N_29593);
nand UO_1175 (O_1175,N_29532,N_29427);
and UO_1176 (O_1176,N_29718,N_29404);
or UO_1177 (O_1177,N_29498,N_29552);
and UO_1178 (O_1178,N_29547,N_29185);
nand UO_1179 (O_1179,N_29720,N_29377);
nor UO_1180 (O_1180,N_29446,N_29678);
nand UO_1181 (O_1181,N_29851,N_29987);
xnor UO_1182 (O_1182,N_29496,N_29343);
and UO_1183 (O_1183,N_29533,N_29106);
nor UO_1184 (O_1184,N_29086,N_29431);
or UO_1185 (O_1185,N_29448,N_29508);
and UO_1186 (O_1186,N_29196,N_29501);
or UO_1187 (O_1187,N_29820,N_29591);
xnor UO_1188 (O_1188,N_29487,N_29626);
nor UO_1189 (O_1189,N_29785,N_29617);
or UO_1190 (O_1190,N_29703,N_29591);
nand UO_1191 (O_1191,N_29973,N_29621);
nand UO_1192 (O_1192,N_29957,N_29288);
xnor UO_1193 (O_1193,N_29786,N_29040);
xor UO_1194 (O_1194,N_29074,N_29996);
nor UO_1195 (O_1195,N_29618,N_29069);
nor UO_1196 (O_1196,N_29117,N_29848);
nand UO_1197 (O_1197,N_29771,N_29025);
nor UO_1198 (O_1198,N_29619,N_29228);
nor UO_1199 (O_1199,N_29607,N_29671);
nand UO_1200 (O_1200,N_29963,N_29462);
xor UO_1201 (O_1201,N_29009,N_29147);
nor UO_1202 (O_1202,N_29392,N_29280);
and UO_1203 (O_1203,N_29888,N_29570);
nand UO_1204 (O_1204,N_29723,N_29051);
nor UO_1205 (O_1205,N_29702,N_29672);
xnor UO_1206 (O_1206,N_29316,N_29941);
nor UO_1207 (O_1207,N_29788,N_29723);
and UO_1208 (O_1208,N_29746,N_29971);
xnor UO_1209 (O_1209,N_29771,N_29353);
xor UO_1210 (O_1210,N_29329,N_29365);
nand UO_1211 (O_1211,N_29047,N_29273);
or UO_1212 (O_1212,N_29969,N_29115);
and UO_1213 (O_1213,N_29012,N_29890);
nand UO_1214 (O_1214,N_29011,N_29463);
nand UO_1215 (O_1215,N_29386,N_29733);
or UO_1216 (O_1216,N_29882,N_29215);
nand UO_1217 (O_1217,N_29773,N_29844);
nor UO_1218 (O_1218,N_29722,N_29154);
or UO_1219 (O_1219,N_29759,N_29779);
and UO_1220 (O_1220,N_29748,N_29635);
nor UO_1221 (O_1221,N_29983,N_29596);
nand UO_1222 (O_1222,N_29017,N_29027);
or UO_1223 (O_1223,N_29180,N_29458);
xnor UO_1224 (O_1224,N_29463,N_29949);
xor UO_1225 (O_1225,N_29491,N_29757);
nor UO_1226 (O_1226,N_29529,N_29390);
xnor UO_1227 (O_1227,N_29119,N_29957);
nand UO_1228 (O_1228,N_29921,N_29831);
nand UO_1229 (O_1229,N_29118,N_29741);
or UO_1230 (O_1230,N_29042,N_29499);
nand UO_1231 (O_1231,N_29430,N_29312);
nand UO_1232 (O_1232,N_29245,N_29829);
and UO_1233 (O_1233,N_29115,N_29138);
xnor UO_1234 (O_1234,N_29420,N_29354);
or UO_1235 (O_1235,N_29941,N_29738);
xnor UO_1236 (O_1236,N_29933,N_29659);
or UO_1237 (O_1237,N_29119,N_29088);
nand UO_1238 (O_1238,N_29370,N_29443);
or UO_1239 (O_1239,N_29889,N_29525);
nor UO_1240 (O_1240,N_29757,N_29423);
nor UO_1241 (O_1241,N_29691,N_29701);
or UO_1242 (O_1242,N_29476,N_29255);
or UO_1243 (O_1243,N_29592,N_29765);
xor UO_1244 (O_1244,N_29971,N_29539);
xnor UO_1245 (O_1245,N_29139,N_29394);
and UO_1246 (O_1246,N_29013,N_29341);
and UO_1247 (O_1247,N_29985,N_29642);
or UO_1248 (O_1248,N_29499,N_29555);
nor UO_1249 (O_1249,N_29035,N_29106);
xor UO_1250 (O_1250,N_29585,N_29650);
nor UO_1251 (O_1251,N_29884,N_29912);
and UO_1252 (O_1252,N_29820,N_29461);
or UO_1253 (O_1253,N_29745,N_29008);
or UO_1254 (O_1254,N_29032,N_29451);
nand UO_1255 (O_1255,N_29868,N_29728);
nor UO_1256 (O_1256,N_29453,N_29568);
or UO_1257 (O_1257,N_29202,N_29960);
nand UO_1258 (O_1258,N_29976,N_29516);
xor UO_1259 (O_1259,N_29817,N_29483);
xnor UO_1260 (O_1260,N_29664,N_29219);
or UO_1261 (O_1261,N_29673,N_29580);
nand UO_1262 (O_1262,N_29129,N_29803);
and UO_1263 (O_1263,N_29724,N_29925);
nor UO_1264 (O_1264,N_29724,N_29324);
xnor UO_1265 (O_1265,N_29614,N_29086);
and UO_1266 (O_1266,N_29250,N_29454);
xor UO_1267 (O_1267,N_29995,N_29105);
xnor UO_1268 (O_1268,N_29237,N_29044);
nor UO_1269 (O_1269,N_29801,N_29031);
xnor UO_1270 (O_1270,N_29017,N_29422);
nand UO_1271 (O_1271,N_29187,N_29131);
xnor UO_1272 (O_1272,N_29010,N_29355);
nor UO_1273 (O_1273,N_29008,N_29467);
nor UO_1274 (O_1274,N_29349,N_29306);
and UO_1275 (O_1275,N_29177,N_29584);
nand UO_1276 (O_1276,N_29330,N_29340);
xor UO_1277 (O_1277,N_29630,N_29640);
xnor UO_1278 (O_1278,N_29099,N_29783);
xor UO_1279 (O_1279,N_29453,N_29753);
nor UO_1280 (O_1280,N_29442,N_29406);
and UO_1281 (O_1281,N_29408,N_29496);
nor UO_1282 (O_1282,N_29661,N_29809);
or UO_1283 (O_1283,N_29792,N_29082);
nor UO_1284 (O_1284,N_29809,N_29330);
nor UO_1285 (O_1285,N_29363,N_29049);
and UO_1286 (O_1286,N_29336,N_29550);
and UO_1287 (O_1287,N_29929,N_29758);
xor UO_1288 (O_1288,N_29075,N_29850);
or UO_1289 (O_1289,N_29462,N_29619);
nand UO_1290 (O_1290,N_29774,N_29707);
and UO_1291 (O_1291,N_29496,N_29707);
nor UO_1292 (O_1292,N_29647,N_29898);
xor UO_1293 (O_1293,N_29276,N_29256);
xor UO_1294 (O_1294,N_29033,N_29517);
xnor UO_1295 (O_1295,N_29293,N_29885);
nand UO_1296 (O_1296,N_29280,N_29984);
or UO_1297 (O_1297,N_29328,N_29571);
nand UO_1298 (O_1298,N_29733,N_29700);
xor UO_1299 (O_1299,N_29313,N_29383);
or UO_1300 (O_1300,N_29506,N_29163);
nand UO_1301 (O_1301,N_29521,N_29687);
xnor UO_1302 (O_1302,N_29752,N_29267);
and UO_1303 (O_1303,N_29608,N_29383);
or UO_1304 (O_1304,N_29118,N_29128);
nand UO_1305 (O_1305,N_29358,N_29008);
or UO_1306 (O_1306,N_29407,N_29516);
xnor UO_1307 (O_1307,N_29828,N_29702);
or UO_1308 (O_1308,N_29525,N_29812);
nor UO_1309 (O_1309,N_29076,N_29991);
xor UO_1310 (O_1310,N_29208,N_29690);
and UO_1311 (O_1311,N_29394,N_29876);
and UO_1312 (O_1312,N_29333,N_29313);
nor UO_1313 (O_1313,N_29983,N_29967);
nor UO_1314 (O_1314,N_29298,N_29273);
or UO_1315 (O_1315,N_29504,N_29099);
nor UO_1316 (O_1316,N_29885,N_29184);
or UO_1317 (O_1317,N_29056,N_29910);
nand UO_1318 (O_1318,N_29099,N_29345);
nor UO_1319 (O_1319,N_29506,N_29973);
nor UO_1320 (O_1320,N_29456,N_29880);
xor UO_1321 (O_1321,N_29150,N_29845);
xor UO_1322 (O_1322,N_29539,N_29063);
or UO_1323 (O_1323,N_29878,N_29954);
nand UO_1324 (O_1324,N_29940,N_29935);
xnor UO_1325 (O_1325,N_29188,N_29691);
xnor UO_1326 (O_1326,N_29985,N_29495);
and UO_1327 (O_1327,N_29279,N_29300);
or UO_1328 (O_1328,N_29011,N_29777);
xnor UO_1329 (O_1329,N_29696,N_29674);
nor UO_1330 (O_1330,N_29226,N_29022);
nand UO_1331 (O_1331,N_29295,N_29080);
xnor UO_1332 (O_1332,N_29890,N_29263);
xnor UO_1333 (O_1333,N_29789,N_29231);
or UO_1334 (O_1334,N_29052,N_29251);
or UO_1335 (O_1335,N_29456,N_29996);
nor UO_1336 (O_1336,N_29523,N_29695);
or UO_1337 (O_1337,N_29626,N_29414);
xnor UO_1338 (O_1338,N_29040,N_29578);
nand UO_1339 (O_1339,N_29972,N_29608);
xor UO_1340 (O_1340,N_29773,N_29252);
or UO_1341 (O_1341,N_29757,N_29857);
or UO_1342 (O_1342,N_29410,N_29088);
nor UO_1343 (O_1343,N_29251,N_29733);
or UO_1344 (O_1344,N_29288,N_29355);
nand UO_1345 (O_1345,N_29333,N_29351);
and UO_1346 (O_1346,N_29412,N_29954);
xor UO_1347 (O_1347,N_29789,N_29311);
xnor UO_1348 (O_1348,N_29893,N_29308);
nor UO_1349 (O_1349,N_29222,N_29372);
or UO_1350 (O_1350,N_29269,N_29825);
xor UO_1351 (O_1351,N_29328,N_29128);
nor UO_1352 (O_1352,N_29046,N_29928);
nor UO_1353 (O_1353,N_29937,N_29437);
nand UO_1354 (O_1354,N_29950,N_29851);
and UO_1355 (O_1355,N_29478,N_29367);
nand UO_1356 (O_1356,N_29697,N_29244);
and UO_1357 (O_1357,N_29527,N_29510);
nor UO_1358 (O_1358,N_29127,N_29134);
nor UO_1359 (O_1359,N_29247,N_29712);
or UO_1360 (O_1360,N_29143,N_29677);
and UO_1361 (O_1361,N_29969,N_29290);
xnor UO_1362 (O_1362,N_29047,N_29415);
and UO_1363 (O_1363,N_29738,N_29164);
and UO_1364 (O_1364,N_29857,N_29393);
or UO_1365 (O_1365,N_29239,N_29405);
nand UO_1366 (O_1366,N_29570,N_29342);
nor UO_1367 (O_1367,N_29820,N_29001);
xor UO_1368 (O_1368,N_29870,N_29276);
or UO_1369 (O_1369,N_29612,N_29163);
and UO_1370 (O_1370,N_29963,N_29845);
xnor UO_1371 (O_1371,N_29504,N_29012);
nand UO_1372 (O_1372,N_29230,N_29725);
xor UO_1373 (O_1373,N_29842,N_29599);
or UO_1374 (O_1374,N_29179,N_29104);
nand UO_1375 (O_1375,N_29130,N_29139);
and UO_1376 (O_1376,N_29022,N_29380);
or UO_1377 (O_1377,N_29181,N_29294);
nor UO_1378 (O_1378,N_29116,N_29822);
or UO_1379 (O_1379,N_29273,N_29116);
and UO_1380 (O_1380,N_29291,N_29994);
nand UO_1381 (O_1381,N_29331,N_29228);
xnor UO_1382 (O_1382,N_29249,N_29481);
xor UO_1383 (O_1383,N_29501,N_29664);
xor UO_1384 (O_1384,N_29611,N_29208);
nor UO_1385 (O_1385,N_29759,N_29383);
xor UO_1386 (O_1386,N_29743,N_29871);
xnor UO_1387 (O_1387,N_29967,N_29090);
xor UO_1388 (O_1388,N_29988,N_29845);
or UO_1389 (O_1389,N_29158,N_29786);
nor UO_1390 (O_1390,N_29543,N_29384);
or UO_1391 (O_1391,N_29046,N_29347);
and UO_1392 (O_1392,N_29369,N_29886);
and UO_1393 (O_1393,N_29364,N_29940);
or UO_1394 (O_1394,N_29137,N_29850);
and UO_1395 (O_1395,N_29331,N_29572);
xor UO_1396 (O_1396,N_29166,N_29421);
and UO_1397 (O_1397,N_29994,N_29648);
nand UO_1398 (O_1398,N_29355,N_29551);
nor UO_1399 (O_1399,N_29195,N_29474);
or UO_1400 (O_1400,N_29419,N_29786);
or UO_1401 (O_1401,N_29326,N_29759);
nor UO_1402 (O_1402,N_29129,N_29276);
nor UO_1403 (O_1403,N_29051,N_29467);
nand UO_1404 (O_1404,N_29976,N_29191);
or UO_1405 (O_1405,N_29593,N_29363);
nor UO_1406 (O_1406,N_29900,N_29591);
nand UO_1407 (O_1407,N_29987,N_29170);
nor UO_1408 (O_1408,N_29884,N_29115);
nand UO_1409 (O_1409,N_29793,N_29542);
nor UO_1410 (O_1410,N_29122,N_29987);
and UO_1411 (O_1411,N_29685,N_29647);
nand UO_1412 (O_1412,N_29869,N_29188);
nand UO_1413 (O_1413,N_29375,N_29007);
and UO_1414 (O_1414,N_29032,N_29640);
and UO_1415 (O_1415,N_29963,N_29623);
xor UO_1416 (O_1416,N_29151,N_29870);
xnor UO_1417 (O_1417,N_29119,N_29844);
or UO_1418 (O_1418,N_29118,N_29213);
xnor UO_1419 (O_1419,N_29298,N_29723);
xnor UO_1420 (O_1420,N_29817,N_29330);
and UO_1421 (O_1421,N_29920,N_29051);
nand UO_1422 (O_1422,N_29818,N_29993);
and UO_1423 (O_1423,N_29304,N_29853);
and UO_1424 (O_1424,N_29915,N_29152);
nor UO_1425 (O_1425,N_29476,N_29354);
nand UO_1426 (O_1426,N_29494,N_29214);
nor UO_1427 (O_1427,N_29173,N_29840);
or UO_1428 (O_1428,N_29360,N_29655);
xor UO_1429 (O_1429,N_29696,N_29285);
and UO_1430 (O_1430,N_29642,N_29391);
or UO_1431 (O_1431,N_29798,N_29001);
and UO_1432 (O_1432,N_29106,N_29316);
nor UO_1433 (O_1433,N_29975,N_29529);
nand UO_1434 (O_1434,N_29976,N_29821);
or UO_1435 (O_1435,N_29323,N_29765);
or UO_1436 (O_1436,N_29638,N_29953);
nor UO_1437 (O_1437,N_29726,N_29772);
nor UO_1438 (O_1438,N_29083,N_29907);
or UO_1439 (O_1439,N_29056,N_29642);
or UO_1440 (O_1440,N_29132,N_29127);
xnor UO_1441 (O_1441,N_29605,N_29621);
and UO_1442 (O_1442,N_29886,N_29553);
and UO_1443 (O_1443,N_29236,N_29842);
xor UO_1444 (O_1444,N_29936,N_29778);
nor UO_1445 (O_1445,N_29926,N_29713);
or UO_1446 (O_1446,N_29000,N_29579);
xnor UO_1447 (O_1447,N_29516,N_29841);
xnor UO_1448 (O_1448,N_29314,N_29802);
xor UO_1449 (O_1449,N_29936,N_29791);
xnor UO_1450 (O_1450,N_29915,N_29960);
nor UO_1451 (O_1451,N_29155,N_29487);
and UO_1452 (O_1452,N_29617,N_29339);
and UO_1453 (O_1453,N_29540,N_29229);
xor UO_1454 (O_1454,N_29608,N_29124);
nor UO_1455 (O_1455,N_29450,N_29692);
xnor UO_1456 (O_1456,N_29899,N_29519);
xor UO_1457 (O_1457,N_29854,N_29985);
nor UO_1458 (O_1458,N_29171,N_29641);
nor UO_1459 (O_1459,N_29602,N_29869);
or UO_1460 (O_1460,N_29312,N_29685);
or UO_1461 (O_1461,N_29888,N_29318);
or UO_1462 (O_1462,N_29013,N_29200);
or UO_1463 (O_1463,N_29365,N_29209);
nand UO_1464 (O_1464,N_29192,N_29017);
and UO_1465 (O_1465,N_29817,N_29717);
nor UO_1466 (O_1466,N_29409,N_29244);
or UO_1467 (O_1467,N_29396,N_29652);
nand UO_1468 (O_1468,N_29941,N_29831);
nor UO_1469 (O_1469,N_29965,N_29932);
and UO_1470 (O_1470,N_29163,N_29181);
xor UO_1471 (O_1471,N_29955,N_29470);
nor UO_1472 (O_1472,N_29650,N_29060);
nor UO_1473 (O_1473,N_29020,N_29879);
nor UO_1474 (O_1474,N_29563,N_29847);
xnor UO_1475 (O_1475,N_29310,N_29388);
and UO_1476 (O_1476,N_29968,N_29134);
xnor UO_1477 (O_1477,N_29213,N_29881);
nand UO_1478 (O_1478,N_29873,N_29458);
or UO_1479 (O_1479,N_29120,N_29331);
nand UO_1480 (O_1480,N_29758,N_29656);
nand UO_1481 (O_1481,N_29912,N_29610);
xnor UO_1482 (O_1482,N_29932,N_29373);
and UO_1483 (O_1483,N_29790,N_29167);
and UO_1484 (O_1484,N_29153,N_29870);
nor UO_1485 (O_1485,N_29343,N_29193);
xnor UO_1486 (O_1486,N_29230,N_29541);
or UO_1487 (O_1487,N_29034,N_29884);
nand UO_1488 (O_1488,N_29793,N_29340);
nand UO_1489 (O_1489,N_29764,N_29944);
and UO_1490 (O_1490,N_29484,N_29307);
nor UO_1491 (O_1491,N_29395,N_29018);
nor UO_1492 (O_1492,N_29166,N_29499);
and UO_1493 (O_1493,N_29013,N_29231);
or UO_1494 (O_1494,N_29533,N_29048);
xor UO_1495 (O_1495,N_29609,N_29864);
and UO_1496 (O_1496,N_29058,N_29925);
nor UO_1497 (O_1497,N_29257,N_29328);
and UO_1498 (O_1498,N_29794,N_29323);
and UO_1499 (O_1499,N_29119,N_29164);
nor UO_1500 (O_1500,N_29650,N_29471);
xnor UO_1501 (O_1501,N_29429,N_29948);
nand UO_1502 (O_1502,N_29064,N_29740);
nor UO_1503 (O_1503,N_29280,N_29303);
nand UO_1504 (O_1504,N_29170,N_29576);
nand UO_1505 (O_1505,N_29604,N_29151);
nand UO_1506 (O_1506,N_29907,N_29723);
nand UO_1507 (O_1507,N_29698,N_29675);
nand UO_1508 (O_1508,N_29898,N_29102);
xnor UO_1509 (O_1509,N_29063,N_29005);
nand UO_1510 (O_1510,N_29306,N_29106);
or UO_1511 (O_1511,N_29134,N_29882);
nor UO_1512 (O_1512,N_29587,N_29581);
xor UO_1513 (O_1513,N_29060,N_29721);
or UO_1514 (O_1514,N_29051,N_29096);
and UO_1515 (O_1515,N_29266,N_29763);
and UO_1516 (O_1516,N_29173,N_29070);
nand UO_1517 (O_1517,N_29920,N_29731);
nand UO_1518 (O_1518,N_29957,N_29032);
xnor UO_1519 (O_1519,N_29900,N_29626);
or UO_1520 (O_1520,N_29181,N_29775);
or UO_1521 (O_1521,N_29113,N_29611);
and UO_1522 (O_1522,N_29073,N_29997);
and UO_1523 (O_1523,N_29323,N_29573);
and UO_1524 (O_1524,N_29198,N_29221);
and UO_1525 (O_1525,N_29183,N_29740);
and UO_1526 (O_1526,N_29659,N_29259);
or UO_1527 (O_1527,N_29720,N_29429);
nor UO_1528 (O_1528,N_29581,N_29521);
and UO_1529 (O_1529,N_29544,N_29612);
xor UO_1530 (O_1530,N_29389,N_29821);
xnor UO_1531 (O_1531,N_29272,N_29421);
xnor UO_1532 (O_1532,N_29620,N_29094);
xnor UO_1533 (O_1533,N_29749,N_29306);
or UO_1534 (O_1534,N_29553,N_29491);
and UO_1535 (O_1535,N_29965,N_29750);
xor UO_1536 (O_1536,N_29419,N_29058);
or UO_1537 (O_1537,N_29967,N_29667);
nor UO_1538 (O_1538,N_29651,N_29094);
or UO_1539 (O_1539,N_29937,N_29163);
and UO_1540 (O_1540,N_29896,N_29837);
or UO_1541 (O_1541,N_29853,N_29768);
and UO_1542 (O_1542,N_29723,N_29598);
nor UO_1543 (O_1543,N_29148,N_29285);
and UO_1544 (O_1544,N_29612,N_29703);
and UO_1545 (O_1545,N_29163,N_29019);
nand UO_1546 (O_1546,N_29641,N_29602);
nand UO_1547 (O_1547,N_29821,N_29147);
or UO_1548 (O_1548,N_29283,N_29225);
and UO_1549 (O_1549,N_29188,N_29920);
nand UO_1550 (O_1550,N_29552,N_29590);
xor UO_1551 (O_1551,N_29808,N_29562);
xnor UO_1552 (O_1552,N_29039,N_29701);
nor UO_1553 (O_1553,N_29691,N_29971);
nor UO_1554 (O_1554,N_29098,N_29908);
xor UO_1555 (O_1555,N_29935,N_29354);
nand UO_1556 (O_1556,N_29169,N_29011);
nor UO_1557 (O_1557,N_29999,N_29362);
nand UO_1558 (O_1558,N_29054,N_29793);
xnor UO_1559 (O_1559,N_29444,N_29376);
and UO_1560 (O_1560,N_29423,N_29043);
and UO_1561 (O_1561,N_29899,N_29425);
xnor UO_1562 (O_1562,N_29416,N_29850);
xor UO_1563 (O_1563,N_29197,N_29139);
and UO_1564 (O_1564,N_29834,N_29195);
and UO_1565 (O_1565,N_29571,N_29094);
or UO_1566 (O_1566,N_29147,N_29804);
and UO_1567 (O_1567,N_29114,N_29267);
or UO_1568 (O_1568,N_29343,N_29149);
nand UO_1569 (O_1569,N_29891,N_29535);
nand UO_1570 (O_1570,N_29550,N_29569);
xnor UO_1571 (O_1571,N_29831,N_29610);
nand UO_1572 (O_1572,N_29448,N_29909);
nand UO_1573 (O_1573,N_29990,N_29666);
xnor UO_1574 (O_1574,N_29036,N_29390);
nand UO_1575 (O_1575,N_29301,N_29230);
nor UO_1576 (O_1576,N_29073,N_29249);
nand UO_1577 (O_1577,N_29044,N_29208);
nor UO_1578 (O_1578,N_29989,N_29214);
and UO_1579 (O_1579,N_29595,N_29887);
nor UO_1580 (O_1580,N_29405,N_29992);
and UO_1581 (O_1581,N_29929,N_29006);
or UO_1582 (O_1582,N_29613,N_29356);
nor UO_1583 (O_1583,N_29612,N_29312);
nor UO_1584 (O_1584,N_29094,N_29205);
nand UO_1585 (O_1585,N_29458,N_29908);
xnor UO_1586 (O_1586,N_29089,N_29945);
xor UO_1587 (O_1587,N_29161,N_29344);
or UO_1588 (O_1588,N_29305,N_29958);
nand UO_1589 (O_1589,N_29333,N_29603);
or UO_1590 (O_1590,N_29006,N_29721);
nor UO_1591 (O_1591,N_29386,N_29281);
and UO_1592 (O_1592,N_29975,N_29584);
xor UO_1593 (O_1593,N_29037,N_29768);
xnor UO_1594 (O_1594,N_29219,N_29354);
and UO_1595 (O_1595,N_29397,N_29219);
or UO_1596 (O_1596,N_29702,N_29847);
nor UO_1597 (O_1597,N_29364,N_29454);
xnor UO_1598 (O_1598,N_29439,N_29681);
and UO_1599 (O_1599,N_29103,N_29232);
and UO_1600 (O_1600,N_29264,N_29663);
and UO_1601 (O_1601,N_29534,N_29442);
and UO_1602 (O_1602,N_29314,N_29256);
nand UO_1603 (O_1603,N_29046,N_29002);
nand UO_1604 (O_1604,N_29316,N_29267);
xnor UO_1605 (O_1605,N_29381,N_29136);
nor UO_1606 (O_1606,N_29308,N_29036);
or UO_1607 (O_1607,N_29174,N_29202);
xnor UO_1608 (O_1608,N_29484,N_29509);
nor UO_1609 (O_1609,N_29091,N_29881);
and UO_1610 (O_1610,N_29181,N_29135);
or UO_1611 (O_1611,N_29904,N_29082);
or UO_1612 (O_1612,N_29355,N_29661);
or UO_1613 (O_1613,N_29036,N_29516);
and UO_1614 (O_1614,N_29707,N_29019);
xnor UO_1615 (O_1615,N_29078,N_29558);
nor UO_1616 (O_1616,N_29088,N_29577);
nor UO_1617 (O_1617,N_29802,N_29724);
and UO_1618 (O_1618,N_29888,N_29330);
and UO_1619 (O_1619,N_29381,N_29495);
nand UO_1620 (O_1620,N_29537,N_29698);
nand UO_1621 (O_1621,N_29378,N_29792);
nand UO_1622 (O_1622,N_29269,N_29866);
nor UO_1623 (O_1623,N_29653,N_29940);
or UO_1624 (O_1624,N_29419,N_29564);
or UO_1625 (O_1625,N_29165,N_29341);
xnor UO_1626 (O_1626,N_29410,N_29816);
xor UO_1627 (O_1627,N_29582,N_29361);
and UO_1628 (O_1628,N_29017,N_29426);
or UO_1629 (O_1629,N_29553,N_29463);
nor UO_1630 (O_1630,N_29154,N_29586);
nor UO_1631 (O_1631,N_29339,N_29325);
xnor UO_1632 (O_1632,N_29282,N_29345);
nor UO_1633 (O_1633,N_29161,N_29059);
and UO_1634 (O_1634,N_29546,N_29833);
nand UO_1635 (O_1635,N_29369,N_29177);
and UO_1636 (O_1636,N_29684,N_29740);
nand UO_1637 (O_1637,N_29838,N_29778);
or UO_1638 (O_1638,N_29781,N_29473);
xor UO_1639 (O_1639,N_29600,N_29213);
xnor UO_1640 (O_1640,N_29075,N_29498);
nand UO_1641 (O_1641,N_29901,N_29383);
nand UO_1642 (O_1642,N_29587,N_29862);
and UO_1643 (O_1643,N_29663,N_29140);
and UO_1644 (O_1644,N_29731,N_29553);
nand UO_1645 (O_1645,N_29373,N_29683);
and UO_1646 (O_1646,N_29860,N_29405);
xor UO_1647 (O_1647,N_29982,N_29388);
nor UO_1648 (O_1648,N_29903,N_29887);
nor UO_1649 (O_1649,N_29447,N_29532);
nor UO_1650 (O_1650,N_29164,N_29797);
and UO_1651 (O_1651,N_29887,N_29498);
nor UO_1652 (O_1652,N_29072,N_29927);
nor UO_1653 (O_1653,N_29113,N_29248);
nand UO_1654 (O_1654,N_29663,N_29555);
nor UO_1655 (O_1655,N_29094,N_29199);
nand UO_1656 (O_1656,N_29678,N_29493);
and UO_1657 (O_1657,N_29432,N_29884);
xnor UO_1658 (O_1658,N_29186,N_29151);
or UO_1659 (O_1659,N_29075,N_29960);
nor UO_1660 (O_1660,N_29168,N_29038);
and UO_1661 (O_1661,N_29961,N_29988);
xnor UO_1662 (O_1662,N_29600,N_29625);
or UO_1663 (O_1663,N_29462,N_29463);
nor UO_1664 (O_1664,N_29298,N_29724);
nor UO_1665 (O_1665,N_29454,N_29400);
nand UO_1666 (O_1666,N_29092,N_29479);
and UO_1667 (O_1667,N_29658,N_29134);
nand UO_1668 (O_1668,N_29382,N_29251);
xnor UO_1669 (O_1669,N_29957,N_29858);
xor UO_1670 (O_1670,N_29997,N_29704);
nand UO_1671 (O_1671,N_29223,N_29379);
and UO_1672 (O_1672,N_29500,N_29762);
nor UO_1673 (O_1673,N_29929,N_29036);
nor UO_1674 (O_1674,N_29065,N_29768);
xnor UO_1675 (O_1675,N_29983,N_29224);
nor UO_1676 (O_1676,N_29901,N_29118);
or UO_1677 (O_1677,N_29385,N_29785);
xor UO_1678 (O_1678,N_29903,N_29318);
and UO_1679 (O_1679,N_29979,N_29956);
nor UO_1680 (O_1680,N_29248,N_29110);
or UO_1681 (O_1681,N_29788,N_29239);
or UO_1682 (O_1682,N_29661,N_29027);
or UO_1683 (O_1683,N_29550,N_29970);
and UO_1684 (O_1684,N_29328,N_29053);
nor UO_1685 (O_1685,N_29693,N_29239);
xnor UO_1686 (O_1686,N_29348,N_29447);
or UO_1687 (O_1687,N_29047,N_29018);
and UO_1688 (O_1688,N_29640,N_29872);
xor UO_1689 (O_1689,N_29638,N_29875);
and UO_1690 (O_1690,N_29072,N_29656);
and UO_1691 (O_1691,N_29917,N_29512);
and UO_1692 (O_1692,N_29698,N_29322);
nor UO_1693 (O_1693,N_29555,N_29924);
or UO_1694 (O_1694,N_29741,N_29906);
and UO_1695 (O_1695,N_29746,N_29190);
xnor UO_1696 (O_1696,N_29595,N_29669);
nor UO_1697 (O_1697,N_29532,N_29503);
nor UO_1698 (O_1698,N_29044,N_29643);
nor UO_1699 (O_1699,N_29901,N_29599);
or UO_1700 (O_1700,N_29606,N_29903);
or UO_1701 (O_1701,N_29409,N_29969);
nand UO_1702 (O_1702,N_29559,N_29608);
and UO_1703 (O_1703,N_29208,N_29583);
or UO_1704 (O_1704,N_29689,N_29614);
nor UO_1705 (O_1705,N_29488,N_29714);
nor UO_1706 (O_1706,N_29932,N_29463);
nand UO_1707 (O_1707,N_29682,N_29220);
xor UO_1708 (O_1708,N_29321,N_29403);
or UO_1709 (O_1709,N_29212,N_29114);
xor UO_1710 (O_1710,N_29509,N_29708);
and UO_1711 (O_1711,N_29995,N_29206);
nand UO_1712 (O_1712,N_29696,N_29926);
nand UO_1713 (O_1713,N_29180,N_29578);
nand UO_1714 (O_1714,N_29984,N_29520);
or UO_1715 (O_1715,N_29898,N_29879);
and UO_1716 (O_1716,N_29429,N_29325);
xor UO_1717 (O_1717,N_29986,N_29381);
and UO_1718 (O_1718,N_29283,N_29959);
and UO_1719 (O_1719,N_29562,N_29723);
nand UO_1720 (O_1720,N_29780,N_29191);
nand UO_1721 (O_1721,N_29245,N_29871);
xor UO_1722 (O_1722,N_29209,N_29644);
xor UO_1723 (O_1723,N_29986,N_29369);
nor UO_1724 (O_1724,N_29660,N_29473);
and UO_1725 (O_1725,N_29788,N_29369);
nand UO_1726 (O_1726,N_29080,N_29743);
nand UO_1727 (O_1727,N_29457,N_29601);
nand UO_1728 (O_1728,N_29832,N_29897);
and UO_1729 (O_1729,N_29581,N_29841);
or UO_1730 (O_1730,N_29729,N_29022);
and UO_1731 (O_1731,N_29200,N_29250);
nor UO_1732 (O_1732,N_29663,N_29722);
or UO_1733 (O_1733,N_29998,N_29286);
and UO_1734 (O_1734,N_29694,N_29462);
or UO_1735 (O_1735,N_29425,N_29122);
xor UO_1736 (O_1736,N_29792,N_29717);
and UO_1737 (O_1737,N_29141,N_29856);
and UO_1738 (O_1738,N_29224,N_29337);
nand UO_1739 (O_1739,N_29242,N_29948);
xor UO_1740 (O_1740,N_29216,N_29127);
xor UO_1741 (O_1741,N_29651,N_29882);
xor UO_1742 (O_1742,N_29045,N_29967);
and UO_1743 (O_1743,N_29837,N_29212);
nand UO_1744 (O_1744,N_29703,N_29829);
nand UO_1745 (O_1745,N_29421,N_29802);
nor UO_1746 (O_1746,N_29348,N_29064);
and UO_1747 (O_1747,N_29657,N_29972);
or UO_1748 (O_1748,N_29715,N_29730);
and UO_1749 (O_1749,N_29251,N_29998);
and UO_1750 (O_1750,N_29244,N_29930);
nand UO_1751 (O_1751,N_29178,N_29693);
or UO_1752 (O_1752,N_29446,N_29695);
nand UO_1753 (O_1753,N_29304,N_29681);
xnor UO_1754 (O_1754,N_29892,N_29074);
or UO_1755 (O_1755,N_29657,N_29937);
and UO_1756 (O_1756,N_29854,N_29315);
nor UO_1757 (O_1757,N_29983,N_29786);
nand UO_1758 (O_1758,N_29124,N_29074);
or UO_1759 (O_1759,N_29427,N_29898);
nand UO_1760 (O_1760,N_29494,N_29678);
nand UO_1761 (O_1761,N_29450,N_29820);
nor UO_1762 (O_1762,N_29462,N_29504);
xnor UO_1763 (O_1763,N_29421,N_29746);
nor UO_1764 (O_1764,N_29596,N_29195);
and UO_1765 (O_1765,N_29362,N_29749);
nor UO_1766 (O_1766,N_29238,N_29989);
or UO_1767 (O_1767,N_29405,N_29947);
and UO_1768 (O_1768,N_29138,N_29958);
nand UO_1769 (O_1769,N_29816,N_29139);
xor UO_1770 (O_1770,N_29703,N_29592);
nor UO_1771 (O_1771,N_29570,N_29275);
or UO_1772 (O_1772,N_29506,N_29356);
nor UO_1773 (O_1773,N_29248,N_29851);
nand UO_1774 (O_1774,N_29476,N_29263);
and UO_1775 (O_1775,N_29941,N_29731);
nor UO_1776 (O_1776,N_29993,N_29379);
xnor UO_1777 (O_1777,N_29058,N_29963);
nor UO_1778 (O_1778,N_29121,N_29082);
nor UO_1779 (O_1779,N_29572,N_29545);
nand UO_1780 (O_1780,N_29551,N_29016);
or UO_1781 (O_1781,N_29063,N_29299);
or UO_1782 (O_1782,N_29392,N_29965);
nand UO_1783 (O_1783,N_29898,N_29820);
and UO_1784 (O_1784,N_29900,N_29712);
nand UO_1785 (O_1785,N_29923,N_29704);
or UO_1786 (O_1786,N_29668,N_29763);
nand UO_1787 (O_1787,N_29264,N_29679);
nand UO_1788 (O_1788,N_29696,N_29342);
nor UO_1789 (O_1789,N_29141,N_29251);
nor UO_1790 (O_1790,N_29817,N_29999);
nand UO_1791 (O_1791,N_29949,N_29474);
nand UO_1792 (O_1792,N_29221,N_29491);
xnor UO_1793 (O_1793,N_29172,N_29711);
and UO_1794 (O_1794,N_29587,N_29371);
or UO_1795 (O_1795,N_29858,N_29663);
nand UO_1796 (O_1796,N_29269,N_29139);
and UO_1797 (O_1797,N_29951,N_29038);
and UO_1798 (O_1798,N_29193,N_29155);
nand UO_1799 (O_1799,N_29421,N_29472);
nand UO_1800 (O_1800,N_29341,N_29261);
nand UO_1801 (O_1801,N_29988,N_29871);
nand UO_1802 (O_1802,N_29030,N_29621);
and UO_1803 (O_1803,N_29006,N_29357);
or UO_1804 (O_1804,N_29048,N_29308);
xor UO_1805 (O_1805,N_29305,N_29154);
or UO_1806 (O_1806,N_29860,N_29145);
nor UO_1807 (O_1807,N_29658,N_29451);
or UO_1808 (O_1808,N_29792,N_29388);
nor UO_1809 (O_1809,N_29037,N_29792);
or UO_1810 (O_1810,N_29828,N_29463);
nand UO_1811 (O_1811,N_29896,N_29108);
or UO_1812 (O_1812,N_29859,N_29337);
nand UO_1813 (O_1813,N_29023,N_29827);
xnor UO_1814 (O_1814,N_29384,N_29798);
xnor UO_1815 (O_1815,N_29318,N_29379);
nor UO_1816 (O_1816,N_29243,N_29504);
xnor UO_1817 (O_1817,N_29325,N_29763);
nand UO_1818 (O_1818,N_29489,N_29421);
or UO_1819 (O_1819,N_29416,N_29378);
nand UO_1820 (O_1820,N_29357,N_29417);
nand UO_1821 (O_1821,N_29290,N_29272);
nand UO_1822 (O_1822,N_29084,N_29362);
xnor UO_1823 (O_1823,N_29475,N_29902);
xnor UO_1824 (O_1824,N_29208,N_29039);
or UO_1825 (O_1825,N_29718,N_29890);
nor UO_1826 (O_1826,N_29107,N_29411);
nor UO_1827 (O_1827,N_29934,N_29251);
and UO_1828 (O_1828,N_29783,N_29328);
or UO_1829 (O_1829,N_29682,N_29452);
nand UO_1830 (O_1830,N_29668,N_29033);
and UO_1831 (O_1831,N_29948,N_29003);
and UO_1832 (O_1832,N_29157,N_29211);
nand UO_1833 (O_1833,N_29422,N_29123);
nor UO_1834 (O_1834,N_29626,N_29269);
nor UO_1835 (O_1835,N_29729,N_29257);
and UO_1836 (O_1836,N_29036,N_29188);
or UO_1837 (O_1837,N_29945,N_29918);
and UO_1838 (O_1838,N_29064,N_29208);
xor UO_1839 (O_1839,N_29861,N_29567);
xnor UO_1840 (O_1840,N_29755,N_29117);
xor UO_1841 (O_1841,N_29944,N_29822);
or UO_1842 (O_1842,N_29232,N_29295);
or UO_1843 (O_1843,N_29572,N_29950);
or UO_1844 (O_1844,N_29172,N_29265);
or UO_1845 (O_1845,N_29032,N_29174);
nor UO_1846 (O_1846,N_29106,N_29079);
and UO_1847 (O_1847,N_29951,N_29029);
nand UO_1848 (O_1848,N_29649,N_29248);
nor UO_1849 (O_1849,N_29430,N_29790);
or UO_1850 (O_1850,N_29925,N_29568);
and UO_1851 (O_1851,N_29571,N_29039);
or UO_1852 (O_1852,N_29665,N_29481);
xor UO_1853 (O_1853,N_29837,N_29590);
nand UO_1854 (O_1854,N_29361,N_29640);
nor UO_1855 (O_1855,N_29661,N_29017);
and UO_1856 (O_1856,N_29908,N_29405);
xnor UO_1857 (O_1857,N_29406,N_29781);
or UO_1858 (O_1858,N_29046,N_29562);
nor UO_1859 (O_1859,N_29279,N_29176);
and UO_1860 (O_1860,N_29232,N_29055);
nor UO_1861 (O_1861,N_29618,N_29797);
xnor UO_1862 (O_1862,N_29947,N_29834);
xnor UO_1863 (O_1863,N_29097,N_29393);
nand UO_1864 (O_1864,N_29387,N_29539);
nor UO_1865 (O_1865,N_29370,N_29130);
xnor UO_1866 (O_1866,N_29034,N_29464);
xor UO_1867 (O_1867,N_29784,N_29185);
nor UO_1868 (O_1868,N_29562,N_29585);
nor UO_1869 (O_1869,N_29857,N_29436);
nand UO_1870 (O_1870,N_29097,N_29054);
xor UO_1871 (O_1871,N_29415,N_29301);
nand UO_1872 (O_1872,N_29465,N_29544);
nor UO_1873 (O_1873,N_29442,N_29024);
or UO_1874 (O_1874,N_29919,N_29626);
nor UO_1875 (O_1875,N_29764,N_29627);
or UO_1876 (O_1876,N_29428,N_29878);
nor UO_1877 (O_1877,N_29942,N_29067);
xor UO_1878 (O_1878,N_29611,N_29432);
nand UO_1879 (O_1879,N_29549,N_29339);
and UO_1880 (O_1880,N_29148,N_29522);
or UO_1881 (O_1881,N_29425,N_29278);
or UO_1882 (O_1882,N_29553,N_29440);
or UO_1883 (O_1883,N_29071,N_29470);
nand UO_1884 (O_1884,N_29745,N_29756);
nor UO_1885 (O_1885,N_29972,N_29678);
nor UO_1886 (O_1886,N_29481,N_29149);
xnor UO_1887 (O_1887,N_29055,N_29364);
xor UO_1888 (O_1888,N_29898,N_29750);
or UO_1889 (O_1889,N_29998,N_29083);
and UO_1890 (O_1890,N_29861,N_29740);
and UO_1891 (O_1891,N_29954,N_29334);
and UO_1892 (O_1892,N_29021,N_29340);
nor UO_1893 (O_1893,N_29064,N_29626);
and UO_1894 (O_1894,N_29536,N_29079);
or UO_1895 (O_1895,N_29651,N_29158);
xor UO_1896 (O_1896,N_29029,N_29385);
nor UO_1897 (O_1897,N_29051,N_29496);
or UO_1898 (O_1898,N_29870,N_29677);
nor UO_1899 (O_1899,N_29164,N_29405);
and UO_1900 (O_1900,N_29045,N_29952);
nand UO_1901 (O_1901,N_29369,N_29368);
xor UO_1902 (O_1902,N_29911,N_29704);
nand UO_1903 (O_1903,N_29907,N_29267);
xor UO_1904 (O_1904,N_29766,N_29397);
xor UO_1905 (O_1905,N_29745,N_29083);
or UO_1906 (O_1906,N_29455,N_29353);
or UO_1907 (O_1907,N_29248,N_29490);
xnor UO_1908 (O_1908,N_29894,N_29165);
and UO_1909 (O_1909,N_29238,N_29958);
xnor UO_1910 (O_1910,N_29588,N_29039);
or UO_1911 (O_1911,N_29185,N_29839);
or UO_1912 (O_1912,N_29646,N_29027);
nand UO_1913 (O_1913,N_29483,N_29721);
nand UO_1914 (O_1914,N_29270,N_29035);
or UO_1915 (O_1915,N_29229,N_29556);
nand UO_1916 (O_1916,N_29000,N_29229);
nor UO_1917 (O_1917,N_29474,N_29883);
nand UO_1918 (O_1918,N_29193,N_29310);
nand UO_1919 (O_1919,N_29652,N_29558);
or UO_1920 (O_1920,N_29472,N_29796);
or UO_1921 (O_1921,N_29376,N_29966);
and UO_1922 (O_1922,N_29782,N_29390);
nand UO_1923 (O_1923,N_29947,N_29058);
xnor UO_1924 (O_1924,N_29338,N_29919);
nand UO_1925 (O_1925,N_29282,N_29878);
nor UO_1926 (O_1926,N_29378,N_29901);
xor UO_1927 (O_1927,N_29760,N_29845);
or UO_1928 (O_1928,N_29503,N_29600);
or UO_1929 (O_1929,N_29393,N_29977);
nand UO_1930 (O_1930,N_29688,N_29194);
nand UO_1931 (O_1931,N_29484,N_29294);
and UO_1932 (O_1932,N_29730,N_29242);
xnor UO_1933 (O_1933,N_29060,N_29415);
nand UO_1934 (O_1934,N_29722,N_29322);
nor UO_1935 (O_1935,N_29615,N_29476);
nor UO_1936 (O_1936,N_29101,N_29981);
nor UO_1937 (O_1937,N_29917,N_29314);
and UO_1938 (O_1938,N_29521,N_29885);
and UO_1939 (O_1939,N_29010,N_29699);
xnor UO_1940 (O_1940,N_29923,N_29062);
nor UO_1941 (O_1941,N_29593,N_29341);
and UO_1942 (O_1942,N_29391,N_29310);
xor UO_1943 (O_1943,N_29309,N_29701);
nor UO_1944 (O_1944,N_29784,N_29306);
and UO_1945 (O_1945,N_29837,N_29282);
nor UO_1946 (O_1946,N_29670,N_29233);
or UO_1947 (O_1947,N_29449,N_29865);
nor UO_1948 (O_1948,N_29778,N_29351);
and UO_1949 (O_1949,N_29031,N_29866);
and UO_1950 (O_1950,N_29432,N_29351);
nand UO_1951 (O_1951,N_29349,N_29283);
and UO_1952 (O_1952,N_29943,N_29048);
and UO_1953 (O_1953,N_29183,N_29531);
xnor UO_1954 (O_1954,N_29324,N_29899);
nand UO_1955 (O_1955,N_29881,N_29037);
or UO_1956 (O_1956,N_29426,N_29504);
xnor UO_1957 (O_1957,N_29034,N_29841);
xor UO_1958 (O_1958,N_29712,N_29862);
nor UO_1959 (O_1959,N_29947,N_29539);
nor UO_1960 (O_1960,N_29251,N_29223);
or UO_1961 (O_1961,N_29674,N_29332);
nand UO_1962 (O_1962,N_29881,N_29834);
xor UO_1963 (O_1963,N_29715,N_29599);
or UO_1964 (O_1964,N_29427,N_29885);
and UO_1965 (O_1965,N_29172,N_29139);
or UO_1966 (O_1966,N_29854,N_29995);
nand UO_1967 (O_1967,N_29548,N_29938);
nand UO_1968 (O_1968,N_29430,N_29781);
and UO_1969 (O_1969,N_29969,N_29413);
and UO_1970 (O_1970,N_29815,N_29290);
nand UO_1971 (O_1971,N_29525,N_29048);
nor UO_1972 (O_1972,N_29623,N_29476);
xor UO_1973 (O_1973,N_29713,N_29161);
xor UO_1974 (O_1974,N_29461,N_29883);
or UO_1975 (O_1975,N_29817,N_29574);
and UO_1976 (O_1976,N_29333,N_29585);
and UO_1977 (O_1977,N_29418,N_29923);
xor UO_1978 (O_1978,N_29421,N_29232);
xnor UO_1979 (O_1979,N_29568,N_29026);
or UO_1980 (O_1980,N_29539,N_29029);
or UO_1981 (O_1981,N_29628,N_29062);
xor UO_1982 (O_1982,N_29560,N_29621);
and UO_1983 (O_1983,N_29662,N_29527);
nand UO_1984 (O_1984,N_29222,N_29009);
or UO_1985 (O_1985,N_29593,N_29265);
or UO_1986 (O_1986,N_29478,N_29510);
nand UO_1987 (O_1987,N_29899,N_29972);
xnor UO_1988 (O_1988,N_29631,N_29983);
or UO_1989 (O_1989,N_29092,N_29510);
or UO_1990 (O_1990,N_29463,N_29577);
nand UO_1991 (O_1991,N_29306,N_29134);
or UO_1992 (O_1992,N_29594,N_29956);
nand UO_1993 (O_1993,N_29437,N_29028);
nand UO_1994 (O_1994,N_29218,N_29846);
xnor UO_1995 (O_1995,N_29065,N_29369);
or UO_1996 (O_1996,N_29088,N_29494);
or UO_1997 (O_1997,N_29783,N_29787);
nand UO_1998 (O_1998,N_29066,N_29883);
nor UO_1999 (O_1999,N_29597,N_29162);
and UO_2000 (O_2000,N_29584,N_29790);
xor UO_2001 (O_2001,N_29039,N_29577);
xor UO_2002 (O_2002,N_29210,N_29802);
nor UO_2003 (O_2003,N_29393,N_29954);
xnor UO_2004 (O_2004,N_29464,N_29503);
nand UO_2005 (O_2005,N_29479,N_29216);
xnor UO_2006 (O_2006,N_29596,N_29437);
xor UO_2007 (O_2007,N_29239,N_29967);
xor UO_2008 (O_2008,N_29018,N_29501);
nor UO_2009 (O_2009,N_29139,N_29576);
or UO_2010 (O_2010,N_29539,N_29169);
nand UO_2011 (O_2011,N_29937,N_29486);
or UO_2012 (O_2012,N_29201,N_29735);
nor UO_2013 (O_2013,N_29554,N_29167);
nor UO_2014 (O_2014,N_29448,N_29620);
nand UO_2015 (O_2015,N_29503,N_29373);
nand UO_2016 (O_2016,N_29591,N_29178);
nand UO_2017 (O_2017,N_29723,N_29909);
and UO_2018 (O_2018,N_29176,N_29152);
xor UO_2019 (O_2019,N_29115,N_29604);
nand UO_2020 (O_2020,N_29842,N_29002);
nand UO_2021 (O_2021,N_29511,N_29778);
and UO_2022 (O_2022,N_29047,N_29104);
xnor UO_2023 (O_2023,N_29563,N_29560);
xor UO_2024 (O_2024,N_29300,N_29055);
nor UO_2025 (O_2025,N_29647,N_29267);
xor UO_2026 (O_2026,N_29148,N_29097);
or UO_2027 (O_2027,N_29630,N_29079);
nand UO_2028 (O_2028,N_29555,N_29438);
nor UO_2029 (O_2029,N_29365,N_29971);
or UO_2030 (O_2030,N_29302,N_29722);
nand UO_2031 (O_2031,N_29644,N_29897);
nand UO_2032 (O_2032,N_29573,N_29562);
and UO_2033 (O_2033,N_29518,N_29853);
and UO_2034 (O_2034,N_29556,N_29773);
nor UO_2035 (O_2035,N_29729,N_29016);
and UO_2036 (O_2036,N_29211,N_29861);
and UO_2037 (O_2037,N_29480,N_29474);
and UO_2038 (O_2038,N_29584,N_29373);
nand UO_2039 (O_2039,N_29742,N_29119);
and UO_2040 (O_2040,N_29440,N_29847);
xnor UO_2041 (O_2041,N_29472,N_29522);
and UO_2042 (O_2042,N_29240,N_29200);
xnor UO_2043 (O_2043,N_29860,N_29193);
nor UO_2044 (O_2044,N_29735,N_29422);
and UO_2045 (O_2045,N_29427,N_29796);
or UO_2046 (O_2046,N_29587,N_29092);
or UO_2047 (O_2047,N_29121,N_29299);
nor UO_2048 (O_2048,N_29361,N_29404);
xor UO_2049 (O_2049,N_29222,N_29973);
xnor UO_2050 (O_2050,N_29538,N_29341);
xor UO_2051 (O_2051,N_29188,N_29056);
and UO_2052 (O_2052,N_29999,N_29616);
nand UO_2053 (O_2053,N_29338,N_29995);
and UO_2054 (O_2054,N_29867,N_29916);
xor UO_2055 (O_2055,N_29719,N_29245);
xnor UO_2056 (O_2056,N_29174,N_29837);
xor UO_2057 (O_2057,N_29551,N_29116);
nand UO_2058 (O_2058,N_29537,N_29202);
nand UO_2059 (O_2059,N_29968,N_29876);
or UO_2060 (O_2060,N_29894,N_29998);
and UO_2061 (O_2061,N_29732,N_29210);
and UO_2062 (O_2062,N_29920,N_29232);
xor UO_2063 (O_2063,N_29605,N_29337);
nor UO_2064 (O_2064,N_29104,N_29847);
and UO_2065 (O_2065,N_29194,N_29584);
nand UO_2066 (O_2066,N_29029,N_29698);
nor UO_2067 (O_2067,N_29217,N_29227);
or UO_2068 (O_2068,N_29907,N_29904);
or UO_2069 (O_2069,N_29331,N_29027);
nand UO_2070 (O_2070,N_29942,N_29880);
nand UO_2071 (O_2071,N_29206,N_29277);
and UO_2072 (O_2072,N_29345,N_29199);
and UO_2073 (O_2073,N_29427,N_29589);
xor UO_2074 (O_2074,N_29022,N_29092);
xor UO_2075 (O_2075,N_29602,N_29656);
or UO_2076 (O_2076,N_29925,N_29204);
and UO_2077 (O_2077,N_29039,N_29022);
and UO_2078 (O_2078,N_29472,N_29788);
xnor UO_2079 (O_2079,N_29217,N_29317);
xnor UO_2080 (O_2080,N_29266,N_29713);
xnor UO_2081 (O_2081,N_29553,N_29939);
xor UO_2082 (O_2082,N_29584,N_29750);
or UO_2083 (O_2083,N_29278,N_29959);
or UO_2084 (O_2084,N_29049,N_29157);
or UO_2085 (O_2085,N_29587,N_29594);
nor UO_2086 (O_2086,N_29963,N_29193);
and UO_2087 (O_2087,N_29656,N_29534);
nor UO_2088 (O_2088,N_29895,N_29932);
nand UO_2089 (O_2089,N_29283,N_29331);
and UO_2090 (O_2090,N_29626,N_29131);
nor UO_2091 (O_2091,N_29262,N_29618);
and UO_2092 (O_2092,N_29232,N_29513);
nand UO_2093 (O_2093,N_29983,N_29542);
nor UO_2094 (O_2094,N_29912,N_29234);
nand UO_2095 (O_2095,N_29588,N_29935);
nand UO_2096 (O_2096,N_29607,N_29271);
or UO_2097 (O_2097,N_29655,N_29139);
or UO_2098 (O_2098,N_29020,N_29963);
or UO_2099 (O_2099,N_29232,N_29606);
nand UO_2100 (O_2100,N_29650,N_29324);
nor UO_2101 (O_2101,N_29792,N_29786);
xor UO_2102 (O_2102,N_29418,N_29790);
and UO_2103 (O_2103,N_29247,N_29480);
nand UO_2104 (O_2104,N_29141,N_29427);
xor UO_2105 (O_2105,N_29220,N_29508);
xnor UO_2106 (O_2106,N_29102,N_29088);
nor UO_2107 (O_2107,N_29354,N_29411);
nand UO_2108 (O_2108,N_29716,N_29560);
nor UO_2109 (O_2109,N_29808,N_29201);
nor UO_2110 (O_2110,N_29380,N_29484);
nand UO_2111 (O_2111,N_29947,N_29723);
nand UO_2112 (O_2112,N_29784,N_29087);
and UO_2113 (O_2113,N_29575,N_29607);
and UO_2114 (O_2114,N_29564,N_29335);
and UO_2115 (O_2115,N_29939,N_29466);
or UO_2116 (O_2116,N_29163,N_29671);
nor UO_2117 (O_2117,N_29109,N_29480);
xnor UO_2118 (O_2118,N_29542,N_29977);
or UO_2119 (O_2119,N_29082,N_29009);
and UO_2120 (O_2120,N_29555,N_29450);
xor UO_2121 (O_2121,N_29373,N_29357);
xnor UO_2122 (O_2122,N_29817,N_29274);
nor UO_2123 (O_2123,N_29891,N_29174);
or UO_2124 (O_2124,N_29010,N_29393);
and UO_2125 (O_2125,N_29954,N_29448);
nand UO_2126 (O_2126,N_29274,N_29670);
nand UO_2127 (O_2127,N_29696,N_29168);
or UO_2128 (O_2128,N_29665,N_29026);
or UO_2129 (O_2129,N_29171,N_29722);
or UO_2130 (O_2130,N_29399,N_29051);
and UO_2131 (O_2131,N_29710,N_29638);
and UO_2132 (O_2132,N_29406,N_29706);
or UO_2133 (O_2133,N_29597,N_29681);
and UO_2134 (O_2134,N_29804,N_29731);
nor UO_2135 (O_2135,N_29001,N_29864);
nand UO_2136 (O_2136,N_29033,N_29426);
nand UO_2137 (O_2137,N_29594,N_29735);
nand UO_2138 (O_2138,N_29575,N_29085);
nor UO_2139 (O_2139,N_29448,N_29103);
and UO_2140 (O_2140,N_29179,N_29178);
and UO_2141 (O_2141,N_29851,N_29882);
or UO_2142 (O_2142,N_29198,N_29412);
xnor UO_2143 (O_2143,N_29585,N_29383);
xor UO_2144 (O_2144,N_29943,N_29286);
xor UO_2145 (O_2145,N_29697,N_29433);
nor UO_2146 (O_2146,N_29048,N_29774);
or UO_2147 (O_2147,N_29766,N_29162);
nor UO_2148 (O_2148,N_29373,N_29456);
xor UO_2149 (O_2149,N_29887,N_29048);
nor UO_2150 (O_2150,N_29511,N_29063);
or UO_2151 (O_2151,N_29500,N_29014);
and UO_2152 (O_2152,N_29152,N_29873);
xor UO_2153 (O_2153,N_29007,N_29314);
nand UO_2154 (O_2154,N_29787,N_29193);
nor UO_2155 (O_2155,N_29732,N_29996);
or UO_2156 (O_2156,N_29866,N_29611);
and UO_2157 (O_2157,N_29081,N_29759);
and UO_2158 (O_2158,N_29805,N_29355);
or UO_2159 (O_2159,N_29167,N_29958);
nor UO_2160 (O_2160,N_29119,N_29385);
or UO_2161 (O_2161,N_29509,N_29355);
xnor UO_2162 (O_2162,N_29614,N_29595);
xnor UO_2163 (O_2163,N_29289,N_29398);
nor UO_2164 (O_2164,N_29687,N_29995);
nand UO_2165 (O_2165,N_29217,N_29767);
or UO_2166 (O_2166,N_29664,N_29719);
nor UO_2167 (O_2167,N_29583,N_29598);
nand UO_2168 (O_2168,N_29881,N_29466);
xnor UO_2169 (O_2169,N_29100,N_29151);
nand UO_2170 (O_2170,N_29157,N_29027);
nand UO_2171 (O_2171,N_29394,N_29805);
xnor UO_2172 (O_2172,N_29811,N_29913);
xnor UO_2173 (O_2173,N_29468,N_29533);
or UO_2174 (O_2174,N_29508,N_29050);
nor UO_2175 (O_2175,N_29145,N_29848);
nor UO_2176 (O_2176,N_29169,N_29979);
or UO_2177 (O_2177,N_29920,N_29223);
nand UO_2178 (O_2178,N_29797,N_29553);
nor UO_2179 (O_2179,N_29374,N_29729);
and UO_2180 (O_2180,N_29463,N_29146);
xor UO_2181 (O_2181,N_29009,N_29872);
nand UO_2182 (O_2182,N_29816,N_29688);
and UO_2183 (O_2183,N_29050,N_29389);
nand UO_2184 (O_2184,N_29735,N_29122);
and UO_2185 (O_2185,N_29139,N_29663);
nor UO_2186 (O_2186,N_29763,N_29687);
xnor UO_2187 (O_2187,N_29891,N_29354);
nand UO_2188 (O_2188,N_29729,N_29445);
nand UO_2189 (O_2189,N_29162,N_29748);
nor UO_2190 (O_2190,N_29361,N_29428);
and UO_2191 (O_2191,N_29112,N_29101);
or UO_2192 (O_2192,N_29883,N_29081);
xor UO_2193 (O_2193,N_29047,N_29819);
or UO_2194 (O_2194,N_29102,N_29034);
xnor UO_2195 (O_2195,N_29837,N_29005);
xnor UO_2196 (O_2196,N_29457,N_29141);
or UO_2197 (O_2197,N_29904,N_29929);
or UO_2198 (O_2198,N_29636,N_29649);
nand UO_2199 (O_2199,N_29711,N_29665);
and UO_2200 (O_2200,N_29631,N_29286);
nor UO_2201 (O_2201,N_29604,N_29423);
and UO_2202 (O_2202,N_29789,N_29089);
nand UO_2203 (O_2203,N_29628,N_29406);
and UO_2204 (O_2204,N_29335,N_29938);
xor UO_2205 (O_2205,N_29649,N_29424);
or UO_2206 (O_2206,N_29413,N_29531);
nor UO_2207 (O_2207,N_29874,N_29947);
xnor UO_2208 (O_2208,N_29756,N_29589);
xnor UO_2209 (O_2209,N_29795,N_29019);
xnor UO_2210 (O_2210,N_29146,N_29175);
and UO_2211 (O_2211,N_29741,N_29931);
nand UO_2212 (O_2212,N_29099,N_29732);
xnor UO_2213 (O_2213,N_29494,N_29685);
or UO_2214 (O_2214,N_29477,N_29280);
nand UO_2215 (O_2215,N_29023,N_29490);
nor UO_2216 (O_2216,N_29764,N_29007);
and UO_2217 (O_2217,N_29953,N_29698);
nor UO_2218 (O_2218,N_29611,N_29391);
nand UO_2219 (O_2219,N_29365,N_29181);
or UO_2220 (O_2220,N_29156,N_29820);
xor UO_2221 (O_2221,N_29546,N_29209);
xor UO_2222 (O_2222,N_29581,N_29304);
or UO_2223 (O_2223,N_29877,N_29607);
or UO_2224 (O_2224,N_29325,N_29302);
and UO_2225 (O_2225,N_29819,N_29044);
and UO_2226 (O_2226,N_29129,N_29873);
or UO_2227 (O_2227,N_29873,N_29977);
xnor UO_2228 (O_2228,N_29843,N_29768);
xor UO_2229 (O_2229,N_29451,N_29831);
and UO_2230 (O_2230,N_29990,N_29591);
or UO_2231 (O_2231,N_29659,N_29235);
xor UO_2232 (O_2232,N_29232,N_29504);
nor UO_2233 (O_2233,N_29980,N_29896);
xnor UO_2234 (O_2234,N_29357,N_29019);
nand UO_2235 (O_2235,N_29855,N_29433);
or UO_2236 (O_2236,N_29752,N_29106);
nor UO_2237 (O_2237,N_29218,N_29171);
nor UO_2238 (O_2238,N_29209,N_29058);
or UO_2239 (O_2239,N_29121,N_29761);
or UO_2240 (O_2240,N_29820,N_29504);
xor UO_2241 (O_2241,N_29319,N_29037);
nor UO_2242 (O_2242,N_29913,N_29874);
or UO_2243 (O_2243,N_29517,N_29285);
nand UO_2244 (O_2244,N_29767,N_29171);
xnor UO_2245 (O_2245,N_29798,N_29247);
nand UO_2246 (O_2246,N_29007,N_29550);
or UO_2247 (O_2247,N_29510,N_29364);
nand UO_2248 (O_2248,N_29513,N_29093);
xor UO_2249 (O_2249,N_29823,N_29599);
nand UO_2250 (O_2250,N_29296,N_29224);
or UO_2251 (O_2251,N_29650,N_29784);
nand UO_2252 (O_2252,N_29577,N_29031);
and UO_2253 (O_2253,N_29221,N_29153);
and UO_2254 (O_2254,N_29441,N_29756);
or UO_2255 (O_2255,N_29667,N_29393);
nor UO_2256 (O_2256,N_29350,N_29773);
xnor UO_2257 (O_2257,N_29347,N_29523);
xnor UO_2258 (O_2258,N_29337,N_29134);
xor UO_2259 (O_2259,N_29677,N_29983);
and UO_2260 (O_2260,N_29801,N_29090);
or UO_2261 (O_2261,N_29148,N_29848);
or UO_2262 (O_2262,N_29141,N_29037);
and UO_2263 (O_2263,N_29419,N_29271);
and UO_2264 (O_2264,N_29797,N_29559);
xnor UO_2265 (O_2265,N_29202,N_29396);
or UO_2266 (O_2266,N_29373,N_29834);
nand UO_2267 (O_2267,N_29048,N_29966);
nand UO_2268 (O_2268,N_29144,N_29568);
nor UO_2269 (O_2269,N_29501,N_29259);
and UO_2270 (O_2270,N_29231,N_29958);
nand UO_2271 (O_2271,N_29629,N_29600);
nor UO_2272 (O_2272,N_29936,N_29949);
nand UO_2273 (O_2273,N_29916,N_29795);
nor UO_2274 (O_2274,N_29181,N_29742);
xnor UO_2275 (O_2275,N_29023,N_29440);
and UO_2276 (O_2276,N_29072,N_29497);
nor UO_2277 (O_2277,N_29679,N_29726);
nand UO_2278 (O_2278,N_29793,N_29278);
nor UO_2279 (O_2279,N_29796,N_29444);
or UO_2280 (O_2280,N_29300,N_29739);
and UO_2281 (O_2281,N_29461,N_29127);
or UO_2282 (O_2282,N_29692,N_29807);
and UO_2283 (O_2283,N_29802,N_29858);
nand UO_2284 (O_2284,N_29814,N_29630);
or UO_2285 (O_2285,N_29706,N_29868);
nand UO_2286 (O_2286,N_29441,N_29889);
xnor UO_2287 (O_2287,N_29738,N_29864);
xnor UO_2288 (O_2288,N_29979,N_29952);
nor UO_2289 (O_2289,N_29181,N_29081);
nand UO_2290 (O_2290,N_29855,N_29114);
xor UO_2291 (O_2291,N_29353,N_29226);
xor UO_2292 (O_2292,N_29898,N_29582);
or UO_2293 (O_2293,N_29973,N_29366);
nand UO_2294 (O_2294,N_29015,N_29599);
nand UO_2295 (O_2295,N_29721,N_29340);
nand UO_2296 (O_2296,N_29365,N_29908);
and UO_2297 (O_2297,N_29522,N_29320);
or UO_2298 (O_2298,N_29999,N_29874);
nand UO_2299 (O_2299,N_29070,N_29964);
xor UO_2300 (O_2300,N_29499,N_29531);
and UO_2301 (O_2301,N_29103,N_29542);
or UO_2302 (O_2302,N_29730,N_29975);
xor UO_2303 (O_2303,N_29084,N_29034);
nand UO_2304 (O_2304,N_29732,N_29550);
or UO_2305 (O_2305,N_29154,N_29434);
and UO_2306 (O_2306,N_29495,N_29871);
nand UO_2307 (O_2307,N_29727,N_29587);
or UO_2308 (O_2308,N_29631,N_29173);
nand UO_2309 (O_2309,N_29589,N_29592);
or UO_2310 (O_2310,N_29798,N_29217);
xnor UO_2311 (O_2311,N_29712,N_29219);
xnor UO_2312 (O_2312,N_29592,N_29687);
nand UO_2313 (O_2313,N_29161,N_29846);
or UO_2314 (O_2314,N_29602,N_29573);
or UO_2315 (O_2315,N_29645,N_29170);
and UO_2316 (O_2316,N_29234,N_29407);
or UO_2317 (O_2317,N_29677,N_29468);
xnor UO_2318 (O_2318,N_29475,N_29582);
nand UO_2319 (O_2319,N_29385,N_29205);
and UO_2320 (O_2320,N_29985,N_29418);
or UO_2321 (O_2321,N_29582,N_29552);
or UO_2322 (O_2322,N_29945,N_29572);
nor UO_2323 (O_2323,N_29234,N_29603);
nand UO_2324 (O_2324,N_29270,N_29667);
nor UO_2325 (O_2325,N_29941,N_29612);
and UO_2326 (O_2326,N_29108,N_29153);
or UO_2327 (O_2327,N_29971,N_29200);
nand UO_2328 (O_2328,N_29271,N_29074);
and UO_2329 (O_2329,N_29965,N_29849);
nand UO_2330 (O_2330,N_29792,N_29273);
or UO_2331 (O_2331,N_29760,N_29613);
nor UO_2332 (O_2332,N_29221,N_29087);
xnor UO_2333 (O_2333,N_29006,N_29759);
xor UO_2334 (O_2334,N_29801,N_29644);
or UO_2335 (O_2335,N_29563,N_29620);
nand UO_2336 (O_2336,N_29385,N_29208);
nand UO_2337 (O_2337,N_29184,N_29138);
nand UO_2338 (O_2338,N_29573,N_29069);
xnor UO_2339 (O_2339,N_29465,N_29747);
nor UO_2340 (O_2340,N_29741,N_29246);
nand UO_2341 (O_2341,N_29285,N_29686);
or UO_2342 (O_2342,N_29304,N_29249);
xor UO_2343 (O_2343,N_29196,N_29771);
and UO_2344 (O_2344,N_29540,N_29028);
nand UO_2345 (O_2345,N_29992,N_29894);
nor UO_2346 (O_2346,N_29252,N_29602);
nand UO_2347 (O_2347,N_29713,N_29322);
xor UO_2348 (O_2348,N_29483,N_29319);
xor UO_2349 (O_2349,N_29017,N_29291);
and UO_2350 (O_2350,N_29466,N_29889);
nor UO_2351 (O_2351,N_29409,N_29738);
nor UO_2352 (O_2352,N_29907,N_29145);
xnor UO_2353 (O_2353,N_29705,N_29225);
nand UO_2354 (O_2354,N_29267,N_29154);
nor UO_2355 (O_2355,N_29347,N_29713);
nor UO_2356 (O_2356,N_29027,N_29343);
nor UO_2357 (O_2357,N_29344,N_29899);
xor UO_2358 (O_2358,N_29853,N_29144);
nor UO_2359 (O_2359,N_29336,N_29988);
xnor UO_2360 (O_2360,N_29038,N_29187);
and UO_2361 (O_2361,N_29951,N_29690);
nor UO_2362 (O_2362,N_29547,N_29313);
xor UO_2363 (O_2363,N_29382,N_29587);
nand UO_2364 (O_2364,N_29481,N_29522);
or UO_2365 (O_2365,N_29286,N_29529);
and UO_2366 (O_2366,N_29588,N_29628);
nor UO_2367 (O_2367,N_29074,N_29464);
and UO_2368 (O_2368,N_29438,N_29601);
or UO_2369 (O_2369,N_29435,N_29571);
and UO_2370 (O_2370,N_29363,N_29285);
xor UO_2371 (O_2371,N_29713,N_29991);
and UO_2372 (O_2372,N_29167,N_29593);
nor UO_2373 (O_2373,N_29325,N_29601);
xnor UO_2374 (O_2374,N_29058,N_29653);
and UO_2375 (O_2375,N_29426,N_29779);
or UO_2376 (O_2376,N_29650,N_29130);
or UO_2377 (O_2377,N_29145,N_29188);
xnor UO_2378 (O_2378,N_29754,N_29071);
xnor UO_2379 (O_2379,N_29788,N_29580);
or UO_2380 (O_2380,N_29802,N_29052);
nor UO_2381 (O_2381,N_29190,N_29103);
nor UO_2382 (O_2382,N_29078,N_29456);
and UO_2383 (O_2383,N_29381,N_29654);
nand UO_2384 (O_2384,N_29162,N_29244);
nor UO_2385 (O_2385,N_29122,N_29531);
nand UO_2386 (O_2386,N_29434,N_29316);
or UO_2387 (O_2387,N_29094,N_29621);
xor UO_2388 (O_2388,N_29275,N_29295);
nand UO_2389 (O_2389,N_29413,N_29845);
and UO_2390 (O_2390,N_29660,N_29409);
nor UO_2391 (O_2391,N_29310,N_29649);
and UO_2392 (O_2392,N_29537,N_29108);
and UO_2393 (O_2393,N_29600,N_29143);
and UO_2394 (O_2394,N_29914,N_29317);
nor UO_2395 (O_2395,N_29788,N_29810);
nor UO_2396 (O_2396,N_29843,N_29687);
and UO_2397 (O_2397,N_29212,N_29537);
xnor UO_2398 (O_2398,N_29465,N_29605);
or UO_2399 (O_2399,N_29706,N_29570);
nand UO_2400 (O_2400,N_29237,N_29130);
nand UO_2401 (O_2401,N_29526,N_29080);
or UO_2402 (O_2402,N_29020,N_29821);
and UO_2403 (O_2403,N_29284,N_29537);
nand UO_2404 (O_2404,N_29243,N_29240);
and UO_2405 (O_2405,N_29926,N_29365);
xnor UO_2406 (O_2406,N_29869,N_29261);
and UO_2407 (O_2407,N_29247,N_29057);
nand UO_2408 (O_2408,N_29169,N_29126);
and UO_2409 (O_2409,N_29004,N_29755);
or UO_2410 (O_2410,N_29481,N_29215);
and UO_2411 (O_2411,N_29279,N_29867);
nor UO_2412 (O_2412,N_29462,N_29917);
nor UO_2413 (O_2413,N_29971,N_29471);
and UO_2414 (O_2414,N_29724,N_29765);
nor UO_2415 (O_2415,N_29252,N_29950);
xnor UO_2416 (O_2416,N_29970,N_29807);
nand UO_2417 (O_2417,N_29905,N_29662);
xor UO_2418 (O_2418,N_29221,N_29826);
xnor UO_2419 (O_2419,N_29734,N_29652);
nand UO_2420 (O_2420,N_29353,N_29770);
nand UO_2421 (O_2421,N_29441,N_29975);
nor UO_2422 (O_2422,N_29416,N_29118);
and UO_2423 (O_2423,N_29362,N_29055);
and UO_2424 (O_2424,N_29597,N_29343);
or UO_2425 (O_2425,N_29294,N_29278);
nor UO_2426 (O_2426,N_29459,N_29230);
and UO_2427 (O_2427,N_29473,N_29323);
and UO_2428 (O_2428,N_29762,N_29516);
nor UO_2429 (O_2429,N_29162,N_29119);
or UO_2430 (O_2430,N_29843,N_29914);
nor UO_2431 (O_2431,N_29147,N_29444);
or UO_2432 (O_2432,N_29999,N_29412);
xnor UO_2433 (O_2433,N_29515,N_29020);
nand UO_2434 (O_2434,N_29211,N_29356);
and UO_2435 (O_2435,N_29029,N_29716);
and UO_2436 (O_2436,N_29055,N_29188);
xnor UO_2437 (O_2437,N_29838,N_29715);
and UO_2438 (O_2438,N_29020,N_29909);
nor UO_2439 (O_2439,N_29999,N_29250);
or UO_2440 (O_2440,N_29885,N_29618);
and UO_2441 (O_2441,N_29582,N_29598);
nand UO_2442 (O_2442,N_29741,N_29427);
and UO_2443 (O_2443,N_29548,N_29524);
or UO_2444 (O_2444,N_29533,N_29389);
and UO_2445 (O_2445,N_29681,N_29446);
nor UO_2446 (O_2446,N_29604,N_29486);
nor UO_2447 (O_2447,N_29883,N_29953);
and UO_2448 (O_2448,N_29846,N_29452);
xor UO_2449 (O_2449,N_29674,N_29472);
nor UO_2450 (O_2450,N_29149,N_29161);
nand UO_2451 (O_2451,N_29709,N_29571);
or UO_2452 (O_2452,N_29026,N_29390);
and UO_2453 (O_2453,N_29814,N_29922);
xnor UO_2454 (O_2454,N_29574,N_29255);
or UO_2455 (O_2455,N_29246,N_29260);
nor UO_2456 (O_2456,N_29683,N_29693);
or UO_2457 (O_2457,N_29594,N_29892);
and UO_2458 (O_2458,N_29296,N_29092);
and UO_2459 (O_2459,N_29893,N_29825);
xnor UO_2460 (O_2460,N_29848,N_29876);
xor UO_2461 (O_2461,N_29302,N_29494);
xnor UO_2462 (O_2462,N_29291,N_29099);
and UO_2463 (O_2463,N_29926,N_29585);
xor UO_2464 (O_2464,N_29273,N_29431);
nor UO_2465 (O_2465,N_29506,N_29139);
xor UO_2466 (O_2466,N_29802,N_29989);
xor UO_2467 (O_2467,N_29734,N_29319);
or UO_2468 (O_2468,N_29327,N_29722);
nand UO_2469 (O_2469,N_29009,N_29925);
nor UO_2470 (O_2470,N_29875,N_29944);
xor UO_2471 (O_2471,N_29344,N_29545);
and UO_2472 (O_2472,N_29624,N_29780);
nor UO_2473 (O_2473,N_29733,N_29079);
or UO_2474 (O_2474,N_29786,N_29330);
or UO_2475 (O_2475,N_29725,N_29038);
nor UO_2476 (O_2476,N_29177,N_29449);
xor UO_2477 (O_2477,N_29707,N_29115);
and UO_2478 (O_2478,N_29920,N_29605);
and UO_2479 (O_2479,N_29989,N_29611);
xnor UO_2480 (O_2480,N_29011,N_29970);
nand UO_2481 (O_2481,N_29635,N_29346);
or UO_2482 (O_2482,N_29459,N_29349);
or UO_2483 (O_2483,N_29116,N_29647);
and UO_2484 (O_2484,N_29891,N_29158);
nor UO_2485 (O_2485,N_29886,N_29222);
or UO_2486 (O_2486,N_29426,N_29193);
nand UO_2487 (O_2487,N_29300,N_29529);
nand UO_2488 (O_2488,N_29139,N_29462);
or UO_2489 (O_2489,N_29991,N_29817);
and UO_2490 (O_2490,N_29729,N_29643);
and UO_2491 (O_2491,N_29451,N_29612);
and UO_2492 (O_2492,N_29805,N_29617);
nor UO_2493 (O_2493,N_29175,N_29914);
xnor UO_2494 (O_2494,N_29569,N_29666);
nand UO_2495 (O_2495,N_29365,N_29476);
xnor UO_2496 (O_2496,N_29753,N_29937);
or UO_2497 (O_2497,N_29447,N_29185);
and UO_2498 (O_2498,N_29089,N_29693);
nor UO_2499 (O_2499,N_29037,N_29039);
and UO_2500 (O_2500,N_29996,N_29967);
nor UO_2501 (O_2501,N_29802,N_29509);
nor UO_2502 (O_2502,N_29507,N_29209);
or UO_2503 (O_2503,N_29374,N_29458);
nor UO_2504 (O_2504,N_29234,N_29405);
xor UO_2505 (O_2505,N_29250,N_29893);
nand UO_2506 (O_2506,N_29120,N_29974);
xnor UO_2507 (O_2507,N_29196,N_29862);
xor UO_2508 (O_2508,N_29598,N_29301);
nor UO_2509 (O_2509,N_29904,N_29268);
or UO_2510 (O_2510,N_29394,N_29073);
nand UO_2511 (O_2511,N_29674,N_29047);
or UO_2512 (O_2512,N_29149,N_29017);
or UO_2513 (O_2513,N_29204,N_29763);
xor UO_2514 (O_2514,N_29237,N_29688);
xnor UO_2515 (O_2515,N_29653,N_29152);
xnor UO_2516 (O_2516,N_29147,N_29059);
nor UO_2517 (O_2517,N_29231,N_29320);
or UO_2518 (O_2518,N_29598,N_29139);
nor UO_2519 (O_2519,N_29358,N_29904);
and UO_2520 (O_2520,N_29875,N_29104);
or UO_2521 (O_2521,N_29581,N_29227);
and UO_2522 (O_2522,N_29247,N_29168);
xnor UO_2523 (O_2523,N_29346,N_29747);
xnor UO_2524 (O_2524,N_29191,N_29190);
nor UO_2525 (O_2525,N_29462,N_29962);
xor UO_2526 (O_2526,N_29459,N_29378);
xnor UO_2527 (O_2527,N_29680,N_29250);
xnor UO_2528 (O_2528,N_29992,N_29670);
nor UO_2529 (O_2529,N_29748,N_29918);
or UO_2530 (O_2530,N_29692,N_29236);
and UO_2531 (O_2531,N_29310,N_29270);
xor UO_2532 (O_2532,N_29248,N_29861);
and UO_2533 (O_2533,N_29040,N_29044);
or UO_2534 (O_2534,N_29353,N_29809);
nand UO_2535 (O_2535,N_29637,N_29554);
nor UO_2536 (O_2536,N_29244,N_29043);
or UO_2537 (O_2537,N_29651,N_29545);
or UO_2538 (O_2538,N_29412,N_29377);
and UO_2539 (O_2539,N_29534,N_29468);
and UO_2540 (O_2540,N_29194,N_29878);
xor UO_2541 (O_2541,N_29227,N_29605);
nand UO_2542 (O_2542,N_29542,N_29969);
nand UO_2543 (O_2543,N_29715,N_29539);
nand UO_2544 (O_2544,N_29496,N_29380);
and UO_2545 (O_2545,N_29681,N_29267);
nand UO_2546 (O_2546,N_29355,N_29265);
and UO_2547 (O_2547,N_29260,N_29850);
xor UO_2548 (O_2548,N_29838,N_29677);
nor UO_2549 (O_2549,N_29092,N_29900);
or UO_2550 (O_2550,N_29219,N_29437);
nand UO_2551 (O_2551,N_29976,N_29744);
or UO_2552 (O_2552,N_29344,N_29082);
and UO_2553 (O_2553,N_29791,N_29956);
xnor UO_2554 (O_2554,N_29100,N_29113);
and UO_2555 (O_2555,N_29307,N_29478);
or UO_2556 (O_2556,N_29442,N_29330);
or UO_2557 (O_2557,N_29215,N_29904);
nand UO_2558 (O_2558,N_29672,N_29620);
or UO_2559 (O_2559,N_29292,N_29108);
nor UO_2560 (O_2560,N_29195,N_29439);
nor UO_2561 (O_2561,N_29739,N_29718);
nor UO_2562 (O_2562,N_29470,N_29632);
xnor UO_2563 (O_2563,N_29507,N_29568);
nor UO_2564 (O_2564,N_29564,N_29882);
xnor UO_2565 (O_2565,N_29771,N_29567);
or UO_2566 (O_2566,N_29955,N_29821);
and UO_2567 (O_2567,N_29035,N_29880);
or UO_2568 (O_2568,N_29463,N_29722);
and UO_2569 (O_2569,N_29662,N_29794);
xnor UO_2570 (O_2570,N_29000,N_29323);
or UO_2571 (O_2571,N_29046,N_29137);
xnor UO_2572 (O_2572,N_29743,N_29447);
xor UO_2573 (O_2573,N_29035,N_29233);
or UO_2574 (O_2574,N_29977,N_29019);
nor UO_2575 (O_2575,N_29092,N_29280);
nand UO_2576 (O_2576,N_29069,N_29066);
nand UO_2577 (O_2577,N_29771,N_29605);
xnor UO_2578 (O_2578,N_29985,N_29813);
and UO_2579 (O_2579,N_29668,N_29957);
xor UO_2580 (O_2580,N_29689,N_29734);
nand UO_2581 (O_2581,N_29150,N_29177);
and UO_2582 (O_2582,N_29814,N_29518);
or UO_2583 (O_2583,N_29124,N_29438);
and UO_2584 (O_2584,N_29622,N_29495);
and UO_2585 (O_2585,N_29337,N_29890);
xnor UO_2586 (O_2586,N_29637,N_29614);
xnor UO_2587 (O_2587,N_29292,N_29791);
and UO_2588 (O_2588,N_29654,N_29010);
nor UO_2589 (O_2589,N_29118,N_29781);
nand UO_2590 (O_2590,N_29210,N_29445);
or UO_2591 (O_2591,N_29226,N_29838);
xor UO_2592 (O_2592,N_29582,N_29857);
nor UO_2593 (O_2593,N_29893,N_29235);
nand UO_2594 (O_2594,N_29374,N_29305);
or UO_2595 (O_2595,N_29514,N_29171);
and UO_2596 (O_2596,N_29939,N_29170);
and UO_2597 (O_2597,N_29217,N_29152);
and UO_2598 (O_2598,N_29862,N_29636);
nand UO_2599 (O_2599,N_29383,N_29946);
nand UO_2600 (O_2600,N_29369,N_29749);
and UO_2601 (O_2601,N_29667,N_29453);
or UO_2602 (O_2602,N_29877,N_29288);
nand UO_2603 (O_2603,N_29018,N_29648);
nor UO_2604 (O_2604,N_29201,N_29360);
nor UO_2605 (O_2605,N_29847,N_29670);
or UO_2606 (O_2606,N_29247,N_29187);
or UO_2607 (O_2607,N_29086,N_29860);
and UO_2608 (O_2608,N_29220,N_29306);
nor UO_2609 (O_2609,N_29788,N_29060);
and UO_2610 (O_2610,N_29703,N_29658);
and UO_2611 (O_2611,N_29453,N_29939);
xor UO_2612 (O_2612,N_29131,N_29129);
xnor UO_2613 (O_2613,N_29395,N_29516);
and UO_2614 (O_2614,N_29987,N_29479);
xnor UO_2615 (O_2615,N_29716,N_29222);
xor UO_2616 (O_2616,N_29185,N_29427);
and UO_2617 (O_2617,N_29131,N_29779);
nand UO_2618 (O_2618,N_29575,N_29715);
and UO_2619 (O_2619,N_29346,N_29529);
nor UO_2620 (O_2620,N_29432,N_29740);
nor UO_2621 (O_2621,N_29297,N_29825);
nand UO_2622 (O_2622,N_29964,N_29489);
nand UO_2623 (O_2623,N_29782,N_29401);
nand UO_2624 (O_2624,N_29573,N_29682);
nor UO_2625 (O_2625,N_29640,N_29867);
and UO_2626 (O_2626,N_29632,N_29000);
and UO_2627 (O_2627,N_29487,N_29906);
nand UO_2628 (O_2628,N_29485,N_29208);
xnor UO_2629 (O_2629,N_29405,N_29012);
nor UO_2630 (O_2630,N_29976,N_29106);
nor UO_2631 (O_2631,N_29577,N_29780);
nand UO_2632 (O_2632,N_29279,N_29154);
nand UO_2633 (O_2633,N_29375,N_29992);
nor UO_2634 (O_2634,N_29689,N_29655);
or UO_2635 (O_2635,N_29777,N_29489);
and UO_2636 (O_2636,N_29055,N_29199);
xor UO_2637 (O_2637,N_29994,N_29629);
and UO_2638 (O_2638,N_29550,N_29075);
and UO_2639 (O_2639,N_29398,N_29985);
nor UO_2640 (O_2640,N_29795,N_29310);
or UO_2641 (O_2641,N_29064,N_29750);
nor UO_2642 (O_2642,N_29288,N_29093);
nor UO_2643 (O_2643,N_29263,N_29007);
nand UO_2644 (O_2644,N_29703,N_29934);
and UO_2645 (O_2645,N_29727,N_29243);
and UO_2646 (O_2646,N_29901,N_29917);
and UO_2647 (O_2647,N_29557,N_29380);
nand UO_2648 (O_2648,N_29853,N_29220);
xnor UO_2649 (O_2649,N_29300,N_29093);
and UO_2650 (O_2650,N_29580,N_29157);
and UO_2651 (O_2651,N_29237,N_29455);
nand UO_2652 (O_2652,N_29851,N_29281);
nand UO_2653 (O_2653,N_29030,N_29681);
and UO_2654 (O_2654,N_29112,N_29181);
nand UO_2655 (O_2655,N_29783,N_29889);
and UO_2656 (O_2656,N_29207,N_29511);
xnor UO_2657 (O_2657,N_29607,N_29058);
and UO_2658 (O_2658,N_29385,N_29167);
nor UO_2659 (O_2659,N_29844,N_29897);
nor UO_2660 (O_2660,N_29075,N_29980);
and UO_2661 (O_2661,N_29855,N_29548);
xnor UO_2662 (O_2662,N_29652,N_29167);
or UO_2663 (O_2663,N_29075,N_29524);
nand UO_2664 (O_2664,N_29993,N_29402);
xnor UO_2665 (O_2665,N_29671,N_29131);
and UO_2666 (O_2666,N_29461,N_29690);
xor UO_2667 (O_2667,N_29483,N_29503);
nand UO_2668 (O_2668,N_29925,N_29372);
xor UO_2669 (O_2669,N_29873,N_29721);
xor UO_2670 (O_2670,N_29646,N_29153);
nand UO_2671 (O_2671,N_29850,N_29740);
xnor UO_2672 (O_2672,N_29403,N_29949);
and UO_2673 (O_2673,N_29245,N_29394);
and UO_2674 (O_2674,N_29771,N_29557);
and UO_2675 (O_2675,N_29065,N_29497);
and UO_2676 (O_2676,N_29212,N_29123);
or UO_2677 (O_2677,N_29402,N_29570);
xnor UO_2678 (O_2678,N_29068,N_29942);
and UO_2679 (O_2679,N_29623,N_29390);
xor UO_2680 (O_2680,N_29567,N_29187);
and UO_2681 (O_2681,N_29456,N_29287);
and UO_2682 (O_2682,N_29837,N_29881);
nand UO_2683 (O_2683,N_29043,N_29057);
and UO_2684 (O_2684,N_29800,N_29447);
nand UO_2685 (O_2685,N_29220,N_29487);
and UO_2686 (O_2686,N_29666,N_29183);
nor UO_2687 (O_2687,N_29927,N_29143);
nor UO_2688 (O_2688,N_29132,N_29883);
nor UO_2689 (O_2689,N_29301,N_29178);
nor UO_2690 (O_2690,N_29601,N_29854);
and UO_2691 (O_2691,N_29869,N_29993);
xnor UO_2692 (O_2692,N_29856,N_29304);
nand UO_2693 (O_2693,N_29130,N_29959);
and UO_2694 (O_2694,N_29593,N_29269);
nor UO_2695 (O_2695,N_29132,N_29689);
and UO_2696 (O_2696,N_29752,N_29273);
nor UO_2697 (O_2697,N_29932,N_29219);
or UO_2698 (O_2698,N_29714,N_29468);
nor UO_2699 (O_2699,N_29925,N_29537);
nor UO_2700 (O_2700,N_29582,N_29851);
xnor UO_2701 (O_2701,N_29456,N_29492);
and UO_2702 (O_2702,N_29096,N_29106);
and UO_2703 (O_2703,N_29929,N_29820);
and UO_2704 (O_2704,N_29695,N_29064);
or UO_2705 (O_2705,N_29789,N_29848);
nor UO_2706 (O_2706,N_29684,N_29608);
or UO_2707 (O_2707,N_29180,N_29102);
or UO_2708 (O_2708,N_29368,N_29887);
or UO_2709 (O_2709,N_29783,N_29292);
xnor UO_2710 (O_2710,N_29440,N_29697);
or UO_2711 (O_2711,N_29630,N_29642);
nor UO_2712 (O_2712,N_29764,N_29418);
or UO_2713 (O_2713,N_29099,N_29839);
or UO_2714 (O_2714,N_29003,N_29435);
or UO_2715 (O_2715,N_29870,N_29631);
and UO_2716 (O_2716,N_29552,N_29570);
or UO_2717 (O_2717,N_29516,N_29323);
nand UO_2718 (O_2718,N_29346,N_29398);
nor UO_2719 (O_2719,N_29182,N_29578);
nand UO_2720 (O_2720,N_29517,N_29891);
xnor UO_2721 (O_2721,N_29584,N_29497);
or UO_2722 (O_2722,N_29279,N_29945);
xnor UO_2723 (O_2723,N_29366,N_29788);
and UO_2724 (O_2724,N_29394,N_29270);
xor UO_2725 (O_2725,N_29152,N_29817);
nor UO_2726 (O_2726,N_29081,N_29984);
and UO_2727 (O_2727,N_29313,N_29857);
xnor UO_2728 (O_2728,N_29725,N_29698);
xnor UO_2729 (O_2729,N_29708,N_29472);
and UO_2730 (O_2730,N_29093,N_29255);
nor UO_2731 (O_2731,N_29403,N_29470);
xor UO_2732 (O_2732,N_29785,N_29373);
or UO_2733 (O_2733,N_29076,N_29575);
and UO_2734 (O_2734,N_29264,N_29588);
xnor UO_2735 (O_2735,N_29790,N_29279);
nand UO_2736 (O_2736,N_29672,N_29105);
xnor UO_2737 (O_2737,N_29497,N_29233);
and UO_2738 (O_2738,N_29506,N_29560);
nand UO_2739 (O_2739,N_29605,N_29442);
nor UO_2740 (O_2740,N_29270,N_29729);
or UO_2741 (O_2741,N_29829,N_29156);
or UO_2742 (O_2742,N_29496,N_29460);
or UO_2743 (O_2743,N_29654,N_29792);
nand UO_2744 (O_2744,N_29387,N_29116);
nand UO_2745 (O_2745,N_29158,N_29597);
or UO_2746 (O_2746,N_29856,N_29834);
nor UO_2747 (O_2747,N_29843,N_29716);
and UO_2748 (O_2748,N_29551,N_29501);
nand UO_2749 (O_2749,N_29765,N_29679);
nand UO_2750 (O_2750,N_29051,N_29230);
or UO_2751 (O_2751,N_29016,N_29407);
nand UO_2752 (O_2752,N_29698,N_29346);
xnor UO_2753 (O_2753,N_29213,N_29299);
or UO_2754 (O_2754,N_29740,N_29723);
nand UO_2755 (O_2755,N_29409,N_29650);
xnor UO_2756 (O_2756,N_29060,N_29337);
or UO_2757 (O_2757,N_29318,N_29247);
xnor UO_2758 (O_2758,N_29276,N_29835);
and UO_2759 (O_2759,N_29369,N_29916);
nor UO_2760 (O_2760,N_29441,N_29795);
xnor UO_2761 (O_2761,N_29806,N_29720);
and UO_2762 (O_2762,N_29005,N_29373);
xor UO_2763 (O_2763,N_29416,N_29651);
and UO_2764 (O_2764,N_29858,N_29417);
nor UO_2765 (O_2765,N_29894,N_29181);
and UO_2766 (O_2766,N_29330,N_29983);
or UO_2767 (O_2767,N_29933,N_29180);
xnor UO_2768 (O_2768,N_29027,N_29181);
or UO_2769 (O_2769,N_29815,N_29355);
nor UO_2770 (O_2770,N_29894,N_29546);
nand UO_2771 (O_2771,N_29371,N_29215);
nor UO_2772 (O_2772,N_29321,N_29862);
nand UO_2773 (O_2773,N_29356,N_29415);
or UO_2774 (O_2774,N_29711,N_29622);
nand UO_2775 (O_2775,N_29872,N_29468);
nand UO_2776 (O_2776,N_29362,N_29156);
nand UO_2777 (O_2777,N_29923,N_29153);
and UO_2778 (O_2778,N_29614,N_29613);
nand UO_2779 (O_2779,N_29649,N_29315);
xnor UO_2780 (O_2780,N_29790,N_29761);
nor UO_2781 (O_2781,N_29260,N_29986);
and UO_2782 (O_2782,N_29047,N_29715);
xnor UO_2783 (O_2783,N_29714,N_29705);
or UO_2784 (O_2784,N_29279,N_29188);
or UO_2785 (O_2785,N_29129,N_29999);
nor UO_2786 (O_2786,N_29036,N_29838);
nand UO_2787 (O_2787,N_29816,N_29709);
or UO_2788 (O_2788,N_29296,N_29311);
nor UO_2789 (O_2789,N_29140,N_29252);
xnor UO_2790 (O_2790,N_29063,N_29986);
nand UO_2791 (O_2791,N_29697,N_29710);
nand UO_2792 (O_2792,N_29571,N_29313);
nor UO_2793 (O_2793,N_29589,N_29018);
and UO_2794 (O_2794,N_29253,N_29652);
nand UO_2795 (O_2795,N_29528,N_29717);
nor UO_2796 (O_2796,N_29120,N_29798);
nor UO_2797 (O_2797,N_29258,N_29217);
xor UO_2798 (O_2798,N_29137,N_29386);
and UO_2799 (O_2799,N_29340,N_29681);
xnor UO_2800 (O_2800,N_29686,N_29012);
or UO_2801 (O_2801,N_29706,N_29906);
nand UO_2802 (O_2802,N_29801,N_29117);
nor UO_2803 (O_2803,N_29662,N_29371);
nand UO_2804 (O_2804,N_29221,N_29011);
xor UO_2805 (O_2805,N_29460,N_29163);
nand UO_2806 (O_2806,N_29092,N_29741);
nand UO_2807 (O_2807,N_29345,N_29291);
or UO_2808 (O_2808,N_29719,N_29462);
nand UO_2809 (O_2809,N_29008,N_29506);
or UO_2810 (O_2810,N_29108,N_29678);
nand UO_2811 (O_2811,N_29744,N_29105);
nor UO_2812 (O_2812,N_29657,N_29986);
or UO_2813 (O_2813,N_29712,N_29296);
and UO_2814 (O_2814,N_29394,N_29763);
and UO_2815 (O_2815,N_29484,N_29662);
xor UO_2816 (O_2816,N_29527,N_29907);
and UO_2817 (O_2817,N_29740,N_29292);
or UO_2818 (O_2818,N_29042,N_29346);
nor UO_2819 (O_2819,N_29892,N_29380);
or UO_2820 (O_2820,N_29869,N_29717);
xnor UO_2821 (O_2821,N_29148,N_29761);
and UO_2822 (O_2822,N_29955,N_29868);
or UO_2823 (O_2823,N_29302,N_29082);
and UO_2824 (O_2824,N_29153,N_29106);
xnor UO_2825 (O_2825,N_29066,N_29683);
and UO_2826 (O_2826,N_29827,N_29915);
nor UO_2827 (O_2827,N_29337,N_29551);
or UO_2828 (O_2828,N_29976,N_29046);
xor UO_2829 (O_2829,N_29993,N_29291);
or UO_2830 (O_2830,N_29863,N_29855);
nor UO_2831 (O_2831,N_29460,N_29770);
xor UO_2832 (O_2832,N_29142,N_29454);
or UO_2833 (O_2833,N_29973,N_29959);
nor UO_2834 (O_2834,N_29884,N_29850);
or UO_2835 (O_2835,N_29684,N_29855);
and UO_2836 (O_2836,N_29486,N_29647);
nor UO_2837 (O_2837,N_29392,N_29196);
xor UO_2838 (O_2838,N_29488,N_29319);
or UO_2839 (O_2839,N_29517,N_29334);
xor UO_2840 (O_2840,N_29707,N_29062);
nand UO_2841 (O_2841,N_29804,N_29339);
and UO_2842 (O_2842,N_29918,N_29782);
nor UO_2843 (O_2843,N_29051,N_29689);
or UO_2844 (O_2844,N_29060,N_29486);
and UO_2845 (O_2845,N_29493,N_29708);
or UO_2846 (O_2846,N_29107,N_29690);
or UO_2847 (O_2847,N_29312,N_29702);
nand UO_2848 (O_2848,N_29520,N_29032);
and UO_2849 (O_2849,N_29544,N_29476);
nor UO_2850 (O_2850,N_29414,N_29182);
and UO_2851 (O_2851,N_29614,N_29057);
nor UO_2852 (O_2852,N_29610,N_29624);
and UO_2853 (O_2853,N_29018,N_29365);
and UO_2854 (O_2854,N_29936,N_29140);
or UO_2855 (O_2855,N_29642,N_29358);
nor UO_2856 (O_2856,N_29534,N_29072);
nand UO_2857 (O_2857,N_29092,N_29072);
nor UO_2858 (O_2858,N_29046,N_29391);
or UO_2859 (O_2859,N_29641,N_29210);
and UO_2860 (O_2860,N_29947,N_29247);
and UO_2861 (O_2861,N_29937,N_29088);
and UO_2862 (O_2862,N_29944,N_29163);
and UO_2863 (O_2863,N_29383,N_29039);
nor UO_2864 (O_2864,N_29904,N_29621);
xor UO_2865 (O_2865,N_29353,N_29460);
or UO_2866 (O_2866,N_29894,N_29521);
xnor UO_2867 (O_2867,N_29124,N_29885);
nand UO_2868 (O_2868,N_29488,N_29434);
and UO_2869 (O_2869,N_29664,N_29120);
or UO_2870 (O_2870,N_29605,N_29180);
nor UO_2871 (O_2871,N_29878,N_29131);
nor UO_2872 (O_2872,N_29850,N_29101);
nand UO_2873 (O_2873,N_29441,N_29405);
or UO_2874 (O_2874,N_29522,N_29973);
or UO_2875 (O_2875,N_29383,N_29491);
and UO_2876 (O_2876,N_29508,N_29244);
xnor UO_2877 (O_2877,N_29664,N_29824);
xor UO_2878 (O_2878,N_29521,N_29205);
or UO_2879 (O_2879,N_29853,N_29049);
xnor UO_2880 (O_2880,N_29846,N_29834);
nor UO_2881 (O_2881,N_29058,N_29907);
nand UO_2882 (O_2882,N_29529,N_29820);
xnor UO_2883 (O_2883,N_29986,N_29112);
and UO_2884 (O_2884,N_29706,N_29314);
nor UO_2885 (O_2885,N_29799,N_29061);
nand UO_2886 (O_2886,N_29525,N_29592);
xnor UO_2887 (O_2887,N_29737,N_29660);
nand UO_2888 (O_2888,N_29210,N_29877);
nor UO_2889 (O_2889,N_29847,N_29085);
or UO_2890 (O_2890,N_29716,N_29345);
and UO_2891 (O_2891,N_29631,N_29172);
and UO_2892 (O_2892,N_29991,N_29516);
xor UO_2893 (O_2893,N_29429,N_29805);
xor UO_2894 (O_2894,N_29993,N_29801);
nand UO_2895 (O_2895,N_29358,N_29958);
nor UO_2896 (O_2896,N_29291,N_29507);
and UO_2897 (O_2897,N_29383,N_29871);
and UO_2898 (O_2898,N_29770,N_29327);
and UO_2899 (O_2899,N_29258,N_29681);
xnor UO_2900 (O_2900,N_29839,N_29487);
and UO_2901 (O_2901,N_29484,N_29515);
xnor UO_2902 (O_2902,N_29911,N_29673);
nor UO_2903 (O_2903,N_29169,N_29625);
nand UO_2904 (O_2904,N_29981,N_29433);
nor UO_2905 (O_2905,N_29107,N_29850);
nand UO_2906 (O_2906,N_29515,N_29351);
nand UO_2907 (O_2907,N_29621,N_29477);
xor UO_2908 (O_2908,N_29895,N_29530);
xnor UO_2909 (O_2909,N_29702,N_29169);
or UO_2910 (O_2910,N_29500,N_29132);
nor UO_2911 (O_2911,N_29944,N_29234);
and UO_2912 (O_2912,N_29859,N_29159);
xnor UO_2913 (O_2913,N_29937,N_29128);
nor UO_2914 (O_2914,N_29961,N_29666);
and UO_2915 (O_2915,N_29601,N_29389);
nand UO_2916 (O_2916,N_29668,N_29298);
or UO_2917 (O_2917,N_29753,N_29186);
and UO_2918 (O_2918,N_29354,N_29436);
nor UO_2919 (O_2919,N_29959,N_29674);
nand UO_2920 (O_2920,N_29008,N_29273);
nand UO_2921 (O_2921,N_29399,N_29597);
nand UO_2922 (O_2922,N_29166,N_29360);
nand UO_2923 (O_2923,N_29116,N_29777);
or UO_2924 (O_2924,N_29361,N_29501);
or UO_2925 (O_2925,N_29029,N_29310);
xor UO_2926 (O_2926,N_29660,N_29281);
and UO_2927 (O_2927,N_29268,N_29054);
and UO_2928 (O_2928,N_29545,N_29232);
nor UO_2929 (O_2929,N_29383,N_29002);
and UO_2930 (O_2930,N_29860,N_29472);
nor UO_2931 (O_2931,N_29763,N_29412);
and UO_2932 (O_2932,N_29873,N_29445);
and UO_2933 (O_2933,N_29340,N_29433);
nand UO_2934 (O_2934,N_29147,N_29291);
or UO_2935 (O_2935,N_29403,N_29878);
or UO_2936 (O_2936,N_29783,N_29689);
nand UO_2937 (O_2937,N_29907,N_29852);
or UO_2938 (O_2938,N_29837,N_29672);
nand UO_2939 (O_2939,N_29940,N_29144);
and UO_2940 (O_2940,N_29058,N_29318);
and UO_2941 (O_2941,N_29049,N_29569);
xnor UO_2942 (O_2942,N_29537,N_29151);
nand UO_2943 (O_2943,N_29196,N_29320);
xor UO_2944 (O_2944,N_29231,N_29465);
or UO_2945 (O_2945,N_29064,N_29094);
xor UO_2946 (O_2946,N_29481,N_29384);
or UO_2947 (O_2947,N_29755,N_29785);
nand UO_2948 (O_2948,N_29240,N_29064);
or UO_2949 (O_2949,N_29861,N_29958);
or UO_2950 (O_2950,N_29225,N_29526);
nand UO_2951 (O_2951,N_29691,N_29298);
nand UO_2952 (O_2952,N_29095,N_29748);
nand UO_2953 (O_2953,N_29972,N_29288);
xor UO_2954 (O_2954,N_29642,N_29076);
or UO_2955 (O_2955,N_29344,N_29711);
xor UO_2956 (O_2956,N_29409,N_29402);
nor UO_2957 (O_2957,N_29083,N_29851);
or UO_2958 (O_2958,N_29345,N_29230);
xor UO_2959 (O_2959,N_29034,N_29290);
nor UO_2960 (O_2960,N_29840,N_29141);
or UO_2961 (O_2961,N_29271,N_29317);
or UO_2962 (O_2962,N_29454,N_29988);
nor UO_2963 (O_2963,N_29089,N_29385);
and UO_2964 (O_2964,N_29241,N_29361);
xor UO_2965 (O_2965,N_29374,N_29833);
or UO_2966 (O_2966,N_29694,N_29060);
nand UO_2967 (O_2967,N_29399,N_29098);
and UO_2968 (O_2968,N_29021,N_29621);
nand UO_2969 (O_2969,N_29533,N_29815);
and UO_2970 (O_2970,N_29491,N_29226);
and UO_2971 (O_2971,N_29110,N_29864);
xor UO_2972 (O_2972,N_29374,N_29581);
and UO_2973 (O_2973,N_29047,N_29379);
xnor UO_2974 (O_2974,N_29944,N_29135);
nand UO_2975 (O_2975,N_29586,N_29696);
or UO_2976 (O_2976,N_29805,N_29837);
xor UO_2977 (O_2977,N_29870,N_29766);
nor UO_2978 (O_2978,N_29779,N_29240);
nand UO_2979 (O_2979,N_29485,N_29259);
nor UO_2980 (O_2980,N_29517,N_29152);
nor UO_2981 (O_2981,N_29923,N_29632);
or UO_2982 (O_2982,N_29076,N_29602);
or UO_2983 (O_2983,N_29532,N_29416);
or UO_2984 (O_2984,N_29680,N_29715);
nor UO_2985 (O_2985,N_29919,N_29750);
nand UO_2986 (O_2986,N_29166,N_29375);
or UO_2987 (O_2987,N_29354,N_29697);
nand UO_2988 (O_2988,N_29137,N_29050);
and UO_2989 (O_2989,N_29758,N_29591);
nor UO_2990 (O_2990,N_29199,N_29843);
nand UO_2991 (O_2991,N_29008,N_29214);
nor UO_2992 (O_2992,N_29979,N_29023);
nand UO_2993 (O_2993,N_29818,N_29305);
xor UO_2994 (O_2994,N_29428,N_29432);
xnor UO_2995 (O_2995,N_29431,N_29038);
or UO_2996 (O_2996,N_29758,N_29434);
nor UO_2997 (O_2997,N_29435,N_29838);
nor UO_2998 (O_2998,N_29144,N_29910);
nor UO_2999 (O_2999,N_29551,N_29302);
or UO_3000 (O_3000,N_29338,N_29385);
and UO_3001 (O_3001,N_29860,N_29800);
or UO_3002 (O_3002,N_29830,N_29051);
nor UO_3003 (O_3003,N_29014,N_29296);
nor UO_3004 (O_3004,N_29367,N_29030);
and UO_3005 (O_3005,N_29575,N_29027);
xnor UO_3006 (O_3006,N_29056,N_29921);
nor UO_3007 (O_3007,N_29605,N_29283);
nand UO_3008 (O_3008,N_29654,N_29477);
or UO_3009 (O_3009,N_29314,N_29878);
nor UO_3010 (O_3010,N_29838,N_29561);
nand UO_3011 (O_3011,N_29751,N_29959);
nor UO_3012 (O_3012,N_29965,N_29722);
or UO_3013 (O_3013,N_29814,N_29198);
nor UO_3014 (O_3014,N_29370,N_29483);
or UO_3015 (O_3015,N_29545,N_29368);
xnor UO_3016 (O_3016,N_29389,N_29326);
or UO_3017 (O_3017,N_29271,N_29087);
nor UO_3018 (O_3018,N_29131,N_29566);
nand UO_3019 (O_3019,N_29040,N_29798);
nor UO_3020 (O_3020,N_29526,N_29953);
nand UO_3021 (O_3021,N_29670,N_29225);
or UO_3022 (O_3022,N_29185,N_29128);
or UO_3023 (O_3023,N_29043,N_29265);
or UO_3024 (O_3024,N_29963,N_29918);
xnor UO_3025 (O_3025,N_29798,N_29293);
and UO_3026 (O_3026,N_29348,N_29742);
nor UO_3027 (O_3027,N_29768,N_29482);
xor UO_3028 (O_3028,N_29401,N_29857);
nand UO_3029 (O_3029,N_29435,N_29811);
or UO_3030 (O_3030,N_29586,N_29957);
or UO_3031 (O_3031,N_29645,N_29061);
or UO_3032 (O_3032,N_29872,N_29579);
and UO_3033 (O_3033,N_29936,N_29830);
nand UO_3034 (O_3034,N_29285,N_29786);
xnor UO_3035 (O_3035,N_29417,N_29303);
xnor UO_3036 (O_3036,N_29511,N_29637);
and UO_3037 (O_3037,N_29063,N_29255);
nor UO_3038 (O_3038,N_29546,N_29390);
xor UO_3039 (O_3039,N_29050,N_29914);
xnor UO_3040 (O_3040,N_29270,N_29940);
xnor UO_3041 (O_3041,N_29085,N_29747);
nand UO_3042 (O_3042,N_29178,N_29155);
nor UO_3043 (O_3043,N_29179,N_29701);
or UO_3044 (O_3044,N_29872,N_29149);
and UO_3045 (O_3045,N_29666,N_29185);
xor UO_3046 (O_3046,N_29728,N_29994);
nor UO_3047 (O_3047,N_29675,N_29076);
xor UO_3048 (O_3048,N_29350,N_29454);
xnor UO_3049 (O_3049,N_29813,N_29236);
nand UO_3050 (O_3050,N_29828,N_29846);
xor UO_3051 (O_3051,N_29236,N_29901);
or UO_3052 (O_3052,N_29033,N_29736);
nand UO_3053 (O_3053,N_29895,N_29872);
xnor UO_3054 (O_3054,N_29577,N_29356);
xor UO_3055 (O_3055,N_29235,N_29193);
nor UO_3056 (O_3056,N_29776,N_29254);
or UO_3057 (O_3057,N_29896,N_29759);
nor UO_3058 (O_3058,N_29101,N_29218);
or UO_3059 (O_3059,N_29175,N_29430);
xnor UO_3060 (O_3060,N_29191,N_29983);
nor UO_3061 (O_3061,N_29586,N_29418);
xnor UO_3062 (O_3062,N_29023,N_29759);
xnor UO_3063 (O_3063,N_29456,N_29922);
or UO_3064 (O_3064,N_29901,N_29097);
nand UO_3065 (O_3065,N_29033,N_29172);
and UO_3066 (O_3066,N_29893,N_29866);
and UO_3067 (O_3067,N_29935,N_29641);
or UO_3068 (O_3068,N_29124,N_29087);
xnor UO_3069 (O_3069,N_29069,N_29097);
or UO_3070 (O_3070,N_29649,N_29707);
or UO_3071 (O_3071,N_29124,N_29623);
nor UO_3072 (O_3072,N_29557,N_29631);
and UO_3073 (O_3073,N_29324,N_29755);
and UO_3074 (O_3074,N_29447,N_29536);
nor UO_3075 (O_3075,N_29906,N_29512);
or UO_3076 (O_3076,N_29789,N_29712);
nand UO_3077 (O_3077,N_29587,N_29132);
or UO_3078 (O_3078,N_29982,N_29780);
nor UO_3079 (O_3079,N_29028,N_29868);
nor UO_3080 (O_3080,N_29133,N_29529);
or UO_3081 (O_3081,N_29917,N_29347);
xor UO_3082 (O_3082,N_29295,N_29788);
xor UO_3083 (O_3083,N_29021,N_29265);
nand UO_3084 (O_3084,N_29509,N_29705);
or UO_3085 (O_3085,N_29381,N_29039);
nor UO_3086 (O_3086,N_29324,N_29428);
or UO_3087 (O_3087,N_29961,N_29867);
nor UO_3088 (O_3088,N_29667,N_29876);
nor UO_3089 (O_3089,N_29714,N_29976);
and UO_3090 (O_3090,N_29138,N_29523);
or UO_3091 (O_3091,N_29134,N_29654);
or UO_3092 (O_3092,N_29509,N_29201);
or UO_3093 (O_3093,N_29562,N_29454);
nand UO_3094 (O_3094,N_29786,N_29479);
xnor UO_3095 (O_3095,N_29086,N_29730);
or UO_3096 (O_3096,N_29932,N_29677);
and UO_3097 (O_3097,N_29203,N_29725);
or UO_3098 (O_3098,N_29494,N_29970);
xor UO_3099 (O_3099,N_29002,N_29141);
and UO_3100 (O_3100,N_29156,N_29964);
xor UO_3101 (O_3101,N_29262,N_29385);
and UO_3102 (O_3102,N_29527,N_29923);
and UO_3103 (O_3103,N_29313,N_29533);
or UO_3104 (O_3104,N_29099,N_29258);
xor UO_3105 (O_3105,N_29501,N_29893);
xor UO_3106 (O_3106,N_29709,N_29553);
nor UO_3107 (O_3107,N_29286,N_29535);
and UO_3108 (O_3108,N_29087,N_29770);
or UO_3109 (O_3109,N_29468,N_29575);
and UO_3110 (O_3110,N_29738,N_29538);
or UO_3111 (O_3111,N_29572,N_29042);
or UO_3112 (O_3112,N_29251,N_29864);
or UO_3113 (O_3113,N_29472,N_29811);
and UO_3114 (O_3114,N_29664,N_29346);
nand UO_3115 (O_3115,N_29452,N_29693);
nand UO_3116 (O_3116,N_29394,N_29757);
or UO_3117 (O_3117,N_29662,N_29077);
nand UO_3118 (O_3118,N_29804,N_29551);
xor UO_3119 (O_3119,N_29434,N_29024);
or UO_3120 (O_3120,N_29219,N_29739);
or UO_3121 (O_3121,N_29828,N_29169);
xor UO_3122 (O_3122,N_29708,N_29125);
nand UO_3123 (O_3123,N_29201,N_29982);
or UO_3124 (O_3124,N_29181,N_29660);
or UO_3125 (O_3125,N_29071,N_29776);
nand UO_3126 (O_3126,N_29697,N_29888);
and UO_3127 (O_3127,N_29597,N_29241);
and UO_3128 (O_3128,N_29919,N_29361);
xnor UO_3129 (O_3129,N_29161,N_29225);
or UO_3130 (O_3130,N_29639,N_29184);
and UO_3131 (O_3131,N_29237,N_29888);
or UO_3132 (O_3132,N_29649,N_29528);
nor UO_3133 (O_3133,N_29503,N_29877);
and UO_3134 (O_3134,N_29971,N_29806);
or UO_3135 (O_3135,N_29780,N_29887);
or UO_3136 (O_3136,N_29099,N_29792);
nand UO_3137 (O_3137,N_29200,N_29382);
xnor UO_3138 (O_3138,N_29127,N_29875);
xnor UO_3139 (O_3139,N_29197,N_29749);
nand UO_3140 (O_3140,N_29846,N_29322);
nand UO_3141 (O_3141,N_29633,N_29340);
and UO_3142 (O_3142,N_29645,N_29799);
xor UO_3143 (O_3143,N_29602,N_29530);
xnor UO_3144 (O_3144,N_29531,N_29580);
and UO_3145 (O_3145,N_29911,N_29038);
or UO_3146 (O_3146,N_29163,N_29605);
or UO_3147 (O_3147,N_29609,N_29824);
or UO_3148 (O_3148,N_29297,N_29643);
nand UO_3149 (O_3149,N_29001,N_29581);
and UO_3150 (O_3150,N_29759,N_29159);
xnor UO_3151 (O_3151,N_29050,N_29003);
nand UO_3152 (O_3152,N_29738,N_29102);
nor UO_3153 (O_3153,N_29439,N_29008);
and UO_3154 (O_3154,N_29122,N_29966);
xnor UO_3155 (O_3155,N_29924,N_29641);
xor UO_3156 (O_3156,N_29509,N_29481);
nor UO_3157 (O_3157,N_29561,N_29078);
nor UO_3158 (O_3158,N_29902,N_29364);
nor UO_3159 (O_3159,N_29949,N_29278);
xor UO_3160 (O_3160,N_29712,N_29838);
or UO_3161 (O_3161,N_29504,N_29776);
nor UO_3162 (O_3162,N_29143,N_29443);
or UO_3163 (O_3163,N_29192,N_29404);
xor UO_3164 (O_3164,N_29228,N_29526);
and UO_3165 (O_3165,N_29174,N_29671);
nand UO_3166 (O_3166,N_29004,N_29264);
xnor UO_3167 (O_3167,N_29803,N_29628);
nor UO_3168 (O_3168,N_29318,N_29568);
xnor UO_3169 (O_3169,N_29305,N_29605);
nand UO_3170 (O_3170,N_29454,N_29030);
nand UO_3171 (O_3171,N_29315,N_29873);
nand UO_3172 (O_3172,N_29804,N_29480);
and UO_3173 (O_3173,N_29563,N_29364);
nand UO_3174 (O_3174,N_29271,N_29739);
and UO_3175 (O_3175,N_29320,N_29592);
xnor UO_3176 (O_3176,N_29949,N_29874);
and UO_3177 (O_3177,N_29519,N_29106);
nand UO_3178 (O_3178,N_29677,N_29984);
and UO_3179 (O_3179,N_29263,N_29384);
nor UO_3180 (O_3180,N_29487,N_29788);
nand UO_3181 (O_3181,N_29878,N_29172);
and UO_3182 (O_3182,N_29917,N_29131);
or UO_3183 (O_3183,N_29610,N_29506);
and UO_3184 (O_3184,N_29728,N_29359);
and UO_3185 (O_3185,N_29102,N_29843);
nor UO_3186 (O_3186,N_29173,N_29996);
nand UO_3187 (O_3187,N_29844,N_29010);
nor UO_3188 (O_3188,N_29779,N_29472);
xnor UO_3189 (O_3189,N_29327,N_29970);
nand UO_3190 (O_3190,N_29628,N_29642);
and UO_3191 (O_3191,N_29760,N_29784);
nand UO_3192 (O_3192,N_29800,N_29601);
nor UO_3193 (O_3193,N_29025,N_29193);
and UO_3194 (O_3194,N_29346,N_29107);
xor UO_3195 (O_3195,N_29834,N_29750);
nand UO_3196 (O_3196,N_29258,N_29808);
xnor UO_3197 (O_3197,N_29305,N_29342);
nor UO_3198 (O_3198,N_29798,N_29509);
nor UO_3199 (O_3199,N_29254,N_29387);
xor UO_3200 (O_3200,N_29972,N_29674);
and UO_3201 (O_3201,N_29522,N_29597);
and UO_3202 (O_3202,N_29010,N_29539);
xnor UO_3203 (O_3203,N_29344,N_29251);
nor UO_3204 (O_3204,N_29223,N_29521);
and UO_3205 (O_3205,N_29219,N_29012);
nand UO_3206 (O_3206,N_29535,N_29432);
or UO_3207 (O_3207,N_29474,N_29653);
nor UO_3208 (O_3208,N_29038,N_29019);
or UO_3209 (O_3209,N_29537,N_29662);
and UO_3210 (O_3210,N_29666,N_29145);
xnor UO_3211 (O_3211,N_29559,N_29763);
xnor UO_3212 (O_3212,N_29202,N_29348);
nand UO_3213 (O_3213,N_29388,N_29087);
or UO_3214 (O_3214,N_29819,N_29855);
or UO_3215 (O_3215,N_29382,N_29295);
and UO_3216 (O_3216,N_29479,N_29608);
xor UO_3217 (O_3217,N_29289,N_29990);
nand UO_3218 (O_3218,N_29645,N_29280);
nor UO_3219 (O_3219,N_29305,N_29496);
nor UO_3220 (O_3220,N_29703,N_29904);
or UO_3221 (O_3221,N_29009,N_29181);
and UO_3222 (O_3222,N_29722,N_29950);
and UO_3223 (O_3223,N_29144,N_29425);
nand UO_3224 (O_3224,N_29115,N_29118);
and UO_3225 (O_3225,N_29491,N_29681);
nand UO_3226 (O_3226,N_29518,N_29752);
or UO_3227 (O_3227,N_29734,N_29541);
xnor UO_3228 (O_3228,N_29001,N_29751);
nor UO_3229 (O_3229,N_29046,N_29689);
nor UO_3230 (O_3230,N_29769,N_29764);
nand UO_3231 (O_3231,N_29085,N_29756);
nand UO_3232 (O_3232,N_29318,N_29991);
nor UO_3233 (O_3233,N_29192,N_29030);
and UO_3234 (O_3234,N_29120,N_29652);
or UO_3235 (O_3235,N_29151,N_29700);
and UO_3236 (O_3236,N_29295,N_29586);
nand UO_3237 (O_3237,N_29550,N_29624);
or UO_3238 (O_3238,N_29181,N_29684);
xor UO_3239 (O_3239,N_29226,N_29404);
nor UO_3240 (O_3240,N_29466,N_29852);
xor UO_3241 (O_3241,N_29787,N_29516);
or UO_3242 (O_3242,N_29989,N_29618);
nor UO_3243 (O_3243,N_29737,N_29671);
nor UO_3244 (O_3244,N_29766,N_29637);
nor UO_3245 (O_3245,N_29279,N_29489);
nor UO_3246 (O_3246,N_29711,N_29842);
nor UO_3247 (O_3247,N_29809,N_29581);
and UO_3248 (O_3248,N_29483,N_29473);
nor UO_3249 (O_3249,N_29625,N_29825);
nand UO_3250 (O_3250,N_29012,N_29229);
xnor UO_3251 (O_3251,N_29333,N_29996);
and UO_3252 (O_3252,N_29084,N_29951);
and UO_3253 (O_3253,N_29658,N_29957);
nor UO_3254 (O_3254,N_29012,N_29713);
nor UO_3255 (O_3255,N_29981,N_29308);
nand UO_3256 (O_3256,N_29654,N_29099);
and UO_3257 (O_3257,N_29932,N_29735);
xnor UO_3258 (O_3258,N_29617,N_29355);
nor UO_3259 (O_3259,N_29036,N_29980);
or UO_3260 (O_3260,N_29192,N_29923);
nand UO_3261 (O_3261,N_29610,N_29175);
or UO_3262 (O_3262,N_29042,N_29036);
nand UO_3263 (O_3263,N_29977,N_29177);
nor UO_3264 (O_3264,N_29567,N_29555);
or UO_3265 (O_3265,N_29119,N_29048);
nand UO_3266 (O_3266,N_29784,N_29617);
or UO_3267 (O_3267,N_29176,N_29996);
and UO_3268 (O_3268,N_29989,N_29251);
or UO_3269 (O_3269,N_29728,N_29439);
or UO_3270 (O_3270,N_29638,N_29275);
and UO_3271 (O_3271,N_29657,N_29709);
and UO_3272 (O_3272,N_29045,N_29653);
nor UO_3273 (O_3273,N_29568,N_29205);
nand UO_3274 (O_3274,N_29972,N_29063);
nor UO_3275 (O_3275,N_29728,N_29216);
nor UO_3276 (O_3276,N_29231,N_29701);
xnor UO_3277 (O_3277,N_29885,N_29146);
and UO_3278 (O_3278,N_29416,N_29302);
and UO_3279 (O_3279,N_29707,N_29370);
nand UO_3280 (O_3280,N_29321,N_29515);
xor UO_3281 (O_3281,N_29263,N_29222);
xor UO_3282 (O_3282,N_29968,N_29211);
nand UO_3283 (O_3283,N_29997,N_29088);
and UO_3284 (O_3284,N_29705,N_29384);
or UO_3285 (O_3285,N_29911,N_29022);
nand UO_3286 (O_3286,N_29159,N_29172);
or UO_3287 (O_3287,N_29493,N_29065);
nor UO_3288 (O_3288,N_29905,N_29337);
and UO_3289 (O_3289,N_29727,N_29036);
and UO_3290 (O_3290,N_29702,N_29499);
nand UO_3291 (O_3291,N_29296,N_29172);
and UO_3292 (O_3292,N_29828,N_29673);
or UO_3293 (O_3293,N_29258,N_29590);
nor UO_3294 (O_3294,N_29013,N_29737);
nor UO_3295 (O_3295,N_29457,N_29035);
nand UO_3296 (O_3296,N_29111,N_29381);
or UO_3297 (O_3297,N_29359,N_29604);
nand UO_3298 (O_3298,N_29065,N_29601);
and UO_3299 (O_3299,N_29598,N_29147);
and UO_3300 (O_3300,N_29662,N_29907);
nand UO_3301 (O_3301,N_29212,N_29319);
nor UO_3302 (O_3302,N_29305,N_29528);
nor UO_3303 (O_3303,N_29174,N_29516);
or UO_3304 (O_3304,N_29139,N_29544);
nand UO_3305 (O_3305,N_29646,N_29835);
and UO_3306 (O_3306,N_29555,N_29519);
xor UO_3307 (O_3307,N_29072,N_29743);
nand UO_3308 (O_3308,N_29273,N_29569);
nand UO_3309 (O_3309,N_29629,N_29848);
or UO_3310 (O_3310,N_29838,N_29926);
nor UO_3311 (O_3311,N_29155,N_29301);
and UO_3312 (O_3312,N_29920,N_29545);
or UO_3313 (O_3313,N_29886,N_29649);
and UO_3314 (O_3314,N_29453,N_29982);
and UO_3315 (O_3315,N_29547,N_29133);
and UO_3316 (O_3316,N_29367,N_29037);
nand UO_3317 (O_3317,N_29758,N_29970);
and UO_3318 (O_3318,N_29100,N_29694);
nor UO_3319 (O_3319,N_29363,N_29620);
and UO_3320 (O_3320,N_29546,N_29371);
xnor UO_3321 (O_3321,N_29907,N_29834);
nor UO_3322 (O_3322,N_29986,N_29008);
nand UO_3323 (O_3323,N_29784,N_29180);
and UO_3324 (O_3324,N_29456,N_29766);
and UO_3325 (O_3325,N_29523,N_29727);
nand UO_3326 (O_3326,N_29757,N_29844);
and UO_3327 (O_3327,N_29853,N_29874);
and UO_3328 (O_3328,N_29680,N_29338);
xnor UO_3329 (O_3329,N_29826,N_29751);
or UO_3330 (O_3330,N_29048,N_29512);
nor UO_3331 (O_3331,N_29230,N_29849);
nor UO_3332 (O_3332,N_29619,N_29512);
nor UO_3333 (O_3333,N_29125,N_29955);
xnor UO_3334 (O_3334,N_29948,N_29321);
nand UO_3335 (O_3335,N_29816,N_29879);
nor UO_3336 (O_3336,N_29278,N_29932);
xnor UO_3337 (O_3337,N_29601,N_29579);
or UO_3338 (O_3338,N_29431,N_29284);
nor UO_3339 (O_3339,N_29623,N_29745);
or UO_3340 (O_3340,N_29220,N_29283);
or UO_3341 (O_3341,N_29618,N_29719);
and UO_3342 (O_3342,N_29134,N_29150);
nor UO_3343 (O_3343,N_29789,N_29279);
or UO_3344 (O_3344,N_29585,N_29851);
nor UO_3345 (O_3345,N_29735,N_29302);
xor UO_3346 (O_3346,N_29924,N_29823);
and UO_3347 (O_3347,N_29853,N_29971);
or UO_3348 (O_3348,N_29033,N_29337);
or UO_3349 (O_3349,N_29674,N_29971);
nor UO_3350 (O_3350,N_29604,N_29699);
xor UO_3351 (O_3351,N_29130,N_29584);
nand UO_3352 (O_3352,N_29494,N_29658);
xnor UO_3353 (O_3353,N_29895,N_29149);
nand UO_3354 (O_3354,N_29103,N_29958);
xor UO_3355 (O_3355,N_29812,N_29861);
or UO_3356 (O_3356,N_29463,N_29241);
xnor UO_3357 (O_3357,N_29145,N_29174);
nand UO_3358 (O_3358,N_29054,N_29993);
nor UO_3359 (O_3359,N_29190,N_29233);
and UO_3360 (O_3360,N_29906,N_29751);
or UO_3361 (O_3361,N_29425,N_29581);
or UO_3362 (O_3362,N_29463,N_29394);
nor UO_3363 (O_3363,N_29486,N_29644);
or UO_3364 (O_3364,N_29045,N_29533);
or UO_3365 (O_3365,N_29365,N_29647);
nor UO_3366 (O_3366,N_29091,N_29889);
nand UO_3367 (O_3367,N_29292,N_29280);
or UO_3368 (O_3368,N_29877,N_29257);
xnor UO_3369 (O_3369,N_29301,N_29266);
xnor UO_3370 (O_3370,N_29380,N_29697);
and UO_3371 (O_3371,N_29076,N_29056);
nor UO_3372 (O_3372,N_29226,N_29546);
nor UO_3373 (O_3373,N_29495,N_29752);
or UO_3374 (O_3374,N_29090,N_29831);
nand UO_3375 (O_3375,N_29884,N_29247);
nor UO_3376 (O_3376,N_29535,N_29927);
and UO_3377 (O_3377,N_29818,N_29505);
or UO_3378 (O_3378,N_29965,N_29942);
or UO_3379 (O_3379,N_29211,N_29489);
or UO_3380 (O_3380,N_29711,N_29552);
xnor UO_3381 (O_3381,N_29060,N_29659);
and UO_3382 (O_3382,N_29731,N_29835);
nand UO_3383 (O_3383,N_29928,N_29528);
and UO_3384 (O_3384,N_29521,N_29224);
and UO_3385 (O_3385,N_29971,N_29586);
nand UO_3386 (O_3386,N_29978,N_29644);
and UO_3387 (O_3387,N_29818,N_29942);
nand UO_3388 (O_3388,N_29912,N_29014);
nand UO_3389 (O_3389,N_29886,N_29326);
and UO_3390 (O_3390,N_29251,N_29712);
or UO_3391 (O_3391,N_29131,N_29855);
and UO_3392 (O_3392,N_29556,N_29029);
and UO_3393 (O_3393,N_29805,N_29204);
nand UO_3394 (O_3394,N_29576,N_29358);
xnor UO_3395 (O_3395,N_29792,N_29887);
xor UO_3396 (O_3396,N_29285,N_29159);
and UO_3397 (O_3397,N_29501,N_29641);
and UO_3398 (O_3398,N_29414,N_29274);
xor UO_3399 (O_3399,N_29709,N_29147);
or UO_3400 (O_3400,N_29255,N_29617);
nand UO_3401 (O_3401,N_29192,N_29261);
and UO_3402 (O_3402,N_29218,N_29088);
xnor UO_3403 (O_3403,N_29805,N_29953);
nor UO_3404 (O_3404,N_29414,N_29565);
xor UO_3405 (O_3405,N_29139,N_29785);
xor UO_3406 (O_3406,N_29052,N_29036);
and UO_3407 (O_3407,N_29334,N_29474);
xnor UO_3408 (O_3408,N_29536,N_29048);
nand UO_3409 (O_3409,N_29329,N_29415);
nor UO_3410 (O_3410,N_29528,N_29491);
or UO_3411 (O_3411,N_29102,N_29444);
and UO_3412 (O_3412,N_29227,N_29332);
nor UO_3413 (O_3413,N_29858,N_29969);
xnor UO_3414 (O_3414,N_29159,N_29793);
xor UO_3415 (O_3415,N_29087,N_29499);
or UO_3416 (O_3416,N_29258,N_29090);
or UO_3417 (O_3417,N_29668,N_29287);
or UO_3418 (O_3418,N_29793,N_29221);
nor UO_3419 (O_3419,N_29970,N_29935);
nor UO_3420 (O_3420,N_29523,N_29681);
or UO_3421 (O_3421,N_29850,N_29072);
xor UO_3422 (O_3422,N_29802,N_29639);
and UO_3423 (O_3423,N_29311,N_29857);
xor UO_3424 (O_3424,N_29735,N_29747);
and UO_3425 (O_3425,N_29486,N_29681);
xor UO_3426 (O_3426,N_29161,N_29648);
and UO_3427 (O_3427,N_29742,N_29939);
nor UO_3428 (O_3428,N_29086,N_29764);
nor UO_3429 (O_3429,N_29632,N_29667);
and UO_3430 (O_3430,N_29007,N_29855);
and UO_3431 (O_3431,N_29002,N_29547);
and UO_3432 (O_3432,N_29019,N_29915);
nor UO_3433 (O_3433,N_29020,N_29338);
nor UO_3434 (O_3434,N_29917,N_29969);
or UO_3435 (O_3435,N_29244,N_29971);
nand UO_3436 (O_3436,N_29683,N_29390);
and UO_3437 (O_3437,N_29559,N_29207);
xor UO_3438 (O_3438,N_29985,N_29824);
and UO_3439 (O_3439,N_29867,N_29636);
and UO_3440 (O_3440,N_29389,N_29635);
nand UO_3441 (O_3441,N_29109,N_29282);
xor UO_3442 (O_3442,N_29487,N_29341);
nor UO_3443 (O_3443,N_29538,N_29912);
and UO_3444 (O_3444,N_29450,N_29060);
nand UO_3445 (O_3445,N_29737,N_29824);
nand UO_3446 (O_3446,N_29679,N_29773);
nand UO_3447 (O_3447,N_29679,N_29124);
nor UO_3448 (O_3448,N_29731,N_29231);
or UO_3449 (O_3449,N_29955,N_29797);
or UO_3450 (O_3450,N_29203,N_29015);
nand UO_3451 (O_3451,N_29817,N_29060);
and UO_3452 (O_3452,N_29128,N_29139);
and UO_3453 (O_3453,N_29800,N_29187);
nor UO_3454 (O_3454,N_29591,N_29802);
nor UO_3455 (O_3455,N_29936,N_29994);
nor UO_3456 (O_3456,N_29839,N_29071);
xor UO_3457 (O_3457,N_29493,N_29595);
or UO_3458 (O_3458,N_29012,N_29312);
or UO_3459 (O_3459,N_29422,N_29326);
and UO_3460 (O_3460,N_29524,N_29226);
nor UO_3461 (O_3461,N_29380,N_29310);
xnor UO_3462 (O_3462,N_29399,N_29560);
xor UO_3463 (O_3463,N_29638,N_29315);
nand UO_3464 (O_3464,N_29691,N_29578);
nand UO_3465 (O_3465,N_29242,N_29963);
xor UO_3466 (O_3466,N_29355,N_29459);
or UO_3467 (O_3467,N_29259,N_29813);
nor UO_3468 (O_3468,N_29566,N_29111);
nor UO_3469 (O_3469,N_29133,N_29212);
or UO_3470 (O_3470,N_29854,N_29663);
xnor UO_3471 (O_3471,N_29250,N_29652);
nand UO_3472 (O_3472,N_29186,N_29683);
and UO_3473 (O_3473,N_29085,N_29278);
or UO_3474 (O_3474,N_29655,N_29128);
nand UO_3475 (O_3475,N_29248,N_29563);
or UO_3476 (O_3476,N_29875,N_29877);
or UO_3477 (O_3477,N_29098,N_29068);
xnor UO_3478 (O_3478,N_29002,N_29882);
nor UO_3479 (O_3479,N_29118,N_29090);
and UO_3480 (O_3480,N_29441,N_29151);
xor UO_3481 (O_3481,N_29003,N_29341);
xnor UO_3482 (O_3482,N_29089,N_29329);
xor UO_3483 (O_3483,N_29105,N_29521);
or UO_3484 (O_3484,N_29334,N_29449);
or UO_3485 (O_3485,N_29064,N_29104);
and UO_3486 (O_3486,N_29863,N_29945);
xor UO_3487 (O_3487,N_29537,N_29289);
xor UO_3488 (O_3488,N_29897,N_29431);
xnor UO_3489 (O_3489,N_29921,N_29136);
nand UO_3490 (O_3490,N_29971,N_29794);
and UO_3491 (O_3491,N_29960,N_29069);
nand UO_3492 (O_3492,N_29497,N_29765);
and UO_3493 (O_3493,N_29151,N_29899);
and UO_3494 (O_3494,N_29857,N_29305);
nor UO_3495 (O_3495,N_29068,N_29956);
and UO_3496 (O_3496,N_29507,N_29007);
xnor UO_3497 (O_3497,N_29126,N_29125);
nor UO_3498 (O_3498,N_29487,N_29831);
and UO_3499 (O_3499,N_29147,N_29596);
endmodule