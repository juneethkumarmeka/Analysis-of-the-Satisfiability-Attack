module basic_1000_10000_1500_100_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_97,In_749);
nand U1 (N_1,In_397,In_216);
or U2 (N_2,In_825,In_170);
or U3 (N_3,In_722,In_500);
nor U4 (N_4,In_910,In_537);
or U5 (N_5,In_769,In_795);
nor U6 (N_6,In_912,In_871);
nand U7 (N_7,In_328,In_411);
xnor U8 (N_8,In_876,In_259);
nor U9 (N_9,In_800,In_830);
nand U10 (N_10,In_937,In_599);
nor U11 (N_11,In_592,In_736);
nor U12 (N_12,In_196,In_396);
nand U13 (N_13,In_545,In_956);
nor U14 (N_14,In_447,In_782);
nand U15 (N_15,In_883,In_509);
nor U16 (N_16,In_843,In_174);
or U17 (N_17,In_460,In_383);
nand U18 (N_18,In_289,In_542);
or U19 (N_19,In_631,In_718);
or U20 (N_20,In_12,In_898);
nand U21 (N_21,In_728,In_819);
nor U22 (N_22,In_483,In_400);
and U23 (N_23,In_760,In_868);
and U24 (N_24,In_475,In_821);
or U25 (N_25,In_245,In_671);
nand U26 (N_26,In_637,In_829);
and U27 (N_27,In_859,In_319);
nand U28 (N_28,In_850,In_504);
nand U29 (N_29,In_979,In_371);
or U30 (N_30,In_22,In_226);
and U31 (N_31,In_163,In_762);
nor U32 (N_32,In_812,In_561);
nand U33 (N_33,In_961,In_523);
and U34 (N_34,In_484,In_392);
nor U35 (N_35,In_747,In_982);
nand U36 (N_36,In_298,In_354);
or U37 (N_37,In_972,In_564);
or U38 (N_38,In_835,In_607);
nor U39 (N_39,In_838,In_881);
and U40 (N_40,In_546,In_175);
and U41 (N_41,In_75,In_647);
nor U42 (N_42,In_58,In_306);
nor U43 (N_43,In_33,In_326);
or U44 (N_44,In_697,In_53);
nand U45 (N_45,In_709,In_330);
and U46 (N_46,In_863,In_449);
or U47 (N_47,In_290,In_781);
and U48 (N_48,In_42,In_414);
or U49 (N_49,In_322,In_200);
and U50 (N_50,In_969,In_717);
xnor U51 (N_51,In_359,In_468);
nand U52 (N_52,In_737,In_38);
and U53 (N_53,In_846,In_69);
or U54 (N_54,In_195,In_182);
nand U55 (N_55,In_344,In_403);
nor U56 (N_56,In_650,In_817);
nor U57 (N_57,In_249,In_572);
and U58 (N_58,In_896,In_528);
nor U59 (N_59,In_673,In_375);
nor U60 (N_60,In_792,In_530);
nor U61 (N_61,In_402,In_466);
and U62 (N_62,In_649,In_930);
or U63 (N_63,In_101,In_852);
or U64 (N_64,In_629,In_343);
nor U65 (N_65,In_352,In_511);
nand U66 (N_66,In_373,In_329);
or U67 (N_67,In_615,In_774);
nand U68 (N_68,In_52,In_254);
or U69 (N_69,In_278,In_95);
or U70 (N_70,In_531,In_155);
nand U71 (N_71,In_444,In_809);
and U72 (N_72,In_418,In_297);
nor U73 (N_73,In_25,In_560);
and U74 (N_74,In_712,In_136);
nor U75 (N_75,In_492,In_146);
nand U76 (N_76,In_268,In_574);
nor U77 (N_77,In_513,In_235);
and U78 (N_78,In_684,In_177);
nand U79 (N_79,In_655,In_860);
nor U80 (N_80,In_653,In_312);
or U81 (N_81,In_368,In_695);
or U82 (N_82,In_630,In_794);
or U83 (N_83,In_462,In_968);
nand U84 (N_84,In_166,In_144);
xnor U85 (N_85,In_395,In_508);
nand U86 (N_86,In_743,In_331);
and U87 (N_87,In_291,In_744);
nand U88 (N_88,In_159,In_596);
and U89 (N_89,In_944,In_148);
nand U90 (N_90,In_798,In_349);
or U91 (N_91,In_457,In_748);
and U92 (N_92,In_40,In_44);
nand U93 (N_93,In_490,In_597);
nand U94 (N_94,In_233,In_640);
or U95 (N_95,In_217,In_454);
or U96 (N_96,In_582,In_141);
nand U97 (N_97,In_435,In_686);
nor U98 (N_98,In_1,In_559);
nand U99 (N_99,In_273,In_156);
or U100 (N_100,N_14,In_690);
nor U101 (N_101,In_20,In_773);
nand U102 (N_102,In_365,In_606);
nand U103 (N_103,In_91,In_147);
nand U104 (N_104,In_142,In_427);
xor U105 (N_105,In_23,In_771);
nor U106 (N_106,In_525,N_2);
and U107 (N_107,N_78,In_237);
and U108 (N_108,In_699,In_301);
nand U109 (N_109,In_557,In_279);
nand U110 (N_110,In_303,N_19);
nand U111 (N_111,In_106,In_369);
and U112 (N_112,In_394,In_866);
or U113 (N_113,In_520,In_393);
or U114 (N_114,In_317,N_31);
nor U115 (N_115,In_884,In_121);
nand U116 (N_116,In_952,In_936);
and U117 (N_117,In_120,In_378);
or U118 (N_118,In_849,In_307);
or U119 (N_119,In_433,In_676);
nor U120 (N_120,In_446,In_935);
and U121 (N_121,In_925,In_797);
or U122 (N_122,In_151,In_85);
or U123 (N_123,In_929,In_502);
and U124 (N_124,N_13,In_818);
or U125 (N_125,In_46,In_730);
or U126 (N_126,In_419,In_527);
nor U127 (N_127,In_11,In_953);
or U128 (N_128,In_927,In_598);
nor U129 (N_129,In_602,In_239);
nor U130 (N_130,In_976,In_16);
or U131 (N_131,In_108,In_39);
nand U132 (N_132,In_720,In_612);
nor U133 (N_133,In_84,N_88);
nor U134 (N_134,In_315,In_864);
nand U135 (N_135,N_49,In_996);
nor U136 (N_136,In_872,In_350);
nand U137 (N_137,In_495,In_325);
nor U138 (N_138,In_501,In_337);
nand U139 (N_139,In_779,In_130);
and U140 (N_140,In_198,In_295);
nand U141 (N_141,In_215,N_17);
nor U142 (N_142,In_918,In_455);
and U143 (N_143,In_841,In_478);
nand U144 (N_144,In_932,In_68);
and U145 (N_145,In_32,In_900);
or U146 (N_146,In_288,In_664);
nand U147 (N_147,In_206,In_905);
or U148 (N_148,In_406,In_113);
nand U149 (N_149,In_138,In_831);
nor U150 (N_150,In_933,In_128);
nor U151 (N_151,In_78,In_994);
and U152 (N_152,In_242,In_429);
or U153 (N_153,In_659,In_210);
or U154 (N_154,N_64,In_152);
nor U155 (N_155,In_86,In_669);
nor U156 (N_156,In_745,In_993);
nor U157 (N_157,In_710,In_417);
or U158 (N_158,In_549,In_687);
and U159 (N_159,In_26,In_90);
and U160 (N_160,In_983,N_52);
or U161 (N_161,In_625,In_274);
nand U162 (N_162,N_22,In_309);
and U163 (N_163,N_9,In_844);
nor U164 (N_164,In_981,In_584);
nor U165 (N_165,In_674,In_480);
nand U166 (N_166,In_593,In_256);
nand U167 (N_167,N_56,In_610);
nand U168 (N_168,N_62,In_639);
and U169 (N_169,In_974,N_45);
nor U170 (N_170,In_102,In_536);
nor U171 (N_171,In_636,In_139);
or U172 (N_172,In_305,In_180);
nand U173 (N_173,In_758,In_401);
and U174 (N_174,In_802,In_558);
or U175 (N_175,N_53,N_30);
and U176 (N_176,In_264,In_158);
nand U177 (N_177,In_556,In_390);
nor U178 (N_178,In_928,In_336);
nand U179 (N_179,In_914,N_75);
or U180 (N_180,In_284,N_32);
nor U181 (N_181,In_185,In_742);
and U182 (N_182,In_547,In_704);
nor U183 (N_183,In_551,In_188);
nor U184 (N_184,In_469,In_618);
or U185 (N_185,N_48,In_725);
and U186 (N_186,In_764,N_38);
and U187 (N_187,In_585,In_241);
and U188 (N_188,In_342,In_497);
or U189 (N_189,In_660,In_608);
nor U190 (N_190,In_258,In_260);
and U191 (N_191,In_765,In_988);
nor U192 (N_192,In_110,In_755);
and U193 (N_193,In_27,In_432);
nor U194 (N_194,N_23,In_589);
nor U195 (N_195,N_10,In_275);
nand U196 (N_196,In_895,In_796);
and U197 (N_197,In_958,In_470);
nand U198 (N_198,In_362,In_515);
nand U199 (N_199,In_338,In_57);
and U200 (N_200,In_201,In_202);
and U201 (N_201,In_897,In_964);
nand U202 (N_202,N_182,In_247);
nand U203 (N_203,In_950,In_287);
nor U204 (N_204,In_127,N_185);
nor U205 (N_205,In_145,In_778);
nor U206 (N_206,N_82,In_197);
nor U207 (N_207,In_735,In_565);
nor U208 (N_208,N_24,In_203);
and U209 (N_209,In_116,N_195);
and U210 (N_210,In_685,In_334);
and U211 (N_211,In_316,N_150);
nor U212 (N_212,In_100,In_665);
and U213 (N_213,In_232,In_999);
nor U214 (N_214,In_277,In_601);
nor U215 (N_215,In_757,N_163);
nand U216 (N_216,N_181,In_842);
xnor U217 (N_217,In_439,In_496);
nor U218 (N_218,N_140,In_923);
or U219 (N_219,In_135,In_548);
and U220 (N_220,In_696,In_571);
or U221 (N_221,In_761,In_41);
or U222 (N_222,In_476,In_516);
or U223 (N_223,In_399,In_398);
nor U224 (N_224,In_253,N_84);
nor U225 (N_225,N_151,In_739);
nor U226 (N_226,In_555,In_357);
nand U227 (N_227,In_211,In_966);
nor U228 (N_228,In_759,In_766);
nand U229 (N_229,In_705,In_17);
or U230 (N_230,In_93,In_791);
and U231 (N_231,N_125,In_387);
nand U232 (N_232,In_31,N_108);
nand U233 (N_233,In_207,N_142);
and U234 (N_234,In_991,N_138);
xor U235 (N_235,In_244,N_166);
or U236 (N_236,In_213,In_834);
nand U237 (N_237,In_886,In_753);
or U238 (N_238,N_93,N_177);
xor U239 (N_239,N_101,In_348);
or U240 (N_240,In_21,In_729);
nand U241 (N_241,In_575,In_892);
and U242 (N_242,N_190,In_865);
or U243 (N_243,In_304,In_689);
and U244 (N_244,In_230,In_553);
or U245 (N_245,In_486,In_916);
nor U246 (N_246,In_702,In_472);
and U247 (N_247,In_990,N_103);
or U248 (N_248,In_915,In_190);
or U249 (N_249,In_236,In_828);
and U250 (N_250,In_998,In_566);
nand U251 (N_251,In_430,In_358);
nand U252 (N_252,In_889,In_627);
or U253 (N_253,In_0,In_420);
or U254 (N_254,In_436,In_815);
or U255 (N_255,In_543,In_36);
nor U256 (N_256,N_172,N_11);
nand U257 (N_257,In_124,In_82);
or U258 (N_258,In_171,In_6);
or U259 (N_259,In_464,N_6);
or U260 (N_260,In_780,N_94);
nand U261 (N_261,N_137,In_262);
xnor U262 (N_262,In_481,In_807);
nor U263 (N_263,In_388,In_66);
or U264 (N_264,In_657,In_111);
nor U265 (N_265,In_54,In_839);
or U266 (N_266,N_147,In_347);
xor U267 (N_267,In_806,In_594);
xnor U268 (N_268,In_134,In_805);
or U269 (N_269,N_171,N_67);
or U270 (N_270,N_129,In_827);
nor U271 (N_271,N_118,In_521);
nor U272 (N_272,In_873,In_228);
and U273 (N_273,In_512,In_59);
nand U274 (N_274,In_678,N_18);
or U275 (N_275,In_443,In_356);
and U276 (N_276,In_614,In_30);
and U277 (N_277,In_353,In_482);
and U278 (N_278,In_672,In_568);
nand U279 (N_279,In_510,N_65);
nor U280 (N_280,In_29,In_526);
nand U281 (N_281,In_72,In_783);
or U282 (N_282,In_931,In_24);
and U283 (N_283,In_224,In_711);
nand U284 (N_284,In_89,In_114);
or U285 (N_285,N_89,In_28);
or U286 (N_286,In_65,N_174);
or U287 (N_287,In_70,In_726);
or U288 (N_288,In_76,In_246);
and U289 (N_289,In_341,In_376);
nand U290 (N_290,In_445,In_532);
or U291 (N_291,In_267,In_112);
nand U292 (N_292,N_144,N_46);
or U293 (N_293,In_220,In_219);
nor U294 (N_294,In_77,In_724);
nor U295 (N_295,In_173,In_281);
or U296 (N_296,In_734,In_300);
and U297 (N_297,In_14,In_441);
nand U298 (N_298,N_55,In_943);
nand U299 (N_299,N_127,N_130);
nor U300 (N_300,In_586,In_768);
nand U301 (N_301,N_28,In_719);
nand U302 (N_302,In_541,In_977);
nand U303 (N_303,N_291,In_345);
or U304 (N_304,In_662,In_652);
and U305 (N_305,In_56,In_634);
or U306 (N_306,In_540,N_102);
or U307 (N_307,N_180,In_503);
nand U308 (N_308,N_189,In_855);
or U309 (N_309,In_364,In_212);
and U310 (N_310,N_139,In_756);
nor U311 (N_311,N_109,In_692);
nor U312 (N_312,In_117,In_194);
or U313 (N_313,In_311,In_271);
nor U314 (N_314,In_485,In_183);
and U315 (N_315,In_938,In_878);
nor U316 (N_316,In_448,In_310);
nor U317 (N_317,N_205,In_885);
nor U318 (N_318,In_787,In_962);
nand U319 (N_319,N_98,In_869);
or U320 (N_320,N_209,N_95);
or U321 (N_321,N_41,In_64);
nor U322 (N_322,In_813,In_980);
and U323 (N_323,In_833,N_60);
or U324 (N_324,In_456,N_105);
nand U325 (N_325,In_721,In_494);
or U326 (N_326,In_880,In_940);
nand U327 (N_327,In_716,In_491);
nor U328 (N_328,N_215,In_161);
and U329 (N_329,In_189,In_870);
nand U330 (N_330,N_219,In_477);
and U331 (N_331,N_238,N_197);
and U332 (N_332,In_221,N_253);
or U333 (N_333,In_479,In_733);
and U334 (N_334,In_79,N_112);
and U335 (N_335,In_48,N_96);
or U336 (N_336,N_155,N_107);
or U337 (N_337,In_374,In_837);
or U338 (N_338,In_554,N_222);
or U339 (N_339,N_200,In_908);
and U340 (N_340,In_851,N_87);
nor U341 (N_341,N_210,In_296);
or U342 (N_342,N_201,In_913);
nand U343 (N_343,In_656,N_162);
nor U344 (N_344,N_20,In_83);
and U345 (N_345,In_770,In_604);
nor U346 (N_346,In_382,N_226);
nand U347 (N_347,In_562,N_74);
and U348 (N_348,In_715,N_218);
nand U349 (N_349,In_891,N_231);
or U350 (N_350,In_569,N_211);
nand U351 (N_351,N_39,In_680);
nor U352 (N_352,In_641,In_984);
nand U353 (N_353,In_363,In_985);
or U354 (N_354,N_265,In_240);
and U355 (N_355,N_120,In_626);
nor U356 (N_356,N_117,In_847);
or U357 (N_357,N_186,In_590);
nand U358 (N_358,In_164,In_738);
and U359 (N_359,N_91,N_51);
or U360 (N_360,In_600,In_621);
nor U361 (N_361,In_587,N_132);
or U362 (N_362,In_119,In_693);
nor U363 (N_363,N_16,In_208);
and U364 (N_364,N_164,N_235);
nor U365 (N_365,In_461,In_438);
nor U366 (N_366,In_205,N_42);
nor U367 (N_367,N_35,In_645);
nand U368 (N_368,N_224,In_804);
or U369 (N_369,In_204,In_663);
nand U370 (N_370,In_285,N_83);
and U371 (N_371,In_820,N_81);
or U372 (N_372,In_920,In_661);
nor U373 (N_373,In_965,In_10);
and U374 (N_374,In_708,N_232);
nor U375 (N_375,N_79,In_514);
and U376 (N_376,N_179,In_917);
nand U377 (N_377,In_622,In_67);
nand U378 (N_378,In_499,In_8);
nor U379 (N_379,In_370,N_50);
nand U380 (N_380,In_654,In_71);
and U381 (N_381,In_47,In_723);
or U382 (N_382,In_423,N_193);
nor U383 (N_383,N_233,In_675);
xor U384 (N_384,N_0,In_955);
and U385 (N_385,In_619,In_179);
nand U386 (N_386,In_313,N_192);
nor U387 (N_387,In_377,In_519);
nor U388 (N_388,In_225,In_366);
or U389 (N_389,In_963,N_4);
nand U390 (N_390,In_939,In_123);
or U391 (N_391,In_172,In_405);
and U392 (N_392,In_416,In_168);
nand U393 (N_393,N_61,N_77);
and U394 (N_394,In_181,In_854);
or U395 (N_395,In_507,N_5);
nand U396 (N_396,N_156,In_154);
and U397 (N_397,In_875,In_570);
or U398 (N_398,In_971,In_270);
and U399 (N_399,In_442,N_227);
xnor U400 (N_400,In_103,N_383);
nor U401 (N_401,N_212,N_364);
and U402 (N_402,In_35,In_577);
or U403 (N_403,In_465,N_100);
nand U404 (N_404,N_249,N_111);
or U405 (N_405,In_104,In_628);
nand U406 (N_406,In_617,In_882);
or U407 (N_407,N_256,N_274);
and U408 (N_408,In_648,N_298);
nand U409 (N_409,In_934,N_350);
nand U410 (N_410,N_339,N_239);
and U411 (N_411,N_183,N_187);
and U412 (N_412,N_334,In_493);
nand U413 (N_413,In_624,N_304);
nand U414 (N_414,N_143,In_945);
and U415 (N_415,In_997,In_184);
or U416 (N_416,N_397,In_37);
nor U417 (N_417,In_360,N_242);
and U418 (N_418,In_583,N_237);
xor U419 (N_419,N_25,N_208);
or U420 (N_420,In_970,N_1);
nand U421 (N_421,N_260,In_13);
nor U422 (N_422,N_160,N_283);
or U423 (N_423,In_61,In_458);
and U424 (N_424,N_338,N_340);
and U425 (N_425,N_234,N_203);
and U426 (N_426,N_216,N_251);
nand U427 (N_427,N_168,In_98);
or U428 (N_428,In_257,In_380);
and U429 (N_429,In_74,In_73);
or U430 (N_430,N_191,N_376);
nor U431 (N_431,In_763,N_159);
nor U432 (N_432,In_453,N_348);
and U433 (N_433,N_271,N_76);
or U434 (N_434,In_186,N_199);
nor U435 (N_435,N_354,N_290);
and U436 (N_436,In_899,In_167);
nand U437 (N_437,In_518,N_169);
nor U438 (N_438,In_836,N_393);
xnor U439 (N_439,In_412,N_358);
nor U440 (N_440,In_772,In_49);
nand U441 (N_441,N_264,N_153);
nand U442 (N_442,In_434,N_297);
nor U443 (N_443,N_278,In_799);
nand U444 (N_444,N_167,In_498);
and U445 (N_445,N_299,N_40);
and U446 (N_446,In_995,N_27);
nor U447 (N_447,N_71,N_33);
nand U448 (N_448,In_276,In_901);
nor U449 (N_449,In_3,In_251);
nor U450 (N_450,In_580,In_238);
or U451 (N_451,N_289,In_909);
and U452 (N_452,N_316,In_428);
and U453 (N_453,In_713,N_8);
or U454 (N_454,N_245,In_632);
or U455 (N_455,In_125,In_750);
nand U456 (N_456,In_776,In_578);
and U457 (N_457,In_814,In_157);
nor U458 (N_458,In_234,In_682);
and U459 (N_459,N_99,In_292);
xnor U460 (N_460,In_822,In_978);
nand U461 (N_461,N_341,In_529);
or U462 (N_462,N_361,In_50);
or U463 (N_463,In_524,In_137);
nor U464 (N_464,In_280,N_15);
and U465 (N_465,N_252,In_450);
or U466 (N_466,In_118,N_225);
nand U467 (N_467,In_751,In_333);
nand U468 (N_468,N_21,In_209);
nand U469 (N_469,In_591,In_80);
nor U470 (N_470,In_143,In_691);
nor U471 (N_471,N_196,In_698);
nand U472 (N_472,In_266,In_947);
and U473 (N_473,In_214,N_247);
and U474 (N_474,In_272,In_283);
or U475 (N_475,N_214,N_284);
xnor U476 (N_476,N_318,N_141);
and U477 (N_477,N_327,N_323);
nor U478 (N_478,In_231,N_309);
nand U479 (N_479,In_355,N_126);
nor U480 (N_480,In_340,N_80);
or U481 (N_481,N_360,In_613);
nor U482 (N_482,N_396,N_377);
or U483 (N_483,In_563,N_286);
nand U484 (N_484,In_440,In_243);
nor U485 (N_485,In_987,N_336);
and U486 (N_486,In_906,N_365);
xnor U487 (N_487,In_165,In_385);
nand U488 (N_488,In_302,N_58);
or U489 (N_489,N_204,In_389);
nand U490 (N_490,N_243,N_70);
and U491 (N_491,N_388,N_250);
and U492 (N_492,N_26,In_19);
or U493 (N_493,In_620,N_395);
and U494 (N_494,N_198,In_45);
nor U495 (N_495,N_157,N_375);
and U496 (N_496,In_609,In_951);
nand U497 (N_497,N_154,N_344);
nor U498 (N_498,In_107,N_254);
and U499 (N_499,N_300,N_276);
nor U500 (N_500,In_192,N_275);
nor U501 (N_501,N_221,In_109);
and U502 (N_502,In_643,N_63);
or U503 (N_503,N_229,In_153);
nor U504 (N_504,In_823,In_706);
or U505 (N_505,N_255,N_115);
or U506 (N_506,N_310,In_299);
nor U507 (N_507,N_461,In_677);
nand U508 (N_508,N_385,N_427);
nor U509 (N_509,N_241,N_43);
nand U510 (N_510,In_87,N_362);
or U511 (N_511,N_330,In_94);
and U512 (N_512,In_848,N_90);
or U513 (N_513,N_295,In_921);
or U514 (N_514,In_658,N_455);
or U515 (N_515,In_579,In_989);
and U516 (N_516,In_874,N_442);
nand U517 (N_517,In_261,N_355);
and U518 (N_518,N_411,In_616);
or U519 (N_519,N_47,In_623);
and U520 (N_520,N_470,In_741);
nand U521 (N_521,In_150,In_856);
nor U522 (N_522,In_321,N_418);
nand U523 (N_523,In_867,In_960);
nor U524 (N_524,N_29,N_146);
and U525 (N_525,N_417,In_642);
nor U526 (N_526,N_440,In_332);
and U527 (N_527,N_445,N_366);
nand U528 (N_528,N_346,N_206);
or U529 (N_529,N_477,N_175);
nand U530 (N_530,N_478,N_259);
nand U531 (N_531,N_282,In_576);
nor U532 (N_532,N_457,N_401);
nor U533 (N_533,N_479,N_400);
and U534 (N_534,In_140,N_424);
nor U535 (N_535,In_694,N_421);
nor U536 (N_536,In_487,N_321);
nor U537 (N_537,N_301,N_268);
and U538 (N_538,N_448,In_973);
and U539 (N_539,In_407,N_374);
or U540 (N_540,In_894,In_60);
or U541 (N_541,In_911,N_389);
or U542 (N_542,N_165,N_353);
and U543 (N_543,In_538,N_439);
nand U544 (N_544,N_428,In_603);
or U545 (N_545,N_266,In_679);
nand U546 (N_546,N_430,N_443);
or U547 (N_547,N_463,N_392);
or U548 (N_548,In_811,In_149);
nand U549 (N_549,In_902,N_272);
or U550 (N_550,In_505,In_784);
and U551 (N_551,N_472,In_926);
or U552 (N_552,In_473,N_314);
nor U553 (N_553,N_460,In_688);
or U554 (N_554,N_450,In_919);
nand U555 (N_555,N_122,N_458);
nand U556 (N_556,In_408,In_187);
or U557 (N_557,N_408,N_145);
nand U558 (N_558,In_415,In_904);
and U559 (N_559,N_329,In_824);
nand U560 (N_560,In_263,In_890);
nor U561 (N_561,N_294,In_4);
nand U562 (N_562,N_34,N_114);
or U563 (N_563,In_269,In_162);
and U564 (N_564,In_948,N_465);
nand U565 (N_565,N_373,In_732);
nand U566 (N_566,N_57,In_635);
nand U567 (N_567,N_453,N_494);
and U568 (N_568,N_467,N_288);
nand U569 (N_569,N_312,N_482);
nand U570 (N_570,In_115,In_506);
nor U571 (N_571,N_356,N_369);
and U572 (N_572,N_337,In_327);
nor U573 (N_573,N_409,In_320);
and U574 (N_574,N_258,In_746);
nand U575 (N_575,N_496,N_384);
nand U576 (N_576,In_409,In_459);
and U577 (N_577,In_522,In_752);
nor U578 (N_578,In_122,In_294);
and U579 (N_579,N_452,In_858);
and U580 (N_580,N_170,In_853);
nand U581 (N_581,In_573,In_703);
nand U582 (N_582,In_701,N_415);
nand U583 (N_583,In_467,N_498);
nor U584 (N_584,In_218,In_941);
nand U585 (N_585,N_474,N_335);
or U586 (N_586,N_69,In_421);
nand U587 (N_587,N_497,In_34);
nand U588 (N_588,In_790,In_740);
nor U589 (N_589,N_342,In_7);
or U590 (N_590,N_473,N_422);
and U591 (N_591,N_446,In_133);
or U592 (N_592,In_426,N_444);
and U593 (N_593,In_788,N_352);
or U594 (N_594,N_404,N_499);
and U595 (N_595,N_308,N_263);
nor U596 (N_596,N_236,N_485);
or U597 (N_597,N_416,N_419);
or U598 (N_598,In_43,N_287);
xnor U599 (N_599,In_199,N_277);
or U600 (N_600,N_326,N_503);
or U601 (N_601,N_518,N_536);
and U602 (N_602,N_511,In_55);
nand U603 (N_603,N_184,In_431);
nand U604 (N_604,N_128,N_584);
and U605 (N_605,N_390,N_123);
nand U606 (N_606,N_223,N_423);
or U607 (N_607,N_548,N_593);
and U608 (N_608,In_857,N_113);
nor U609 (N_609,N_333,N_513);
or U610 (N_610,In_132,N_176);
nor U611 (N_611,In_63,N_320);
or U612 (N_612,N_583,In_605);
nor U613 (N_613,N_386,N_522);
or U614 (N_614,N_406,In_893);
nand U615 (N_615,In_877,N_563);
or U616 (N_616,N_519,In_437);
nand U617 (N_617,N_213,N_578);
or U618 (N_618,In_178,N_525);
nand U619 (N_619,In_223,In_451);
or U620 (N_620,In_957,N_596);
nand U621 (N_621,N_580,N_431);
or U622 (N_622,N_567,In_81);
or U623 (N_623,N_468,N_106);
and U624 (N_624,In_949,N_562);
and U625 (N_625,N_487,N_549);
and U626 (N_626,N_194,N_305);
nand U627 (N_627,In_588,N_573);
and U628 (N_628,N_331,In_651);
nand U629 (N_629,N_92,N_257);
nand U630 (N_630,N_217,N_124);
or U631 (N_631,In_638,N_261);
nor U632 (N_632,N_528,In_611);
or U633 (N_633,In_670,In_99);
and U634 (N_634,In_384,N_68);
nor U635 (N_635,In_731,N_437);
and U636 (N_636,N_292,N_207);
nor U637 (N_637,N_509,In_424);
nor U638 (N_638,In_785,N_381);
and U639 (N_639,N_515,In_633);
nor U640 (N_640,N_557,N_273);
or U641 (N_641,N_405,N_378);
nand U642 (N_642,In_62,N_582);
or U643 (N_643,In_808,In_18);
nand U644 (N_644,N_484,N_441);
nand U645 (N_645,N_398,In_975);
or U646 (N_646,N_97,N_425);
or U647 (N_647,In_314,In_840);
or U648 (N_648,N_558,N_152);
nor U649 (N_649,N_501,In_410);
or U650 (N_650,N_37,In_489);
and U651 (N_651,N_315,In_131);
nand U652 (N_652,In_667,N_280);
nor U653 (N_653,In_544,N_502);
and U654 (N_654,In_265,In_946);
nor U655 (N_655,N_454,N_85);
nor U656 (N_656,N_476,N_402);
and U657 (N_657,N_178,N_570);
nor U658 (N_658,N_391,N_54);
xnor U659 (N_659,N_119,N_306);
nor U660 (N_660,In_222,N_506);
nor U661 (N_661,In_861,In_367);
or U662 (N_662,N_527,N_173);
nor U663 (N_663,N_134,In_845);
and U664 (N_664,In_668,In_681);
nor U665 (N_665,N_544,N_36);
and U666 (N_666,N_554,N_86);
nand U667 (N_667,In_308,N_493);
nand U668 (N_668,In_372,In_552);
nand U669 (N_669,N_574,N_542);
or U670 (N_670,N_436,N_279);
nor U671 (N_671,In_954,In_227);
and U672 (N_672,N_262,N_565);
nand U673 (N_673,N_387,N_538);
and U674 (N_674,N_394,N_597);
and U675 (N_675,In_786,N_512);
and U676 (N_676,N_568,In_700);
and U677 (N_677,In_105,N_302);
nand U678 (N_678,N_413,N_426);
or U679 (N_679,In_707,N_576);
nor U680 (N_680,In_775,N_104);
nand U681 (N_681,In_683,N_486);
nor U682 (N_682,In_826,N_559);
and U683 (N_683,In_539,N_370);
and U684 (N_684,N_566,N_267);
or U685 (N_685,In_229,In_887);
or U686 (N_686,N_545,In_425);
nand U687 (N_687,N_399,N_293);
nand U688 (N_688,N_379,N_368);
or U689 (N_689,N_481,N_325);
xnor U690 (N_690,In_986,N_581);
nor U691 (N_691,N_551,N_495);
nor U692 (N_692,In_96,In_15);
nor U693 (N_693,N_564,N_188);
nor U694 (N_694,N_449,N_7);
nand U695 (N_695,In_92,In_535);
nor U696 (N_696,N_307,N_475);
or U697 (N_697,In_967,N_311);
or U698 (N_698,In_879,N_148);
nand U699 (N_699,In_351,In_88);
xor U700 (N_700,N_673,N_533);
nor U701 (N_701,In_942,N_459);
or U702 (N_702,N_555,N_447);
nand U703 (N_703,In_339,In_255);
or U704 (N_704,N_681,In_191);
nand U705 (N_705,N_688,N_136);
and U706 (N_706,In_992,In_252);
and U707 (N_707,N_303,N_537);
and U708 (N_708,N_619,In_595);
and U709 (N_709,In_816,N_116);
nand U710 (N_710,N_438,N_650);
or U711 (N_711,In_452,N_466);
and U712 (N_712,In_386,N_618);
and U713 (N_713,N_432,In_666);
nand U714 (N_714,N_319,N_532);
or U715 (N_715,N_547,N_131);
or U716 (N_716,N_553,N_464);
nor U717 (N_717,N_491,In_567);
xor U718 (N_718,In_346,In_361);
or U719 (N_719,N_407,N_516);
nand U720 (N_720,In_581,N_634);
nor U721 (N_721,N_380,N_642);
and U722 (N_722,N_372,N_490);
nor U723 (N_723,In_2,N_646);
and U724 (N_724,N_691,N_552);
nand U725 (N_725,In_714,N_615);
nor U726 (N_726,N_662,N_220);
or U727 (N_727,In_832,N_674);
nor U728 (N_728,In_422,N_328);
nand U729 (N_729,N_592,N_676);
or U730 (N_730,N_135,N_666);
nand U731 (N_731,N_332,In_404);
nor U732 (N_732,N_456,N_281);
or U733 (N_733,N_664,N_492);
nor U734 (N_734,N_202,In_169);
nand U735 (N_735,N_686,N_683);
and U736 (N_736,N_604,N_343);
nand U737 (N_737,N_571,N_609);
nor U738 (N_738,In_471,N_623);
or U739 (N_739,N_367,N_641);
and U740 (N_740,N_651,N_577);
or U741 (N_741,In_533,N_541);
and U742 (N_742,N_149,N_543);
nand U743 (N_743,In_862,N_667);
nor U744 (N_744,N_520,In_903);
nor U745 (N_745,N_680,In_727);
nand U746 (N_746,N_612,N_526);
or U747 (N_747,N_679,N_661);
or U748 (N_748,N_644,N_639);
or U749 (N_749,N_617,N_462);
and U750 (N_750,N_610,N_626);
xor U751 (N_751,N_483,N_605);
nand U752 (N_752,N_607,In_176);
or U753 (N_753,In_293,N_671);
nand U754 (N_754,N_633,N_603);
nand U755 (N_755,N_694,N_434);
and U756 (N_756,N_285,N_625);
or U757 (N_757,In_922,N_587);
nor U758 (N_758,N_640,N_382);
nand U759 (N_759,N_363,N_685);
or U760 (N_760,N_471,In_282);
and U761 (N_761,N_351,N_628);
and U762 (N_762,N_534,N_110);
and U763 (N_763,N_508,In_463);
nand U764 (N_764,In_9,N_521);
nand U765 (N_765,In_888,N_621);
nand U766 (N_766,N_624,N_347);
or U767 (N_767,N_480,N_652);
and U768 (N_768,In_413,N_697);
and U769 (N_769,N_66,N_572);
nand U770 (N_770,N_357,N_313);
nor U771 (N_771,N_645,N_72);
nor U772 (N_772,N_627,N_529);
nand U773 (N_773,N_270,N_420);
nand U774 (N_774,N_349,In_959);
and U775 (N_775,In_534,N_296);
nand U776 (N_776,N_629,N_591);
and U777 (N_777,N_158,N_658);
nor U778 (N_778,N_698,N_569);
or U779 (N_779,N_657,N_632);
xnor U780 (N_780,N_489,N_678);
and U781 (N_781,N_601,In_51);
nand U782 (N_782,N_246,In_810);
nor U783 (N_783,N_550,In_286);
nand U784 (N_784,N_539,N_692);
xor U785 (N_785,N_659,N_44);
nand U786 (N_786,In_907,N_648);
nor U787 (N_787,N_599,N_696);
or U788 (N_788,N_602,N_689);
or U789 (N_789,N_324,N_595);
nor U790 (N_790,N_677,N_121);
nand U791 (N_791,N_244,N_649);
and U792 (N_792,In_250,N_613);
nor U793 (N_793,N_684,N_643);
or U794 (N_794,In_793,N_608);
or U795 (N_795,N_505,N_556);
and U796 (N_796,N_523,N_322);
nand U797 (N_797,N_630,N_412);
nand U798 (N_798,N_514,N_575);
or U799 (N_799,N_611,N_500);
or U800 (N_800,N_647,N_747);
nand U801 (N_801,In_391,N_782);
nand U802 (N_802,N_230,N_638);
and U803 (N_803,N_783,N_775);
nand U804 (N_804,N_777,N_161);
and U805 (N_805,N_726,In_474);
nand U806 (N_806,N_743,N_718);
and U807 (N_807,N_790,N_561);
nand U808 (N_808,N_248,N_675);
and U809 (N_809,N_797,N_716);
and U810 (N_810,N_762,N_737);
nor U811 (N_811,N_656,N_589);
and U812 (N_812,N_748,N_779);
nand U813 (N_813,In_644,N_636);
and U814 (N_814,N_763,N_750);
or U815 (N_815,N_724,N_240);
nor U816 (N_816,N_706,N_620);
nor U817 (N_817,N_690,N_780);
nand U818 (N_818,In_803,N_798);
nor U819 (N_819,N_655,N_414);
and U820 (N_820,N_732,N_792);
nand U821 (N_821,In_777,N_435);
and U822 (N_822,N_764,N_717);
nand U823 (N_823,In_517,N_614);
nand U824 (N_824,N_725,N_622);
nand U825 (N_825,N_665,N_785);
or U826 (N_826,In_924,N_693);
nor U827 (N_827,In_646,In_789);
and U828 (N_828,N_517,N_653);
nand U829 (N_829,N_540,N_712);
nand U830 (N_830,N_687,N_768);
nor U831 (N_831,N_73,N_429);
nand U832 (N_832,N_588,N_469);
nand U833 (N_833,N_531,In_126);
and U834 (N_834,N_269,N_637);
and U835 (N_835,N_507,In_335);
nor U836 (N_836,N_769,N_433);
nand U837 (N_837,N_733,N_739);
nand U838 (N_838,N_371,N_746);
and U839 (N_839,N_546,N_713);
nor U840 (N_840,N_585,N_669);
and U841 (N_841,N_12,N_699);
and U842 (N_842,N_668,N_794);
or U843 (N_843,In_323,N_710);
nor U844 (N_844,N_715,In_488);
nor U845 (N_845,N_789,N_317);
nor U846 (N_846,N_793,In_318);
nand U847 (N_847,N_767,N_345);
or U848 (N_848,In_129,N_403);
nor U849 (N_849,N_719,N_761);
or U850 (N_850,N_722,N_773);
or U851 (N_851,N_730,In_324);
nand U852 (N_852,N_787,N_720);
and U853 (N_853,N_738,In_248);
nand U854 (N_854,N_616,N_654);
or U855 (N_855,N_741,N_759);
and U856 (N_856,N_771,N_781);
nand U857 (N_857,In_160,N_765);
nand U858 (N_858,N_776,N_742);
or U859 (N_859,N_590,N_749);
nand U860 (N_860,N_714,N_703);
nand U861 (N_861,N_701,N_707);
or U862 (N_862,In_767,N_682);
nor U863 (N_863,N_488,N_734);
and U864 (N_864,N_766,N_736);
and U865 (N_865,N_791,N_711);
and U866 (N_866,N_560,N_727);
nand U867 (N_867,In_193,In_381);
nand U868 (N_868,N_228,In_5);
or U869 (N_869,N_510,N_133);
and U870 (N_870,N_451,In_754);
nor U871 (N_871,N_740,N_731);
and U872 (N_872,N_744,N_702);
and U873 (N_873,N_586,N_729);
or U874 (N_874,N_535,N_670);
nand U875 (N_875,N_756,N_774);
or U876 (N_876,N_753,N_709);
and U877 (N_877,N_663,N_660);
or U878 (N_878,In_550,In_801);
and U879 (N_879,N_723,N_757);
nor U880 (N_880,N_786,In_379);
and U881 (N_881,N_799,N_59);
nand U882 (N_882,N_359,N_755);
nor U883 (N_883,N_784,N_3);
and U884 (N_884,N_631,N_705);
nand U885 (N_885,N_795,N_600);
nor U886 (N_886,N_704,N_796);
or U887 (N_887,N_758,N_760);
and U888 (N_888,N_410,N_524);
or U889 (N_889,N_700,N_728);
nor U890 (N_890,N_672,N_579);
nor U891 (N_891,N_772,N_708);
or U892 (N_892,N_695,N_788);
nand U893 (N_893,N_594,N_752);
or U894 (N_894,N_598,N_754);
or U895 (N_895,N_751,N_504);
or U896 (N_896,N_778,N_770);
nand U897 (N_897,N_745,N_530);
nand U898 (N_898,N_606,N_735);
or U899 (N_899,N_721,N_635);
or U900 (N_900,N_804,N_826);
and U901 (N_901,N_834,N_866);
xnor U902 (N_902,N_878,N_853);
nor U903 (N_903,N_806,N_812);
nor U904 (N_904,N_844,N_801);
or U905 (N_905,N_876,N_899);
and U906 (N_906,N_859,N_820);
nand U907 (N_907,N_847,N_815);
nand U908 (N_908,N_817,N_857);
nor U909 (N_909,N_851,N_884);
nor U910 (N_910,N_809,N_814);
xor U911 (N_911,N_839,N_807);
and U912 (N_912,N_827,N_863);
nor U913 (N_913,N_852,N_808);
and U914 (N_914,N_861,N_842);
nor U915 (N_915,N_886,N_805);
xnor U916 (N_916,N_818,N_836);
and U917 (N_917,N_896,N_832);
and U918 (N_918,N_864,N_854);
xnor U919 (N_919,N_877,N_823);
nand U920 (N_920,N_813,N_870);
or U921 (N_921,N_849,N_858);
nand U922 (N_922,N_895,N_891);
nand U923 (N_923,N_838,N_897);
nand U924 (N_924,N_824,N_888);
nand U925 (N_925,N_872,N_843);
and U926 (N_926,N_883,N_874);
xnor U927 (N_927,N_890,N_892);
nand U928 (N_928,N_810,N_893);
nor U929 (N_929,N_830,N_880);
and U930 (N_930,N_885,N_865);
xor U931 (N_931,N_862,N_837);
nand U932 (N_932,N_831,N_879);
nand U933 (N_933,N_882,N_833);
nand U934 (N_934,N_875,N_828);
nor U935 (N_935,N_869,N_845);
nand U936 (N_936,N_829,N_856);
or U937 (N_937,N_819,N_889);
or U938 (N_938,N_840,N_873);
and U939 (N_939,N_821,N_848);
nand U940 (N_940,N_825,N_898);
nor U941 (N_941,N_816,N_860);
nor U942 (N_942,N_855,N_868);
and U943 (N_943,N_850,N_802);
and U944 (N_944,N_800,N_894);
nand U945 (N_945,N_803,N_811);
and U946 (N_946,N_867,N_835);
nor U947 (N_947,N_871,N_887);
nor U948 (N_948,N_846,N_881);
nand U949 (N_949,N_822,N_841);
nor U950 (N_950,N_815,N_830);
nor U951 (N_951,N_862,N_827);
or U952 (N_952,N_894,N_876);
or U953 (N_953,N_829,N_844);
or U954 (N_954,N_861,N_837);
nor U955 (N_955,N_825,N_841);
nand U956 (N_956,N_839,N_880);
and U957 (N_957,N_899,N_856);
and U958 (N_958,N_875,N_855);
nor U959 (N_959,N_891,N_807);
nor U960 (N_960,N_845,N_890);
nand U961 (N_961,N_895,N_867);
and U962 (N_962,N_813,N_841);
nand U963 (N_963,N_886,N_833);
nor U964 (N_964,N_838,N_867);
nand U965 (N_965,N_837,N_869);
xnor U966 (N_966,N_867,N_863);
and U967 (N_967,N_860,N_843);
and U968 (N_968,N_815,N_803);
nor U969 (N_969,N_837,N_823);
or U970 (N_970,N_842,N_888);
nor U971 (N_971,N_898,N_857);
and U972 (N_972,N_814,N_863);
nand U973 (N_973,N_816,N_844);
nand U974 (N_974,N_808,N_830);
nor U975 (N_975,N_854,N_895);
and U976 (N_976,N_856,N_838);
and U977 (N_977,N_865,N_843);
nor U978 (N_978,N_835,N_802);
nor U979 (N_979,N_891,N_892);
and U980 (N_980,N_862,N_805);
nand U981 (N_981,N_829,N_837);
or U982 (N_982,N_801,N_891);
nor U983 (N_983,N_828,N_855);
nor U984 (N_984,N_865,N_812);
nand U985 (N_985,N_851,N_827);
or U986 (N_986,N_846,N_899);
and U987 (N_987,N_832,N_880);
and U988 (N_988,N_883,N_870);
and U989 (N_989,N_848,N_815);
nand U990 (N_990,N_877,N_832);
and U991 (N_991,N_832,N_887);
nand U992 (N_992,N_852,N_894);
nand U993 (N_993,N_880,N_823);
or U994 (N_994,N_861,N_870);
and U995 (N_995,N_860,N_819);
xor U996 (N_996,N_851,N_847);
nand U997 (N_997,N_820,N_806);
nand U998 (N_998,N_890,N_858);
and U999 (N_999,N_874,N_812);
or U1000 (N_1000,N_935,N_955);
xnor U1001 (N_1001,N_989,N_987);
xor U1002 (N_1002,N_972,N_945);
or U1003 (N_1003,N_940,N_957);
nor U1004 (N_1004,N_963,N_999);
and U1005 (N_1005,N_905,N_934);
or U1006 (N_1006,N_946,N_914);
and U1007 (N_1007,N_931,N_926);
nor U1008 (N_1008,N_920,N_968);
nand U1009 (N_1009,N_921,N_908);
nor U1010 (N_1010,N_936,N_943);
and U1011 (N_1011,N_991,N_982);
and U1012 (N_1012,N_938,N_953);
and U1013 (N_1013,N_964,N_962);
nand U1014 (N_1014,N_924,N_994);
or U1015 (N_1015,N_960,N_928);
and U1016 (N_1016,N_930,N_937);
nand U1017 (N_1017,N_941,N_907);
and U1018 (N_1018,N_958,N_998);
or U1019 (N_1019,N_913,N_912);
nand U1020 (N_1020,N_904,N_971);
nand U1021 (N_1021,N_927,N_922);
nand U1022 (N_1022,N_902,N_978);
or U1023 (N_1023,N_903,N_970);
or U1024 (N_1024,N_967,N_911);
xor U1025 (N_1025,N_980,N_939);
or U1026 (N_1026,N_969,N_929);
nor U1027 (N_1027,N_952,N_944);
and U1028 (N_1028,N_981,N_948);
or U1029 (N_1029,N_950,N_906);
and U1030 (N_1030,N_925,N_974);
nand U1031 (N_1031,N_984,N_995);
nand U1032 (N_1032,N_932,N_933);
and U1033 (N_1033,N_973,N_909);
or U1034 (N_1034,N_992,N_917);
or U1035 (N_1035,N_947,N_956);
or U1036 (N_1036,N_986,N_951);
nand U1037 (N_1037,N_975,N_961);
nor U1038 (N_1038,N_949,N_990);
nand U1039 (N_1039,N_910,N_915);
and U1040 (N_1040,N_993,N_954);
nor U1041 (N_1041,N_900,N_985);
nor U1042 (N_1042,N_923,N_983);
or U1043 (N_1043,N_996,N_979);
and U1044 (N_1044,N_959,N_942);
and U1045 (N_1045,N_966,N_997);
or U1046 (N_1046,N_919,N_916);
and U1047 (N_1047,N_988,N_918);
nand U1048 (N_1048,N_977,N_901);
nand U1049 (N_1049,N_965,N_976);
nand U1050 (N_1050,N_918,N_966);
nor U1051 (N_1051,N_918,N_954);
and U1052 (N_1052,N_904,N_942);
and U1053 (N_1053,N_962,N_922);
or U1054 (N_1054,N_927,N_942);
nor U1055 (N_1055,N_907,N_942);
nand U1056 (N_1056,N_929,N_924);
and U1057 (N_1057,N_946,N_900);
and U1058 (N_1058,N_996,N_940);
nor U1059 (N_1059,N_985,N_908);
and U1060 (N_1060,N_975,N_973);
and U1061 (N_1061,N_973,N_981);
nand U1062 (N_1062,N_913,N_988);
nor U1063 (N_1063,N_964,N_941);
nand U1064 (N_1064,N_927,N_994);
nor U1065 (N_1065,N_942,N_905);
nand U1066 (N_1066,N_978,N_901);
nand U1067 (N_1067,N_933,N_953);
and U1068 (N_1068,N_976,N_920);
and U1069 (N_1069,N_968,N_956);
nor U1070 (N_1070,N_988,N_949);
or U1071 (N_1071,N_909,N_980);
nor U1072 (N_1072,N_971,N_945);
and U1073 (N_1073,N_957,N_973);
and U1074 (N_1074,N_901,N_998);
nand U1075 (N_1075,N_996,N_930);
and U1076 (N_1076,N_903,N_935);
nor U1077 (N_1077,N_991,N_987);
nor U1078 (N_1078,N_932,N_920);
xnor U1079 (N_1079,N_907,N_946);
nand U1080 (N_1080,N_957,N_937);
nand U1081 (N_1081,N_978,N_983);
nor U1082 (N_1082,N_934,N_901);
or U1083 (N_1083,N_986,N_938);
nor U1084 (N_1084,N_922,N_982);
or U1085 (N_1085,N_916,N_909);
or U1086 (N_1086,N_980,N_948);
nor U1087 (N_1087,N_976,N_901);
nand U1088 (N_1088,N_902,N_909);
nand U1089 (N_1089,N_902,N_967);
nand U1090 (N_1090,N_995,N_997);
or U1091 (N_1091,N_973,N_984);
nand U1092 (N_1092,N_933,N_995);
nor U1093 (N_1093,N_974,N_919);
nand U1094 (N_1094,N_972,N_902);
and U1095 (N_1095,N_979,N_928);
or U1096 (N_1096,N_904,N_943);
nor U1097 (N_1097,N_949,N_961);
and U1098 (N_1098,N_921,N_927);
nor U1099 (N_1099,N_939,N_970);
or U1100 (N_1100,N_1043,N_1004);
and U1101 (N_1101,N_1009,N_1090);
or U1102 (N_1102,N_1002,N_1029);
nand U1103 (N_1103,N_1024,N_1019);
nor U1104 (N_1104,N_1008,N_1099);
and U1105 (N_1105,N_1053,N_1007);
or U1106 (N_1106,N_1087,N_1049);
nor U1107 (N_1107,N_1026,N_1015);
nor U1108 (N_1108,N_1094,N_1072);
nor U1109 (N_1109,N_1017,N_1045);
nand U1110 (N_1110,N_1042,N_1073);
nand U1111 (N_1111,N_1016,N_1037);
nand U1112 (N_1112,N_1020,N_1082);
and U1113 (N_1113,N_1050,N_1000);
nor U1114 (N_1114,N_1003,N_1080);
nand U1115 (N_1115,N_1083,N_1071);
nand U1116 (N_1116,N_1051,N_1081);
and U1117 (N_1117,N_1011,N_1010);
nand U1118 (N_1118,N_1091,N_1014);
nand U1119 (N_1119,N_1054,N_1028);
and U1120 (N_1120,N_1034,N_1040);
nand U1121 (N_1121,N_1075,N_1013);
nand U1122 (N_1122,N_1032,N_1077);
nor U1123 (N_1123,N_1060,N_1079);
nor U1124 (N_1124,N_1064,N_1031);
nor U1125 (N_1125,N_1068,N_1027);
or U1126 (N_1126,N_1067,N_1046);
or U1127 (N_1127,N_1089,N_1058);
and U1128 (N_1128,N_1076,N_1063);
nand U1129 (N_1129,N_1059,N_1078);
nand U1130 (N_1130,N_1023,N_1074);
and U1131 (N_1131,N_1012,N_1093);
and U1132 (N_1132,N_1069,N_1039);
nor U1133 (N_1133,N_1036,N_1018);
and U1134 (N_1134,N_1052,N_1088);
or U1135 (N_1135,N_1033,N_1025);
or U1136 (N_1136,N_1055,N_1095);
nand U1137 (N_1137,N_1022,N_1085);
and U1138 (N_1138,N_1061,N_1057);
nand U1139 (N_1139,N_1066,N_1044);
and U1140 (N_1140,N_1097,N_1048);
and U1141 (N_1141,N_1006,N_1056);
and U1142 (N_1142,N_1047,N_1021);
and U1143 (N_1143,N_1092,N_1041);
nor U1144 (N_1144,N_1070,N_1038);
nor U1145 (N_1145,N_1084,N_1086);
nand U1146 (N_1146,N_1098,N_1035);
nand U1147 (N_1147,N_1096,N_1062);
nor U1148 (N_1148,N_1005,N_1030);
nor U1149 (N_1149,N_1001,N_1065);
and U1150 (N_1150,N_1042,N_1017);
and U1151 (N_1151,N_1029,N_1090);
nand U1152 (N_1152,N_1036,N_1074);
nor U1153 (N_1153,N_1096,N_1094);
or U1154 (N_1154,N_1008,N_1078);
and U1155 (N_1155,N_1074,N_1013);
and U1156 (N_1156,N_1044,N_1048);
nor U1157 (N_1157,N_1022,N_1044);
nand U1158 (N_1158,N_1096,N_1055);
nor U1159 (N_1159,N_1084,N_1037);
and U1160 (N_1160,N_1004,N_1026);
nor U1161 (N_1161,N_1002,N_1047);
nor U1162 (N_1162,N_1089,N_1048);
and U1163 (N_1163,N_1081,N_1060);
or U1164 (N_1164,N_1089,N_1031);
and U1165 (N_1165,N_1088,N_1004);
and U1166 (N_1166,N_1058,N_1027);
and U1167 (N_1167,N_1005,N_1043);
nor U1168 (N_1168,N_1023,N_1002);
nand U1169 (N_1169,N_1021,N_1057);
and U1170 (N_1170,N_1042,N_1000);
nor U1171 (N_1171,N_1090,N_1017);
or U1172 (N_1172,N_1086,N_1035);
nor U1173 (N_1173,N_1085,N_1091);
nand U1174 (N_1174,N_1067,N_1019);
and U1175 (N_1175,N_1018,N_1017);
nand U1176 (N_1176,N_1036,N_1073);
nor U1177 (N_1177,N_1038,N_1069);
or U1178 (N_1178,N_1063,N_1006);
and U1179 (N_1179,N_1063,N_1027);
and U1180 (N_1180,N_1051,N_1007);
nand U1181 (N_1181,N_1075,N_1082);
or U1182 (N_1182,N_1078,N_1062);
nand U1183 (N_1183,N_1040,N_1027);
and U1184 (N_1184,N_1083,N_1007);
xnor U1185 (N_1185,N_1006,N_1077);
and U1186 (N_1186,N_1096,N_1022);
or U1187 (N_1187,N_1085,N_1098);
and U1188 (N_1188,N_1011,N_1001);
nand U1189 (N_1189,N_1050,N_1041);
and U1190 (N_1190,N_1038,N_1013);
nor U1191 (N_1191,N_1030,N_1056);
nor U1192 (N_1192,N_1077,N_1013);
nor U1193 (N_1193,N_1021,N_1031);
nor U1194 (N_1194,N_1071,N_1053);
or U1195 (N_1195,N_1044,N_1094);
or U1196 (N_1196,N_1002,N_1019);
nor U1197 (N_1197,N_1070,N_1091);
nand U1198 (N_1198,N_1015,N_1050);
or U1199 (N_1199,N_1039,N_1081);
or U1200 (N_1200,N_1150,N_1137);
nand U1201 (N_1201,N_1169,N_1129);
and U1202 (N_1202,N_1106,N_1153);
and U1203 (N_1203,N_1156,N_1184);
and U1204 (N_1204,N_1182,N_1109);
and U1205 (N_1205,N_1118,N_1114);
xnor U1206 (N_1206,N_1119,N_1177);
or U1207 (N_1207,N_1195,N_1197);
and U1208 (N_1208,N_1194,N_1180);
nor U1209 (N_1209,N_1152,N_1117);
nand U1210 (N_1210,N_1136,N_1105);
or U1211 (N_1211,N_1189,N_1142);
and U1212 (N_1212,N_1173,N_1110);
nand U1213 (N_1213,N_1161,N_1102);
nand U1214 (N_1214,N_1128,N_1123);
xnor U1215 (N_1215,N_1126,N_1146);
and U1216 (N_1216,N_1159,N_1107);
or U1217 (N_1217,N_1187,N_1163);
and U1218 (N_1218,N_1183,N_1155);
and U1219 (N_1219,N_1148,N_1196);
nor U1220 (N_1220,N_1134,N_1141);
or U1221 (N_1221,N_1135,N_1112);
nand U1222 (N_1222,N_1175,N_1113);
nand U1223 (N_1223,N_1143,N_1190);
nand U1224 (N_1224,N_1132,N_1198);
and U1225 (N_1225,N_1125,N_1160);
nor U1226 (N_1226,N_1104,N_1166);
and U1227 (N_1227,N_1101,N_1178);
nand U1228 (N_1228,N_1124,N_1199);
nor U1229 (N_1229,N_1191,N_1120);
or U1230 (N_1230,N_1140,N_1192);
nor U1231 (N_1231,N_1176,N_1122);
nor U1232 (N_1232,N_1144,N_1103);
nand U1233 (N_1233,N_1147,N_1158);
and U1234 (N_1234,N_1130,N_1174);
nand U1235 (N_1235,N_1164,N_1127);
nand U1236 (N_1236,N_1149,N_1165);
and U1237 (N_1237,N_1138,N_1186);
nor U1238 (N_1238,N_1172,N_1139);
and U1239 (N_1239,N_1193,N_1131);
nor U1240 (N_1240,N_1170,N_1133);
and U1241 (N_1241,N_1121,N_1108);
or U1242 (N_1242,N_1157,N_1188);
or U1243 (N_1243,N_1116,N_1181);
or U1244 (N_1244,N_1179,N_1167);
nand U1245 (N_1245,N_1168,N_1100);
and U1246 (N_1246,N_1145,N_1185);
nor U1247 (N_1247,N_1115,N_1171);
or U1248 (N_1248,N_1151,N_1154);
and U1249 (N_1249,N_1111,N_1162);
xnor U1250 (N_1250,N_1187,N_1141);
or U1251 (N_1251,N_1145,N_1120);
nand U1252 (N_1252,N_1121,N_1166);
and U1253 (N_1253,N_1198,N_1157);
and U1254 (N_1254,N_1160,N_1190);
or U1255 (N_1255,N_1186,N_1160);
or U1256 (N_1256,N_1177,N_1127);
and U1257 (N_1257,N_1101,N_1183);
or U1258 (N_1258,N_1175,N_1164);
nor U1259 (N_1259,N_1147,N_1169);
nand U1260 (N_1260,N_1165,N_1127);
and U1261 (N_1261,N_1148,N_1124);
nor U1262 (N_1262,N_1176,N_1151);
nand U1263 (N_1263,N_1119,N_1132);
or U1264 (N_1264,N_1109,N_1187);
or U1265 (N_1265,N_1142,N_1176);
and U1266 (N_1266,N_1112,N_1196);
or U1267 (N_1267,N_1118,N_1179);
or U1268 (N_1268,N_1111,N_1169);
or U1269 (N_1269,N_1150,N_1108);
nor U1270 (N_1270,N_1166,N_1193);
nand U1271 (N_1271,N_1167,N_1195);
nand U1272 (N_1272,N_1148,N_1134);
nand U1273 (N_1273,N_1169,N_1101);
nor U1274 (N_1274,N_1195,N_1115);
nor U1275 (N_1275,N_1164,N_1187);
nor U1276 (N_1276,N_1162,N_1108);
nand U1277 (N_1277,N_1107,N_1199);
nand U1278 (N_1278,N_1169,N_1137);
nor U1279 (N_1279,N_1178,N_1115);
nand U1280 (N_1280,N_1170,N_1102);
or U1281 (N_1281,N_1112,N_1107);
nor U1282 (N_1282,N_1164,N_1167);
and U1283 (N_1283,N_1119,N_1134);
or U1284 (N_1284,N_1190,N_1179);
xnor U1285 (N_1285,N_1198,N_1131);
nor U1286 (N_1286,N_1123,N_1108);
nand U1287 (N_1287,N_1155,N_1198);
nand U1288 (N_1288,N_1138,N_1128);
nor U1289 (N_1289,N_1148,N_1164);
or U1290 (N_1290,N_1119,N_1121);
xor U1291 (N_1291,N_1111,N_1191);
nor U1292 (N_1292,N_1185,N_1176);
nor U1293 (N_1293,N_1135,N_1138);
or U1294 (N_1294,N_1121,N_1147);
and U1295 (N_1295,N_1157,N_1125);
nand U1296 (N_1296,N_1101,N_1119);
nand U1297 (N_1297,N_1171,N_1173);
nor U1298 (N_1298,N_1132,N_1160);
nor U1299 (N_1299,N_1142,N_1175);
nor U1300 (N_1300,N_1272,N_1260);
or U1301 (N_1301,N_1242,N_1236);
and U1302 (N_1302,N_1227,N_1281);
and U1303 (N_1303,N_1238,N_1234);
and U1304 (N_1304,N_1254,N_1252);
or U1305 (N_1305,N_1244,N_1228);
nor U1306 (N_1306,N_1299,N_1226);
and U1307 (N_1307,N_1231,N_1294);
xnor U1308 (N_1308,N_1213,N_1205);
or U1309 (N_1309,N_1290,N_1284);
or U1310 (N_1310,N_1298,N_1249);
and U1311 (N_1311,N_1258,N_1202);
nor U1312 (N_1312,N_1225,N_1235);
and U1313 (N_1313,N_1223,N_1253);
nand U1314 (N_1314,N_1207,N_1212);
and U1315 (N_1315,N_1275,N_1243);
and U1316 (N_1316,N_1206,N_1222);
nor U1317 (N_1317,N_1224,N_1204);
xor U1318 (N_1318,N_1285,N_1218);
and U1319 (N_1319,N_1266,N_1269);
nor U1320 (N_1320,N_1240,N_1229);
nand U1321 (N_1321,N_1246,N_1289);
and U1322 (N_1322,N_1201,N_1247);
nor U1323 (N_1323,N_1257,N_1248);
or U1324 (N_1324,N_1276,N_1220);
nor U1325 (N_1325,N_1268,N_1209);
nand U1326 (N_1326,N_1297,N_1283);
and U1327 (N_1327,N_1288,N_1286);
nand U1328 (N_1328,N_1291,N_1264);
and U1329 (N_1329,N_1200,N_1278);
nor U1330 (N_1330,N_1219,N_1265);
nor U1331 (N_1331,N_1263,N_1279);
and U1332 (N_1332,N_1261,N_1282);
nor U1333 (N_1333,N_1255,N_1280);
and U1334 (N_1334,N_1262,N_1295);
xnor U1335 (N_1335,N_1274,N_1251);
nor U1336 (N_1336,N_1277,N_1250);
nor U1337 (N_1337,N_1256,N_1259);
nor U1338 (N_1338,N_1214,N_1267);
and U1339 (N_1339,N_1296,N_1203);
nand U1340 (N_1340,N_1287,N_1230);
nand U1341 (N_1341,N_1273,N_1239);
and U1342 (N_1342,N_1210,N_1241);
and U1343 (N_1343,N_1217,N_1292);
or U1344 (N_1344,N_1221,N_1270);
and U1345 (N_1345,N_1215,N_1233);
nor U1346 (N_1346,N_1237,N_1216);
or U1347 (N_1347,N_1271,N_1211);
or U1348 (N_1348,N_1245,N_1232);
nor U1349 (N_1349,N_1208,N_1293);
xnor U1350 (N_1350,N_1238,N_1229);
nand U1351 (N_1351,N_1262,N_1202);
nand U1352 (N_1352,N_1289,N_1226);
or U1353 (N_1353,N_1273,N_1298);
nor U1354 (N_1354,N_1225,N_1288);
or U1355 (N_1355,N_1289,N_1206);
and U1356 (N_1356,N_1250,N_1241);
and U1357 (N_1357,N_1246,N_1288);
or U1358 (N_1358,N_1222,N_1249);
nand U1359 (N_1359,N_1288,N_1222);
nor U1360 (N_1360,N_1222,N_1239);
nand U1361 (N_1361,N_1262,N_1266);
nor U1362 (N_1362,N_1260,N_1274);
and U1363 (N_1363,N_1243,N_1244);
and U1364 (N_1364,N_1279,N_1202);
and U1365 (N_1365,N_1277,N_1236);
or U1366 (N_1366,N_1252,N_1280);
or U1367 (N_1367,N_1249,N_1279);
xor U1368 (N_1368,N_1239,N_1200);
nor U1369 (N_1369,N_1287,N_1234);
or U1370 (N_1370,N_1274,N_1269);
nand U1371 (N_1371,N_1258,N_1227);
or U1372 (N_1372,N_1257,N_1261);
nor U1373 (N_1373,N_1256,N_1265);
and U1374 (N_1374,N_1221,N_1205);
or U1375 (N_1375,N_1200,N_1247);
nor U1376 (N_1376,N_1250,N_1276);
xor U1377 (N_1377,N_1267,N_1228);
nor U1378 (N_1378,N_1291,N_1239);
nand U1379 (N_1379,N_1246,N_1276);
or U1380 (N_1380,N_1248,N_1267);
nand U1381 (N_1381,N_1230,N_1282);
and U1382 (N_1382,N_1228,N_1236);
and U1383 (N_1383,N_1235,N_1215);
nor U1384 (N_1384,N_1247,N_1216);
nor U1385 (N_1385,N_1226,N_1293);
nand U1386 (N_1386,N_1268,N_1243);
nor U1387 (N_1387,N_1204,N_1262);
and U1388 (N_1388,N_1238,N_1276);
nor U1389 (N_1389,N_1282,N_1256);
or U1390 (N_1390,N_1215,N_1217);
nand U1391 (N_1391,N_1235,N_1290);
or U1392 (N_1392,N_1210,N_1217);
nand U1393 (N_1393,N_1229,N_1281);
nand U1394 (N_1394,N_1220,N_1225);
and U1395 (N_1395,N_1246,N_1224);
or U1396 (N_1396,N_1272,N_1265);
nand U1397 (N_1397,N_1227,N_1205);
and U1398 (N_1398,N_1217,N_1203);
xor U1399 (N_1399,N_1203,N_1216);
nor U1400 (N_1400,N_1393,N_1365);
nand U1401 (N_1401,N_1397,N_1372);
and U1402 (N_1402,N_1359,N_1399);
nor U1403 (N_1403,N_1392,N_1317);
or U1404 (N_1404,N_1394,N_1389);
or U1405 (N_1405,N_1322,N_1374);
nand U1406 (N_1406,N_1324,N_1315);
nand U1407 (N_1407,N_1368,N_1348);
nand U1408 (N_1408,N_1351,N_1302);
nor U1409 (N_1409,N_1335,N_1371);
nor U1410 (N_1410,N_1316,N_1307);
nor U1411 (N_1411,N_1332,N_1308);
nand U1412 (N_1412,N_1391,N_1354);
nand U1413 (N_1413,N_1367,N_1369);
or U1414 (N_1414,N_1344,N_1336);
and U1415 (N_1415,N_1396,N_1349);
and U1416 (N_1416,N_1370,N_1343);
and U1417 (N_1417,N_1323,N_1358);
and U1418 (N_1418,N_1366,N_1310);
or U1419 (N_1419,N_1311,N_1360);
and U1420 (N_1420,N_1363,N_1353);
and U1421 (N_1421,N_1352,N_1319);
or U1422 (N_1422,N_1334,N_1320);
or U1423 (N_1423,N_1395,N_1330);
nor U1424 (N_1424,N_1381,N_1305);
or U1425 (N_1425,N_1340,N_1333);
or U1426 (N_1426,N_1314,N_1312);
and U1427 (N_1427,N_1376,N_1357);
nor U1428 (N_1428,N_1345,N_1300);
nor U1429 (N_1429,N_1385,N_1398);
and U1430 (N_1430,N_1380,N_1388);
or U1431 (N_1431,N_1378,N_1346);
nand U1432 (N_1432,N_1341,N_1306);
nand U1433 (N_1433,N_1364,N_1304);
nor U1434 (N_1434,N_1362,N_1375);
and U1435 (N_1435,N_1301,N_1325);
nand U1436 (N_1436,N_1321,N_1356);
nand U1437 (N_1437,N_1309,N_1318);
or U1438 (N_1438,N_1384,N_1303);
or U1439 (N_1439,N_1390,N_1350);
and U1440 (N_1440,N_1327,N_1387);
nor U1441 (N_1441,N_1377,N_1337);
and U1442 (N_1442,N_1382,N_1326);
nor U1443 (N_1443,N_1338,N_1328);
and U1444 (N_1444,N_1383,N_1331);
or U1445 (N_1445,N_1373,N_1361);
nand U1446 (N_1446,N_1339,N_1347);
or U1447 (N_1447,N_1313,N_1386);
or U1448 (N_1448,N_1342,N_1379);
nor U1449 (N_1449,N_1329,N_1355);
or U1450 (N_1450,N_1314,N_1387);
and U1451 (N_1451,N_1386,N_1357);
or U1452 (N_1452,N_1303,N_1371);
and U1453 (N_1453,N_1388,N_1305);
and U1454 (N_1454,N_1392,N_1308);
and U1455 (N_1455,N_1348,N_1374);
or U1456 (N_1456,N_1327,N_1399);
or U1457 (N_1457,N_1355,N_1318);
or U1458 (N_1458,N_1319,N_1337);
or U1459 (N_1459,N_1353,N_1313);
or U1460 (N_1460,N_1349,N_1383);
or U1461 (N_1461,N_1362,N_1309);
nand U1462 (N_1462,N_1347,N_1308);
nand U1463 (N_1463,N_1326,N_1306);
and U1464 (N_1464,N_1386,N_1332);
nor U1465 (N_1465,N_1399,N_1328);
nand U1466 (N_1466,N_1318,N_1340);
or U1467 (N_1467,N_1307,N_1309);
nand U1468 (N_1468,N_1325,N_1350);
nand U1469 (N_1469,N_1322,N_1324);
nand U1470 (N_1470,N_1333,N_1395);
nor U1471 (N_1471,N_1321,N_1389);
and U1472 (N_1472,N_1361,N_1358);
nand U1473 (N_1473,N_1309,N_1351);
nand U1474 (N_1474,N_1359,N_1391);
or U1475 (N_1475,N_1396,N_1334);
or U1476 (N_1476,N_1323,N_1301);
nor U1477 (N_1477,N_1356,N_1341);
nor U1478 (N_1478,N_1382,N_1349);
or U1479 (N_1479,N_1337,N_1333);
xnor U1480 (N_1480,N_1359,N_1372);
or U1481 (N_1481,N_1371,N_1323);
and U1482 (N_1482,N_1385,N_1360);
nand U1483 (N_1483,N_1379,N_1343);
and U1484 (N_1484,N_1359,N_1351);
and U1485 (N_1485,N_1342,N_1319);
nor U1486 (N_1486,N_1385,N_1322);
nor U1487 (N_1487,N_1335,N_1317);
or U1488 (N_1488,N_1393,N_1362);
and U1489 (N_1489,N_1386,N_1392);
nand U1490 (N_1490,N_1321,N_1302);
xnor U1491 (N_1491,N_1327,N_1313);
and U1492 (N_1492,N_1312,N_1327);
nor U1493 (N_1493,N_1379,N_1397);
nand U1494 (N_1494,N_1332,N_1337);
and U1495 (N_1495,N_1368,N_1358);
and U1496 (N_1496,N_1340,N_1334);
nand U1497 (N_1497,N_1349,N_1321);
nor U1498 (N_1498,N_1307,N_1388);
nor U1499 (N_1499,N_1312,N_1359);
xnor U1500 (N_1500,N_1428,N_1406);
and U1501 (N_1501,N_1401,N_1438);
and U1502 (N_1502,N_1404,N_1411);
and U1503 (N_1503,N_1444,N_1471);
or U1504 (N_1504,N_1493,N_1446);
nor U1505 (N_1505,N_1447,N_1482);
and U1506 (N_1506,N_1451,N_1449);
nor U1507 (N_1507,N_1488,N_1454);
nor U1508 (N_1508,N_1407,N_1494);
nor U1509 (N_1509,N_1417,N_1486);
and U1510 (N_1510,N_1436,N_1437);
nor U1511 (N_1511,N_1485,N_1459);
nand U1512 (N_1512,N_1418,N_1467);
nand U1513 (N_1513,N_1452,N_1443);
or U1514 (N_1514,N_1435,N_1415);
or U1515 (N_1515,N_1472,N_1490);
nand U1516 (N_1516,N_1463,N_1480);
or U1517 (N_1517,N_1461,N_1403);
or U1518 (N_1518,N_1483,N_1464);
or U1519 (N_1519,N_1413,N_1432);
nor U1520 (N_1520,N_1455,N_1400);
nand U1521 (N_1521,N_1499,N_1450);
and U1522 (N_1522,N_1465,N_1495);
nand U1523 (N_1523,N_1429,N_1478);
xor U1524 (N_1524,N_1422,N_1484);
or U1525 (N_1525,N_1414,N_1434);
nor U1526 (N_1526,N_1445,N_1416);
nand U1527 (N_1527,N_1466,N_1410);
nor U1528 (N_1528,N_1473,N_1412);
xor U1529 (N_1529,N_1409,N_1456);
nor U1530 (N_1530,N_1421,N_1408);
or U1531 (N_1531,N_1439,N_1491);
and U1532 (N_1532,N_1487,N_1427);
or U1533 (N_1533,N_1497,N_1453);
or U1534 (N_1534,N_1460,N_1423);
nand U1535 (N_1535,N_1492,N_1479);
nor U1536 (N_1536,N_1468,N_1405);
xnor U1537 (N_1537,N_1470,N_1474);
nor U1538 (N_1538,N_1425,N_1433);
or U1539 (N_1539,N_1477,N_1426);
and U1540 (N_1540,N_1442,N_1448);
nand U1541 (N_1541,N_1420,N_1440);
or U1542 (N_1542,N_1424,N_1419);
and U1543 (N_1543,N_1458,N_1462);
nand U1544 (N_1544,N_1475,N_1431);
or U1545 (N_1545,N_1481,N_1476);
or U1546 (N_1546,N_1496,N_1498);
nand U1547 (N_1547,N_1402,N_1457);
nor U1548 (N_1548,N_1489,N_1441);
nor U1549 (N_1549,N_1469,N_1430);
nand U1550 (N_1550,N_1447,N_1410);
nand U1551 (N_1551,N_1443,N_1459);
or U1552 (N_1552,N_1417,N_1401);
nor U1553 (N_1553,N_1481,N_1460);
and U1554 (N_1554,N_1406,N_1413);
nor U1555 (N_1555,N_1428,N_1468);
and U1556 (N_1556,N_1471,N_1448);
nand U1557 (N_1557,N_1496,N_1400);
and U1558 (N_1558,N_1435,N_1402);
nor U1559 (N_1559,N_1418,N_1446);
nor U1560 (N_1560,N_1472,N_1475);
nor U1561 (N_1561,N_1450,N_1455);
nor U1562 (N_1562,N_1490,N_1437);
and U1563 (N_1563,N_1478,N_1450);
or U1564 (N_1564,N_1436,N_1440);
nor U1565 (N_1565,N_1441,N_1412);
or U1566 (N_1566,N_1429,N_1442);
and U1567 (N_1567,N_1485,N_1448);
nor U1568 (N_1568,N_1462,N_1498);
and U1569 (N_1569,N_1493,N_1461);
nor U1570 (N_1570,N_1493,N_1464);
and U1571 (N_1571,N_1446,N_1481);
or U1572 (N_1572,N_1487,N_1479);
or U1573 (N_1573,N_1422,N_1459);
and U1574 (N_1574,N_1453,N_1456);
nor U1575 (N_1575,N_1449,N_1495);
and U1576 (N_1576,N_1413,N_1400);
or U1577 (N_1577,N_1478,N_1414);
nor U1578 (N_1578,N_1455,N_1475);
nor U1579 (N_1579,N_1404,N_1499);
or U1580 (N_1580,N_1440,N_1435);
and U1581 (N_1581,N_1456,N_1497);
nand U1582 (N_1582,N_1406,N_1436);
and U1583 (N_1583,N_1430,N_1438);
nand U1584 (N_1584,N_1493,N_1467);
nor U1585 (N_1585,N_1445,N_1415);
and U1586 (N_1586,N_1432,N_1436);
nand U1587 (N_1587,N_1485,N_1425);
or U1588 (N_1588,N_1409,N_1458);
or U1589 (N_1589,N_1480,N_1450);
nand U1590 (N_1590,N_1444,N_1493);
or U1591 (N_1591,N_1437,N_1430);
and U1592 (N_1592,N_1415,N_1438);
nor U1593 (N_1593,N_1496,N_1415);
nor U1594 (N_1594,N_1445,N_1468);
nand U1595 (N_1595,N_1420,N_1449);
nand U1596 (N_1596,N_1407,N_1446);
or U1597 (N_1597,N_1495,N_1401);
nor U1598 (N_1598,N_1478,N_1432);
and U1599 (N_1599,N_1477,N_1428);
nor U1600 (N_1600,N_1557,N_1526);
nand U1601 (N_1601,N_1536,N_1569);
or U1602 (N_1602,N_1590,N_1556);
nor U1603 (N_1603,N_1598,N_1525);
nor U1604 (N_1604,N_1563,N_1530);
or U1605 (N_1605,N_1517,N_1550);
nand U1606 (N_1606,N_1565,N_1549);
and U1607 (N_1607,N_1580,N_1593);
nand U1608 (N_1608,N_1578,N_1513);
and U1609 (N_1609,N_1551,N_1523);
or U1610 (N_1610,N_1524,N_1540);
nand U1611 (N_1611,N_1559,N_1576);
nor U1612 (N_1612,N_1543,N_1542);
nor U1613 (N_1613,N_1555,N_1511);
nor U1614 (N_1614,N_1588,N_1591);
and U1615 (N_1615,N_1509,N_1500);
and U1616 (N_1616,N_1561,N_1599);
nor U1617 (N_1617,N_1594,N_1586);
nor U1618 (N_1618,N_1538,N_1582);
and U1619 (N_1619,N_1583,N_1539);
nor U1620 (N_1620,N_1515,N_1546);
nor U1621 (N_1621,N_1537,N_1579);
or U1622 (N_1622,N_1519,N_1584);
nor U1623 (N_1623,N_1572,N_1568);
xor U1624 (N_1624,N_1544,N_1558);
or U1625 (N_1625,N_1512,N_1547);
and U1626 (N_1626,N_1554,N_1552);
or U1627 (N_1627,N_1507,N_1592);
or U1628 (N_1628,N_1520,N_1529);
and U1629 (N_1629,N_1506,N_1531);
nand U1630 (N_1630,N_1570,N_1503);
nand U1631 (N_1631,N_1566,N_1502);
nand U1632 (N_1632,N_1535,N_1587);
nand U1633 (N_1633,N_1527,N_1514);
or U1634 (N_1634,N_1585,N_1510);
nor U1635 (N_1635,N_1571,N_1589);
and U1636 (N_1636,N_1581,N_1567);
and U1637 (N_1637,N_1516,N_1553);
nand U1638 (N_1638,N_1505,N_1595);
nor U1639 (N_1639,N_1508,N_1528);
and U1640 (N_1640,N_1574,N_1532);
and U1641 (N_1641,N_1560,N_1575);
nor U1642 (N_1642,N_1518,N_1562);
or U1643 (N_1643,N_1521,N_1504);
and U1644 (N_1644,N_1534,N_1545);
nand U1645 (N_1645,N_1596,N_1573);
or U1646 (N_1646,N_1533,N_1541);
or U1647 (N_1647,N_1501,N_1522);
or U1648 (N_1648,N_1564,N_1548);
or U1649 (N_1649,N_1577,N_1597);
and U1650 (N_1650,N_1588,N_1573);
or U1651 (N_1651,N_1576,N_1512);
and U1652 (N_1652,N_1562,N_1542);
and U1653 (N_1653,N_1535,N_1519);
nand U1654 (N_1654,N_1574,N_1520);
or U1655 (N_1655,N_1548,N_1536);
or U1656 (N_1656,N_1508,N_1584);
and U1657 (N_1657,N_1581,N_1593);
nor U1658 (N_1658,N_1595,N_1545);
nor U1659 (N_1659,N_1540,N_1590);
nor U1660 (N_1660,N_1515,N_1514);
nor U1661 (N_1661,N_1500,N_1556);
or U1662 (N_1662,N_1523,N_1557);
nand U1663 (N_1663,N_1551,N_1557);
and U1664 (N_1664,N_1505,N_1583);
nor U1665 (N_1665,N_1553,N_1559);
nand U1666 (N_1666,N_1562,N_1525);
and U1667 (N_1667,N_1505,N_1594);
and U1668 (N_1668,N_1518,N_1550);
nor U1669 (N_1669,N_1566,N_1521);
or U1670 (N_1670,N_1531,N_1563);
nor U1671 (N_1671,N_1524,N_1545);
nor U1672 (N_1672,N_1596,N_1560);
or U1673 (N_1673,N_1519,N_1580);
and U1674 (N_1674,N_1546,N_1562);
or U1675 (N_1675,N_1597,N_1510);
nand U1676 (N_1676,N_1500,N_1505);
nor U1677 (N_1677,N_1522,N_1534);
nor U1678 (N_1678,N_1593,N_1569);
and U1679 (N_1679,N_1510,N_1522);
and U1680 (N_1680,N_1545,N_1516);
and U1681 (N_1681,N_1522,N_1560);
or U1682 (N_1682,N_1530,N_1534);
and U1683 (N_1683,N_1541,N_1593);
or U1684 (N_1684,N_1589,N_1585);
or U1685 (N_1685,N_1577,N_1587);
or U1686 (N_1686,N_1553,N_1539);
nor U1687 (N_1687,N_1577,N_1551);
or U1688 (N_1688,N_1591,N_1549);
and U1689 (N_1689,N_1558,N_1557);
and U1690 (N_1690,N_1544,N_1529);
nand U1691 (N_1691,N_1553,N_1555);
and U1692 (N_1692,N_1511,N_1592);
and U1693 (N_1693,N_1506,N_1523);
nor U1694 (N_1694,N_1583,N_1578);
xor U1695 (N_1695,N_1573,N_1589);
and U1696 (N_1696,N_1586,N_1562);
or U1697 (N_1697,N_1509,N_1574);
nand U1698 (N_1698,N_1500,N_1585);
and U1699 (N_1699,N_1544,N_1520);
nor U1700 (N_1700,N_1681,N_1659);
nor U1701 (N_1701,N_1615,N_1637);
nand U1702 (N_1702,N_1635,N_1638);
or U1703 (N_1703,N_1607,N_1612);
nand U1704 (N_1704,N_1668,N_1621);
nand U1705 (N_1705,N_1649,N_1682);
nor U1706 (N_1706,N_1632,N_1611);
nand U1707 (N_1707,N_1650,N_1605);
and U1708 (N_1708,N_1695,N_1680);
nor U1709 (N_1709,N_1608,N_1692);
and U1710 (N_1710,N_1620,N_1656);
xor U1711 (N_1711,N_1662,N_1685);
nor U1712 (N_1712,N_1669,N_1660);
nand U1713 (N_1713,N_1661,N_1636);
nand U1714 (N_1714,N_1600,N_1625);
nand U1715 (N_1715,N_1653,N_1672);
or U1716 (N_1716,N_1698,N_1618);
or U1717 (N_1717,N_1679,N_1694);
nor U1718 (N_1718,N_1642,N_1699);
nor U1719 (N_1719,N_1604,N_1671);
and U1720 (N_1720,N_1657,N_1691);
and U1721 (N_1721,N_1696,N_1693);
nor U1722 (N_1722,N_1687,N_1655);
or U1723 (N_1723,N_1676,N_1629);
nand U1724 (N_1724,N_1627,N_1675);
or U1725 (N_1725,N_1648,N_1614);
nor U1726 (N_1726,N_1677,N_1644);
and U1727 (N_1727,N_1643,N_1664);
or U1728 (N_1728,N_1678,N_1623);
and U1729 (N_1729,N_1686,N_1603);
nand U1730 (N_1730,N_1606,N_1613);
and U1731 (N_1731,N_1652,N_1633);
nand U1732 (N_1732,N_1658,N_1651);
or U1733 (N_1733,N_1631,N_1690);
nor U1734 (N_1734,N_1639,N_1602);
or U1735 (N_1735,N_1647,N_1684);
nor U1736 (N_1736,N_1674,N_1641);
nand U1737 (N_1737,N_1624,N_1610);
and U1738 (N_1738,N_1688,N_1628);
nand U1739 (N_1739,N_1673,N_1645);
and U1740 (N_1740,N_1663,N_1667);
and U1741 (N_1741,N_1665,N_1640);
or U1742 (N_1742,N_1601,N_1616);
nand U1743 (N_1743,N_1609,N_1670);
or U1744 (N_1744,N_1654,N_1617);
nand U1745 (N_1745,N_1697,N_1622);
and U1746 (N_1746,N_1646,N_1689);
nor U1747 (N_1747,N_1630,N_1619);
and U1748 (N_1748,N_1634,N_1683);
and U1749 (N_1749,N_1666,N_1626);
nor U1750 (N_1750,N_1614,N_1654);
nand U1751 (N_1751,N_1698,N_1629);
nand U1752 (N_1752,N_1656,N_1629);
nor U1753 (N_1753,N_1600,N_1697);
or U1754 (N_1754,N_1665,N_1693);
nand U1755 (N_1755,N_1632,N_1606);
or U1756 (N_1756,N_1649,N_1687);
or U1757 (N_1757,N_1662,N_1670);
nand U1758 (N_1758,N_1608,N_1676);
nand U1759 (N_1759,N_1696,N_1692);
nand U1760 (N_1760,N_1693,N_1609);
or U1761 (N_1761,N_1675,N_1666);
nand U1762 (N_1762,N_1607,N_1671);
nand U1763 (N_1763,N_1629,N_1630);
nor U1764 (N_1764,N_1680,N_1638);
or U1765 (N_1765,N_1639,N_1614);
nand U1766 (N_1766,N_1664,N_1630);
nor U1767 (N_1767,N_1690,N_1609);
or U1768 (N_1768,N_1684,N_1622);
nor U1769 (N_1769,N_1647,N_1633);
or U1770 (N_1770,N_1609,N_1652);
or U1771 (N_1771,N_1600,N_1688);
or U1772 (N_1772,N_1612,N_1684);
and U1773 (N_1773,N_1620,N_1621);
xnor U1774 (N_1774,N_1630,N_1642);
or U1775 (N_1775,N_1604,N_1621);
and U1776 (N_1776,N_1671,N_1653);
or U1777 (N_1777,N_1647,N_1615);
and U1778 (N_1778,N_1637,N_1648);
or U1779 (N_1779,N_1649,N_1677);
or U1780 (N_1780,N_1679,N_1618);
and U1781 (N_1781,N_1658,N_1674);
xnor U1782 (N_1782,N_1600,N_1689);
or U1783 (N_1783,N_1623,N_1654);
or U1784 (N_1784,N_1646,N_1657);
or U1785 (N_1785,N_1678,N_1672);
nor U1786 (N_1786,N_1609,N_1691);
and U1787 (N_1787,N_1619,N_1624);
or U1788 (N_1788,N_1629,N_1686);
or U1789 (N_1789,N_1666,N_1672);
nand U1790 (N_1790,N_1665,N_1681);
or U1791 (N_1791,N_1667,N_1630);
and U1792 (N_1792,N_1614,N_1604);
nor U1793 (N_1793,N_1628,N_1613);
nor U1794 (N_1794,N_1691,N_1673);
nand U1795 (N_1795,N_1604,N_1686);
and U1796 (N_1796,N_1633,N_1675);
or U1797 (N_1797,N_1694,N_1619);
or U1798 (N_1798,N_1631,N_1627);
nand U1799 (N_1799,N_1632,N_1600);
nor U1800 (N_1800,N_1795,N_1748);
or U1801 (N_1801,N_1756,N_1737);
or U1802 (N_1802,N_1776,N_1774);
or U1803 (N_1803,N_1762,N_1719);
nand U1804 (N_1804,N_1751,N_1742);
nor U1805 (N_1805,N_1732,N_1796);
nor U1806 (N_1806,N_1726,N_1786);
xor U1807 (N_1807,N_1703,N_1701);
xor U1808 (N_1808,N_1713,N_1799);
or U1809 (N_1809,N_1790,N_1782);
or U1810 (N_1810,N_1753,N_1708);
nand U1811 (N_1811,N_1768,N_1746);
nor U1812 (N_1812,N_1760,N_1764);
and U1813 (N_1813,N_1789,N_1715);
nand U1814 (N_1814,N_1787,N_1709);
nor U1815 (N_1815,N_1717,N_1705);
or U1816 (N_1816,N_1712,N_1783);
nand U1817 (N_1817,N_1793,N_1788);
nor U1818 (N_1818,N_1711,N_1725);
and U1819 (N_1819,N_1785,N_1765);
nor U1820 (N_1820,N_1754,N_1707);
or U1821 (N_1821,N_1733,N_1759);
and U1822 (N_1822,N_1784,N_1700);
or U1823 (N_1823,N_1743,N_1797);
nor U1824 (N_1824,N_1798,N_1763);
or U1825 (N_1825,N_1720,N_1724);
and U1826 (N_1826,N_1739,N_1749);
or U1827 (N_1827,N_1716,N_1738);
and U1828 (N_1828,N_1704,N_1791);
nand U1829 (N_1829,N_1710,N_1777);
and U1830 (N_1830,N_1731,N_1730);
or U1831 (N_1831,N_1778,N_1767);
and U1832 (N_1832,N_1781,N_1727);
nor U1833 (N_1833,N_1714,N_1750);
nand U1834 (N_1834,N_1757,N_1747);
or U1835 (N_1835,N_1758,N_1766);
and U1836 (N_1836,N_1761,N_1773);
nand U1837 (N_1837,N_1741,N_1735);
nand U1838 (N_1838,N_1734,N_1772);
nor U1839 (N_1839,N_1718,N_1792);
nand U1840 (N_1840,N_1775,N_1779);
or U1841 (N_1841,N_1794,N_1736);
nor U1842 (N_1842,N_1721,N_1752);
or U1843 (N_1843,N_1780,N_1744);
nor U1844 (N_1844,N_1728,N_1723);
nand U1845 (N_1845,N_1771,N_1702);
nand U1846 (N_1846,N_1706,N_1755);
nand U1847 (N_1847,N_1745,N_1769);
and U1848 (N_1848,N_1740,N_1729);
nor U1849 (N_1849,N_1770,N_1722);
and U1850 (N_1850,N_1768,N_1787);
nand U1851 (N_1851,N_1734,N_1751);
nor U1852 (N_1852,N_1786,N_1734);
nand U1853 (N_1853,N_1712,N_1794);
nand U1854 (N_1854,N_1742,N_1716);
or U1855 (N_1855,N_1746,N_1793);
and U1856 (N_1856,N_1742,N_1749);
nor U1857 (N_1857,N_1726,N_1731);
nor U1858 (N_1858,N_1783,N_1776);
and U1859 (N_1859,N_1775,N_1746);
nor U1860 (N_1860,N_1751,N_1772);
and U1861 (N_1861,N_1707,N_1796);
nor U1862 (N_1862,N_1714,N_1790);
nor U1863 (N_1863,N_1771,N_1732);
or U1864 (N_1864,N_1716,N_1706);
xnor U1865 (N_1865,N_1717,N_1711);
nand U1866 (N_1866,N_1774,N_1796);
or U1867 (N_1867,N_1753,N_1714);
nor U1868 (N_1868,N_1773,N_1738);
nor U1869 (N_1869,N_1727,N_1711);
nor U1870 (N_1870,N_1778,N_1715);
nand U1871 (N_1871,N_1708,N_1710);
or U1872 (N_1872,N_1762,N_1792);
nor U1873 (N_1873,N_1720,N_1731);
nor U1874 (N_1874,N_1733,N_1792);
or U1875 (N_1875,N_1729,N_1771);
or U1876 (N_1876,N_1788,N_1742);
or U1877 (N_1877,N_1777,N_1767);
or U1878 (N_1878,N_1780,N_1714);
and U1879 (N_1879,N_1755,N_1763);
or U1880 (N_1880,N_1745,N_1767);
or U1881 (N_1881,N_1708,N_1795);
and U1882 (N_1882,N_1798,N_1744);
or U1883 (N_1883,N_1736,N_1756);
or U1884 (N_1884,N_1729,N_1777);
or U1885 (N_1885,N_1792,N_1753);
and U1886 (N_1886,N_1770,N_1775);
nand U1887 (N_1887,N_1744,N_1778);
and U1888 (N_1888,N_1793,N_1708);
nand U1889 (N_1889,N_1727,N_1795);
or U1890 (N_1890,N_1790,N_1783);
and U1891 (N_1891,N_1701,N_1729);
and U1892 (N_1892,N_1748,N_1734);
or U1893 (N_1893,N_1746,N_1782);
or U1894 (N_1894,N_1775,N_1717);
and U1895 (N_1895,N_1770,N_1774);
or U1896 (N_1896,N_1729,N_1761);
nand U1897 (N_1897,N_1794,N_1735);
and U1898 (N_1898,N_1779,N_1703);
nor U1899 (N_1899,N_1702,N_1746);
and U1900 (N_1900,N_1853,N_1877);
or U1901 (N_1901,N_1828,N_1813);
and U1902 (N_1902,N_1830,N_1896);
and U1903 (N_1903,N_1851,N_1850);
or U1904 (N_1904,N_1894,N_1807);
nand U1905 (N_1905,N_1800,N_1820);
nor U1906 (N_1906,N_1869,N_1875);
or U1907 (N_1907,N_1801,N_1890);
nand U1908 (N_1908,N_1834,N_1855);
nand U1909 (N_1909,N_1865,N_1848);
nand U1910 (N_1910,N_1808,N_1847);
or U1911 (N_1911,N_1872,N_1868);
or U1912 (N_1912,N_1831,N_1876);
nand U1913 (N_1913,N_1889,N_1841);
and U1914 (N_1914,N_1884,N_1859);
nand U1915 (N_1915,N_1852,N_1866);
nor U1916 (N_1916,N_1898,N_1893);
nor U1917 (N_1917,N_1871,N_1888);
or U1918 (N_1918,N_1839,N_1817);
and U1919 (N_1919,N_1837,N_1892);
and U1920 (N_1920,N_1881,N_1819);
nor U1921 (N_1921,N_1854,N_1845);
nor U1922 (N_1922,N_1815,N_1823);
nand U1923 (N_1923,N_1874,N_1829);
or U1924 (N_1924,N_1849,N_1861);
or U1925 (N_1925,N_1833,N_1887);
nor U1926 (N_1926,N_1899,N_1822);
nand U1927 (N_1927,N_1836,N_1816);
nand U1928 (N_1928,N_1840,N_1863);
or U1929 (N_1929,N_1803,N_1856);
nand U1930 (N_1930,N_1844,N_1897);
nand U1931 (N_1931,N_1826,N_1818);
nor U1932 (N_1932,N_1810,N_1882);
nand U1933 (N_1933,N_1824,N_1804);
nor U1934 (N_1934,N_1891,N_1864);
or U1935 (N_1935,N_1832,N_1862);
and U1936 (N_1936,N_1802,N_1809);
nand U1937 (N_1937,N_1835,N_1879);
nand U1938 (N_1938,N_1873,N_1885);
and U1939 (N_1939,N_1886,N_1895);
nand U1940 (N_1940,N_1811,N_1838);
nor U1941 (N_1941,N_1821,N_1880);
nor U1942 (N_1942,N_1860,N_1883);
nand U1943 (N_1943,N_1814,N_1842);
and U1944 (N_1944,N_1858,N_1806);
or U1945 (N_1945,N_1843,N_1878);
and U1946 (N_1946,N_1805,N_1867);
and U1947 (N_1947,N_1857,N_1870);
nand U1948 (N_1948,N_1846,N_1812);
nand U1949 (N_1949,N_1827,N_1825);
nor U1950 (N_1950,N_1804,N_1823);
and U1951 (N_1951,N_1818,N_1832);
and U1952 (N_1952,N_1818,N_1835);
nor U1953 (N_1953,N_1806,N_1840);
nor U1954 (N_1954,N_1806,N_1803);
and U1955 (N_1955,N_1817,N_1851);
nand U1956 (N_1956,N_1809,N_1842);
nor U1957 (N_1957,N_1879,N_1887);
and U1958 (N_1958,N_1883,N_1881);
nor U1959 (N_1959,N_1836,N_1803);
nor U1960 (N_1960,N_1842,N_1876);
or U1961 (N_1961,N_1858,N_1875);
and U1962 (N_1962,N_1887,N_1854);
nand U1963 (N_1963,N_1858,N_1882);
nand U1964 (N_1964,N_1885,N_1882);
and U1965 (N_1965,N_1819,N_1879);
nand U1966 (N_1966,N_1803,N_1895);
or U1967 (N_1967,N_1823,N_1895);
nand U1968 (N_1968,N_1889,N_1829);
or U1969 (N_1969,N_1842,N_1865);
or U1970 (N_1970,N_1864,N_1888);
xnor U1971 (N_1971,N_1854,N_1823);
nand U1972 (N_1972,N_1840,N_1844);
nand U1973 (N_1973,N_1894,N_1841);
or U1974 (N_1974,N_1842,N_1806);
and U1975 (N_1975,N_1873,N_1834);
nor U1976 (N_1976,N_1819,N_1812);
or U1977 (N_1977,N_1870,N_1896);
nand U1978 (N_1978,N_1805,N_1830);
nor U1979 (N_1979,N_1834,N_1845);
nand U1980 (N_1980,N_1854,N_1847);
or U1981 (N_1981,N_1864,N_1885);
and U1982 (N_1982,N_1815,N_1893);
nand U1983 (N_1983,N_1893,N_1842);
nand U1984 (N_1984,N_1884,N_1826);
nor U1985 (N_1985,N_1885,N_1898);
and U1986 (N_1986,N_1811,N_1835);
or U1987 (N_1987,N_1887,N_1897);
nand U1988 (N_1988,N_1807,N_1841);
nor U1989 (N_1989,N_1827,N_1888);
or U1990 (N_1990,N_1841,N_1829);
nor U1991 (N_1991,N_1895,N_1864);
nand U1992 (N_1992,N_1822,N_1814);
nand U1993 (N_1993,N_1829,N_1883);
nor U1994 (N_1994,N_1840,N_1877);
xnor U1995 (N_1995,N_1813,N_1823);
nand U1996 (N_1996,N_1863,N_1823);
nand U1997 (N_1997,N_1852,N_1833);
and U1998 (N_1998,N_1820,N_1843);
nor U1999 (N_1999,N_1898,N_1829);
nand U2000 (N_2000,N_1991,N_1957);
or U2001 (N_2001,N_1933,N_1903);
or U2002 (N_2002,N_1900,N_1941);
and U2003 (N_2003,N_1969,N_1923);
and U2004 (N_2004,N_1997,N_1986);
nand U2005 (N_2005,N_1976,N_1950);
xnor U2006 (N_2006,N_1987,N_1982);
nor U2007 (N_2007,N_1929,N_1928);
nor U2008 (N_2008,N_1983,N_1980);
nor U2009 (N_2009,N_1959,N_1994);
and U2010 (N_2010,N_1936,N_1953);
xor U2011 (N_2011,N_1901,N_1934);
nor U2012 (N_2012,N_1967,N_1975);
and U2013 (N_2013,N_1974,N_1960);
and U2014 (N_2014,N_1968,N_1920);
nand U2015 (N_2015,N_1902,N_1979);
or U2016 (N_2016,N_1984,N_1944);
nor U2017 (N_2017,N_1954,N_1907);
nor U2018 (N_2018,N_1942,N_1981);
or U2019 (N_2019,N_1955,N_1932);
or U2020 (N_2020,N_1949,N_1905);
or U2021 (N_2021,N_1916,N_1925);
and U2022 (N_2022,N_1921,N_1912);
and U2023 (N_2023,N_1952,N_1963);
or U2024 (N_2024,N_1922,N_1938);
nand U2025 (N_2025,N_1966,N_1904);
nor U2026 (N_2026,N_1972,N_1985);
nand U2027 (N_2027,N_1927,N_1909);
or U2028 (N_2028,N_1992,N_1937);
and U2029 (N_2029,N_1948,N_1951);
nor U2030 (N_2030,N_1993,N_1917);
and U2031 (N_2031,N_1945,N_1971);
nor U2032 (N_2032,N_1964,N_1930);
and U2033 (N_2033,N_1965,N_1918);
and U2034 (N_2034,N_1939,N_1970);
nor U2035 (N_2035,N_1935,N_1946);
and U2036 (N_2036,N_1908,N_1956);
and U2037 (N_2037,N_1911,N_1915);
and U2038 (N_2038,N_1988,N_1940);
and U2039 (N_2039,N_1926,N_1999);
or U2040 (N_2040,N_1962,N_1998);
nand U2041 (N_2041,N_1931,N_1973);
and U2042 (N_2042,N_1914,N_1924);
or U2043 (N_2043,N_1990,N_1906);
xor U2044 (N_2044,N_1995,N_1910);
and U2045 (N_2045,N_1958,N_1978);
nand U2046 (N_2046,N_1989,N_1996);
and U2047 (N_2047,N_1947,N_1977);
or U2048 (N_2048,N_1961,N_1913);
nand U2049 (N_2049,N_1943,N_1919);
nand U2050 (N_2050,N_1965,N_1933);
nor U2051 (N_2051,N_1939,N_1943);
nand U2052 (N_2052,N_1945,N_1988);
nand U2053 (N_2053,N_1948,N_1979);
or U2054 (N_2054,N_1902,N_1968);
or U2055 (N_2055,N_1900,N_1974);
nor U2056 (N_2056,N_1948,N_1940);
or U2057 (N_2057,N_1968,N_1977);
or U2058 (N_2058,N_1965,N_1911);
or U2059 (N_2059,N_1913,N_1909);
or U2060 (N_2060,N_1984,N_1995);
or U2061 (N_2061,N_1913,N_1956);
and U2062 (N_2062,N_1957,N_1978);
nand U2063 (N_2063,N_1962,N_1947);
nand U2064 (N_2064,N_1909,N_1955);
or U2065 (N_2065,N_1927,N_1991);
nor U2066 (N_2066,N_1908,N_1918);
or U2067 (N_2067,N_1962,N_1983);
or U2068 (N_2068,N_1937,N_1940);
nor U2069 (N_2069,N_1948,N_1967);
nand U2070 (N_2070,N_1925,N_1997);
nor U2071 (N_2071,N_1916,N_1946);
nor U2072 (N_2072,N_1916,N_1900);
and U2073 (N_2073,N_1950,N_1957);
or U2074 (N_2074,N_1934,N_1912);
nand U2075 (N_2075,N_1975,N_1933);
and U2076 (N_2076,N_1996,N_1981);
nand U2077 (N_2077,N_1915,N_1922);
and U2078 (N_2078,N_1944,N_1999);
nand U2079 (N_2079,N_1932,N_1963);
and U2080 (N_2080,N_1945,N_1990);
nor U2081 (N_2081,N_1971,N_1927);
or U2082 (N_2082,N_1910,N_1916);
and U2083 (N_2083,N_1970,N_1952);
nor U2084 (N_2084,N_1951,N_1991);
and U2085 (N_2085,N_1942,N_1904);
and U2086 (N_2086,N_1949,N_1962);
nor U2087 (N_2087,N_1993,N_1905);
or U2088 (N_2088,N_1921,N_1949);
and U2089 (N_2089,N_1933,N_1989);
nand U2090 (N_2090,N_1901,N_1969);
nor U2091 (N_2091,N_1935,N_1920);
nand U2092 (N_2092,N_1932,N_1931);
and U2093 (N_2093,N_1956,N_1985);
nor U2094 (N_2094,N_1904,N_1941);
nor U2095 (N_2095,N_1989,N_1916);
and U2096 (N_2096,N_1942,N_1911);
or U2097 (N_2097,N_1963,N_1990);
xnor U2098 (N_2098,N_1997,N_1903);
and U2099 (N_2099,N_1993,N_1944);
or U2100 (N_2100,N_2003,N_2061);
nor U2101 (N_2101,N_2063,N_2051);
nand U2102 (N_2102,N_2094,N_2073);
and U2103 (N_2103,N_2014,N_2052);
or U2104 (N_2104,N_2067,N_2041);
or U2105 (N_2105,N_2008,N_2070);
nand U2106 (N_2106,N_2028,N_2066);
or U2107 (N_2107,N_2012,N_2060);
or U2108 (N_2108,N_2077,N_2057);
or U2109 (N_2109,N_2015,N_2097);
or U2110 (N_2110,N_2075,N_2044);
nor U2111 (N_2111,N_2042,N_2024);
and U2112 (N_2112,N_2085,N_2099);
and U2113 (N_2113,N_2022,N_2021);
and U2114 (N_2114,N_2025,N_2084);
or U2115 (N_2115,N_2026,N_2053);
nor U2116 (N_2116,N_2038,N_2092);
nor U2117 (N_2117,N_2032,N_2091);
nor U2118 (N_2118,N_2019,N_2034);
and U2119 (N_2119,N_2027,N_2082);
or U2120 (N_2120,N_2029,N_2031);
nand U2121 (N_2121,N_2083,N_2006);
nand U2122 (N_2122,N_2056,N_2072);
or U2123 (N_2123,N_2096,N_2002);
xor U2124 (N_2124,N_2048,N_2071);
or U2125 (N_2125,N_2047,N_2069);
nand U2126 (N_2126,N_2074,N_2087);
nor U2127 (N_2127,N_2030,N_2009);
or U2128 (N_2128,N_2000,N_2076);
and U2129 (N_2129,N_2078,N_2046);
nor U2130 (N_2130,N_2058,N_2004);
and U2131 (N_2131,N_2055,N_2086);
and U2132 (N_2132,N_2098,N_2039);
or U2133 (N_2133,N_2081,N_2059);
and U2134 (N_2134,N_2043,N_2033);
nor U2135 (N_2135,N_2020,N_2093);
or U2136 (N_2136,N_2010,N_2016);
nor U2137 (N_2137,N_2064,N_2089);
and U2138 (N_2138,N_2036,N_2045);
and U2139 (N_2139,N_2023,N_2011);
or U2140 (N_2140,N_2017,N_2088);
nand U2141 (N_2141,N_2054,N_2062);
or U2142 (N_2142,N_2037,N_2079);
nor U2143 (N_2143,N_2018,N_2040);
or U2144 (N_2144,N_2001,N_2035);
and U2145 (N_2145,N_2090,N_2080);
nor U2146 (N_2146,N_2065,N_2005);
nor U2147 (N_2147,N_2007,N_2049);
and U2148 (N_2148,N_2095,N_2068);
and U2149 (N_2149,N_2050,N_2013);
nor U2150 (N_2150,N_2064,N_2069);
nor U2151 (N_2151,N_2017,N_2015);
nand U2152 (N_2152,N_2004,N_2010);
and U2153 (N_2153,N_2091,N_2038);
nor U2154 (N_2154,N_2001,N_2007);
nand U2155 (N_2155,N_2089,N_2054);
nor U2156 (N_2156,N_2067,N_2039);
or U2157 (N_2157,N_2071,N_2054);
nand U2158 (N_2158,N_2077,N_2045);
nor U2159 (N_2159,N_2094,N_2007);
or U2160 (N_2160,N_2088,N_2030);
and U2161 (N_2161,N_2016,N_2000);
nor U2162 (N_2162,N_2051,N_2035);
or U2163 (N_2163,N_2053,N_2035);
or U2164 (N_2164,N_2083,N_2041);
nor U2165 (N_2165,N_2054,N_2038);
nand U2166 (N_2166,N_2045,N_2035);
and U2167 (N_2167,N_2067,N_2049);
nand U2168 (N_2168,N_2010,N_2005);
or U2169 (N_2169,N_2055,N_2004);
nor U2170 (N_2170,N_2049,N_2053);
nor U2171 (N_2171,N_2030,N_2029);
and U2172 (N_2172,N_2070,N_2007);
and U2173 (N_2173,N_2039,N_2033);
or U2174 (N_2174,N_2040,N_2082);
or U2175 (N_2175,N_2036,N_2072);
and U2176 (N_2176,N_2000,N_2023);
or U2177 (N_2177,N_2070,N_2035);
or U2178 (N_2178,N_2069,N_2001);
nand U2179 (N_2179,N_2047,N_2086);
and U2180 (N_2180,N_2082,N_2070);
and U2181 (N_2181,N_2093,N_2075);
nand U2182 (N_2182,N_2070,N_2024);
or U2183 (N_2183,N_2080,N_2060);
nor U2184 (N_2184,N_2046,N_2039);
or U2185 (N_2185,N_2098,N_2073);
nand U2186 (N_2186,N_2041,N_2032);
xor U2187 (N_2187,N_2090,N_2051);
xnor U2188 (N_2188,N_2066,N_2082);
nand U2189 (N_2189,N_2018,N_2033);
or U2190 (N_2190,N_2082,N_2093);
nand U2191 (N_2191,N_2081,N_2010);
nor U2192 (N_2192,N_2075,N_2028);
nor U2193 (N_2193,N_2028,N_2049);
nor U2194 (N_2194,N_2017,N_2001);
and U2195 (N_2195,N_2059,N_2091);
nand U2196 (N_2196,N_2055,N_2048);
and U2197 (N_2197,N_2058,N_2013);
nand U2198 (N_2198,N_2076,N_2002);
nor U2199 (N_2199,N_2095,N_2013);
or U2200 (N_2200,N_2175,N_2168);
nor U2201 (N_2201,N_2167,N_2149);
xnor U2202 (N_2202,N_2112,N_2189);
xnor U2203 (N_2203,N_2177,N_2156);
and U2204 (N_2204,N_2181,N_2114);
or U2205 (N_2205,N_2188,N_2134);
nor U2206 (N_2206,N_2120,N_2117);
or U2207 (N_2207,N_2146,N_2148);
or U2208 (N_2208,N_2138,N_2109);
and U2209 (N_2209,N_2105,N_2152);
nor U2210 (N_2210,N_2108,N_2164);
nand U2211 (N_2211,N_2158,N_2136);
and U2212 (N_2212,N_2187,N_2123);
or U2213 (N_2213,N_2192,N_2185);
or U2214 (N_2214,N_2125,N_2115);
and U2215 (N_2215,N_2100,N_2174);
and U2216 (N_2216,N_2197,N_2124);
nand U2217 (N_2217,N_2127,N_2166);
xor U2218 (N_2218,N_2129,N_2137);
or U2219 (N_2219,N_2104,N_2107);
or U2220 (N_2220,N_2122,N_2119);
nor U2221 (N_2221,N_2155,N_2102);
nand U2222 (N_2222,N_2179,N_2111);
nand U2223 (N_2223,N_2199,N_2147);
nand U2224 (N_2224,N_2196,N_2191);
or U2225 (N_2225,N_2132,N_2171);
xor U2226 (N_2226,N_2140,N_2110);
xnor U2227 (N_2227,N_2153,N_2178);
or U2228 (N_2228,N_2128,N_2194);
nand U2229 (N_2229,N_2101,N_2113);
or U2230 (N_2230,N_2195,N_2103);
or U2231 (N_2231,N_2106,N_2165);
xor U2232 (N_2232,N_2154,N_2130);
nor U2233 (N_2233,N_2198,N_2170);
nand U2234 (N_2234,N_2159,N_2116);
or U2235 (N_2235,N_2184,N_2169);
and U2236 (N_2236,N_2172,N_2163);
and U2237 (N_2237,N_2118,N_2142);
nor U2238 (N_2238,N_2150,N_2183);
and U2239 (N_2239,N_2135,N_2176);
and U2240 (N_2240,N_2133,N_2126);
nor U2241 (N_2241,N_2145,N_2144);
or U2242 (N_2242,N_2151,N_2141);
and U2243 (N_2243,N_2131,N_2143);
or U2244 (N_2244,N_2180,N_2190);
xor U2245 (N_2245,N_2157,N_2193);
or U2246 (N_2246,N_2173,N_2139);
or U2247 (N_2247,N_2160,N_2162);
and U2248 (N_2248,N_2186,N_2182);
nand U2249 (N_2249,N_2121,N_2161);
nand U2250 (N_2250,N_2173,N_2154);
nor U2251 (N_2251,N_2126,N_2177);
and U2252 (N_2252,N_2117,N_2102);
nand U2253 (N_2253,N_2133,N_2185);
nand U2254 (N_2254,N_2121,N_2113);
and U2255 (N_2255,N_2188,N_2111);
and U2256 (N_2256,N_2125,N_2144);
nor U2257 (N_2257,N_2179,N_2129);
nor U2258 (N_2258,N_2191,N_2171);
and U2259 (N_2259,N_2126,N_2123);
nand U2260 (N_2260,N_2105,N_2149);
or U2261 (N_2261,N_2181,N_2128);
nor U2262 (N_2262,N_2105,N_2102);
nor U2263 (N_2263,N_2185,N_2174);
nor U2264 (N_2264,N_2102,N_2157);
or U2265 (N_2265,N_2108,N_2180);
or U2266 (N_2266,N_2138,N_2192);
nand U2267 (N_2267,N_2127,N_2117);
and U2268 (N_2268,N_2147,N_2130);
and U2269 (N_2269,N_2144,N_2111);
or U2270 (N_2270,N_2155,N_2194);
and U2271 (N_2271,N_2183,N_2125);
nor U2272 (N_2272,N_2110,N_2158);
nor U2273 (N_2273,N_2170,N_2157);
and U2274 (N_2274,N_2186,N_2168);
and U2275 (N_2275,N_2179,N_2130);
and U2276 (N_2276,N_2162,N_2153);
nor U2277 (N_2277,N_2177,N_2123);
or U2278 (N_2278,N_2186,N_2124);
nor U2279 (N_2279,N_2196,N_2182);
xor U2280 (N_2280,N_2192,N_2195);
nor U2281 (N_2281,N_2132,N_2155);
and U2282 (N_2282,N_2112,N_2197);
and U2283 (N_2283,N_2133,N_2106);
xnor U2284 (N_2284,N_2138,N_2126);
nand U2285 (N_2285,N_2129,N_2128);
nand U2286 (N_2286,N_2181,N_2189);
nor U2287 (N_2287,N_2163,N_2162);
nand U2288 (N_2288,N_2135,N_2170);
or U2289 (N_2289,N_2147,N_2139);
nor U2290 (N_2290,N_2109,N_2142);
nand U2291 (N_2291,N_2100,N_2146);
and U2292 (N_2292,N_2156,N_2198);
nand U2293 (N_2293,N_2139,N_2186);
nor U2294 (N_2294,N_2144,N_2159);
and U2295 (N_2295,N_2163,N_2193);
and U2296 (N_2296,N_2122,N_2191);
nand U2297 (N_2297,N_2141,N_2117);
or U2298 (N_2298,N_2128,N_2146);
and U2299 (N_2299,N_2102,N_2176);
and U2300 (N_2300,N_2299,N_2259);
nor U2301 (N_2301,N_2291,N_2264);
nor U2302 (N_2302,N_2245,N_2288);
and U2303 (N_2303,N_2208,N_2252);
nor U2304 (N_2304,N_2257,N_2236);
or U2305 (N_2305,N_2235,N_2258);
nand U2306 (N_2306,N_2224,N_2206);
nor U2307 (N_2307,N_2241,N_2289);
nor U2308 (N_2308,N_2227,N_2268);
nand U2309 (N_2309,N_2207,N_2263);
nor U2310 (N_2310,N_2298,N_2271);
or U2311 (N_2311,N_2203,N_2261);
nand U2312 (N_2312,N_2210,N_2242);
or U2313 (N_2313,N_2221,N_2286);
nor U2314 (N_2314,N_2211,N_2234);
nand U2315 (N_2315,N_2250,N_2269);
nor U2316 (N_2316,N_2213,N_2248);
or U2317 (N_2317,N_2243,N_2214);
nand U2318 (N_2318,N_2246,N_2287);
nor U2319 (N_2319,N_2231,N_2270);
nand U2320 (N_2320,N_2228,N_2247);
nor U2321 (N_2321,N_2223,N_2201);
nand U2322 (N_2322,N_2220,N_2239);
and U2323 (N_2323,N_2283,N_2249);
nand U2324 (N_2324,N_2273,N_2297);
nand U2325 (N_2325,N_2215,N_2255);
nor U2326 (N_2326,N_2205,N_2222);
and U2327 (N_2327,N_2233,N_2294);
or U2328 (N_2328,N_2262,N_2279);
nor U2329 (N_2329,N_2238,N_2232);
nor U2330 (N_2330,N_2284,N_2229);
nand U2331 (N_2331,N_2251,N_2265);
and U2332 (N_2332,N_2290,N_2277);
or U2333 (N_2333,N_2292,N_2230);
and U2334 (N_2334,N_2240,N_2296);
nand U2335 (N_2335,N_2209,N_2253);
nor U2336 (N_2336,N_2272,N_2216);
nor U2337 (N_2337,N_2225,N_2212);
and U2338 (N_2338,N_2280,N_2278);
nand U2339 (N_2339,N_2200,N_2295);
nand U2340 (N_2340,N_2266,N_2218);
or U2341 (N_2341,N_2202,N_2267);
or U2342 (N_2342,N_2219,N_2276);
xnor U2343 (N_2343,N_2226,N_2260);
nor U2344 (N_2344,N_2254,N_2217);
or U2345 (N_2345,N_2237,N_2285);
or U2346 (N_2346,N_2256,N_2274);
nor U2347 (N_2347,N_2275,N_2244);
nand U2348 (N_2348,N_2281,N_2204);
nand U2349 (N_2349,N_2293,N_2282);
nand U2350 (N_2350,N_2248,N_2293);
nor U2351 (N_2351,N_2227,N_2231);
nand U2352 (N_2352,N_2264,N_2283);
or U2353 (N_2353,N_2211,N_2287);
and U2354 (N_2354,N_2299,N_2260);
or U2355 (N_2355,N_2223,N_2248);
or U2356 (N_2356,N_2291,N_2289);
or U2357 (N_2357,N_2247,N_2232);
or U2358 (N_2358,N_2251,N_2283);
nand U2359 (N_2359,N_2280,N_2202);
or U2360 (N_2360,N_2264,N_2215);
nor U2361 (N_2361,N_2208,N_2287);
nor U2362 (N_2362,N_2264,N_2234);
or U2363 (N_2363,N_2222,N_2245);
and U2364 (N_2364,N_2214,N_2225);
or U2365 (N_2365,N_2258,N_2208);
and U2366 (N_2366,N_2260,N_2231);
and U2367 (N_2367,N_2223,N_2242);
nand U2368 (N_2368,N_2224,N_2207);
nor U2369 (N_2369,N_2288,N_2215);
nor U2370 (N_2370,N_2282,N_2226);
nor U2371 (N_2371,N_2291,N_2200);
or U2372 (N_2372,N_2274,N_2269);
nand U2373 (N_2373,N_2299,N_2200);
nand U2374 (N_2374,N_2238,N_2262);
and U2375 (N_2375,N_2232,N_2258);
nor U2376 (N_2376,N_2208,N_2253);
nor U2377 (N_2377,N_2298,N_2265);
and U2378 (N_2378,N_2217,N_2226);
nor U2379 (N_2379,N_2266,N_2224);
xnor U2380 (N_2380,N_2243,N_2209);
nand U2381 (N_2381,N_2206,N_2242);
nor U2382 (N_2382,N_2241,N_2266);
nor U2383 (N_2383,N_2237,N_2216);
xor U2384 (N_2384,N_2220,N_2284);
or U2385 (N_2385,N_2225,N_2224);
or U2386 (N_2386,N_2219,N_2213);
nor U2387 (N_2387,N_2209,N_2272);
nor U2388 (N_2388,N_2237,N_2284);
nand U2389 (N_2389,N_2291,N_2287);
nand U2390 (N_2390,N_2222,N_2282);
and U2391 (N_2391,N_2246,N_2251);
nor U2392 (N_2392,N_2280,N_2235);
nor U2393 (N_2393,N_2230,N_2205);
nand U2394 (N_2394,N_2284,N_2228);
and U2395 (N_2395,N_2261,N_2230);
and U2396 (N_2396,N_2200,N_2265);
or U2397 (N_2397,N_2211,N_2296);
and U2398 (N_2398,N_2208,N_2204);
or U2399 (N_2399,N_2202,N_2283);
nand U2400 (N_2400,N_2308,N_2392);
and U2401 (N_2401,N_2393,N_2324);
and U2402 (N_2402,N_2378,N_2330);
or U2403 (N_2403,N_2345,N_2390);
nand U2404 (N_2404,N_2369,N_2368);
nor U2405 (N_2405,N_2374,N_2375);
and U2406 (N_2406,N_2348,N_2363);
nor U2407 (N_2407,N_2349,N_2354);
nand U2408 (N_2408,N_2323,N_2342);
or U2409 (N_2409,N_2351,N_2394);
or U2410 (N_2410,N_2322,N_2358);
and U2411 (N_2411,N_2361,N_2373);
or U2412 (N_2412,N_2327,N_2352);
nand U2413 (N_2413,N_2371,N_2300);
or U2414 (N_2414,N_2320,N_2376);
nor U2415 (N_2415,N_2332,N_2353);
nand U2416 (N_2416,N_2344,N_2396);
nor U2417 (N_2417,N_2313,N_2318);
nand U2418 (N_2418,N_2382,N_2389);
and U2419 (N_2419,N_2339,N_2381);
or U2420 (N_2420,N_2334,N_2359);
nor U2421 (N_2421,N_2367,N_2379);
nor U2422 (N_2422,N_2364,N_2329);
and U2423 (N_2423,N_2302,N_2316);
or U2424 (N_2424,N_2325,N_2386);
and U2425 (N_2425,N_2317,N_2346);
and U2426 (N_2426,N_2328,N_2365);
nand U2427 (N_2427,N_2338,N_2380);
nand U2428 (N_2428,N_2357,N_2388);
and U2429 (N_2429,N_2350,N_2310);
nand U2430 (N_2430,N_2312,N_2304);
nand U2431 (N_2431,N_2397,N_2336);
nor U2432 (N_2432,N_2319,N_2311);
or U2433 (N_2433,N_2387,N_2340);
or U2434 (N_2434,N_2372,N_2301);
and U2435 (N_2435,N_2399,N_2362);
nor U2436 (N_2436,N_2333,N_2315);
nor U2437 (N_2437,N_2314,N_2343);
or U2438 (N_2438,N_2398,N_2335);
or U2439 (N_2439,N_2307,N_2395);
nand U2440 (N_2440,N_2326,N_2356);
nor U2441 (N_2441,N_2384,N_2385);
or U2442 (N_2442,N_2337,N_2391);
nand U2443 (N_2443,N_2331,N_2355);
and U2444 (N_2444,N_2347,N_2303);
nor U2445 (N_2445,N_2305,N_2321);
or U2446 (N_2446,N_2341,N_2306);
or U2447 (N_2447,N_2370,N_2309);
nand U2448 (N_2448,N_2383,N_2377);
nand U2449 (N_2449,N_2360,N_2366);
and U2450 (N_2450,N_2336,N_2368);
or U2451 (N_2451,N_2352,N_2326);
and U2452 (N_2452,N_2390,N_2365);
nand U2453 (N_2453,N_2399,N_2355);
and U2454 (N_2454,N_2358,N_2308);
and U2455 (N_2455,N_2321,N_2383);
and U2456 (N_2456,N_2304,N_2347);
nand U2457 (N_2457,N_2372,N_2318);
or U2458 (N_2458,N_2367,N_2322);
or U2459 (N_2459,N_2366,N_2314);
or U2460 (N_2460,N_2342,N_2356);
xor U2461 (N_2461,N_2389,N_2342);
and U2462 (N_2462,N_2372,N_2393);
nand U2463 (N_2463,N_2373,N_2362);
and U2464 (N_2464,N_2330,N_2364);
nand U2465 (N_2465,N_2385,N_2315);
nor U2466 (N_2466,N_2366,N_2373);
nand U2467 (N_2467,N_2396,N_2381);
nand U2468 (N_2468,N_2379,N_2323);
or U2469 (N_2469,N_2303,N_2388);
nand U2470 (N_2470,N_2349,N_2346);
and U2471 (N_2471,N_2348,N_2317);
and U2472 (N_2472,N_2303,N_2376);
nand U2473 (N_2473,N_2385,N_2326);
nand U2474 (N_2474,N_2345,N_2326);
or U2475 (N_2475,N_2385,N_2310);
nor U2476 (N_2476,N_2368,N_2302);
xnor U2477 (N_2477,N_2328,N_2313);
and U2478 (N_2478,N_2348,N_2393);
nand U2479 (N_2479,N_2373,N_2305);
and U2480 (N_2480,N_2306,N_2344);
and U2481 (N_2481,N_2309,N_2375);
nor U2482 (N_2482,N_2355,N_2384);
xor U2483 (N_2483,N_2356,N_2338);
or U2484 (N_2484,N_2364,N_2309);
and U2485 (N_2485,N_2398,N_2385);
nor U2486 (N_2486,N_2322,N_2384);
or U2487 (N_2487,N_2336,N_2370);
nor U2488 (N_2488,N_2364,N_2356);
nand U2489 (N_2489,N_2388,N_2336);
or U2490 (N_2490,N_2364,N_2352);
nand U2491 (N_2491,N_2368,N_2399);
and U2492 (N_2492,N_2399,N_2383);
and U2493 (N_2493,N_2302,N_2389);
and U2494 (N_2494,N_2393,N_2303);
or U2495 (N_2495,N_2341,N_2369);
or U2496 (N_2496,N_2303,N_2381);
xor U2497 (N_2497,N_2341,N_2315);
and U2498 (N_2498,N_2377,N_2311);
nor U2499 (N_2499,N_2353,N_2360);
nor U2500 (N_2500,N_2426,N_2464);
nand U2501 (N_2501,N_2420,N_2421);
and U2502 (N_2502,N_2484,N_2454);
nand U2503 (N_2503,N_2407,N_2406);
and U2504 (N_2504,N_2437,N_2492);
or U2505 (N_2505,N_2497,N_2483);
nand U2506 (N_2506,N_2455,N_2453);
nor U2507 (N_2507,N_2451,N_2476);
nand U2508 (N_2508,N_2431,N_2466);
or U2509 (N_2509,N_2432,N_2411);
and U2510 (N_2510,N_2465,N_2408);
nand U2511 (N_2511,N_2400,N_2417);
nand U2512 (N_2512,N_2467,N_2418);
nand U2513 (N_2513,N_2419,N_2425);
nand U2514 (N_2514,N_2414,N_2443);
and U2515 (N_2515,N_2422,N_2413);
or U2516 (N_2516,N_2468,N_2459);
nor U2517 (N_2517,N_2428,N_2410);
and U2518 (N_2518,N_2489,N_2445);
or U2519 (N_2519,N_2439,N_2446);
xor U2520 (N_2520,N_2499,N_2441);
nor U2521 (N_2521,N_2491,N_2494);
or U2522 (N_2522,N_2478,N_2474);
nand U2523 (N_2523,N_2462,N_2442);
nand U2524 (N_2524,N_2481,N_2433);
and U2525 (N_2525,N_2436,N_2452);
or U2526 (N_2526,N_2461,N_2429);
xor U2527 (N_2527,N_2470,N_2424);
nor U2528 (N_2528,N_2435,N_2458);
or U2529 (N_2529,N_2477,N_2480);
and U2530 (N_2530,N_2471,N_2479);
nor U2531 (N_2531,N_2415,N_2427);
and U2532 (N_2532,N_2472,N_2493);
nand U2533 (N_2533,N_2486,N_2487);
nor U2534 (N_2534,N_2498,N_2438);
or U2535 (N_2535,N_2403,N_2405);
nor U2536 (N_2536,N_2495,N_2473);
nand U2537 (N_2537,N_2401,N_2412);
or U2538 (N_2538,N_2444,N_2450);
nand U2539 (N_2539,N_2457,N_2490);
and U2540 (N_2540,N_2404,N_2496);
nor U2541 (N_2541,N_2463,N_2447);
nor U2542 (N_2542,N_2416,N_2460);
or U2543 (N_2543,N_2469,N_2434);
nor U2544 (N_2544,N_2440,N_2485);
nor U2545 (N_2545,N_2423,N_2488);
xor U2546 (N_2546,N_2449,N_2448);
and U2547 (N_2547,N_2430,N_2409);
nor U2548 (N_2548,N_2456,N_2402);
and U2549 (N_2549,N_2475,N_2482);
and U2550 (N_2550,N_2412,N_2407);
nor U2551 (N_2551,N_2492,N_2414);
nor U2552 (N_2552,N_2481,N_2450);
and U2553 (N_2553,N_2462,N_2455);
xnor U2554 (N_2554,N_2425,N_2418);
and U2555 (N_2555,N_2483,N_2447);
and U2556 (N_2556,N_2425,N_2435);
or U2557 (N_2557,N_2455,N_2412);
nor U2558 (N_2558,N_2451,N_2427);
nor U2559 (N_2559,N_2435,N_2479);
nor U2560 (N_2560,N_2418,N_2440);
nor U2561 (N_2561,N_2453,N_2423);
nand U2562 (N_2562,N_2498,N_2428);
nand U2563 (N_2563,N_2486,N_2467);
nor U2564 (N_2564,N_2485,N_2446);
and U2565 (N_2565,N_2488,N_2438);
and U2566 (N_2566,N_2419,N_2463);
or U2567 (N_2567,N_2477,N_2466);
and U2568 (N_2568,N_2451,N_2406);
xnor U2569 (N_2569,N_2419,N_2445);
nor U2570 (N_2570,N_2497,N_2467);
and U2571 (N_2571,N_2425,N_2426);
nor U2572 (N_2572,N_2406,N_2462);
or U2573 (N_2573,N_2495,N_2454);
nand U2574 (N_2574,N_2455,N_2475);
xnor U2575 (N_2575,N_2499,N_2465);
and U2576 (N_2576,N_2468,N_2408);
and U2577 (N_2577,N_2467,N_2453);
nor U2578 (N_2578,N_2495,N_2430);
nand U2579 (N_2579,N_2446,N_2445);
nor U2580 (N_2580,N_2444,N_2489);
or U2581 (N_2581,N_2465,N_2425);
and U2582 (N_2582,N_2425,N_2448);
nor U2583 (N_2583,N_2419,N_2471);
xnor U2584 (N_2584,N_2430,N_2406);
or U2585 (N_2585,N_2406,N_2426);
or U2586 (N_2586,N_2414,N_2435);
or U2587 (N_2587,N_2423,N_2460);
or U2588 (N_2588,N_2460,N_2494);
or U2589 (N_2589,N_2491,N_2485);
nor U2590 (N_2590,N_2483,N_2461);
nor U2591 (N_2591,N_2410,N_2448);
and U2592 (N_2592,N_2418,N_2407);
and U2593 (N_2593,N_2453,N_2469);
or U2594 (N_2594,N_2423,N_2462);
or U2595 (N_2595,N_2424,N_2440);
or U2596 (N_2596,N_2440,N_2464);
and U2597 (N_2597,N_2479,N_2424);
or U2598 (N_2598,N_2440,N_2462);
xor U2599 (N_2599,N_2403,N_2431);
nand U2600 (N_2600,N_2536,N_2509);
or U2601 (N_2601,N_2529,N_2581);
and U2602 (N_2602,N_2544,N_2550);
nand U2603 (N_2603,N_2592,N_2586);
nand U2604 (N_2604,N_2541,N_2539);
nor U2605 (N_2605,N_2516,N_2583);
or U2606 (N_2606,N_2500,N_2538);
and U2607 (N_2607,N_2571,N_2563);
nor U2608 (N_2608,N_2528,N_2547);
nor U2609 (N_2609,N_2519,N_2594);
and U2610 (N_2610,N_2590,N_2534);
nand U2611 (N_2611,N_2598,N_2582);
or U2612 (N_2612,N_2537,N_2572);
and U2613 (N_2613,N_2515,N_2559);
nand U2614 (N_2614,N_2520,N_2525);
or U2615 (N_2615,N_2545,N_2578);
nor U2616 (N_2616,N_2530,N_2543);
nand U2617 (N_2617,N_2579,N_2521);
nor U2618 (N_2618,N_2595,N_2570);
and U2619 (N_2619,N_2565,N_2564);
or U2620 (N_2620,N_2555,N_2507);
nor U2621 (N_2621,N_2517,N_2527);
nor U2622 (N_2622,N_2511,N_2526);
and U2623 (N_2623,N_2558,N_2566);
nand U2624 (N_2624,N_2504,N_2593);
nor U2625 (N_2625,N_2502,N_2501);
nand U2626 (N_2626,N_2584,N_2512);
or U2627 (N_2627,N_2532,N_2573);
nor U2628 (N_2628,N_2549,N_2587);
or U2629 (N_2629,N_2518,N_2540);
xor U2630 (N_2630,N_2580,N_2588);
nor U2631 (N_2631,N_2567,N_2569);
or U2632 (N_2632,N_2505,N_2506);
or U2633 (N_2633,N_2554,N_2599);
nor U2634 (N_2634,N_2503,N_2531);
nand U2635 (N_2635,N_2589,N_2542);
and U2636 (N_2636,N_2552,N_2556);
or U2637 (N_2637,N_2577,N_2596);
nor U2638 (N_2638,N_2524,N_2561);
nor U2639 (N_2639,N_2546,N_2562);
nand U2640 (N_2640,N_2575,N_2510);
and U2641 (N_2641,N_2560,N_2523);
nand U2642 (N_2642,N_2557,N_2514);
nor U2643 (N_2643,N_2513,N_2574);
or U2644 (N_2644,N_2535,N_2508);
nand U2645 (N_2645,N_2585,N_2548);
nand U2646 (N_2646,N_2568,N_2553);
or U2647 (N_2647,N_2533,N_2576);
nor U2648 (N_2648,N_2591,N_2522);
and U2649 (N_2649,N_2597,N_2551);
and U2650 (N_2650,N_2587,N_2561);
nand U2651 (N_2651,N_2554,N_2597);
nor U2652 (N_2652,N_2516,N_2584);
nor U2653 (N_2653,N_2579,N_2503);
and U2654 (N_2654,N_2552,N_2550);
nand U2655 (N_2655,N_2522,N_2503);
nand U2656 (N_2656,N_2552,N_2517);
nand U2657 (N_2657,N_2526,N_2510);
or U2658 (N_2658,N_2582,N_2596);
nor U2659 (N_2659,N_2512,N_2524);
nand U2660 (N_2660,N_2574,N_2565);
nand U2661 (N_2661,N_2591,N_2567);
nor U2662 (N_2662,N_2510,N_2532);
nand U2663 (N_2663,N_2537,N_2527);
nand U2664 (N_2664,N_2553,N_2587);
and U2665 (N_2665,N_2591,N_2597);
and U2666 (N_2666,N_2506,N_2526);
and U2667 (N_2667,N_2560,N_2582);
nand U2668 (N_2668,N_2557,N_2524);
nor U2669 (N_2669,N_2506,N_2595);
or U2670 (N_2670,N_2514,N_2561);
nand U2671 (N_2671,N_2544,N_2540);
and U2672 (N_2672,N_2508,N_2531);
nand U2673 (N_2673,N_2501,N_2557);
and U2674 (N_2674,N_2519,N_2544);
and U2675 (N_2675,N_2536,N_2566);
nand U2676 (N_2676,N_2563,N_2589);
nand U2677 (N_2677,N_2587,N_2539);
nand U2678 (N_2678,N_2598,N_2545);
or U2679 (N_2679,N_2548,N_2543);
nand U2680 (N_2680,N_2551,N_2584);
nor U2681 (N_2681,N_2564,N_2576);
and U2682 (N_2682,N_2583,N_2547);
or U2683 (N_2683,N_2598,N_2501);
nor U2684 (N_2684,N_2552,N_2544);
nor U2685 (N_2685,N_2579,N_2519);
nand U2686 (N_2686,N_2508,N_2597);
nor U2687 (N_2687,N_2579,N_2566);
nand U2688 (N_2688,N_2572,N_2587);
and U2689 (N_2689,N_2572,N_2575);
and U2690 (N_2690,N_2590,N_2512);
nor U2691 (N_2691,N_2537,N_2505);
or U2692 (N_2692,N_2529,N_2582);
nor U2693 (N_2693,N_2538,N_2575);
nor U2694 (N_2694,N_2558,N_2579);
and U2695 (N_2695,N_2583,N_2540);
nor U2696 (N_2696,N_2515,N_2547);
or U2697 (N_2697,N_2561,N_2592);
and U2698 (N_2698,N_2552,N_2523);
xnor U2699 (N_2699,N_2519,N_2528);
nand U2700 (N_2700,N_2610,N_2669);
and U2701 (N_2701,N_2633,N_2611);
nor U2702 (N_2702,N_2635,N_2668);
nand U2703 (N_2703,N_2674,N_2698);
and U2704 (N_2704,N_2629,N_2678);
nor U2705 (N_2705,N_2623,N_2636);
or U2706 (N_2706,N_2689,N_2614);
or U2707 (N_2707,N_2631,N_2683);
and U2708 (N_2708,N_2618,N_2682);
nand U2709 (N_2709,N_2673,N_2622);
or U2710 (N_2710,N_2679,N_2606);
nor U2711 (N_2711,N_2665,N_2612);
or U2712 (N_2712,N_2620,N_2648);
nand U2713 (N_2713,N_2677,N_2600);
nor U2714 (N_2714,N_2670,N_2651);
and U2715 (N_2715,N_2630,N_2696);
nor U2716 (N_2716,N_2645,N_2661);
nor U2717 (N_2717,N_2642,N_2615);
nor U2718 (N_2718,N_2602,N_2667);
nor U2719 (N_2719,N_2663,N_2657);
nor U2720 (N_2720,N_2608,N_2647);
or U2721 (N_2721,N_2656,N_2662);
or U2722 (N_2722,N_2639,N_2699);
xor U2723 (N_2723,N_2607,N_2638);
nor U2724 (N_2724,N_2609,N_2685);
nor U2725 (N_2725,N_2643,N_2687);
and U2726 (N_2726,N_2658,N_2693);
nor U2727 (N_2727,N_2688,N_2676);
nand U2728 (N_2728,N_2632,N_2652);
or U2729 (N_2729,N_2641,N_2640);
nor U2730 (N_2730,N_2601,N_2646);
and U2731 (N_2731,N_2695,N_2649);
or U2732 (N_2732,N_2684,N_2634);
or U2733 (N_2733,N_2697,N_2694);
and U2734 (N_2734,N_2681,N_2690);
nand U2735 (N_2735,N_2604,N_2625);
or U2736 (N_2736,N_2654,N_2653);
nand U2737 (N_2737,N_2650,N_2605);
or U2738 (N_2738,N_2680,N_2655);
and U2739 (N_2739,N_2659,N_2619);
nand U2740 (N_2740,N_2627,N_2616);
nand U2741 (N_2741,N_2644,N_2628);
or U2742 (N_2742,N_2672,N_2686);
nand U2743 (N_2743,N_2692,N_2621);
nor U2744 (N_2744,N_2637,N_2603);
and U2745 (N_2745,N_2660,N_2617);
xor U2746 (N_2746,N_2675,N_2664);
nand U2747 (N_2747,N_2624,N_2691);
or U2748 (N_2748,N_2671,N_2613);
and U2749 (N_2749,N_2666,N_2626);
and U2750 (N_2750,N_2630,N_2683);
nor U2751 (N_2751,N_2665,N_2682);
and U2752 (N_2752,N_2650,N_2644);
or U2753 (N_2753,N_2669,N_2628);
nand U2754 (N_2754,N_2659,N_2616);
and U2755 (N_2755,N_2699,N_2606);
nand U2756 (N_2756,N_2635,N_2687);
or U2757 (N_2757,N_2699,N_2684);
nor U2758 (N_2758,N_2663,N_2611);
and U2759 (N_2759,N_2625,N_2609);
nor U2760 (N_2760,N_2653,N_2675);
nor U2761 (N_2761,N_2664,N_2673);
or U2762 (N_2762,N_2654,N_2622);
or U2763 (N_2763,N_2612,N_2644);
and U2764 (N_2764,N_2637,N_2646);
or U2765 (N_2765,N_2632,N_2668);
nand U2766 (N_2766,N_2601,N_2687);
and U2767 (N_2767,N_2641,N_2662);
nor U2768 (N_2768,N_2628,N_2650);
nor U2769 (N_2769,N_2649,N_2686);
and U2770 (N_2770,N_2633,N_2631);
nor U2771 (N_2771,N_2657,N_2670);
nand U2772 (N_2772,N_2659,N_2657);
and U2773 (N_2773,N_2662,N_2618);
and U2774 (N_2774,N_2672,N_2691);
nor U2775 (N_2775,N_2607,N_2612);
or U2776 (N_2776,N_2629,N_2676);
or U2777 (N_2777,N_2692,N_2691);
nand U2778 (N_2778,N_2625,N_2670);
and U2779 (N_2779,N_2661,N_2662);
nand U2780 (N_2780,N_2686,N_2618);
and U2781 (N_2781,N_2687,N_2685);
nand U2782 (N_2782,N_2607,N_2688);
or U2783 (N_2783,N_2610,N_2633);
or U2784 (N_2784,N_2685,N_2603);
and U2785 (N_2785,N_2664,N_2606);
nor U2786 (N_2786,N_2624,N_2699);
and U2787 (N_2787,N_2615,N_2695);
nand U2788 (N_2788,N_2622,N_2665);
or U2789 (N_2789,N_2604,N_2628);
or U2790 (N_2790,N_2608,N_2643);
or U2791 (N_2791,N_2601,N_2605);
and U2792 (N_2792,N_2608,N_2630);
and U2793 (N_2793,N_2697,N_2613);
nor U2794 (N_2794,N_2672,N_2647);
or U2795 (N_2795,N_2619,N_2604);
or U2796 (N_2796,N_2608,N_2665);
or U2797 (N_2797,N_2677,N_2633);
and U2798 (N_2798,N_2691,N_2646);
nand U2799 (N_2799,N_2658,N_2648);
nand U2800 (N_2800,N_2797,N_2723);
nor U2801 (N_2801,N_2756,N_2736);
or U2802 (N_2802,N_2732,N_2784);
nor U2803 (N_2803,N_2777,N_2765);
nand U2804 (N_2804,N_2701,N_2754);
nand U2805 (N_2805,N_2793,N_2792);
nand U2806 (N_2806,N_2752,N_2720);
xor U2807 (N_2807,N_2761,N_2742);
nand U2808 (N_2808,N_2789,N_2748);
or U2809 (N_2809,N_2731,N_2711);
nand U2810 (N_2810,N_2781,N_2700);
or U2811 (N_2811,N_2747,N_2712);
nor U2812 (N_2812,N_2796,N_2729);
and U2813 (N_2813,N_2755,N_2713);
nor U2814 (N_2814,N_2745,N_2778);
and U2815 (N_2815,N_2714,N_2770);
and U2816 (N_2816,N_2790,N_2730);
or U2817 (N_2817,N_2750,N_2725);
or U2818 (N_2818,N_2721,N_2749);
or U2819 (N_2819,N_2716,N_2763);
nor U2820 (N_2820,N_2760,N_2746);
and U2821 (N_2821,N_2740,N_2709);
nor U2822 (N_2822,N_2726,N_2733);
or U2823 (N_2823,N_2785,N_2710);
nor U2824 (N_2824,N_2715,N_2705);
nor U2825 (N_2825,N_2771,N_2708);
nand U2826 (N_2826,N_2718,N_2767);
and U2827 (N_2827,N_2743,N_2786);
and U2828 (N_2828,N_2798,N_2772);
nor U2829 (N_2829,N_2727,N_2758);
nand U2830 (N_2830,N_2799,N_2741);
or U2831 (N_2831,N_2788,N_2764);
nor U2832 (N_2832,N_2769,N_2751);
nand U2833 (N_2833,N_2780,N_2774);
and U2834 (N_2834,N_2744,N_2794);
nand U2835 (N_2835,N_2738,N_2776);
or U2836 (N_2836,N_2779,N_2773);
nand U2837 (N_2837,N_2766,N_2707);
nand U2838 (N_2838,N_2759,N_2737);
xnor U2839 (N_2839,N_2724,N_2722);
and U2840 (N_2840,N_2739,N_2735);
and U2841 (N_2841,N_2703,N_2787);
and U2842 (N_2842,N_2719,N_2783);
or U2843 (N_2843,N_2734,N_2791);
nand U2844 (N_2844,N_2795,N_2762);
nor U2845 (N_2845,N_2753,N_2775);
and U2846 (N_2846,N_2704,N_2757);
and U2847 (N_2847,N_2717,N_2702);
nand U2848 (N_2848,N_2706,N_2768);
or U2849 (N_2849,N_2782,N_2728);
and U2850 (N_2850,N_2787,N_2754);
nand U2851 (N_2851,N_2779,N_2793);
and U2852 (N_2852,N_2702,N_2783);
and U2853 (N_2853,N_2720,N_2776);
nor U2854 (N_2854,N_2795,N_2759);
or U2855 (N_2855,N_2706,N_2753);
and U2856 (N_2856,N_2722,N_2762);
and U2857 (N_2857,N_2757,N_2797);
and U2858 (N_2858,N_2716,N_2702);
and U2859 (N_2859,N_2742,N_2727);
nand U2860 (N_2860,N_2702,N_2779);
and U2861 (N_2861,N_2780,N_2704);
nor U2862 (N_2862,N_2774,N_2791);
nor U2863 (N_2863,N_2748,N_2709);
nor U2864 (N_2864,N_2763,N_2705);
xor U2865 (N_2865,N_2764,N_2779);
or U2866 (N_2866,N_2702,N_2756);
and U2867 (N_2867,N_2717,N_2703);
nor U2868 (N_2868,N_2783,N_2701);
or U2869 (N_2869,N_2750,N_2793);
xnor U2870 (N_2870,N_2729,N_2731);
or U2871 (N_2871,N_2751,N_2759);
and U2872 (N_2872,N_2779,N_2726);
and U2873 (N_2873,N_2753,N_2713);
nand U2874 (N_2874,N_2756,N_2778);
nand U2875 (N_2875,N_2709,N_2764);
nand U2876 (N_2876,N_2704,N_2715);
or U2877 (N_2877,N_2761,N_2743);
nor U2878 (N_2878,N_2754,N_2751);
and U2879 (N_2879,N_2707,N_2725);
nor U2880 (N_2880,N_2770,N_2765);
or U2881 (N_2881,N_2787,N_2705);
nor U2882 (N_2882,N_2701,N_2773);
or U2883 (N_2883,N_2765,N_2729);
nor U2884 (N_2884,N_2794,N_2748);
nor U2885 (N_2885,N_2741,N_2757);
nor U2886 (N_2886,N_2772,N_2763);
or U2887 (N_2887,N_2757,N_2702);
nand U2888 (N_2888,N_2745,N_2726);
nand U2889 (N_2889,N_2723,N_2702);
xnor U2890 (N_2890,N_2744,N_2781);
nor U2891 (N_2891,N_2717,N_2724);
and U2892 (N_2892,N_2720,N_2784);
and U2893 (N_2893,N_2736,N_2787);
nor U2894 (N_2894,N_2787,N_2721);
and U2895 (N_2895,N_2704,N_2707);
nor U2896 (N_2896,N_2773,N_2767);
and U2897 (N_2897,N_2738,N_2775);
or U2898 (N_2898,N_2766,N_2732);
or U2899 (N_2899,N_2723,N_2788);
and U2900 (N_2900,N_2890,N_2881);
and U2901 (N_2901,N_2847,N_2823);
nor U2902 (N_2902,N_2865,N_2864);
or U2903 (N_2903,N_2820,N_2803);
nor U2904 (N_2904,N_2812,N_2888);
and U2905 (N_2905,N_2814,N_2829);
nand U2906 (N_2906,N_2878,N_2813);
or U2907 (N_2907,N_2856,N_2851);
nor U2908 (N_2908,N_2809,N_2882);
nor U2909 (N_2909,N_2853,N_2891);
and U2910 (N_2910,N_2863,N_2862);
nand U2911 (N_2911,N_2869,N_2824);
or U2912 (N_2912,N_2836,N_2806);
xor U2913 (N_2913,N_2840,N_2827);
and U2914 (N_2914,N_2826,N_2858);
nand U2915 (N_2915,N_2874,N_2821);
and U2916 (N_2916,N_2811,N_2831);
and U2917 (N_2917,N_2801,N_2868);
nand U2918 (N_2918,N_2807,N_2884);
and U2919 (N_2919,N_2867,N_2849);
and U2920 (N_2920,N_2854,N_2850);
nor U2921 (N_2921,N_2805,N_2837);
or U2922 (N_2922,N_2838,N_2872);
nand U2923 (N_2923,N_2830,N_2893);
and U2924 (N_2924,N_2841,N_2887);
or U2925 (N_2925,N_2816,N_2886);
and U2926 (N_2926,N_2839,N_2804);
or U2927 (N_2927,N_2898,N_2833);
nand U2928 (N_2928,N_2871,N_2859);
and U2929 (N_2929,N_2818,N_2895);
or U2930 (N_2930,N_2899,N_2835);
and U2931 (N_2931,N_2873,N_2832);
and U2932 (N_2932,N_2845,N_2896);
nand U2933 (N_2933,N_2844,N_2852);
or U2934 (N_2934,N_2857,N_2855);
or U2935 (N_2935,N_2870,N_2883);
and U2936 (N_2936,N_2861,N_2889);
nand U2937 (N_2937,N_2885,N_2822);
or U2938 (N_2938,N_2802,N_2828);
nor U2939 (N_2939,N_2825,N_2875);
and U2940 (N_2940,N_2817,N_2815);
nor U2941 (N_2941,N_2897,N_2810);
nor U2942 (N_2942,N_2800,N_2877);
nand U2943 (N_2943,N_2879,N_2842);
nand U2944 (N_2944,N_2819,N_2880);
and U2945 (N_2945,N_2848,N_2843);
or U2946 (N_2946,N_2894,N_2846);
nand U2947 (N_2947,N_2808,N_2860);
nand U2948 (N_2948,N_2892,N_2834);
or U2949 (N_2949,N_2876,N_2866);
nand U2950 (N_2950,N_2870,N_2810);
or U2951 (N_2951,N_2821,N_2851);
nor U2952 (N_2952,N_2895,N_2853);
or U2953 (N_2953,N_2821,N_2895);
nor U2954 (N_2954,N_2862,N_2880);
or U2955 (N_2955,N_2883,N_2877);
nand U2956 (N_2956,N_2851,N_2808);
and U2957 (N_2957,N_2803,N_2809);
or U2958 (N_2958,N_2874,N_2873);
nor U2959 (N_2959,N_2839,N_2871);
or U2960 (N_2960,N_2819,N_2897);
nand U2961 (N_2961,N_2869,N_2851);
or U2962 (N_2962,N_2815,N_2857);
or U2963 (N_2963,N_2800,N_2811);
nor U2964 (N_2964,N_2807,N_2817);
and U2965 (N_2965,N_2889,N_2885);
and U2966 (N_2966,N_2832,N_2847);
nor U2967 (N_2967,N_2810,N_2832);
nor U2968 (N_2968,N_2884,N_2892);
nand U2969 (N_2969,N_2862,N_2871);
nor U2970 (N_2970,N_2857,N_2804);
or U2971 (N_2971,N_2813,N_2828);
and U2972 (N_2972,N_2802,N_2827);
and U2973 (N_2973,N_2885,N_2855);
and U2974 (N_2974,N_2818,N_2809);
and U2975 (N_2975,N_2854,N_2827);
nand U2976 (N_2976,N_2828,N_2868);
or U2977 (N_2977,N_2891,N_2855);
nor U2978 (N_2978,N_2882,N_2864);
or U2979 (N_2979,N_2825,N_2862);
nor U2980 (N_2980,N_2839,N_2879);
nand U2981 (N_2981,N_2814,N_2894);
or U2982 (N_2982,N_2861,N_2883);
nor U2983 (N_2983,N_2837,N_2829);
and U2984 (N_2984,N_2862,N_2870);
nand U2985 (N_2985,N_2891,N_2828);
nand U2986 (N_2986,N_2847,N_2872);
or U2987 (N_2987,N_2844,N_2867);
xnor U2988 (N_2988,N_2882,N_2872);
nor U2989 (N_2989,N_2814,N_2877);
nand U2990 (N_2990,N_2811,N_2892);
and U2991 (N_2991,N_2861,N_2869);
and U2992 (N_2992,N_2844,N_2837);
xor U2993 (N_2993,N_2807,N_2847);
or U2994 (N_2994,N_2838,N_2808);
nand U2995 (N_2995,N_2865,N_2869);
or U2996 (N_2996,N_2896,N_2816);
or U2997 (N_2997,N_2834,N_2870);
nor U2998 (N_2998,N_2872,N_2893);
or U2999 (N_2999,N_2856,N_2838);
or U3000 (N_3000,N_2919,N_2944);
or U3001 (N_3001,N_2941,N_2918);
or U3002 (N_3002,N_2951,N_2913);
nand U3003 (N_3003,N_2992,N_2930);
or U3004 (N_3004,N_2987,N_2915);
nand U3005 (N_3005,N_2972,N_2957);
nand U3006 (N_3006,N_2947,N_2923);
nor U3007 (N_3007,N_2904,N_2960);
or U3008 (N_3008,N_2973,N_2953);
nor U3009 (N_3009,N_2924,N_2950);
nor U3010 (N_3010,N_2978,N_2909);
nor U3011 (N_3011,N_2917,N_2959);
xnor U3012 (N_3012,N_2990,N_2928);
nand U3013 (N_3013,N_2977,N_2916);
nor U3014 (N_3014,N_2908,N_2949);
xor U3015 (N_3015,N_2965,N_2989);
nand U3016 (N_3016,N_2932,N_2991);
nand U3017 (N_3017,N_2933,N_2921);
nand U3018 (N_3018,N_2926,N_2963);
nand U3019 (N_3019,N_2998,N_2912);
and U3020 (N_3020,N_2938,N_2961);
and U3021 (N_3021,N_2900,N_2970);
nand U3022 (N_3022,N_2993,N_2962);
and U3023 (N_3023,N_2925,N_2903);
nor U3024 (N_3024,N_2948,N_2939);
and U3025 (N_3025,N_2907,N_2964);
nand U3026 (N_3026,N_2979,N_2955);
and U3027 (N_3027,N_2968,N_2914);
and U3028 (N_3028,N_2942,N_2901);
nand U3029 (N_3029,N_2988,N_2980);
and U3030 (N_3030,N_2935,N_2995);
nor U3031 (N_3031,N_2986,N_2958);
or U3032 (N_3032,N_2952,N_2911);
nor U3033 (N_3033,N_2945,N_2985);
and U3034 (N_3034,N_2974,N_2984);
nand U3035 (N_3035,N_2975,N_2976);
nor U3036 (N_3036,N_2931,N_2967);
nor U3037 (N_3037,N_2943,N_2906);
nand U3038 (N_3038,N_2929,N_2971);
nand U3039 (N_3039,N_2940,N_2920);
or U3040 (N_3040,N_2910,N_2905);
and U3041 (N_3041,N_2994,N_2999);
nand U3042 (N_3042,N_2937,N_2936);
nand U3043 (N_3043,N_2922,N_2902);
nor U3044 (N_3044,N_2966,N_2954);
xnor U3045 (N_3045,N_2982,N_2983);
and U3046 (N_3046,N_2946,N_2927);
or U3047 (N_3047,N_2981,N_2934);
or U3048 (N_3048,N_2969,N_2997);
nand U3049 (N_3049,N_2956,N_2996);
nor U3050 (N_3050,N_2970,N_2966);
or U3051 (N_3051,N_2965,N_2956);
or U3052 (N_3052,N_2958,N_2956);
nor U3053 (N_3053,N_2918,N_2917);
and U3054 (N_3054,N_2952,N_2996);
nor U3055 (N_3055,N_2935,N_2978);
and U3056 (N_3056,N_2958,N_2906);
nand U3057 (N_3057,N_2982,N_2991);
or U3058 (N_3058,N_2968,N_2959);
nand U3059 (N_3059,N_2947,N_2907);
and U3060 (N_3060,N_2953,N_2967);
and U3061 (N_3061,N_2915,N_2965);
nor U3062 (N_3062,N_2936,N_2959);
and U3063 (N_3063,N_2993,N_2930);
nand U3064 (N_3064,N_2978,N_2988);
nor U3065 (N_3065,N_2940,N_2967);
and U3066 (N_3066,N_2989,N_2939);
nand U3067 (N_3067,N_2977,N_2959);
nor U3068 (N_3068,N_2961,N_2977);
and U3069 (N_3069,N_2907,N_2940);
and U3070 (N_3070,N_2934,N_2914);
nor U3071 (N_3071,N_2974,N_2987);
nor U3072 (N_3072,N_2958,N_2971);
or U3073 (N_3073,N_2947,N_2914);
nand U3074 (N_3074,N_2950,N_2928);
or U3075 (N_3075,N_2951,N_2924);
nand U3076 (N_3076,N_2955,N_2942);
nor U3077 (N_3077,N_2977,N_2991);
and U3078 (N_3078,N_2988,N_2900);
and U3079 (N_3079,N_2933,N_2978);
nor U3080 (N_3080,N_2966,N_2926);
nor U3081 (N_3081,N_2977,N_2979);
and U3082 (N_3082,N_2978,N_2959);
xnor U3083 (N_3083,N_2910,N_2988);
nor U3084 (N_3084,N_2930,N_2902);
nor U3085 (N_3085,N_2958,N_2936);
and U3086 (N_3086,N_2960,N_2987);
and U3087 (N_3087,N_2963,N_2967);
and U3088 (N_3088,N_2991,N_2902);
nand U3089 (N_3089,N_2997,N_2968);
or U3090 (N_3090,N_2901,N_2909);
and U3091 (N_3091,N_2921,N_2988);
nor U3092 (N_3092,N_2923,N_2922);
nand U3093 (N_3093,N_2962,N_2949);
nand U3094 (N_3094,N_2903,N_2952);
xor U3095 (N_3095,N_2932,N_2903);
and U3096 (N_3096,N_2912,N_2933);
and U3097 (N_3097,N_2968,N_2916);
or U3098 (N_3098,N_2983,N_2944);
or U3099 (N_3099,N_2945,N_2924);
or U3100 (N_3100,N_3011,N_3002);
or U3101 (N_3101,N_3091,N_3040);
nor U3102 (N_3102,N_3020,N_3030);
nor U3103 (N_3103,N_3043,N_3034);
or U3104 (N_3104,N_3061,N_3046);
or U3105 (N_3105,N_3098,N_3042);
or U3106 (N_3106,N_3082,N_3057);
and U3107 (N_3107,N_3048,N_3092);
or U3108 (N_3108,N_3050,N_3028);
and U3109 (N_3109,N_3053,N_3024);
nand U3110 (N_3110,N_3023,N_3003);
nand U3111 (N_3111,N_3086,N_3041);
nand U3112 (N_3112,N_3036,N_3087);
nand U3113 (N_3113,N_3083,N_3060);
nor U3114 (N_3114,N_3007,N_3063);
and U3115 (N_3115,N_3035,N_3045);
nor U3116 (N_3116,N_3068,N_3084);
and U3117 (N_3117,N_3051,N_3096);
and U3118 (N_3118,N_3081,N_3099);
or U3119 (N_3119,N_3052,N_3015);
nand U3120 (N_3120,N_3014,N_3025);
nor U3121 (N_3121,N_3064,N_3016);
nand U3122 (N_3122,N_3038,N_3027);
nand U3123 (N_3123,N_3010,N_3018);
nor U3124 (N_3124,N_3076,N_3072);
and U3125 (N_3125,N_3095,N_3039);
nand U3126 (N_3126,N_3067,N_3047);
or U3127 (N_3127,N_3013,N_3062);
or U3128 (N_3128,N_3026,N_3090);
and U3129 (N_3129,N_3001,N_3000);
or U3130 (N_3130,N_3073,N_3004);
nand U3131 (N_3131,N_3080,N_3066);
or U3132 (N_3132,N_3032,N_3009);
or U3133 (N_3133,N_3021,N_3078);
or U3134 (N_3134,N_3088,N_3085);
and U3135 (N_3135,N_3079,N_3097);
or U3136 (N_3136,N_3071,N_3093);
nand U3137 (N_3137,N_3069,N_3077);
nor U3138 (N_3138,N_3008,N_3058);
and U3139 (N_3139,N_3056,N_3022);
nand U3140 (N_3140,N_3044,N_3005);
nor U3141 (N_3141,N_3075,N_3049);
and U3142 (N_3142,N_3059,N_3033);
xor U3143 (N_3143,N_3094,N_3065);
nand U3144 (N_3144,N_3029,N_3006);
nand U3145 (N_3145,N_3070,N_3017);
or U3146 (N_3146,N_3089,N_3074);
and U3147 (N_3147,N_3054,N_3055);
and U3148 (N_3148,N_3031,N_3037);
or U3149 (N_3149,N_3019,N_3012);
nor U3150 (N_3150,N_3087,N_3066);
and U3151 (N_3151,N_3025,N_3028);
nand U3152 (N_3152,N_3037,N_3002);
and U3153 (N_3153,N_3001,N_3024);
nand U3154 (N_3154,N_3033,N_3087);
and U3155 (N_3155,N_3093,N_3003);
or U3156 (N_3156,N_3088,N_3044);
nor U3157 (N_3157,N_3017,N_3080);
or U3158 (N_3158,N_3050,N_3014);
nor U3159 (N_3159,N_3006,N_3017);
nor U3160 (N_3160,N_3010,N_3015);
nand U3161 (N_3161,N_3078,N_3032);
nand U3162 (N_3162,N_3079,N_3019);
nand U3163 (N_3163,N_3086,N_3040);
or U3164 (N_3164,N_3026,N_3050);
or U3165 (N_3165,N_3033,N_3048);
nor U3166 (N_3166,N_3028,N_3051);
nor U3167 (N_3167,N_3015,N_3012);
and U3168 (N_3168,N_3041,N_3064);
nand U3169 (N_3169,N_3021,N_3026);
nand U3170 (N_3170,N_3030,N_3068);
nor U3171 (N_3171,N_3073,N_3042);
or U3172 (N_3172,N_3013,N_3051);
or U3173 (N_3173,N_3074,N_3090);
or U3174 (N_3174,N_3043,N_3056);
or U3175 (N_3175,N_3051,N_3068);
nand U3176 (N_3176,N_3083,N_3041);
nand U3177 (N_3177,N_3098,N_3077);
or U3178 (N_3178,N_3036,N_3030);
nand U3179 (N_3179,N_3014,N_3082);
and U3180 (N_3180,N_3085,N_3050);
nor U3181 (N_3181,N_3057,N_3019);
or U3182 (N_3182,N_3093,N_3042);
nand U3183 (N_3183,N_3087,N_3015);
nand U3184 (N_3184,N_3050,N_3012);
or U3185 (N_3185,N_3040,N_3018);
and U3186 (N_3186,N_3058,N_3075);
and U3187 (N_3187,N_3057,N_3028);
nor U3188 (N_3188,N_3079,N_3023);
or U3189 (N_3189,N_3075,N_3040);
nor U3190 (N_3190,N_3024,N_3018);
nand U3191 (N_3191,N_3099,N_3072);
nor U3192 (N_3192,N_3028,N_3014);
nand U3193 (N_3193,N_3039,N_3052);
and U3194 (N_3194,N_3011,N_3027);
or U3195 (N_3195,N_3071,N_3039);
nand U3196 (N_3196,N_3032,N_3012);
xor U3197 (N_3197,N_3045,N_3065);
or U3198 (N_3198,N_3091,N_3068);
nand U3199 (N_3199,N_3034,N_3060);
or U3200 (N_3200,N_3142,N_3141);
nor U3201 (N_3201,N_3191,N_3115);
nor U3202 (N_3202,N_3124,N_3164);
or U3203 (N_3203,N_3155,N_3194);
nor U3204 (N_3204,N_3190,N_3111);
and U3205 (N_3205,N_3117,N_3160);
nand U3206 (N_3206,N_3113,N_3154);
nand U3207 (N_3207,N_3184,N_3179);
and U3208 (N_3208,N_3143,N_3180);
nand U3209 (N_3209,N_3168,N_3135);
and U3210 (N_3210,N_3101,N_3197);
or U3211 (N_3211,N_3116,N_3193);
and U3212 (N_3212,N_3167,N_3169);
and U3213 (N_3213,N_3196,N_3118);
nand U3214 (N_3214,N_3120,N_3173);
or U3215 (N_3215,N_3125,N_3134);
or U3216 (N_3216,N_3156,N_3165);
or U3217 (N_3217,N_3102,N_3105);
or U3218 (N_3218,N_3103,N_3177);
nand U3219 (N_3219,N_3159,N_3138);
nor U3220 (N_3220,N_3171,N_3178);
or U3221 (N_3221,N_3136,N_3140);
nor U3222 (N_3222,N_3137,N_3199);
nor U3223 (N_3223,N_3133,N_3185);
nor U3224 (N_3224,N_3128,N_3176);
nand U3225 (N_3225,N_3183,N_3153);
xnor U3226 (N_3226,N_3112,N_3148);
or U3227 (N_3227,N_3186,N_3139);
or U3228 (N_3228,N_3181,N_3130);
nor U3229 (N_3229,N_3129,N_3157);
or U3230 (N_3230,N_3161,N_3158);
and U3231 (N_3231,N_3107,N_3150);
nor U3232 (N_3232,N_3109,N_3172);
nand U3233 (N_3233,N_3121,N_3119);
nand U3234 (N_3234,N_3110,N_3188);
nand U3235 (N_3235,N_3187,N_3174);
nor U3236 (N_3236,N_3100,N_3198);
nand U3237 (N_3237,N_3146,N_3152);
and U3238 (N_3238,N_3149,N_3127);
nand U3239 (N_3239,N_3192,N_3126);
or U3240 (N_3240,N_3175,N_3123);
and U3241 (N_3241,N_3147,N_3163);
nand U3242 (N_3242,N_3122,N_3144);
or U3243 (N_3243,N_3108,N_3114);
nand U3244 (N_3244,N_3166,N_3195);
nand U3245 (N_3245,N_3106,N_3132);
and U3246 (N_3246,N_3151,N_3182);
or U3247 (N_3247,N_3145,N_3189);
or U3248 (N_3248,N_3104,N_3131);
xor U3249 (N_3249,N_3162,N_3170);
nand U3250 (N_3250,N_3131,N_3138);
or U3251 (N_3251,N_3140,N_3159);
nor U3252 (N_3252,N_3140,N_3160);
or U3253 (N_3253,N_3131,N_3114);
nor U3254 (N_3254,N_3137,N_3138);
nand U3255 (N_3255,N_3179,N_3165);
nand U3256 (N_3256,N_3187,N_3146);
or U3257 (N_3257,N_3190,N_3156);
nand U3258 (N_3258,N_3173,N_3159);
or U3259 (N_3259,N_3151,N_3171);
nor U3260 (N_3260,N_3113,N_3122);
and U3261 (N_3261,N_3138,N_3162);
nor U3262 (N_3262,N_3145,N_3171);
or U3263 (N_3263,N_3147,N_3139);
nor U3264 (N_3264,N_3169,N_3154);
nor U3265 (N_3265,N_3150,N_3170);
and U3266 (N_3266,N_3185,N_3149);
nand U3267 (N_3267,N_3107,N_3197);
nor U3268 (N_3268,N_3134,N_3126);
and U3269 (N_3269,N_3147,N_3198);
or U3270 (N_3270,N_3179,N_3151);
or U3271 (N_3271,N_3164,N_3134);
or U3272 (N_3272,N_3134,N_3141);
and U3273 (N_3273,N_3118,N_3149);
and U3274 (N_3274,N_3156,N_3136);
or U3275 (N_3275,N_3118,N_3170);
and U3276 (N_3276,N_3107,N_3118);
nor U3277 (N_3277,N_3199,N_3118);
and U3278 (N_3278,N_3109,N_3123);
nor U3279 (N_3279,N_3156,N_3178);
and U3280 (N_3280,N_3192,N_3107);
nor U3281 (N_3281,N_3158,N_3108);
and U3282 (N_3282,N_3161,N_3186);
nand U3283 (N_3283,N_3158,N_3133);
or U3284 (N_3284,N_3142,N_3174);
and U3285 (N_3285,N_3142,N_3157);
and U3286 (N_3286,N_3186,N_3127);
or U3287 (N_3287,N_3104,N_3119);
nor U3288 (N_3288,N_3168,N_3162);
and U3289 (N_3289,N_3196,N_3105);
nor U3290 (N_3290,N_3156,N_3171);
nand U3291 (N_3291,N_3184,N_3186);
and U3292 (N_3292,N_3128,N_3181);
or U3293 (N_3293,N_3153,N_3135);
nand U3294 (N_3294,N_3134,N_3181);
nor U3295 (N_3295,N_3101,N_3175);
nand U3296 (N_3296,N_3195,N_3171);
nor U3297 (N_3297,N_3175,N_3116);
and U3298 (N_3298,N_3173,N_3145);
or U3299 (N_3299,N_3141,N_3119);
nor U3300 (N_3300,N_3297,N_3276);
nor U3301 (N_3301,N_3257,N_3273);
nor U3302 (N_3302,N_3205,N_3224);
and U3303 (N_3303,N_3258,N_3294);
nor U3304 (N_3304,N_3209,N_3238);
nor U3305 (N_3305,N_3261,N_3259);
nand U3306 (N_3306,N_3225,N_3260);
and U3307 (N_3307,N_3208,N_3240);
and U3308 (N_3308,N_3287,N_3242);
or U3309 (N_3309,N_3229,N_3206);
nor U3310 (N_3310,N_3256,N_3289);
and U3311 (N_3311,N_3280,N_3252);
and U3312 (N_3312,N_3239,N_3200);
and U3313 (N_3313,N_3223,N_3274);
nor U3314 (N_3314,N_3275,N_3207);
and U3315 (N_3315,N_3285,N_3216);
and U3316 (N_3316,N_3266,N_3268);
and U3317 (N_3317,N_3211,N_3288);
or U3318 (N_3318,N_3254,N_3228);
or U3319 (N_3319,N_3226,N_3299);
nor U3320 (N_3320,N_3210,N_3241);
nand U3321 (N_3321,N_3269,N_3230);
or U3322 (N_3322,N_3233,N_3227);
nor U3323 (N_3323,N_3246,N_3296);
or U3324 (N_3324,N_3215,N_3267);
or U3325 (N_3325,N_3231,N_3286);
and U3326 (N_3326,N_3284,N_3250);
nand U3327 (N_3327,N_3219,N_3248);
nor U3328 (N_3328,N_3237,N_3277);
or U3329 (N_3329,N_3235,N_3247);
nor U3330 (N_3330,N_3243,N_3220);
nand U3331 (N_3331,N_3214,N_3201);
nor U3332 (N_3332,N_3281,N_3222);
nand U3333 (N_3333,N_3295,N_3283);
nand U3334 (N_3334,N_3204,N_3272);
or U3335 (N_3335,N_3232,N_3264);
nor U3336 (N_3336,N_3221,N_3202);
and U3337 (N_3337,N_3282,N_3278);
nand U3338 (N_3338,N_3290,N_3298);
xor U3339 (N_3339,N_3249,N_3279);
or U3340 (N_3340,N_3271,N_3253);
nor U3341 (N_3341,N_3218,N_3203);
nand U3342 (N_3342,N_3244,N_3234);
and U3343 (N_3343,N_3265,N_3213);
nor U3344 (N_3344,N_3262,N_3270);
nor U3345 (N_3345,N_3217,N_3251);
and U3346 (N_3346,N_3212,N_3263);
or U3347 (N_3347,N_3291,N_3293);
nand U3348 (N_3348,N_3245,N_3292);
nand U3349 (N_3349,N_3255,N_3236);
nand U3350 (N_3350,N_3256,N_3241);
and U3351 (N_3351,N_3261,N_3254);
or U3352 (N_3352,N_3222,N_3285);
nor U3353 (N_3353,N_3262,N_3247);
or U3354 (N_3354,N_3246,N_3285);
nor U3355 (N_3355,N_3276,N_3257);
nor U3356 (N_3356,N_3209,N_3297);
nand U3357 (N_3357,N_3259,N_3293);
nor U3358 (N_3358,N_3267,N_3249);
or U3359 (N_3359,N_3241,N_3272);
and U3360 (N_3360,N_3288,N_3278);
nand U3361 (N_3361,N_3206,N_3231);
or U3362 (N_3362,N_3224,N_3262);
or U3363 (N_3363,N_3286,N_3241);
or U3364 (N_3364,N_3236,N_3237);
or U3365 (N_3365,N_3250,N_3242);
nand U3366 (N_3366,N_3261,N_3267);
or U3367 (N_3367,N_3272,N_3243);
xor U3368 (N_3368,N_3293,N_3285);
and U3369 (N_3369,N_3213,N_3280);
or U3370 (N_3370,N_3270,N_3255);
and U3371 (N_3371,N_3293,N_3252);
or U3372 (N_3372,N_3224,N_3230);
or U3373 (N_3373,N_3264,N_3223);
nor U3374 (N_3374,N_3237,N_3214);
nand U3375 (N_3375,N_3200,N_3276);
nor U3376 (N_3376,N_3219,N_3225);
or U3377 (N_3377,N_3292,N_3260);
nand U3378 (N_3378,N_3201,N_3253);
nor U3379 (N_3379,N_3264,N_3206);
and U3380 (N_3380,N_3211,N_3246);
nor U3381 (N_3381,N_3211,N_3226);
nand U3382 (N_3382,N_3259,N_3286);
nand U3383 (N_3383,N_3249,N_3223);
nand U3384 (N_3384,N_3255,N_3250);
nand U3385 (N_3385,N_3277,N_3243);
xor U3386 (N_3386,N_3250,N_3249);
nand U3387 (N_3387,N_3277,N_3205);
and U3388 (N_3388,N_3251,N_3289);
or U3389 (N_3389,N_3263,N_3296);
nor U3390 (N_3390,N_3236,N_3299);
or U3391 (N_3391,N_3289,N_3286);
nand U3392 (N_3392,N_3270,N_3231);
nand U3393 (N_3393,N_3291,N_3231);
and U3394 (N_3394,N_3294,N_3249);
nand U3395 (N_3395,N_3299,N_3294);
nor U3396 (N_3396,N_3271,N_3250);
nand U3397 (N_3397,N_3206,N_3296);
nor U3398 (N_3398,N_3260,N_3230);
nor U3399 (N_3399,N_3292,N_3272);
or U3400 (N_3400,N_3326,N_3310);
nor U3401 (N_3401,N_3359,N_3353);
nand U3402 (N_3402,N_3355,N_3388);
nand U3403 (N_3403,N_3352,N_3313);
xor U3404 (N_3404,N_3368,N_3373);
or U3405 (N_3405,N_3354,N_3374);
nor U3406 (N_3406,N_3340,N_3312);
nand U3407 (N_3407,N_3362,N_3363);
nor U3408 (N_3408,N_3319,N_3398);
nor U3409 (N_3409,N_3346,N_3307);
and U3410 (N_3410,N_3330,N_3311);
nand U3411 (N_3411,N_3348,N_3391);
or U3412 (N_3412,N_3357,N_3304);
or U3413 (N_3413,N_3360,N_3338);
and U3414 (N_3414,N_3397,N_3314);
nor U3415 (N_3415,N_3308,N_3320);
nor U3416 (N_3416,N_3393,N_3335);
or U3417 (N_3417,N_3392,N_3370);
xnor U3418 (N_3418,N_3331,N_3358);
nor U3419 (N_3419,N_3336,N_3316);
or U3420 (N_3420,N_3377,N_3364);
nor U3421 (N_3421,N_3379,N_3317);
nand U3422 (N_3422,N_3387,N_3396);
or U3423 (N_3423,N_3356,N_3386);
and U3424 (N_3424,N_3375,N_3361);
and U3425 (N_3425,N_3347,N_3380);
or U3426 (N_3426,N_3329,N_3301);
and U3427 (N_3427,N_3385,N_3306);
nor U3428 (N_3428,N_3321,N_3327);
nand U3429 (N_3429,N_3376,N_3365);
and U3430 (N_3430,N_3341,N_3344);
nor U3431 (N_3431,N_3324,N_3332);
and U3432 (N_3432,N_3372,N_3305);
xnor U3433 (N_3433,N_3309,N_3384);
nand U3434 (N_3434,N_3378,N_3333);
nor U3435 (N_3435,N_3315,N_3366);
or U3436 (N_3436,N_3334,N_3371);
nand U3437 (N_3437,N_3399,N_3350);
nor U3438 (N_3438,N_3381,N_3369);
or U3439 (N_3439,N_3343,N_3318);
nor U3440 (N_3440,N_3303,N_3367);
nor U3441 (N_3441,N_3325,N_3390);
and U3442 (N_3442,N_3339,N_3323);
nor U3443 (N_3443,N_3389,N_3383);
nor U3444 (N_3444,N_3337,N_3345);
and U3445 (N_3445,N_3342,N_3322);
and U3446 (N_3446,N_3300,N_3351);
nand U3447 (N_3447,N_3302,N_3394);
or U3448 (N_3448,N_3328,N_3382);
or U3449 (N_3449,N_3395,N_3349);
nand U3450 (N_3450,N_3375,N_3329);
and U3451 (N_3451,N_3338,N_3365);
and U3452 (N_3452,N_3391,N_3310);
and U3453 (N_3453,N_3349,N_3310);
or U3454 (N_3454,N_3381,N_3367);
nand U3455 (N_3455,N_3363,N_3367);
nor U3456 (N_3456,N_3394,N_3367);
and U3457 (N_3457,N_3341,N_3330);
or U3458 (N_3458,N_3328,N_3347);
and U3459 (N_3459,N_3376,N_3326);
and U3460 (N_3460,N_3313,N_3343);
and U3461 (N_3461,N_3381,N_3319);
nor U3462 (N_3462,N_3364,N_3320);
and U3463 (N_3463,N_3351,N_3334);
nor U3464 (N_3464,N_3384,N_3348);
nand U3465 (N_3465,N_3386,N_3379);
nor U3466 (N_3466,N_3342,N_3385);
or U3467 (N_3467,N_3325,N_3310);
nor U3468 (N_3468,N_3305,N_3398);
nand U3469 (N_3469,N_3372,N_3330);
nor U3470 (N_3470,N_3300,N_3324);
and U3471 (N_3471,N_3373,N_3326);
nand U3472 (N_3472,N_3340,N_3360);
or U3473 (N_3473,N_3328,N_3384);
or U3474 (N_3474,N_3381,N_3309);
nor U3475 (N_3475,N_3386,N_3327);
xnor U3476 (N_3476,N_3325,N_3356);
nor U3477 (N_3477,N_3340,N_3334);
and U3478 (N_3478,N_3323,N_3377);
or U3479 (N_3479,N_3302,N_3326);
nor U3480 (N_3480,N_3380,N_3393);
xor U3481 (N_3481,N_3300,N_3312);
or U3482 (N_3482,N_3370,N_3303);
nand U3483 (N_3483,N_3364,N_3342);
xnor U3484 (N_3484,N_3386,N_3323);
and U3485 (N_3485,N_3335,N_3332);
nor U3486 (N_3486,N_3304,N_3390);
and U3487 (N_3487,N_3314,N_3300);
or U3488 (N_3488,N_3360,N_3366);
and U3489 (N_3489,N_3304,N_3318);
nand U3490 (N_3490,N_3311,N_3309);
nand U3491 (N_3491,N_3321,N_3372);
nand U3492 (N_3492,N_3321,N_3343);
nand U3493 (N_3493,N_3306,N_3330);
and U3494 (N_3494,N_3316,N_3357);
or U3495 (N_3495,N_3356,N_3349);
and U3496 (N_3496,N_3337,N_3336);
or U3497 (N_3497,N_3381,N_3361);
nand U3498 (N_3498,N_3341,N_3333);
nand U3499 (N_3499,N_3309,N_3366);
nand U3500 (N_3500,N_3440,N_3485);
nand U3501 (N_3501,N_3450,N_3421);
nand U3502 (N_3502,N_3408,N_3461);
and U3503 (N_3503,N_3413,N_3488);
and U3504 (N_3504,N_3458,N_3424);
or U3505 (N_3505,N_3427,N_3460);
and U3506 (N_3506,N_3415,N_3425);
nand U3507 (N_3507,N_3482,N_3467);
nand U3508 (N_3508,N_3405,N_3400);
or U3509 (N_3509,N_3464,N_3484);
nor U3510 (N_3510,N_3428,N_3471);
or U3511 (N_3511,N_3445,N_3456);
and U3512 (N_3512,N_3468,N_3419);
nand U3513 (N_3513,N_3420,N_3431);
or U3514 (N_3514,N_3406,N_3443);
and U3515 (N_3515,N_3469,N_3414);
and U3516 (N_3516,N_3491,N_3483);
and U3517 (N_3517,N_3496,N_3418);
or U3518 (N_3518,N_3490,N_3470);
or U3519 (N_3519,N_3474,N_3410);
and U3520 (N_3520,N_3486,N_3439);
and U3521 (N_3521,N_3442,N_3452);
or U3522 (N_3522,N_3479,N_3416);
nor U3523 (N_3523,N_3459,N_3473);
nand U3524 (N_3524,N_3407,N_3478);
nor U3525 (N_3525,N_3423,N_3417);
and U3526 (N_3526,N_3465,N_3476);
and U3527 (N_3527,N_3437,N_3487);
or U3528 (N_3528,N_3433,N_3454);
and U3529 (N_3529,N_3436,N_3475);
nor U3530 (N_3530,N_3497,N_3426);
and U3531 (N_3531,N_3477,N_3480);
and U3532 (N_3532,N_3489,N_3455);
or U3533 (N_3533,N_3457,N_3498);
nand U3534 (N_3534,N_3449,N_3401);
and U3535 (N_3535,N_3494,N_3409);
nor U3536 (N_3536,N_3481,N_3462);
or U3537 (N_3537,N_3472,N_3435);
nand U3538 (N_3538,N_3429,N_3412);
nand U3539 (N_3539,N_3403,N_3404);
and U3540 (N_3540,N_3430,N_3492);
or U3541 (N_3541,N_3422,N_3499);
nor U3542 (N_3542,N_3432,N_3434);
nand U3543 (N_3543,N_3453,N_3446);
and U3544 (N_3544,N_3438,N_3493);
nor U3545 (N_3545,N_3448,N_3447);
nor U3546 (N_3546,N_3444,N_3411);
and U3547 (N_3547,N_3466,N_3463);
nor U3548 (N_3548,N_3402,N_3495);
or U3549 (N_3549,N_3451,N_3441);
nand U3550 (N_3550,N_3404,N_3433);
nor U3551 (N_3551,N_3480,N_3487);
nand U3552 (N_3552,N_3427,N_3410);
nand U3553 (N_3553,N_3430,N_3439);
and U3554 (N_3554,N_3467,N_3435);
or U3555 (N_3555,N_3446,N_3499);
nand U3556 (N_3556,N_3480,N_3499);
or U3557 (N_3557,N_3451,N_3416);
nor U3558 (N_3558,N_3463,N_3400);
nand U3559 (N_3559,N_3492,N_3461);
and U3560 (N_3560,N_3434,N_3448);
nor U3561 (N_3561,N_3466,N_3419);
and U3562 (N_3562,N_3435,N_3481);
nor U3563 (N_3563,N_3458,N_3441);
nand U3564 (N_3564,N_3467,N_3445);
nand U3565 (N_3565,N_3446,N_3406);
nand U3566 (N_3566,N_3465,N_3417);
and U3567 (N_3567,N_3432,N_3417);
nand U3568 (N_3568,N_3463,N_3488);
nand U3569 (N_3569,N_3489,N_3498);
nand U3570 (N_3570,N_3438,N_3404);
nand U3571 (N_3571,N_3482,N_3433);
xnor U3572 (N_3572,N_3409,N_3468);
nand U3573 (N_3573,N_3470,N_3400);
nor U3574 (N_3574,N_3401,N_3403);
nor U3575 (N_3575,N_3473,N_3454);
or U3576 (N_3576,N_3485,N_3449);
or U3577 (N_3577,N_3406,N_3461);
or U3578 (N_3578,N_3489,N_3467);
and U3579 (N_3579,N_3487,N_3414);
and U3580 (N_3580,N_3409,N_3467);
nand U3581 (N_3581,N_3408,N_3448);
nor U3582 (N_3582,N_3460,N_3474);
nand U3583 (N_3583,N_3404,N_3436);
nor U3584 (N_3584,N_3412,N_3472);
or U3585 (N_3585,N_3460,N_3491);
or U3586 (N_3586,N_3425,N_3468);
or U3587 (N_3587,N_3425,N_3481);
nor U3588 (N_3588,N_3450,N_3466);
and U3589 (N_3589,N_3468,N_3485);
nor U3590 (N_3590,N_3495,N_3444);
and U3591 (N_3591,N_3409,N_3416);
and U3592 (N_3592,N_3485,N_3495);
or U3593 (N_3593,N_3459,N_3481);
nor U3594 (N_3594,N_3401,N_3407);
and U3595 (N_3595,N_3401,N_3400);
nand U3596 (N_3596,N_3423,N_3435);
nand U3597 (N_3597,N_3404,N_3458);
nor U3598 (N_3598,N_3438,N_3498);
or U3599 (N_3599,N_3439,N_3460);
nor U3600 (N_3600,N_3589,N_3526);
or U3601 (N_3601,N_3561,N_3515);
and U3602 (N_3602,N_3502,N_3500);
and U3603 (N_3603,N_3555,N_3522);
nor U3604 (N_3604,N_3575,N_3568);
or U3605 (N_3605,N_3563,N_3552);
nand U3606 (N_3606,N_3533,N_3536);
nand U3607 (N_3607,N_3543,N_3534);
nand U3608 (N_3608,N_3540,N_3514);
nor U3609 (N_3609,N_3516,N_3544);
or U3610 (N_3610,N_3505,N_3545);
and U3611 (N_3611,N_3523,N_3569);
nand U3612 (N_3612,N_3509,N_3588);
or U3613 (N_3613,N_3504,N_3554);
or U3614 (N_3614,N_3530,N_3524);
or U3615 (N_3615,N_3513,N_3587);
xnor U3616 (N_3616,N_3518,N_3586);
or U3617 (N_3617,N_3538,N_3598);
nor U3618 (N_3618,N_3594,N_3584);
or U3619 (N_3619,N_3550,N_3542);
and U3620 (N_3620,N_3508,N_3501);
and U3621 (N_3621,N_3559,N_3507);
and U3622 (N_3622,N_3592,N_3581);
nor U3623 (N_3623,N_3573,N_3539);
nand U3624 (N_3624,N_3570,N_3517);
nand U3625 (N_3625,N_3510,N_3557);
and U3626 (N_3626,N_3549,N_3503);
nand U3627 (N_3627,N_3566,N_3585);
or U3628 (N_3628,N_3565,N_3551);
nand U3629 (N_3629,N_3558,N_3519);
and U3630 (N_3630,N_3564,N_3511);
nor U3631 (N_3631,N_3571,N_3577);
nand U3632 (N_3632,N_3580,N_3553);
nor U3633 (N_3633,N_3579,N_3572);
nand U3634 (N_3634,N_3531,N_3529);
and U3635 (N_3635,N_3527,N_3597);
nor U3636 (N_3636,N_3591,N_3547);
or U3637 (N_3637,N_3582,N_3595);
or U3638 (N_3638,N_3593,N_3520);
xor U3639 (N_3639,N_3576,N_3574);
or U3640 (N_3640,N_3562,N_3583);
nor U3641 (N_3641,N_3556,N_3567);
nand U3642 (N_3642,N_3578,N_3512);
nand U3643 (N_3643,N_3599,N_3537);
nand U3644 (N_3644,N_3541,N_3532);
and U3645 (N_3645,N_3548,N_3506);
and U3646 (N_3646,N_3596,N_3521);
and U3647 (N_3647,N_3528,N_3535);
or U3648 (N_3648,N_3546,N_3525);
nor U3649 (N_3649,N_3590,N_3560);
and U3650 (N_3650,N_3519,N_3525);
and U3651 (N_3651,N_3510,N_3523);
or U3652 (N_3652,N_3506,N_3559);
or U3653 (N_3653,N_3533,N_3528);
nor U3654 (N_3654,N_3558,N_3566);
nand U3655 (N_3655,N_3558,N_3589);
nand U3656 (N_3656,N_3505,N_3579);
nand U3657 (N_3657,N_3536,N_3552);
and U3658 (N_3658,N_3572,N_3529);
nand U3659 (N_3659,N_3539,N_3556);
nand U3660 (N_3660,N_3508,N_3555);
nor U3661 (N_3661,N_3556,N_3538);
or U3662 (N_3662,N_3523,N_3594);
nand U3663 (N_3663,N_3540,N_3568);
and U3664 (N_3664,N_3563,N_3545);
nand U3665 (N_3665,N_3563,N_3511);
nand U3666 (N_3666,N_3572,N_3557);
nor U3667 (N_3667,N_3563,N_3597);
nor U3668 (N_3668,N_3508,N_3519);
nor U3669 (N_3669,N_3564,N_3537);
and U3670 (N_3670,N_3546,N_3527);
or U3671 (N_3671,N_3503,N_3578);
or U3672 (N_3672,N_3555,N_3532);
or U3673 (N_3673,N_3574,N_3598);
and U3674 (N_3674,N_3503,N_3531);
or U3675 (N_3675,N_3596,N_3532);
and U3676 (N_3676,N_3503,N_3547);
nand U3677 (N_3677,N_3590,N_3527);
nand U3678 (N_3678,N_3508,N_3542);
and U3679 (N_3679,N_3504,N_3528);
nor U3680 (N_3680,N_3581,N_3582);
and U3681 (N_3681,N_3585,N_3549);
and U3682 (N_3682,N_3517,N_3559);
and U3683 (N_3683,N_3518,N_3516);
nor U3684 (N_3684,N_3574,N_3553);
or U3685 (N_3685,N_3510,N_3548);
and U3686 (N_3686,N_3575,N_3534);
nand U3687 (N_3687,N_3528,N_3522);
nor U3688 (N_3688,N_3594,N_3533);
or U3689 (N_3689,N_3509,N_3559);
nand U3690 (N_3690,N_3570,N_3580);
and U3691 (N_3691,N_3533,N_3539);
or U3692 (N_3692,N_3592,N_3582);
nand U3693 (N_3693,N_3576,N_3545);
or U3694 (N_3694,N_3579,N_3504);
or U3695 (N_3695,N_3554,N_3579);
and U3696 (N_3696,N_3557,N_3532);
nor U3697 (N_3697,N_3502,N_3552);
and U3698 (N_3698,N_3553,N_3577);
and U3699 (N_3699,N_3520,N_3541);
or U3700 (N_3700,N_3698,N_3629);
nand U3701 (N_3701,N_3628,N_3643);
or U3702 (N_3702,N_3666,N_3631);
or U3703 (N_3703,N_3665,N_3684);
nand U3704 (N_3704,N_3675,N_3606);
nand U3705 (N_3705,N_3625,N_3634);
xor U3706 (N_3706,N_3621,N_3679);
nand U3707 (N_3707,N_3689,N_3630);
and U3708 (N_3708,N_3640,N_3607);
nor U3709 (N_3709,N_3641,N_3657);
or U3710 (N_3710,N_3618,N_3610);
and U3711 (N_3711,N_3697,N_3623);
and U3712 (N_3712,N_3619,N_3680);
or U3713 (N_3713,N_3636,N_3635);
nor U3714 (N_3714,N_3661,N_3674);
and U3715 (N_3715,N_3622,N_3627);
nand U3716 (N_3716,N_3603,N_3696);
nand U3717 (N_3717,N_3681,N_3649);
nor U3718 (N_3718,N_3695,N_3650);
nand U3719 (N_3719,N_3652,N_3656);
nor U3720 (N_3720,N_3609,N_3671);
or U3721 (N_3721,N_3678,N_3692);
or U3722 (N_3722,N_3672,N_3617);
nand U3723 (N_3723,N_3653,N_3601);
nand U3724 (N_3724,N_3655,N_3615);
and U3725 (N_3725,N_3647,N_3626);
nand U3726 (N_3726,N_3600,N_3658);
nor U3727 (N_3727,N_3668,N_3673);
or U3728 (N_3728,N_3604,N_3687);
nand U3729 (N_3729,N_3693,N_3645);
nor U3730 (N_3730,N_3659,N_3667);
and U3731 (N_3731,N_3613,N_3691);
nand U3732 (N_3732,N_3639,N_3614);
nor U3733 (N_3733,N_3648,N_3677);
nor U3734 (N_3734,N_3620,N_3664);
and U3735 (N_3735,N_3685,N_3663);
nor U3736 (N_3736,N_3690,N_3669);
xnor U3737 (N_3737,N_3660,N_3632);
nand U3738 (N_3738,N_3654,N_3608);
nor U3739 (N_3739,N_3611,N_3612);
nand U3740 (N_3740,N_3686,N_3633);
or U3741 (N_3741,N_3644,N_3646);
and U3742 (N_3742,N_3638,N_3642);
nand U3743 (N_3743,N_3694,N_3682);
and U3744 (N_3744,N_3616,N_3605);
or U3745 (N_3745,N_3602,N_3637);
nor U3746 (N_3746,N_3662,N_3683);
or U3747 (N_3747,N_3676,N_3670);
or U3748 (N_3748,N_3699,N_3688);
nor U3749 (N_3749,N_3624,N_3651);
or U3750 (N_3750,N_3660,N_3622);
nand U3751 (N_3751,N_3602,N_3634);
nand U3752 (N_3752,N_3621,N_3624);
and U3753 (N_3753,N_3659,N_3676);
xnor U3754 (N_3754,N_3606,N_3699);
and U3755 (N_3755,N_3689,N_3626);
and U3756 (N_3756,N_3699,N_3638);
nor U3757 (N_3757,N_3639,N_3697);
and U3758 (N_3758,N_3609,N_3652);
and U3759 (N_3759,N_3650,N_3642);
and U3760 (N_3760,N_3628,N_3678);
nor U3761 (N_3761,N_3600,N_3686);
nor U3762 (N_3762,N_3656,N_3614);
nor U3763 (N_3763,N_3673,N_3633);
and U3764 (N_3764,N_3619,N_3666);
or U3765 (N_3765,N_3685,N_3610);
or U3766 (N_3766,N_3677,N_3614);
or U3767 (N_3767,N_3648,N_3643);
and U3768 (N_3768,N_3690,N_3644);
and U3769 (N_3769,N_3675,N_3662);
nand U3770 (N_3770,N_3626,N_3634);
nor U3771 (N_3771,N_3673,N_3623);
or U3772 (N_3772,N_3684,N_3674);
nor U3773 (N_3773,N_3694,N_3642);
nor U3774 (N_3774,N_3687,N_3695);
and U3775 (N_3775,N_3685,N_3604);
nor U3776 (N_3776,N_3676,N_3616);
xnor U3777 (N_3777,N_3674,N_3640);
nor U3778 (N_3778,N_3686,N_3681);
or U3779 (N_3779,N_3608,N_3614);
and U3780 (N_3780,N_3697,N_3681);
and U3781 (N_3781,N_3620,N_3658);
and U3782 (N_3782,N_3643,N_3650);
or U3783 (N_3783,N_3646,N_3670);
and U3784 (N_3784,N_3661,N_3644);
or U3785 (N_3785,N_3613,N_3624);
nor U3786 (N_3786,N_3617,N_3690);
or U3787 (N_3787,N_3601,N_3621);
and U3788 (N_3788,N_3632,N_3696);
or U3789 (N_3789,N_3688,N_3671);
nand U3790 (N_3790,N_3686,N_3668);
or U3791 (N_3791,N_3694,N_3629);
nand U3792 (N_3792,N_3675,N_3626);
or U3793 (N_3793,N_3649,N_3659);
or U3794 (N_3794,N_3691,N_3651);
xnor U3795 (N_3795,N_3644,N_3610);
and U3796 (N_3796,N_3640,N_3645);
nand U3797 (N_3797,N_3601,N_3648);
nand U3798 (N_3798,N_3682,N_3688);
nand U3799 (N_3799,N_3657,N_3619);
nand U3800 (N_3800,N_3781,N_3763);
nor U3801 (N_3801,N_3792,N_3757);
nor U3802 (N_3802,N_3770,N_3779);
and U3803 (N_3803,N_3725,N_3798);
and U3804 (N_3804,N_3794,N_3704);
or U3805 (N_3805,N_3773,N_3761);
nand U3806 (N_3806,N_3769,N_3743);
or U3807 (N_3807,N_3724,N_3739);
xor U3808 (N_3808,N_3742,N_3722);
nor U3809 (N_3809,N_3787,N_3728);
and U3810 (N_3810,N_3786,N_3741);
nand U3811 (N_3811,N_3712,N_3727);
nor U3812 (N_3812,N_3780,N_3784);
nor U3813 (N_3813,N_3726,N_3789);
nand U3814 (N_3814,N_3710,N_3716);
nor U3815 (N_3815,N_3777,N_3721);
and U3816 (N_3816,N_3783,N_3796);
nor U3817 (N_3817,N_3747,N_3745);
and U3818 (N_3818,N_3740,N_3731);
or U3819 (N_3819,N_3701,N_3799);
or U3820 (N_3820,N_3776,N_3746);
and U3821 (N_3821,N_3713,N_3775);
or U3822 (N_3822,N_3702,N_3749);
nor U3823 (N_3823,N_3730,N_3760);
or U3824 (N_3824,N_3772,N_3790);
and U3825 (N_3825,N_3720,N_3766);
and U3826 (N_3826,N_3737,N_3765);
or U3827 (N_3827,N_3729,N_3778);
or U3828 (N_3828,N_3764,N_3756);
and U3829 (N_3829,N_3793,N_3706);
xnor U3830 (N_3830,N_3703,N_3791);
or U3831 (N_3831,N_3758,N_3759);
nor U3832 (N_3832,N_3782,N_3762);
nor U3833 (N_3833,N_3797,N_3768);
nand U3834 (N_3834,N_3717,N_3715);
or U3835 (N_3835,N_3708,N_3732);
nand U3836 (N_3836,N_3774,N_3707);
or U3837 (N_3837,N_3736,N_3735);
nand U3838 (N_3838,N_3711,N_3700);
and U3839 (N_3839,N_3788,N_3748);
and U3840 (N_3840,N_3785,N_3714);
nand U3841 (N_3841,N_3723,N_3754);
and U3842 (N_3842,N_3752,N_3767);
nand U3843 (N_3843,N_3733,N_3709);
or U3844 (N_3844,N_3719,N_3750);
nand U3845 (N_3845,N_3734,N_3718);
nor U3846 (N_3846,N_3705,N_3751);
nor U3847 (N_3847,N_3738,N_3771);
or U3848 (N_3848,N_3753,N_3795);
or U3849 (N_3849,N_3744,N_3755);
or U3850 (N_3850,N_3711,N_3729);
or U3851 (N_3851,N_3718,N_3754);
nand U3852 (N_3852,N_3749,N_3733);
nand U3853 (N_3853,N_3783,N_3788);
nor U3854 (N_3854,N_3722,N_3720);
nand U3855 (N_3855,N_3797,N_3712);
nor U3856 (N_3856,N_3741,N_3743);
or U3857 (N_3857,N_3751,N_3731);
or U3858 (N_3858,N_3710,N_3738);
or U3859 (N_3859,N_3759,N_3783);
nand U3860 (N_3860,N_3703,N_3787);
or U3861 (N_3861,N_3733,N_3721);
xnor U3862 (N_3862,N_3709,N_3742);
or U3863 (N_3863,N_3740,N_3738);
nor U3864 (N_3864,N_3701,N_3705);
and U3865 (N_3865,N_3774,N_3728);
or U3866 (N_3866,N_3744,N_3737);
xnor U3867 (N_3867,N_3701,N_3747);
nor U3868 (N_3868,N_3747,N_3744);
nor U3869 (N_3869,N_3789,N_3759);
or U3870 (N_3870,N_3752,N_3732);
and U3871 (N_3871,N_3794,N_3772);
and U3872 (N_3872,N_3755,N_3790);
nor U3873 (N_3873,N_3768,N_3738);
nand U3874 (N_3874,N_3706,N_3752);
nand U3875 (N_3875,N_3791,N_3705);
or U3876 (N_3876,N_3792,N_3782);
nor U3877 (N_3877,N_3795,N_3702);
nor U3878 (N_3878,N_3769,N_3717);
nand U3879 (N_3879,N_3750,N_3790);
nor U3880 (N_3880,N_3797,N_3729);
nor U3881 (N_3881,N_3793,N_3708);
nor U3882 (N_3882,N_3700,N_3768);
nand U3883 (N_3883,N_3713,N_3790);
and U3884 (N_3884,N_3736,N_3721);
nor U3885 (N_3885,N_3704,N_3784);
nand U3886 (N_3886,N_3754,N_3793);
or U3887 (N_3887,N_3761,N_3710);
nand U3888 (N_3888,N_3711,N_3741);
and U3889 (N_3889,N_3787,N_3710);
and U3890 (N_3890,N_3731,N_3772);
nand U3891 (N_3891,N_3772,N_3749);
and U3892 (N_3892,N_3770,N_3707);
or U3893 (N_3893,N_3770,N_3763);
and U3894 (N_3894,N_3734,N_3742);
or U3895 (N_3895,N_3781,N_3703);
nand U3896 (N_3896,N_3797,N_3749);
or U3897 (N_3897,N_3737,N_3752);
and U3898 (N_3898,N_3730,N_3724);
or U3899 (N_3899,N_3797,N_3719);
or U3900 (N_3900,N_3807,N_3806);
nor U3901 (N_3901,N_3883,N_3870);
or U3902 (N_3902,N_3852,N_3829);
or U3903 (N_3903,N_3826,N_3859);
nor U3904 (N_3904,N_3862,N_3853);
nand U3905 (N_3905,N_3864,N_3863);
nor U3906 (N_3906,N_3860,N_3810);
nor U3907 (N_3907,N_3830,N_3805);
nand U3908 (N_3908,N_3816,N_3840);
nor U3909 (N_3909,N_3831,N_3801);
nor U3910 (N_3910,N_3874,N_3868);
nor U3911 (N_3911,N_3812,N_3843);
and U3912 (N_3912,N_3872,N_3848);
nor U3913 (N_3913,N_3893,N_3881);
nor U3914 (N_3914,N_3842,N_3808);
nor U3915 (N_3915,N_3809,N_3824);
nand U3916 (N_3916,N_3819,N_3835);
or U3917 (N_3917,N_3866,N_3895);
nor U3918 (N_3918,N_3856,N_3855);
and U3919 (N_3919,N_3837,N_3833);
and U3920 (N_3920,N_3804,N_3851);
nand U3921 (N_3921,N_3823,N_3890);
nand U3922 (N_3922,N_3877,N_3821);
nor U3923 (N_3923,N_3879,N_3818);
or U3924 (N_3924,N_3839,N_3867);
nand U3925 (N_3925,N_3846,N_3886);
xor U3926 (N_3926,N_3827,N_3894);
and U3927 (N_3927,N_3802,N_3884);
nor U3928 (N_3928,N_3878,N_3876);
or U3929 (N_3929,N_3825,N_3845);
nand U3930 (N_3930,N_3897,N_3813);
or U3931 (N_3931,N_3869,N_3811);
nand U3932 (N_3932,N_3822,N_3880);
or U3933 (N_3933,N_3820,N_3803);
or U3934 (N_3934,N_3844,N_3832);
nor U3935 (N_3935,N_3836,N_3861);
nor U3936 (N_3936,N_3849,N_3815);
nor U3937 (N_3937,N_3873,N_3898);
or U3938 (N_3938,N_3834,N_3857);
nand U3939 (N_3939,N_3896,N_3885);
or U3940 (N_3940,N_3854,N_3850);
or U3941 (N_3941,N_3887,N_3800);
nand U3942 (N_3942,N_3882,N_3891);
or U3943 (N_3943,N_3841,N_3899);
nand U3944 (N_3944,N_3828,N_3814);
nor U3945 (N_3945,N_3888,N_3889);
nand U3946 (N_3946,N_3838,N_3858);
xnor U3947 (N_3947,N_3865,N_3892);
or U3948 (N_3948,N_3847,N_3875);
nand U3949 (N_3949,N_3817,N_3871);
or U3950 (N_3950,N_3863,N_3894);
nand U3951 (N_3951,N_3884,N_3809);
or U3952 (N_3952,N_3889,N_3835);
nor U3953 (N_3953,N_3888,N_3825);
and U3954 (N_3954,N_3899,N_3852);
nand U3955 (N_3955,N_3889,N_3895);
nor U3956 (N_3956,N_3824,N_3837);
or U3957 (N_3957,N_3832,N_3852);
nand U3958 (N_3958,N_3877,N_3896);
nor U3959 (N_3959,N_3813,N_3824);
nor U3960 (N_3960,N_3864,N_3875);
xnor U3961 (N_3961,N_3806,N_3879);
or U3962 (N_3962,N_3871,N_3881);
nand U3963 (N_3963,N_3837,N_3874);
nor U3964 (N_3964,N_3817,N_3883);
or U3965 (N_3965,N_3891,N_3826);
and U3966 (N_3966,N_3897,N_3804);
nor U3967 (N_3967,N_3837,N_3866);
or U3968 (N_3968,N_3823,N_3869);
nor U3969 (N_3969,N_3852,N_3867);
or U3970 (N_3970,N_3828,N_3895);
and U3971 (N_3971,N_3813,N_3891);
xor U3972 (N_3972,N_3852,N_3889);
and U3973 (N_3973,N_3872,N_3811);
nor U3974 (N_3974,N_3831,N_3840);
or U3975 (N_3975,N_3838,N_3863);
and U3976 (N_3976,N_3821,N_3898);
nand U3977 (N_3977,N_3870,N_3806);
nor U3978 (N_3978,N_3831,N_3815);
or U3979 (N_3979,N_3858,N_3859);
nor U3980 (N_3980,N_3833,N_3821);
nor U3981 (N_3981,N_3862,N_3834);
and U3982 (N_3982,N_3839,N_3870);
nor U3983 (N_3983,N_3826,N_3827);
nor U3984 (N_3984,N_3809,N_3882);
or U3985 (N_3985,N_3801,N_3845);
nor U3986 (N_3986,N_3838,N_3862);
nor U3987 (N_3987,N_3823,N_3883);
nor U3988 (N_3988,N_3824,N_3873);
nor U3989 (N_3989,N_3840,N_3856);
nand U3990 (N_3990,N_3873,N_3856);
and U3991 (N_3991,N_3867,N_3885);
or U3992 (N_3992,N_3894,N_3824);
nand U3993 (N_3993,N_3836,N_3838);
or U3994 (N_3994,N_3837,N_3802);
or U3995 (N_3995,N_3842,N_3888);
and U3996 (N_3996,N_3873,N_3852);
and U3997 (N_3997,N_3808,N_3818);
nor U3998 (N_3998,N_3818,N_3850);
nand U3999 (N_3999,N_3821,N_3874);
nor U4000 (N_4000,N_3946,N_3916);
nand U4001 (N_4001,N_3901,N_3943);
or U4002 (N_4002,N_3975,N_3922);
nand U4003 (N_4003,N_3990,N_3981);
nand U4004 (N_4004,N_3920,N_3991);
nor U4005 (N_4005,N_3951,N_3998);
nand U4006 (N_4006,N_3987,N_3928);
xor U4007 (N_4007,N_3953,N_3950);
nand U4008 (N_4008,N_3918,N_3942);
nand U4009 (N_4009,N_3944,N_3908);
nand U4010 (N_4010,N_3911,N_3973);
or U4011 (N_4011,N_3917,N_3939);
nand U4012 (N_4012,N_3978,N_3979);
or U4013 (N_4013,N_3924,N_3933);
or U4014 (N_4014,N_3929,N_3997);
nand U4015 (N_4015,N_3996,N_3915);
and U4016 (N_4016,N_3960,N_3926);
and U4017 (N_4017,N_3954,N_3966);
nand U4018 (N_4018,N_3941,N_3925);
nor U4019 (N_4019,N_3900,N_3972);
and U4020 (N_4020,N_3994,N_3989);
nand U4021 (N_4021,N_3927,N_3965);
and U4022 (N_4022,N_3913,N_3935);
and U4023 (N_4023,N_3938,N_3984);
nor U4024 (N_4024,N_3907,N_3903);
nor U4025 (N_4025,N_3932,N_3985);
and U4026 (N_4026,N_3952,N_3977);
or U4027 (N_4027,N_3963,N_3976);
or U4028 (N_4028,N_3959,N_3919);
and U4029 (N_4029,N_3995,N_3986);
nor U4030 (N_4030,N_3910,N_3962);
nor U4031 (N_4031,N_3923,N_3969);
nor U4032 (N_4032,N_3914,N_3988);
nor U4033 (N_4033,N_3999,N_3930);
nand U4034 (N_4034,N_3980,N_3968);
nor U4035 (N_4035,N_3912,N_3948);
nor U4036 (N_4036,N_3993,N_3909);
or U4037 (N_4037,N_3934,N_3936);
or U4038 (N_4038,N_3964,N_3931);
nor U4039 (N_4039,N_3957,N_3992);
and U4040 (N_4040,N_3906,N_3902);
xnor U4041 (N_4041,N_3905,N_3940);
and U4042 (N_4042,N_3971,N_3945);
nor U4043 (N_4043,N_3921,N_3974);
or U4044 (N_4044,N_3970,N_3983);
or U4045 (N_4045,N_3982,N_3904);
nand U4046 (N_4046,N_3956,N_3958);
nor U4047 (N_4047,N_3955,N_3947);
nor U4048 (N_4048,N_3961,N_3949);
or U4049 (N_4049,N_3937,N_3967);
nand U4050 (N_4050,N_3929,N_3910);
or U4051 (N_4051,N_3941,N_3909);
nor U4052 (N_4052,N_3997,N_3989);
nand U4053 (N_4053,N_3955,N_3985);
or U4054 (N_4054,N_3982,N_3918);
or U4055 (N_4055,N_3913,N_3946);
nor U4056 (N_4056,N_3992,N_3940);
and U4057 (N_4057,N_3921,N_3976);
nor U4058 (N_4058,N_3912,N_3965);
or U4059 (N_4059,N_3972,N_3904);
and U4060 (N_4060,N_3921,N_3905);
and U4061 (N_4061,N_3923,N_3949);
nor U4062 (N_4062,N_3920,N_3958);
nor U4063 (N_4063,N_3985,N_3986);
or U4064 (N_4064,N_3936,N_3908);
or U4065 (N_4065,N_3902,N_3952);
or U4066 (N_4066,N_3972,N_3955);
nor U4067 (N_4067,N_3931,N_3941);
or U4068 (N_4068,N_3957,N_3989);
xnor U4069 (N_4069,N_3997,N_3936);
nor U4070 (N_4070,N_3954,N_3904);
or U4071 (N_4071,N_3924,N_3949);
nand U4072 (N_4072,N_3938,N_3967);
nor U4073 (N_4073,N_3967,N_3961);
nand U4074 (N_4074,N_3949,N_3912);
and U4075 (N_4075,N_3991,N_3981);
nor U4076 (N_4076,N_3924,N_3908);
or U4077 (N_4077,N_3902,N_3997);
and U4078 (N_4078,N_3910,N_3969);
and U4079 (N_4079,N_3935,N_3909);
or U4080 (N_4080,N_3980,N_3941);
nor U4081 (N_4081,N_3924,N_3911);
nor U4082 (N_4082,N_3923,N_3993);
or U4083 (N_4083,N_3971,N_3900);
or U4084 (N_4084,N_3911,N_3932);
nor U4085 (N_4085,N_3922,N_3968);
xor U4086 (N_4086,N_3972,N_3980);
nand U4087 (N_4087,N_3985,N_3965);
nand U4088 (N_4088,N_3915,N_3912);
nand U4089 (N_4089,N_3949,N_3969);
nor U4090 (N_4090,N_3917,N_3962);
and U4091 (N_4091,N_3986,N_3939);
or U4092 (N_4092,N_3991,N_3964);
nor U4093 (N_4093,N_3998,N_3915);
nand U4094 (N_4094,N_3973,N_3986);
nand U4095 (N_4095,N_3916,N_3936);
nand U4096 (N_4096,N_3933,N_3940);
nor U4097 (N_4097,N_3985,N_3915);
or U4098 (N_4098,N_3920,N_3936);
and U4099 (N_4099,N_3948,N_3999);
and U4100 (N_4100,N_4063,N_4076);
nor U4101 (N_4101,N_4079,N_4011);
or U4102 (N_4102,N_4036,N_4095);
nor U4103 (N_4103,N_4078,N_4097);
or U4104 (N_4104,N_4071,N_4058);
and U4105 (N_4105,N_4062,N_4023);
nand U4106 (N_4106,N_4088,N_4042);
or U4107 (N_4107,N_4093,N_4047);
nor U4108 (N_4108,N_4030,N_4094);
or U4109 (N_4109,N_4007,N_4070);
nand U4110 (N_4110,N_4082,N_4085);
nand U4111 (N_4111,N_4067,N_4020);
nor U4112 (N_4112,N_4018,N_4039);
nand U4113 (N_4113,N_4084,N_4053);
or U4114 (N_4114,N_4098,N_4002);
and U4115 (N_4115,N_4035,N_4092);
or U4116 (N_4116,N_4019,N_4081);
nor U4117 (N_4117,N_4048,N_4027);
nor U4118 (N_4118,N_4012,N_4038);
and U4119 (N_4119,N_4046,N_4024);
and U4120 (N_4120,N_4060,N_4000);
and U4121 (N_4121,N_4010,N_4009);
nor U4122 (N_4122,N_4026,N_4069);
nor U4123 (N_4123,N_4074,N_4087);
and U4124 (N_4124,N_4059,N_4031);
nor U4125 (N_4125,N_4003,N_4029);
or U4126 (N_4126,N_4001,N_4080);
nand U4127 (N_4127,N_4025,N_4013);
nand U4128 (N_4128,N_4056,N_4044);
nor U4129 (N_4129,N_4066,N_4054);
nor U4130 (N_4130,N_4086,N_4016);
and U4131 (N_4131,N_4065,N_4057);
and U4132 (N_4132,N_4005,N_4043);
nand U4133 (N_4133,N_4015,N_4061);
nor U4134 (N_4134,N_4089,N_4073);
and U4135 (N_4135,N_4099,N_4041);
nand U4136 (N_4136,N_4055,N_4008);
and U4137 (N_4137,N_4049,N_4033);
or U4138 (N_4138,N_4006,N_4064);
and U4139 (N_4139,N_4052,N_4034);
and U4140 (N_4140,N_4017,N_4014);
and U4141 (N_4141,N_4077,N_4050);
nor U4142 (N_4142,N_4068,N_4091);
nand U4143 (N_4143,N_4072,N_4021);
nand U4144 (N_4144,N_4022,N_4096);
nand U4145 (N_4145,N_4090,N_4051);
nor U4146 (N_4146,N_4040,N_4037);
nor U4147 (N_4147,N_4075,N_4045);
or U4148 (N_4148,N_4028,N_4083);
or U4149 (N_4149,N_4032,N_4004);
or U4150 (N_4150,N_4075,N_4099);
and U4151 (N_4151,N_4095,N_4031);
and U4152 (N_4152,N_4025,N_4021);
nand U4153 (N_4153,N_4025,N_4092);
nand U4154 (N_4154,N_4017,N_4024);
nor U4155 (N_4155,N_4053,N_4070);
nor U4156 (N_4156,N_4049,N_4001);
nor U4157 (N_4157,N_4043,N_4036);
or U4158 (N_4158,N_4068,N_4074);
nor U4159 (N_4159,N_4018,N_4087);
or U4160 (N_4160,N_4074,N_4000);
or U4161 (N_4161,N_4066,N_4045);
nor U4162 (N_4162,N_4005,N_4033);
or U4163 (N_4163,N_4079,N_4087);
nand U4164 (N_4164,N_4043,N_4095);
nor U4165 (N_4165,N_4096,N_4058);
nor U4166 (N_4166,N_4082,N_4051);
nor U4167 (N_4167,N_4017,N_4025);
nand U4168 (N_4168,N_4073,N_4061);
nor U4169 (N_4169,N_4061,N_4077);
nor U4170 (N_4170,N_4025,N_4048);
or U4171 (N_4171,N_4097,N_4022);
nor U4172 (N_4172,N_4072,N_4008);
nand U4173 (N_4173,N_4060,N_4049);
or U4174 (N_4174,N_4001,N_4028);
nand U4175 (N_4175,N_4075,N_4084);
nor U4176 (N_4176,N_4038,N_4020);
nand U4177 (N_4177,N_4095,N_4072);
nand U4178 (N_4178,N_4035,N_4056);
and U4179 (N_4179,N_4029,N_4019);
or U4180 (N_4180,N_4025,N_4044);
or U4181 (N_4181,N_4053,N_4077);
and U4182 (N_4182,N_4050,N_4054);
and U4183 (N_4183,N_4008,N_4024);
nor U4184 (N_4184,N_4041,N_4068);
or U4185 (N_4185,N_4063,N_4044);
nand U4186 (N_4186,N_4082,N_4062);
nor U4187 (N_4187,N_4014,N_4040);
or U4188 (N_4188,N_4018,N_4073);
and U4189 (N_4189,N_4050,N_4017);
or U4190 (N_4190,N_4030,N_4006);
or U4191 (N_4191,N_4053,N_4026);
nor U4192 (N_4192,N_4068,N_4073);
and U4193 (N_4193,N_4076,N_4077);
nor U4194 (N_4194,N_4067,N_4037);
nor U4195 (N_4195,N_4066,N_4026);
or U4196 (N_4196,N_4048,N_4023);
nor U4197 (N_4197,N_4099,N_4044);
or U4198 (N_4198,N_4095,N_4006);
and U4199 (N_4199,N_4049,N_4084);
and U4200 (N_4200,N_4120,N_4114);
nor U4201 (N_4201,N_4180,N_4139);
nor U4202 (N_4202,N_4165,N_4132);
and U4203 (N_4203,N_4174,N_4135);
nor U4204 (N_4204,N_4117,N_4129);
or U4205 (N_4205,N_4103,N_4195);
nand U4206 (N_4206,N_4185,N_4191);
nand U4207 (N_4207,N_4145,N_4107);
and U4208 (N_4208,N_4164,N_4163);
or U4209 (N_4209,N_4196,N_4141);
nand U4210 (N_4210,N_4136,N_4162);
and U4211 (N_4211,N_4170,N_4108);
nand U4212 (N_4212,N_4101,N_4110);
nor U4213 (N_4213,N_4143,N_4118);
nand U4214 (N_4214,N_4125,N_4144);
nor U4215 (N_4215,N_4121,N_4167);
nor U4216 (N_4216,N_4116,N_4154);
nand U4217 (N_4217,N_4173,N_4178);
and U4218 (N_4218,N_4169,N_4193);
nand U4219 (N_4219,N_4183,N_4142);
or U4220 (N_4220,N_4199,N_4155);
or U4221 (N_4221,N_4159,N_4160);
nand U4222 (N_4222,N_4179,N_4190);
nor U4223 (N_4223,N_4157,N_4194);
xnor U4224 (N_4224,N_4152,N_4187);
and U4225 (N_4225,N_4124,N_4112);
or U4226 (N_4226,N_4153,N_4113);
and U4227 (N_4227,N_4133,N_4106);
or U4228 (N_4228,N_4122,N_4188);
and U4229 (N_4229,N_4147,N_4181);
nor U4230 (N_4230,N_4140,N_4128);
nand U4231 (N_4231,N_4161,N_4197);
or U4232 (N_4232,N_4111,N_4176);
nor U4233 (N_4233,N_4115,N_4134);
nor U4234 (N_4234,N_4172,N_4150);
or U4235 (N_4235,N_4104,N_4166);
nand U4236 (N_4236,N_4184,N_4100);
nor U4237 (N_4237,N_4127,N_4158);
nand U4238 (N_4238,N_4131,N_4168);
nand U4239 (N_4239,N_4148,N_4137);
and U4240 (N_4240,N_4189,N_4151);
xor U4241 (N_4241,N_4109,N_4156);
xnor U4242 (N_4242,N_4123,N_4119);
and U4243 (N_4243,N_4102,N_4138);
nand U4244 (N_4244,N_4192,N_4105);
and U4245 (N_4245,N_4126,N_4146);
or U4246 (N_4246,N_4171,N_4175);
or U4247 (N_4247,N_4186,N_4177);
nor U4248 (N_4248,N_4149,N_4198);
nand U4249 (N_4249,N_4182,N_4130);
and U4250 (N_4250,N_4175,N_4129);
and U4251 (N_4251,N_4128,N_4192);
nor U4252 (N_4252,N_4102,N_4174);
nand U4253 (N_4253,N_4189,N_4176);
and U4254 (N_4254,N_4125,N_4103);
and U4255 (N_4255,N_4164,N_4121);
nor U4256 (N_4256,N_4183,N_4128);
nor U4257 (N_4257,N_4108,N_4109);
and U4258 (N_4258,N_4188,N_4125);
nand U4259 (N_4259,N_4177,N_4195);
nand U4260 (N_4260,N_4128,N_4121);
nor U4261 (N_4261,N_4140,N_4141);
nor U4262 (N_4262,N_4135,N_4120);
or U4263 (N_4263,N_4102,N_4103);
nand U4264 (N_4264,N_4123,N_4157);
or U4265 (N_4265,N_4182,N_4163);
or U4266 (N_4266,N_4189,N_4134);
nor U4267 (N_4267,N_4183,N_4109);
nand U4268 (N_4268,N_4123,N_4115);
and U4269 (N_4269,N_4151,N_4198);
and U4270 (N_4270,N_4161,N_4153);
and U4271 (N_4271,N_4134,N_4101);
xnor U4272 (N_4272,N_4162,N_4140);
or U4273 (N_4273,N_4180,N_4152);
xor U4274 (N_4274,N_4179,N_4141);
nor U4275 (N_4275,N_4102,N_4129);
and U4276 (N_4276,N_4131,N_4112);
nand U4277 (N_4277,N_4174,N_4186);
and U4278 (N_4278,N_4172,N_4182);
nor U4279 (N_4279,N_4149,N_4129);
or U4280 (N_4280,N_4184,N_4175);
nor U4281 (N_4281,N_4132,N_4172);
xnor U4282 (N_4282,N_4156,N_4176);
nand U4283 (N_4283,N_4181,N_4190);
or U4284 (N_4284,N_4146,N_4133);
or U4285 (N_4285,N_4104,N_4158);
xor U4286 (N_4286,N_4123,N_4186);
and U4287 (N_4287,N_4189,N_4100);
xor U4288 (N_4288,N_4193,N_4126);
or U4289 (N_4289,N_4159,N_4150);
or U4290 (N_4290,N_4137,N_4147);
and U4291 (N_4291,N_4186,N_4166);
and U4292 (N_4292,N_4105,N_4117);
nor U4293 (N_4293,N_4190,N_4105);
nor U4294 (N_4294,N_4145,N_4117);
and U4295 (N_4295,N_4130,N_4123);
and U4296 (N_4296,N_4105,N_4131);
nand U4297 (N_4297,N_4127,N_4184);
and U4298 (N_4298,N_4151,N_4133);
and U4299 (N_4299,N_4180,N_4128);
or U4300 (N_4300,N_4259,N_4286);
and U4301 (N_4301,N_4205,N_4248);
or U4302 (N_4302,N_4221,N_4284);
or U4303 (N_4303,N_4234,N_4237);
or U4304 (N_4304,N_4223,N_4207);
and U4305 (N_4305,N_4203,N_4268);
nor U4306 (N_4306,N_4204,N_4288);
nand U4307 (N_4307,N_4231,N_4241);
nand U4308 (N_4308,N_4295,N_4230);
or U4309 (N_4309,N_4272,N_4242);
and U4310 (N_4310,N_4264,N_4219);
nor U4311 (N_4311,N_4252,N_4208);
and U4312 (N_4312,N_4249,N_4227);
and U4313 (N_4313,N_4271,N_4293);
and U4314 (N_4314,N_4246,N_4258);
nand U4315 (N_4315,N_4222,N_4245);
or U4316 (N_4316,N_4253,N_4228);
and U4317 (N_4317,N_4263,N_4250);
or U4318 (N_4318,N_4298,N_4282);
nor U4319 (N_4319,N_4266,N_4233);
nor U4320 (N_4320,N_4239,N_4218);
nor U4321 (N_4321,N_4201,N_4238);
and U4322 (N_4322,N_4278,N_4275);
nand U4323 (N_4323,N_4251,N_4274);
nand U4324 (N_4324,N_4206,N_4285);
nor U4325 (N_4325,N_4214,N_4279);
and U4326 (N_4326,N_4247,N_4297);
nand U4327 (N_4327,N_4273,N_4290);
nor U4328 (N_4328,N_4236,N_4225);
xor U4329 (N_4329,N_4232,N_4210);
nand U4330 (N_4330,N_4296,N_4289);
nor U4331 (N_4331,N_4209,N_4240);
and U4332 (N_4332,N_4226,N_4260);
nor U4333 (N_4333,N_4292,N_4235);
nor U4334 (N_4334,N_4287,N_4262);
and U4335 (N_4335,N_4212,N_4265);
nor U4336 (N_4336,N_4256,N_4254);
and U4337 (N_4337,N_4217,N_4255);
nor U4338 (N_4338,N_4244,N_4283);
nor U4339 (N_4339,N_4243,N_4229);
or U4340 (N_4340,N_4299,N_4270);
and U4341 (N_4341,N_4280,N_4267);
or U4342 (N_4342,N_4281,N_4291);
nor U4343 (N_4343,N_4220,N_4276);
nand U4344 (N_4344,N_4213,N_4224);
and U4345 (N_4345,N_4269,N_4202);
xnor U4346 (N_4346,N_4294,N_4211);
or U4347 (N_4347,N_4261,N_4215);
or U4348 (N_4348,N_4216,N_4200);
or U4349 (N_4349,N_4257,N_4277);
and U4350 (N_4350,N_4211,N_4277);
nor U4351 (N_4351,N_4239,N_4224);
or U4352 (N_4352,N_4205,N_4256);
nand U4353 (N_4353,N_4264,N_4276);
and U4354 (N_4354,N_4205,N_4269);
or U4355 (N_4355,N_4236,N_4231);
or U4356 (N_4356,N_4299,N_4202);
and U4357 (N_4357,N_4262,N_4258);
nand U4358 (N_4358,N_4264,N_4240);
or U4359 (N_4359,N_4217,N_4263);
and U4360 (N_4360,N_4273,N_4231);
or U4361 (N_4361,N_4244,N_4261);
nor U4362 (N_4362,N_4278,N_4258);
nand U4363 (N_4363,N_4218,N_4266);
nand U4364 (N_4364,N_4241,N_4273);
and U4365 (N_4365,N_4207,N_4297);
or U4366 (N_4366,N_4280,N_4269);
or U4367 (N_4367,N_4241,N_4227);
nand U4368 (N_4368,N_4261,N_4235);
and U4369 (N_4369,N_4262,N_4227);
nor U4370 (N_4370,N_4219,N_4271);
and U4371 (N_4371,N_4233,N_4200);
nor U4372 (N_4372,N_4216,N_4220);
nand U4373 (N_4373,N_4267,N_4214);
xnor U4374 (N_4374,N_4251,N_4293);
nand U4375 (N_4375,N_4258,N_4203);
nor U4376 (N_4376,N_4232,N_4205);
and U4377 (N_4377,N_4277,N_4210);
nor U4378 (N_4378,N_4217,N_4221);
and U4379 (N_4379,N_4284,N_4203);
nand U4380 (N_4380,N_4259,N_4221);
and U4381 (N_4381,N_4294,N_4203);
nor U4382 (N_4382,N_4245,N_4289);
nand U4383 (N_4383,N_4294,N_4252);
nand U4384 (N_4384,N_4292,N_4290);
nor U4385 (N_4385,N_4287,N_4209);
nor U4386 (N_4386,N_4214,N_4266);
nor U4387 (N_4387,N_4245,N_4299);
nand U4388 (N_4388,N_4212,N_4214);
and U4389 (N_4389,N_4223,N_4258);
and U4390 (N_4390,N_4277,N_4222);
nor U4391 (N_4391,N_4277,N_4206);
nand U4392 (N_4392,N_4272,N_4273);
and U4393 (N_4393,N_4291,N_4234);
nand U4394 (N_4394,N_4288,N_4289);
or U4395 (N_4395,N_4288,N_4228);
nor U4396 (N_4396,N_4202,N_4251);
or U4397 (N_4397,N_4208,N_4292);
xnor U4398 (N_4398,N_4295,N_4244);
xnor U4399 (N_4399,N_4239,N_4265);
nor U4400 (N_4400,N_4347,N_4369);
xnor U4401 (N_4401,N_4362,N_4381);
or U4402 (N_4402,N_4331,N_4388);
xnor U4403 (N_4403,N_4380,N_4336);
and U4404 (N_4404,N_4389,N_4335);
or U4405 (N_4405,N_4393,N_4313);
nor U4406 (N_4406,N_4329,N_4361);
nand U4407 (N_4407,N_4317,N_4303);
or U4408 (N_4408,N_4376,N_4333);
xor U4409 (N_4409,N_4364,N_4324);
or U4410 (N_4410,N_4308,N_4343);
or U4411 (N_4411,N_4326,N_4372);
and U4412 (N_4412,N_4345,N_4391);
nand U4413 (N_4413,N_4398,N_4390);
or U4414 (N_4414,N_4358,N_4310);
or U4415 (N_4415,N_4371,N_4378);
nor U4416 (N_4416,N_4344,N_4319);
and U4417 (N_4417,N_4307,N_4366);
nor U4418 (N_4418,N_4340,N_4332);
or U4419 (N_4419,N_4305,N_4351);
nor U4420 (N_4420,N_4387,N_4382);
or U4421 (N_4421,N_4383,N_4367);
and U4422 (N_4422,N_4322,N_4373);
or U4423 (N_4423,N_4346,N_4323);
nor U4424 (N_4424,N_4301,N_4396);
and U4425 (N_4425,N_4370,N_4363);
nor U4426 (N_4426,N_4309,N_4360);
or U4427 (N_4427,N_4315,N_4385);
and U4428 (N_4428,N_4316,N_4328);
nor U4429 (N_4429,N_4392,N_4395);
nand U4430 (N_4430,N_4374,N_4327);
nor U4431 (N_4431,N_4334,N_4330);
or U4432 (N_4432,N_4356,N_4312);
and U4433 (N_4433,N_4379,N_4314);
nand U4434 (N_4434,N_4338,N_4342);
or U4435 (N_4435,N_4320,N_4384);
or U4436 (N_4436,N_4357,N_4397);
nand U4437 (N_4437,N_4311,N_4321);
nand U4438 (N_4438,N_4352,N_4350);
or U4439 (N_4439,N_4304,N_4365);
nor U4440 (N_4440,N_4337,N_4302);
and U4441 (N_4441,N_4377,N_4353);
nand U4442 (N_4442,N_4300,N_4341);
nor U4443 (N_4443,N_4375,N_4368);
and U4444 (N_4444,N_4349,N_4386);
or U4445 (N_4445,N_4394,N_4318);
or U4446 (N_4446,N_4339,N_4354);
or U4447 (N_4447,N_4325,N_4355);
or U4448 (N_4448,N_4306,N_4348);
nand U4449 (N_4449,N_4399,N_4359);
nand U4450 (N_4450,N_4378,N_4383);
and U4451 (N_4451,N_4338,N_4308);
nor U4452 (N_4452,N_4343,N_4342);
nand U4453 (N_4453,N_4375,N_4369);
nor U4454 (N_4454,N_4394,N_4380);
nand U4455 (N_4455,N_4320,N_4376);
nand U4456 (N_4456,N_4371,N_4350);
and U4457 (N_4457,N_4354,N_4302);
nand U4458 (N_4458,N_4378,N_4358);
and U4459 (N_4459,N_4318,N_4374);
and U4460 (N_4460,N_4358,N_4319);
and U4461 (N_4461,N_4358,N_4395);
nor U4462 (N_4462,N_4378,N_4317);
nor U4463 (N_4463,N_4374,N_4376);
nor U4464 (N_4464,N_4384,N_4343);
nor U4465 (N_4465,N_4368,N_4367);
nor U4466 (N_4466,N_4370,N_4329);
or U4467 (N_4467,N_4394,N_4383);
nor U4468 (N_4468,N_4324,N_4366);
nor U4469 (N_4469,N_4337,N_4309);
or U4470 (N_4470,N_4397,N_4347);
or U4471 (N_4471,N_4317,N_4321);
nor U4472 (N_4472,N_4329,N_4319);
nor U4473 (N_4473,N_4363,N_4353);
nor U4474 (N_4474,N_4336,N_4385);
nand U4475 (N_4475,N_4360,N_4383);
nand U4476 (N_4476,N_4378,N_4345);
or U4477 (N_4477,N_4368,N_4328);
and U4478 (N_4478,N_4308,N_4345);
and U4479 (N_4479,N_4311,N_4396);
nand U4480 (N_4480,N_4349,N_4355);
xor U4481 (N_4481,N_4380,N_4357);
xor U4482 (N_4482,N_4353,N_4351);
nor U4483 (N_4483,N_4326,N_4321);
nor U4484 (N_4484,N_4382,N_4374);
and U4485 (N_4485,N_4386,N_4395);
nand U4486 (N_4486,N_4315,N_4352);
and U4487 (N_4487,N_4304,N_4331);
or U4488 (N_4488,N_4383,N_4371);
nor U4489 (N_4489,N_4324,N_4307);
nor U4490 (N_4490,N_4370,N_4352);
nand U4491 (N_4491,N_4316,N_4394);
nand U4492 (N_4492,N_4376,N_4357);
and U4493 (N_4493,N_4394,N_4354);
and U4494 (N_4494,N_4328,N_4321);
nor U4495 (N_4495,N_4384,N_4365);
nand U4496 (N_4496,N_4373,N_4366);
nand U4497 (N_4497,N_4334,N_4354);
nor U4498 (N_4498,N_4369,N_4313);
or U4499 (N_4499,N_4354,N_4337);
and U4500 (N_4500,N_4404,N_4452);
and U4501 (N_4501,N_4488,N_4413);
or U4502 (N_4502,N_4497,N_4463);
or U4503 (N_4503,N_4468,N_4480);
and U4504 (N_4504,N_4430,N_4442);
nand U4505 (N_4505,N_4475,N_4420);
nand U4506 (N_4506,N_4427,N_4426);
and U4507 (N_4507,N_4472,N_4464);
and U4508 (N_4508,N_4402,N_4489);
nand U4509 (N_4509,N_4437,N_4492);
or U4510 (N_4510,N_4428,N_4462);
nand U4511 (N_4511,N_4458,N_4481);
or U4512 (N_4512,N_4499,N_4438);
nand U4513 (N_4513,N_4453,N_4439);
and U4514 (N_4514,N_4403,N_4471);
xnor U4515 (N_4515,N_4423,N_4401);
nor U4516 (N_4516,N_4498,N_4478);
or U4517 (N_4517,N_4432,N_4417);
and U4518 (N_4518,N_4474,N_4418);
nor U4519 (N_4519,N_4440,N_4409);
or U4520 (N_4520,N_4429,N_4450);
and U4521 (N_4521,N_4479,N_4467);
nor U4522 (N_4522,N_4460,N_4448);
and U4523 (N_4523,N_4411,N_4425);
nand U4524 (N_4524,N_4424,N_4491);
nand U4525 (N_4525,N_4459,N_4444);
nor U4526 (N_4526,N_4451,N_4414);
or U4527 (N_4527,N_4457,N_4434);
nor U4528 (N_4528,N_4476,N_4449);
or U4529 (N_4529,N_4456,N_4484);
or U4530 (N_4530,N_4455,N_4405);
nor U4531 (N_4531,N_4461,N_4407);
or U4532 (N_4532,N_4493,N_4495);
nor U4533 (N_4533,N_4415,N_4441);
nand U4534 (N_4534,N_4485,N_4422);
and U4535 (N_4535,N_4469,N_4416);
or U4536 (N_4536,N_4465,N_4431);
nand U4537 (N_4537,N_4410,N_4482);
and U4538 (N_4538,N_4412,N_4483);
and U4539 (N_4539,N_4490,N_4447);
nand U4540 (N_4540,N_4445,N_4436);
or U4541 (N_4541,N_4406,N_4408);
nor U4542 (N_4542,N_4419,N_4443);
nor U4543 (N_4543,N_4433,N_4400);
nand U4544 (N_4544,N_4435,N_4477);
or U4545 (N_4545,N_4446,N_4487);
nor U4546 (N_4546,N_4486,N_4473);
nand U4547 (N_4547,N_4454,N_4470);
and U4548 (N_4548,N_4496,N_4466);
nand U4549 (N_4549,N_4494,N_4421);
nor U4550 (N_4550,N_4424,N_4461);
nand U4551 (N_4551,N_4400,N_4495);
and U4552 (N_4552,N_4468,N_4410);
nand U4553 (N_4553,N_4464,N_4405);
nor U4554 (N_4554,N_4417,N_4473);
or U4555 (N_4555,N_4474,N_4492);
and U4556 (N_4556,N_4400,N_4476);
nor U4557 (N_4557,N_4448,N_4456);
nand U4558 (N_4558,N_4435,N_4407);
nor U4559 (N_4559,N_4402,N_4418);
and U4560 (N_4560,N_4464,N_4483);
nor U4561 (N_4561,N_4440,N_4422);
xor U4562 (N_4562,N_4472,N_4461);
nor U4563 (N_4563,N_4456,N_4445);
nand U4564 (N_4564,N_4463,N_4472);
nand U4565 (N_4565,N_4478,N_4434);
and U4566 (N_4566,N_4477,N_4484);
xor U4567 (N_4567,N_4419,N_4465);
nor U4568 (N_4568,N_4494,N_4467);
or U4569 (N_4569,N_4499,N_4489);
nand U4570 (N_4570,N_4425,N_4459);
nor U4571 (N_4571,N_4443,N_4432);
nand U4572 (N_4572,N_4442,N_4423);
nor U4573 (N_4573,N_4405,N_4432);
or U4574 (N_4574,N_4489,N_4429);
and U4575 (N_4575,N_4441,N_4472);
and U4576 (N_4576,N_4421,N_4482);
and U4577 (N_4577,N_4404,N_4408);
xnor U4578 (N_4578,N_4435,N_4425);
nand U4579 (N_4579,N_4487,N_4420);
and U4580 (N_4580,N_4427,N_4458);
and U4581 (N_4581,N_4451,N_4457);
and U4582 (N_4582,N_4471,N_4401);
or U4583 (N_4583,N_4484,N_4472);
nand U4584 (N_4584,N_4485,N_4420);
or U4585 (N_4585,N_4484,N_4411);
and U4586 (N_4586,N_4409,N_4457);
or U4587 (N_4587,N_4436,N_4412);
or U4588 (N_4588,N_4420,N_4456);
and U4589 (N_4589,N_4403,N_4476);
or U4590 (N_4590,N_4453,N_4426);
or U4591 (N_4591,N_4434,N_4479);
and U4592 (N_4592,N_4410,N_4458);
and U4593 (N_4593,N_4424,N_4417);
or U4594 (N_4594,N_4447,N_4492);
and U4595 (N_4595,N_4470,N_4474);
and U4596 (N_4596,N_4493,N_4488);
nor U4597 (N_4597,N_4406,N_4492);
and U4598 (N_4598,N_4483,N_4478);
xnor U4599 (N_4599,N_4435,N_4409);
or U4600 (N_4600,N_4510,N_4552);
nand U4601 (N_4601,N_4554,N_4542);
and U4602 (N_4602,N_4505,N_4543);
or U4603 (N_4603,N_4539,N_4567);
and U4604 (N_4604,N_4514,N_4516);
and U4605 (N_4605,N_4531,N_4578);
or U4606 (N_4606,N_4507,N_4597);
or U4607 (N_4607,N_4544,N_4557);
nor U4608 (N_4608,N_4534,N_4559);
or U4609 (N_4609,N_4560,N_4571);
and U4610 (N_4610,N_4537,N_4535);
or U4611 (N_4611,N_4529,N_4593);
or U4612 (N_4612,N_4532,N_4547);
or U4613 (N_4613,N_4503,N_4591);
nand U4614 (N_4614,N_4568,N_4595);
nand U4615 (N_4615,N_4588,N_4540);
and U4616 (N_4616,N_4582,N_4580);
and U4617 (N_4617,N_4563,N_4570);
nand U4618 (N_4618,N_4584,N_4528);
xnor U4619 (N_4619,N_4576,N_4587);
nand U4620 (N_4620,N_4521,N_4579);
and U4621 (N_4621,N_4558,N_4596);
or U4622 (N_4622,N_4565,N_4577);
and U4623 (N_4623,N_4530,N_4574);
or U4624 (N_4624,N_4517,N_4511);
or U4625 (N_4625,N_4590,N_4501);
nor U4626 (N_4626,N_4562,N_4555);
nor U4627 (N_4627,N_4551,N_4541);
or U4628 (N_4628,N_4500,N_4548);
and U4629 (N_4629,N_4556,N_4564);
or U4630 (N_4630,N_4524,N_4575);
or U4631 (N_4631,N_4589,N_4550);
or U4632 (N_4632,N_4598,N_4520);
or U4633 (N_4633,N_4549,N_4509);
and U4634 (N_4634,N_4599,N_4527);
nor U4635 (N_4635,N_4586,N_4523);
nand U4636 (N_4636,N_4519,N_4506);
nand U4637 (N_4637,N_4594,N_4504);
nand U4638 (N_4638,N_4512,N_4515);
or U4639 (N_4639,N_4566,N_4522);
nand U4640 (N_4640,N_4585,N_4572);
or U4641 (N_4641,N_4533,N_4553);
nor U4642 (N_4642,N_4573,N_4561);
and U4643 (N_4643,N_4513,N_4502);
and U4644 (N_4644,N_4518,N_4525);
nand U4645 (N_4645,N_4508,N_4545);
or U4646 (N_4646,N_4538,N_4569);
and U4647 (N_4647,N_4536,N_4592);
xor U4648 (N_4648,N_4583,N_4546);
nor U4649 (N_4649,N_4526,N_4581);
nand U4650 (N_4650,N_4500,N_4585);
or U4651 (N_4651,N_4581,N_4523);
and U4652 (N_4652,N_4552,N_4566);
or U4653 (N_4653,N_4568,N_4585);
nor U4654 (N_4654,N_4537,N_4578);
and U4655 (N_4655,N_4506,N_4526);
nor U4656 (N_4656,N_4514,N_4535);
xor U4657 (N_4657,N_4503,N_4570);
or U4658 (N_4658,N_4508,N_4595);
or U4659 (N_4659,N_4574,N_4566);
nor U4660 (N_4660,N_4500,N_4517);
nand U4661 (N_4661,N_4510,N_4501);
nand U4662 (N_4662,N_4581,N_4569);
and U4663 (N_4663,N_4535,N_4548);
nand U4664 (N_4664,N_4561,N_4544);
nand U4665 (N_4665,N_4591,N_4564);
nor U4666 (N_4666,N_4538,N_4587);
or U4667 (N_4667,N_4538,N_4554);
and U4668 (N_4668,N_4514,N_4508);
and U4669 (N_4669,N_4557,N_4596);
or U4670 (N_4670,N_4502,N_4574);
nor U4671 (N_4671,N_4566,N_4539);
or U4672 (N_4672,N_4552,N_4567);
nor U4673 (N_4673,N_4514,N_4580);
nand U4674 (N_4674,N_4544,N_4579);
or U4675 (N_4675,N_4538,N_4510);
nand U4676 (N_4676,N_4527,N_4557);
and U4677 (N_4677,N_4538,N_4512);
or U4678 (N_4678,N_4564,N_4555);
nand U4679 (N_4679,N_4558,N_4578);
nand U4680 (N_4680,N_4590,N_4500);
nor U4681 (N_4681,N_4520,N_4534);
and U4682 (N_4682,N_4519,N_4588);
or U4683 (N_4683,N_4502,N_4541);
nor U4684 (N_4684,N_4516,N_4521);
nor U4685 (N_4685,N_4506,N_4537);
nand U4686 (N_4686,N_4572,N_4520);
nor U4687 (N_4687,N_4527,N_4568);
and U4688 (N_4688,N_4560,N_4500);
and U4689 (N_4689,N_4593,N_4575);
nand U4690 (N_4690,N_4590,N_4593);
and U4691 (N_4691,N_4547,N_4548);
or U4692 (N_4692,N_4583,N_4564);
or U4693 (N_4693,N_4566,N_4596);
nand U4694 (N_4694,N_4554,N_4567);
nand U4695 (N_4695,N_4560,N_4592);
nand U4696 (N_4696,N_4584,N_4560);
or U4697 (N_4697,N_4578,N_4597);
nand U4698 (N_4698,N_4537,N_4595);
nand U4699 (N_4699,N_4514,N_4549);
nand U4700 (N_4700,N_4692,N_4621);
and U4701 (N_4701,N_4608,N_4620);
nand U4702 (N_4702,N_4627,N_4651);
xor U4703 (N_4703,N_4618,N_4677);
nand U4704 (N_4704,N_4676,N_4614);
and U4705 (N_4705,N_4639,N_4673);
or U4706 (N_4706,N_4669,N_4600);
nor U4707 (N_4707,N_4632,N_4693);
nand U4708 (N_4708,N_4668,N_4654);
and U4709 (N_4709,N_4666,N_4671);
xor U4710 (N_4710,N_4605,N_4682);
nor U4711 (N_4711,N_4635,N_4606);
or U4712 (N_4712,N_4603,N_4672);
nand U4713 (N_4713,N_4681,N_4643);
nand U4714 (N_4714,N_4616,N_4661);
or U4715 (N_4715,N_4619,N_4629);
nor U4716 (N_4716,N_4644,N_4656);
nor U4717 (N_4717,N_4684,N_4630);
nand U4718 (N_4718,N_4645,N_4689);
or U4719 (N_4719,N_4653,N_4691);
and U4720 (N_4720,N_4695,N_4663);
nor U4721 (N_4721,N_4607,N_4665);
nand U4722 (N_4722,N_4655,N_4680);
and U4723 (N_4723,N_4660,N_4612);
nor U4724 (N_4724,N_4688,N_4658);
or U4725 (N_4725,N_4610,N_4694);
nand U4726 (N_4726,N_4641,N_4687);
nor U4727 (N_4727,N_4678,N_4623);
and U4728 (N_4728,N_4613,N_4690);
xnor U4729 (N_4729,N_4631,N_4657);
or U4730 (N_4730,N_4647,N_4675);
and U4731 (N_4731,N_4662,N_4622);
or U4732 (N_4732,N_4637,N_4696);
nand U4733 (N_4733,N_4624,N_4633);
nand U4734 (N_4734,N_4626,N_4650);
nand U4735 (N_4735,N_4667,N_4636);
nand U4736 (N_4736,N_4615,N_4611);
nand U4737 (N_4737,N_4697,N_4617);
xor U4738 (N_4738,N_4634,N_4648);
nor U4739 (N_4739,N_4646,N_4679);
and U4740 (N_4740,N_4628,N_4670);
and U4741 (N_4741,N_4664,N_4642);
or U4742 (N_4742,N_4698,N_4625);
and U4743 (N_4743,N_4674,N_4640);
nand U4744 (N_4744,N_4609,N_4659);
nor U4745 (N_4745,N_4685,N_4601);
nand U4746 (N_4746,N_4683,N_4699);
and U4747 (N_4747,N_4649,N_4604);
nor U4748 (N_4748,N_4602,N_4652);
and U4749 (N_4749,N_4686,N_4638);
and U4750 (N_4750,N_4644,N_4628);
xnor U4751 (N_4751,N_4604,N_4641);
and U4752 (N_4752,N_4681,N_4651);
and U4753 (N_4753,N_4607,N_4658);
or U4754 (N_4754,N_4674,N_4697);
or U4755 (N_4755,N_4608,N_4613);
or U4756 (N_4756,N_4645,N_4619);
and U4757 (N_4757,N_4600,N_4698);
or U4758 (N_4758,N_4605,N_4629);
nor U4759 (N_4759,N_4678,N_4637);
and U4760 (N_4760,N_4601,N_4639);
and U4761 (N_4761,N_4646,N_4662);
nand U4762 (N_4762,N_4661,N_4697);
and U4763 (N_4763,N_4672,N_4610);
nor U4764 (N_4764,N_4608,N_4614);
or U4765 (N_4765,N_4692,N_4629);
nand U4766 (N_4766,N_4692,N_4649);
and U4767 (N_4767,N_4693,N_4657);
or U4768 (N_4768,N_4640,N_4690);
nand U4769 (N_4769,N_4617,N_4634);
or U4770 (N_4770,N_4623,N_4643);
nand U4771 (N_4771,N_4680,N_4681);
and U4772 (N_4772,N_4615,N_4601);
nor U4773 (N_4773,N_4610,N_4656);
and U4774 (N_4774,N_4613,N_4603);
nand U4775 (N_4775,N_4600,N_4611);
and U4776 (N_4776,N_4679,N_4655);
or U4777 (N_4777,N_4641,N_4647);
nor U4778 (N_4778,N_4660,N_4641);
nand U4779 (N_4779,N_4623,N_4690);
and U4780 (N_4780,N_4673,N_4616);
and U4781 (N_4781,N_4640,N_4693);
nor U4782 (N_4782,N_4606,N_4613);
or U4783 (N_4783,N_4618,N_4662);
nor U4784 (N_4784,N_4609,N_4627);
nor U4785 (N_4785,N_4648,N_4606);
and U4786 (N_4786,N_4612,N_4676);
nand U4787 (N_4787,N_4631,N_4686);
nand U4788 (N_4788,N_4636,N_4670);
xnor U4789 (N_4789,N_4620,N_4676);
nor U4790 (N_4790,N_4673,N_4629);
and U4791 (N_4791,N_4606,N_4631);
nand U4792 (N_4792,N_4610,N_4692);
or U4793 (N_4793,N_4624,N_4662);
or U4794 (N_4794,N_4698,N_4658);
nand U4795 (N_4795,N_4695,N_4682);
and U4796 (N_4796,N_4659,N_4622);
or U4797 (N_4797,N_4643,N_4640);
nand U4798 (N_4798,N_4694,N_4615);
and U4799 (N_4799,N_4601,N_4691);
nor U4800 (N_4800,N_4705,N_4749);
and U4801 (N_4801,N_4723,N_4789);
and U4802 (N_4802,N_4707,N_4704);
xor U4803 (N_4803,N_4791,N_4725);
nand U4804 (N_4804,N_4708,N_4790);
or U4805 (N_4805,N_4719,N_4779);
nor U4806 (N_4806,N_4793,N_4729);
nand U4807 (N_4807,N_4737,N_4766);
nor U4808 (N_4808,N_4746,N_4754);
nor U4809 (N_4809,N_4787,N_4764);
nand U4810 (N_4810,N_4717,N_4777);
and U4811 (N_4811,N_4752,N_4714);
or U4812 (N_4812,N_4785,N_4773);
or U4813 (N_4813,N_4736,N_4711);
and U4814 (N_4814,N_4731,N_4796);
nor U4815 (N_4815,N_4722,N_4776);
and U4816 (N_4816,N_4733,N_4772);
or U4817 (N_4817,N_4724,N_4727);
nor U4818 (N_4818,N_4716,N_4763);
or U4819 (N_4819,N_4732,N_4703);
nand U4820 (N_4820,N_4758,N_4799);
and U4821 (N_4821,N_4784,N_4743);
or U4822 (N_4822,N_4715,N_4726);
or U4823 (N_4823,N_4751,N_4797);
nand U4824 (N_4824,N_4788,N_4794);
and U4825 (N_4825,N_4701,N_4783);
and U4826 (N_4826,N_4769,N_4710);
and U4827 (N_4827,N_4742,N_4780);
and U4828 (N_4828,N_4760,N_4795);
and U4829 (N_4829,N_4712,N_4798);
and U4830 (N_4830,N_4745,N_4753);
and U4831 (N_4831,N_4768,N_4767);
xor U4832 (N_4832,N_4755,N_4792);
nor U4833 (N_4833,N_4774,N_4735);
nor U4834 (N_4834,N_4747,N_4759);
nand U4835 (N_4835,N_4782,N_4718);
or U4836 (N_4836,N_4770,N_4786);
nand U4837 (N_4837,N_4702,N_4744);
and U4838 (N_4838,N_4709,N_4700);
and U4839 (N_4839,N_4775,N_4756);
and U4840 (N_4840,N_4721,N_4738);
and U4841 (N_4841,N_4739,N_4778);
and U4842 (N_4842,N_4762,N_4750);
nand U4843 (N_4843,N_4734,N_4765);
or U4844 (N_4844,N_4706,N_4741);
nor U4845 (N_4845,N_4728,N_4720);
or U4846 (N_4846,N_4761,N_4771);
nand U4847 (N_4847,N_4748,N_4713);
and U4848 (N_4848,N_4757,N_4730);
nor U4849 (N_4849,N_4740,N_4781);
nor U4850 (N_4850,N_4724,N_4712);
or U4851 (N_4851,N_4730,N_4736);
nor U4852 (N_4852,N_4749,N_4730);
and U4853 (N_4853,N_4788,N_4712);
and U4854 (N_4854,N_4739,N_4737);
or U4855 (N_4855,N_4764,N_4730);
nor U4856 (N_4856,N_4751,N_4736);
nand U4857 (N_4857,N_4716,N_4735);
and U4858 (N_4858,N_4788,N_4731);
and U4859 (N_4859,N_4709,N_4772);
or U4860 (N_4860,N_4724,N_4749);
and U4861 (N_4861,N_4789,N_4796);
and U4862 (N_4862,N_4709,N_4762);
and U4863 (N_4863,N_4765,N_4778);
nand U4864 (N_4864,N_4791,N_4753);
nor U4865 (N_4865,N_4769,N_4775);
and U4866 (N_4866,N_4700,N_4742);
or U4867 (N_4867,N_4797,N_4793);
or U4868 (N_4868,N_4799,N_4794);
or U4869 (N_4869,N_4722,N_4751);
or U4870 (N_4870,N_4751,N_4725);
nand U4871 (N_4871,N_4761,N_4701);
nand U4872 (N_4872,N_4723,N_4786);
nor U4873 (N_4873,N_4779,N_4799);
and U4874 (N_4874,N_4754,N_4769);
nor U4875 (N_4875,N_4748,N_4712);
nor U4876 (N_4876,N_4727,N_4790);
and U4877 (N_4877,N_4769,N_4782);
nand U4878 (N_4878,N_4747,N_4760);
or U4879 (N_4879,N_4729,N_4769);
xnor U4880 (N_4880,N_4748,N_4786);
or U4881 (N_4881,N_4726,N_4783);
nor U4882 (N_4882,N_4765,N_4768);
or U4883 (N_4883,N_4795,N_4790);
xnor U4884 (N_4884,N_4707,N_4786);
nand U4885 (N_4885,N_4710,N_4751);
nand U4886 (N_4886,N_4702,N_4709);
nor U4887 (N_4887,N_4787,N_4768);
or U4888 (N_4888,N_4785,N_4722);
and U4889 (N_4889,N_4751,N_4794);
or U4890 (N_4890,N_4764,N_4755);
nor U4891 (N_4891,N_4733,N_4706);
or U4892 (N_4892,N_4786,N_4795);
nor U4893 (N_4893,N_4789,N_4795);
and U4894 (N_4894,N_4777,N_4716);
or U4895 (N_4895,N_4718,N_4750);
and U4896 (N_4896,N_4735,N_4793);
or U4897 (N_4897,N_4728,N_4783);
nor U4898 (N_4898,N_4719,N_4725);
nor U4899 (N_4899,N_4740,N_4731);
and U4900 (N_4900,N_4837,N_4852);
and U4901 (N_4901,N_4834,N_4872);
nand U4902 (N_4902,N_4862,N_4889);
nand U4903 (N_4903,N_4861,N_4808);
nor U4904 (N_4904,N_4870,N_4836);
nand U4905 (N_4905,N_4880,N_4894);
and U4906 (N_4906,N_4863,N_4801);
nor U4907 (N_4907,N_4841,N_4840);
nor U4908 (N_4908,N_4887,N_4812);
nand U4909 (N_4909,N_4856,N_4886);
nand U4910 (N_4910,N_4855,N_4883);
nor U4911 (N_4911,N_4811,N_4857);
and U4912 (N_4912,N_4888,N_4893);
nor U4913 (N_4913,N_4802,N_4867);
or U4914 (N_4914,N_4831,N_4830);
nor U4915 (N_4915,N_4869,N_4897);
or U4916 (N_4916,N_4821,N_4824);
nand U4917 (N_4917,N_4876,N_4810);
or U4918 (N_4918,N_4844,N_4819);
or U4919 (N_4919,N_4890,N_4875);
nand U4920 (N_4920,N_4820,N_4842);
nor U4921 (N_4921,N_4832,N_4829);
and U4922 (N_4922,N_4828,N_4881);
or U4923 (N_4923,N_4892,N_4823);
or U4924 (N_4924,N_4846,N_4859);
or U4925 (N_4925,N_4848,N_4898);
and U4926 (N_4926,N_4845,N_4874);
nand U4927 (N_4927,N_4827,N_4866);
nor U4928 (N_4928,N_4864,N_4813);
and U4929 (N_4929,N_4838,N_4835);
nand U4930 (N_4930,N_4851,N_4882);
and U4931 (N_4931,N_4826,N_4809);
and U4932 (N_4932,N_4873,N_4816);
and U4933 (N_4933,N_4896,N_4879);
and U4934 (N_4934,N_4868,N_4860);
nand U4935 (N_4935,N_4884,N_4817);
and U4936 (N_4936,N_4858,N_4899);
xnor U4937 (N_4937,N_4833,N_4843);
or U4938 (N_4938,N_4885,N_4877);
nand U4939 (N_4939,N_4850,N_4822);
or U4940 (N_4940,N_4805,N_4839);
nand U4941 (N_4941,N_4818,N_4871);
nand U4942 (N_4942,N_4849,N_4815);
and U4943 (N_4943,N_4891,N_4800);
and U4944 (N_4944,N_4854,N_4804);
or U4945 (N_4945,N_4878,N_4895);
or U4946 (N_4946,N_4847,N_4825);
nor U4947 (N_4947,N_4803,N_4853);
nand U4948 (N_4948,N_4814,N_4806);
nand U4949 (N_4949,N_4865,N_4807);
nor U4950 (N_4950,N_4847,N_4840);
or U4951 (N_4951,N_4898,N_4839);
or U4952 (N_4952,N_4885,N_4814);
nand U4953 (N_4953,N_4810,N_4829);
and U4954 (N_4954,N_4872,N_4873);
nor U4955 (N_4955,N_4837,N_4847);
or U4956 (N_4956,N_4806,N_4826);
or U4957 (N_4957,N_4857,N_4869);
or U4958 (N_4958,N_4877,N_4865);
and U4959 (N_4959,N_4801,N_4854);
nor U4960 (N_4960,N_4888,N_4862);
or U4961 (N_4961,N_4853,N_4851);
and U4962 (N_4962,N_4850,N_4863);
or U4963 (N_4963,N_4824,N_4861);
and U4964 (N_4964,N_4839,N_4894);
or U4965 (N_4965,N_4864,N_4822);
nor U4966 (N_4966,N_4857,N_4897);
and U4967 (N_4967,N_4858,N_4889);
xnor U4968 (N_4968,N_4885,N_4831);
nor U4969 (N_4969,N_4844,N_4875);
or U4970 (N_4970,N_4869,N_4876);
and U4971 (N_4971,N_4862,N_4803);
and U4972 (N_4972,N_4899,N_4879);
nor U4973 (N_4973,N_4879,N_4844);
or U4974 (N_4974,N_4883,N_4814);
and U4975 (N_4975,N_4849,N_4881);
or U4976 (N_4976,N_4890,N_4884);
and U4977 (N_4977,N_4872,N_4850);
nor U4978 (N_4978,N_4875,N_4832);
and U4979 (N_4979,N_4890,N_4824);
nor U4980 (N_4980,N_4806,N_4873);
or U4981 (N_4981,N_4838,N_4842);
and U4982 (N_4982,N_4899,N_4866);
or U4983 (N_4983,N_4886,N_4827);
nor U4984 (N_4984,N_4892,N_4884);
or U4985 (N_4985,N_4815,N_4834);
nand U4986 (N_4986,N_4884,N_4877);
and U4987 (N_4987,N_4805,N_4881);
or U4988 (N_4988,N_4804,N_4860);
and U4989 (N_4989,N_4821,N_4854);
nor U4990 (N_4990,N_4857,N_4851);
nor U4991 (N_4991,N_4883,N_4852);
or U4992 (N_4992,N_4885,N_4817);
and U4993 (N_4993,N_4852,N_4816);
or U4994 (N_4994,N_4894,N_4810);
and U4995 (N_4995,N_4806,N_4801);
nand U4996 (N_4996,N_4899,N_4882);
nor U4997 (N_4997,N_4803,N_4822);
nor U4998 (N_4998,N_4853,N_4899);
nor U4999 (N_4999,N_4831,N_4812);
nand U5000 (N_5000,N_4945,N_4991);
nand U5001 (N_5001,N_4927,N_4985);
and U5002 (N_5002,N_4993,N_4944);
and U5003 (N_5003,N_4917,N_4942);
nor U5004 (N_5004,N_4987,N_4941);
nand U5005 (N_5005,N_4905,N_4926);
or U5006 (N_5006,N_4957,N_4933);
nor U5007 (N_5007,N_4947,N_4940);
and U5008 (N_5008,N_4952,N_4983);
and U5009 (N_5009,N_4977,N_4998);
or U5010 (N_5010,N_4999,N_4978);
nor U5011 (N_5011,N_4912,N_4907);
and U5012 (N_5012,N_4943,N_4996);
nand U5013 (N_5013,N_4980,N_4958);
nor U5014 (N_5014,N_4913,N_4939);
nor U5015 (N_5015,N_4931,N_4992);
nor U5016 (N_5016,N_4922,N_4916);
or U5017 (N_5017,N_4936,N_4915);
nand U5018 (N_5018,N_4935,N_4904);
and U5019 (N_5019,N_4901,N_4918);
nand U5020 (N_5020,N_4997,N_4911);
nand U5021 (N_5021,N_4966,N_4989);
nor U5022 (N_5022,N_4932,N_4990);
or U5023 (N_5023,N_4994,N_4950);
nor U5024 (N_5024,N_4900,N_4923);
xnor U5025 (N_5025,N_4961,N_4908);
and U5026 (N_5026,N_4930,N_4971);
and U5027 (N_5027,N_4954,N_4903);
nor U5028 (N_5028,N_4948,N_4968);
nand U5029 (N_5029,N_4959,N_4919);
nand U5030 (N_5030,N_4969,N_4986);
nand U5031 (N_5031,N_4960,N_4937);
nand U5032 (N_5032,N_4921,N_4910);
and U5033 (N_5033,N_4963,N_4973);
nand U5034 (N_5034,N_4953,N_4909);
and U5035 (N_5035,N_4979,N_4951);
or U5036 (N_5036,N_4928,N_4949);
nand U5037 (N_5037,N_4955,N_4995);
nand U5038 (N_5038,N_4988,N_4984);
or U5039 (N_5039,N_4974,N_4962);
nand U5040 (N_5040,N_4964,N_4906);
nor U5041 (N_5041,N_4970,N_4967);
or U5042 (N_5042,N_4920,N_4976);
nand U5043 (N_5043,N_4924,N_4975);
nand U5044 (N_5044,N_4929,N_4972);
or U5045 (N_5045,N_4938,N_4902);
nor U5046 (N_5046,N_4925,N_4956);
nand U5047 (N_5047,N_4965,N_4934);
or U5048 (N_5048,N_4914,N_4982);
and U5049 (N_5049,N_4981,N_4946);
nor U5050 (N_5050,N_4978,N_4998);
or U5051 (N_5051,N_4928,N_4941);
or U5052 (N_5052,N_4990,N_4902);
nand U5053 (N_5053,N_4916,N_4948);
nor U5054 (N_5054,N_4914,N_4962);
or U5055 (N_5055,N_4994,N_4965);
or U5056 (N_5056,N_4905,N_4934);
or U5057 (N_5057,N_4975,N_4950);
or U5058 (N_5058,N_4969,N_4914);
nand U5059 (N_5059,N_4930,N_4900);
or U5060 (N_5060,N_4901,N_4977);
and U5061 (N_5061,N_4976,N_4915);
nand U5062 (N_5062,N_4916,N_4908);
and U5063 (N_5063,N_4902,N_4995);
or U5064 (N_5064,N_4970,N_4999);
or U5065 (N_5065,N_4919,N_4987);
or U5066 (N_5066,N_4989,N_4981);
nor U5067 (N_5067,N_4986,N_4975);
nor U5068 (N_5068,N_4912,N_4986);
nor U5069 (N_5069,N_4945,N_4952);
or U5070 (N_5070,N_4921,N_4965);
and U5071 (N_5071,N_4938,N_4978);
and U5072 (N_5072,N_4975,N_4955);
and U5073 (N_5073,N_4997,N_4910);
nor U5074 (N_5074,N_4951,N_4993);
and U5075 (N_5075,N_4958,N_4909);
nor U5076 (N_5076,N_4947,N_4950);
or U5077 (N_5077,N_4993,N_4937);
and U5078 (N_5078,N_4949,N_4919);
and U5079 (N_5079,N_4930,N_4980);
and U5080 (N_5080,N_4940,N_4974);
nor U5081 (N_5081,N_4909,N_4979);
nor U5082 (N_5082,N_4957,N_4916);
nor U5083 (N_5083,N_4920,N_4970);
and U5084 (N_5084,N_4974,N_4930);
xor U5085 (N_5085,N_4932,N_4960);
and U5086 (N_5086,N_4927,N_4954);
and U5087 (N_5087,N_4940,N_4933);
and U5088 (N_5088,N_4987,N_4985);
xnor U5089 (N_5089,N_4997,N_4950);
or U5090 (N_5090,N_4939,N_4923);
nor U5091 (N_5091,N_4966,N_4906);
or U5092 (N_5092,N_4962,N_4935);
or U5093 (N_5093,N_4912,N_4970);
or U5094 (N_5094,N_4916,N_4919);
nand U5095 (N_5095,N_4962,N_4921);
nand U5096 (N_5096,N_4989,N_4924);
nand U5097 (N_5097,N_4914,N_4939);
nor U5098 (N_5098,N_4978,N_4920);
and U5099 (N_5099,N_4902,N_4993);
nand U5100 (N_5100,N_5019,N_5093);
and U5101 (N_5101,N_5020,N_5070);
nand U5102 (N_5102,N_5037,N_5012);
or U5103 (N_5103,N_5087,N_5061);
nand U5104 (N_5104,N_5035,N_5091);
nand U5105 (N_5105,N_5045,N_5011);
and U5106 (N_5106,N_5076,N_5071);
nand U5107 (N_5107,N_5024,N_5090);
or U5108 (N_5108,N_5022,N_5034);
or U5109 (N_5109,N_5082,N_5009);
nor U5110 (N_5110,N_5050,N_5077);
nand U5111 (N_5111,N_5029,N_5028);
nand U5112 (N_5112,N_5072,N_5062);
or U5113 (N_5113,N_5041,N_5096);
and U5114 (N_5114,N_5006,N_5079);
nor U5115 (N_5115,N_5094,N_5051);
and U5116 (N_5116,N_5081,N_5088);
nand U5117 (N_5117,N_5005,N_5064);
nor U5118 (N_5118,N_5057,N_5016);
nor U5119 (N_5119,N_5010,N_5047);
nor U5120 (N_5120,N_5049,N_5092);
and U5121 (N_5121,N_5089,N_5030);
and U5122 (N_5122,N_5053,N_5052);
and U5123 (N_5123,N_5069,N_5073);
and U5124 (N_5124,N_5067,N_5066);
and U5125 (N_5125,N_5084,N_5000);
and U5126 (N_5126,N_5058,N_5074);
nand U5127 (N_5127,N_5098,N_5039);
and U5128 (N_5128,N_5038,N_5097);
and U5129 (N_5129,N_5059,N_5099);
and U5130 (N_5130,N_5083,N_5060);
nor U5131 (N_5131,N_5032,N_5003);
or U5132 (N_5132,N_5031,N_5044);
nor U5133 (N_5133,N_5055,N_5040);
and U5134 (N_5134,N_5065,N_5015);
and U5135 (N_5135,N_5008,N_5017);
nor U5136 (N_5136,N_5007,N_5004);
or U5137 (N_5137,N_5033,N_5048);
nand U5138 (N_5138,N_5046,N_5068);
and U5139 (N_5139,N_5001,N_5021);
nor U5140 (N_5140,N_5080,N_5025);
and U5141 (N_5141,N_5013,N_5026);
or U5142 (N_5142,N_5086,N_5056);
nand U5143 (N_5143,N_5023,N_5063);
and U5144 (N_5144,N_5095,N_5085);
or U5145 (N_5145,N_5027,N_5075);
nor U5146 (N_5146,N_5036,N_5043);
nor U5147 (N_5147,N_5018,N_5002);
nand U5148 (N_5148,N_5014,N_5054);
nand U5149 (N_5149,N_5078,N_5042);
nor U5150 (N_5150,N_5027,N_5093);
and U5151 (N_5151,N_5044,N_5016);
nand U5152 (N_5152,N_5024,N_5068);
or U5153 (N_5153,N_5061,N_5065);
and U5154 (N_5154,N_5042,N_5034);
or U5155 (N_5155,N_5009,N_5044);
or U5156 (N_5156,N_5070,N_5086);
and U5157 (N_5157,N_5064,N_5032);
nor U5158 (N_5158,N_5005,N_5085);
nand U5159 (N_5159,N_5001,N_5019);
or U5160 (N_5160,N_5033,N_5056);
nor U5161 (N_5161,N_5054,N_5012);
and U5162 (N_5162,N_5053,N_5039);
and U5163 (N_5163,N_5007,N_5022);
nor U5164 (N_5164,N_5015,N_5080);
and U5165 (N_5165,N_5084,N_5086);
or U5166 (N_5166,N_5026,N_5052);
and U5167 (N_5167,N_5097,N_5012);
or U5168 (N_5168,N_5092,N_5025);
and U5169 (N_5169,N_5001,N_5071);
or U5170 (N_5170,N_5019,N_5027);
and U5171 (N_5171,N_5032,N_5041);
or U5172 (N_5172,N_5093,N_5072);
nand U5173 (N_5173,N_5045,N_5063);
nand U5174 (N_5174,N_5011,N_5000);
and U5175 (N_5175,N_5038,N_5023);
nor U5176 (N_5176,N_5019,N_5061);
or U5177 (N_5177,N_5095,N_5078);
nor U5178 (N_5178,N_5012,N_5000);
or U5179 (N_5179,N_5070,N_5067);
nand U5180 (N_5180,N_5047,N_5040);
and U5181 (N_5181,N_5091,N_5020);
and U5182 (N_5182,N_5068,N_5035);
and U5183 (N_5183,N_5044,N_5053);
nand U5184 (N_5184,N_5054,N_5092);
nand U5185 (N_5185,N_5015,N_5009);
and U5186 (N_5186,N_5036,N_5001);
or U5187 (N_5187,N_5062,N_5046);
nand U5188 (N_5188,N_5092,N_5038);
nor U5189 (N_5189,N_5070,N_5017);
nand U5190 (N_5190,N_5054,N_5033);
or U5191 (N_5191,N_5053,N_5002);
and U5192 (N_5192,N_5052,N_5030);
and U5193 (N_5193,N_5081,N_5092);
nand U5194 (N_5194,N_5070,N_5042);
nand U5195 (N_5195,N_5035,N_5056);
or U5196 (N_5196,N_5048,N_5043);
nor U5197 (N_5197,N_5023,N_5056);
nand U5198 (N_5198,N_5080,N_5001);
nor U5199 (N_5199,N_5083,N_5098);
nor U5200 (N_5200,N_5180,N_5128);
xnor U5201 (N_5201,N_5155,N_5181);
nand U5202 (N_5202,N_5194,N_5167);
or U5203 (N_5203,N_5150,N_5147);
nor U5204 (N_5204,N_5108,N_5107);
nand U5205 (N_5205,N_5159,N_5101);
or U5206 (N_5206,N_5100,N_5149);
nor U5207 (N_5207,N_5140,N_5179);
nor U5208 (N_5208,N_5175,N_5168);
nor U5209 (N_5209,N_5176,N_5178);
nor U5210 (N_5210,N_5169,N_5127);
nand U5211 (N_5211,N_5191,N_5102);
nand U5212 (N_5212,N_5189,N_5133);
nor U5213 (N_5213,N_5134,N_5142);
nand U5214 (N_5214,N_5170,N_5186);
and U5215 (N_5215,N_5109,N_5113);
or U5216 (N_5216,N_5177,N_5192);
and U5217 (N_5217,N_5145,N_5112);
xor U5218 (N_5218,N_5158,N_5197);
and U5219 (N_5219,N_5132,N_5154);
or U5220 (N_5220,N_5104,N_5123);
and U5221 (N_5221,N_5115,N_5184);
and U5222 (N_5222,N_5137,N_5156);
and U5223 (N_5223,N_5129,N_5152);
or U5224 (N_5224,N_5146,N_5117);
and U5225 (N_5225,N_5124,N_5114);
nor U5226 (N_5226,N_5122,N_5187);
or U5227 (N_5227,N_5118,N_5195);
nor U5228 (N_5228,N_5153,N_5144);
nand U5229 (N_5229,N_5139,N_5130);
or U5230 (N_5230,N_5106,N_5166);
and U5231 (N_5231,N_5141,N_5105);
or U5232 (N_5232,N_5135,N_5116);
and U5233 (N_5233,N_5120,N_5157);
nand U5234 (N_5234,N_5126,N_5143);
nor U5235 (N_5235,N_5162,N_5185);
and U5236 (N_5236,N_5171,N_5161);
and U5237 (N_5237,N_5196,N_5138);
nand U5238 (N_5238,N_5190,N_5136);
nor U5239 (N_5239,N_5163,N_5174);
nand U5240 (N_5240,N_5164,N_5111);
nor U5241 (N_5241,N_5183,N_5103);
and U5242 (N_5242,N_5165,N_5148);
nand U5243 (N_5243,N_5131,N_5193);
nand U5244 (N_5244,N_5173,N_5172);
nor U5245 (N_5245,N_5198,N_5160);
nor U5246 (N_5246,N_5151,N_5119);
nand U5247 (N_5247,N_5182,N_5125);
nand U5248 (N_5248,N_5110,N_5199);
and U5249 (N_5249,N_5188,N_5121);
nand U5250 (N_5250,N_5105,N_5195);
and U5251 (N_5251,N_5160,N_5124);
nand U5252 (N_5252,N_5134,N_5112);
nor U5253 (N_5253,N_5156,N_5142);
nor U5254 (N_5254,N_5169,N_5148);
nor U5255 (N_5255,N_5178,N_5105);
nor U5256 (N_5256,N_5115,N_5164);
nand U5257 (N_5257,N_5191,N_5184);
or U5258 (N_5258,N_5141,N_5186);
or U5259 (N_5259,N_5151,N_5130);
and U5260 (N_5260,N_5154,N_5153);
nand U5261 (N_5261,N_5185,N_5145);
nor U5262 (N_5262,N_5116,N_5173);
and U5263 (N_5263,N_5169,N_5185);
xnor U5264 (N_5264,N_5178,N_5199);
nor U5265 (N_5265,N_5162,N_5197);
nor U5266 (N_5266,N_5108,N_5145);
and U5267 (N_5267,N_5143,N_5177);
or U5268 (N_5268,N_5164,N_5123);
nor U5269 (N_5269,N_5148,N_5143);
or U5270 (N_5270,N_5123,N_5100);
and U5271 (N_5271,N_5162,N_5142);
xor U5272 (N_5272,N_5116,N_5161);
or U5273 (N_5273,N_5104,N_5141);
or U5274 (N_5274,N_5118,N_5153);
nor U5275 (N_5275,N_5172,N_5117);
nor U5276 (N_5276,N_5110,N_5115);
and U5277 (N_5277,N_5158,N_5176);
and U5278 (N_5278,N_5189,N_5129);
nand U5279 (N_5279,N_5117,N_5165);
nor U5280 (N_5280,N_5114,N_5147);
nand U5281 (N_5281,N_5113,N_5171);
and U5282 (N_5282,N_5146,N_5103);
nor U5283 (N_5283,N_5157,N_5191);
nor U5284 (N_5284,N_5154,N_5115);
nand U5285 (N_5285,N_5134,N_5165);
or U5286 (N_5286,N_5123,N_5198);
nand U5287 (N_5287,N_5128,N_5183);
or U5288 (N_5288,N_5122,N_5151);
or U5289 (N_5289,N_5193,N_5155);
or U5290 (N_5290,N_5101,N_5156);
nand U5291 (N_5291,N_5182,N_5160);
and U5292 (N_5292,N_5161,N_5179);
or U5293 (N_5293,N_5133,N_5174);
nor U5294 (N_5294,N_5108,N_5160);
nand U5295 (N_5295,N_5144,N_5186);
nand U5296 (N_5296,N_5121,N_5111);
nand U5297 (N_5297,N_5139,N_5117);
nand U5298 (N_5298,N_5165,N_5105);
or U5299 (N_5299,N_5186,N_5115);
nand U5300 (N_5300,N_5238,N_5262);
nand U5301 (N_5301,N_5216,N_5258);
or U5302 (N_5302,N_5245,N_5236);
nor U5303 (N_5303,N_5280,N_5277);
and U5304 (N_5304,N_5234,N_5239);
nor U5305 (N_5305,N_5235,N_5213);
nand U5306 (N_5306,N_5291,N_5279);
and U5307 (N_5307,N_5287,N_5275);
nand U5308 (N_5308,N_5210,N_5225);
nand U5309 (N_5309,N_5250,N_5290);
and U5310 (N_5310,N_5267,N_5282);
or U5311 (N_5311,N_5272,N_5222);
or U5312 (N_5312,N_5233,N_5284);
and U5313 (N_5313,N_5221,N_5237);
nand U5314 (N_5314,N_5251,N_5220);
nand U5315 (N_5315,N_5281,N_5231);
nor U5316 (N_5316,N_5283,N_5246);
nand U5317 (N_5317,N_5298,N_5259);
or U5318 (N_5318,N_5202,N_5241);
and U5319 (N_5319,N_5200,N_5212);
and U5320 (N_5320,N_5209,N_5226);
and U5321 (N_5321,N_5203,N_5295);
or U5322 (N_5322,N_5296,N_5261);
nand U5323 (N_5323,N_5269,N_5242);
nor U5324 (N_5324,N_5276,N_5265);
nand U5325 (N_5325,N_5297,N_5228);
or U5326 (N_5326,N_5255,N_5208);
nor U5327 (N_5327,N_5299,N_5292);
nor U5328 (N_5328,N_5227,N_5217);
nand U5329 (N_5329,N_5252,N_5278);
and U5330 (N_5330,N_5201,N_5268);
or U5331 (N_5331,N_5293,N_5243);
or U5332 (N_5332,N_5256,N_5247);
or U5333 (N_5333,N_5285,N_5214);
nand U5334 (N_5334,N_5218,N_5288);
and U5335 (N_5335,N_5229,N_5206);
nor U5336 (N_5336,N_5232,N_5240);
nor U5337 (N_5337,N_5264,N_5248);
nor U5338 (N_5338,N_5230,N_5253);
nand U5339 (N_5339,N_5257,N_5263);
nand U5340 (N_5340,N_5273,N_5205);
xor U5341 (N_5341,N_5219,N_5274);
nand U5342 (N_5342,N_5223,N_5270);
or U5343 (N_5343,N_5254,N_5289);
nand U5344 (N_5344,N_5224,N_5207);
and U5345 (N_5345,N_5266,N_5211);
or U5346 (N_5346,N_5271,N_5204);
and U5347 (N_5347,N_5215,N_5249);
nand U5348 (N_5348,N_5260,N_5244);
or U5349 (N_5349,N_5286,N_5294);
nor U5350 (N_5350,N_5282,N_5270);
nor U5351 (N_5351,N_5260,N_5229);
nand U5352 (N_5352,N_5234,N_5262);
and U5353 (N_5353,N_5270,N_5267);
nand U5354 (N_5354,N_5216,N_5283);
or U5355 (N_5355,N_5283,N_5267);
nor U5356 (N_5356,N_5244,N_5270);
and U5357 (N_5357,N_5288,N_5273);
and U5358 (N_5358,N_5238,N_5272);
and U5359 (N_5359,N_5278,N_5230);
and U5360 (N_5360,N_5225,N_5261);
nand U5361 (N_5361,N_5273,N_5265);
nand U5362 (N_5362,N_5262,N_5233);
and U5363 (N_5363,N_5252,N_5285);
or U5364 (N_5364,N_5243,N_5288);
and U5365 (N_5365,N_5282,N_5235);
nand U5366 (N_5366,N_5220,N_5270);
nor U5367 (N_5367,N_5204,N_5298);
or U5368 (N_5368,N_5277,N_5236);
and U5369 (N_5369,N_5296,N_5293);
or U5370 (N_5370,N_5272,N_5274);
and U5371 (N_5371,N_5240,N_5243);
and U5372 (N_5372,N_5247,N_5214);
nor U5373 (N_5373,N_5217,N_5257);
and U5374 (N_5374,N_5209,N_5262);
nor U5375 (N_5375,N_5200,N_5218);
nand U5376 (N_5376,N_5266,N_5257);
nor U5377 (N_5377,N_5276,N_5217);
or U5378 (N_5378,N_5298,N_5231);
or U5379 (N_5379,N_5237,N_5263);
nand U5380 (N_5380,N_5295,N_5275);
nor U5381 (N_5381,N_5248,N_5262);
and U5382 (N_5382,N_5287,N_5227);
nand U5383 (N_5383,N_5240,N_5206);
or U5384 (N_5384,N_5258,N_5239);
and U5385 (N_5385,N_5216,N_5210);
nor U5386 (N_5386,N_5258,N_5233);
and U5387 (N_5387,N_5205,N_5217);
nand U5388 (N_5388,N_5221,N_5250);
nor U5389 (N_5389,N_5296,N_5219);
nand U5390 (N_5390,N_5283,N_5239);
nand U5391 (N_5391,N_5275,N_5204);
nor U5392 (N_5392,N_5228,N_5235);
or U5393 (N_5393,N_5260,N_5280);
nand U5394 (N_5394,N_5209,N_5260);
or U5395 (N_5395,N_5265,N_5208);
or U5396 (N_5396,N_5208,N_5271);
or U5397 (N_5397,N_5284,N_5287);
or U5398 (N_5398,N_5272,N_5216);
or U5399 (N_5399,N_5226,N_5248);
nand U5400 (N_5400,N_5314,N_5320);
nor U5401 (N_5401,N_5303,N_5328);
or U5402 (N_5402,N_5329,N_5358);
or U5403 (N_5403,N_5307,N_5334);
or U5404 (N_5404,N_5313,N_5368);
or U5405 (N_5405,N_5374,N_5344);
and U5406 (N_5406,N_5353,N_5365);
and U5407 (N_5407,N_5355,N_5361);
nor U5408 (N_5408,N_5388,N_5386);
or U5409 (N_5409,N_5336,N_5362);
nand U5410 (N_5410,N_5311,N_5341);
nor U5411 (N_5411,N_5327,N_5308);
nor U5412 (N_5412,N_5384,N_5349);
and U5413 (N_5413,N_5339,N_5376);
or U5414 (N_5414,N_5345,N_5318);
and U5415 (N_5415,N_5338,N_5330);
nand U5416 (N_5416,N_5323,N_5385);
nor U5417 (N_5417,N_5387,N_5393);
nand U5418 (N_5418,N_5380,N_5326);
and U5419 (N_5419,N_5397,N_5305);
nor U5420 (N_5420,N_5371,N_5300);
nand U5421 (N_5421,N_5373,N_5315);
xnor U5422 (N_5422,N_5348,N_5390);
and U5423 (N_5423,N_5394,N_5302);
nand U5424 (N_5424,N_5398,N_5331);
and U5425 (N_5425,N_5350,N_5322);
nor U5426 (N_5426,N_5379,N_5378);
nand U5427 (N_5427,N_5316,N_5391);
nor U5428 (N_5428,N_5333,N_5360);
or U5429 (N_5429,N_5366,N_5346);
nand U5430 (N_5430,N_5306,N_5377);
nor U5431 (N_5431,N_5312,N_5351);
nor U5432 (N_5432,N_5301,N_5382);
nor U5433 (N_5433,N_5340,N_5342);
and U5434 (N_5434,N_5337,N_5364);
nor U5435 (N_5435,N_5399,N_5372);
and U5436 (N_5436,N_5325,N_5343);
nor U5437 (N_5437,N_5319,N_5347);
and U5438 (N_5438,N_5324,N_5367);
nor U5439 (N_5439,N_5392,N_5359);
nand U5440 (N_5440,N_5370,N_5369);
nor U5441 (N_5441,N_5309,N_5383);
and U5442 (N_5442,N_5304,N_5363);
and U5443 (N_5443,N_5356,N_5375);
and U5444 (N_5444,N_5335,N_5396);
nand U5445 (N_5445,N_5381,N_5354);
nand U5446 (N_5446,N_5395,N_5332);
xnor U5447 (N_5447,N_5310,N_5321);
or U5448 (N_5448,N_5352,N_5317);
nand U5449 (N_5449,N_5389,N_5357);
nor U5450 (N_5450,N_5348,N_5303);
or U5451 (N_5451,N_5356,N_5368);
and U5452 (N_5452,N_5308,N_5307);
or U5453 (N_5453,N_5326,N_5362);
nand U5454 (N_5454,N_5304,N_5311);
nand U5455 (N_5455,N_5346,N_5303);
and U5456 (N_5456,N_5354,N_5372);
nor U5457 (N_5457,N_5396,N_5305);
or U5458 (N_5458,N_5364,N_5323);
nand U5459 (N_5459,N_5375,N_5388);
nand U5460 (N_5460,N_5355,N_5382);
nor U5461 (N_5461,N_5378,N_5351);
nor U5462 (N_5462,N_5313,N_5322);
nand U5463 (N_5463,N_5337,N_5347);
and U5464 (N_5464,N_5351,N_5303);
nor U5465 (N_5465,N_5396,N_5321);
or U5466 (N_5466,N_5365,N_5317);
and U5467 (N_5467,N_5311,N_5336);
nor U5468 (N_5468,N_5327,N_5367);
or U5469 (N_5469,N_5343,N_5371);
nand U5470 (N_5470,N_5363,N_5323);
or U5471 (N_5471,N_5389,N_5390);
nor U5472 (N_5472,N_5384,N_5357);
nor U5473 (N_5473,N_5306,N_5398);
xnor U5474 (N_5474,N_5341,N_5393);
nand U5475 (N_5475,N_5310,N_5345);
or U5476 (N_5476,N_5382,N_5357);
or U5477 (N_5477,N_5338,N_5376);
nand U5478 (N_5478,N_5300,N_5305);
xnor U5479 (N_5479,N_5310,N_5358);
and U5480 (N_5480,N_5335,N_5374);
and U5481 (N_5481,N_5357,N_5350);
nor U5482 (N_5482,N_5387,N_5350);
and U5483 (N_5483,N_5388,N_5368);
or U5484 (N_5484,N_5392,N_5352);
and U5485 (N_5485,N_5350,N_5372);
nand U5486 (N_5486,N_5349,N_5313);
or U5487 (N_5487,N_5353,N_5327);
and U5488 (N_5488,N_5399,N_5344);
nand U5489 (N_5489,N_5367,N_5381);
or U5490 (N_5490,N_5380,N_5367);
and U5491 (N_5491,N_5388,N_5315);
or U5492 (N_5492,N_5367,N_5334);
and U5493 (N_5493,N_5315,N_5391);
or U5494 (N_5494,N_5323,N_5313);
nor U5495 (N_5495,N_5399,N_5355);
and U5496 (N_5496,N_5399,N_5338);
xnor U5497 (N_5497,N_5330,N_5340);
nand U5498 (N_5498,N_5303,N_5368);
or U5499 (N_5499,N_5352,N_5300);
nand U5500 (N_5500,N_5441,N_5445);
nor U5501 (N_5501,N_5411,N_5432);
and U5502 (N_5502,N_5497,N_5425);
nand U5503 (N_5503,N_5403,N_5480);
and U5504 (N_5504,N_5485,N_5412);
nor U5505 (N_5505,N_5422,N_5469);
nand U5506 (N_5506,N_5465,N_5494);
nand U5507 (N_5507,N_5484,N_5461);
nand U5508 (N_5508,N_5451,N_5434);
and U5509 (N_5509,N_5456,N_5401);
or U5510 (N_5510,N_5452,N_5466);
and U5511 (N_5511,N_5433,N_5447);
nand U5512 (N_5512,N_5459,N_5492);
nor U5513 (N_5513,N_5431,N_5428);
nand U5514 (N_5514,N_5487,N_5458);
xor U5515 (N_5515,N_5474,N_5440);
nand U5516 (N_5516,N_5442,N_5410);
nor U5517 (N_5517,N_5439,N_5409);
and U5518 (N_5518,N_5430,N_5438);
nor U5519 (N_5519,N_5478,N_5423);
or U5520 (N_5520,N_5473,N_5464);
nor U5521 (N_5521,N_5470,N_5468);
nand U5522 (N_5522,N_5402,N_5449);
or U5523 (N_5523,N_5499,N_5455);
nor U5524 (N_5524,N_5475,N_5496);
or U5525 (N_5525,N_5426,N_5407);
nand U5526 (N_5526,N_5408,N_5454);
or U5527 (N_5527,N_5437,N_5463);
and U5528 (N_5528,N_5435,N_5453);
and U5529 (N_5529,N_5405,N_5400);
nand U5530 (N_5530,N_5419,N_5482);
nand U5531 (N_5531,N_5424,N_5413);
nor U5532 (N_5532,N_5476,N_5489);
nor U5533 (N_5533,N_5444,N_5490);
nand U5534 (N_5534,N_5479,N_5429);
nor U5535 (N_5535,N_5443,N_5477);
or U5536 (N_5536,N_5498,N_5427);
nand U5537 (N_5537,N_5421,N_5495);
nor U5538 (N_5538,N_5462,N_5417);
nand U5539 (N_5539,N_5416,N_5493);
or U5540 (N_5540,N_5486,N_5460);
or U5541 (N_5541,N_5481,N_5414);
and U5542 (N_5542,N_5472,N_5491);
or U5543 (N_5543,N_5406,N_5448);
and U5544 (N_5544,N_5446,N_5404);
nand U5545 (N_5545,N_5471,N_5483);
and U5546 (N_5546,N_5415,N_5467);
or U5547 (N_5547,N_5488,N_5457);
nand U5548 (N_5548,N_5450,N_5436);
nor U5549 (N_5549,N_5418,N_5420);
and U5550 (N_5550,N_5410,N_5448);
or U5551 (N_5551,N_5404,N_5457);
or U5552 (N_5552,N_5400,N_5426);
nor U5553 (N_5553,N_5489,N_5492);
and U5554 (N_5554,N_5455,N_5430);
and U5555 (N_5555,N_5492,N_5438);
nor U5556 (N_5556,N_5496,N_5480);
nand U5557 (N_5557,N_5441,N_5443);
nand U5558 (N_5558,N_5446,N_5487);
or U5559 (N_5559,N_5465,N_5412);
nor U5560 (N_5560,N_5447,N_5432);
nand U5561 (N_5561,N_5447,N_5470);
nand U5562 (N_5562,N_5429,N_5447);
nand U5563 (N_5563,N_5467,N_5440);
or U5564 (N_5564,N_5424,N_5447);
and U5565 (N_5565,N_5497,N_5456);
nand U5566 (N_5566,N_5477,N_5447);
nor U5567 (N_5567,N_5424,N_5462);
nor U5568 (N_5568,N_5465,N_5410);
nor U5569 (N_5569,N_5429,N_5488);
nor U5570 (N_5570,N_5404,N_5422);
and U5571 (N_5571,N_5447,N_5490);
nand U5572 (N_5572,N_5445,N_5466);
nor U5573 (N_5573,N_5477,N_5469);
or U5574 (N_5574,N_5460,N_5467);
and U5575 (N_5575,N_5462,N_5433);
nor U5576 (N_5576,N_5446,N_5477);
xor U5577 (N_5577,N_5436,N_5477);
and U5578 (N_5578,N_5454,N_5432);
nand U5579 (N_5579,N_5459,N_5491);
nand U5580 (N_5580,N_5424,N_5458);
and U5581 (N_5581,N_5412,N_5432);
nand U5582 (N_5582,N_5434,N_5401);
and U5583 (N_5583,N_5459,N_5415);
nor U5584 (N_5584,N_5495,N_5489);
and U5585 (N_5585,N_5423,N_5425);
and U5586 (N_5586,N_5489,N_5453);
nor U5587 (N_5587,N_5488,N_5426);
nand U5588 (N_5588,N_5405,N_5498);
and U5589 (N_5589,N_5432,N_5493);
nand U5590 (N_5590,N_5432,N_5478);
nand U5591 (N_5591,N_5422,N_5412);
and U5592 (N_5592,N_5410,N_5408);
and U5593 (N_5593,N_5450,N_5466);
nor U5594 (N_5594,N_5406,N_5488);
or U5595 (N_5595,N_5421,N_5480);
and U5596 (N_5596,N_5418,N_5403);
nand U5597 (N_5597,N_5463,N_5492);
nand U5598 (N_5598,N_5478,N_5490);
nand U5599 (N_5599,N_5485,N_5495);
nand U5600 (N_5600,N_5555,N_5587);
nand U5601 (N_5601,N_5570,N_5536);
nand U5602 (N_5602,N_5580,N_5518);
or U5603 (N_5603,N_5503,N_5520);
nor U5604 (N_5604,N_5532,N_5540);
nor U5605 (N_5605,N_5509,N_5523);
or U5606 (N_5606,N_5524,N_5565);
or U5607 (N_5607,N_5557,N_5586);
and U5608 (N_5608,N_5569,N_5514);
and U5609 (N_5609,N_5581,N_5527);
and U5610 (N_5610,N_5547,N_5559);
nand U5611 (N_5611,N_5575,N_5571);
nor U5612 (N_5612,N_5543,N_5583);
and U5613 (N_5613,N_5566,N_5572);
nor U5614 (N_5614,N_5528,N_5592);
nand U5615 (N_5615,N_5576,N_5539);
nand U5616 (N_5616,N_5545,N_5541);
and U5617 (N_5617,N_5549,N_5568);
nand U5618 (N_5618,N_5567,N_5594);
nand U5619 (N_5619,N_5548,N_5506);
or U5620 (N_5620,N_5582,N_5554);
or U5621 (N_5621,N_5551,N_5538);
or U5622 (N_5622,N_5501,N_5517);
nand U5623 (N_5623,N_5537,N_5530);
or U5624 (N_5624,N_5553,N_5525);
nor U5625 (N_5625,N_5516,N_5510);
and U5626 (N_5626,N_5574,N_5508);
nor U5627 (N_5627,N_5552,N_5561);
or U5628 (N_5628,N_5529,N_5526);
and U5629 (N_5629,N_5550,N_5534);
nand U5630 (N_5630,N_5546,N_5579);
nor U5631 (N_5631,N_5596,N_5585);
nor U5632 (N_5632,N_5584,N_5533);
or U5633 (N_5633,N_5502,N_5505);
nor U5634 (N_5634,N_5500,N_5512);
and U5635 (N_5635,N_5544,N_5597);
nor U5636 (N_5636,N_5519,N_5511);
and U5637 (N_5637,N_5598,N_5578);
or U5638 (N_5638,N_5558,N_5589);
nor U5639 (N_5639,N_5591,N_5588);
and U5640 (N_5640,N_5515,N_5562);
nand U5641 (N_5641,N_5595,N_5564);
or U5642 (N_5642,N_5590,N_5599);
nor U5643 (N_5643,N_5542,N_5560);
and U5644 (N_5644,N_5521,N_5593);
or U5645 (N_5645,N_5531,N_5577);
nor U5646 (N_5646,N_5535,N_5504);
nand U5647 (N_5647,N_5513,N_5563);
or U5648 (N_5648,N_5556,N_5507);
and U5649 (N_5649,N_5522,N_5573);
nand U5650 (N_5650,N_5521,N_5538);
or U5651 (N_5651,N_5556,N_5517);
nor U5652 (N_5652,N_5500,N_5551);
nor U5653 (N_5653,N_5577,N_5526);
or U5654 (N_5654,N_5542,N_5510);
or U5655 (N_5655,N_5544,N_5560);
nand U5656 (N_5656,N_5544,N_5580);
xnor U5657 (N_5657,N_5558,N_5591);
and U5658 (N_5658,N_5501,N_5526);
or U5659 (N_5659,N_5538,N_5596);
nor U5660 (N_5660,N_5520,N_5536);
nand U5661 (N_5661,N_5581,N_5584);
nor U5662 (N_5662,N_5566,N_5596);
or U5663 (N_5663,N_5513,N_5552);
nand U5664 (N_5664,N_5599,N_5519);
or U5665 (N_5665,N_5523,N_5517);
xnor U5666 (N_5666,N_5553,N_5516);
and U5667 (N_5667,N_5590,N_5541);
or U5668 (N_5668,N_5588,N_5525);
or U5669 (N_5669,N_5525,N_5573);
nor U5670 (N_5670,N_5507,N_5573);
xor U5671 (N_5671,N_5560,N_5581);
or U5672 (N_5672,N_5501,N_5536);
xnor U5673 (N_5673,N_5560,N_5537);
and U5674 (N_5674,N_5548,N_5521);
nor U5675 (N_5675,N_5574,N_5586);
or U5676 (N_5676,N_5597,N_5593);
nor U5677 (N_5677,N_5514,N_5593);
or U5678 (N_5678,N_5529,N_5578);
and U5679 (N_5679,N_5504,N_5570);
nor U5680 (N_5680,N_5511,N_5537);
or U5681 (N_5681,N_5558,N_5581);
nor U5682 (N_5682,N_5500,N_5562);
and U5683 (N_5683,N_5559,N_5566);
or U5684 (N_5684,N_5578,N_5570);
or U5685 (N_5685,N_5533,N_5553);
nand U5686 (N_5686,N_5596,N_5574);
nor U5687 (N_5687,N_5570,N_5592);
and U5688 (N_5688,N_5535,N_5589);
nand U5689 (N_5689,N_5546,N_5591);
nor U5690 (N_5690,N_5536,N_5533);
nand U5691 (N_5691,N_5522,N_5535);
and U5692 (N_5692,N_5520,N_5554);
nor U5693 (N_5693,N_5592,N_5580);
or U5694 (N_5694,N_5503,N_5586);
nor U5695 (N_5695,N_5518,N_5538);
nand U5696 (N_5696,N_5535,N_5594);
xor U5697 (N_5697,N_5597,N_5522);
and U5698 (N_5698,N_5542,N_5515);
and U5699 (N_5699,N_5548,N_5591);
or U5700 (N_5700,N_5627,N_5673);
and U5701 (N_5701,N_5622,N_5638);
and U5702 (N_5702,N_5642,N_5679);
nand U5703 (N_5703,N_5606,N_5637);
and U5704 (N_5704,N_5662,N_5672);
and U5705 (N_5705,N_5665,N_5625);
or U5706 (N_5706,N_5621,N_5676);
nor U5707 (N_5707,N_5615,N_5623);
nand U5708 (N_5708,N_5678,N_5616);
and U5709 (N_5709,N_5674,N_5683);
or U5710 (N_5710,N_5653,N_5641);
or U5711 (N_5711,N_5652,N_5689);
nor U5712 (N_5712,N_5608,N_5670);
nor U5713 (N_5713,N_5695,N_5669);
and U5714 (N_5714,N_5635,N_5660);
or U5715 (N_5715,N_5655,N_5697);
nor U5716 (N_5716,N_5640,N_5656);
nand U5717 (N_5717,N_5691,N_5643);
or U5718 (N_5718,N_5610,N_5630);
nor U5719 (N_5719,N_5647,N_5646);
and U5720 (N_5720,N_5618,N_5696);
nor U5721 (N_5721,N_5684,N_5667);
or U5722 (N_5722,N_5602,N_5657);
or U5723 (N_5723,N_5694,N_5686);
or U5724 (N_5724,N_5659,N_5663);
nand U5725 (N_5725,N_5620,N_5648);
nor U5726 (N_5726,N_5631,N_5645);
or U5727 (N_5727,N_5675,N_5613);
and U5728 (N_5728,N_5668,N_5639);
nand U5729 (N_5729,N_5628,N_5690);
nor U5730 (N_5730,N_5603,N_5685);
or U5731 (N_5731,N_5633,N_5666);
or U5732 (N_5732,N_5692,N_5601);
xnor U5733 (N_5733,N_5614,N_5612);
or U5734 (N_5734,N_5664,N_5682);
or U5735 (N_5735,N_5680,N_5626);
and U5736 (N_5736,N_5699,N_5693);
nand U5737 (N_5737,N_5617,N_5600);
and U5738 (N_5738,N_5671,N_5619);
nor U5739 (N_5739,N_5687,N_5611);
and U5740 (N_5740,N_5681,N_5607);
nor U5741 (N_5741,N_5609,N_5698);
nand U5742 (N_5742,N_5624,N_5650);
and U5743 (N_5743,N_5636,N_5654);
and U5744 (N_5744,N_5634,N_5651);
and U5745 (N_5745,N_5629,N_5649);
nand U5746 (N_5746,N_5604,N_5644);
or U5747 (N_5747,N_5688,N_5658);
nand U5748 (N_5748,N_5632,N_5605);
and U5749 (N_5749,N_5677,N_5661);
and U5750 (N_5750,N_5609,N_5613);
nand U5751 (N_5751,N_5658,N_5627);
and U5752 (N_5752,N_5677,N_5644);
or U5753 (N_5753,N_5678,N_5611);
or U5754 (N_5754,N_5656,N_5668);
or U5755 (N_5755,N_5607,N_5686);
nand U5756 (N_5756,N_5675,N_5663);
nor U5757 (N_5757,N_5672,N_5657);
nand U5758 (N_5758,N_5621,N_5674);
and U5759 (N_5759,N_5657,N_5610);
and U5760 (N_5760,N_5623,N_5619);
or U5761 (N_5761,N_5684,N_5658);
xor U5762 (N_5762,N_5661,N_5604);
xor U5763 (N_5763,N_5671,N_5611);
or U5764 (N_5764,N_5632,N_5674);
and U5765 (N_5765,N_5615,N_5656);
and U5766 (N_5766,N_5679,N_5677);
or U5767 (N_5767,N_5637,N_5629);
nand U5768 (N_5768,N_5652,N_5667);
or U5769 (N_5769,N_5643,N_5611);
nand U5770 (N_5770,N_5677,N_5675);
nor U5771 (N_5771,N_5698,N_5680);
and U5772 (N_5772,N_5688,N_5654);
and U5773 (N_5773,N_5669,N_5615);
and U5774 (N_5774,N_5666,N_5665);
and U5775 (N_5775,N_5628,N_5656);
nor U5776 (N_5776,N_5611,N_5668);
nor U5777 (N_5777,N_5683,N_5660);
nor U5778 (N_5778,N_5649,N_5603);
or U5779 (N_5779,N_5678,N_5603);
or U5780 (N_5780,N_5659,N_5655);
and U5781 (N_5781,N_5636,N_5602);
nor U5782 (N_5782,N_5605,N_5684);
or U5783 (N_5783,N_5685,N_5670);
or U5784 (N_5784,N_5615,N_5686);
and U5785 (N_5785,N_5669,N_5693);
nand U5786 (N_5786,N_5657,N_5653);
nand U5787 (N_5787,N_5653,N_5629);
nand U5788 (N_5788,N_5642,N_5683);
or U5789 (N_5789,N_5661,N_5603);
nand U5790 (N_5790,N_5668,N_5641);
or U5791 (N_5791,N_5665,N_5651);
and U5792 (N_5792,N_5601,N_5666);
nor U5793 (N_5793,N_5645,N_5677);
nor U5794 (N_5794,N_5620,N_5639);
or U5795 (N_5795,N_5630,N_5642);
or U5796 (N_5796,N_5612,N_5698);
nand U5797 (N_5797,N_5643,N_5625);
nor U5798 (N_5798,N_5698,N_5603);
nor U5799 (N_5799,N_5607,N_5653);
nor U5800 (N_5800,N_5786,N_5778);
nand U5801 (N_5801,N_5735,N_5783);
nand U5802 (N_5802,N_5775,N_5729);
or U5803 (N_5803,N_5741,N_5701);
nand U5804 (N_5804,N_5766,N_5763);
nor U5805 (N_5805,N_5710,N_5739);
nand U5806 (N_5806,N_5734,N_5757);
and U5807 (N_5807,N_5762,N_5780);
and U5808 (N_5808,N_5746,N_5707);
nand U5809 (N_5809,N_5726,N_5787);
nor U5810 (N_5810,N_5720,N_5719);
nor U5811 (N_5811,N_5718,N_5714);
nor U5812 (N_5812,N_5737,N_5736);
nor U5813 (N_5813,N_5785,N_5788);
nand U5814 (N_5814,N_5703,N_5721);
and U5815 (N_5815,N_5700,N_5754);
nand U5816 (N_5816,N_5761,N_5769);
or U5817 (N_5817,N_5705,N_5752);
and U5818 (N_5818,N_5793,N_5740);
nor U5819 (N_5819,N_5794,N_5776);
nor U5820 (N_5820,N_5744,N_5795);
or U5821 (N_5821,N_5773,N_5723);
and U5822 (N_5822,N_5756,N_5731);
nand U5823 (N_5823,N_5709,N_5704);
or U5824 (N_5824,N_5742,N_5706);
nor U5825 (N_5825,N_5765,N_5747);
nor U5826 (N_5826,N_5722,N_5751);
or U5827 (N_5827,N_5784,N_5712);
nand U5828 (N_5828,N_5724,N_5792);
nor U5829 (N_5829,N_5799,N_5713);
and U5830 (N_5830,N_5750,N_5758);
nand U5831 (N_5831,N_5725,N_5716);
and U5832 (N_5832,N_5755,N_5791);
nor U5833 (N_5833,N_5745,N_5702);
xnor U5834 (N_5834,N_5733,N_5753);
or U5835 (N_5835,N_5796,N_5711);
nor U5836 (N_5836,N_5782,N_5790);
nand U5837 (N_5837,N_5743,N_5759);
nand U5838 (N_5838,N_5708,N_5770);
nand U5839 (N_5839,N_5789,N_5764);
nand U5840 (N_5840,N_5760,N_5728);
xnor U5841 (N_5841,N_5748,N_5774);
nor U5842 (N_5842,N_5777,N_5732);
or U5843 (N_5843,N_5767,N_5749);
nor U5844 (N_5844,N_5715,N_5771);
or U5845 (N_5845,N_5738,N_5768);
nand U5846 (N_5846,N_5779,N_5727);
xnor U5847 (N_5847,N_5717,N_5730);
nand U5848 (N_5848,N_5798,N_5781);
nor U5849 (N_5849,N_5772,N_5797);
or U5850 (N_5850,N_5767,N_5790);
nand U5851 (N_5851,N_5724,N_5711);
or U5852 (N_5852,N_5772,N_5708);
nand U5853 (N_5853,N_5713,N_5727);
or U5854 (N_5854,N_5770,N_5718);
xor U5855 (N_5855,N_5799,N_5754);
and U5856 (N_5856,N_5717,N_5753);
xor U5857 (N_5857,N_5740,N_5747);
or U5858 (N_5858,N_5770,N_5725);
nor U5859 (N_5859,N_5735,N_5736);
nor U5860 (N_5860,N_5756,N_5723);
nor U5861 (N_5861,N_5773,N_5762);
nand U5862 (N_5862,N_5799,N_5743);
and U5863 (N_5863,N_5736,N_5777);
nor U5864 (N_5864,N_5718,N_5721);
and U5865 (N_5865,N_5745,N_5725);
and U5866 (N_5866,N_5782,N_5700);
or U5867 (N_5867,N_5797,N_5760);
nand U5868 (N_5868,N_5731,N_5785);
nand U5869 (N_5869,N_5791,N_5729);
and U5870 (N_5870,N_5724,N_5775);
nand U5871 (N_5871,N_5718,N_5755);
and U5872 (N_5872,N_5772,N_5765);
nor U5873 (N_5873,N_5747,N_5795);
or U5874 (N_5874,N_5760,N_5790);
and U5875 (N_5875,N_5724,N_5743);
or U5876 (N_5876,N_5718,N_5778);
or U5877 (N_5877,N_5797,N_5707);
nor U5878 (N_5878,N_5707,N_5744);
nand U5879 (N_5879,N_5782,N_5722);
and U5880 (N_5880,N_5761,N_5716);
and U5881 (N_5881,N_5769,N_5749);
nor U5882 (N_5882,N_5738,N_5792);
nand U5883 (N_5883,N_5715,N_5738);
or U5884 (N_5884,N_5763,N_5738);
or U5885 (N_5885,N_5716,N_5798);
nand U5886 (N_5886,N_5719,N_5741);
nor U5887 (N_5887,N_5788,N_5729);
nor U5888 (N_5888,N_5782,N_5709);
or U5889 (N_5889,N_5773,N_5702);
nand U5890 (N_5890,N_5791,N_5793);
and U5891 (N_5891,N_5794,N_5753);
nand U5892 (N_5892,N_5782,N_5705);
nor U5893 (N_5893,N_5735,N_5754);
nor U5894 (N_5894,N_5786,N_5744);
nand U5895 (N_5895,N_5709,N_5735);
xor U5896 (N_5896,N_5786,N_5795);
or U5897 (N_5897,N_5784,N_5744);
nor U5898 (N_5898,N_5764,N_5721);
nor U5899 (N_5899,N_5770,N_5720);
nand U5900 (N_5900,N_5874,N_5808);
and U5901 (N_5901,N_5870,N_5803);
nor U5902 (N_5902,N_5856,N_5836);
nor U5903 (N_5903,N_5809,N_5844);
and U5904 (N_5904,N_5854,N_5812);
or U5905 (N_5905,N_5866,N_5857);
nand U5906 (N_5906,N_5817,N_5823);
or U5907 (N_5907,N_5828,N_5816);
xor U5908 (N_5908,N_5889,N_5864);
and U5909 (N_5909,N_5883,N_5894);
nand U5910 (N_5910,N_5881,N_5859);
and U5911 (N_5911,N_5861,N_5867);
nor U5912 (N_5912,N_5813,N_5820);
and U5913 (N_5913,N_5834,N_5830);
and U5914 (N_5914,N_5878,N_5818);
nor U5915 (N_5915,N_5835,N_5827);
xor U5916 (N_5916,N_5855,N_5877);
nor U5917 (N_5917,N_5829,N_5806);
nor U5918 (N_5918,N_5839,N_5893);
nand U5919 (N_5919,N_5884,N_5862);
and U5920 (N_5920,N_5851,N_5843);
and U5921 (N_5921,N_5852,N_5846);
and U5922 (N_5922,N_5802,N_5892);
and U5923 (N_5923,N_5825,N_5837);
nor U5924 (N_5924,N_5807,N_5819);
or U5925 (N_5925,N_5868,N_5800);
nor U5926 (N_5926,N_5850,N_5871);
nor U5927 (N_5927,N_5833,N_5886);
nor U5928 (N_5928,N_5853,N_5826);
and U5929 (N_5929,N_5815,N_5863);
xor U5930 (N_5930,N_5869,N_5896);
or U5931 (N_5931,N_5885,N_5814);
or U5932 (N_5932,N_5804,N_5880);
nor U5933 (N_5933,N_5898,N_5821);
and U5934 (N_5934,N_5831,N_5888);
nor U5935 (N_5935,N_5838,N_5811);
nand U5936 (N_5936,N_5847,N_5842);
and U5937 (N_5937,N_5882,N_5845);
and U5938 (N_5938,N_5848,N_5890);
and U5939 (N_5939,N_5824,N_5897);
xor U5940 (N_5940,N_5872,N_5849);
or U5941 (N_5941,N_5873,N_5895);
nor U5942 (N_5942,N_5860,N_5879);
nor U5943 (N_5943,N_5876,N_5858);
nor U5944 (N_5944,N_5810,N_5840);
or U5945 (N_5945,N_5832,N_5801);
nor U5946 (N_5946,N_5875,N_5865);
nand U5947 (N_5947,N_5891,N_5899);
nand U5948 (N_5948,N_5805,N_5822);
xnor U5949 (N_5949,N_5887,N_5841);
nand U5950 (N_5950,N_5852,N_5899);
nand U5951 (N_5951,N_5846,N_5890);
or U5952 (N_5952,N_5853,N_5846);
nand U5953 (N_5953,N_5839,N_5880);
nor U5954 (N_5954,N_5880,N_5897);
nand U5955 (N_5955,N_5849,N_5851);
nand U5956 (N_5956,N_5881,N_5847);
xnor U5957 (N_5957,N_5863,N_5857);
or U5958 (N_5958,N_5853,N_5856);
nor U5959 (N_5959,N_5818,N_5884);
or U5960 (N_5960,N_5822,N_5821);
nor U5961 (N_5961,N_5851,N_5897);
nand U5962 (N_5962,N_5874,N_5838);
nor U5963 (N_5963,N_5819,N_5832);
nor U5964 (N_5964,N_5888,N_5856);
nand U5965 (N_5965,N_5826,N_5889);
and U5966 (N_5966,N_5859,N_5843);
and U5967 (N_5967,N_5893,N_5898);
nor U5968 (N_5968,N_5871,N_5820);
nor U5969 (N_5969,N_5879,N_5859);
and U5970 (N_5970,N_5819,N_5818);
or U5971 (N_5971,N_5870,N_5843);
and U5972 (N_5972,N_5807,N_5809);
and U5973 (N_5973,N_5868,N_5877);
nor U5974 (N_5974,N_5856,N_5805);
or U5975 (N_5975,N_5858,N_5842);
nand U5976 (N_5976,N_5830,N_5816);
or U5977 (N_5977,N_5850,N_5842);
nand U5978 (N_5978,N_5818,N_5842);
and U5979 (N_5979,N_5853,N_5807);
and U5980 (N_5980,N_5856,N_5891);
nor U5981 (N_5981,N_5818,N_5800);
nand U5982 (N_5982,N_5826,N_5871);
and U5983 (N_5983,N_5837,N_5818);
or U5984 (N_5984,N_5875,N_5891);
and U5985 (N_5985,N_5889,N_5830);
and U5986 (N_5986,N_5866,N_5824);
nor U5987 (N_5987,N_5865,N_5823);
nand U5988 (N_5988,N_5826,N_5825);
and U5989 (N_5989,N_5897,N_5817);
nor U5990 (N_5990,N_5865,N_5877);
or U5991 (N_5991,N_5846,N_5837);
and U5992 (N_5992,N_5895,N_5887);
nor U5993 (N_5993,N_5862,N_5854);
nand U5994 (N_5994,N_5816,N_5896);
nand U5995 (N_5995,N_5809,N_5869);
nand U5996 (N_5996,N_5896,N_5860);
nor U5997 (N_5997,N_5898,N_5823);
nor U5998 (N_5998,N_5810,N_5879);
and U5999 (N_5999,N_5807,N_5801);
nor U6000 (N_6000,N_5945,N_5904);
and U6001 (N_6001,N_5981,N_5973);
and U6002 (N_6002,N_5978,N_5962);
or U6003 (N_6003,N_5928,N_5949);
nor U6004 (N_6004,N_5926,N_5914);
or U6005 (N_6005,N_5985,N_5944);
nor U6006 (N_6006,N_5942,N_5956);
and U6007 (N_6007,N_5916,N_5990);
and U6008 (N_6008,N_5964,N_5900);
nand U6009 (N_6009,N_5902,N_5923);
or U6010 (N_6010,N_5940,N_5908);
and U6011 (N_6011,N_5922,N_5954);
or U6012 (N_6012,N_5984,N_5930);
or U6013 (N_6013,N_5911,N_5957);
nor U6014 (N_6014,N_5971,N_5934);
nor U6015 (N_6015,N_5909,N_5929);
and U6016 (N_6016,N_5991,N_5999);
xor U6017 (N_6017,N_5938,N_5966);
nor U6018 (N_6018,N_5969,N_5913);
or U6019 (N_6019,N_5967,N_5963);
and U6020 (N_6020,N_5952,N_5997);
nor U6021 (N_6021,N_5958,N_5994);
or U6022 (N_6022,N_5974,N_5917);
and U6023 (N_6023,N_5968,N_5987);
nor U6024 (N_6024,N_5931,N_5943);
and U6025 (N_6025,N_5937,N_5983);
nor U6026 (N_6026,N_5959,N_5920);
nor U6027 (N_6027,N_5933,N_5960);
nand U6028 (N_6028,N_5951,N_5992);
or U6029 (N_6029,N_5993,N_5918);
and U6030 (N_6030,N_5905,N_5948);
and U6031 (N_6031,N_5915,N_5979);
nand U6032 (N_6032,N_5972,N_5907);
and U6033 (N_6033,N_5996,N_5976);
or U6034 (N_6034,N_5924,N_5965);
and U6035 (N_6035,N_5947,N_5977);
and U6036 (N_6036,N_5998,N_5939);
and U6037 (N_6037,N_5910,N_5953);
nand U6038 (N_6038,N_5932,N_5989);
and U6039 (N_6039,N_5980,N_5927);
nor U6040 (N_6040,N_5912,N_5925);
xor U6041 (N_6041,N_5970,N_5921);
and U6042 (N_6042,N_5906,N_5982);
nor U6043 (N_6043,N_5901,N_5995);
nor U6044 (N_6044,N_5955,N_5936);
nand U6045 (N_6045,N_5975,N_5946);
nand U6046 (N_6046,N_5950,N_5903);
or U6047 (N_6047,N_5935,N_5986);
nor U6048 (N_6048,N_5988,N_5941);
nand U6049 (N_6049,N_5919,N_5961);
and U6050 (N_6050,N_5940,N_5949);
and U6051 (N_6051,N_5931,N_5946);
nand U6052 (N_6052,N_5998,N_5962);
nor U6053 (N_6053,N_5913,N_5910);
nand U6054 (N_6054,N_5902,N_5922);
or U6055 (N_6055,N_5909,N_5992);
or U6056 (N_6056,N_5953,N_5935);
nor U6057 (N_6057,N_5980,N_5964);
xnor U6058 (N_6058,N_5992,N_5980);
nand U6059 (N_6059,N_5992,N_5907);
and U6060 (N_6060,N_5985,N_5927);
or U6061 (N_6061,N_5909,N_5931);
and U6062 (N_6062,N_5925,N_5983);
nand U6063 (N_6063,N_5989,N_5980);
and U6064 (N_6064,N_5958,N_5956);
and U6065 (N_6065,N_5982,N_5951);
or U6066 (N_6066,N_5901,N_5900);
or U6067 (N_6067,N_5906,N_5931);
nand U6068 (N_6068,N_5911,N_5905);
nor U6069 (N_6069,N_5905,N_5970);
nor U6070 (N_6070,N_5994,N_5998);
nor U6071 (N_6071,N_5987,N_5967);
nor U6072 (N_6072,N_5915,N_5905);
nor U6073 (N_6073,N_5939,N_5935);
nand U6074 (N_6074,N_5950,N_5994);
and U6075 (N_6075,N_5955,N_5986);
nor U6076 (N_6076,N_5909,N_5957);
and U6077 (N_6077,N_5963,N_5988);
and U6078 (N_6078,N_5926,N_5996);
nand U6079 (N_6079,N_5980,N_5919);
or U6080 (N_6080,N_5992,N_5916);
nand U6081 (N_6081,N_5918,N_5916);
and U6082 (N_6082,N_5941,N_5980);
or U6083 (N_6083,N_5920,N_5970);
xor U6084 (N_6084,N_5982,N_5996);
and U6085 (N_6085,N_5916,N_5993);
and U6086 (N_6086,N_5958,N_5963);
or U6087 (N_6087,N_5993,N_5956);
nand U6088 (N_6088,N_5995,N_5967);
and U6089 (N_6089,N_5959,N_5907);
and U6090 (N_6090,N_5920,N_5949);
nand U6091 (N_6091,N_5980,N_5931);
nand U6092 (N_6092,N_5966,N_5956);
and U6093 (N_6093,N_5984,N_5921);
xnor U6094 (N_6094,N_5928,N_5906);
nor U6095 (N_6095,N_5930,N_5988);
and U6096 (N_6096,N_5965,N_5964);
nor U6097 (N_6097,N_5974,N_5998);
and U6098 (N_6098,N_5940,N_5913);
nand U6099 (N_6099,N_5962,N_5972);
or U6100 (N_6100,N_6084,N_6015);
or U6101 (N_6101,N_6079,N_6029);
and U6102 (N_6102,N_6060,N_6051);
nor U6103 (N_6103,N_6038,N_6021);
or U6104 (N_6104,N_6075,N_6032);
or U6105 (N_6105,N_6050,N_6013);
nor U6106 (N_6106,N_6018,N_6000);
and U6107 (N_6107,N_6007,N_6086);
and U6108 (N_6108,N_6031,N_6076);
or U6109 (N_6109,N_6057,N_6061);
nand U6110 (N_6110,N_6054,N_6055);
nor U6111 (N_6111,N_6040,N_6099);
nor U6112 (N_6112,N_6002,N_6011);
or U6113 (N_6113,N_6005,N_6059);
and U6114 (N_6114,N_6098,N_6043);
nor U6115 (N_6115,N_6081,N_6096);
nand U6116 (N_6116,N_6068,N_6049);
xor U6117 (N_6117,N_6080,N_6083);
nand U6118 (N_6118,N_6034,N_6027);
nor U6119 (N_6119,N_6019,N_6062);
or U6120 (N_6120,N_6036,N_6093);
and U6121 (N_6121,N_6078,N_6012);
or U6122 (N_6122,N_6010,N_6016);
nor U6123 (N_6123,N_6046,N_6052);
or U6124 (N_6124,N_6003,N_6094);
and U6125 (N_6125,N_6020,N_6033);
nor U6126 (N_6126,N_6077,N_6071);
or U6127 (N_6127,N_6072,N_6066);
nand U6128 (N_6128,N_6095,N_6047);
nor U6129 (N_6129,N_6025,N_6069);
and U6130 (N_6130,N_6039,N_6091);
and U6131 (N_6131,N_6008,N_6088);
or U6132 (N_6132,N_6085,N_6067);
and U6133 (N_6133,N_6006,N_6053);
nand U6134 (N_6134,N_6063,N_6065);
nand U6135 (N_6135,N_6082,N_6097);
nor U6136 (N_6136,N_6090,N_6014);
and U6137 (N_6137,N_6023,N_6064);
nand U6138 (N_6138,N_6073,N_6037);
and U6139 (N_6139,N_6009,N_6017);
nor U6140 (N_6140,N_6041,N_6074);
nand U6141 (N_6141,N_6056,N_6045);
or U6142 (N_6142,N_6042,N_6028);
nor U6143 (N_6143,N_6026,N_6022);
nor U6144 (N_6144,N_6024,N_6035);
or U6145 (N_6145,N_6070,N_6087);
nor U6146 (N_6146,N_6048,N_6030);
nand U6147 (N_6147,N_6089,N_6092);
or U6148 (N_6148,N_6001,N_6044);
nor U6149 (N_6149,N_6004,N_6058);
and U6150 (N_6150,N_6095,N_6000);
or U6151 (N_6151,N_6006,N_6036);
or U6152 (N_6152,N_6055,N_6061);
and U6153 (N_6153,N_6027,N_6042);
or U6154 (N_6154,N_6000,N_6064);
nor U6155 (N_6155,N_6085,N_6070);
nand U6156 (N_6156,N_6056,N_6058);
and U6157 (N_6157,N_6002,N_6026);
nor U6158 (N_6158,N_6084,N_6011);
and U6159 (N_6159,N_6071,N_6046);
or U6160 (N_6160,N_6019,N_6074);
and U6161 (N_6161,N_6065,N_6025);
nor U6162 (N_6162,N_6024,N_6031);
nor U6163 (N_6163,N_6047,N_6036);
and U6164 (N_6164,N_6006,N_6019);
nand U6165 (N_6165,N_6087,N_6001);
or U6166 (N_6166,N_6074,N_6024);
or U6167 (N_6167,N_6033,N_6011);
nand U6168 (N_6168,N_6010,N_6071);
or U6169 (N_6169,N_6036,N_6077);
or U6170 (N_6170,N_6036,N_6014);
nor U6171 (N_6171,N_6096,N_6044);
or U6172 (N_6172,N_6046,N_6049);
or U6173 (N_6173,N_6000,N_6061);
nor U6174 (N_6174,N_6038,N_6060);
or U6175 (N_6175,N_6024,N_6071);
nand U6176 (N_6176,N_6087,N_6010);
nor U6177 (N_6177,N_6041,N_6023);
nand U6178 (N_6178,N_6049,N_6067);
nor U6179 (N_6179,N_6066,N_6053);
or U6180 (N_6180,N_6098,N_6070);
or U6181 (N_6181,N_6080,N_6042);
and U6182 (N_6182,N_6010,N_6090);
nor U6183 (N_6183,N_6059,N_6054);
nor U6184 (N_6184,N_6041,N_6065);
nand U6185 (N_6185,N_6094,N_6052);
and U6186 (N_6186,N_6097,N_6031);
or U6187 (N_6187,N_6016,N_6096);
or U6188 (N_6188,N_6037,N_6079);
and U6189 (N_6189,N_6071,N_6045);
nor U6190 (N_6190,N_6026,N_6040);
and U6191 (N_6191,N_6007,N_6045);
or U6192 (N_6192,N_6001,N_6089);
nand U6193 (N_6193,N_6092,N_6069);
or U6194 (N_6194,N_6022,N_6048);
or U6195 (N_6195,N_6050,N_6004);
or U6196 (N_6196,N_6059,N_6094);
nor U6197 (N_6197,N_6068,N_6020);
or U6198 (N_6198,N_6021,N_6087);
nand U6199 (N_6199,N_6030,N_6047);
and U6200 (N_6200,N_6170,N_6174);
and U6201 (N_6201,N_6190,N_6119);
nor U6202 (N_6202,N_6124,N_6149);
and U6203 (N_6203,N_6179,N_6144);
and U6204 (N_6204,N_6150,N_6164);
or U6205 (N_6205,N_6192,N_6126);
nor U6206 (N_6206,N_6152,N_6133);
nand U6207 (N_6207,N_6187,N_6109);
and U6208 (N_6208,N_6198,N_6116);
nor U6209 (N_6209,N_6113,N_6110);
and U6210 (N_6210,N_6121,N_6108);
nor U6211 (N_6211,N_6193,N_6196);
nand U6212 (N_6212,N_6194,N_6111);
or U6213 (N_6213,N_6162,N_6145);
nand U6214 (N_6214,N_6186,N_6157);
nand U6215 (N_6215,N_6153,N_6141);
nor U6216 (N_6216,N_6182,N_6171);
nand U6217 (N_6217,N_6167,N_6163);
or U6218 (N_6218,N_6168,N_6103);
and U6219 (N_6219,N_6173,N_6178);
nor U6220 (N_6220,N_6137,N_6105);
nor U6221 (N_6221,N_6134,N_6166);
nand U6222 (N_6222,N_6129,N_6120);
nand U6223 (N_6223,N_6197,N_6132);
and U6224 (N_6224,N_6156,N_6183);
nor U6225 (N_6225,N_6147,N_6158);
nor U6226 (N_6226,N_6101,N_6131);
and U6227 (N_6227,N_6115,N_6180);
or U6228 (N_6228,N_6154,N_6102);
and U6229 (N_6229,N_6161,N_6114);
nand U6230 (N_6230,N_6130,N_6135);
and U6231 (N_6231,N_6155,N_6142);
nand U6232 (N_6232,N_6128,N_6177);
and U6233 (N_6233,N_6112,N_6175);
and U6234 (N_6234,N_6123,N_6148);
nand U6235 (N_6235,N_6176,N_6195);
nor U6236 (N_6236,N_6146,N_6160);
or U6237 (N_6237,N_6181,N_6143);
nor U6238 (N_6238,N_6139,N_6165);
nand U6239 (N_6239,N_6136,N_6191);
and U6240 (N_6240,N_6100,N_6140);
or U6241 (N_6241,N_6159,N_6117);
and U6242 (N_6242,N_6185,N_6169);
or U6243 (N_6243,N_6138,N_6106);
nand U6244 (N_6244,N_6104,N_6118);
and U6245 (N_6245,N_6199,N_6188);
and U6246 (N_6246,N_6127,N_6184);
or U6247 (N_6247,N_6107,N_6189);
nand U6248 (N_6248,N_6122,N_6125);
and U6249 (N_6249,N_6151,N_6172);
nor U6250 (N_6250,N_6127,N_6189);
xnor U6251 (N_6251,N_6138,N_6179);
or U6252 (N_6252,N_6161,N_6159);
nor U6253 (N_6253,N_6156,N_6187);
nand U6254 (N_6254,N_6197,N_6128);
and U6255 (N_6255,N_6145,N_6189);
nor U6256 (N_6256,N_6191,N_6124);
nor U6257 (N_6257,N_6135,N_6128);
and U6258 (N_6258,N_6118,N_6129);
and U6259 (N_6259,N_6168,N_6143);
nand U6260 (N_6260,N_6169,N_6161);
nor U6261 (N_6261,N_6170,N_6141);
or U6262 (N_6262,N_6114,N_6125);
nand U6263 (N_6263,N_6150,N_6131);
nand U6264 (N_6264,N_6163,N_6155);
or U6265 (N_6265,N_6124,N_6140);
xnor U6266 (N_6266,N_6114,N_6199);
nor U6267 (N_6267,N_6179,N_6162);
or U6268 (N_6268,N_6128,N_6149);
or U6269 (N_6269,N_6197,N_6130);
nand U6270 (N_6270,N_6147,N_6129);
nor U6271 (N_6271,N_6127,N_6193);
and U6272 (N_6272,N_6116,N_6114);
nand U6273 (N_6273,N_6100,N_6174);
nand U6274 (N_6274,N_6115,N_6183);
and U6275 (N_6275,N_6154,N_6181);
or U6276 (N_6276,N_6194,N_6199);
nand U6277 (N_6277,N_6106,N_6150);
and U6278 (N_6278,N_6176,N_6168);
and U6279 (N_6279,N_6129,N_6172);
or U6280 (N_6280,N_6139,N_6102);
or U6281 (N_6281,N_6140,N_6179);
or U6282 (N_6282,N_6114,N_6132);
and U6283 (N_6283,N_6180,N_6117);
and U6284 (N_6284,N_6166,N_6173);
nor U6285 (N_6285,N_6156,N_6151);
nor U6286 (N_6286,N_6119,N_6137);
nor U6287 (N_6287,N_6156,N_6166);
and U6288 (N_6288,N_6159,N_6176);
nand U6289 (N_6289,N_6190,N_6184);
nor U6290 (N_6290,N_6134,N_6156);
nand U6291 (N_6291,N_6139,N_6109);
nand U6292 (N_6292,N_6160,N_6199);
nor U6293 (N_6293,N_6176,N_6141);
and U6294 (N_6294,N_6167,N_6186);
nor U6295 (N_6295,N_6125,N_6108);
nand U6296 (N_6296,N_6139,N_6172);
nor U6297 (N_6297,N_6151,N_6108);
nand U6298 (N_6298,N_6168,N_6191);
xnor U6299 (N_6299,N_6126,N_6107);
and U6300 (N_6300,N_6206,N_6269);
nand U6301 (N_6301,N_6231,N_6270);
nor U6302 (N_6302,N_6210,N_6226);
nand U6303 (N_6303,N_6291,N_6295);
nand U6304 (N_6304,N_6222,N_6228);
nand U6305 (N_6305,N_6240,N_6277);
and U6306 (N_6306,N_6225,N_6266);
nand U6307 (N_6307,N_6262,N_6268);
nor U6308 (N_6308,N_6215,N_6282);
and U6309 (N_6309,N_6246,N_6257);
or U6310 (N_6310,N_6209,N_6289);
or U6311 (N_6311,N_6212,N_6217);
nor U6312 (N_6312,N_6208,N_6230);
nand U6313 (N_6313,N_6211,N_6281);
and U6314 (N_6314,N_6216,N_6241);
or U6315 (N_6315,N_6213,N_6293);
nand U6316 (N_6316,N_6292,N_6273);
and U6317 (N_6317,N_6261,N_6214);
nand U6318 (N_6318,N_6258,N_6201);
or U6319 (N_6319,N_6267,N_6233);
nor U6320 (N_6320,N_6204,N_6223);
and U6321 (N_6321,N_6254,N_6252);
nor U6322 (N_6322,N_6232,N_6263);
nor U6323 (N_6323,N_6237,N_6274);
nor U6324 (N_6324,N_6284,N_6294);
or U6325 (N_6325,N_6242,N_6243);
nor U6326 (N_6326,N_6247,N_6288);
nor U6327 (N_6327,N_6219,N_6259);
or U6328 (N_6328,N_6224,N_6283);
and U6329 (N_6329,N_6256,N_6296);
or U6330 (N_6330,N_6265,N_6220);
or U6331 (N_6331,N_6275,N_6264);
nand U6332 (N_6332,N_6290,N_6271);
nand U6333 (N_6333,N_6235,N_6205);
nor U6334 (N_6334,N_6272,N_6221);
nand U6335 (N_6335,N_6245,N_6203);
nor U6336 (N_6336,N_6297,N_6260);
or U6337 (N_6337,N_6279,N_6202);
and U6338 (N_6338,N_6207,N_6248);
nand U6339 (N_6339,N_6286,N_6227);
and U6340 (N_6340,N_6251,N_6238);
xnor U6341 (N_6341,N_6250,N_6299);
and U6342 (N_6342,N_6276,N_6236);
and U6343 (N_6343,N_6287,N_6244);
and U6344 (N_6344,N_6298,N_6255);
or U6345 (N_6345,N_6253,N_6234);
xor U6346 (N_6346,N_6278,N_6200);
or U6347 (N_6347,N_6249,N_6280);
and U6348 (N_6348,N_6218,N_6229);
nand U6349 (N_6349,N_6285,N_6239);
and U6350 (N_6350,N_6206,N_6246);
nand U6351 (N_6351,N_6285,N_6207);
nand U6352 (N_6352,N_6210,N_6289);
nor U6353 (N_6353,N_6204,N_6271);
or U6354 (N_6354,N_6284,N_6282);
nand U6355 (N_6355,N_6246,N_6230);
and U6356 (N_6356,N_6252,N_6226);
and U6357 (N_6357,N_6263,N_6296);
xor U6358 (N_6358,N_6299,N_6212);
and U6359 (N_6359,N_6254,N_6205);
nand U6360 (N_6360,N_6242,N_6281);
or U6361 (N_6361,N_6247,N_6270);
or U6362 (N_6362,N_6279,N_6226);
or U6363 (N_6363,N_6213,N_6206);
or U6364 (N_6364,N_6212,N_6202);
and U6365 (N_6365,N_6293,N_6264);
nand U6366 (N_6366,N_6297,N_6227);
or U6367 (N_6367,N_6284,N_6218);
nand U6368 (N_6368,N_6225,N_6203);
nor U6369 (N_6369,N_6205,N_6259);
nand U6370 (N_6370,N_6237,N_6291);
nand U6371 (N_6371,N_6238,N_6256);
nand U6372 (N_6372,N_6261,N_6209);
or U6373 (N_6373,N_6223,N_6212);
nor U6374 (N_6374,N_6236,N_6210);
nand U6375 (N_6375,N_6269,N_6265);
nand U6376 (N_6376,N_6208,N_6247);
or U6377 (N_6377,N_6230,N_6247);
or U6378 (N_6378,N_6215,N_6294);
nor U6379 (N_6379,N_6222,N_6262);
xnor U6380 (N_6380,N_6277,N_6248);
nor U6381 (N_6381,N_6284,N_6229);
xor U6382 (N_6382,N_6206,N_6293);
or U6383 (N_6383,N_6269,N_6219);
and U6384 (N_6384,N_6221,N_6223);
nor U6385 (N_6385,N_6221,N_6280);
and U6386 (N_6386,N_6246,N_6266);
nand U6387 (N_6387,N_6266,N_6261);
nand U6388 (N_6388,N_6248,N_6274);
and U6389 (N_6389,N_6210,N_6275);
or U6390 (N_6390,N_6280,N_6283);
or U6391 (N_6391,N_6258,N_6243);
and U6392 (N_6392,N_6295,N_6254);
nor U6393 (N_6393,N_6274,N_6250);
and U6394 (N_6394,N_6285,N_6206);
or U6395 (N_6395,N_6221,N_6229);
nor U6396 (N_6396,N_6295,N_6251);
nand U6397 (N_6397,N_6201,N_6244);
nand U6398 (N_6398,N_6240,N_6256);
or U6399 (N_6399,N_6264,N_6291);
and U6400 (N_6400,N_6388,N_6371);
nand U6401 (N_6401,N_6315,N_6393);
nor U6402 (N_6402,N_6320,N_6310);
and U6403 (N_6403,N_6351,N_6394);
nand U6404 (N_6404,N_6342,N_6346);
nand U6405 (N_6405,N_6329,N_6328);
nor U6406 (N_6406,N_6395,N_6331);
and U6407 (N_6407,N_6312,N_6398);
nor U6408 (N_6408,N_6304,N_6349);
and U6409 (N_6409,N_6327,N_6381);
or U6410 (N_6410,N_6372,N_6314);
nor U6411 (N_6411,N_6316,N_6319);
and U6412 (N_6412,N_6309,N_6399);
or U6413 (N_6413,N_6353,N_6308);
or U6414 (N_6414,N_6389,N_6332);
nand U6415 (N_6415,N_6352,N_6369);
or U6416 (N_6416,N_6337,N_6334);
nor U6417 (N_6417,N_6361,N_6326);
or U6418 (N_6418,N_6311,N_6300);
xor U6419 (N_6419,N_6373,N_6366);
nor U6420 (N_6420,N_6339,N_6385);
or U6421 (N_6421,N_6306,N_6362);
and U6422 (N_6422,N_6324,N_6325);
nor U6423 (N_6423,N_6391,N_6365);
nor U6424 (N_6424,N_6379,N_6375);
or U6425 (N_6425,N_6364,N_6344);
nand U6426 (N_6426,N_6397,N_6336);
nand U6427 (N_6427,N_6370,N_6343);
nand U6428 (N_6428,N_6322,N_6358);
nand U6429 (N_6429,N_6387,N_6355);
or U6430 (N_6430,N_6377,N_6390);
or U6431 (N_6431,N_6350,N_6348);
xor U6432 (N_6432,N_6376,N_6357);
and U6433 (N_6433,N_6321,N_6347);
xor U6434 (N_6434,N_6307,N_6305);
or U6435 (N_6435,N_6367,N_6302);
nand U6436 (N_6436,N_6354,N_6386);
or U6437 (N_6437,N_6333,N_6360);
nor U6438 (N_6438,N_6318,N_6356);
nor U6439 (N_6439,N_6374,N_6330);
and U6440 (N_6440,N_6301,N_6335);
or U6441 (N_6441,N_6340,N_6323);
and U6442 (N_6442,N_6396,N_6368);
nor U6443 (N_6443,N_6317,N_6380);
nand U6444 (N_6444,N_6303,N_6383);
or U6445 (N_6445,N_6341,N_6382);
nor U6446 (N_6446,N_6392,N_6378);
or U6447 (N_6447,N_6313,N_6345);
nor U6448 (N_6448,N_6359,N_6363);
or U6449 (N_6449,N_6338,N_6384);
or U6450 (N_6450,N_6309,N_6343);
or U6451 (N_6451,N_6324,N_6331);
nand U6452 (N_6452,N_6385,N_6355);
or U6453 (N_6453,N_6346,N_6354);
nor U6454 (N_6454,N_6363,N_6393);
and U6455 (N_6455,N_6351,N_6313);
nand U6456 (N_6456,N_6385,N_6304);
xor U6457 (N_6457,N_6372,N_6306);
nor U6458 (N_6458,N_6356,N_6368);
or U6459 (N_6459,N_6339,N_6396);
xnor U6460 (N_6460,N_6357,N_6397);
nor U6461 (N_6461,N_6359,N_6382);
nor U6462 (N_6462,N_6356,N_6336);
or U6463 (N_6463,N_6325,N_6306);
and U6464 (N_6464,N_6366,N_6339);
nand U6465 (N_6465,N_6310,N_6318);
nand U6466 (N_6466,N_6332,N_6369);
and U6467 (N_6467,N_6301,N_6384);
or U6468 (N_6468,N_6364,N_6366);
or U6469 (N_6469,N_6349,N_6341);
nand U6470 (N_6470,N_6366,N_6361);
or U6471 (N_6471,N_6343,N_6390);
nor U6472 (N_6472,N_6332,N_6306);
nor U6473 (N_6473,N_6359,N_6332);
and U6474 (N_6474,N_6315,N_6316);
nor U6475 (N_6475,N_6324,N_6385);
or U6476 (N_6476,N_6366,N_6385);
or U6477 (N_6477,N_6342,N_6334);
and U6478 (N_6478,N_6322,N_6304);
and U6479 (N_6479,N_6347,N_6382);
nand U6480 (N_6480,N_6349,N_6351);
nor U6481 (N_6481,N_6364,N_6314);
and U6482 (N_6482,N_6382,N_6370);
nand U6483 (N_6483,N_6354,N_6307);
nor U6484 (N_6484,N_6339,N_6321);
nor U6485 (N_6485,N_6378,N_6384);
nand U6486 (N_6486,N_6311,N_6324);
nand U6487 (N_6487,N_6317,N_6301);
nand U6488 (N_6488,N_6370,N_6339);
nor U6489 (N_6489,N_6355,N_6313);
nand U6490 (N_6490,N_6385,N_6391);
nor U6491 (N_6491,N_6375,N_6394);
and U6492 (N_6492,N_6359,N_6325);
nor U6493 (N_6493,N_6340,N_6382);
nor U6494 (N_6494,N_6390,N_6305);
and U6495 (N_6495,N_6386,N_6312);
nor U6496 (N_6496,N_6308,N_6315);
nand U6497 (N_6497,N_6384,N_6335);
nand U6498 (N_6498,N_6309,N_6330);
nand U6499 (N_6499,N_6375,N_6367);
xnor U6500 (N_6500,N_6410,N_6425);
nor U6501 (N_6501,N_6481,N_6435);
or U6502 (N_6502,N_6486,N_6429);
xnor U6503 (N_6503,N_6427,N_6472);
or U6504 (N_6504,N_6467,N_6406);
or U6505 (N_6505,N_6430,N_6475);
or U6506 (N_6506,N_6454,N_6484);
or U6507 (N_6507,N_6488,N_6468);
or U6508 (N_6508,N_6424,N_6447);
nand U6509 (N_6509,N_6401,N_6449);
and U6510 (N_6510,N_6434,N_6412);
or U6511 (N_6511,N_6411,N_6407);
or U6512 (N_6512,N_6440,N_6498);
nor U6513 (N_6513,N_6493,N_6460);
nor U6514 (N_6514,N_6409,N_6426);
nor U6515 (N_6515,N_6418,N_6497);
and U6516 (N_6516,N_6428,N_6471);
nand U6517 (N_6517,N_6431,N_6451);
nor U6518 (N_6518,N_6495,N_6455);
nor U6519 (N_6519,N_6402,N_6496);
or U6520 (N_6520,N_6469,N_6414);
nor U6521 (N_6521,N_6459,N_6405);
and U6522 (N_6522,N_6444,N_6461);
nand U6523 (N_6523,N_6479,N_6480);
nor U6524 (N_6524,N_6490,N_6437);
nor U6525 (N_6525,N_6417,N_6487);
nand U6526 (N_6526,N_6453,N_6457);
or U6527 (N_6527,N_6420,N_6445);
or U6528 (N_6528,N_6422,N_6491);
or U6529 (N_6529,N_6452,N_6408);
nor U6530 (N_6530,N_6438,N_6466);
and U6531 (N_6531,N_6470,N_6483);
nor U6532 (N_6532,N_6439,N_6450);
and U6533 (N_6533,N_6458,N_6404);
nand U6534 (N_6534,N_6462,N_6477);
nor U6535 (N_6535,N_6416,N_6423);
nand U6536 (N_6536,N_6478,N_6415);
nand U6537 (N_6537,N_6441,N_6456);
or U6538 (N_6538,N_6492,N_6400);
or U6539 (N_6539,N_6465,N_6419);
nor U6540 (N_6540,N_6436,N_6482);
nand U6541 (N_6541,N_6433,N_6485);
or U6542 (N_6542,N_6413,N_6464);
and U6543 (N_6543,N_6448,N_6494);
nor U6544 (N_6544,N_6499,N_6443);
nand U6545 (N_6545,N_6489,N_6442);
nor U6546 (N_6546,N_6463,N_6476);
nand U6547 (N_6547,N_6421,N_6474);
and U6548 (N_6548,N_6473,N_6403);
nand U6549 (N_6549,N_6432,N_6446);
or U6550 (N_6550,N_6419,N_6427);
and U6551 (N_6551,N_6499,N_6452);
and U6552 (N_6552,N_6403,N_6498);
nor U6553 (N_6553,N_6437,N_6478);
nand U6554 (N_6554,N_6402,N_6438);
nand U6555 (N_6555,N_6422,N_6442);
nor U6556 (N_6556,N_6410,N_6402);
or U6557 (N_6557,N_6469,N_6430);
or U6558 (N_6558,N_6428,N_6480);
and U6559 (N_6559,N_6425,N_6439);
nand U6560 (N_6560,N_6487,N_6491);
and U6561 (N_6561,N_6436,N_6430);
and U6562 (N_6562,N_6485,N_6438);
or U6563 (N_6563,N_6403,N_6406);
nor U6564 (N_6564,N_6406,N_6497);
or U6565 (N_6565,N_6461,N_6439);
nor U6566 (N_6566,N_6424,N_6489);
or U6567 (N_6567,N_6471,N_6446);
nor U6568 (N_6568,N_6433,N_6468);
nor U6569 (N_6569,N_6444,N_6424);
and U6570 (N_6570,N_6447,N_6455);
or U6571 (N_6571,N_6428,N_6438);
and U6572 (N_6572,N_6420,N_6489);
nand U6573 (N_6573,N_6430,N_6460);
or U6574 (N_6574,N_6414,N_6463);
and U6575 (N_6575,N_6423,N_6498);
or U6576 (N_6576,N_6409,N_6435);
nor U6577 (N_6577,N_6423,N_6430);
and U6578 (N_6578,N_6423,N_6462);
and U6579 (N_6579,N_6404,N_6444);
nand U6580 (N_6580,N_6485,N_6428);
or U6581 (N_6581,N_6431,N_6463);
nand U6582 (N_6582,N_6475,N_6423);
nor U6583 (N_6583,N_6499,N_6459);
or U6584 (N_6584,N_6420,N_6470);
nand U6585 (N_6585,N_6440,N_6481);
nand U6586 (N_6586,N_6465,N_6450);
nor U6587 (N_6587,N_6465,N_6464);
nor U6588 (N_6588,N_6461,N_6452);
nor U6589 (N_6589,N_6410,N_6443);
nand U6590 (N_6590,N_6425,N_6433);
and U6591 (N_6591,N_6465,N_6413);
nor U6592 (N_6592,N_6483,N_6418);
and U6593 (N_6593,N_6417,N_6418);
and U6594 (N_6594,N_6402,N_6431);
or U6595 (N_6595,N_6469,N_6452);
or U6596 (N_6596,N_6467,N_6437);
nand U6597 (N_6597,N_6468,N_6480);
and U6598 (N_6598,N_6457,N_6447);
and U6599 (N_6599,N_6416,N_6493);
and U6600 (N_6600,N_6569,N_6563);
or U6601 (N_6601,N_6579,N_6582);
nor U6602 (N_6602,N_6517,N_6504);
and U6603 (N_6603,N_6521,N_6585);
or U6604 (N_6604,N_6509,N_6541);
or U6605 (N_6605,N_6540,N_6571);
nand U6606 (N_6606,N_6502,N_6568);
and U6607 (N_6607,N_6512,N_6548);
xnor U6608 (N_6608,N_6599,N_6583);
or U6609 (N_6609,N_6574,N_6515);
xnor U6610 (N_6610,N_6565,N_6566);
xnor U6611 (N_6611,N_6543,N_6501);
and U6612 (N_6612,N_6511,N_6529);
nor U6613 (N_6613,N_6553,N_6518);
or U6614 (N_6614,N_6577,N_6552);
nand U6615 (N_6615,N_6523,N_6576);
nand U6616 (N_6616,N_6537,N_6557);
or U6617 (N_6617,N_6573,N_6575);
or U6618 (N_6618,N_6564,N_6596);
nor U6619 (N_6619,N_6578,N_6527);
and U6620 (N_6620,N_6545,N_6547);
nand U6621 (N_6621,N_6500,N_6567);
and U6622 (N_6622,N_6591,N_6595);
and U6623 (N_6623,N_6589,N_6514);
or U6624 (N_6624,N_6520,N_6590);
or U6625 (N_6625,N_6522,N_6528);
and U6626 (N_6626,N_6594,N_6533);
nor U6627 (N_6627,N_6546,N_6538);
and U6628 (N_6628,N_6516,N_6560);
and U6629 (N_6629,N_6513,N_6572);
and U6630 (N_6630,N_6586,N_6539);
nand U6631 (N_6631,N_6530,N_6580);
and U6632 (N_6632,N_6551,N_6554);
nand U6633 (N_6633,N_6534,N_6561);
xor U6634 (N_6634,N_6556,N_6584);
nor U6635 (N_6635,N_6555,N_6593);
nand U6636 (N_6636,N_6581,N_6503);
or U6637 (N_6637,N_6592,N_6544);
nor U6638 (N_6638,N_6550,N_6597);
or U6639 (N_6639,N_6505,N_6525);
or U6640 (N_6640,N_6562,N_6542);
nor U6641 (N_6641,N_6558,N_6587);
and U6642 (N_6642,N_6536,N_6510);
and U6643 (N_6643,N_6559,N_6519);
and U6644 (N_6644,N_6598,N_6526);
nor U6645 (N_6645,N_6532,N_6531);
nor U6646 (N_6646,N_6524,N_6506);
nor U6647 (N_6647,N_6535,N_6570);
or U6648 (N_6648,N_6508,N_6588);
and U6649 (N_6649,N_6507,N_6549);
and U6650 (N_6650,N_6554,N_6581);
or U6651 (N_6651,N_6545,N_6523);
nand U6652 (N_6652,N_6504,N_6536);
and U6653 (N_6653,N_6552,N_6554);
and U6654 (N_6654,N_6596,N_6580);
nor U6655 (N_6655,N_6521,N_6599);
nor U6656 (N_6656,N_6599,N_6568);
nand U6657 (N_6657,N_6599,N_6580);
or U6658 (N_6658,N_6586,N_6597);
nand U6659 (N_6659,N_6587,N_6535);
nor U6660 (N_6660,N_6517,N_6580);
nor U6661 (N_6661,N_6500,N_6531);
xor U6662 (N_6662,N_6593,N_6502);
nand U6663 (N_6663,N_6586,N_6550);
nand U6664 (N_6664,N_6550,N_6551);
and U6665 (N_6665,N_6599,N_6535);
nor U6666 (N_6666,N_6534,N_6506);
and U6667 (N_6667,N_6523,N_6505);
nor U6668 (N_6668,N_6538,N_6560);
and U6669 (N_6669,N_6502,N_6569);
and U6670 (N_6670,N_6523,N_6543);
and U6671 (N_6671,N_6542,N_6530);
or U6672 (N_6672,N_6516,N_6549);
nand U6673 (N_6673,N_6566,N_6536);
nor U6674 (N_6674,N_6502,N_6595);
nand U6675 (N_6675,N_6558,N_6512);
or U6676 (N_6676,N_6542,N_6521);
xor U6677 (N_6677,N_6570,N_6599);
nand U6678 (N_6678,N_6592,N_6506);
nand U6679 (N_6679,N_6565,N_6531);
and U6680 (N_6680,N_6566,N_6520);
nand U6681 (N_6681,N_6556,N_6598);
or U6682 (N_6682,N_6564,N_6563);
nand U6683 (N_6683,N_6536,N_6543);
nor U6684 (N_6684,N_6559,N_6500);
or U6685 (N_6685,N_6528,N_6541);
nand U6686 (N_6686,N_6591,N_6572);
nor U6687 (N_6687,N_6500,N_6514);
or U6688 (N_6688,N_6536,N_6593);
nor U6689 (N_6689,N_6532,N_6593);
nand U6690 (N_6690,N_6580,N_6561);
nor U6691 (N_6691,N_6567,N_6597);
nor U6692 (N_6692,N_6505,N_6582);
nor U6693 (N_6693,N_6518,N_6543);
and U6694 (N_6694,N_6503,N_6591);
nand U6695 (N_6695,N_6543,N_6540);
nor U6696 (N_6696,N_6586,N_6521);
nor U6697 (N_6697,N_6533,N_6531);
xor U6698 (N_6698,N_6597,N_6587);
nor U6699 (N_6699,N_6500,N_6590);
nand U6700 (N_6700,N_6607,N_6602);
and U6701 (N_6701,N_6613,N_6600);
nor U6702 (N_6702,N_6687,N_6625);
nand U6703 (N_6703,N_6666,N_6608);
nor U6704 (N_6704,N_6655,N_6648);
nor U6705 (N_6705,N_6684,N_6699);
nand U6706 (N_6706,N_6642,N_6689);
or U6707 (N_6707,N_6672,N_6665);
nand U6708 (N_6708,N_6634,N_6616);
nor U6709 (N_6709,N_6670,N_6653);
and U6710 (N_6710,N_6627,N_6603);
nand U6711 (N_6711,N_6685,N_6614);
nor U6712 (N_6712,N_6694,N_6698);
nand U6713 (N_6713,N_6606,N_6645);
or U6714 (N_6714,N_6695,N_6667);
or U6715 (N_6715,N_6674,N_6641);
or U6716 (N_6716,N_6662,N_6619);
xnor U6717 (N_6717,N_6649,N_6656);
and U6718 (N_6718,N_6664,N_6673);
or U6719 (N_6719,N_6654,N_6647);
nand U6720 (N_6720,N_6679,N_6660);
or U6721 (N_6721,N_6651,N_6636);
and U6722 (N_6722,N_6693,N_6610);
xnor U6723 (N_6723,N_6611,N_6630);
and U6724 (N_6724,N_6609,N_6601);
nor U6725 (N_6725,N_6640,N_6697);
or U6726 (N_6726,N_6663,N_6618);
and U6727 (N_6727,N_6632,N_6623);
and U6728 (N_6728,N_6643,N_6646);
or U6729 (N_6729,N_6678,N_6624);
or U6730 (N_6730,N_6621,N_6604);
nor U6731 (N_6731,N_6657,N_6605);
and U6732 (N_6732,N_6676,N_6675);
or U6733 (N_6733,N_6637,N_6682);
and U6734 (N_6734,N_6671,N_6677);
nand U6735 (N_6735,N_6681,N_6617);
nand U6736 (N_6736,N_6691,N_6668);
nand U6737 (N_6737,N_6612,N_6652);
xor U6738 (N_6738,N_6661,N_6631);
and U6739 (N_6739,N_6620,N_6622);
or U6740 (N_6740,N_6659,N_6690);
nor U6741 (N_6741,N_6639,N_6658);
or U6742 (N_6742,N_6669,N_6680);
or U6743 (N_6743,N_6686,N_6644);
nor U6744 (N_6744,N_6628,N_6626);
and U6745 (N_6745,N_6692,N_6635);
or U6746 (N_6746,N_6638,N_6696);
or U6747 (N_6747,N_6615,N_6650);
nor U6748 (N_6748,N_6688,N_6683);
nand U6749 (N_6749,N_6629,N_6633);
and U6750 (N_6750,N_6684,N_6673);
nand U6751 (N_6751,N_6620,N_6659);
or U6752 (N_6752,N_6614,N_6695);
or U6753 (N_6753,N_6620,N_6666);
and U6754 (N_6754,N_6636,N_6609);
nor U6755 (N_6755,N_6651,N_6606);
nor U6756 (N_6756,N_6607,N_6681);
and U6757 (N_6757,N_6679,N_6688);
or U6758 (N_6758,N_6634,N_6662);
and U6759 (N_6759,N_6642,N_6603);
nand U6760 (N_6760,N_6677,N_6618);
and U6761 (N_6761,N_6604,N_6661);
or U6762 (N_6762,N_6669,N_6678);
or U6763 (N_6763,N_6633,N_6636);
and U6764 (N_6764,N_6639,N_6621);
nand U6765 (N_6765,N_6659,N_6671);
and U6766 (N_6766,N_6684,N_6650);
nand U6767 (N_6767,N_6623,N_6603);
or U6768 (N_6768,N_6671,N_6680);
and U6769 (N_6769,N_6600,N_6629);
nand U6770 (N_6770,N_6686,N_6660);
xor U6771 (N_6771,N_6642,N_6660);
or U6772 (N_6772,N_6671,N_6683);
xor U6773 (N_6773,N_6650,N_6606);
nand U6774 (N_6774,N_6696,N_6614);
or U6775 (N_6775,N_6665,N_6682);
nor U6776 (N_6776,N_6663,N_6696);
and U6777 (N_6777,N_6692,N_6647);
nand U6778 (N_6778,N_6615,N_6619);
and U6779 (N_6779,N_6643,N_6627);
xnor U6780 (N_6780,N_6603,N_6641);
and U6781 (N_6781,N_6619,N_6625);
and U6782 (N_6782,N_6655,N_6632);
nand U6783 (N_6783,N_6610,N_6640);
and U6784 (N_6784,N_6656,N_6652);
nor U6785 (N_6785,N_6696,N_6643);
nor U6786 (N_6786,N_6658,N_6642);
and U6787 (N_6787,N_6605,N_6667);
nor U6788 (N_6788,N_6615,N_6608);
nor U6789 (N_6789,N_6614,N_6624);
and U6790 (N_6790,N_6651,N_6653);
and U6791 (N_6791,N_6689,N_6651);
nand U6792 (N_6792,N_6606,N_6661);
or U6793 (N_6793,N_6660,N_6676);
or U6794 (N_6794,N_6688,N_6685);
nor U6795 (N_6795,N_6693,N_6682);
nor U6796 (N_6796,N_6695,N_6607);
and U6797 (N_6797,N_6643,N_6677);
and U6798 (N_6798,N_6612,N_6654);
xor U6799 (N_6799,N_6630,N_6672);
nand U6800 (N_6800,N_6726,N_6741);
or U6801 (N_6801,N_6734,N_6754);
and U6802 (N_6802,N_6700,N_6718);
xnor U6803 (N_6803,N_6765,N_6783);
or U6804 (N_6804,N_6715,N_6757);
and U6805 (N_6805,N_6736,N_6753);
nand U6806 (N_6806,N_6787,N_6772);
or U6807 (N_6807,N_6740,N_6723);
nand U6808 (N_6808,N_6775,N_6746);
nor U6809 (N_6809,N_6792,N_6789);
nor U6810 (N_6810,N_6763,N_6760);
nor U6811 (N_6811,N_6719,N_6724);
nand U6812 (N_6812,N_6786,N_6797);
or U6813 (N_6813,N_6785,N_6749);
or U6814 (N_6814,N_6793,N_6705);
nand U6815 (N_6815,N_6766,N_6742);
or U6816 (N_6816,N_6764,N_6791);
and U6817 (N_6817,N_6717,N_6762);
nand U6818 (N_6818,N_6771,N_6761);
or U6819 (N_6819,N_6767,N_6790);
and U6820 (N_6820,N_6779,N_6710);
nor U6821 (N_6821,N_6768,N_6777);
or U6822 (N_6822,N_6725,N_6769);
or U6823 (N_6823,N_6732,N_6704);
or U6824 (N_6824,N_6773,N_6751);
nand U6825 (N_6825,N_6702,N_6713);
nor U6826 (N_6826,N_6730,N_6712);
xnor U6827 (N_6827,N_6796,N_6747);
nand U6828 (N_6828,N_6728,N_6759);
nor U6829 (N_6829,N_6714,N_6756);
and U6830 (N_6830,N_6798,N_6706);
and U6831 (N_6831,N_6794,N_6745);
nand U6832 (N_6832,N_6774,N_6770);
nor U6833 (N_6833,N_6758,N_6752);
nand U6834 (N_6834,N_6729,N_6716);
nand U6835 (N_6835,N_6750,N_6707);
nand U6836 (N_6836,N_6711,N_6776);
or U6837 (N_6837,N_6755,N_6737);
and U6838 (N_6838,N_6743,N_6784);
or U6839 (N_6839,N_6781,N_6739);
nand U6840 (N_6840,N_6782,N_6795);
or U6841 (N_6841,N_6738,N_6748);
nor U6842 (N_6842,N_6722,N_6744);
nand U6843 (N_6843,N_6780,N_6735);
nor U6844 (N_6844,N_6720,N_6731);
nor U6845 (N_6845,N_6799,N_6709);
nand U6846 (N_6846,N_6721,N_6708);
and U6847 (N_6847,N_6778,N_6733);
or U6848 (N_6848,N_6703,N_6701);
nand U6849 (N_6849,N_6727,N_6788);
nand U6850 (N_6850,N_6774,N_6799);
nand U6851 (N_6851,N_6791,N_6705);
and U6852 (N_6852,N_6759,N_6712);
or U6853 (N_6853,N_6746,N_6737);
and U6854 (N_6854,N_6748,N_6784);
nor U6855 (N_6855,N_6742,N_6784);
and U6856 (N_6856,N_6749,N_6717);
nand U6857 (N_6857,N_6736,N_6727);
nor U6858 (N_6858,N_6789,N_6771);
and U6859 (N_6859,N_6722,N_6700);
nand U6860 (N_6860,N_6704,N_6710);
nor U6861 (N_6861,N_6783,N_6779);
nand U6862 (N_6862,N_6771,N_6744);
nand U6863 (N_6863,N_6779,N_6752);
nor U6864 (N_6864,N_6709,N_6737);
or U6865 (N_6865,N_6747,N_6716);
and U6866 (N_6866,N_6786,N_6766);
nand U6867 (N_6867,N_6736,N_6718);
nand U6868 (N_6868,N_6756,N_6713);
nor U6869 (N_6869,N_6703,N_6708);
and U6870 (N_6870,N_6749,N_6783);
nand U6871 (N_6871,N_6739,N_6708);
and U6872 (N_6872,N_6704,N_6780);
or U6873 (N_6873,N_6734,N_6751);
nand U6874 (N_6874,N_6780,N_6737);
and U6875 (N_6875,N_6768,N_6798);
or U6876 (N_6876,N_6796,N_6784);
nor U6877 (N_6877,N_6726,N_6769);
nor U6878 (N_6878,N_6782,N_6731);
and U6879 (N_6879,N_6775,N_6728);
nor U6880 (N_6880,N_6714,N_6748);
or U6881 (N_6881,N_6759,N_6705);
xor U6882 (N_6882,N_6702,N_6743);
and U6883 (N_6883,N_6750,N_6757);
and U6884 (N_6884,N_6722,N_6729);
xnor U6885 (N_6885,N_6744,N_6776);
or U6886 (N_6886,N_6700,N_6721);
and U6887 (N_6887,N_6788,N_6794);
nor U6888 (N_6888,N_6722,N_6749);
nand U6889 (N_6889,N_6701,N_6749);
nand U6890 (N_6890,N_6702,N_6751);
nand U6891 (N_6891,N_6725,N_6793);
and U6892 (N_6892,N_6737,N_6750);
nor U6893 (N_6893,N_6742,N_6765);
nand U6894 (N_6894,N_6700,N_6758);
and U6895 (N_6895,N_6749,N_6792);
nor U6896 (N_6896,N_6719,N_6756);
nand U6897 (N_6897,N_6717,N_6791);
xor U6898 (N_6898,N_6706,N_6720);
and U6899 (N_6899,N_6709,N_6739);
nor U6900 (N_6900,N_6809,N_6839);
xnor U6901 (N_6901,N_6866,N_6870);
and U6902 (N_6902,N_6878,N_6880);
nand U6903 (N_6903,N_6823,N_6825);
or U6904 (N_6904,N_6837,N_6844);
or U6905 (N_6905,N_6861,N_6896);
and U6906 (N_6906,N_6800,N_6852);
nor U6907 (N_6907,N_6891,N_6897);
or U6908 (N_6908,N_6864,N_6846);
nand U6909 (N_6909,N_6831,N_6835);
or U6910 (N_6910,N_6860,N_6848);
and U6911 (N_6911,N_6819,N_6805);
and U6912 (N_6912,N_6893,N_6817);
xor U6913 (N_6913,N_6890,N_6879);
and U6914 (N_6914,N_6851,N_6874);
or U6915 (N_6915,N_6873,N_6838);
nor U6916 (N_6916,N_6826,N_6820);
or U6917 (N_6917,N_6898,N_6857);
or U6918 (N_6918,N_6806,N_6840);
or U6919 (N_6919,N_6843,N_6853);
or U6920 (N_6920,N_6884,N_6824);
or U6921 (N_6921,N_6892,N_6849);
or U6922 (N_6922,N_6810,N_6854);
and U6923 (N_6923,N_6859,N_6808);
nand U6924 (N_6924,N_6876,N_6801);
nand U6925 (N_6925,N_6829,N_6822);
nor U6926 (N_6926,N_6877,N_6813);
nand U6927 (N_6927,N_6804,N_6803);
or U6928 (N_6928,N_6887,N_6899);
nor U6929 (N_6929,N_6847,N_6871);
or U6930 (N_6930,N_6882,N_6885);
and U6931 (N_6931,N_6888,N_6842);
nand U6932 (N_6932,N_6895,N_6812);
nand U6933 (N_6933,N_6836,N_6865);
or U6934 (N_6934,N_6832,N_6889);
and U6935 (N_6935,N_6833,N_6856);
nand U6936 (N_6936,N_6894,N_6845);
or U6937 (N_6937,N_6834,N_6811);
nand U6938 (N_6938,N_6875,N_6862);
nor U6939 (N_6939,N_6886,N_6841);
or U6940 (N_6940,N_6815,N_6818);
and U6941 (N_6941,N_6863,N_6802);
nand U6942 (N_6942,N_6828,N_6850);
nor U6943 (N_6943,N_6821,N_6827);
nor U6944 (N_6944,N_6814,N_6869);
or U6945 (N_6945,N_6807,N_6868);
or U6946 (N_6946,N_6858,N_6830);
nor U6947 (N_6947,N_6867,N_6855);
nor U6948 (N_6948,N_6881,N_6872);
or U6949 (N_6949,N_6816,N_6883);
or U6950 (N_6950,N_6844,N_6892);
and U6951 (N_6951,N_6839,N_6890);
nand U6952 (N_6952,N_6881,N_6867);
or U6953 (N_6953,N_6867,N_6826);
nand U6954 (N_6954,N_6896,N_6801);
nand U6955 (N_6955,N_6806,N_6837);
nand U6956 (N_6956,N_6840,N_6891);
nand U6957 (N_6957,N_6845,N_6851);
and U6958 (N_6958,N_6834,N_6823);
nand U6959 (N_6959,N_6857,N_6870);
and U6960 (N_6960,N_6847,N_6822);
or U6961 (N_6961,N_6843,N_6811);
nand U6962 (N_6962,N_6844,N_6896);
nand U6963 (N_6963,N_6883,N_6811);
xor U6964 (N_6964,N_6890,N_6817);
and U6965 (N_6965,N_6828,N_6806);
and U6966 (N_6966,N_6880,N_6825);
and U6967 (N_6967,N_6827,N_6862);
or U6968 (N_6968,N_6850,N_6884);
or U6969 (N_6969,N_6828,N_6846);
and U6970 (N_6970,N_6830,N_6823);
or U6971 (N_6971,N_6820,N_6872);
and U6972 (N_6972,N_6897,N_6877);
or U6973 (N_6973,N_6834,N_6802);
nor U6974 (N_6974,N_6806,N_6864);
nor U6975 (N_6975,N_6859,N_6890);
nand U6976 (N_6976,N_6881,N_6866);
and U6977 (N_6977,N_6813,N_6865);
nand U6978 (N_6978,N_6819,N_6893);
or U6979 (N_6979,N_6899,N_6808);
or U6980 (N_6980,N_6839,N_6881);
nand U6981 (N_6981,N_6830,N_6846);
nand U6982 (N_6982,N_6883,N_6823);
or U6983 (N_6983,N_6846,N_6845);
and U6984 (N_6984,N_6808,N_6847);
or U6985 (N_6985,N_6875,N_6863);
nor U6986 (N_6986,N_6899,N_6879);
nor U6987 (N_6987,N_6801,N_6808);
or U6988 (N_6988,N_6895,N_6837);
nand U6989 (N_6989,N_6807,N_6840);
and U6990 (N_6990,N_6893,N_6875);
and U6991 (N_6991,N_6839,N_6870);
nand U6992 (N_6992,N_6882,N_6866);
and U6993 (N_6993,N_6819,N_6848);
or U6994 (N_6994,N_6812,N_6833);
nor U6995 (N_6995,N_6858,N_6831);
nand U6996 (N_6996,N_6892,N_6874);
or U6997 (N_6997,N_6818,N_6838);
xor U6998 (N_6998,N_6825,N_6856);
nand U6999 (N_6999,N_6888,N_6848);
nor U7000 (N_7000,N_6973,N_6961);
nor U7001 (N_7001,N_6907,N_6993);
nor U7002 (N_7002,N_6969,N_6918);
and U7003 (N_7003,N_6930,N_6950);
and U7004 (N_7004,N_6999,N_6921);
nand U7005 (N_7005,N_6992,N_6932);
and U7006 (N_7006,N_6946,N_6922);
nor U7007 (N_7007,N_6958,N_6957);
and U7008 (N_7008,N_6994,N_6929);
nand U7009 (N_7009,N_6963,N_6997);
or U7010 (N_7010,N_6986,N_6980);
or U7011 (N_7011,N_6928,N_6967);
nor U7012 (N_7012,N_6987,N_6971);
nor U7013 (N_7013,N_6923,N_6966);
nor U7014 (N_7014,N_6903,N_6960);
and U7015 (N_7015,N_6955,N_6925);
and U7016 (N_7016,N_6968,N_6952);
and U7017 (N_7017,N_6924,N_6965);
and U7018 (N_7018,N_6991,N_6976);
or U7019 (N_7019,N_6954,N_6981);
nand U7020 (N_7020,N_6998,N_6972);
nand U7021 (N_7021,N_6945,N_6990);
nor U7022 (N_7022,N_6975,N_6905);
nand U7023 (N_7023,N_6989,N_6917);
and U7024 (N_7024,N_6953,N_6939);
nor U7025 (N_7025,N_6926,N_6943);
xnor U7026 (N_7026,N_6977,N_6906);
or U7027 (N_7027,N_6974,N_6916);
or U7028 (N_7028,N_6948,N_6910);
or U7029 (N_7029,N_6941,N_6913);
nor U7030 (N_7030,N_6951,N_6988);
and U7031 (N_7031,N_6900,N_6931);
nor U7032 (N_7032,N_6911,N_6949);
and U7033 (N_7033,N_6933,N_6944);
or U7034 (N_7034,N_6914,N_6984);
or U7035 (N_7035,N_6962,N_6959);
and U7036 (N_7036,N_6985,N_6964);
and U7037 (N_7037,N_6970,N_6979);
or U7038 (N_7038,N_6908,N_6982);
or U7039 (N_7039,N_6936,N_6956);
nor U7040 (N_7040,N_6934,N_6942);
nor U7041 (N_7041,N_6912,N_6947);
and U7042 (N_7042,N_6909,N_6902);
nor U7043 (N_7043,N_6937,N_6927);
or U7044 (N_7044,N_6996,N_6919);
xor U7045 (N_7045,N_6978,N_6983);
and U7046 (N_7046,N_6915,N_6901);
and U7047 (N_7047,N_6995,N_6920);
and U7048 (N_7048,N_6938,N_6935);
or U7049 (N_7049,N_6904,N_6940);
nor U7050 (N_7050,N_6907,N_6966);
and U7051 (N_7051,N_6902,N_6924);
or U7052 (N_7052,N_6983,N_6911);
nor U7053 (N_7053,N_6958,N_6997);
and U7054 (N_7054,N_6931,N_6933);
and U7055 (N_7055,N_6940,N_6906);
and U7056 (N_7056,N_6982,N_6936);
and U7057 (N_7057,N_6952,N_6905);
or U7058 (N_7058,N_6966,N_6928);
and U7059 (N_7059,N_6952,N_6972);
or U7060 (N_7060,N_6942,N_6945);
nand U7061 (N_7061,N_6925,N_6967);
nand U7062 (N_7062,N_6907,N_6995);
xnor U7063 (N_7063,N_6919,N_6990);
and U7064 (N_7064,N_6987,N_6940);
and U7065 (N_7065,N_6905,N_6995);
nor U7066 (N_7066,N_6946,N_6960);
nor U7067 (N_7067,N_6900,N_6925);
nand U7068 (N_7068,N_6912,N_6995);
and U7069 (N_7069,N_6979,N_6901);
or U7070 (N_7070,N_6917,N_6933);
xnor U7071 (N_7071,N_6906,N_6950);
xnor U7072 (N_7072,N_6906,N_6958);
xor U7073 (N_7073,N_6980,N_6966);
or U7074 (N_7074,N_6948,N_6972);
and U7075 (N_7075,N_6962,N_6997);
nand U7076 (N_7076,N_6935,N_6912);
and U7077 (N_7077,N_6957,N_6908);
nor U7078 (N_7078,N_6993,N_6917);
xor U7079 (N_7079,N_6978,N_6935);
xor U7080 (N_7080,N_6932,N_6940);
and U7081 (N_7081,N_6964,N_6942);
nor U7082 (N_7082,N_6957,N_6931);
nand U7083 (N_7083,N_6943,N_6972);
nand U7084 (N_7084,N_6978,N_6946);
and U7085 (N_7085,N_6940,N_6963);
or U7086 (N_7086,N_6989,N_6901);
nand U7087 (N_7087,N_6927,N_6919);
and U7088 (N_7088,N_6902,N_6916);
or U7089 (N_7089,N_6986,N_6921);
or U7090 (N_7090,N_6975,N_6974);
or U7091 (N_7091,N_6994,N_6961);
nand U7092 (N_7092,N_6922,N_6909);
nor U7093 (N_7093,N_6929,N_6971);
nand U7094 (N_7094,N_6954,N_6959);
or U7095 (N_7095,N_6985,N_6918);
xnor U7096 (N_7096,N_6928,N_6910);
or U7097 (N_7097,N_6926,N_6936);
nand U7098 (N_7098,N_6962,N_6976);
nor U7099 (N_7099,N_6988,N_6933);
nor U7100 (N_7100,N_7074,N_7078);
and U7101 (N_7101,N_7055,N_7023);
and U7102 (N_7102,N_7026,N_7084);
and U7103 (N_7103,N_7041,N_7021);
nand U7104 (N_7104,N_7000,N_7099);
nand U7105 (N_7105,N_7058,N_7088);
nor U7106 (N_7106,N_7095,N_7009);
and U7107 (N_7107,N_7012,N_7077);
nand U7108 (N_7108,N_7073,N_7025);
or U7109 (N_7109,N_7090,N_7039);
nor U7110 (N_7110,N_7019,N_7079);
nand U7111 (N_7111,N_7043,N_7014);
nand U7112 (N_7112,N_7052,N_7002);
and U7113 (N_7113,N_7049,N_7071);
and U7114 (N_7114,N_7020,N_7046);
and U7115 (N_7115,N_7072,N_7034);
or U7116 (N_7116,N_7007,N_7094);
nor U7117 (N_7117,N_7017,N_7011);
and U7118 (N_7118,N_7008,N_7086);
or U7119 (N_7119,N_7044,N_7063);
and U7120 (N_7120,N_7013,N_7054);
and U7121 (N_7121,N_7018,N_7062);
nand U7122 (N_7122,N_7075,N_7010);
and U7123 (N_7123,N_7089,N_7040);
nand U7124 (N_7124,N_7001,N_7061);
and U7125 (N_7125,N_7057,N_7045);
or U7126 (N_7126,N_7065,N_7087);
nor U7127 (N_7127,N_7081,N_7024);
nand U7128 (N_7128,N_7083,N_7027);
or U7129 (N_7129,N_7029,N_7037);
nand U7130 (N_7130,N_7035,N_7036);
and U7131 (N_7131,N_7031,N_7097);
or U7132 (N_7132,N_7033,N_7048);
and U7133 (N_7133,N_7006,N_7082);
nand U7134 (N_7134,N_7070,N_7051);
and U7135 (N_7135,N_7047,N_7004);
nor U7136 (N_7136,N_7053,N_7060);
nand U7137 (N_7137,N_7080,N_7098);
and U7138 (N_7138,N_7038,N_7022);
or U7139 (N_7139,N_7093,N_7092);
nor U7140 (N_7140,N_7032,N_7003);
nand U7141 (N_7141,N_7068,N_7067);
or U7142 (N_7142,N_7030,N_7028);
nand U7143 (N_7143,N_7096,N_7059);
or U7144 (N_7144,N_7050,N_7076);
and U7145 (N_7145,N_7005,N_7085);
and U7146 (N_7146,N_7042,N_7066);
nor U7147 (N_7147,N_7069,N_7064);
or U7148 (N_7148,N_7016,N_7056);
nand U7149 (N_7149,N_7015,N_7091);
nand U7150 (N_7150,N_7026,N_7029);
or U7151 (N_7151,N_7096,N_7053);
and U7152 (N_7152,N_7012,N_7049);
or U7153 (N_7153,N_7018,N_7007);
nor U7154 (N_7154,N_7067,N_7089);
nor U7155 (N_7155,N_7043,N_7045);
nor U7156 (N_7156,N_7017,N_7094);
nand U7157 (N_7157,N_7073,N_7007);
nor U7158 (N_7158,N_7062,N_7029);
nand U7159 (N_7159,N_7015,N_7071);
nor U7160 (N_7160,N_7008,N_7029);
nand U7161 (N_7161,N_7014,N_7083);
nor U7162 (N_7162,N_7044,N_7004);
nand U7163 (N_7163,N_7000,N_7045);
or U7164 (N_7164,N_7072,N_7042);
nand U7165 (N_7165,N_7037,N_7011);
or U7166 (N_7166,N_7026,N_7054);
and U7167 (N_7167,N_7091,N_7050);
nand U7168 (N_7168,N_7039,N_7036);
and U7169 (N_7169,N_7055,N_7080);
nand U7170 (N_7170,N_7076,N_7082);
nand U7171 (N_7171,N_7084,N_7078);
nand U7172 (N_7172,N_7002,N_7033);
or U7173 (N_7173,N_7064,N_7077);
nor U7174 (N_7174,N_7008,N_7076);
nor U7175 (N_7175,N_7035,N_7044);
and U7176 (N_7176,N_7026,N_7095);
nand U7177 (N_7177,N_7061,N_7040);
nand U7178 (N_7178,N_7098,N_7001);
nor U7179 (N_7179,N_7074,N_7059);
nand U7180 (N_7180,N_7008,N_7090);
and U7181 (N_7181,N_7018,N_7024);
nand U7182 (N_7182,N_7086,N_7015);
and U7183 (N_7183,N_7078,N_7002);
nor U7184 (N_7184,N_7093,N_7003);
and U7185 (N_7185,N_7086,N_7052);
or U7186 (N_7186,N_7054,N_7059);
or U7187 (N_7187,N_7031,N_7074);
and U7188 (N_7188,N_7037,N_7010);
nand U7189 (N_7189,N_7078,N_7053);
or U7190 (N_7190,N_7071,N_7003);
nor U7191 (N_7191,N_7054,N_7032);
nor U7192 (N_7192,N_7009,N_7024);
and U7193 (N_7193,N_7000,N_7071);
nor U7194 (N_7194,N_7070,N_7048);
and U7195 (N_7195,N_7062,N_7073);
nor U7196 (N_7196,N_7036,N_7021);
nor U7197 (N_7197,N_7048,N_7078);
and U7198 (N_7198,N_7034,N_7028);
or U7199 (N_7199,N_7095,N_7003);
and U7200 (N_7200,N_7183,N_7180);
or U7201 (N_7201,N_7169,N_7152);
or U7202 (N_7202,N_7155,N_7161);
nor U7203 (N_7203,N_7191,N_7194);
or U7204 (N_7204,N_7168,N_7144);
and U7205 (N_7205,N_7113,N_7189);
and U7206 (N_7206,N_7198,N_7172);
or U7207 (N_7207,N_7125,N_7186);
nand U7208 (N_7208,N_7137,N_7139);
nand U7209 (N_7209,N_7112,N_7181);
or U7210 (N_7210,N_7164,N_7149);
xnor U7211 (N_7211,N_7146,N_7178);
nand U7212 (N_7212,N_7167,N_7123);
or U7213 (N_7213,N_7156,N_7175);
nor U7214 (N_7214,N_7143,N_7153);
and U7215 (N_7215,N_7114,N_7159);
and U7216 (N_7216,N_7130,N_7134);
nor U7217 (N_7217,N_7106,N_7118);
or U7218 (N_7218,N_7195,N_7188);
and U7219 (N_7219,N_7111,N_7136);
or U7220 (N_7220,N_7101,N_7122);
and U7221 (N_7221,N_7109,N_7197);
nor U7222 (N_7222,N_7133,N_7174);
and U7223 (N_7223,N_7105,N_7115);
nor U7224 (N_7224,N_7128,N_7102);
or U7225 (N_7225,N_7163,N_7100);
nand U7226 (N_7226,N_7170,N_7150);
nand U7227 (N_7227,N_7185,N_7148);
nand U7228 (N_7228,N_7179,N_7132);
xnor U7229 (N_7229,N_7187,N_7196);
nand U7230 (N_7230,N_7147,N_7135);
nor U7231 (N_7231,N_7199,N_7154);
nand U7232 (N_7232,N_7117,N_7110);
nor U7233 (N_7233,N_7107,N_7177);
nor U7234 (N_7234,N_7124,N_7121);
nand U7235 (N_7235,N_7141,N_7165);
or U7236 (N_7236,N_7127,N_7157);
or U7237 (N_7237,N_7119,N_7126);
nor U7238 (N_7238,N_7142,N_7176);
nand U7239 (N_7239,N_7162,N_7192);
or U7240 (N_7240,N_7140,N_7151);
and U7241 (N_7241,N_7145,N_7193);
or U7242 (N_7242,N_7160,N_7120);
nor U7243 (N_7243,N_7158,N_7103);
nor U7244 (N_7244,N_7131,N_7182);
or U7245 (N_7245,N_7190,N_7129);
and U7246 (N_7246,N_7184,N_7116);
and U7247 (N_7247,N_7104,N_7171);
nor U7248 (N_7248,N_7108,N_7166);
nor U7249 (N_7249,N_7173,N_7138);
nand U7250 (N_7250,N_7136,N_7163);
and U7251 (N_7251,N_7175,N_7108);
xnor U7252 (N_7252,N_7151,N_7191);
nand U7253 (N_7253,N_7141,N_7191);
or U7254 (N_7254,N_7197,N_7178);
or U7255 (N_7255,N_7174,N_7179);
nor U7256 (N_7256,N_7155,N_7126);
nand U7257 (N_7257,N_7172,N_7195);
and U7258 (N_7258,N_7183,N_7157);
and U7259 (N_7259,N_7102,N_7151);
or U7260 (N_7260,N_7172,N_7124);
nor U7261 (N_7261,N_7122,N_7109);
and U7262 (N_7262,N_7111,N_7158);
and U7263 (N_7263,N_7189,N_7158);
and U7264 (N_7264,N_7156,N_7193);
nand U7265 (N_7265,N_7165,N_7183);
and U7266 (N_7266,N_7101,N_7125);
nand U7267 (N_7267,N_7128,N_7184);
or U7268 (N_7268,N_7131,N_7189);
nor U7269 (N_7269,N_7146,N_7124);
nor U7270 (N_7270,N_7109,N_7160);
or U7271 (N_7271,N_7194,N_7144);
nand U7272 (N_7272,N_7191,N_7192);
nor U7273 (N_7273,N_7124,N_7176);
or U7274 (N_7274,N_7180,N_7169);
or U7275 (N_7275,N_7125,N_7134);
nor U7276 (N_7276,N_7139,N_7150);
nor U7277 (N_7277,N_7102,N_7107);
or U7278 (N_7278,N_7147,N_7169);
nor U7279 (N_7279,N_7109,N_7150);
nand U7280 (N_7280,N_7108,N_7137);
or U7281 (N_7281,N_7179,N_7102);
and U7282 (N_7282,N_7154,N_7124);
xor U7283 (N_7283,N_7132,N_7154);
nand U7284 (N_7284,N_7171,N_7150);
nand U7285 (N_7285,N_7197,N_7174);
nor U7286 (N_7286,N_7138,N_7177);
nand U7287 (N_7287,N_7110,N_7162);
nor U7288 (N_7288,N_7193,N_7131);
nand U7289 (N_7289,N_7161,N_7153);
nand U7290 (N_7290,N_7193,N_7183);
and U7291 (N_7291,N_7125,N_7130);
nand U7292 (N_7292,N_7154,N_7121);
nor U7293 (N_7293,N_7120,N_7178);
nand U7294 (N_7294,N_7127,N_7152);
xor U7295 (N_7295,N_7148,N_7156);
or U7296 (N_7296,N_7152,N_7145);
nor U7297 (N_7297,N_7175,N_7183);
or U7298 (N_7298,N_7172,N_7152);
or U7299 (N_7299,N_7161,N_7136);
nand U7300 (N_7300,N_7281,N_7264);
and U7301 (N_7301,N_7257,N_7255);
nor U7302 (N_7302,N_7222,N_7288);
nand U7303 (N_7303,N_7250,N_7291);
nor U7304 (N_7304,N_7251,N_7277);
or U7305 (N_7305,N_7276,N_7227);
nor U7306 (N_7306,N_7203,N_7258);
nor U7307 (N_7307,N_7240,N_7210);
and U7308 (N_7308,N_7298,N_7272);
or U7309 (N_7309,N_7287,N_7217);
nor U7310 (N_7310,N_7228,N_7231);
xnor U7311 (N_7311,N_7234,N_7242);
nor U7312 (N_7312,N_7273,N_7285);
and U7313 (N_7313,N_7214,N_7260);
nor U7314 (N_7314,N_7219,N_7224);
nor U7315 (N_7315,N_7235,N_7201);
or U7316 (N_7316,N_7283,N_7244);
and U7317 (N_7317,N_7241,N_7202);
or U7318 (N_7318,N_7218,N_7247);
or U7319 (N_7319,N_7233,N_7211);
or U7320 (N_7320,N_7230,N_7236);
nand U7321 (N_7321,N_7200,N_7295);
or U7322 (N_7322,N_7263,N_7282);
or U7323 (N_7323,N_7271,N_7293);
and U7324 (N_7324,N_7289,N_7296);
nand U7325 (N_7325,N_7239,N_7238);
nor U7326 (N_7326,N_7254,N_7280);
nor U7327 (N_7327,N_7265,N_7237);
and U7328 (N_7328,N_7248,N_7223);
and U7329 (N_7329,N_7286,N_7253);
and U7330 (N_7330,N_7220,N_7205);
and U7331 (N_7331,N_7294,N_7207);
nand U7332 (N_7332,N_7229,N_7204);
and U7333 (N_7333,N_7275,N_7270);
nor U7334 (N_7334,N_7259,N_7245);
and U7335 (N_7335,N_7292,N_7284);
nand U7336 (N_7336,N_7215,N_7278);
or U7337 (N_7337,N_7297,N_7266);
and U7338 (N_7338,N_7290,N_7274);
nor U7339 (N_7339,N_7213,N_7221);
nor U7340 (N_7340,N_7262,N_7243);
and U7341 (N_7341,N_7249,N_7279);
nor U7342 (N_7342,N_7226,N_7269);
and U7343 (N_7343,N_7256,N_7209);
or U7344 (N_7344,N_7246,N_7252);
and U7345 (N_7345,N_7216,N_7232);
or U7346 (N_7346,N_7206,N_7208);
nor U7347 (N_7347,N_7268,N_7299);
nand U7348 (N_7348,N_7261,N_7225);
or U7349 (N_7349,N_7267,N_7212);
nor U7350 (N_7350,N_7294,N_7247);
and U7351 (N_7351,N_7292,N_7280);
nor U7352 (N_7352,N_7221,N_7218);
nor U7353 (N_7353,N_7200,N_7233);
nor U7354 (N_7354,N_7213,N_7207);
and U7355 (N_7355,N_7276,N_7212);
nor U7356 (N_7356,N_7251,N_7261);
and U7357 (N_7357,N_7227,N_7268);
nor U7358 (N_7358,N_7248,N_7295);
nor U7359 (N_7359,N_7202,N_7221);
nor U7360 (N_7360,N_7257,N_7281);
or U7361 (N_7361,N_7279,N_7299);
and U7362 (N_7362,N_7265,N_7204);
nor U7363 (N_7363,N_7235,N_7286);
or U7364 (N_7364,N_7225,N_7217);
or U7365 (N_7365,N_7243,N_7272);
and U7366 (N_7366,N_7226,N_7243);
nand U7367 (N_7367,N_7259,N_7272);
and U7368 (N_7368,N_7271,N_7205);
or U7369 (N_7369,N_7257,N_7237);
xor U7370 (N_7370,N_7202,N_7242);
nor U7371 (N_7371,N_7201,N_7244);
and U7372 (N_7372,N_7219,N_7208);
and U7373 (N_7373,N_7242,N_7239);
nand U7374 (N_7374,N_7255,N_7200);
or U7375 (N_7375,N_7236,N_7261);
nor U7376 (N_7376,N_7291,N_7275);
nand U7377 (N_7377,N_7215,N_7211);
or U7378 (N_7378,N_7233,N_7296);
nand U7379 (N_7379,N_7283,N_7220);
nand U7380 (N_7380,N_7259,N_7237);
or U7381 (N_7381,N_7293,N_7232);
nand U7382 (N_7382,N_7211,N_7296);
and U7383 (N_7383,N_7260,N_7267);
nand U7384 (N_7384,N_7210,N_7291);
xor U7385 (N_7385,N_7203,N_7229);
or U7386 (N_7386,N_7292,N_7201);
xnor U7387 (N_7387,N_7285,N_7255);
nand U7388 (N_7388,N_7247,N_7251);
or U7389 (N_7389,N_7250,N_7248);
nor U7390 (N_7390,N_7223,N_7288);
and U7391 (N_7391,N_7265,N_7220);
nand U7392 (N_7392,N_7267,N_7289);
or U7393 (N_7393,N_7296,N_7292);
and U7394 (N_7394,N_7299,N_7278);
or U7395 (N_7395,N_7201,N_7245);
nor U7396 (N_7396,N_7255,N_7269);
nor U7397 (N_7397,N_7202,N_7214);
or U7398 (N_7398,N_7270,N_7281);
and U7399 (N_7399,N_7278,N_7294);
or U7400 (N_7400,N_7359,N_7358);
or U7401 (N_7401,N_7336,N_7327);
nand U7402 (N_7402,N_7390,N_7360);
or U7403 (N_7403,N_7352,N_7307);
nand U7404 (N_7404,N_7338,N_7373);
or U7405 (N_7405,N_7389,N_7320);
nand U7406 (N_7406,N_7308,N_7345);
and U7407 (N_7407,N_7372,N_7374);
nand U7408 (N_7408,N_7381,N_7326);
nand U7409 (N_7409,N_7334,N_7365);
or U7410 (N_7410,N_7387,N_7391);
nor U7411 (N_7411,N_7343,N_7313);
nand U7412 (N_7412,N_7323,N_7393);
and U7413 (N_7413,N_7318,N_7310);
nor U7414 (N_7414,N_7368,N_7377);
and U7415 (N_7415,N_7363,N_7328);
and U7416 (N_7416,N_7302,N_7331);
and U7417 (N_7417,N_7347,N_7300);
and U7418 (N_7418,N_7366,N_7329);
or U7419 (N_7419,N_7395,N_7399);
xor U7420 (N_7420,N_7398,N_7333);
and U7421 (N_7421,N_7335,N_7354);
nor U7422 (N_7422,N_7305,N_7380);
nor U7423 (N_7423,N_7386,N_7341);
or U7424 (N_7424,N_7361,N_7304);
or U7425 (N_7425,N_7309,N_7324);
nand U7426 (N_7426,N_7357,N_7376);
nand U7427 (N_7427,N_7371,N_7351);
nor U7428 (N_7428,N_7332,N_7350);
or U7429 (N_7429,N_7317,N_7364);
and U7430 (N_7430,N_7316,N_7301);
or U7431 (N_7431,N_7385,N_7383);
nor U7432 (N_7432,N_7394,N_7375);
nand U7433 (N_7433,N_7355,N_7382);
nand U7434 (N_7434,N_7342,N_7396);
and U7435 (N_7435,N_7312,N_7362);
nor U7436 (N_7436,N_7344,N_7349);
nand U7437 (N_7437,N_7337,N_7397);
or U7438 (N_7438,N_7322,N_7346);
nor U7439 (N_7439,N_7367,N_7303);
or U7440 (N_7440,N_7348,N_7314);
nand U7441 (N_7441,N_7315,N_7370);
or U7442 (N_7442,N_7369,N_7356);
nand U7443 (N_7443,N_7306,N_7379);
nor U7444 (N_7444,N_7325,N_7319);
nor U7445 (N_7445,N_7311,N_7340);
or U7446 (N_7446,N_7339,N_7321);
or U7447 (N_7447,N_7378,N_7392);
nand U7448 (N_7448,N_7353,N_7330);
and U7449 (N_7449,N_7388,N_7384);
nand U7450 (N_7450,N_7355,N_7338);
and U7451 (N_7451,N_7322,N_7313);
or U7452 (N_7452,N_7341,N_7339);
and U7453 (N_7453,N_7388,N_7373);
or U7454 (N_7454,N_7384,N_7337);
nor U7455 (N_7455,N_7310,N_7370);
or U7456 (N_7456,N_7391,N_7351);
or U7457 (N_7457,N_7363,N_7348);
and U7458 (N_7458,N_7397,N_7345);
or U7459 (N_7459,N_7315,N_7300);
nor U7460 (N_7460,N_7366,N_7303);
xor U7461 (N_7461,N_7326,N_7318);
and U7462 (N_7462,N_7356,N_7365);
nand U7463 (N_7463,N_7346,N_7339);
or U7464 (N_7464,N_7370,N_7380);
nand U7465 (N_7465,N_7374,N_7378);
or U7466 (N_7466,N_7329,N_7355);
nor U7467 (N_7467,N_7354,N_7321);
nand U7468 (N_7468,N_7378,N_7339);
and U7469 (N_7469,N_7300,N_7346);
or U7470 (N_7470,N_7383,N_7316);
nand U7471 (N_7471,N_7361,N_7319);
nand U7472 (N_7472,N_7341,N_7329);
nor U7473 (N_7473,N_7388,N_7350);
or U7474 (N_7474,N_7374,N_7331);
or U7475 (N_7475,N_7341,N_7314);
or U7476 (N_7476,N_7348,N_7351);
and U7477 (N_7477,N_7358,N_7398);
nand U7478 (N_7478,N_7301,N_7317);
nor U7479 (N_7479,N_7385,N_7345);
and U7480 (N_7480,N_7320,N_7381);
nand U7481 (N_7481,N_7300,N_7320);
and U7482 (N_7482,N_7344,N_7304);
and U7483 (N_7483,N_7389,N_7350);
nand U7484 (N_7484,N_7345,N_7303);
and U7485 (N_7485,N_7345,N_7383);
xnor U7486 (N_7486,N_7398,N_7350);
or U7487 (N_7487,N_7378,N_7357);
xnor U7488 (N_7488,N_7312,N_7354);
and U7489 (N_7489,N_7352,N_7389);
or U7490 (N_7490,N_7347,N_7398);
or U7491 (N_7491,N_7373,N_7384);
nor U7492 (N_7492,N_7323,N_7385);
and U7493 (N_7493,N_7336,N_7371);
nor U7494 (N_7494,N_7304,N_7363);
nor U7495 (N_7495,N_7386,N_7344);
nand U7496 (N_7496,N_7388,N_7334);
nand U7497 (N_7497,N_7386,N_7309);
nor U7498 (N_7498,N_7341,N_7354);
and U7499 (N_7499,N_7381,N_7360);
nand U7500 (N_7500,N_7449,N_7425);
nand U7501 (N_7501,N_7406,N_7453);
nand U7502 (N_7502,N_7458,N_7421);
and U7503 (N_7503,N_7497,N_7435);
and U7504 (N_7504,N_7447,N_7422);
and U7505 (N_7505,N_7482,N_7401);
nor U7506 (N_7506,N_7484,N_7436);
and U7507 (N_7507,N_7411,N_7410);
nand U7508 (N_7508,N_7439,N_7414);
nor U7509 (N_7509,N_7491,N_7479);
or U7510 (N_7510,N_7465,N_7461);
and U7511 (N_7511,N_7485,N_7487);
nand U7512 (N_7512,N_7496,N_7460);
nor U7513 (N_7513,N_7418,N_7454);
nor U7514 (N_7514,N_7444,N_7452);
nand U7515 (N_7515,N_7499,N_7405);
nand U7516 (N_7516,N_7478,N_7407);
nor U7517 (N_7517,N_7416,N_7403);
and U7518 (N_7518,N_7420,N_7433);
and U7519 (N_7519,N_7486,N_7481);
xor U7520 (N_7520,N_7427,N_7451);
xor U7521 (N_7521,N_7480,N_7415);
and U7522 (N_7522,N_7493,N_7477);
nor U7523 (N_7523,N_7471,N_7476);
nor U7524 (N_7524,N_7426,N_7489);
or U7525 (N_7525,N_7463,N_7498);
xnor U7526 (N_7526,N_7429,N_7442);
nand U7527 (N_7527,N_7431,N_7492);
nand U7528 (N_7528,N_7443,N_7472);
nor U7529 (N_7529,N_7400,N_7432);
and U7530 (N_7530,N_7474,N_7470);
or U7531 (N_7531,N_7495,N_7445);
and U7532 (N_7532,N_7448,N_7490);
nand U7533 (N_7533,N_7409,N_7438);
and U7534 (N_7534,N_7467,N_7404);
nand U7535 (N_7535,N_7456,N_7473);
or U7536 (N_7536,N_7412,N_7455);
and U7537 (N_7537,N_7464,N_7468);
nand U7538 (N_7538,N_7413,N_7488);
nand U7539 (N_7539,N_7446,N_7437);
and U7540 (N_7540,N_7475,N_7430);
and U7541 (N_7541,N_7469,N_7462);
and U7542 (N_7542,N_7428,N_7459);
or U7543 (N_7543,N_7434,N_7419);
and U7544 (N_7544,N_7423,N_7402);
or U7545 (N_7545,N_7441,N_7466);
nor U7546 (N_7546,N_7424,N_7408);
or U7547 (N_7547,N_7457,N_7494);
or U7548 (N_7548,N_7417,N_7483);
nand U7549 (N_7549,N_7440,N_7450);
and U7550 (N_7550,N_7456,N_7492);
nor U7551 (N_7551,N_7487,N_7438);
nor U7552 (N_7552,N_7462,N_7454);
nand U7553 (N_7553,N_7478,N_7459);
nand U7554 (N_7554,N_7490,N_7411);
and U7555 (N_7555,N_7429,N_7476);
and U7556 (N_7556,N_7446,N_7407);
nand U7557 (N_7557,N_7491,N_7481);
and U7558 (N_7558,N_7421,N_7427);
nor U7559 (N_7559,N_7435,N_7476);
nand U7560 (N_7560,N_7487,N_7427);
nor U7561 (N_7561,N_7411,N_7492);
nand U7562 (N_7562,N_7467,N_7431);
xnor U7563 (N_7563,N_7454,N_7435);
nor U7564 (N_7564,N_7493,N_7451);
nand U7565 (N_7565,N_7404,N_7478);
nand U7566 (N_7566,N_7487,N_7419);
nand U7567 (N_7567,N_7414,N_7433);
nand U7568 (N_7568,N_7458,N_7449);
or U7569 (N_7569,N_7403,N_7455);
nand U7570 (N_7570,N_7488,N_7479);
and U7571 (N_7571,N_7434,N_7482);
nor U7572 (N_7572,N_7427,N_7406);
nor U7573 (N_7573,N_7423,N_7418);
nand U7574 (N_7574,N_7467,N_7475);
nand U7575 (N_7575,N_7430,N_7474);
or U7576 (N_7576,N_7407,N_7486);
and U7577 (N_7577,N_7488,N_7493);
nor U7578 (N_7578,N_7407,N_7448);
or U7579 (N_7579,N_7463,N_7483);
nand U7580 (N_7580,N_7440,N_7429);
nor U7581 (N_7581,N_7442,N_7443);
and U7582 (N_7582,N_7459,N_7449);
or U7583 (N_7583,N_7455,N_7440);
and U7584 (N_7584,N_7437,N_7422);
nor U7585 (N_7585,N_7448,N_7444);
or U7586 (N_7586,N_7416,N_7404);
nand U7587 (N_7587,N_7451,N_7494);
nor U7588 (N_7588,N_7456,N_7495);
or U7589 (N_7589,N_7477,N_7472);
and U7590 (N_7590,N_7435,N_7494);
nor U7591 (N_7591,N_7476,N_7472);
and U7592 (N_7592,N_7480,N_7495);
and U7593 (N_7593,N_7499,N_7442);
nand U7594 (N_7594,N_7455,N_7492);
nand U7595 (N_7595,N_7441,N_7488);
nor U7596 (N_7596,N_7469,N_7415);
or U7597 (N_7597,N_7481,N_7466);
nor U7598 (N_7598,N_7418,N_7403);
nand U7599 (N_7599,N_7491,N_7496);
or U7600 (N_7600,N_7586,N_7535);
or U7601 (N_7601,N_7577,N_7505);
or U7602 (N_7602,N_7539,N_7529);
or U7603 (N_7603,N_7572,N_7544);
or U7604 (N_7604,N_7531,N_7502);
and U7605 (N_7605,N_7545,N_7579);
nor U7606 (N_7606,N_7590,N_7508);
nand U7607 (N_7607,N_7582,N_7588);
nor U7608 (N_7608,N_7525,N_7526);
and U7609 (N_7609,N_7589,N_7559);
or U7610 (N_7610,N_7514,N_7536);
nor U7611 (N_7611,N_7511,N_7533);
or U7612 (N_7612,N_7520,N_7542);
or U7613 (N_7613,N_7575,N_7538);
or U7614 (N_7614,N_7598,N_7595);
nor U7615 (N_7615,N_7571,N_7563);
and U7616 (N_7616,N_7509,N_7537);
or U7617 (N_7617,N_7557,N_7599);
or U7618 (N_7618,N_7528,N_7596);
nor U7619 (N_7619,N_7510,N_7521);
and U7620 (N_7620,N_7556,N_7594);
nor U7621 (N_7621,N_7513,N_7551);
nor U7622 (N_7622,N_7500,N_7562);
xor U7623 (N_7623,N_7517,N_7541);
or U7624 (N_7624,N_7552,N_7518);
and U7625 (N_7625,N_7532,N_7506);
nor U7626 (N_7626,N_7553,N_7585);
nor U7627 (N_7627,N_7555,N_7581);
nand U7628 (N_7628,N_7522,N_7527);
nand U7629 (N_7629,N_7560,N_7591);
or U7630 (N_7630,N_7543,N_7550);
or U7631 (N_7631,N_7549,N_7570);
nand U7632 (N_7632,N_7573,N_7584);
nor U7633 (N_7633,N_7567,N_7597);
or U7634 (N_7634,N_7501,N_7578);
and U7635 (N_7635,N_7530,N_7524);
nand U7636 (N_7636,N_7558,N_7507);
nand U7637 (N_7637,N_7565,N_7548);
or U7638 (N_7638,N_7503,N_7580);
and U7639 (N_7639,N_7576,N_7546);
and U7640 (N_7640,N_7561,N_7547);
and U7641 (N_7641,N_7574,N_7566);
and U7642 (N_7642,N_7568,N_7534);
and U7643 (N_7643,N_7593,N_7569);
or U7644 (N_7644,N_7504,N_7564);
nor U7645 (N_7645,N_7523,N_7516);
nor U7646 (N_7646,N_7583,N_7554);
or U7647 (N_7647,N_7592,N_7512);
nor U7648 (N_7648,N_7540,N_7587);
nor U7649 (N_7649,N_7519,N_7515);
nand U7650 (N_7650,N_7599,N_7545);
or U7651 (N_7651,N_7588,N_7565);
nand U7652 (N_7652,N_7590,N_7581);
nor U7653 (N_7653,N_7585,N_7594);
nand U7654 (N_7654,N_7531,N_7563);
nor U7655 (N_7655,N_7592,N_7558);
and U7656 (N_7656,N_7506,N_7593);
nor U7657 (N_7657,N_7523,N_7588);
nor U7658 (N_7658,N_7532,N_7552);
or U7659 (N_7659,N_7523,N_7585);
and U7660 (N_7660,N_7532,N_7534);
and U7661 (N_7661,N_7512,N_7539);
and U7662 (N_7662,N_7548,N_7580);
or U7663 (N_7663,N_7526,N_7585);
nand U7664 (N_7664,N_7591,N_7556);
nor U7665 (N_7665,N_7523,N_7569);
nor U7666 (N_7666,N_7535,N_7503);
or U7667 (N_7667,N_7515,N_7555);
nor U7668 (N_7668,N_7501,N_7560);
and U7669 (N_7669,N_7558,N_7598);
or U7670 (N_7670,N_7521,N_7513);
nand U7671 (N_7671,N_7512,N_7553);
or U7672 (N_7672,N_7556,N_7506);
or U7673 (N_7673,N_7540,N_7561);
nand U7674 (N_7674,N_7505,N_7547);
nand U7675 (N_7675,N_7501,N_7565);
and U7676 (N_7676,N_7577,N_7587);
or U7677 (N_7677,N_7589,N_7517);
nor U7678 (N_7678,N_7535,N_7532);
or U7679 (N_7679,N_7551,N_7552);
nand U7680 (N_7680,N_7556,N_7565);
nor U7681 (N_7681,N_7591,N_7540);
nor U7682 (N_7682,N_7557,N_7548);
or U7683 (N_7683,N_7565,N_7526);
and U7684 (N_7684,N_7581,N_7516);
nor U7685 (N_7685,N_7507,N_7526);
and U7686 (N_7686,N_7598,N_7556);
nor U7687 (N_7687,N_7590,N_7579);
nand U7688 (N_7688,N_7519,N_7548);
and U7689 (N_7689,N_7527,N_7510);
and U7690 (N_7690,N_7568,N_7504);
or U7691 (N_7691,N_7546,N_7539);
and U7692 (N_7692,N_7561,N_7515);
xnor U7693 (N_7693,N_7522,N_7567);
or U7694 (N_7694,N_7532,N_7503);
and U7695 (N_7695,N_7503,N_7549);
or U7696 (N_7696,N_7515,N_7593);
and U7697 (N_7697,N_7509,N_7596);
nor U7698 (N_7698,N_7566,N_7503);
and U7699 (N_7699,N_7509,N_7538);
and U7700 (N_7700,N_7653,N_7698);
nor U7701 (N_7701,N_7681,N_7688);
and U7702 (N_7702,N_7657,N_7638);
or U7703 (N_7703,N_7650,N_7669);
nor U7704 (N_7704,N_7623,N_7608);
or U7705 (N_7705,N_7654,N_7685);
nand U7706 (N_7706,N_7675,N_7601);
nand U7707 (N_7707,N_7602,N_7677);
and U7708 (N_7708,N_7635,N_7600);
nor U7709 (N_7709,N_7614,N_7663);
nand U7710 (N_7710,N_7691,N_7619);
and U7711 (N_7711,N_7649,N_7617);
xnor U7712 (N_7712,N_7613,N_7692);
or U7713 (N_7713,N_7660,N_7620);
or U7714 (N_7714,N_7626,N_7690);
or U7715 (N_7715,N_7629,N_7670);
or U7716 (N_7716,N_7616,N_7651);
nand U7717 (N_7717,N_7645,N_7695);
or U7718 (N_7718,N_7680,N_7665);
nand U7719 (N_7719,N_7612,N_7643);
and U7720 (N_7720,N_7609,N_7622);
nor U7721 (N_7721,N_7667,N_7672);
or U7722 (N_7722,N_7696,N_7636);
nor U7723 (N_7723,N_7687,N_7673);
nand U7724 (N_7724,N_7684,N_7659);
or U7725 (N_7725,N_7694,N_7634);
xnor U7726 (N_7726,N_7674,N_7644);
and U7727 (N_7727,N_7640,N_7624);
nor U7728 (N_7728,N_7604,N_7605);
or U7729 (N_7729,N_7631,N_7686);
nor U7730 (N_7730,N_7607,N_7628);
nor U7731 (N_7731,N_7656,N_7641);
nand U7732 (N_7732,N_7664,N_7661);
or U7733 (N_7733,N_7633,N_7642);
and U7734 (N_7734,N_7632,N_7621);
or U7735 (N_7735,N_7671,N_7615);
or U7736 (N_7736,N_7627,N_7697);
nand U7737 (N_7737,N_7610,N_7652);
nor U7738 (N_7738,N_7689,N_7666);
or U7739 (N_7739,N_7647,N_7618);
nand U7740 (N_7740,N_7639,N_7603);
or U7741 (N_7741,N_7625,N_7679);
or U7742 (N_7742,N_7682,N_7699);
and U7743 (N_7743,N_7658,N_7630);
or U7744 (N_7744,N_7606,N_7676);
and U7745 (N_7745,N_7668,N_7662);
nand U7746 (N_7746,N_7683,N_7693);
or U7747 (N_7747,N_7655,N_7646);
and U7748 (N_7748,N_7611,N_7648);
nor U7749 (N_7749,N_7637,N_7678);
and U7750 (N_7750,N_7600,N_7637);
nor U7751 (N_7751,N_7621,N_7653);
nor U7752 (N_7752,N_7622,N_7635);
nand U7753 (N_7753,N_7637,N_7640);
nand U7754 (N_7754,N_7631,N_7695);
nor U7755 (N_7755,N_7661,N_7669);
and U7756 (N_7756,N_7697,N_7657);
and U7757 (N_7757,N_7647,N_7601);
or U7758 (N_7758,N_7674,N_7648);
or U7759 (N_7759,N_7614,N_7628);
or U7760 (N_7760,N_7692,N_7654);
nand U7761 (N_7761,N_7685,N_7646);
and U7762 (N_7762,N_7607,N_7602);
nand U7763 (N_7763,N_7623,N_7672);
nand U7764 (N_7764,N_7608,N_7670);
nand U7765 (N_7765,N_7646,N_7622);
nor U7766 (N_7766,N_7625,N_7659);
and U7767 (N_7767,N_7637,N_7604);
and U7768 (N_7768,N_7695,N_7600);
or U7769 (N_7769,N_7601,N_7603);
nor U7770 (N_7770,N_7695,N_7613);
and U7771 (N_7771,N_7688,N_7614);
nand U7772 (N_7772,N_7613,N_7665);
or U7773 (N_7773,N_7618,N_7610);
and U7774 (N_7774,N_7618,N_7609);
nand U7775 (N_7775,N_7620,N_7605);
nand U7776 (N_7776,N_7648,N_7644);
or U7777 (N_7777,N_7663,N_7639);
nor U7778 (N_7778,N_7655,N_7622);
nand U7779 (N_7779,N_7652,N_7607);
nand U7780 (N_7780,N_7693,N_7690);
nor U7781 (N_7781,N_7644,N_7695);
or U7782 (N_7782,N_7602,N_7627);
nand U7783 (N_7783,N_7603,N_7692);
nor U7784 (N_7784,N_7696,N_7669);
nand U7785 (N_7785,N_7601,N_7635);
or U7786 (N_7786,N_7631,N_7617);
nor U7787 (N_7787,N_7642,N_7694);
nor U7788 (N_7788,N_7605,N_7652);
nand U7789 (N_7789,N_7618,N_7613);
nand U7790 (N_7790,N_7628,N_7610);
nor U7791 (N_7791,N_7637,N_7669);
nor U7792 (N_7792,N_7658,N_7628);
nand U7793 (N_7793,N_7604,N_7655);
nor U7794 (N_7794,N_7637,N_7676);
nand U7795 (N_7795,N_7661,N_7699);
nand U7796 (N_7796,N_7680,N_7634);
and U7797 (N_7797,N_7618,N_7694);
and U7798 (N_7798,N_7661,N_7680);
or U7799 (N_7799,N_7639,N_7643);
nor U7800 (N_7800,N_7709,N_7721);
nor U7801 (N_7801,N_7754,N_7776);
nand U7802 (N_7802,N_7775,N_7717);
nand U7803 (N_7803,N_7711,N_7761);
or U7804 (N_7804,N_7798,N_7746);
or U7805 (N_7805,N_7741,N_7778);
nand U7806 (N_7806,N_7724,N_7765);
nor U7807 (N_7807,N_7705,N_7793);
and U7808 (N_7808,N_7730,N_7769);
and U7809 (N_7809,N_7757,N_7787);
nand U7810 (N_7810,N_7700,N_7743);
or U7811 (N_7811,N_7773,N_7722);
nand U7812 (N_7812,N_7751,N_7726);
nand U7813 (N_7813,N_7745,N_7794);
and U7814 (N_7814,N_7771,N_7748);
nor U7815 (N_7815,N_7752,N_7718);
and U7816 (N_7816,N_7767,N_7782);
and U7817 (N_7817,N_7796,N_7768);
and U7818 (N_7818,N_7733,N_7783);
and U7819 (N_7819,N_7728,N_7715);
nand U7820 (N_7820,N_7790,N_7753);
nor U7821 (N_7821,N_7779,N_7760);
nor U7822 (N_7822,N_7714,N_7788);
nand U7823 (N_7823,N_7762,N_7750);
nand U7824 (N_7824,N_7723,N_7719);
nand U7825 (N_7825,N_7799,N_7732);
and U7826 (N_7826,N_7742,N_7755);
or U7827 (N_7827,N_7786,N_7702);
xnor U7828 (N_7828,N_7784,N_7701);
nand U7829 (N_7829,N_7797,N_7747);
nor U7830 (N_7830,N_7772,N_7792);
nor U7831 (N_7831,N_7791,N_7710);
nand U7832 (N_7832,N_7770,N_7720);
nand U7833 (N_7833,N_7763,N_7774);
and U7834 (N_7834,N_7764,N_7766);
and U7835 (N_7835,N_7738,N_7713);
or U7836 (N_7836,N_7780,N_7781);
nand U7837 (N_7837,N_7735,N_7725);
nand U7838 (N_7838,N_7758,N_7739);
nand U7839 (N_7839,N_7789,N_7785);
or U7840 (N_7840,N_7740,N_7737);
and U7841 (N_7841,N_7731,N_7736);
nand U7842 (N_7842,N_7795,N_7749);
nor U7843 (N_7843,N_7708,N_7707);
nand U7844 (N_7844,N_7706,N_7703);
or U7845 (N_7845,N_7727,N_7759);
nor U7846 (N_7846,N_7777,N_7734);
and U7847 (N_7847,N_7716,N_7712);
or U7848 (N_7848,N_7704,N_7729);
and U7849 (N_7849,N_7756,N_7744);
nand U7850 (N_7850,N_7724,N_7725);
nor U7851 (N_7851,N_7733,N_7779);
nand U7852 (N_7852,N_7704,N_7717);
nor U7853 (N_7853,N_7750,N_7785);
or U7854 (N_7854,N_7772,N_7702);
or U7855 (N_7855,N_7738,N_7785);
nor U7856 (N_7856,N_7759,N_7704);
nor U7857 (N_7857,N_7769,N_7748);
xor U7858 (N_7858,N_7766,N_7799);
and U7859 (N_7859,N_7730,N_7742);
nand U7860 (N_7860,N_7741,N_7773);
or U7861 (N_7861,N_7794,N_7774);
and U7862 (N_7862,N_7759,N_7762);
or U7863 (N_7863,N_7792,N_7786);
and U7864 (N_7864,N_7738,N_7771);
and U7865 (N_7865,N_7794,N_7787);
or U7866 (N_7866,N_7745,N_7752);
nor U7867 (N_7867,N_7720,N_7706);
nor U7868 (N_7868,N_7718,N_7701);
and U7869 (N_7869,N_7713,N_7703);
and U7870 (N_7870,N_7788,N_7723);
nand U7871 (N_7871,N_7797,N_7756);
or U7872 (N_7872,N_7732,N_7713);
nand U7873 (N_7873,N_7770,N_7763);
nand U7874 (N_7874,N_7713,N_7721);
and U7875 (N_7875,N_7712,N_7721);
nand U7876 (N_7876,N_7765,N_7722);
nand U7877 (N_7877,N_7743,N_7734);
and U7878 (N_7878,N_7766,N_7719);
and U7879 (N_7879,N_7777,N_7787);
or U7880 (N_7880,N_7772,N_7713);
and U7881 (N_7881,N_7766,N_7794);
and U7882 (N_7882,N_7772,N_7739);
nand U7883 (N_7883,N_7720,N_7724);
nor U7884 (N_7884,N_7731,N_7793);
nand U7885 (N_7885,N_7730,N_7719);
and U7886 (N_7886,N_7700,N_7722);
or U7887 (N_7887,N_7709,N_7763);
nand U7888 (N_7888,N_7772,N_7793);
nand U7889 (N_7889,N_7795,N_7774);
or U7890 (N_7890,N_7735,N_7762);
nand U7891 (N_7891,N_7707,N_7780);
or U7892 (N_7892,N_7701,N_7756);
nand U7893 (N_7893,N_7736,N_7780);
or U7894 (N_7894,N_7786,N_7704);
and U7895 (N_7895,N_7708,N_7781);
or U7896 (N_7896,N_7708,N_7721);
nand U7897 (N_7897,N_7779,N_7771);
and U7898 (N_7898,N_7713,N_7710);
or U7899 (N_7899,N_7701,N_7745);
or U7900 (N_7900,N_7809,N_7802);
nand U7901 (N_7901,N_7864,N_7878);
xnor U7902 (N_7902,N_7835,N_7873);
nand U7903 (N_7903,N_7896,N_7876);
nor U7904 (N_7904,N_7895,N_7803);
nor U7905 (N_7905,N_7885,N_7890);
or U7906 (N_7906,N_7879,N_7869);
or U7907 (N_7907,N_7826,N_7807);
nor U7908 (N_7908,N_7867,N_7813);
or U7909 (N_7909,N_7814,N_7829);
nand U7910 (N_7910,N_7801,N_7881);
nand U7911 (N_7911,N_7868,N_7870);
nor U7912 (N_7912,N_7817,N_7863);
or U7913 (N_7913,N_7845,N_7841);
and U7914 (N_7914,N_7816,N_7836);
nor U7915 (N_7915,N_7893,N_7842);
nor U7916 (N_7916,N_7861,N_7874);
nand U7917 (N_7917,N_7860,N_7818);
nor U7918 (N_7918,N_7833,N_7837);
and U7919 (N_7919,N_7828,N_7849);
and U7920 (N_7920,N_7827,N_7871);
or U7921 (N_7921,N_7865,N_7851);
or U7922 (N_7922,N_7875,N_7853);
and U7923 (N_7923,N_7825,N_7854);
nand U7924 (N_7924,N_7810,N_7886);
or U7925 (N_7925,N_7891,N_7832);
nand U7926 (N_7926,N_7858,N_7823);
or U7927 (N_7927,N_7811,N_7899);
nor U7928 (N_7928,N_7848,N_7872);
nor U7929 (N_7929,N_7824,N_7859);
and U7930 (N_7930,N_7897,N_7847);
nand U7931 (N_7931,N_7880,N_7806);
nand U7932 (N_7932,N_7819,N_7883);
or U7933 (N_7933,N_7884,N_7804);
and U7934 (N_7934,N_7834,N_7850);
nor U7935 (N_7935,N_7831,N_7846);
nor U7936 (N_7936,N_7830,N_7820);
nand U7937 (N_7937,N_7805,N_7855);
or U7938 (N_7938,N_7856,N_7857);
or U7939 (N_7939,N_7877,N_7888);
and U7940 (N_7940,N_7815,N_7840);
or U7941 (N_7941,N_7894,N_7844);
or U7942 (N_7942,N_7838,N_7889);
nor U7943 (N_7943,N_7822,N_7862);
nand U7944 (N_7944,N_7898,N_7843);
or U7945 (N_7945,N_7852,N_7887);
nor U7946 (N_7946,N_7812,N_7892);
nand U7947 (N_7947,N_7808,N_7839);
xor U7948 (N_7948,N_7821,N_7800);
nor U7949 (N_7949,N_7882,N_7866);
and U7950 (N_7950,N_7873,N_7884);
nand U7951 (N_7951,N_7872,N_7899);
and U7952 (N_7952,N_7812,N_7821);
nor U7953 (N_7953,N_7803,N_7856);
nor U7954 (N_7954,N_7854,N_7856);
or U7955 (N_7955,N_7896,N_7839);
nor U7956 (N_7956,N_7801,N_7844);
and U7957 (N_7957,N_7848,N_7871);
or U7958 (N_7958,N_7821,N_7809);
and U7959 (N_7959,N_7891,N_7800);
and U7960 (N_7960,N_7891,N_7846);
nand U7961 (N_7961,N_7800,N_7812);
nand U7962 (N_7962,N_7884,N_7801);
and U7963 (N_7963,N_7807,N_7839);
nand U7964 (N_7964,N_7844,N_7853);
nand U7965 (N_7965,N_7818,N_7880);
nand U7966 (N_7966,N_7811,N_7826);
nor U7967 (N_7967,N_7837,N_7883);
and U7968 (N_7968,N_7818,N_7875);
and U7969 (N_7969,N_7835,N_7844);
nand U7970 (N_7970,N_7837,N_7803);
or U7971 (N_7971,N_7893,N_7875);
xor U7972 (N_7972,N_7884,N_7894);
or U7973 (N_7973,N_7852,N_7833);
and U7974 (N_7974,N_7898,N_7867);
nand U7975 (N_7975,N_7895,N_7811);
nand U7976 (N_7976,N_7813,N_7849);
and U7977 (N_7977,N_7859,N_7819);
and U7978 (N_7978,N_7834,N_7886);
nor U7979 (N_7979,N_7895,N_7835);
or U7980 (N_7980,N_7856,N_7868);
xor U7981 (N_7981,N_7808,N_7847);
nor U7982 (N_7982,N_7848,N_7843);
and U7983 (N_7983,N_7819,N_7882);
or U7984 (N_7984,N_7899,N_7873);
or U7985 (N_7985,N_7826,N_7808);
nor U7986 (N_7986,N_7864,N_7854);
nand U7987 (N_7987,N_7877,N_7827);
nand U7988 (N_7988,N_7855,N_7809);
and U7989 (N_7989,N_7872,N_7884);
nand U7990 (N_7990,N_7846,N_7804);
nand U7991 (N_7991,N_7859,N_7874);
nand U7992 (N_7992,N_7881,N_7819);
nor U7993 (N_7993,N_7890,N_7830);
and U7994 (N_7994,N_7845,N_7869);
and U7995 (N_7995,N_7838,N_7874);
and U7996 (N_7996,N_7885,N_7851);
and U7997 (N_7997,N_7882,N_7801);
and U7998 (N_7998,N_7820,N_7840);
nand U7999 (N_7999,N_7886,N_7897);
nand U8000 (N_8000,N_7900,N_7967);
nor U8001 (N_8001,N_7990,N_7980);
or U8002 (N_8002,N_7915,N_7905);
or U8003 (N_8003,N_7998,N_7959);
or U8004 (N_8004,N_7952,N_7983);
and U8005 (N_8005,N_7927,N_7932);
or U8006 (N_8006,N_7933,N_7995);
nor U8007 (N_8007,N_7924,N_7951);
nor U8008 (N_8008,N_7907,N_7955);
nand U8009 (N_8009,N_7961,N_7934);
nor U8010 (N_8010,N_7936,N_7992);
nand U8011 (N_8011,N_7908,N_7965);
xor U8012 (N_8012,N_7984,N_7968);
nor U8013 (N_8013,N_7975,N_7991);
nand U8014 (N_8014,N_7914,N_7943);
and U8015 (N_8015,N_7910,N_7994);
xnor U8016 (N_8016,N_7942,N_7938);
nor U8017 (N_8017,N_7977,N_7997);
nand U8018 (N_8018,N_7903,N_7957);
and U8019 (N_8019,N_7950,N_7970);
and U8020 (N_8020,N_7989,N_7960);
and U8021 (N_8021,N_7911,N_7945);
or U8022 (N_8022,N_7976,N_7921);
or U8023 (N_8023,N_7913,N_7941);
or U8024 (N_8024,N_7901,N_7981);
nand U8025 (N_8025,N_7904,N_7935);
and U8026 (N_8026,N_7917,N_7931);
nor U8027 (N_8027,N_7956,N_7971);
nor U8028 (N_8028,N_7906,N_7918);
or U8029 (N_8029,N_7946,N_7972);
and U8030 (N_8030,N_7979,N_7948);
and U8031 (N_8031,N_7925,N_7930);
or U8032 (N_8032,N_7944,N_7922);
nor U8033 (N_8033,N_7929,N_7987);
or U8034 (N_8034,N_7947,N_7988);
nand U8035 (N_8035,N_7909,N_7964);
or U8036 (N_8036,N_7966,N_7996);
or U8037 (N_8037,N_7920,N_7949);
nor U8038 (N_8038,N_7963,N_7986);
or U8039 (N_8039,N_7999,N_7937);
and U8040 (N_8040,N_7923,N_7953);
nand U8041 (N_8041,N_7969,N_7954);
and U8042 (N_8042,N_7962,N_7939);
and U8043 (N_8043,N_7916,N_7982);
nor U8044 (N_8044,N_7973,N_7978);
nand U8045 (N_8045,N_7940,N_7928);
or U8046 (N_8046,N_7926,N_7985);
nand U8047 (N_8047,N_7993,N_7974);
and U8048 (N_8048,N_7958,N_7919);
nand U8049 (N_8049,N_7902,N_7912);
or U8050 (N_8050,N_7997,N_7929);
xnor U8051 (N_8051,N_7915,N_7962);
and U8052 (N_8052,N_7921,N_7988);
or U8053 (N_8053,N_7913,N_7962);
and U8054 (N_8054,N_7998,N_7909);
xor U8055 (N_8055,N_7916,N_7965);
nor U8056 (N_8056,N_7900,N_7978);
or U8057 (N_8057,N_7920,N_7964);
or U8058 (N_8058,N_7922,N_7988);
nor U8059 (N_8059,N_7900,N_7980);
or U8060 (N_8060,N_7902,N_7977);
or U8061 (N_8061,N_7972,N_7959);
nor U8062 (N_8062,N_7930,N_7980);
and U8063 (N_8063,N_7978,N_7938);
nand U8064 (N_8064,N_7955,N_7949);
nand U8065 (N_8065,N_7962,N_7927);
nor U8066 (N_8066,N_7939,N_7948);
nor U8067 (N_8067,N_7967,N_7956);
or U8068 (N_8068,N_7974,N_7906);
and U8069 (N_8069,N_7957,N_7900);
nor U8070 (N_8070,N_7994,N_7926);
or U8071 (N_8071,N_7972,N_7950);
nor U8072 (N_8072,N_7929,N_7936);
or U8073 (N_8073,N_7966,N_7947);
nor U8074 (N_8074,N_7936,N_7924);
nor U8075 (N_8075,N_7947,N_7986);
or U8076 (N_8076,N_7994,N_7999);
nand U8077 (N_8077,N_7914,N_7974);
and U8078 (N_8078,N_7993,N_7909);
nor U8079 (N_8079,N_7996,N_7918);
nand U8080 (N_8080,N_7934,N_7910);
or U8081 (N_8081,N_7946,N_7937);
or U8082 (N_8082,N_7968,N_7951);
nor U8083 (N_8083,N_7998,N_7930);
nand U8084 (N_8084,N_7914,N_7978);
nand U8085 (N_8085,N_7944,N_7951);
and U8086 (N_8086,N_7959,N_7939);
and U8087 (N_8087,N_7957,N_7916);
nor U8088 (N_8088,N_7970,N_7904);
and U8089 (N_8089,N_7966,N_7994);
and U8090 (N_8090,N_7909,N_7937);
nor U8091 (N_8091,N_7906,N_7995);
or U8092 (N_8092,N_7903,N_7932);
nor U8093 (N_8093,N_7900,N_7976);
or U8094 (N_8094,N_7928,N_7913);
or U8095 (N_8095,N_7956,N_7906);
nor U8096 (N_8096,N_7940,N_7933);
nand U8097 (N_8097,N_7909,N_7995);
nor U8098 (N_8098,N_7989,N_7997);
and U8099 (N_8099,N_7963,N_7915);
or U8100 (N_8100,N_8082,N_8057);
nor U8101 (N_8101,N_8005,N_8014);
nor U8102 (N_8102,N_8072,N_8068);
nor U8103 (N_8103,N_8094,N_8044);
and U8104 (N_8104,N_8086,N_8066);
xnor U8105 (N_8105,N_8036,N_8037);
nor U8106 (N_8106,N_8000,N_8034);
nor U8107 (N_8107,N_8067,N_8045);
or U8108 (N_8108,N_8070,N_8080);
nor U8109 (N_8109,N_8084,N_8018);
nand U8110 (N_8110,N_8095,N_8056);
and U8111 (N_8111,N_8030,N_8091);
and U8112 (N_8112,N_8029,N_8053);
or U8113 (N_8113,N_8027,N_8017);
or U8114 (N_8114,N_8088,N_8058);
or U8115 (N_8115,N_8071,N_8064);
or U8116 (N_8116,N_8015,N_8033);
or U8117 (N_8117,N_8073,N_8010);
or U8118 (N_8118,N_8042,N_8093);
and U8119 (N_8119,N_8023,N_8047);
nand U8120 (N_8120,N_8008,N_8048);
or U8121 (N_8121,N_8003,N_8032);
nor U8122 (N_8122,N_8096,N_8039);
nand U8123 (N_8123,N_8081,N_8055);
nor U8124 (N_8124,N_8031,N_8009);
nor U8125 (N_8125,N_8085,N_8092);
and U8126 (N_8126,N_8078,N_8074);
or U8127 (N_8127,N_8063,N_8040);
and U8128 (N_8128,N_8035,N_8075);
nor U8129 (N_8129,N_8060,N_8062);
or U8130 (N_8130,N_8043,N_8004);
or U8131 (N_8131,N_8059,N_8099);
and U8132 (N_8132,N_8089,N_8012);
nand U8133 (N_8133,N_8061,N_8001);
nor U8134 (N_8134,N_8069,N_8002);
and U8135 (N_8135,N_8028,N_8041);
nor U8136 (N_8136,N_8025,N_8049);
and U8137 (N_8137,N_8007,N_8079);
nor U8138 (N_8138,N_8021,N_8046);
and U8139 (N_8139,N_8050,N_8083);
and U8140 (N_8140,N_8098,N_8019);
and U8141 (N_8141,N_8016,N_8020);
or U8142 (N_8142,N_8090,N_8052);
and U8143 (N_8143,N_8054,N_8011);
nand U8144 (N_8144,N_8077,N_8024);
and U8145 (N_8145,N_8013,N_8087);
nor U8146 (N_8146,N_8097,N_8038);
or U8147 (N_8147,N_8051,N_8065);
or U8148 (N_8148,N_8076,N_8006);
nor U8149 (N_8149,N_8022,N_8026);
nor U8150 (N_8150,N_8003,N_8012);
nor U8151 (N_8151,N_8058,N_8092);
and U8152 (N_8152,N_8091,N_8079);
and U8153 (N_8153,N_8034,N_8095);
and U8154 (N_8154,N_8086,N_8041);
or U8155 (N_8155,N_8067,N_8021);
nand U8156 (N_8156,N_8059,N_8044);
and U8157 (N_8157,N_8037,N_8010);
and U8158 (N_8158,N_8036,N_8020);
and U8159 (N_8159,N_8098,N_8070);
nand U8160 (N_8160,N_8004,N_8077);
nor U8161 (N_8161,N_8036,N_8027);
or U8162 (N_8162,N_8094,N_8022);
nand U8163 (N_8163,N_8049,N_8047);
nand U8164 (N_8164,N_8070,N_8093);
or U8165 (N_8165,N_8009,N_8003);
or U8166 (N_8166,N_8055,N_8077);
nor U8167 (N_8167,N_8016,N_8090);
nand U8168 (N_8168,N_8048,N_8027);
and U8169 (N_8169,N_8099,N_8027);
nor U8170 (N_8170,N_8039,N_8050);
and U8171 (N_8171,N_8073,N_8034);
and U8172 (N_8172,N_8087,N_8027);
or U8173 (N_8173,N_8059,N_8062);
nand U8174 (N_8174,N_8039,N_8051);
and U8175 (N_8175,N_8069,N_8080);
nand U8176 (N_8176,N_8081,N_8024);
or U8177 (N_8177,N_8028,N_8025);
or U8178 (N_8178,N_8038,N_8071);
or U8179 (N_8179,N_8057,N_8087);
or U8180 (N_8180,N_8062,N_8039);
and U8181 (N_8181,N_8003,N_8059);
and U8182 (N_8182,N_8088,N_8021);
and U8183 (N_8183,N_8070,N_8006);
nand U8184 (N_8184,N_8043,N_8078);
and U8185 (N_8185,N_8044,N_8030);
or U8186 (N_8186,N_8053,N_8065);
or U8187 (N_8187,N_8029,N_8004);
or U8188 (N_8188,N_8012,N_8019);
and U8189 (N_8189,N_8085,N_8020);
and U8190 (N_8190,N_8080,N_8094);
and U8191 (N_8191,N_8086,N_8033);
nand U8192 (N_8192,N_8026,N_8025);
and U8193 (N_8193,N_8014,N_8068);
or U8194 (N_8194,N_8054,N_8056);
nand U8195 (N_8195,N_8019,N_8003);
nand U8196 (N_8196,N_8018,N_8024);
and U8197 (N_8197,N_8096,N_8054);
nor U8198 (N_8198,N_8090,N_8004);
and U8199 (N_8199,N_8070,N_8053);
or U8200 (N_8200,N_8147,N_8168);
nand U8201 (N_8201,N_8182,N_8110);
nor U8202 (N_8202,N_8169,N_8143);
nor U8203 (N_8203,N_8179,N_8197);
and U8204 (N_8204,N_8101,N_8154);
xor U8205 (N_8205,N_8131,N_8142);
nor U8206 (N_8206,N_8151,N_8180);
nor U8207 (N_8207,N_8146,N_8144);
or U8208 (N_8208,N_8170,N_8149);
or U8209 (N_8209,N_8105,N_8164);
nor U8210 (N_8210,N_8145,N_8166);
nand U8211 (N_8211,N_8187,N_8152);
nor U8212 (N_8212,N_8102,N_8132);
or U8213 (N_8213,N_8186,N_8192);
or U8214 (N_8214,N_8108,N_8106);
nor U8215 (N_8215,N_8159,N_8163);
nand U8216 (N_8216,N_8127,N_8117);
and U8217 (N_8217,N_8150,N_8140);
nor U8218 (N_8218,N_8115,N_8174);
nor U8219 (N_8219,N_8194,N_8128);
or U8220 (N_8220,N_8113,N_8122);
nor U8221 (N_8221,N_8171,N_8100);
nor U8222 (N_8222,N_8116,N_8118);
nand U8223 (N_8223,N_8199,N_8167);
and U8224 (N_8224,N_8158,N_8160);
or U8225 (N_8225,N_8157,N_8148);
nand U8226 (N_8226,N_8193,N_8126);
or U8227 (N_8227,N_8121,N_8136);
or U8228 (N_8228,N_8165,N_8181);
and U8229 (N_8229,N_8191,N_8141);
or U8230 (N_8230,N_8119,N_8109);
nand U8231 (N_8231,N_8130,N_8162);
and U8232 (N_8232,N_8155,N_8188);
and U8233 (N_8233,N_8103,N_8112);
nor U8234 (N_8234,N_8190,N_8172);
nand U8235 (N_8235,N_8161,N_8137);
nand U8236 (N_8236,N_8124,N_8153);
nand U8237 (N_8237,N_8114,N_8198);
nor U8238 (N_8238,N_8173,N_8189);
or U8239 (N_8239,N_8175,N_8129);
or U8240 (N_8240,N_8183,N_8184);
and U8241 (N_8241,N_8178,N_8196);
or U8242 (N_8242,N_8125,N_8185);
nor U8243 (N_8243,N_8138,N_8104);
and U8244 (N_8244,N_8135,N_8177);
and U8245 (N_8245,N_8107,N_8133);
and U8246 (N_8246,N_8139,N_8195);
or U8247 (N_8247,N_8120,N_8176);
nor U8248 (N_8248,N_8123,N_8111);
and U8249 (N_8249,N_8134,N_8156);
nor U8250 (N_8250,N_8160,N_8124);
nand U8251 (N_8251,N_8110,N_8158);
or U8252 (N_8252,N_8123,N_8128);
nand U8253 (N_8253,N_8139,N_8168);
or U8254 (N_8254,N_8174,N_8158);
nand U8255 (N_8255,N_8186,N_8124);
and U8256 (N_8256,N_8119,N_8113);
nor U8257 (N_8257,N_8135,N_8120);
and U8258 (N_8258,N_8178,N_8142);
nor U8259 (N_8259,N_8129,N_8195);
and U8260 (N_8260,N_8176,N_8107);
nand U8261 (N_8261,N_8151,N_8144);
nand U8262 (N_8262,N_8123,N_8190);
nand U8263 (N_8263,N_8190,N_8161);
nand U8264 (N_8264,N_8138,N_8151);
or U8265 (N_8265,N_8181,N_8100);
nor U8266 (N_8266,N_8175,N_8168);
or U8267 (N_8267,N_8195,N_8138);
and U8268 (N_8268,N_8167,N_8130);
nand U8269 (N_8269,N_8199,N_8132);
nor U8270 (N_8270,N_8131,N_8100);
nand U8271 (N_8271,N_8186,N_8103);
or U8272 (N_8272,N_8184,N_8102);
or U8273 (N_8273,N_8162,N_8101);
or U8274 (N_8274,N_8148,N_8128);
xor U8275 (N_8275,N_8115,N_8145);
nor U8276 (N_8276,N_8168,N_8146);
and U8277 (N_8277,N_8155,N_8179);
or U8278 (N_8278,N_8168,N_8171);
nand U8279 (N_8279,N_8196,N_8107);
and U8280 (N_8280,N_8131,N_8109);
nor U8281 (N_8281,N_8129,N_8130);
nor U8282 (N_8282,N_8156,N_8161);
or U8283 (N_8283,N_8188,N_8163);
and U8284 (N_8284,N_8167,N_8103);
and U8285 (N_8285,N_8114,N_8186);
nand U8286 (N_8286,N_8131,N_8145);
and U8287 (N_8287,N_8190,N_8196);
and U8288 (N_8288,N_8149,N_8190);
nand U8289 (N_8289,N_8171,N_8119);
nand U8290 (N_8290,N_8188,N_8182);
and U8291 (N_8291,N_8167,N_8120);
and U8292 (N_8292,N_8128,N_8166);
or U8293 (N_8293,N_8117,N_8115);
nand U8294 (N_8294,N_8120,N_8107);
and U8295 (N_8295,N_8139,N_8154);
nand U8296 (N_8296,N_8194,N_8112);
nor U8297 (N_8297,N_8152,N_8100);
nor U8298 (N_8298,N_8174,N_8194);
and U8299 (N_8299,N_8128,N_8131);
nand U8300 (N_8300,N_8242,N_8267);
and U8301 (N_8301,N_8254,N_8200);
xor U8302 (N_8302,N_8291,N_8203);
or U8303 (N_8303,N_8271,N_8255);
or U8304 (N_8304,N_8277,N_8223);
nor U8305 (N_8305,N_8263,N_8275);
nor U8306 (N_8306,N_8296,N_8229);
nand U8307 (N_8307,N_8244,N_8286);
nand U8308 (N_8308,N_8202,N_8232);
and U8309 (N_8309,N_8279,N_8220);
and U8310 (N_8310,N_8234,N_8297);
or U8311 (N_8311,N_8241,N_8273);
nor U8312 (N_8312,N_8228,N_8278);
or U8313 (N_8313,N_8290,N_8250);
xnor U8314 (N_8314,N_8249,N_8221);
xor U8315 (N_8315,N_8239,N_8212);
nor U8316 (N_8316,N_8287,N_8245);
nor U8317 (N_8317,N_8206,N_8237);
and U8318 (N_8318,N_8288,N_8257);
nand U8319 (N_8319,N_8292,N_8270);
nor U8320 (N_8320,N_8238,N_8243);
nor U8321 (N_8321,N_8235,N_8224);
nor U8322 (N_8322,N_8240,N_8215);
nor U8323 (N_8323,N_8272,N_8253);
or U8324 (N_8324,N_8230,N_8205);
or U8325 (N_8325,N_8216,N_8285);
nor U8326 (N_8326,N_8207,N_8280);
or U8327 (N_8327,N_8231,N_8226);
nand U8328 (N_8328,N_8265,N_8227);
nor U8329 (N_8329,N_8259,N_8217);
or U8330 (N_8330,N_8233,N_8219);
nor U8331 (N_8331,N_8264,N_8214);
and U8332 (N_8332,N_8262,N_8261);
or U8333 (N_8333,N_8213,N_8222);
and U8334 (N_8334,N_8284,N_8289);
nor U8335 (N_8335,N_8252,N_8293);
nand U8336 (N_8336,N_8218,N_8246);
and U8337 (N_8337,N_8281,N_8298);
nor U8338 (N_8338,N_8247,N_8204);
and U8339 (N_8339,N_8269,N_8208);
or U8340 (N_8340,N_8225,N_8274);
or U8341 (N_8341,N_8268,N_8258);
or U8342 (N_8342,N_8211,N_8236);
and U8343 (N_8343,N_8260,N_8201);
nor U8344 (N_8344,N_8283,N_8294);
and U8345 (N_8345,N_8266,N_8248);
or U8346 (N_8346,N_8282,N_8209);
or U8347 (N_8347,N_8295,N_8251);
or U8348 (N_8348,N_8276,N_8299);
nor U8349 (N_8349,N_8210,N_8256);
nor U8350 (N_8350,N_8279,N_8294);
or U8351 (N_8351,N_8247,N_8217);
nand U8352 (N_8352,N_8226,N_8240);
nand U8353 (N_8353,N_8243,N_8295);
nor U8354 (N_8354,N_8218,N_8244);
and U8355 (N_8355,N_8284,N_8269);
or U8356 (N_8356,N_8229,N_8264);
and U8357 (N_8357,N_8261,N_8268);
nand U8358 (N_8358,N_8259,N_8238);
or U8359 (N_8359,N_8238,N_8204);
nand U8360 (N_8360,N_8270,N_8296);
and U8361 (N_8361,N_8241,N_8219);
and U8362 (N_8362,N_8247,N_8294);
nand U8363 (N_8363,N_8240,N_8293);
nand U8364 (N_8364,N_8266,N_8210);
nor U8365 (N_8365,N_8200,N_8231);
xor U8366 (N_8366,N_8255,N_8257);
nand U8367 (N_8367,N_8208,N_8284);
nor U8368 (N_8368,N_8242,N_8234);
or U8369 (N_8369,N_8256,N_8209);
or U8370 (N_8370,N_8208,N_8223);
nor U8371 (N_8371,N_8252,N_8235);
nand U8372 (N_8372,N_8274,N_8230);
nor U8373 (N_8373,N_8240,N_8261);
and U8374 (N_8374,N_8233,N_8244);
or U8375 (N_8375,N_8274,N_8269);
and U8376 (N_8376,N_8200,N_8215);
or U8377 (N_8377,N_8268,N_8224);
and U8378 (N_8378,N_8201,N_8286);
and U8379 (N_8379,N_8263,N_8270);
xor U8380 (N_8380,N_8293,N_8284);
nor U8381 (N_8381,N_8201,N_8256);
nor U8382 (N_8382,N_8216,N_8280);
nand U8383 (N_8383,N_8297,N_8249);
or U8384 (N_8384,N_8240,N_8200);
and U8385 (N_8385,N_8213,N_8232);
nor U8386 (N_8386,N_8220,N_8260);
nand U8387 (N_8387,N_8213,N_8286);
nand U8388 (N_8388,N_8266,N_8219);
nor U8389 (N_8389,N_8208,N_8241);
nand U8390 (N_8390,N_8281,N_8265);
nand U8391 (N_8391,N_8294,N_8234);
or U8392 (N_8392,N_8258,N_8291);
xor U8393 (N_8393,N_8229,N_8259);
or U8394 (N_8394,N_8201,N_8288);
nand U8395 (N_8395,N_8293,N_8232);
nand U8396 (N_8396,N_8281,N_8205);
nand U8397 (N_8397,N_8206,N_8202);
nand U8398 (N_8398,N_8225,N_8266);
and U8399 (N_8399,N_8224,N_8247);
and U8400 (N_8400,N_8347,N_8398);
and U8401 (N_8401,N_8383,N_8330);
xor U8402 (N_8402,N_8389,N_8374);
and U8403 (N_8403,N_8328,N_8326);
nand U8404 (N_8404,N_8363,N_8351);
or U8405 (N_8405,N_8341,N_8364);
or U8406 (N_8406,N_8339,N_8302);
nor U8407 (N_8407,N_8349,N_8353);
or U8408 (N_8408,N_8336,N_8392);
nor U8409 (N_8409,N_8354,N_8399);
or U8410 (N_8410,N_8306,N_8322);
or U8411 (N_8411,N_8385,N_8338);
nor U8412 (N_8412,N_8331,N_8321);
and U8413 (N_8413,N_8360,N_8387);
or U8414 (N_8414,N_8344,N_8345);
nand U8415 (N_8415,N_8355,N_8388);
nand U8416 (N_8416,N_8380,N_8396);
nor U8417 (N_8417,N_8348,N_8350);
xnor U8418 (N_8418,N_8371,N_8319);
nand U8419 (N_8419,N_8335,N_8368);
or U8420 (N_8420,N_8362,N_8369);
nor U8421 (N_8421,N_8303,N_8390);
and U8422 (N_8422,N_8300,N_8397);
xor U8423 (N_8423,N_8373,N_8367);
nor U8424 (N_8424,N_8393,N_8308);
nor U8425 (N_8425,N_8394,N_8370);
nor U8426 (N_8426,N_8358,N_8313);
nor U8427 (N_8427,N_8327,N_8312);
nor U8428 (N_8428,N_8384,N_8359);
nor U8429 (N_8429,N_8337,N_8386);
nand U8430 (N_8430,N_8332,N_8379);
nor U8431 (N_8431,N_8391,N_8310);
nor U8432 (N_8432,N_8301,N_8340);
and U8433 (N_8433,N_8304,N_8323);
and U8434 (N_8434,N_8334,N_8317);
nand U8435 (N_8435,N_8365,N_8372);
nand U8436 (N_8436,N_8356,N_8342);
nor U8437 (N_8437,N_8357,N_8346);
and U8438 (N_8438,N_8377,N_8352);
or U8439 (N_8439,N_8366,N_8329);
or U8440 (N_8440,N_8316,N_8311);
and U8441 (N_8441,N_8376,N_8307);
nor U8442 (N_8442,N_8315,N_8320);
or U8443 (N_8443,N_8314,N_8375);
nor U8444 (N_8444,N_8305,N_8361);
nand U8445 (N_8445,N_8318,N_8343);
or U8446 (N_8446,N_8324,N_8381);
nand U8447 (N_8447,N_8333,N_8325);
and U8448 (N_8448,N_8382,N_8395);
nand U8449 (N_8449,N_8378,N_8309);
nor U8450 (N_8450,N_8381,N_8320);
nand U8451 (N_8451,N_8308,N_8365);
or U8452 (N_8452,N_8363,N_8306);
or U8453 (N_8453,N_8384,N_8321);
or U8454 (N_8454,N_8316,N_8307);
and U8455 (N_8455,N_8301,N_8373);
nor U8456 (N_8456,N_8396,N_8369);
nor U8457 (N_8457,N_8312,N_8349);
and U8458 (N_8458,N_8328,N_8325);
nor U8459 (N_8459,N_8338,N_8376);
or U8460 (N_8460,N_8300,N_8306);
nand U8461 (N_8461,N_8352,N_8386);
or U8462 (N_8462,N_8335,N_8365);
or U8463 (N_8463,N_8342,N_8334);
nor U8464 (N_8464,N_8364,N_8351);
nor U8465 (N_8465,N_8353,N_8334);
and U8466 (N_8466,N_8306,N_8368);
nand U8467 (N_8467,N_8356,N_8392);
or U8468 (N_8468,N_8322,N_8397);
nand U8469 (N_8469,N_8317,N_8358);
nand U8470 (N_8470,N_8392,N_8385);
or U8471 (N_8471,N_8302,N_8388);
nand U8472 (N_8472,N_8337,N_8304);
and U8473 (N_8473,N_8311,N_8314);
and U8474 (N_8474,N_8301,N_8303);
nor U8475 (N_8475,N_8301,N_8366);
or U8476 (N_8476,N_8389,N_8344);
and U8477 (N_8477,N_8381,N_8372);
nor U8478 (N_8478,N_8376,N_8345);
nor U8479 (N_8479,N_8391,N_8380);
nand U8480 (N_8480,N_8379,N_8357);
nor U8481 (N_8481,N_8306,N_8337);
nand U8482 (N_8482,N_8361,N_8367);
nand U8483 (N_8483,N_8314,N_8317);
and U8484 (N_8484,N_8300,N_8352);
nand U8485 (N_8485,N_8390,N_8310);
nand U8486 (N_8486,N_8369,N_8341);
nand U8487 (N_8487,N_8301,N_8309);
and U8488 (N_8488,N_8371,N_8394);
nand U8489 (N_8489,N_8379,N_8334);
nand U8490 (N_8490,N_8334,N_8329);
nand U8491 (N_8491,N_8326,N_8354);
nand U8492 (N_8492,N_8370,N_8304);
nand U8493 (N_8493,N_8311,N_8399);
and U8494 (N_8494,N_8329,N_8382);
nand U8495 (N_8495,N_8357,N_8373);
or U8496 (N_8496,N_8310,N_8382);
and U8497 (N_8497,N_8394,N_8302);
nand U8498 (N_8498,N_8344,N_8378);
nor U8499 (N_8499,N_8390,N_8368);
and U8500 (N_8500,N_8421,N_8435);
or U8501 (N_8501,N_8403,N_8433);
and U8502 (N_8502,N_8470,N_8441);
xor U8503 (N_8503,N_8464,N_8465);
and U8504 (N_8504,N_8482,N_8492);
nor U8505 (N_8505,N_8494,N_8461);
and U8506 (N_8506,N_8451,N_8444);
and U8507 (N_8507,N_8424,N_8469);
or U8508 (N_8508,N_8434,N_8453);
and U8509 (N_8509,N_8497,N_8449);
and U8510 (N_8510,N_8445,N_8430);
nor U8511 (N_8511,N_8418,N_8466);
and U8512 (N_8512,N_8416,N_8417);
nor U8513 (N_8513,N_8407,N_8432);
or U8514 (N_8514,N_8414,N_8411);
nand U8515 (N_8515,N_8485,N_8426);
and U8516 (N_8516,N_8436,N_8431);
nor U8517 (N_8517,N_8442,N_8499);
or U8518 (N_8518,N_8439,N_8456);
nand U8519 (N_8519,N_8415,N_8491);
or U8520 (N_8520,N_8475,N_8462);
and U8521 (N_8521,N_8401,N_8472);
nor U8522 (N_8522,N_8458,N_8468);
or U8523 (N_8523,N_8446,N_8425);
nor U8524 (N_8524,N_8438,N_8473);
xor U8525 (N_8525,N_8454,N_8447);
and U8526 (N_8526,N_8413,N_8474);
or U8527 (N_8527,N_8408,N_8423);
or U8528 (N_8528,N_8481,N_8483);
or U8529 (N_8529,N_8402,N_8459);
nand U8530 (N_8530,N_8488,N_8489);
nor U8531 (N_8531,N_8467,N_8427);
nor U8532 (N_8532,N_8463,N_8428);
and U8533 (N_8533,N_8412,N_8471);
nor U8534 (N_8534,N_8419,N_8495);
and U8535 (N_8535,N_8404,N_8410);
or U8536 (N_8536,N_8422,N_8486);
nor U8537 (N_8537,N_8450,N_8409);
nand U8538 (N_8538,N_8477,N_8437);
or U8539 (N_8539,N_8479,N_8452);
and U8540 (N_8540,N_8493,N_8448);
and U8541 (N_8541,N_8476,N_8490);
nand U8542 (N_8542,N_8478,N_8457);
or U8543 (N_8543,N_8440,N_8405);
or U8544 (N_8544,N_8487,N_8406);
nor U8545 (N_8545,N_8400,N_8455);
nand U8546 (N_8546,N_8420,N_8496);
and U8547 (N_8547,N_8443,N_8460);
nor U8548 (N_8548,N_8484,N_8480);
or U8549 (N_8549,N_8429,N_8498);
nand U8550 (N_8550,N_8443,N_8450);
and U8551 (N_8551,N_8460,N_8445);
xor U8552 (N_8552,N_8432,N_8476);
and U8553 (N_8553,N_8492,N_8490);
nor U8554 (N_8554,N_8408,N_8471);
and U8555 (N_8555,N_8413,N_8491);
and U8556 (N_8556,N_8413,N_8443);
nor U8557 (N_8557,N_8428,N_8484);
nor U8558 (N_8558,N_8441,N_8475);
nor U8559 (N_8559,N_8423,N_8437);
nand U8560 (N_8560,N_8419,N_8417);
nand U8561 (N_8561,N_8477,N_8458);
nor U8562 (N_8562,N_8439,N_8437);
nand U8563 (N_8563,N_8432,N_8404);
or U8564 (N_8564,N_8401,N_8468);
or U8565 (N_8565,N_8493,N_8440);
or U8566 (N_8566,N_8432,N_8448);
or U8567 (N_8567,N_8415,N_8436);
and U8568 (N_8568,N_8465,N_8477);
or U8569 (N_8569,N_8481,N_8428);
nand U8570 (N_8570,N_8418,N_8427);
nor U8571 (N_8571,N_8437,N_8400);
and U8572 (N_8572,N_8414,N_8442);
and U8573 (N_8573,N_8466,N_8485);
or U8574 (N_8574,N_8439,N_8415);
nor U8575 (N_8575,N_8400,N_8482);
and U8576 (N_8576,N_8402,N_8498);
and U8577 (N_8577,N_8455,N_8482);
nand U8578 (N_8578,N_8430,N_8410);
or U8579 (N_8579,N_8443,N_8406);
or U8580 (N_8580,N_8473,N_8471);
nor U8581 (N_8581,N_8479,N_8493);
and U8582 (N_8582,N_8470,N_8477);
nand U8583 (N_8583,N_8478,N_8489);
nand U8584 (N_8584,N_8440,N_8459);
nor U8585 (N_8585,N_8436,N_8414);
or U8586 (N_8586,N_8416,N_8476);
nor U8587 (N_8587,N_8419,N_8486);
and U8588 (N_8588,N_8455,N_8408);
and U8589 (N_8589,N_8480,N_8422);
and U8590 (N_8590,N_8474,N_8410);
nor U8591 (N_8591,N_8402,N_8424);
nand U8592 (N_8592,N_8470,N_8418);
nor U8593 (N_8593,N_8484,N_8440);
and U8594 (N_8594,N_8408,N_8453);
or U8595 (N_8595,N_8482,N_8442);
and U8596 (N_8596,N_8480,N_8451);
nor U8597 (N_8597,N_8483,N_8406);
nand U8598 (N_8598,N_8452,N_8469);
nor U8599 (N_8599,N_8429,N_8468);
nand U8600 (N_8600,N_8518,N_8580);
nand U8601 (N_8601,N_8527,N_8504);
nand U8602 (N_8602,N_8555,N_8502);
nand U8603 (N_8603,N_8514,N_8584);
and U8604 (N_8604,N_8548,N_8594);
nor U8605 (N_8605,N_8576,N_8537);
and U8606 (N_8606,N_8585,N_8558);
and U8607 (N_8607,N_8579,N_8525);
and U8608 (N_8608,N_8541,N_8581);
nand U8609 (N_8609,N_8590,N_8534);
or U8610 (N_8610,N_8597,N_8591);
xor U8611 (N_8611,N_8512,N_8589);
and U8612 (N_8612,N_8539,N_8513);
nor U8613 (N_8613,N_8592,N_8554);
and U8614 (N_8614,N_8562,N_8508);
or U8615 (N_8615,N_8578,N_8533);
nand U8616 (N_8616,N_8530,N_8522);
nand U8617 (N_8617,N_8500,N_8549);
nand U8618 (N_8618,N_8511,N_8507);
nor U8619 (N_8619,N_8536,N_8598);
and U8620 (N_8620,N_8552,N_8546);
and U8621 (N_8621,N_8528,N_8599);
nor U8622 (N_8622,N_8595,N_8559);
nand U8623 (N_8623,N_8517,N_8532);
nand U8624 (N_8624,N_8515,N_8545);
and U8625 (N_8625,N_8557,N_8543);
and U8626 (N_8626,N_8501,N_8540);
or U8627 (N_8627,N_8572,N_8587);
and U8628 (N_8628,N_8566,N_8571);
nor U8629 (N_8629,N_8542,N_8596);
and U8630 (N_8630,N_8563,N_8506);
nor U8631 (N_8631,N_8535,N_8538);
nand U8632 (N_8632,N_8575,N_8553);
nor U8633 (N_8633,N_8586,N_8569);
xor U8634 (N_8634,N_8519,N_8510);
nor U8635 (N_8635,N_8524,N_8544);
xnor U8636 (N_8636,N_8573,N_8529);
nor U8637 (N_8637,N_8588,N_8550);
and U8638 (N_8638,N_8577,N_8551);
or U8639 (N_8639,N_8564,N_8570);
nand U8640 (N_8640,N_8521,N_8593);
and U8641 (N_8641,N_8516,N_8574);
and U8642 (N_8642,N_8509,N_8520);
and U8643 (N_8643,N_8583,N_8523);
nor U8644 (N_8644,N_8556,N_8561);
or U8645 (N_8645,N_8560,N_8531);
or U8646 (N_8646,N_8526,N_8565);
nor U8647 (N_8647,N_8505,N_8503);
nor U8648 (N_8648,N_8567,N_8568);
or U8649 (N_8649,N_8547,N_8582);
nand U8650 (N_8650,N_8559,N_8541);
xor U8651 (N_8651,N_8512,N_8553);
and U8652 (N_8652,N_8587,N_8591);
nor U8653 (N_8653,N_8553,N_8532);
or U8654 (N_8654,N_8570,N_8571);
and U8655 (N_8655,N_8564,N_8535);
nand U8656 (N_8656,N_8568,N_8575);
nor U8657 (N_8657,N_8527,N_8544);
nor U8658 (N_8658,N_8524,N_8572);
and U8659 (N_8659,N_8500,N_8591);
nand U8660 (N_8660,N_8517,N_8588);
or U8661 (N_8661,N_8574,N_8515);
or U8662 (N_8662,N_8532,N_8579);
nor U8663 (N_8663,N_8536,N_8503);
nor U8664 (N_8664,N_8578,N_8510);
and U8665 (N_8665,N_8500,N_8581);
nand U8666 (N_8666,N_8528,N_8534);
nor U8667 (N_8667,N_8539,N_8543);
nor U8668 (N_8668,N_8562,N_8563);
and U8669 (N_8669,N_8500,N_8525);
nand U8670 (N_8670,N_8561,N_8532);
nand U8671 (N_8671,N_8576,N_8551);
and U8672 (N_8672,N_8539,N_8550);
nand U8673 (N_8673,N_8567,N_8548);
nor U8674 (N_8674,N_8598,N_8506);
or U8675 (N_8675,N_8545,N_8541);
nand U8676 (N_8676,N_8540,N_8535);
and U8677 (N_8677,N_8548,N_8523);
nand U8678 (N_8678,N_8531,N_8518);
nand U8679 (N_8679,N_8573,N_8534);
nand U8680 (N_8680,N_8525,N_8519);
or U8681 (N_8681,N_8583,N_8506);
and U8682 (N_8682,N_8524,N_8520);
nand U8683 (N_8683,N_8549,N_8585);
or U8684 (N_8684,N_8543,N_8507);
and U8685 (N_8685,N_8564,N_8558);
and U8686 (N_8686,N_8508,N_8587);
nor U8687 (N_8687,N_8519,N_8542);
nor U8688 (N_8688,N_8590,N_8598);
nand U8689 (N_8689,N_8593,N_8580);
nor U8690 (N_8690,N_8573,N_8518);
nor U8691 (N_8691,N_8557,N_8563);
nand U8692 (N_8692,N_8596,N_8510);
and U8693 (N_8693,N_8574,N_8555);
xor U8694 (N_8694,N_8593,N_8514);
nor U8695 (N_8695,N_8580,N_8541);
nor U8696 (N_8696,N_8537,N_8546);
nand U8697 (N_8697,N_8507,N_8584);
nor U8698 (N_8698,N_8505,N_8535);
and U8699 (N_8699,N_8534,N_8505);
nand U8700 (N_8700,N_8628,N_8670);
and U8701 (N_8701,N_8629,N_8631);
and U8702 (N_8702,N_8633,N_8655);
and U8703 (N_8703,N_8681,N_8672);
and U8704 (N_8704,N_8667,N_8649);
and U8705 (N_8705,N_8626,N_8678);
and U8706 (N_8706,N_8627,N_8620);
nor U8707 (N_8707,N_8635,N_8663);
nor U8708 (N_8708,N_8664,N_8619);
and U8709 (N_8709,N_8660,N_8691);
nand U8710 (N_8710,N_8698,N_8695);
and U8711 (N_8711,N_8657,N_8694);
or U8712 (N_8712,N_8675,N_8608);
or U8713 (N_8713,N_8600,N_8682);
and U8714 (N_8714,N_8650,N_8644);
and U8715 (N_8715,N_8640,N_8622);
or U8716 (N_8716,N_8632,N_8683);
nand U8717 (N_8717,N_8686,N_8605);
or U8718 (N_8718,N_8659,N_8636);
or U8719 (N_8719,N_8680,N_8662);
and U8720 (N_8720,N_8647,N_8624);
or U8721 (N_8721,N_8616,N_8641);
nand U8722 (N_8722,N_8625,N_8639);
nand U8723 (N_8723,N_8614,N_8689);
and U8724 (N_8724,N_8658,N_8606);
and U8725 (N_8725,N_8602,N_8654);
nand U8726 (N_8726,N_8688,N_8634);
nor U8727 (N_8727,N_8601,N_8646);
and U8728 (N_8728,N_8656,N_8699);
nor U8729 (N_8729,N_8604,N_8603);
nand U8730 (N_8730,N_8612,N_8697);
and U8731 (N_8731,N_8693,N_8669);
and U8732 (N_8732,N_8623,N_8651);
and U8733 (N_8733,N_8673,N_8615);
nor U8734 (N_8734,N_8611,N_8665);
and U8735 (N_8735,N_8685,N_8645);
or U8736 (N_8736,N_8642,N_8638);
or U8737 (N_8737,N_8676,N_8652);
and U8738 (N_8738,N_8671,N_8692);
nand U8739 (N_8739,N_8637,N_8684);
or U8740 (N_8740,N_8674,N_8668);
and U8741 (N_8741,N_8621,N_8648);
nor U8742 (N_8742,N_8687,N_8630);
and U8743 (N_8743,N_8653,N_8610);
or U8744 (N_8744,N_8661,N_8643);
nor U8745 (N_8745,N_8618,N_8617);
nand U8746 (N_8746,N_8696,N_8679);
nand U8747 (N_8747,N_8666,N_8613);
nor U8748 (N_8748,N_8607,N_8677);
nor U8749 (N_8749,N_8690,N_8609);
nor U8750 (N_8750,N_8657,N_8600);
or U8751 (N_8751,N_8610,N_8621);
and U8752 (N_8752,N_8657,N_8618);
nor U8753 (N_8753,N_8658,N_8663);
and U8754 (N_8754,N_8601,N_8689);
or U8755 (N_8755,N_8603,N_8639);
or U8756 (N_8756,N_8686,N_8649);
and U8757 (N_8757,N_8621,N_8653);
nor U8758 (N_8758,N_8632,N_8602);
or U8759 (N_8759,N_8630,N_8631);
nor U8760 (N_8760,N_8695,N_8692);
and U8761 (N_8761,N_8667,N_8632);
nor U8762 (N_8762,N_8699,N_8662);
and U8763 (N_8763,N_8619,N_8638);
nand U8764 (N_8764,N_8682,N_8651);
nand U8765 (N_8765,N_8602,N_8647);
nor U8766 (N_8766,N_8699,N_8666);
nor U8767 (N_8767,N_8685,N_8625);
and U8768 (N_8768,N_8633,N_8601);
nor U8769 (N_8769,N_8672,N_8640);
and U8770 (N_8770,N_8697,N_8614);
nand U8771 (N_8771,N_8678,N_8681);
and U8772 (N_8772,N_8662,N_8677);
nand U8773 (N_8773,N_8602,N_8680);
nand U8774 (N_8774,N_8693,N_8676);
or U8775 (N_8775,N_8642,N_8644);
xnor U8776 (N_8776,N_8684,N_8624);
nand U8777 (N_8777,N_8637,N_8689);
or U8778 (N_8778,N_8675,N_8620);
nand U8779 (N_8779,N_8698,N_8669);
nand U8780 (N_8780,N_8653,N_8693);
or U8781 (N_8781,N_8652,N_8643);
nand U8782 (N_8782,N_8633,N_8629);
and U8783 (N_8783,N_8646,N_8604);
xor U8784 (N_8784,N_8694,N_8608);
or U8785 (N_8785,N_8697,N_8687);
nor U8786 (N_8786,N_8608,N_8638);
nand U8787 (N_8787,N_8686,N_8606);
or U8788 (N_8788,N_8635,N_8696);
nor U8789 (N_8789,N_8644,N_8677);
nand U8790 (N_8790,N_8633,N_8652);
nand U8791 (N_8791,N_8667,N_8660);
nand U8792 (N_8792,N_8683,N_8606);
nand U8793 (N_8793,N_8687,N_8637);
nand U8794 (N_8794,N_8629,N_8617);
nor U8795 (N_8795,N_8639,N_8657);
nand U8796 (N_8796,N_8656,N_8677);
nand U8797 (N_8797,N_8645,N_8614);
nand U8798 (N_8798,N_8614,N_8684);
nand U8799 (N_8799,N_8684,N_8681);
or U8800 (N_8800,N_8795,N_8772);
nand U8801 (N_8801,N_8764,N_8726);
nor U8802 (N_8802,N_8720,N_8787);
and U8803 (N_8803,N_8760,N_8789);
nor U8804 (N_8804,N_8700,N_8728);
nor U8805 (N_8805,N_8707,N_8703);
nand U8806 (N_8806,N_8775,N_8706);
or U8807 (N_8807,N_8753,N_8763);
nand U8808 (N_8808,N_8732,N_8702);
or U8809 (N_8809,N_8729,N_8757);
or U8810 (N_8810,N_8731,N_8759);
xnor U8811 (N_8811,N_8738,N_8755);
nand U8812 (N_8812,N_8745,N_8774);
nand U8813 (N_8813,N_8712,N_8784);
nor U8814 (N_8814,N_8723,N_8754);
nand U8815 (N_8815,N_8735,N_8771);
or U8816 (N_8816,N_8744,N_8756);
nand U8817 (N_8817,N_8780,N_8783);
and U8818 (N_8818,N_8779,N_8737);
nor U8819 (N_8819,N_8768,N_8746);
nand U8820 (N_8820,N_8721,N_8713);
or U8821 (N_8821,N_8773,N_8796);
or U8822 (N_8822,N_8714,N_8743);
and U8823 (N_8823,N_8769,N_8750);
nand U8824 (N_8824,N_8705,N_8777);
or U8825 (N_8825,N_8798,N_8766);
or U8826 (N_8826,N_8724,N_8782);
nor U8827 (N_8827,N_8749,N_8797);
and U8828 (N_8828,N_8709,N_8733);
nor U8829 (N_8829,N_8727,N_8761);
nand U8830 (N_8830,N_8718,N_8711);
or U8831 (N_8831,N_8719,N_8762);
or U8832 (N_8832,N_8770,N_8791);
and U8833 (N_8833,N_8751,N_8701);
and U8834 (N_8834,N_8799,N_8740);
or U8835 (N_8835,N_8788,N_8715);
or U8836 (N_8836,N_8741,N_8722);
xnor U8837 (N_8837,N_8752,N_8717);
nand U8838 (N_8838,N_8767,N_8704);
nand U8839 (N_8839,N_8794,N_8793);
nand U8840 (N_8840,N_8765,N_8778);
or U8841 (N_8841,N_8708,N_8792);
xor U8842 (N_8842,N_8785,N_8730);
or U8843 (N_8843,N_8725,N_8781);
or U8844 (N_8844,N_8736,N_8776);
nand U8845 (N_8845,N_8734,N_8747);
nor U8846 (N_8846,N_8742,N_8790);
nand U8847 (N_8847,N_8758,N_8739);
nand U8848 (N_8848,N_8710,N_8786);
and U8849 (N_8849,N_8716,N_8748);
nand U8850 (N_8850,N_8770,N_8772);
nand U8851 (N_8851,N_8731,N_8774);
or U8852 (N_8852,N_8722,N_8754);
and U8853 (N_8853,N_8729,N_8746);
nor U8854 (N_8854,N_8794,N_8754);
nor U8855 (N_8855,N_8799,N_8736);
and U8856 (N_8856,N_8753,N_8740);
and U8857 (N_8857,N_8704,N_8784);
or U8858 (N_8858,N_8757,N_8706);
or U8859 (N_8859,N_8755,N_8790);
nand U8860 (N_8860,N_8764,N_8725);
nor U8861 (N_8861,N_8731,N_8778);
nor U8862 (N_8862,N_8724,N_8723);
nor U8863 (N_8863,N_8752,N_8760);
nand U8864 (N_8864,N_8720,N_8763);
or U8865 (N_8865,N_8728,N_8754);
nand U8866 (N_8866,N_8729,N_8739);
and U8867 (N_8867,N_8770,N_8709);
nor U8868 (N_8868,N_8729,N_8717);
xnor U8869 (N_8869,N_8776,N_8715);
nor U8870 (N_8870,N_8712,N_8711);
and U8871 (N_8871,N_8746,N_8725);
xor U8872 (N_8872,N_8776,N_8712);
and U8873 (N_8873,N_8798,N_8775);
nor U8874 (N_8874,N_8741,N_8784);
nor U8875 (N_8875,N_8744,N_8798);
and U8876 (N_8876,N_8779,N_8720);
nand U8877 (N_8877,N_8750,N_8735);
nand U8878 (N_8878,N_8737,N_8754);
nand U8879 (N_8879,N_8736,N_8798);
and U8880 (N_8880,N_8700,N_8747);
nand U8881 (N_8881,N_8738,N_8773);
nor U8882 (N_8882,N_8781,N_8761);
or U8883 (N_8883,N_8716,N_8753);
nor U8884 (N_8884,N_8744,N_8762);
nor U8885 (N_8885,N_8783,N_8709);
or U8886 (N_8886,N_8764,N_8741);
nor U8887 (N_8887,N_8715,N_8775);
nor U8888 (N_8888,N_8742,N_8731);
and U8889 (N_8889,N_8720,N_8788);
and U8890 (N_8890,N_8733,N_8713);
and U8891 (N_8891,N_8779,N_8722);
and U8892 (N_8892,N_8724,N_8702);
nor U8893 (N_8893,N_8785,N_8753);
xor U8894 (N_8894,N_8742,N_8767);
nand U8895 (N_8895,N_8785,N_8738);
or U8896 (N_8896,N_8752,N_8759);
and U8897 (N_8897,N_8715,N_8716);
nor U8898 (N_8898,N_8737,N_8792);
nand U8899 (N_8899,N_8754,N_8786);
or U8900 (N_8900,N_8821,N_8877);
or U8901 (N_8901,N_8862,N_8885);
nand U8902 (N_8902,N_8846,N_8816);
or U8903 (N_8903,N_8853,N_8808);
or U8904 (N_8904,N_8878,N_8888);
nand U8905 (N_8905,N_8887,N_8873);
and U8906 (N_8906,N_8802,N_8811);
nor U8907 (N_8907,N_8832,N_8855);
nand U8908 (N_8908,N_8892,N_8894);
nor U8909 (N_8909,N_8891,N_8874);
nor U8910 (N_8910,N_8897,N_8817);
or U8911 (N_8911,N_8857,N_8809);
or U8912 (N_8912,N_8850,N_8812);
nand U8913 (N_8913,N_8801,N_8818);
nor U8914 (N_8914,N_8860,N_8819);
and U8915 (N_8915,N_8839,N_8833);
nor U8916 (N_8916,N_8814,N_8835);
nand U8917 (N_8917,N_8867,N_8830);
and U8918 (N_8918,N_8806,N_8889);
nor U8919 (N_8919,N_8858,N_8848);
and U8920 (N_8920,N_8856,N_8813);
and U8921 (N_8921,N_8896,N_8803);
and U8922 (N_8922,N_8876,N_8810);
nand U8923 (N_8923,N_8820,N_8845);
nor U8924 (N_8924,N_8834,N_8893);
nand U8925 (N_8925,N_8838,N_8868);
nand U8926 (N_8926,N_8842,N_8840);
and U8927 (N_8927,N_8883,N_8831);
nor U8928 (N_8928,N_8837,N_8805);
and U8929 (N_8929,N_8815,N_8826);
or U8930 (N_8930,N_8865,N_8895);
nand U8931 (N_8931,N_8843,N_8804);
nor U8932 (N_8932,N_8841,N_8824);
or U8933 (N_8933,N_8851,N_8854);
or U8934 (N_8934,N_8886,N_8864);
nor U8935 (N_8935,N_8825,N_8882);
xnor U8936 (N_8936,N_8844,N_8861);
and U8937 (N_8937,N_8823,N_8849);
and U8938 (N_8938,N_8890,N_8822);
or U8939 (N_8939,N_8828,N_8807);
or U8940 (N_8940,N_8827,N_8872);
nand U8941 (N_8941,N_8847,N_8899);
and U8942 (N_8942,N_8898,N_8881);
or U8943 (N_8943,N_8875,N_8863);
nand U8944 (N_8944,N_8859,N_8852);
or U8945 (N_8945,N_8879,N_8871);
and U8946 (N_8946,N_8829,N_8884);
nor U8947 (N_8947,N_8800,N_8869);
nor U8948 (N_8948,N_8866,N_8836);
nor U8949 (N_8949,N_8880,N_8870);
nand U8950 (N_8950,N_8851,N_8829);
nand U8951 (N_8951,N_8865,N_8803);
and U8952 (N_8952,N_8830,N_8826);
and U8953 (N_8953,N_8851,N_8886);
and U8954 (N_8954,N_8863,N_8857);
nand U8955 (N_8955,N_8866,N_8879);
nand U8956 (N_8956,N_8842,N_8834);
nor U8957 (N_8957,N_8823,N_8859);
or U8958 (N_8958,N_8876,N_8853);
and U8959 (N_8959,N_8836,N_8885);
and U8960 (N_8960,N_8808,N_8896);
nand U8961 (N_8961,N_8868,N_8856);
nand U8962 (N_8962,N_8805,N_8856);
xnor U8963 (N_8963,N_8871,N_8896);
nor U8964 (N_8964,N_8803,N_8812);
nand U8965 (N_8965,N_8802,N_8899);
nor U8966 (N_8966,N_8864,N_8882);
or U8967 (N_8967,N_8805,N_8890);
nor U8968 (N_8968,N_8889,N_8890);
nand U8969 (N_8969,N_8838,N_8861);
nand U8970 (N_8970,N_8864,N_8855);
nor U8971 (N_8971,N_8881,N_8897);
xor U8972 (N_8972,N_8876,N_8817);
nand U8973 (N_8973,N_8894,N_8891);
nor U8974 (N_8974,N_8810,N_8805);
or U8975 (N_8975,N_8835,N_8837);
and U8976 (N_8976,N_8862,N_8802);
or U8977 (N_8977,N_8829,N_8864);
xnor U8978 (N_8978,N_8829,N_8869);
nand U8979 (N_8979,N_8847,N_8823);
or U8980 (N_8980,N_8875,N_8836);
and U8981 (N_8981,N_8820,N_8824);
nand U8982 (N_8982,N_8840,N_8838);
or U8983 (N_8983,N_8835,N_8834);
and U8984 (N_8984,N_8820,N_8814);
and U8985 (N_8985,N_8832,N_8882);
nor U8986 (N_8986,N_8889,N_8840);
xnor U8987 (N_8987,N_8877,N_8812);
or U8988 (N_8988,N_8812,N_8863);
nor U8989 (N_8989,N_8875,N_8855);
nand U8990 (N_8990,N_8855,N_8883);
nand U8991 (N_8991,N_8820,N_8871);
nor U8992 (N_8992,N_8832,N_8863);
or U8993 (N_8993,N_8858,N_8828);
and U8994 (N_8994,N_8812,N_8851);
or U8995 (N_8995,N_8870,N_8824);
nor U8996 (N_8996,N_8819,N_8834);
nor U8997 (N_8997,N_8867,N_8899);
nor U8998 (N_8998,N_8842,N_8805);
and U8999 (N_8999,N_8846,N_8879);
nor U9000 (N_9000,N_8973,N_8956);
nand U9001 (N_9001,N_8914,N_8949);
and U9002 (N_9002,N_8947,N_8925);
nor U9003 (N_9003,N_8913,N_8951);
nor U9004 (N_9004,N_8910,N_8982);
nand U9005 (N_9005,N_8983,N_8977);
nand U9006 (N_9006,N_8916,N_8954);
or U9007 (N_9007,N_8904,N_8924);
nand U9008 (N_9008,N_8908,N_8919);
and U9009 (N_9009,N_8979,N_8966);
nand U9010 (N_9010,N_8941,N_8959);
or U9011 (N_9011,N_8986,N_8923);
and U9012 (N_9012,N_8975,N_8920);
nor U9013 (N_9013,N_8970,N_8980);
nor U9014 (N_9014,N_8934,N_8961);
nand U9015 (N_9015,N_8939,N_8903);
nor U9016 (N_9016,N_8957,N_8971);
and U9017 (N_9017,N_8928,N_8902);
nand U9018 (N_9018,N_8968,N_8988);
nor U9019 (N_9019,N_8992,N_8995);
nor U9020 (N_9020,N_8993,N_8915);
xnor U9021 (N_9021,N_8972,N_8948);
and U9022 (N_9022,N_8978,N_8953);
or U9023 (N_9023,N_8944,N_8917);
or U9024 (N_9024,N_8985,N_8935);
xor U9025 (N_9025,N_8960,N_8955);
and U9026 (N_9026,N_8952,N_8931);
xor U9027 (N_9027,N_8907,N_8942);
nand U9028 (N_9028,N_8999,N_8963);
or U9029 (N_9029,N_8922,N_8969);
nor U9030 (N_9030,N_8905,N_8990);
nor U9031 (N_9031,N_8946,N_8906);
nor U9032 (N_9032,N_8984,N_8945);
and U9033 (N_9033,N_8938,N_8940);
nand U9034 (N_9034,N_8921,N_8933);
or U9035 (N_9035,N_8943,N_8930);
nand U9036 (N_9036,N_8998,N_8989);
nand U9037 (N_9037,N_8964,N_8950);
xnor U9038 (N_9038,N_8994,N_8911);
nor U9039 (N_9039,N_8965,N_8997);
nand U9040 (N_9040,N_8991,N_8900);
and U9041 (N_9041,N_8937,N_8958);
nor U9042 (N_9042,N_8987,N_8996);
or U9043 (N_9043,N_8912,N_8909);
and U9044 (N_9044,N_8918,N_8926);
and U9045 (N_9045,N_8974,N_8936);
and U9046 (N_9046,N_8901,N_8932);
nor U9047 (N_9047,N_8927,N_8929);
nand U9048 (N_9048,N_8962,N_8981);
nor U9049 (N_9049,N_8976,N_8967);
nor U9050 (N_9050,N_8952,N_8945);
nand U9051 (N_9051,N_8956,N_8957);
nor U9052 (N_9052,N_8924,N_8940);
nor U9053 (N_9053,N_8979,N_8918);
and U9054 (N_9054,N_8934,N_8945);
or U9055 (N_9055,N_8936,N_8917);
or U9056 (N_9056,N_8922,N_8937);
nand U9057 (N_9057,N_8948,N_8963);
or U9058 (N_9058,N_8929,N_8983);
or U9059 (N_9059,N_8974,N_8913);
xnor U9060 (N_9060,N_8934,N_8946);
and U9061 (N_9061,N_8939,N_8907);
and U9062 (N_9062,N_8974,N_8903);
nor U9063 (N_9063,N_8995,N_8936);
nand U9064 (N_9064,N_8991,N_8979);
xor U9065 (N_9065,N_8977,N_8905);
or U9066 (N_9066,N_8938,N_8941);
nor U9067 (N_9067,N_8952,N_8903);
nand U9068 (N_9068,N_8969,N_8961);
nor U9069 (N_9069,N_8916,N_8936);
nand U9070 (N_9070,N_8921,N_8942);
nor U9071 (N_9071,N_8985,N_8952);
and U9072 (N_9072,N_8980,N_8988);
nor U9073 (N_9073,N_8951,N_8909);
nand U9074 (N_9074,N_8989,N_8924);
nand U9075 (N_9075,N_8905,N_8993);
and U9076 (N_9076,N_8958,N_8905);
nor U9077 (N_9077,N_8907,N_8990);
and U9078 (N_9078,N_8915,N_8953);
or U9079 (N_9079,N_8932,N_8925);
xor U9080 (N_9080,N_8970,N_8953);
or U9081 (N_9081,N_8966,N_8937);
or U9082 (N_9082,N_8900,N_8951);
nor U9083 (N_9083,N_8961,N_8913);
or U9084 (N_9084,N_8969,N_8927);
xor U9085 (N_9085,N_8940,N_8978);
nand U9086 (N_9086,N_8966,N_8968);
nor U9087 (N_9087,N_8962,N_8999);
nand U9088 (N_9088,N_8908,N_8918);
nand U9089 (N_9089,N_8981,N_8928);
or U9090 (N_9090,N_8904,N_8914);
nor U9091 (N_9091,N_8915,N_8964);
nor U9092 (N_9092,N_8931,N_8973);
nand U9093 (N_9093,N_8982,N_8967);
or U9094 (N_9094,N_8906,N_8988);
nand U9095 (N_9095,N_8993,N_8926);
nand U9096 (N_9096,N_8934,N_8936);
nand U9097 (N_9097,N_8935,N_8906);
xnor U9098 (N_9098,N_8940,N_8923);
nand U9099 (N_9099,N_8907,N_8987);
nand U9100 (N_9100,N_9052,N_9072);
or U9101 (N_9101,N_9039,N_9035);
and U9102 (N_9102,N_9053,N_9068);
nand U9103 (N_9103,N_9090,N_9060);
or U9104 (N_9104,N_9089,N_9013);
nor U9105 (N_9105,N_9067,N_9044);
or U9106 (N_9106,N_9088,N_9045);
nand U9107 (N_9107,N_9006,N_9064);
nand U9108 (N_9108,N_9071,N_9086);
or U9109 (N_9109,N_9021,N_9020);
nor U9110 (N_9110,N_9092,N_9085);
or U9111 (N_9111,N_9059,N_9023);
and U9112 (N_9112,N_9094,N_9051);
and U9113 (N_9113,N_9015,N_9018);
or U9114 (N_9114,N_9066,N_9058);
or U9115 (N_9115,N_9003,N_9032);
or U9116 (N_9116,N_9076,N_9091);
and U9117 (N_9117,N_9099,N_9030);
and U9118 (N_9118,N_9082,N_9002);
or U9119 (N_9119,N_9070,N_9056);
and U9120 (N_9120,N_9047,N_9087);
xnor U9121 (N_9121,N_9079,N_9012);
or U9122 (N_9122,N_9098,N_9075);
nand U9123 (N_9123,N_9074,N_9000);
or U9124 (N_9124,N_9029,N_9093);
and U9125 (N_9125,N_9024,N_9050);
nand U9126 (N_9126,N_9010,N_9014);
and U9127 (N_9127,N_9065,N_9054);
nand U9128 (N_9128,N_9034,N_9042);
or U9129 (N_9129,N_9084,N_9016);
nand U9130 (N_9130,N_9033,N_9097);
nand U9131 (N_9131,N_9009,N_9046);
nor U9132 (N_9132,N_9049,N_9031);
or U9133 (N_9133,N_9019,N_9057);
or U9134 (N_9134,N_9040,N_9025);
and U9135 (N_9135,N_9004,N_9062);
nor U9136 (N_9136,N_9043,N_9095);
and U9137 (N_9137,N_9096,N_9036);
nor U9138 (N_9138,N_9037,N_9061);
nor U9139 (N_9139,N_9001,N_9028);
or U9140 (N_9140,N_9048,N_9078);
nand U9141 (N_9141,N_9005,N_9081);
nor U9142 (N_9142,N_9038,N_9077);
or U9143 (N_9143,N_9080,N_9026);
or U9144 (N_9144,N_9055,N_9069);
and U9145 (N_9145,N_9008,N_9022);
nand U9146 (N_9146,N_9017,N_9027);
nand U9147 (N_9147,N_9063,N_9011);
and U9148 (N_9148,N_9007,N_9073);
and U9149 (N_9149,N_9041,N_9083);
nand U9150 (N_9150,N_9065,N_9009);
or U9151 (N_9151,N_9045,N_9046);
nor U9152 (N_9152,N_9004,N_9038);
or U9153 (N_9153,N_9095,N_9096);
nand U9154 (N_9154,N_9003,N_9041);
or U9155 (N_9155,N_9076,N_9050);
and U9156 (N_9156,N_9009,N_9007);
nor U9157 (N_9157,N_9016,N_9024);
and U9158 (N_9158,N_9070,N_9027);
xnor U9159 (N_9159,N_9024,N_9071);
nand U9160 (N_9160,N_9057,N_9020);
xor U9161 (N_9161,N_9017,N_9093);
and U9162 (N_9162,N_9063,N_9088);
and U9163 (N_9163,N_9084,N_9011);
nor U9164 (N_9164,N_9015,N_9072);
nor U9165 (N_9165,N_9037,N_9085);
nand U9166 (N_9166,N_9024,N_9095);
and U9167 (N_9167,N_9006,N_9041);
or U9168 (N_9168,N_9039,N_9089);
nand U9169 (N_9169,N_9005,N_9069);
nand U9170 (N_9170,N_9018,N_9081);
or U9171 (N_9171,N_9035,N_9015);
nand U9172 (N_9172,N_9046,N_9058);
nand U9173 (N_9173,N_9080,N_9033);
or U9174 (N_9174,N_9045,N_9008);
or U9175 (N_9175,N_9061,N_9022);
or U9176 (N_9176,N_9072,N_9038);
and U9177 (N_9177,N_9082,N_9078);
nand U9178 (N_9178,N_9010,N_9065);
nor U9179 (N_9179,N_9011,N_9070);
or U9180 (N_9180,N_9082,N_9070);
or U9181 (N_9181,N_9015,N_9034);
and U9182 (N_9182,N_9011,N_9097);
or U9183 (N_9183,N_9061,N_9066);
nand U9184 (N_9184,N_9092,N_9005);
and U9185 (N_9185,N_9071,N_9041);
nor U9186 (N_9186,N_9001,N_9045);
or U9187 (N_9187,N_9067,N_9019);
nand U9188 (N_9188,N_9030,N_9087);
and U9189 (N_9189,N_9081,N_9045);
and U9190 (N_9190,N_9096,N_9064);
nor U9191 (N_9191,N_9046,N_9020);
nor U9192 (N_9192,N_9031,N_9066);
nor U9193 (N_9193,N_9060,N_9067);
or U9194 (N_9194,N_9043,N_9041);
or U9195 (N_9195,N_9066,N_9040);
nand U9196 (N_9196,N_9018,N_9086);
nor U9197 (N_9197,N_9035,N_9075);
nor U9198 (N_9198,N_9056,N_9061);
or U9199 (N_9199,N_9027,N_9092);
nand U9200 (N_9200,N_9186,N_9177);
or U9201 (N_9201,N_9136,N_9182);
or U9202 (N_9202,N_9125,N_9145);
or U9203 (N_9203,N_9158,N_9105);
nor U9204 (N_9204,N_9174,N_9110);
nand U9205 (N_9205,N_9152,N_9168);
or U9206 (N_9206,N_9199,N_9161);
nand U9207 (N_9207,N_9103,N_9123);
or U9208 (N_9208,N_9102,N_9162);
and U9209 (N_9209,N_9196,N_9115);
nand U9210 (N_9210,N_9189,N_9148);
and U9211 (N_9211,N_9181,N_9124);
and U9212 (N_9212,N_9131,N_9160);
nor U9213 (N_9213,N_9141,N_9137);
nand U9214 (N_9214,N_9116,N_9185);
and U9215 (N_9215,N_9153,N_9172);
or U9216 (N_9216,N_9139,N_9198);
nor U9217 (N_9217,N_9119,N_9173);
nor U9218 (N_9218,N_9171,N_9100);
nand U9219 (N_9219,N_9122,N_9118);
nor U9220 (N_9220,N_9184,N_9166);
and U9221 (N_9221,N_9146,N_9191);
nor U9222 (N_9222,N_9138,N_9121);
nor U9223 (N_9223,N_9150,N_9188);
nand U9224 (N_9224,N_9106,N_9128);
or U9225 (N_9225,N_9135,N_9154);
nand U9226 (N_9226,N_9197,N_9126);
or U9227 (N_9227,N_9194,N_9190);
nor U9228 (N_9228,N_9134,N_9193);
and U9229 (N_9229,N_9112,N_9157);
nand U9230 (N_9230,N_9117,N_9169);
nand U9231 (N_9231,N_9170,N_9143);
nand U9232 (N_9232,N_9159,N_9178);
nor U9233 (N_9233,N_9144,N_9180);
and U9234 (N_9234,N_9113,N_9142);
or U9235 (N_9235,N_9114,N_9195);
and U9236 (N_9236,N_9127,N_9151);
nor U9237 (N_9237,N_9107,N_9130);
xnor U9238 (N_9238,N_9147,N_9101);
and U9239 (N_9239,N_9156,N_9108);
or U9240 (N_9240,N_9163,N_9167);
or U9241 (N_9241,N_9129,N_9140);
or U9242 (N_9242,N_9120,N_9187);
or U9243 (N_9243,N_9104,N_9179);
nand U9244 (N_9244,N_9111,N_9192);
or U9245 (N_9245,N_9149,N_9164);
or U9246 (N_9246,N_9165,N_9132);
or U9247 (N_9247,N_9175,N_9183);
and U9248 (N_9248,N_9155,N_9109);
and U9249 (N_9249,N_9133,N_9176);
and U9250 (N_9250,N_9193,N_9144);
nand U9251 (N_9251,N_9104,N_9182);
and U9252 (N_9252,N_9160,N_9112);
nand U9253 (N_9253,N_9191,N_9156);
nand U9254 (N_9254,N_9103,N_9161);
nand U9255 (N_9255,N_9132,N_9118);
xnor U9256 (N_9256,N_9139,N_9159);
and U9257 (N_9257,N_9102,N_9100);
nand U9258 (N_9258,N_9145,N_9191);
nor U9259 (N_9259,N_9138,N_9103);
nor U9260 (N_9260,N_9100,N_9104);
nand U9261 (N_9261,N_9161,N_9182);
nand U9262 (N_9262,N_9173,N_9134);
nor U9263 (N_9263,N_9164,N_9137);
and U9264 (N_9264,N_9109,N_9162);
and U9265 (N_9265,N_9145,N_9170);
and U9266 (N_9266,N_9179,N_9140);
and U9267 (N_9267,N_9117,N_9142);
nand U9268 (N_9268,N_9108,N_9110);
nor U9269 (N_9269,N_9109,N_9193);
and U9270 (N_9270,N_9197,N_9141);
and U9271 (N_9271,N_9186,N_9132);
or U9272 (N_9272,N_9101,N_9136);
or U9273 (N_9273,N_9164,N_9150);
or U9274 (N_9274,N_9170,N_9119);
nor U9275 (N_9275,N_9132,N_9197);
and U9276 (N_9276,N_9119,N_9165);
nand U9277 (N_9277,N_9158,N_9163);
and U9278 (N_9278,N_9197,N_9142);
or U9279 (N_9279,N_9188,N_9195);
or U9280 (N_9280,N_9164,N_9165);
or U9281 (N_9281,N_9167,N_9182);
nor U9282 (N_9282,N_9119,N_9193);
or U9283 (N_9283,N_9190,N_9131);
nand U9284 (N_9284,N_9134,N_9146);
nand U9285 (N_9285,N_9174,N_9179);
nand U9286 (N_9286,N_9132,N_9133);
or U9287 (N_9287,N_9156,N_9137);
nand U9288 (N_9288,N_9118,N_9161);
nor U9289 (N_9289,N_9129,N_9130);
and U9290 (N_9290,N_9120,N_9173);
and U9291 (N_9291,N_9172,N_9166);
nor U9292 (N_9292,N_9187,N_9152);
and U9293 (N_9293,N_9199,N_9138);
or U9294 (N_9294,N_9107,N_9152);
and U9295 (N_9295,N_9108,N_9132);
nor U9296 (N_9296,N_9195,N_9186);
nor U9297 (N_9297,N_9158,N_9168);
and U9298 (N_9298,N_9152,N_9179);
nand U9299 (N_9299,N_9140,N_9164);
and U9300 (N_9300,N_9234,N_9288);
or U9301 (N_9301,N_9206,N_9233);
and U9302 (N_9302,N_9245,N_9203);
nand U9303 (N_9303,N_9262,N_9296);
or U9304 (N_9304,N_9240,N_9290);
nor U9305 (N_9305,N_9250,N_9269);
nand U9306 (N_9306,N_9292,N_9213);
nor U9307 (N_9307,N_9253,N_9249);
and U9308 (N_9308,N_9252,N_9204);
and U9309 (N_9309,N_9226,N_9216);
and U9310 (N_9310,N_9229,N_9277);
nor U9311 (N_9311,N_9241,N_9220);
or U9312 (N_9312,N_9211,N_9212);
and U9313 (N_9313,N_9210,N_9284);
nor U9314 (N_9314,N_9215,N_9218);
nor U9315 (N_9315,N_9254,N_9223);
nand U9316 (N_9316,N_9294,N_9255);
nor U9317 (N_9317,N_9278,N_9266);
and U9318 (N_9318,N_9231,N_9271);
nand U9319 (N_9319,N_9247,N_9267);
or U9320 (N_9320,N_9244,N_9286);
or U9321 (N_9321,N_9268,N_9258);
nand U9322 (N_9322,N_9217,N_9295);
nand U9323 (N_9323,N_9265,N_9209);
nor U9324 (N_9324,N_9219,N_9270);
nor U9325 (N_9325,N_9259,N_9280);
nand U9326 (N_9326,N_9222,N_9298);
or U9327 (N_9327,N_9297,N_9201);
nand U9328 (N_9328,N_9237,N_9289);
nor U9329 (N_9329,N_9273,N_9251);
and U9330 (N_9330,N_9230,N_9260);
or U9331 (N_9331,N_9236,N_9285);
nor U9332 (N_9332,N_9214,N_9239);
nor U9333 (N_9333,N_9275,N_9225);
and U9334 (N_9334,N_9235,N_9282);
nor U9335 (N_9335,N_9291,N_9232);
and U9336 (N_9336,N_9276,N_9248);
nand U9337 (N_9337,N_9257,N_9263);
nor U9338 (N_9338,N_9279,N_9274);
nand U9339 (N_9339,N_9228,N_9287);
nor U9340 (N_9340,N_9200,N_9242);
nor U9341 (N_9341,N_9221,N_9227);
and U9342 (N_9342,N_9205,N_9207);
xnor U9343 (N_9343,N_9261,N_9238);
nand U9344 (N_9344,N_9202,N_9293);
nor U9345 (N_9345,N_9224,N_9272);
nand U9346 (N_9346,N_9243,N_9299);
nand U9347 (N_9347,N_9256,N_9208);
nand U9348 (N_9348,N_9264,N_9281);
nand U9349 (N_9349,N_9283,N_9246);
nor U9350 (N_9350,N_9291,N_9285);
xnor U9351 (N_9351,N_9233,N_9217);
nand U9352 (N_9352,N_9207,N_9262);
and U9353 (N_9353,N_9255,N_9284);
and U9354 (N_9354,N_9252,N_9250);
nand U9355 (N_9355,N_9208,N_9223);
or U9356 (N_9356,N_9228,N_9296);
or U9357 (N_9357,N_9243,N_9241);
nand U9358 (N_9358,N_9271,N_9232);
nand U9359 (N_9359,N_9203,N_9299);
nand U9360 (N_9360,N_9259,N_9248);
nor U9361 (N_9361,N_9207,N_9200);
nand U9362 (N_9362,N_9258,N_9288);
or U9363 (N_9363,N_9294,N_9202);
nor U9364 (N_9364,N_9260,N_9220);
nand U9365 (N_9365,N_9208,N_9257);
nor U9366 (N_9366,N_9292,N_9291);
and U9367 (N_9367,N_9246,N_9294);
nor U9368 (N_9368,N_9255,N_9240);
nand U9369 (N_9369,N_9292,N_9254);
and U9370 (N_9370,N_9211,N_9263);
nand U9371 (N_9371,N_9291,N_9235);
and U9372 (N_9372,N_9296,N_9209);
nand U9373 (N_9373,N_9274,N_9209);
or U9374 (N_9374,N_9255,N_9257);
or U9375 (N_9375,N_9233,N_9268);
or U9376 (N_9376,N_9269,N_9200);
nor U9377 (N_9377,N_9202,N_9247);
nand U9378 (N_9378,N_9213,N_9294);
nand U9379 (N_9379,N_9275,N_9264);
and U9380 (N_9380,N_9206,N_9288);
nor U9381 (N_9381,N_9294,N_9210);
or U9382 (N_9382,N_9295,N_9216);
nand U9383 (N_9383,N_9215,N_9212);
nand U9384 (N_9384,N_9219,N_9228);
nand U9385 (N_9385,N_9228,N_9275);
nand U9386 (N_9386,N_9216,N_9222);
nand U9387 (N_9387,N_9284,N_9244);
nand U9388 (N_9388,N_9280,N_9292);
or U9389 (N_9389,N_9219,N_9227);
nor U9390 (N_9390,N_9259,N_9296);
or U9391 (N_9391,N_9231,N_9213);
or U9392 (N_9392,N_9275,N_9210);
nor U9393 (N_9393,N_9269,N_9277);
nor U9394 (N_9394,N_9220,N_9234);
nand U9395 (N_9395,N_9229,N_9250);
nand U9396 (N_9396,N_9270,N_9211);
nor U9397 (N_9397,N_9222,N_9254);
nand U9398 (N_9398,N_9278,N_9251);
nand U9399 (N_9399,N_9224,N_9237);
and U9400 (N_9400,N_9367,N_9357);
nand U9401 (N_9401,N_9350,N_9399);
nor U9402 (N_9402,N_9351,N_9312);
nand U9403 (N_9403,N_9331,N_9335);
and U9404 (N_9404,N_9300,N_9328);
nand U9405 (N_9405,N_9398,N_9348);
and U9406 (N_9406,N_9342,N_9333);
or U9407 (N_9407,N_9379,N_9303);
or U9408 (N_9408,N_9356,N_9387);
or U9409 (N_9409,N_9364,N_9346);
nand U9410 (N_9410,N_9395,N_9372);
or U9411 (N_9411,N_9306,N_9338);
nor U9412 (N_9412,N_9377,N_9371);
and U9413 (N_9413,N_9339,N_9370);
or U9414 (N_9414,N_9309,N_9340);
or U9415 (N_9415,N_9362,N_9365);
nor U9416 (N_9416,N_9307,N_9305);
nand U9417 (N_9417,N_9374,N_9323);
or U9418 (N_9418,N_9327,N_9314);
nor U9419 (N_9419,N_9354,N_9373);
nand U9420 (N_9420,N_9366,N_9324);
nand U9421 (N_9421,N_9316,N_9343);
and U9422 (N_9422,N_9326,N_9344);
and U9423 (N_9423,N_9349,N_9353);
xor U9424 (N_9424,N_9341,N_9391);
nor U9425 (N_9425,N_9384,N_9361);
nor U9426 (N_9426,N_9358,N_9393);
nand U9427 (N_9427,N_9359,N_9345);
or U9428 (N_9428,N_9385,N_9388);
nand U9429 (N_9429,N_9389,N_9382);
nand U9430 (N_9430,N_9322,N_9368);
nor U9431 (N_9431,N_9313,N_9317);
and U9432 (N_9432,N_9369,N_9392);
and U9433 (N_9433,N_9383,N_9318);
nor U9434 (N_9434,N_9315,N_9332);
nand U9435 (N_9435,N_9378,N_9360);
nand U9436 (N_9436,N_9397,N_9319);
and U9437 (N_9437,N_9320,N_9330);
and U9438 (N_9438,N_9325,N_9311);
nor U9439 (N_9439,N_9329,N_9380);
nand U9440 (N_9440,N_9394,N_9386);
or U9441 (N_9441,N_9355,N_9302);
nor U9442 (N_9442,N_9334,N_9308);
nand U9443 (N_9443,N_9336,N_9321);
and U9444 (N_9444,N_9310,N_9352);
nor U9445 (N_9445,N_9304,N_9396);
nor U9446 (N_9446,N_9337,N_9376);
nand U9447 (N_9447,N_9301,N_9390);
or U9448 (N_9448,N_9347,N_9363);
or U9449 (N_9449,N_9375,N_9381);
and U9450 (N_9450,N_9339,N_9318);
nor U9451 (N_9451,N_9346,N_9311);
or U9452 (N_9452,N_9385,N_9322);
nor U9453 (N_9453,N_9395,N_9364);
and U9454 (N_9454,N_9321,N_9347);
nand U9455 (N_9455,N_9358,N_9302);
and U9456 (N_9456,N_9349,N_9389);
or U9457 (N_9457,N_9335,N_9355);
nor U9458 (N_9458,N_9368,N_9317);
and U9459 (N_9459,N_9309,N_9354);
nor U9460 (N_9460,N_9382,N_9335);
nor U9461 (N_9461,N_9372,N_9385);
or U9462 (N_9462,N_9341,N_9351);
or U9463 (N_9463,N_9311,N_9371);
and U9464 (N_9464,N_9375,N_9318);
and U9465 (N_9465,N_9331,N_9317);
and U9466 (N_9466,N_9398,N_9358);
or U9467 (N_9467,N_9358,N_9363);
nand U9468 (N_9468,N_9343,N_9309);
nor U9469 (N_9469,N_9368,N_9399);
nand U9470 (N_9470,N_9312,N_9386);
xor U9471 (N_9471,N_9371,N_9387);
nor U9472 (N_9472,N_9396,N_9334);
and U9473 (N_9473,N_9308,N_9385);
xnor U9474 (N_9474,N_9353,N_9391);
nand U9475 (N_9475,N_9337,N_9361);
nand U9476 (N_9476,N_9319,N_9336);
and U9477 (N_9477,N_9378,N_9397);
nor U9478 (N_9478,N_9327,N_9355);
nand U9479 (N_9479,N_9306,N_9347);
nand U9480 (N_9480,N_9333,N_9358);
nand U9481 (N_9481,N_9321,N_9398);
nor U9482 (N_9482,N_9377,N_9392);
nand U9483 (N_9483,N_9369,N_9320);
and U9484 (N_9484,N_9332,N_9375);
and U9485 (N_9485,N_9384,N_9382);
and U9486 (N_9486,N_9349,N_9318);
nand U9487 (N_9487,N_9346,N_9304);
nor U9488 (N_9488,N_9334,N_9343);
xnor U9489 (N_9489,N_9326,N_9331);
and U9490 (N_9490,N_9324,N_9341);
nand U9491 (N_9491,N_9328,N_9374);
nor U9492 (N_9492,N_9347,N_9390);
and U9493 (N_9493,N_9350,N_9389);
nand U9494 (N_9494,N_9324,N_9380);
xor U9495 (N_9495,N_9382,N_9396);
nand U9496 (N_9496,N_9315,N_9310);
and U9497 (N_9497,N_9384,N_9360);
and U9498 (N_9498,N_9348,N_9378);
or U9499 (N_9499,N_9373,N_9343);
or U9500 (N_9500,N_9414,N_9478);
nor U9501 (N_9501,N_9419,N_9484);
and U9502 (N_9502,N_9436,N_9480);
nor U9503 (N_9503,N_9434,N_9468);
nand U9504 (N_9504,N_9499,N_9403);
nand U9505 (N_9505,N_9445,N_9423);
or U9506 (N_9506,N_9416,N_9450);
or U9507 (N_9507,N_9472,N_9459);
nor U9508 (N_9508,N_9481,N_9444);
nand U9509 (N_9509,N_9447,N_9424);
or U9510 (N_9510,N_9498,N_9476);
nand U9511 (N_9511,N_9421,N_9432);
nand U9512 (N_9512,N_9452,N_9428);
xor U9513 (N_9513,N_9443,N_9464);
and U9514 (N_9514,N_9490,N_9494);
and U9515 (N_9515,N_9491,N_9497);
nor U9516 (N_9516,N_9460,N_9470);
nor U9517 (N_9517,N_9448,N_9426);
nor U9518 (N_9518,N_9400,N_9463);
nand U9519 (N_9519,N_9405,N_9429);
and U9520 (N_9520,N_9487,N_9457);
nor U9521 (N_9521,N_9420,N_9454);
nor U9522 (N_9522,N_9465,N_9466);
nor U9523 (N_9523,N_9467,N_9427);
nand U9524 (N_9524,N_9462,N_9458);
and U9525 (N_9525,N_9437,N_9455);
nand U9526 (N_9526,N_9409,N_9412);
or U9527 (N_9527,N_9456,N_9417);
nor U9528 (N_9528,N_9479,N_9492);
and U9529 (N_9529,N_9477,N_9488);
or U9530 (N_9530,N_9408,N_9439);
nor U9531 (N_9531,N_9449,N_9495);
nand U9532 (N_9532,N_9469,N_9413);
nor U9533 (N_9533,N_9410,N_9486);
and U9534 (N_9534,N_9440,N_9402);
nor U9535 (N_9535,N_9415,N_9431);
nand U9536 (N_9536,N_9475,N_9442);
and U9537 (N_9537,N_9438,N_9473);
and U9538 (N_9538,N_9496,N_9474);
and U9539 (N_9539,N_9435,N_9493);
or U9540 (N_9540,N_9433,N_9453);
or U9541 (N_9541,N_9406,N_9483);
nor U9542 (N_9542,N_9407,N_9422);
or U9543 (N_9543,N_9411,N_9485);
nor U9544 (N_9544,N_9430,N_9401);
nor U9545 (N_9545,N_9418,N_9482);
nor U9546 (N_9546,N_9451,N_9446);
and U9547 (N_9547,N_9461,N_9441);
and U9548 (N_9548,N_9489,N_9471);
nand U9549 (N_9549,N_9404,N_9425);
and U9550 (N_9550,N_9463,N_9405);
and U9551 (N_9551,N_9418,N_9413);
nand U9552 (N_9552,N_9470,N_9455);
nor U9553 (N_9553,N_9436,N_9414);
or U9554 (N_9554,N_9427,N_9409);
nand U9555 (N_9555,N_9441,N_9439);
and U9556 (N_9556,N_9403,N_9418);
or U9557 (N_9557,N_9491,N_9448);
nor U9558 (N_9558,N_9415,N_9450);
xor U9559 (N_9559,N_9466,N_9451);
nand U9560 (N_9560,N_9406,N_9481);
nand U9561 (N_9561,N_9468,N_9417);
nor U9562 (N_9562,N_9451,N_9487);
and U9563 (N_9563,N_9431,N_9461);
nand U9564 (N_9564,N_9482,N_9428);
nor U9565 (N_9565,N_9432,N_9428);
nor U9566 (N_9566,N_9418,N_9496);
nor U9567 (N_9567,N_9471,N_9493);
nand U9568 (N_9568,N_9428,N_9480);
nor U9569 (N_9569,N_9436,N_9442);
xnor U9570 (N_9570,N_9446,N_9423);
nor U9571 (N_9571,N_9494,N_9456);
and U9572 (N_9572,N_9401,N_9461);
or U9573 (N_9573,N_9452,N_9420);
and U9574 (N_9574,N_9428,N_9441);
nand U9575 (N_9575,N_9481,N_9401);
nand U9576 (N_9576,N_9484,N_9478);
or U9577 (N_9577,N_9460,N_9456);
or U9578 (N_9578,N_9448,N_9498);
and U9579 (N_9579,N_9406,N_9497);
xnor U9580 (N_9580,N_9455,N_9498);
or U9581 (N_9581,N_9450,N_9456);
or U9582 (N_9582,N_9445,N_9434);
nand U9583 (N_9583,N_9437,N_9416);
nand U9584 (N_9584,N_9435,N_9405);
nand U9585 (N_9585,N_9442,N_9433);
or U9586 (N_9586,N_9405,N_9478);
nor U9587 (N_9587,N_9450,N_9487);
nor U9588 (N_9588,N_9497,N_9405);
and U9589 (N_9589,N_9487,N_9461);
or U9590 (N_9590,N_9455,N_9451);
or U9591 (N_9591,N_9440,N_9400);
nor U9592 (N_9592,N_9477,N_9425);
and U9593 (N_9593,N_9422,N_9493);
nor U9594 (N_9594,N_9416,N_9423);
or U9595 (N_9595,N_9467,N_9473);
or U9596 (N_9596,N_9420,N_9432);
nand U9597 (N_9597,N_9404,N_9417);
and U9598 (N_9598,N_9493,N_9496);
or U9599 (N_9599,N_9461,N_9412);
or U9600 (N_9600,N_9591,N_9515);
and U9601 (N_9601,N_9528,N_9579);
nand U9602 (N_9602,N_9553,N_9534);
nand U9603 (N_9603,N_9551,N_9502);
nor U9604 (N_9604,N_9540,N_9524);
and U9605 (N_9605,N_9529,N_9584);
nand U9606 (N_9606,N_9568,N_9522);
and U9607 (N_9607,N_9550,N_9516);
nor U9608 (N_9608,N_9546,N_9530);
nor U9609 (N_9609,N_9572,N_9535);
nand U9610 (N_9610,N_9590,N_9504);
or U9611 (N_9611,N_9554,N_9526);
and U9612 (N_9612,N_9532,N_9588);
nand U9613 (N_9613,N_9576,N_9506);
nor U9614 (N_9614,N_9527,N_9587);
nand U9615 (N_9615,N_9558,N_9565);
or U9616 (N_9616,N_9557,N_9517);
and U9617 (N_9617,N_9573,N_9585);
nor U9618 (N_9618,N_9536,N_9592);
or U9619 (N_9619,N_9594,N_9549);
nand U9620 (N_9620,N_9544,N_9542);
or U9621 (N_9621,N_9523,N_9577);
and U9622 (N_9622,N_9547,N_9598);
nor U9623 (N_9623,N_9574,N_9580);
xnor U9624 (N_9624,N_9569,N_9548);
nor U9625 (N_9625,N_9539,N_9582);
and U9626 (N_9626,N_9501,N_9509);
nor U9627 (N_9627,N_9567,N_9500);
and U9628 (N_9628,N_9563,N_9520);
or U9629 (N_9629,N_9555,N_9541);
or U9630 (N_9630,N_9533,N_9525);
nand U9631 (N_9631,N_9537,N_9564);
nor U9632 (N_9632,N_9578,N_9519);
nor U9633 (N_9633,N_9559,N_9552);
and U9634 (N_9634,N_9560,N_9562);
nand U9635 (N_9635,N_9586,N_9571);
nor U9636 (N_9636,N_9570,N_9521);
nor U9637 (N_9637,N_9513,N_9543);
nand U9638 (N_9638,N_9583,N_9595);
and U9639 (N_9639,N_9508,N_9545);
or U9640 (N_9640,N_9512,N_9566);
nand U9641 (N_9641,N_9511,N_9597);
and U9642 (N_9642,N_9518,N_9510);
or U9643 (N_9643,N_9531,N_9561);
or U9644 (N_9644,N_9575,N_9599);
or U9645 (N_9645,N_9514,N_9556);
or U9646 (N_9646,N_9503,N_9589);
nand U9647 (N_9647,N_9593,N_9596);
xor U9648 (N_9648,N_9507,N_9581);
nand U9649 (N_9649,N_9505,N_9538);
nor U9650 (N_9650,N_9589,N_9565);
nand U9651 (N_9651,N_9563,N_9559);
or U9652 (N_9652,N_9544,N_9558);
or U9653 (N_9653,N_9570,N_9519);
nor U9654 (N_9654,N_9584,N_9508);
xor U9655 (N_9655,N_9535,N_9505);
or U9656 (N_9656,N_9521,N_9510);
nor U9657 (N_9657,N_9596,N_9530);
nand U9658 (N_9658,N_9528,N_9507);
nand U9659 (N_9659,N_9594,N_9563);
nand U9660 (N_9660,N_9592,N_9594);
nand U9661 (N_9661,N_9550,N_9518);
and U9662 (N_9662,N_9599,N_9573);
nor U9663 (N_9663,N_9528,N_9588);
nand U9664 (N_9664,N_9541,N_9577);
or U9665 (N_9665,N_9557,N_9512);
nor U9666 (N_9666,N_9528,N_9524);
nor U9667 (N_9667,N_9520,N_9544);
nor U9668 (N_9668,N_9564,N_9590);
or U9669 (N_9669,N_9589,N_9511);
nand U9670 (N_9670,N_9542,N_9588);
or U9671 (N_9671,N_9532,N_9557);
nand U9672 (N_9672,N_9565,N_9559);
and U9673 (N_9673,N_9574,N_9565);
nor U9674 (N_9674,N_9584,N_9564);
or U9675 (N_9675,N_9595,N_9505);
or U9676 (N_9676,N_9587,N_9578);
and U9677 (N_9677,N_9506,N_9587);
or U9678 (N_9678,N_9554,N_9595);
and U9679 (N_9679,N_9554,N_9590);
or U9680 (N_9680,N_9515,N_9502);
and U9681 (N_9681,N_9550,N_9513);
and U9682 (N_9682,N_9553,N_9595);
nor U9683 (N_9683,N_9562,N_9579);
or U9684 (N_9684,N_9559,N_9502);
nor U9685 (N_9685,N_9561,N_9552);
nor U9686 (N_9686,N_9520,N_9560);
and U9687 (N_9687,N_9589,N_9533);
or U9688 (N_9688,N_9536,N_9597);
nand U9689 (N_9689,N_9580,N_9578);
nand U9690 (N_9690,N_9524,N_9512);
or U9691 (N_9691,N_9597,N_9539);
nor U9692 (N_9692,N_9554,N_9549);
and U9693 (N_9693,N_9517,N_9567);
nand U9694 (N_9694,N_9595,N_9552);
nor U9695 (N_9695,N_9522,N_9534);
nor U9696 (N_9696,N_9502,N_9521);
and U9697 (N_9697,N_9570,N_9596);
and U9698 (N_9698,N_9569,N_9532);
nor U9699 (N_9699,N_9555,N_9525);
nand U9700 (N_9700,N_9641,N_9612);
and U9701 (N_9701,N_9602,N_9614);
nand U9702 (N_9702,N_9633,N_9675);
or U9703 (N_9703,N_9615,N_9666);
nor U9704 (N_9704,N_9683,N_9684);
nand U9705 (N_9705,N_9674,N_9616);
and U9706 (N_9706,N_9672,N_9622);
or U9707 (N_9707,N_9604,N_9655);
nor U9708 (N_9708,N_9607,N_9664);
or U9709 (N_9709,N_9651,N_9687);
nor U9710 (N_9710,N_9649,N_9673);
or U9711 (N_9711,N_9669,N_9645);
nand U9712 (N_9712,N_9629,N_9685);
or U9713 (N_9713,N_9689,N_9619);
nand U9714 (N_9714,N_9652,N_9606);
nor U9715 (N_9715,N_9671,N_9611);
or U9716 (N_9716,N_9693,N_9659);
nor U9717 (N_9717,N_9625,N_9682);
or U9718 (N_9718,N_9621,N_9624);
nor U9719 (N_9719,N_9608,N_9699);
and U9720 (N_9720,N_9638,N_9697);
nand U9721 (N_9721,N_9617,N_9628);
nand U9722 (N_9722,N_9660,N_9650);
nor U9723 (N_9723,N_9605,N_9636);
and U9724 (N_9724,N_9609,N_9676);
nand U9725 (N_9725,N_9670,N_9620);
and U9726 (N_9726,N_9618,N_9635);
nand U9727 (N_9727,N_9600,N_9698);
nand U9728 (N_9728,N_9632,N_9634);
nor U9729 (N_9729,N_9653,N_9696);
nor U9730 (N_9730,N_9630,N_9623);
nand U9731 (N_9731,N_9679,N_9661);
nand U9732 (N_9732,N_9640,N_9657);
or U9733 (N_9733,N_9613,N_9648);
nor U9734 (N_9734,N_9663,N_9654);
and U9735 (N_9735,N_9610,N_9688);
and U9736 (N_9736,N_9643,N_9692);
nor U9737 (N_9737,N_9695,N_9678);
and U9738 (N_9738,N_9681,N_9656);
and U9739 (N_9739,N_9601,N_9690);
nor U9740 (N_9740,N_9662,N_9647);
or U9741 (N_9741,N_9631,N_9691);
and U9742 (N_9742,N_9627,N_9694);
or U9743 (N_9743,N_9639,N_9603);
nor U9744 (N_9744,N_9642,N_9668);
and U9745 (N_9745,N_9646,N_9626);
or U9746 (N_9746,N_9665,N_9658);
and U9747 (N_9747,N_9680,N_9667);
nand U9748 (N_9748,N_9677,N_9637);
nor U9749 (N_9749,N_9644,N_9686);
nand U9750 (N_9750,N_9676,N_9605);
nor U9751 (N_9751,N_9694,N_9668);
nand U9752 (N_9752,N_9628,N_9654);
or U9753 (N_9753,N_9600,N_9660);
or U9754 (N_9754,N_9696,N_9681);
and U9755 (N_9755,N_9623,N_9603);
nand U9756 (N_9756,N_9623,N_9697);
and U9757 (N_9757,N_9670,N_9605);
and U9758 (N_9758,N_9659,N_9651);
xor U9759 (N_9759,N_9647,N_9689);
nor U9760 (N_9760,N_9689,N_9639);
or U9761 (N_9761,N_9604,N_9661);
nand U9762 (N_9762,N_9602,N_9655);
and U9763 (N_9763,N_9695,N_9652);
or U9764 (N_9764,N_9609,N_9610);
nand U9765 (N_9765,N_9629,N_9690);
nand U9766 (N_9766,N_9627,N_9686);
or U9767 (N_9767,N_9672,N_9682);
or U9768 (N_9768,N_9652,N_9642);
nor U9769 (N_9769,N_9601,N_9657);
nor U9770 (N_9770,N_9645,N_9682);
and U9771 (N_9771,N_9619,N_9670);
and U9772 (N_9772,N_9688,N_9674);
xnor U9773 (N_9773,N_9692,N_9695);
or U9774 (N_9774,N_9658,N_9605);
and U9775 (N_9775,N_9681,N_9674);
nand U9776 (N_9776,N_9617,N_9640);
and U9777 (N_9777,N_9624,N_9644);
nor U9778 (N_9778,N_9603,N_9691);
nor U9779 (N_9779,N_9656,N_9615);
or U9780 (N_9780,N_9699,N_9694);
nand U9781 (N_9781,N_9619,N_9622);
or U9782 (N_9782,N_9657,N_9650);
or U9783 (N_9783,N_9650,N_9663);
and U9784 (N_9784,N_9679,N_9653);
or U9785 (N_9785,N_9675,N_9690);
nand U9786 (N_9786,N_9667,N_9662);
nor U9787 (N_9787,N_9603,N_9618);
and U9788 (N_9788,N_9619,N_9667);
nor U9789 (N_9789,N_9629,N_9696);
xnor U9790 (N_9790,N_9679,N_9621);
nand U9791 (N_9791,N_9606,N_9644);
or U9792 (N_9792,N_9662,N_9675);
nand U9793 (N_9793,N_9690,N_9651);
nor U9794 (N_9794,N_9664,N_9654);
and U9795 (N_9795,N_9635,N_9695);
nor U9796 (N_9796,N_9668,N_9685);
or U9797 (N_9797,N_9646,N_9699);
and U9798 (N_9798,N_9662,N_9615);
and U9799 (N_9799,N_9626,N_9651);
nand U9800 (N_9800,N_9749,N_9721);
nor U9801 (N_9801,N_9733,N_9777);
nor U9802 (N_9802,N_9726,N_9714);
or U9803 (N_9803,N_9720,N_9738);
nand U9804 (N_9804,N_9768,N_9718);
nor U9805 (N_9805,N_9702,N_9745);
or U9806 (N_9806,N_9705,N_9731);
and U9807 (N_9807,N_9753,N_9780);
and U9808 (N_9808,N_9742,N_9703);
xor U9809 (N_9809,N_9744,N_9774);
nand U9810 (N_9810,N_9751,N_9734);
and U9811 (N_9811,N_9760,N_9752);
or U9812 (N_9812,N_9730,N_9724);
or U9813 (N_9813,N_9779,N_9791);
nor U9814 (N_9814,N_9706,N_9773);
nor U9815 (N_9815,N_9769,N_9756);
or U9816 (N_9816,N_9766,N_9750);
nor U9817 (N_9817,N_9743,N_9712);
nor U9818 (N_9818,N_9741,N_9783);
nor U9819 (N_9819,N_9796,N_9717);
or U9820 (N_9820,N_9784,N_9782);
nor U9821 (N_9821,N_9790,N_9740);
or U9822 (N_9822,N_9748,N_9739);
nor U9823 (N_9823,N_9792,N_9785);
or U9824 (N_9824,N_9765,N_9793);
nor U9825 (N_9825,N_9798,N_9797);
or U9826 (N_9826,N_9776,N_9727);
nand U9827 (N_9827,N_9772,N_9719);
nor U9828 (N_9828,N_9755,N_9757);
nor U9829 (N_9829,N_9778,N_9761);
and U9830 (N_9830,N_9775,N_9786);
or U9831 (N_9831,N_9701,N_9716);
nor U9832 (N_9832,N_9747,N_9707);
nand U9833 (N_9833,N_9770,N_9758);
or U9834 (N_9834,N_9735,N_9700);
and U9835 (N_9835,N_9711,N_9736);
and U9836 (N_9836,N_9771,N_9746);
nor U9837 (N_9837,N_9729,N_9764);
or U9838 (N_9838,N_9713,N_9710);
and U9839 (N_9839,N_9762,N_9763);
or U9840 (N_9840,N_9725,N_9767);
or U9841 (N_9841,N_9732,N_9787);
nor U9842 (N_9842,N_9737,N_9723);
nand U9843 (N_9843,N_9759,N_9799);
nor U9844 (N_9844,N_9722,N_9781);
and U9845 (N_9845,N_9754,N_9789);
nand U9846 (N_9846,N_9795,N_9708);
or U9847 (N_9847,N_9728,N_9715);
nor U9848 (N_9848,N_9704,N_9709);
nand U9849 (N_9849,N_9788,N_9794);
nor U9850 (N_9850,N_9752,N_9732);
or U9851 (N_9851,N_9770,N_9775);
and U9852 (N_9852,N_9719,N_9736);
nand U9853 (N_9853,N_9742,N_9708);
nor U9854 (N_9854,N_9760,N_9780);
nand U9855 (N_9855,N_9715,N_9753);
nor U9856 (N_9856,N_9712,N_9753);
and U9857 (N_9857,N_9758,N_9784);
nor U9858 (N_9858,N_9770,N_9784);
nor U9859 (N_9859,N_9737,N_9739);
or U9860 (N_9860,N_9708,N_9719);
nand U9861 (N_9861,N_9734,N_9744);
xnor U9862 (N_9862,N_9764,N_9750);
nand U9863 (N_9863,N_9724,N_9788);
or U9864 (N_9864,N_9785,N_9772);
nand U9865 (N_9865,N_9779,N_9711);
nand U9866 (N_9866,N_9778,N_9747);
and U9867 (N_9867,N_9787,N_9717);
nand U9868 (N_9868,N_9723,N_9751);
nand U9869 (N_9869,N_9793,N_9791);
nand U9870 (N_9870,N_9772,N_9733);
and U9871 (N_9871,N_9796,N_9759);
or U9872 (N_9872,N_9769,N_9764);
and U9873 (N_9873,N_9702,N_9794);
or U9874 (N_9874,N_9744,N_9737);
nand U9875 (N_9875,N_9779,N_9703);
and U9876 (N_9876,N_9793,N_9747);
nand U9877 (N_9877,N_9717,N_9713);
nor U9878 (N_9878,N_9718,N_9783);
nor U9879 (N_9879,N_9745,N_9722);
and U9880 (N_9880,N_9741,N_9702);
and U9881 (N_9881,N_9799,N_9749);
nor U9882 (N_9882,N_9769,N_9762);
and U9883 (N_9883,N_9709,N_9707);
nor U9884 (N_9884,N_9798,N_9788);
and U9885 (N_9885,N_9764,N_9719);
nor U9886 (N_9886,N_9709,N_9711);
and U9887 (N_9887,N_9776,N_9739);
nor U9888 (N_9888,N_9780,N_9793);
or U9889 (N_9889,N_9724,N_9770);
and U9890 (N_9890,N_9768,N_9733);
and U9891 (N_9891,N_9761,N_9748);
nor U9892 (N_9892,N_9786,N_9714);
or U9893 (N_9893,N_9709,N_9791);
or U9894 (N_9894,N_9773,N_9785);
or U9895 (N_9895,N_9703,N_9741);
nand U9896 (N_9896,N_9789,N_9783);
nor U9897 (N_9897,N_9770,N_9705);
or U9898 (N_9898,N_9710,N_9723);
nand U9899 (N_9899,N_9706,N_9759);
and U9900 (N_9900,N_9816,N_9877);
and U9901 (N_9901,N_9819,N_9807);
nand U9902 (N_9902,N_9860,N_9833);
nand U9903 (N_9903,N_9897,N_9804);
nand U9904 (N_9904,N_9891,N_9809);
nand U9905 (N_9905,N_9868,N_9810);
or U9906 (N_9906,N_9822,N_9886);
and U9907 (N_9907,N_9844,N_9888);
or U9908 (N_9908,N_9864,N_9847);
and U9909 (N_9909,N_9838,N_9830);
nor U9910 (N_9910,N_9800,N_9825);
or U9911 (N_9911,N_9852,N_9840);
or U9912 (N_9912,N_9849,N_9873);
or U9913 (N_9913,N_9898,N_9894);
nand U9914 (N_9914,N_9846,N_9889);
nor U9915 (N_9915,N_9890,N_9826);
or U9916 (N_9916,N_9801,N_9812);
nand U9917 (N_9917,N_9892,N_9885);
nor U9918 (N_9918,N_9837,N_9820);
and U9919 (N_9919,N_9842,N_9882);
and U9920 (N_9920,N_9818,N_9845);
and U9921 (N_9921,N_9854,N_9823);
and U9922 (N_9922,N_9874,N_9893);
xnor U9923 (N_9923,N_9853,N_9863);
and U9924 (N_9924,N_9834,N_9858);
nand U9925 (N_9925,N_9857,N_9850);
nand U9926 (N_9926,N_9829,N_9802);
or U9927 (N_9927,N_9875,N_9813);
or U9928 (N_9928,N_9831,N_9867);
nand U9929 (N_9929,N_9871,N_9836);
or U9930 (N_9930,N_9856,N_9815);
nor U9931 (N_9931,N_9861,N_9808);
nand U9932 (N_9932,N_9843,N_9848);
and U9933 (N_9933,N_9835,N_9862);
nor U9934 (N_9934,N_9805,N_9876);
xor U9935 (N_9935,N_9899,N_9806);
xnor U9936 (N_9936,N_9803,N_9865);
and U9937 (N_9937,N_9855,N_9880);
nand U9938 (N_9938,N_9817,N_9866);
nor U9939 (N_9939,N_9881,N_9896);
or U9940 (N_9940,N_9859,N_9895);
nor U9941 (N_9941,N_9878,N_9870);
or U9942 (N_9942,N_9879,N_9814);
nor U9943 (N_9943,N_9883,N_9821);
or U9944 (N_9944,N_9887,N_9824);
nand U9945 (N_9945,N_9841,N_9851);
nand U9946 (N_9946,N_9811,N_9828);
and U9947 (N_9947,N_9869,N_9872);
xnor U9948 (N_9948,N_9832,N_9827);
nor U9949 (N_9949,N_9839,N_9884);
nor U9950 (N_9950,N_9825,N_9887);
nor U9951 (N_9951,N_9806,N_9823);
xor U9952 (N_9952,N_9896,N_9880);
or U9953 (N_9953,N_9877,N_9837);
nor U9954 (N_9954,N_9874,N_9859);
nand U9955 (N_9955,N_9879,N_9809);
and U9956 (N_9956,N_9806,N_9821);
and U9957 (N_9957,N_9821,N_9807);
and U9958 (N_9958,N_9821,N_9805);
nand U9959 (N_9959,N_9810,N_9803);
nand U9960 (N_9960,N_9849,N_9880);
and U9961 (N_9961,N_9866,N_9837);
and U9962 (N_9962,N_9898,N_9849);
nor U9963 (N_9963,N_9834,N_9821);
and U9964 (N_9964,N_9875,N_9856);
nand U9965 (N_9965,N_9817,N_9871);
nor U9966 (N_9966,N_9810,N_9812);
or U9967 (N_9967,N_9842,N_9876);
nand U9968 (N_9968,N_9811,N_9864);
or U9969 (N_9969,N_9803,N_9866);
nor U9970 (N_9970,N_9821,N_9822);
and U9971 (N_9971,N_9825,N_9852);
or U9972 (N_9972,N_9898,N_9806);
and U9973 (N_9973,N_9814,N_9858);
or U9974 (N_9974,N_9884,N_9800);
nor U9975 (N_9975,N_9899,N_9851);
and U9976 (N_9976,N_9847,N_9832);
nand U9977 (N_9977,N_9812,N_9886);
or U9978 (N_9978,N_9875,N_9871);
nor U9979 (N_9979,N_9885,N_9886);
and U9980 (N_9980,N_9814,N_9862);
nor U9981 (N_9981,N_9854,N_9884);
or U9982 (N_9982,N_9823,N_9817);
and U9983 (N_9983,N_9838,N_9833);
xnor U9984 (N_9984,N_9821,N_9830);
and U9985 (N_9985,N_9818,N_9824);
nor U9986 (N_9986,N_9842,N_9854);
and U9987 (N_9987,N_9849,N_9827);
nor U9988 (N_9988,N_9816,N_9823);
nor U9989 (N_9989,N_9849,N_9896);
nand U9990 (N_9990,N_9812,N_9821);
and U9991 (N_9991,N_9889,N_9810);
or U9992 (N_9992,N_9864,N_9895);
and U9993 (N_9993,N_9865,N_9841);
nand U9994 (N_9994,N_9805,N_9827);
or U9995 (N_9995,N_9851,N_9816);
or U9996 (N_9996,N_9845,N_9850);
nor U9997 (N_9997,N_9840,N_9870);
and U9998 (N_9998,N_9885,N_9821);
nor U9999 (N_9999,N_9814,N_9893);
and UO_0 (O_0,N_9932,N_9977);
nor UO_1 (O_1,N_9973,N_9924);
nand UO_2 (O_2,N_9927,N_9905);
nor UO_3 (O_3,N_9926,N_9909);
nand UO_4 (O_4,N_9970,N_9910);
nor UO_5 (O_5,N_9919,N_9993);
and UO_6 (O_6,N_9988,N_9912);
or UO_7 (O_7,N_9964,N_9961);
xor UO_8 (O_8,N_9950,N_9960);
or UO_9 (O_9,N_9922,N_9911);
nand UO_10 (O_10,N_9972,N_9936);
or UO_11 (O_11,N_9906,N_9946);
nand UO_12 (O_12,N_9952,N_9978);
nor UO_13 (O_13,N_9904,N_9996);
and UO_14 (O_14,N_9974,N_9902);
or UO_15 (O_15,N_9981,N_9957);
and UO_16 (O_16,N_9969,N_9998);
or UO_17 (O_17,N_9955,N_9966);
nand UO_18 (O_18,N_9913,N_9908);
or UO_19 (O_19,N_9928,N_9929);
nor UO_20 (O_20,N_9997,N_9959);
nor UO_21 (O_21,N_9933,N_9989);
or UO_22 (O_22,N_9939,N_9907);
nor UO_23 (O_23,N_9938,N_9979);
and UO_24 (O_24,N_9948,N_9903);
and UO_25 (O_25,N_9976,N_9931);
or UO_26 (O_26,N_9940,N_9953);
and UO_27 (O_27,N_9930,N_9968);
nor UO_28 (O_28,N_9967,N_9920);
and UO_29 (O_29,N_9958,N_9925);
and UO_30 (O_30,N_9944,N_9985);
or UO_31 (O_31,N_9986,N_9982);
nor UO_32 (O_32,N_9991,N_9975);
or UO_33 (O_33,N_9980,N_9994);
nor UO_34 (O_34,N_9999,N_9971);
nor UO_35 (O_35,N_9984,N_9917);
or UO_36 (O_36,N_9954,N_9921);
and UO_37 (O_37,N_9949,N_9992);
or UO_38 (O_38,N_9915,N_9941);
nand UO_39 (O_39,N_9937,N_9914);
nand UO_40 (O_40,N_9983,N_9947);
nand UO_41 (O_41,N_9901,N_9951);
nor UO_42 (O_42,N_9990,N_9935);
nor UO_43 (O_43,N_9916,N_9943);
nand UO_44 (O_44,N_9934,N_9965);
nor UO_45 (O_45,N_9918,N_9900);
nor UO_46 (O_46,N_9956,N_9987);
nand UO_47 (O_47,N_9942,N_9963);
nand UO_48 (O_48,N_9923,N_9995);
or UO_49 (O_49,N_9962,N_9945);
nor UO_50 (O_50,N_9971,N_9911);
and UO_51 (O_51,N_9973,N_9994);
nor UO_52 (O_52,N_9923,N_9996);
and UO_53 (O_53,N_9904,N_9924);
and UO_54 (O_54,N_9931,N_9994);
or UO_55 (O_55,N_9902,N_9981);
and UO_56 (O_56,N_9996,N_9952);
or UO_57 (O_57,N_9933,N_9919);
nand UO_58 (O_58,N_9975,N_9942);
and UO_59 (O_59,N_9981,N_9941);
and UO_60 (O_60,N_9944,N_9971);
or UO_61 (O_61,N_9914,N_9944);
nor UO_62 (O_62,N_9941,N_9994);
nand UO_63 (O_63,N_9910,N_9908);
nor UO_64 (O_64,N_9938,N_9934);
and UO_65 (O_65,N_9913,N_9912);
nand UO_66 (O_66,N_9993,N_9990);
nor UO_67 (O_67,N_9909,N_9915);
and UO_68 (O_68,N_9956,N_9955);
nand UO_69 (O_69,N_9942,N_9931);
and UO_70 (O_70,N_9921,N_9925);
and UO_71 (O_71,N_9951,N_9936);
nor UO_72 (O_72,N_9913,N_9934);
nand UO_73 (O_73,N_9914,N_9982);
and UO_74 (O_74,N_9956,N_9949);
nor UO_75 (O_75,N_9921,N_9962);
xor UO_76 (O_76,N_9991,N_9914);
or UO_77 (O_77,N_9993,N_9992);
and UO_78 (O_78,N_9925,N_9939);
and UO_79 (O_79,N_9960,N_9926);
nand UO_80 (O_80,N_9965,N_9959);
nor UO_81 (O_81,N_9977,N_9971);
or UO_82 (O_82,N_9970,N_9923);
nand UO_83 (O_83,N_9968,N_9916);
and UO_84 (O_84,N_9930,N_9942);
and UO_85 (O_85,N_9981,N_9983);
or UO_86 (O_86,N_9981,N_9995);
xnor UO_87 (O_87,N_9910,N_9915);
nand UO_88 (O_88,N_9903,N_9972);
and UO_89 (O_89,N_9955,N_9921);
nand UO_90 (O_90,N_9906,N_9912);
or UO_91 (O_91,N_9910,N_9921);
and UO_92 (O_92,N_9993,N_9933);
nor UO_93 (O_93,N_9924,N_9949);
nand UO_94 (O_94,N_9973,N_9903);
nor UO_95 (O_95,N_9940,N_9925);
or UO_96 (O_96,N_9938,N_9902);
nor UO_97 (O_97,N_9995,N_9931);
nand UO_98 (O_98,N_9930,N_9917);
or UO_99 (O_99,N_9949,N_9931);
nand UO_100 (O_100,N_9953,N_9922);
nor UO_101 (O_101,N_9924,N_9926);
nor UO_102 (O_102,N_9974,N_9957);
nand UO_103 (O_103,N_9970,N_9917);
nand UO_104 (O_104,N_9996,N_9913);
nand UO_105 (O_105,N_9932,N_9960);
and UO_106 (O_106,N_9913,N_9930);
nand UO_107 (O_107,N_9933,N_9975);
or UO_108 (O_108,N_9956,N_9966);
nor UO_109 (O_109,N_9976,N_9935);
nand UO_110 (O_110,N_9927,N_9994);
nor UO_111 (O_111,N_9916,N_9910);
nor UO_112 (O_112,N_9945,N_9983);
nor UO_113 (O_113,N_9988,N_9923);
nor UO_114 (O_114,N_9909,N_9932);
and UO_115 (O_115,N_9970,N_9949);
nand UO_116 (O_116,N_9935,N_9977);
nor UO_117 (O_117,N_9911,N_9906);
and UO_118 (O_118,N_9959,N_9915);
and UO_119 (O_119,N_9932,N_9931);
and UO_120 (O_120,N_9963,N_9929);
nor UO_121 (O_121,N_9924,N_9905);
or UO_122 (O_122,N_9940,N_9966);
nor UO_123 (O_123,N_9963,N_9994);
nand UO_124 (O_124,N_9973,N_9981);
and UO_125 (O_125,N_9927,N_9965);
nor UO_126 (O_126,N_9993,N_9955);
nand UO_127 (O_127,N_9904,N_9915);
or UO_128 (O_128,N_9991,N_9902);
nor UO_129 (O_129,N_9939,N_9959);
or UO_130 (O_130,N_9998,N_9907);
xnor UO_131 (O_131,N_9938,N_9976);
or UO_132 (O_132,N_9930,N_9964);
and UO_133 (O_133,N_9928,N_9952);
or UO_134 (O_134,N_9928,N_9949);
or UO_135 (O_135,N_9947,N_9928);
nand UO_136 (O_136,N_9943,N_9936);
nor UO_137 (O_137,N_9984,N_9931);
nor UO_138 (O_138,N_9907,N_9908);
or UO_139 (O_139,N_9912,N_9909);
and UO_140 (O_140,N_9933,N_9930);
and UO_141 (O_141,N_9928,N_9995);
nor UO_142 (O_142,N_9987,N_9935);
nand UO_143 (O_143,N_9910,N_9955);
or UO_144 (O_144,N_9951,N_9925);
and UO_145 (O_145,N_9919,N_9973);
nor UO_146 (O_146,N_9932,N_9945);
and UO_147 (O_147,N_9926,N_9961);
xor UO_148 (O_148,N_9990,N_9973);
xor UO_149 (O_149,N_9940,N_9924);
nand UO_150 (O_150,N_9985,N_9997);
nand UO_151 (O_151,N_9946,N_9920);
nand UO_152 (O_152,N_9989,N_9976);
nor UO_153 (O_153,N_9905,N_9977);
nor UO_154 (O_154,N_9912,N_9982);
and UO_155 (O_155,N_9959,N_9951);
and UO_156 (O_156,N_9906,N_9989);
and UO_157 (O_157,N_9996,N_9974);
and UO_158 (O_158,N_9941,N_9968);
nor UO_159 (O_159,N_9976,N_9990);
nand UO_160 (O_160,N_9929,N_9909);
nor UO_161 (O_161,N_9911,N_9935);
nand UO_162 (O_162,N_9920,N_9983);
nor UO_163 (O_163,N_9926,N_9984);
nor UO_164 (O_164,N_9906,N_9914);
nand UO_165 (O_165,N_9963,N_9950);
nor UO_166 (O_166,N_9925,N_9968);
nor UO_167 (O_167,N_9991,N_9903);
or UO_168 (O_168,N_9953,N_9920);
nand UO_169 (O_169,N_9975,N_9932);
and UO_170 (O_170,N_9998,N_9950);
or UO_171 (O_171,N_9948,N_9967);
or UO_172 (O_172,N_9929,N_9923);
or UO_173 (O_173,N_9998,N_9932);
nor UO_174 (O_174,N_9984,N_9973);
and UO_175 (O_175,N_9931,N_9988);
nor UO_176 (O_176,N_9917,N_9987);
nor UO_177 (O_177,N_9951,N_9967);
or UO_178 (O_178,N_9942,N_9933);
and UO_179 (O_179,N_9933,N_9958);
and UO_180 (O_180,N_9927,N_9938);
and UO_181 (O_181,N_9979,N_9978);
nand UO_182 (O_182,N_9900,N_9916);
nor UO_183 (O_183,N_9986,N_9978);
nor UO_184 (O_184,N_9951,N_9945);
nand UO_185 (O_185,N_9986,N_9900);
or UO_186 (O_186,N_9976,N_9910);
nor UO_187 (O_187,N_9973,N_9999);
nand UO_188 (O_188,N_9987,N_9988);
nor UO_189 (O_189,N_9957,N_9975);
or UO_190 (O_190,N_9903,N_9912);
nor UO_191 (O_191,N_9927,N_9940);
nor UO_192 (O_192,N_9971,N_9908);
nor UO_193 (O_193,N_9914,N_9953);
xnor UO_194 (O_194,N_9938,N_9973);
and UO_195 (O_195,N_9907,N_9909);
nor UO_196 (O_196,N_9956,N_9965);
or UO_197 (O_197,N_9955,N_9915);
and UO_198 (O_198,N_9951,N_9923);
or UO_199 (O_199,N_9926,N_9908);
and UO_200 (O_200,N_9974,N_9945);
and UO_201 (O_201,N_9942,N_9922);
nor UO_202 (O_202,N_9984,N_9979);
nor UO_203 (O_203,N_9990,N_9936);
nor UO_204 (O_204,N_9958,N_9906);
nand UO_205 (O_205,N_9977,N_9903);
nand UO_206 (O_206,N_9980,N_9961);
or UO_207 (O_207,N_9912,N_9960);
nor UO_208 (O_208,N_9988,N_9906);
or UO_209 (O_209,N_9956,N_9912);
nand UO_210 (O_210,N_9998,N_9904);
or UO_211 (O_211,N_9904,N_9970);
or UO_212 (O_212,N_9927,N_9995);
nand UO_213 (O_213,N_9906,N_9925);
or UO_214 (O_214,N_9959,N_9905);
nor UO_215 (O_215,N_9984,N_9937);
and UO_216 (O_216,N_9920,N_9965);
and UO_217 (O_217,N_9970,N_9929);
nand UO_218 (O_218,N_9961,N_9986);
and UO_219 (O_219,N_9986,N_9979);
and UO_220 (O_220,N_9951,N_9913);
xor UO_221 (O_221,N_9904,N_9919);
and UO_222 (O_222,N_9941,N_9966);
nor UO_223 (O_223,N_9967,N_9932);
and UO_224 (O_224,N_9963,N_9996);
and UO_225 (O_225,N_9901,N_9944);
or UO_226 (O_226,N_9973,N_9995);
nand UO_227 (O_227,N_9903,N_9944);
and UO_228 (O_228,N_9928,N_9914);
or UO_229 (O_229,N_9925,N_9974);
nand UO_230 (O_230,N_9961,N_9978);
and UO_231 (O_231,N_9900,N_9950);
or UO_232 (O_232,N_9992,N_9915);
nand UO_233 (O_233,N_9917,N_9902);
nor UO_234 (O_234,N_9937,N_9998);
nor UO_235 (O_235,N_9945,N_9940);
nor UO_236 (O_236,N_9926,N_9922);
nor UO_237 (O_237,N_9975,N_9997);
nand UO_238 (O_238,N_9994,N_9944);
and UO_239 (O_239,N_9912,N_9966);
and UO_240 (O_240,N_9976,N_9922);
and UO_241 (O_241,N_9966,N_9968);
or UO_242 (O_242,N_9909,N_9979);
nor UO_243 (O_243,N_9989,N_9965);
nor UO_244 (O_244,N_9945,N_9912);
xor UO_245 (O_245,N_9978,N_9926);
nor UO_246 (O_246,N_9972,N_9950);
and UO_247 (O_247,N_9944,N_9984);
and UO_248 (O_248,N_9966,N_9986);
nand UO_249 (O_249,N_9926,N_9992);
and UO_250 (O_250,N_9921,N_9932);
and UO_251 (O_251,N_9995,N_9976);
or UO_252 (O_252,N_9947,N_9993);
or UO_253 (O_253,N_9988,N_9902);
nor UO_254 (O_254,N_9967,N_9930);
nand UO_255 (O_255,N_9958,N_9949);
nand UO_256 (O_256,N_9990,N_9972);
or UO_257 (O_257,N_9996,N_9965);
nor UO_258 (O_258,N_9965,N_9940);
and UO_259 (O_259,N_9970,N_9901);
or UO_260 (O_260,N_9927,N_9925);
nor UO_261 (O_261,N_9974,N_9909);
or UO_262 (O_262,N_9949,N_9977);
or UO_263 (O_263,N_9986,N_9951);
and UO_264 (O_264,N_9968,N_9948);
nand UO_265 (O_265,N_9929,N_9933);
nand UO_266 (O_266,N_9904,N_9993);
nor UO_267 (O_267,N_9921,N_9938);
and UO_268 (O_268,N_9987,N_9966);
or UO_269 (O_269,N_9934,N_9942);
nand UO_270 (O_270,N_9948,N_9943);
nor UO_271 (O_271,N_9926,N_9933);
and UO_272 (O_272,N_9979,N_9944);
nor UO_273 (O_273,N_9973,N_9952);
or UO_274 (O_274,N_9955,N_9980);
or UO_275 (O_275,N_9949,N_9910);
and UO_276 (O_276,N_9948,N_9933);
or UO_277 (O_277,N_9967,N_9952);
or UO_278 (O_278,N_9921,N_9975);
and UO_279 (O_279,N_9917,N_9934);
nand UO_280 (O_280,N_9946,N_9982);
nand UO_281 (O_281,N_9913,N_9921);
and UO_282 (O_282,N_9921,N_9909);
nor UO_283 (O_283,N_9936,N_9950);
nand UO_284 (O_284,N_9926,N_9970);
and UO_285 (O_285,N_9944,N_9966);
and UO_286 (O_286,N_9943,N_9920);
nand UO_287 (O_287,N_9943,N_9901);
or UO_288 (O_288,N_9976,N_9920);
and UO_289 (O_289,N_9903,N_9915);
or UO_290 (O_290,N_9992,N_9945);
xor UO_291 (O_291,N_9921,N_9991);
nor UO_292 (O_292,N_9988,N_9997);
nor UO_293 (O_293,N_9976,N_9954);
or UO_294 (O_294,N_9962,N_9976);
and UO_295 (O_295,N_9968,N_9976);
nand UO_296 (O_296,N_9909,N_9920);
and UO_297 (O_297,N_9955,N_9988);
nor UO_298 (O_298,N_9962,N_9949);
nor UO_299 (O_299,N_9935,N_9962);
nand UO_300 (O_300,N_9949,N_9976);
nor UO_301 (O_301,N_9946,N_9984);
nor UO_302 (O_302,N_9954,N_9925);
nor UO_303 (O_303,N_9907,N_9938);
nand UO_304 (O_304,N_9977,N_9912);
or UO_305 (O_305,N_9913,N_9972);
nor UO_306 (O_306,N_9929,N_9960);
nor UO_307 (O_307,N_9918,N_9968);
and UO_308 (O_308,N_9953,N_9954);
nand UO_309 (O_309,N_9992,N_9960);
and UO_310 (O_310,N_9985,N_9902);
and UO_311 (O_311,N_9964,N_9946);
or UO_312 (O_312,N_9954,N_9988);
nor UO_313 (O_313,N_9924,N_9922);
or UO_314 (O_314,N_9958,N_9971);
nor UO_315 (O_315,N_9990,N_9931);
or UO_316 (O_316,N_9958,N_9991);
nor UO_317 (O_317,N_9927,N_9991);
nor UO_318 (O_318,N_9998,N_9901);
or UO_319 (O_319,N_9942,N_9945);
nor UO_320 (O_320,N_9941,N_9959);
nor UO_321 (O_321,N_9981,N_9919);
nor UO_322 (O_322,N_9957,N_9901);
and UO_323 (O_323,N_9941,N_9989);
and UO_324 (O_324,N_9967,N_9996);
nor UO_325 (O_325,N_9952,N_9992);
and UO_326 (O_326,N_9918,N_9925);
and UO_327 (O_327,N_9943,N_9953);
and UO_328 (O_328,N_9993,N_9949);
nor UO_329 (O_329,N_9944,N_9947);
or UO_330 (O_330,N_9929,N_9976);
nand UO_331 (O_331,N_9998,N_9942);
and UO_332 (O_332,N_9924,N_9998);
or UO_333 (O_333,N_9926,N_9996);
nand UO_334 (O_334,N_9956,N_9970);
nand UO_335 (O_335,N_9954,N_9977);
nand UO_336 (O_336,N_9973,N_9958);
or UO_337 (O_337,N_9966,N_9967);
xnor UO_338 (O_338,N_9965,N_9944);
nor UO_339 (O_339,N_9968,N_9965);
nand UO_340 (O_340,N_9963,N_9958);
or UO_341 (O_341,N_9972,N_9932);
and UO_342 (O_342,N_9988,N_9919);
nor UO_343 (O_343,N_9904,N_9906);
or UO_344 (O_344,N_9996,N_9938);
and UO_345 (O_345,N_9973,N_9989);
and UO_346 (O_346,N_9916,N_9967);
or UO_347 (O_347,N_9948,N_9960);
and UO_348 (O_348,N_9981,N_9935);
and UO_349 (O_349,N_9920,N_9938);
or UO_350 (O_350,N_9967,N_9990);
and UO_351 (O_351,N_9934,N_9952);
nor UO_352 (O_352,N_9955,N_9935);
nor UO_353 (O_353,N_9993,N_9997);
nor UO_354 (O_354,N_9995,N_9934);
nand UO_355 (O_355,N_9990,N_9981);
nand UO_356 (O_356,N_9966,N_9960);
nor UO_357 (O_357,N_9995,N_9925);
nand UO_358 (O_358,N_9932,N_9906);
or UO_359 (O_359,N_9946,N_9974);
xor UO_360 (O_360,N_9999,N_9934);
nor UO_361 (O_361,N_9927,N_9915);
nand UO_362 (O_362,N_9968,N_9949);
or UO_363 (O_363,N_9968,N_9931);
and UO_364 (O_364,N_9941,N_9920);
and UO_365 (O_365,N_9903,N_9919);
and UO_366 (O_366,N_9904,N_9923);
or UO_367 (O_367,N_9913,N_9960);
nand UO_368 (O_368,N_9928,N_9978);
or UO_369 (O_369,N_9978,N_9975);
and UO_370 (O_370,N_9971,N_9955);
nor UO_371 (O_371,N_9905,N_9931);
nor UO_372 (O_372,N_9987,N_9942);
nand UO_373 (O_373,N_9915,N_9934);
nand UO_374 (O_374,N_9949,N_9965);
nor UO_375 (O_375,N_9935,N_9902);
nand UO_376 (O_376,N_9940,N_9958);
or UO_377 (O_377,N_9917,N_9949);
or UO_378 (O_378,N_9975,N_9967);
and UO_379 (O_379,N_9998,N_9986);
nand UO_380 (O_380,N_9965,N_9982);
nor UO_381 (O_381,N_9907,N_9912);
or UO_382 (O_382,N_9911,N_9929);
nor UO_383 (O_383,N_9945,N_9923);
nand UO_384 (O_384,N_9989,N_9975);
or UO_385 (O_385,N_9906,N_9930);
or UO_386 (O_386,N_9951,N_9920);
nor UO_387 (O_387,N_9958,N_9953);
nor UO_388 (O_388,N_9933,N_9949);
or UO_389 (O_389,N_9904,N_9971);
and UO_390 (O_390,N_9943,N_9981);
xor UO_391 (O_391,N_9982,N_9996);
and UO_392 (O_392,N_9961,N_9996);
nor UO_393 (O_393,N_9911,N_9960);
or UO_394 (O_394,N_9992,N_9950);
or UO_395 (O_395,N_9967,N_9931);
xor UO_396 (O_396,N_9968,N_9953);
and UO_397 (O_397,N_9907,N_9945);
or UO_398 (O_398,N_9904,N_9984);
xor UO_399 (O_399,N_9907,N_9914);
nand UO_400 (O_400,N_9980,N_9901);
and UO_401 (O_401,N_9946,N_9905);
nor UO_402 (O_402,N_9994,N_9910);
nand UO_403 (O_403,N_9987,N_9951);
or UO_404 (O_404,N_9901,N_9912);
or UO_405 (O_405,N_9937,N_9978);
and UO_406 (O_406,N_9995,N_9970);
nor UO_407 (O_407,N_9938,N_9994);
and UO_408 (O_408,N_9951,N_9988);
and UO_409 (O_409,N_9994,N_9997);
nor UO_410 (O_410,N_9913,N_9903);
nand UO_411 (O_411,N_9986,N_9954);
nand UO_412 (O_412,N_9924,N_9951);
nand UO_413 (O_413,N_9991,N_9970);
or UO_414 (O_414,N_9951,N_9948);
and UO_415 (O_415,N_9900,N_9974);
or UO_416 (O_416,N_9986,N_9958);
nand UO_417 (O_417,N_9979,N_9988);
xnor UO_418 (O_418,N_9951,N_9978);
nor UO_419 (O_419,N_9959,N_9913);
nand UO_420 (O_420,N_9915,N_9937);
or UO_421 (O_421,N_9938,N_9909);
and UO_422 (O_422,N_9931,N_9980);
nor UO_423 (O_423,N_9927,N_9961);
and UO_424 (O_424,N_9998,N_9968);
or UO_425 (O_425,N_9981,N_9945);
and UO_426 (O_426,N_9913,N_9917);
nand UO_427 (O_427,N_9992,N_9994);
nand UO_428 (O_428,N_9998,N_9988);
nand UO_429 (O_429,N_9924,N_9912);
nor UO_430 (O_430,N_9996,N_9922);
and UO_431 (O_431,N_9988,N_9973);
and UO_432 (O_432,N_9955,N_9978);
or UO_433 (O_433,N_9943,N_9932);
or UO_434 (O_434,N_9976,N_9994);
or UO_435 (O_435,N_9990,N_9980);
and UO_436 (O_436,N_9966,N_9973);
and UO_437 (O_437,N_9964,N_9996);
xnor UO_438 (O_438,N_9959,N_9920);
and UO_439 (O_439,N_9920,N_9942);
nor UO_440 (O_440,N_9961,N_9924);
nand UO_441 (O_441,N_9968,N_9922);
nor UO_442 (O_442,N_9911,N_9983);
nand UO_443 (O_443,N_9926,N_9901);
or UO_444 (O_444,N_9985,N_9956);
and UO_445 (O_445,N_9946,N_9940);
and UO_446 (O_446,N_9960,N_9910);
nand UO_447 (O_447,N_9985,N_9984);
xnor UO_448 (O_448,N_9960,N_9921);
and UO_449 (O_449,N_9900,N_9934);
xor UO_450 (O_450,N_9950,N_9970);
and UO_451 (O_451,N_9983,N_9923);
nor UO_452 (O_452,N_9990,N_9937);
nor UO_453 (O_453,N_9989,N_9987);
or UO_454 (O_454,N_9997,N_9916);
nand UO_455 (O_455,N_9990,N_9965);
and UO_456 (O_456,N_9958,N_9966);
nand UO_457 (O_457,N_9969,N_9939);
nand UO_458 (O_458,N_9964,N_9991);
and UO_459 (O_459,N_9931,N_9935);
nor UO_460 (O_460,N_9905,N_9923);
or UO_461 (O_461,N_9991,N_9900);
and UO_462 (O_462,N_9988,N_9926);
nor UO_463 (O_463,N_9970,N_9915);
or UO_464 (O_464,N_9977,N_9983);
or UO_465 (O_465,N_9958,N_9996);
nand UO_466 (O_466,N_9917,N_9980);
or UO_467 (O_467,N_9956,N_9957);
nor UO_468 (O_468,N_9977,N_9937);
and UO_469 (O_469,N_9973,N_9913);
xor UO_470 (O_470,N_9901,N_9942);
and UO_471 (O_471,N_9965,N_9984);
and UO_472 (O_472,N_9957,N_9967);
or UO_473 (O_473,N_9929,N_9921);
nand UO_474 (O_474,N_9938,N_9957);
nand UO_475 (O_475,N_9962,N_9974);
or UO_476 (O_476,N_9968,N_9907);
and UO_477 (O_477,N_9951,N_9958);
nand UO_478 (O_478,N_9961,N_9979);
and UO_479 (O_479,N_9963,N_9936);
nand UO_480 (O_480,N_9993,N_9915);
or UO_481 (O_481,N_9981,N_9976);
xor UO_482 (O_482,N_9932,N_9963);
and UO_483 (O_483,N_9987,N_9925);
or UO_484 (O_484,N_9950,N_9943);
and UO_485 (O_485,N_9938,N_9999);
and UO_486 (O_486,N_9992,N_9988);
nor UO_487 (O_487,N_9959,N_9963);
nor UO_488 (O_488,N_9937,N_9924);
nand UO_489 (O_489,N_9922,N_9906);
and UO_490 (O_490,N_9984,N_9927);
nand UO_491 (O_491,N_9917,N_9985);
nand UO_492 (O_492,N_9961,N_9951);
nor UO_493 (O_493,N_9933,N_9900);
nand UO_494 (O_494,N_9986,N_9941);
nand UO_495 (O_495,N_9989,N_9912);
nor UO_496 (O_496,N_9900,N_9992);
nor UO_497 (O_497,N_9903,N_9927);
nor UO_498 (O_498,N_9978,N_9923);
and UO_499 (O_499,N_9969,N_9908);
and UO_500 (O_500,N_9989,N_9953);
or UO_501 (O_501,N_9932,N_9958);
or UO_502 (O_502,N_9930,N_9976);
nor UO_503 (O_503,N_9982,N_9998);
or UO_504 (O_504,N_9978,N_9980);
nand UO_505 (O_505,N_9990,N_9961);
nor UO_506 (O_506,N_9970,N_9990);
nand UO_507 (O_507,N_9943,N_9962);
or UO_508 (O_508,N_9946,N_9959);
or UO_509 (O_509,N_9991,N_9969);
and UO_510 (O_510,N_9997,N_9969);
or UO_511 (O_511,N_9964,N_9980);
and UO_512 (O_512,N_9944,N_9963);
and UO_513 (O_513,N_9966,N_9936);
or UO_514 (O_514,N_9978,N_9920);
or UO_515 (O_515,N_9908,N_9927);
xnor UO_516 (O_516,N_9934,N_9988);
or UO_517 (O_517,N_9932,N_9910);
nor UO_518 (O_518,N_9973,N_9923);
and UO_519 (O_519,N_9930,N_9995);
and UO_520 (O_520,N_9992,N_9907);
and UO_521 (O_521,N_9966,N_9978);
nor UO_522 (O_522,N_9950,N_9959);
or UO_523 (O_523,N_9959,N_9943);
and UO_524 (O_524,N_9947,N_9907);
or UO_525 (O_525,N_9983,N_9949);
and UO_526 (O_526,N_9994,N_9956);
nand UO_527 (O_527,N_9948,N_9958);
nor UO_528 (O_528,N_9961,N_9939);
nor UO_529 (O_529,N_9945,N_9988);
and UO_530 (O_530,N_9945,N_9977);
nor UO_531 (O_531,N_9936,N_9910);
nand UO_532 (O_532,N_9939,N_9910);
and UO_533 (O_533,N_9906,N_9964);
or UO_534 (O_534,N_9953,N_9941);
and UO_535 (O_535,N_9977,N_9938);
or UO_536 (O_536,N_9918,N_9948);
and UO_537 (O_537,N_9912,N_9935);
or UO_538 (O_538,N_9916,N_9960);
or UO_539 (O_539,N_9932,N_9914);
and UO_540 (O_540,N_9962,N_9999);
and UO_541 (O_541,N_9925,N_9908);
or UO_542 (O_542,N_9994,N_9993);
or UO_543 (O_543,N_9972,N_9951);
nand UO_544 (O_544,N_9906,N_9968);
nor UO_545 (O_545,N_9932,N_9952);
xor UO_546 (O_546,N_9959,N_9929);
or UO_547 (O_547,N_9946,N_9938);
nor UO_548 (O_548,N_9909,N_9983);
or UO_549 (O_549,N_9977,N_9940);
or UO_550 (O_550,N_9916,N_9930);
or UO_551 (O_551,N_9903,N_9943);
or UO_552 (O_552,N_9973,N_9925);
and UO_553 (O_553,N_9942,N_9900);
nand UO_554 (O_554,N_9926,N_9951);
nor UO_555 (O_555,N_9927,N_9982);
and UO_556 (O_556,N_9923,N_9980);
and UO_557 (O_557,N_9970,N_9959);
nor UO_558 (O_558,N_9985,N_9921);
or UO_559 (O_559,N_9995,N_9921);
nor UO_560 (O_560,N_9954,N_9904);
and UO_561 (O_561,N_9908,N_9922);
or UO_562 (O_562,N_9905,N_9929);
and UO_563 (O_563,N_9924,N_9970);
nor UO_564 (O_564,N_9920,N_9990);
or UO_565 (O_565,N_9954,N_9932);
and UO_566 (O_566,N_9979,N_9971);
and UO_567 (O_567,N_9973,N_9930);
or UO_568 (O_568,N_9901,N_9985);
nor UO_569 (O_569,N_9994,N_9900);
or UO_570 (O_570,N_9914,N_9951);
nor UO_571 (O_571,N_9997,N_9947);
and UO_572 (O_572,N_9988,N_9936);
or UO_573 (O_573,N_9936,N_9954);
or UO_574 (O_574,N_9980,N_9949);
and UO_575 (O_575,N_9968,N_9924);
nand UO_576 (O_576,N_9992,N_9951);
nor UO_577 (O_577,N_9996,N_9917);
nand UO_578 (O_578,N_9915,N_9919);
or UO_579 (O_579,N_9971,N_9964);
and UO_580 (O_580,N_9978,N_9941);
and UO_581 (O_581,N_9906,N_9999);
nand UO_582 (O_582,N_9900,N_9941);
and UO_583 (O_583,N_9955,N_9901);
nor UO_584 (O_584,N_9907,N_9983);
nor UO_585 (O_585,N_9920,N_9979);
nand UO_586 (O_586,N_9969,N_9950);
or UO_587 (O_587,N_9985,N_9928);
and UO_588 (O_588,N_9981,N_9908);
and UO_589 (O_589,N_9928,N_9988);
or UO_590 (O_590,N_9933,N_9937);
and UO_591 (O_591,N_9930,N_9948);
nor UO_592 (O_592,N_9984,N_9933);
nor UO_593 (O_593,N_9986,N_9937);
and UO_594 (O_594,N_9959,N_9911);
nor UO_595 (O_595,N_9904,N_9941);
nand UO_596 (O_596,N_9967,N_9968);
or UO_597 (O_597,N_9971,N_9976);
xor UO_598 (O_598,N_9910,N_9929);
nand UO_599 (O_599,N_9946,N_9925);
and UO_600 (O_600,N_9905,N_9957);
or UO_601 (O_601,N_9962,N_9911);
nor UO_602 (O_602,N_9906,N_9956);
and UO_603 (O_603,N_9988,N_9920);
xor UO_604 (O_604,N_9986,N_9938);
or UO_605 (O_605,N_9907,N_9979);
or UO_606 (O_606,N_9930,N_9910);
and UO_607 (O_607,N_9936,N_9917);
or UO_608 (O_608,N_9934,N_9935);
and UO_609 (O_609,N_9951,N_9906);
or UO_610 (O_610,N_9932,N_9997);
nor UO_611 (O_611,N_9920,N_9932);
or UO_612 (O_612,N_9994,N_9962);
nand UO_613 (O_613,N_9965,N_9999);
nor UO_614 (O_614,N_9954,N_9980);
or UO_615 (O_615,N_9900,N_9997);
or UO_616 (O_616,N_9996,N_9960);
or UO_617 (O_617,N_9932,N_9988);
nor UO_618 (O_618,N_9957,N_9983);
or UO_619 (O_619,N_9931,N_9936);
or UO_620 (O_620,N_9920,N_9901);
nor UO_621 (O_621,N_9926,N_9911);
nor UO_622 (O_622,N_9993,N_9938);
nand UO_623 (O_623,N_9990,N_9954);
or UO_624 (O_624,N_9954,N_9993);
nand UO_625 (O_625,N_9953,N_9993);
nand UO_626 (O_626,N_9979,N_9973);
or UO_627 (O_627,N_9921,N_9940);
nor UO_628 (O_628,N_9978,N_9927);
nand UO_629 (O_629,N_9943,N_9977);
nand UO_630 (O_630,N_9941,N_9956);
and UO_631 (O_631,N_9941,N_9934);
or UO_632 (O_632,N_9904,N_9974);
or UO_633 (O_633,N_9970,N_9903);
nand UO_634 (O_634,N_9929,N_9913);
and UO_635 (O_635,N_9907,N_9948);
or UO_636 (O_636,N_9968,N_9989);
nor UO_637 (O_637,N_9998,N_9921);
nor UO_638 (O_638,N_9950,N_9926);
nand UO_639 (O_639,N_9906,N_9954);
nor UO_640 (O_640,N_9939,N_9927);
and UO_641 (O_641,N_9990,N_9960);
or UO_642 (O_642,N_9922,N_9990);
nand UO_643 (O_643,N_9978,N_9938);
nor UO_644 (O_644,N_9977,N_9976);
and UO_645 (O_645,N_9904,N_9920);
or UO_646 (O_646,N_9959,N_9958);
nor UO_647 (O_647,N_9947,N_9974);
or UO_648 (O_648,N_9931,N_9986);
nor UO_649 (O_649,N_9961,N_9946);
nor UO_650 (O_650,N_9943,N_9969);
nand UO_651 (O_651,N_9962,N_9903);
nand UO_652 (O_652,N_9962,N_9908);
nor UO_653 (O_653,N_9945,N_9903);
and UO_654 (O_654,N_9929,N_9986);
or UO_655 (O_655,N_9956,N_9976);
nor UO_656 (O_656,N_9902,N_9968);
nand UO_657 (O_657,N_9904,N_9909);
nor UO_658 (O_658,N_9954,N_9927);
nand UO_659 (O_659,N_9988,N_9966);
nor UO_660 (O_660,N_9990,N_9998);
nor UO_661 (O_661,N_9936,N_9981);
and UO_662 (O_662,N_9940,N_9929);
nand UO_663 (O_663,N_9948,N_9993);
nor UO_664 (O_664,N_9997,N_9953);
and UO_665 (O_665,N_9906,N_9978);
or UO_666 (O_666,N_9968,N_9938);
nor UO_667 (O_667,N_9968,N_9970);
nor UO_668 (O_668,N_9914,N_9961);
nand UO_669 (O_669,N_9975,N_9994);
nand UO_670 (O_670,N_9983,N_9924);
nor UO_671 (O_671,N_9903,N_9950);
or UO_672 (O_672,N_9953,N_9996);
or UO_673 (O_673,N_9982,N_9921);
or UO_674 (O_674,N_9991,N_9944);
nor UO_675 (O_675,N_9916,N_9926);
nor UO_676 (O_676,N_9953,N_9978);
nand UO_677 (O_677,N_9989,N_9979);
and UO_678 (O_678,N_9924,N_9971);
nor UO_679 (O_679,N_9923,N_9902);
nor UO_680 (O_680,N_9948,N_9913);
nor UO_681 (O_681,N_9928,N_9964);
or UO_682 (O_682,N_9973,N_9991);
and UO_683 (O_683,N_9983,N_9955);
nor UO_684 (O_684,N_9999,N_9959);
and UO_685 (O_685,N_9919,N_9924);
nor UO_686 (O_686,N_9921,N_9979);
or UO_687 (O_687,N_9906,N_9937);
and UO_688 (O_688,N_9965,N_9972);
xor UO_689 (O_689,N_9939,N_9974);
and UO_690 (O_690,N_9925,N_9977);
nand UO_691 (O_691,N_9902,N_9966);
nor UO_692 (O_692,N_9957,N_9979);
nor UO_693 (O_693,N_9906,N_9997);
nor UO_694 (O_694,N_9975,N_9983);
nor UO_695 (O_695,N_9920,N_9984);
or UO_696 (O_696,N_9933,N_9950);
nor UO_697 (O_697,N_9936,N_9940);
nor UO_698 (O_698,N_9955,N_9924);
or UO_699 (O_699,N_9938,N_9917);
or UO_700 (O_700,N_9954,N_9991);
or UO_701 (O_701,N_9928,N_9910);
nand UO_702 (O_702,N_9942,N_9924);
and UO_703 (O_703,N_9987,N_9954);
and UO_704 (O_704,N_9925,N_9970);
xor UO_705 (O_705,N_9999,N_9910);
nand UO_706 (O_706,N_9926,N_9937);
xnor UO_707 (O_707,N_9929,N_9930);
nor UO_708 (O_708,N_9959,N_9955);
nor UO_709 (O_709,N_9921,N_9981);
and UO_710 (O_710,N_9947,N_9953);
xnor UO_711 (O_711,N_9988,N_9933);
or UO_712 (O_712,N_9940,N_9961);
nor UO_713 (O_713,N_9981,N_9998);
nand UO_714 (O_714,N_9962,N_9963);
nand UO_715 (O_715,N_9974,N_9936);
or UO_716 (O_716,N_9913,N_9975);
and UO_717 (O_717,N_9945,N_9953);
nand UO_718 (O_718,N_9977,N_9990);
nand UO_719 (O_719,N_9969,N_9971);
nor UO_720 (O_720,N_9995,N_9935);
nor UO_721 (O_721,N_9932,N_9913);
and UO_722 (O_722,N_9931,N_9998);
nor UO_723 (O_723,N_9900,N_9952);
nor UO_724 (O_724,N_9985,N_9990);
nor UO_725 (O_725,N_9924,N_9990);
nor UO_726 (O_726,N_9987,N_9958);
nor UO_727 (O_727,N_9964,N_9968);
nand UO_728 (O_728,N_9964,N_9932);
or UO_729 (O_729,N_9966,N_9954);
nand UO_730 (O_730,N_9932,N_9949);
nor UO_731 (O_731,N_9926,N_9918);
nand UO_732 (O_732,N_9904,N_9989);
nand UO_733 (O_733,N_9967,N_9918);
nand UO_734 (O_734,N_9951,N_9995);
nor UO_735 (O_735,N_9954,N_9926);
nand UO_736 (O_736,N_9979,N_9931);
nor UO_737 (O_737,N_9925,N_9909);
or UO_738 (O_738,N_9957,N_9970);
or UO_739 (O_739,N_9975,N_9964);
nor UO_740 (O_740,N_9968,N_9980);
or UO_741 (O_741,N_9969,N_9911);
or UO_742 (O_742,N_9970,N_9976);
nand UO_743 (O_743,N_9947,N_9962);
nand UO_744 (O_744,N_9945,N_9909);
nand UO_745 (O_745,N_9910,N_9950);
or UO_746 (O_746,N_9932,N_9966);
nor UO_747 (O_747,N_9910,N_9912);
nand UO_748 (O_748,N_9907,N_9991);
or UO_749 (O_749,N_9913,N_9906);
and UO_750 (O_750,N_9975,N_9901);
and UO_751 (O_751,N_9916,N_9903);
nor UO_752 (O_752,N_9917,N_9956);
or UO_753 (O_753,N_9973,N_9918);
or UO_754 (O_754,N_9991,N_9981);
nor UO_755 (O_755,N_9915,N_9964);
nand UO_756 (O_756,N_9949,N_9929);
and UO_757 (O_757,N_9995,N_9958);
nand UO_758 (O_758,N_9975,N_9939);
or UO_759 (O_759,N_9948,N_9926);
or UO_760 (O_760,N_9967,N_9973);
or UO_761 (O_761,N_9920,N_9964);
nor UO_762 (O_762,N_9994,N_9937);
or UO_763 (O_763,N_9969,N_9993);
and UO_764 (O_764,N_9964,N_9969);
nand UO_765 (O_765,N_9964,N_9995);
nand UO_766 (O_766,N_9967,N_9924);
and UO_767 (O_767,N_9972,N_9911);
nor UO_768 (O_768,N_9980,N_9969);
nand UO_769 (O_769,N_9961,N_9958);
and UO_770 (O_770,N_9996,N_9916);
xor UO_771 (O_771,N_9998,N_9994);
and UO_772 (O_772,N_9988,N_9908);
and UO_773 (O_773,N_9990,N_9969);
and UO_774 (O_774,N_9995,N_9978);
or UO_775 (O_775,N_9955,N_9937);
or UO_776 (O_776,N_9985,N_9991);
nor UO_777 (O_777,N_9916,N_9972);
nor UO_778 (O_778,N_9963,N_9906);
and UO_779 (O_779,N_9982,N_9995);
xnor UO_780 (O_780,N_9914,N_9925);
or UO_781 (O_781,N_9941,N_9988);
nor UO_782 (O_782,N_9901,N_9968);
nand UO_783 (O_783,N_9913,N_9998);
nand UO_784 (O_784,N_9945,N_9991);
xnor UO_785 (O_785,N_9924,N_9952);
nor UO_786 (O_786,N_9901,N_9989);
and UO_787 (O_787,N_9969,N_9956);
or UO_788 (O_788,N_9948,N_9914);
and UO_789 (O_789,N_9959,N_9968);
or UO_790 (O_790,N_9999,N_9916);
and UO_791 (O_791,N_9932,N_9978);
nand UO_792 (O_792,N_9980,N_9984);
or UO_793 (O_793,N_9909,N_9922);
and UO_794 (O_794,N_9990,N_9909);
nand UO_795 (O_795,N_9965,N_9963);
or UO_796 (O_796,N_9920,N_9933);
or UO_797 (O_797,N_9949,N_9995);
nand UO_798 (O_798,N_9935,N_9964);
and UO_799 (O_799,N_9989,N_9960);
nor UO_800 (O_800,N_9970,N_9907);
or UO_801 (O_801,N_9935,N_9910);
and UO_802 (O_802,N_9986,N_9967);
or UO_803 (O_803,N_9940,N_9900);
nand UO_804 (O_804,N_9919,N_9957);
nor UO_805 (O_805,N_9966,N_9991);
and UO_806 (O_806,N_9995,N_9989);
nor UO_807 (O_807,N_9902,N_9934);
or UO_808 (O_808,N_9912,N_9939);
and UO_809 (O_809,N_9940,N_9949);
nand UO_810 (O_810,N_9905,N_9900);
nand UO_811 (O_811,N_9940,N_9984);
nor UO_812 (O_812,N_9953,N_9934);
nand UO_813 (O_813,N_9998,N_9917);
nand UO_814 (O_814,N_9999,N_9918);
or UO_815 (O_815,N_9918,N_9904);
or UO_816 (O_816,N_9926,N_9913);
nor UO_817 (O_817,N_9964,N_9905);
and UO_818 (O_818,N_9972,N_9973);
nand UO_819 (O_819,N_9963,N_9926);
xnor UO_820 (O_820,N_9973,N_9902);
or UO_821 (O_821,N_9925,N_9949);
nor UO_822 (O_822,N_9999,N_9987);
and UO_823 (O_823,N_9971,N_9948);
and UO_824 (O_824,N_9936,N_9905);
or UO_825 (O_825,N_9998,N_9965);
and UO_826 (O_826,N_9948,N_9919);
or UO_827 (O_827,N_9959,N_9924);
nand UO_828 (O_828,N_9955,N_9938);
and UO_829 (O_829,N_9944,N_9921);
or UO_830 (O_830,N_9944,N_9995);
and UO_831 (O_831,N_9907,N_9951);
or UO_832 (O_832,N_9961,N_9922);
nor UO_833 (O_833,N_9948,N_9974);
nor UO_834 (O_834,N_9901,N_9995);
nand UO_835 (O_835,N_9998,N_9987);
nand UO_836 (O_836,N_9917,N_9974);
and UO_837 (O_837,N_9940,N_9901);
or UO_838 (O_838,N_9928,N_9984);
and UO_839 (O_839,N_9971,N_9963);
nand UO_840 (O_840,N_9963,N_9943);
and UO_841 (O_841,N_9909,N_9988);
nand UO_842 (O_842,N_9980,N_9985);
nor UO_843 (O_843,N_9921,N_9939);
nor UO_844 (O_844,N_9977,N_9936);
or UO_845 (O_845,N_9957,N_9988);
or UO_846 (O_846,N_9900,N_9965);
and UO_847 (O_847,N_9907,N_9973);
or UO_848 (O_848,N_9952,N_9950);
nand UO_849 (O_849,N_9929,N_9927);
nand UO_850 (O_850,N_9982,N_9952);
and UO_851 (O_851,N_9962,N_9969);
nand UO_852 (O_852,N_9957,N_9969);
nand UO_853 (O_853,N_9910,N_9981);
nand UO_854 (O_854,N_9911,N_9917);
nand UO_855 (O_855,N_9975,N_9918);
nand UO_856 (O_856,N_9930,N_9926);
nand UO_857 (O_857,N_9986,N_9971);
or UO_858 (O_858,N_9968,N_9913);
and UO_859 (O_859,N_9952,N_9922);
and UO_860 (O_860,N_9993,N_9989);
and UO_861 (O_861,N_9959,N_9949);
or UO_862 (O_862,N_9922,N_9919);
and UO_863 (O_863,N_9939,N_9909);
xnor UO_864 (O_864,N_9920,N_9975);
and UO_865 (O_865,N_9955,N_9951);
nor UO_866 (O_866,N_9908,N_9904);
and UO_867 (O_867,N_9900,N_9961);
or UO_868 (O_868,N_9966,N_9997);
or UO_869 (O_869,N_9928,N_9909);
or UO_870 (O_870,N_9942,N_9969);
and UO_871 (O_871,N_9995,N_9953);
or UO_872 (O_872,N_9922,N_9995);
nor UO_873 (O_873,N_9952,N_9953);
and UO_874 (O_874,N_9929,N_9985);
nand UO_875 (O_875,N_9953,N_9962);
or UO_876 (O_876,N_9976,N_9967);
and UO_877 (O_877,N_9939,N_9933);
nand UO_878 (O_878,N_9939,N_9900);
nor UO_879 (O_879,N_9921,N_9945);
nor UO_880 (O_880,N_9936,N_9933);
nand UO_881 (O_881,N_9999,N_9953);
or UO_882 (O_882,N_9990,N_9984);
nand UO_883 (O_883,N_9930,N_9919);
nor UO_884 (O_884,N_9914,N_9957);
and UO_885 (O_885,N_9985,N_9900);
or UO_886 (O_886,N_9983,N_9938);
nand UO_887 (O_887,N_9910,N_9948);
nand UO_888 (O_888,N_9992,N_9990);
nor UO_889 (O_889,N_9943,N_9946);
nand UO_890 (O_890,N_9968,N_9911);
nor UO_891 (O_891,N_9960,N_9991);
nor UO_892 (O_892,N_9904,N_9900);
or UO_893 (O_893,N_9954,N_9923);
nand UO_894 (O_894,N_9999,N_9966);
and UO_895 (O_895,N_9939,N_9997);
or UO_896 (O_896,N_9951,N_9911);
nor UO_897 (O_897,N_9975,N_9941);
and UO_898 (O_898,N_9930,N_9925);
or UO_899 (O_899,N_9905,N_9951);
nor UO_900 (O_900,N_9966,N_9965);
nand UO_901 (O_901,N_9935,N_9907);
nand UO_902 (O_902,N_9941,N_9980);
and UO_903 (O_903,N_9983,N_9984);
nor UO_904 (O_904,N_9968,N_9945);
or UO_905 (O_905,N_9957,N_9913);
or UO_906 (O_906,N_9973,N_9954);
and UO_907 (O_907,N_9979,N_9946);
and UO_908 (O_908,N_9949,N_9952);
nor UO_909 (O_909,N_9901,N_9977);
and UO_910 (O_910,N_9943,N_9955);
and UO_911 (O_911,N_9944,N_9929);
nand UO_912 (O_912,N_9951,N_9973);
nand UO_913 (O_913,N_9965,N_9945);
or UO_914 (O_914,N_9921,N_9994);
or UO_915 (O_915,N_9931,N_9955);
nand UO_916 (O_916,N_9997,N_9951);
nand UO_917 (O_917,N_9998,N_9963);
and UO_918 (O_918,N_9989,N_9962);
nand UO_919 (O_919,N_9925,N_9980);
and UO_920 (O_920,N_9907,N_9922);
nand UO_921 (O_921,N_9961,N_9929);
and UO_922 (O_922,N_9971,N_9934);
and UO_923 (O_923,N_9906,N_9918);
and UO_924 (O_924,N_9972,N_9912);
and UO_925 (O_925,N_9960,N_9957);
or UO_926 (O_926,N_9935,N_9922);
nor UO_927 (O_927,N_9905,N_9950);
nor UO_928 (O_928,N_9982,N_9993);
nor UO_929 (O_929,N_9914,N_9945);
and UO_930 (O_930,N_9920,N_9992);
or UO_931 (O_931,N_9997,N_9961);
xor UO_932 (O_932,N_9942,N_9962);
nor UO_933 (O_933,N_9993,N_9974);
xor UO_934 (O_934,N_9947,N_9973);
or UO_935 (O_935,N_9953,N_9988);
or UO_936 (O_936,N_9914,N_9973);
and UO_937 (O_937,N_9902,N_9948);
or UO_938 (O_938,N_9943,N_9980);
and UO_939 (O_939,N_9987,N_9969);
and UO_940 (O_940,N_9979,N_9928);
nor UO_941 (O_941,N_9912,N_9934);
or UO_942 (O_942,N_9944,N_9939);
or UO_943 (O_943,N_9986,N_9972);
nand UO_944 (O_944,N_9931,N_9987);
or UO_945 (O_945,N_9914,N_9970);
nor UO_946 (O_946,N_9972,N_9926);
nand UO_947 (O_947,N_9970,N_9999);
or UO_948 (O_948,N_9976,N_9969);
nand UO_949 (O_949,N_9910,N_9904);
nand UO_950 (O_950,N_9963,N_9939);
or UO_951 (O_951,N_9915,N_9981);
and UO_952 (O_952,N_9945,N_9930);
nor UO_953 (O_953,N_9938,N_9937);
or UO_954 (O_954,N_9965,N_9901);
nand UO_955 (O_955,N_9927,N_9936);
or UO_956 (O_956,N_9959,N_9922);
and UO_957 (O_957,N_9977,N_9959);
and UO_958 (O_958,N_9909,N_9985);
and UO_959 (O_959,N_9952,N_9966);
and UO_960 (O_960,N_9980,N_9940);
or UO_961 (O_961,N_9991,N_9931);
or UO_962 (O_962,N_9951,N_9990);
or UO_963 (O_963,N_9939,N_9934);
nand UO_964 (O_964,N_9929,N_9951);
and UO_965 (O_965,N_9964,N_9901);
nor UO_966 (O_966,N_9927,N_9943);
nand UO_967 (O_967,N_9957,N_9973);
nand UO_968 (O_968,N_9919,N_9918);
and UO_969 (O_969,N_9960,N_9938);
nor UO_970 (O_970,N_9929,N_9998);
nand UO_971 (O_971,N_9949,N_9937);
nor UO_972 (O_972,N_9901,N_9961);
or UO_973 (O_973,N_9949,N_9981);
or UO_974 (O_974,N_9963,N_9979);
or UO_975 (O_975,N_9977,N_9955);
and UO_976 (O_976,N_9909,N_9989);
nor UO_977 (O_977,N_9928,N_9999);
or UO_978 (O_978,N_9914,N_9990);
or UO_979 (O_979,N_9945,N_9931);
nor UO_980 (O_980,N_9908,N_9992);
and UO_981 (O_981,N_9950,N_9942);
or UO_982 (O_982,N_9948,N_9940);
nor UO_983 (O_983,N_9990,N_9963);
nor UO_984 (O_984,N_9920,N_9917);
or UO_985 (O_985,N_9972,N_9927);
nand UO_986 (O_986,N_9927,N_9976);
and UO_987 (O_987,N_9942,N_9951);
and UO_988 (O_988,N_9935,N_9901);
and UO_989 (O_989,N_9956,N_9916);
and UO_990 (O_990,N_9943,N_9928);
and UO_991 (O_991,N_9964,N_9934);
nor UO_992 (O_992,N_9995,N_9920);
and UO_993 (O_993,N_9928,N_9976);
nor UO_994 (O_994,N_9940,N_9987);
nor UO_995 (O_995,N_9952,N_9987);
or UO_996 (O_996,N_9994,N_9942);
or UO_997 (O_997,N_9919,N_9998);
or UO_998 (O_998,N_9912,N_9936);
and UO_999 (O_999,N_9911,N_9966);
or UO_1000 (O_1000,N_9975,N_9931);
nor UO_1001 (O_1001,N_9986,N_9983);
nand UO_1002 (O_1002,N_9917,N_9951);
and UO_1003 (O_1003,N_9969,N_9909);
or UO_1004 (O_1004,N_9946,N_9988);
and UO_1005 (O_1005,N_9972,N_9977);
xnor UO_1006 (O_1006,N_9979,N_9999);
nor UO_1007 (O_1007,N_9966,N_9957);
and UO_1008 (O_1008,N_9993,N_9914);
and UO_1009 (O_1009,N_9988,N_9962);
or UO_1010 (O_1010,N_9986,N_9956);
and UO_1011 (O_1011,N_9923,N_9921);
xnor UO_1012 (O_1012,N_9948,N_9995);
and UO_1013 (O_1013,N_9960,N_9980);
or UO_1014 (O_1014,N_9996,N_9939);
and UO_1015 (O_1015,N_9900,N_9936);
and UO_1016 (O_1016,N_9975,N_9976);
and UO_1017 (O_1017,N_9915,N_9975);
nand UO_1018 (O_1018,N_9950,N_9974);
and UO_1019 (O_1019,N_9996,N_9956);
and UO_1020 (O_1020,N_9959,N_9967);
nand UO_1021 (O_1021,N_9925,N_9994);
or UO_1022 (O_1022,N_9993,N_9922);
and UO_1023 (O_1023,N_9902,N_9906);
nor UO_1024 (O_1024,N_9990,N_9971);
and UO_1025 (O_1025,N_9968,N_9983);
or UO_1026 (O_1026,N_9962,N_9997);
nand UO_1027 (O_1027,N_9922,N_9949);
or UO_1028 (O_1028,N_9904,N_9914);
and UO_1029 (O_1029,N_9975,N_9970);
nand UO_1030 (O_1030,N_9953,N_9910);
or UO_1031 (O_1031,N_9952,N_9923);
or UO_1032 (O_1032,N_9967,N_9928);
xor UO_1033 (O_1033,N_9954,N_9919);
nand UO_1034 (O_1034,N_9928,N_9940);
or UO_1035 (O_1035,N_9908,N_9903);
and UO_1036 (O_1036,N_9973,N_9934);
nand UO_1037 (O_1037,N_9971,N_9949);
or UO_1038 (O_1038,N_9968,N_9905);
nor UO_1039 (O_1039,N_9933,N_9915);
or UO_1040 (O_1040,N_9944,N_9981);
or UO_1041 (O_1041,N_9956,N_9946);
nand UO_1042 (O_1042,N_9971,N_9998);
nor UO_1043 (O_1043,N_9991,N_9984);
xor UO_1044 (O_1044,N_9969,N_9904);
or UO_1045 (O_1045,N_9930,N_9950);
nor UO_1046 (O_1046,N_9959,N_9983);
nor UO_1047 (O_1047,N_9994,N_9911);
nor UO_1048 (O_1048,N_9901,N_9948);
and UO_1049 (O_1049,N_9909,N_9978);
nor UO_1050 (O_1050,N_9999,N_9951);
and UO_1051 (O_1051,N_9934,N_9990);
or UO_1052 (O_1052,N_9981,N_9940);
nand UO_1053 (O_1053,N_9917,N_9991);
xor UO_1054 (O_1054,N_9921,N_9906);
and UO_1055 (O_1055,N_9967,N_9927);
or UO_1056 (O_1056,N_9916,N_9957);
nor UO_1057 (O_1057,N_9969,N_9922);
and UO_1058 (O_1058,N_9908,N_9955);
or UO_1059 (O_1059,N_9962,N_9993);
nand UO_1060 (O_1060,N_9943,N_9968);
and UO_1061 (O_1061,N_9943,N_9957);
or UO_1062 (O_1062,N_9959,N_9907);
nor UO_1063 (O_1063,N_9994,N_9985);
or UO_1064 (O_1064,N_9950,N_9945);
or UO_1065 (O_1065,N_9927,N_9900);
and UO_1066 (O_1066,N_9916,N_9939);
or UO_1067 (O_1067,N_9959,N_9934);
nor UO_1068 (O_1068,N_9910,N_9906);
and UO_1069 (O_1069,N_9952,N_9941);
and UO_1070 (O_1070,N_9966,N_9993);
nor UO_1071 (O_1071,N_9972,N_9966);
nand UO_1072 (O_1072,N_9977,N_9920);
nand UO_1073 (O_1073,N_9922,N_9943);
or UO_1074 (O_1074,N_9962,N_9922);
nand UO_1075 (O_1075,N_9965,N_9979);
nand UO_1076 (O_1076,N_9965,N_9974);
nor UO_1077 (O_1077,N_9957,N_9968);
nor UO_1078 (O_1078,N_9913,N_9900);
or UO_1079 (O_1079,N_9976,N_9974);
nor UO_1080 (O_1080,N_9952,N_9961);
nor UO_1081 (O_1081,N_9940,N_9954);
nor UO_1082 (O_1082,N_9986,N_9918);
nor UO_1083 (O_1083,N_9998,N_9908);
nand UO_1084 (O_1084,N_9979,N_9906);
nand UO_1085 (O_1085,N_9936,N_9964);
nand UO_1086 (O_1086,N_9970,N_9973);
and UO_1087 (O_1087,N_9987,N_9997);
nor UO_1088 (O_1088,N_9975,N_9927);
nor UO_1089 (O_1089,N_9968,N_9926);
and UO_1090 (O_1090,N_9904,N_9986);
nor UO_1091 (O_1091,N_9933,N_9997);
nor UO_1092 (O_1092,N_9920,N_9936);
or UO_1093 (O_1093,N_9971,N_9987);
and UO_1094 (O_1094,N_9999,N_9956);
xnor UO_1095 (O_1095,N_9933,N_9996);
or UO_1096 (O_1096,N_9902,N_9943);
nand UO_1097 (O_1097,N_9963,N_9991);
nor UO_1098 (O_1098,N_9987,N_9919);
nor UO_1099 (O_1099,N_9935,N_9972);
nor UO_1100 (O_1100,N_9903,N_9976);
nand UO_1101 (O_1101,N_9941,N_9974);
and UO_1102 (O_1102,N_9985,N_9942);
xor UO_1103 (O_1103,N_9934,N_9925);
and UO_1104 (O_1104,N_9929,N_9990);
nand UO_1105 (O_1105,N_9974,N_9931);
xor UO_1106 (O_1106,N_9922,N_9913);
nor UO_1107 (O_1107,N_9924,N_9914);
and UO_1108 (O_1108,N_9988,N_9921);
nand UO_1109 (O_1109,N_9977,N_9918);
nand UO_1110 (O_1110,N_9918,N_9947);
nor UO_1111 (O_1111,N_9980,N_9979);
and UO_1112 (O_1112,N_9960,N_9907);
nor UO_1113 (O_1113,N_9902,N_9950);
nand UO_1114 (O_1114,N_9909,N_9957);
nor UO_1115 (O_1115,N_9962,N_9973);
and UO_1116 (O_1116,N_9923,N_9955);
nand UO_1117 (O_1117,N_9987,N_9905);
or UO_1118 (O_1118,N_9933,N_9931);
and UO_1119 (O_1119,N_9964,N_9950);
nand UO_1120 (O_1120,N_9953,N_9927);
nor UO_1121 (O_1121,N_9999,N_9957);
nand UO_1122 (O_1122,N_9908,N_9957);
or UO_1123 (O_1123,N_9941,N_9991);
nor UO_1124 (O_1124,N_9949,N_9989);
nand UO_1125 (O_1125,N_9987,N_9910);
or UO_1126 (O_1126,N_9960,N_9986);
and UO_1127 (O_1127,N_9999,N_9945);
or UO_1128 (O_1128,N_9975,N_9934);
nor UO_1129 (O_1129,N_9909,N_9942);
xor UO_1130 (O_1130,N_9962,N_9940);
or UO_1131 (O_1131,N_9913,N_9995);
nor UO_1132 (O_1132,N_9983,N_9980);
xnor UO_1133 (O_1133,N_9905,N_9928);
and UO_1134 (O_1134,N_9903,N_9974);
nor UO_1135 (O_1135,N_9946,N_9962);
or UO_1136 (O_1136,N_9954,N_9900);
and UO_1137 (O_1137,N_9939,N_9929);
nand UO_1138 (O_1138,N_9936,N_9929);
nor UO_1139 (O_1139,N_9975,N_9999);
and UO_1140 (O_1140,N_9977,N_9944);
nor UO_1141 (O_1141,N_9959,N_9992);
and UO_1142 (O_1142,N_9966,N_9939);
nor UO_1143 (O_1143,N_9995,N_9943);
nand UO_1144 (O_1144,N_9903,N_9967);
nor UO_1145 (O_1145,N_9958,N_9982);
nor UO_1146 (O_1146,N_9953,N_9905);
and UO_1147 (O_1147,N_9961,N_9902);
nor UO_1148 (O_1148,N_9996,N_9944);
nand UO_1149 (O_1149,N_9962,N_9936);
and UO_1150 (O_1150,N_9903,N_9954);
nand UO_1151 (O_1151,N_9951,N_9983);
nor UO_1152 (O_1152,N_9979,N_9926);
or UO_1153 (O_1153,N_9918,N_9998);
or UO_1154 (O_1154,N_9907,N_9963);
and UO_1155 (O_1155,N_9972,N_9915);
nor UO_1156 (O_1156,N_9993,N_9924);
or UO_1157 (O_1157,N_9944,N_9978);
or UO_1158 (O_1158,N_9973,N_9982);
and UO_1159 (O_1159,N_9919,N_9926);
nor UO_1160 (O_1160,N_9951,N_9943);
or UO_1161 (O_1161,N_9949,N_9935);
or UO_1162 (O_1162,N_9936,N_9973);
nand UO_1163 (O_1163,N_9993,N_9977);
or UO_1164 (O_1164,N_9907,N_9933);
nor UO_1165 (O_1165,N_9939,N_9986);
or UO_1166 (O_1166,N_9913,N_9964);
and UO_1167 (O_1167,N_9963,N_9904);
nor UO_1168 (O_1168,N_9953,N_9906);
xnor UO_1169 (O_1169,N_9956,N_9967);
nand UO_1170 (O_1170,N_9915,N_9928);
and UO_1171 (O_1171,N_9943,N_9912);
nor UO_1172 (O_1172,N_9986,N_9905);
nand UO_1173 (O_1173,N_9960,N_9959);
or UO_1174 (O_1174,N_9940,N_9959);
nor UO_1175 (O_1175,N_9972,N_9923);
or UO_1176 (O_1176,N_9952,N_9981);
nand UO_1177 (O_1177,N_9920,N_9922);
or UO_1178 (O_1178,N_9911,N_9925);
or UO_1179 (O_1179,N_9992,N_9958);
and UO_1180 (O_1180,N_9935,N_9954);
and UO_1181 (O_1181,N_9912,N_9973);
xor UO_1182 (O_1182,N_9949,N_9914);
nand UO_1183 (O_1183,N_9924,N_9999);
and UO_1184 (O_1184,N_9989,N_9926);
and UO_1185 (O_1185,N_9938,N_9914);
nor UO_1186 (O_1186,N_9975,N_9961);
nand UO_1187 (O_1187,N_9905,N_9904);
or UO_1188 (O_1188,N_9958,N_9985);
nor UO_1189 (O_1189,N_9985,N_9968);
nand UO_1190 (O_1190,N_9905,N_9974);
and UO_1191 (O_1191,N_9958,N_9928);
and UO_1192 (O_1192,N_9948,N_9957);
nor UO_1193 (O_1193,N_9942,N_9907);
nor UO_1194 (O_1194,N_9906,N_9994);
and UO_1195 (O_1195,N_9974,N_9983);
and UO_1196 (O_1196,N_9949,N_9900);
and UO_1197 (O_1197,N_9986,N_9985);
and UO_1198 (O_1198,N_9946,N_9915);
nor UO_1199 (O_1199,N_9970,N_9971);
and UO_1200 (O_1200,N_9978,N_9939);
nor UO_1201 (O_1201,N_9951,N_9953);
nand UO_1202 (O_1202,N_9962,N_9913);
or UO_1203 (O_1203,N_9976,N_9973);
nor UO_1204 (O_1204,N_9934,N_9963);
nand UO_1205 (O_1205,N_9903,N_9929);
nand UO_1206 (O_1206,N_9919,N_9967);
nor UO_1207 (O_1207,N_9919,N_9952);
and UO_1208 (O_1208,N_9960,N_9969);
xor UO_1209 (O_1209,N_9993,N_9985);
nor UO_1210 (O_1210,N_9999,N_9946);
or UO_1211 (O_1211,N_9992,N_9917);
and UO_1212 (O_1212,N_9951,N_9904);
nor UO_1213 (O_1213,N_9916,N_9989);
and UO_1214 (O_1214,N_9914,N_9960);
nand UO_1215 (O_1215,N_9986,N_9934);
or UO_1216 (O_1216,N_9951,N_9946);
xnor UO_1217 (O_1217,N_9967,N_9921);
or UO_1218 (O_1218,N_9927,N_9916);
nor UO_1219 (O_1219,N_9911,N_9933);
and UO_1220 (O_1220,N_9943,N_9986);
nor UO_1221 (O_1221,N_9977,N_9992);
nand UO_1222 (O_1222,N_9921,N_9919);
and UO_1223 (O_1223,N_9901,N_9928);
nor UO_1224 (O_1224,N_9919,N_9911);
or UO_1225 (O_1225,N_9963,N_9948);
nand UO_1226 (O_1226,N_9912,N_9944);
nor UO_1227 (O_1227,N_9971,N_9915);
nor UO_1228 (O_1228,N_9992,N_9997);
and UO_1229 (O_1229,N_9918,N_9945);
or UO_1230 (O_1230,N_9991,N_9901);
and UO_1231 (O_1231,N_9910,N_9931);
and UO_1232 (O_1232,N_9910,N_9938);
nor UO_1233 (O_1233,N_9962,N_9926);
xnor UO_1234 (O_1234,N_9953,N_9917);
nor UO_1235 (O_1235,N_9936,N_9947);
nand UO_1236 (O_1236,N_9906,N_9973);
nor UO_1237 (O_1237,N_9977,N_9970);
or UO_1238 (O_1238,N_9968,N_9932);
nand UO_1239 (O_1239,N_9942,N_9960);
or UO_1240 (O_1240,N_9973,N_9942);
xor UO_1241 (O_1241,N_9997,N_9983);
nor UO_1242 (O_1242,N_9978,N_9972);
or UO_1243 (O_1243,N_9945,N_9984);
nor UO_1244 (O_1244,N_9935,N_9943);
or UO_1245 (O_1245,N_9987,N_9943);
or UO_1246 (O_1246,N_9938,N_9961);
xor UO_1247 (O_1247,N_9984,N_9911);
nand UO_1248 (O_1248,N_9923,N_9975);
nor UO_1249 (O_1249,N_9934,N_9944);
nand UO_1250 (O_1250,N_9994,N_9958);
nor UO_1251 (O_1251,N_9957,N_9984);
and UO_1252 (O_1252,N_9972,N_9959);
nand UO_1253 (O_1253,N_9985,N_9999);
and UO_1254 (O_1254,N_9983,N_9912);
or UO_1255 (O_1255,N_9979,N_9949);
nand UO_1256 (O_1256,N_9977,N_9908);
and UO_1257 (O_1257,N_9911,N_9977);
or UO_1258 (O_1258,N_9944,N_9976);
xor UO_1259 (O_1259,N_9962,N_9917);
and UO_1260 (O_1260,N_9916,N_9958);
nor UO_1261 (O_1261,N_9911,N_9944);
xor UO_1262 (O_1262,N_9993,N_9964);
nor UO_1263 (O_1263,N_9955,N_9975);
or UO_1264 (O_1264,N_9957,N_9924);
or UO_1265 (O_1265,N_9975,N_9906);
or UO_1266 (O_1266,N_9950,N_9978);
nor UO_1267 (O_1267,N_9918,N_9978);
or UO_1268 (O_1268,N_9934,N_9948);
nor UO_1269 (O_1269,N_9966,N_9906);
nand UO_1270 (O_1270,N_9932,N_9987);
and UO_1271 (O_1271,N_9921,N_9953);
and UO_1272 (O_1272,N_9988,N_9968);
nand UO_1273 (O_1273,N_9938,N_9997);
or UO_1274 (O_1274,N_9963,N_9966);
and UO_1275 (O_1275,N_9909,N_9940);
and UO_1276 (O_1276,N_9926,N_9993);
nor UO_1277 (O_1277,N_9955,N_9940);
nand UO_1278 (O_1278,N_9927,N_9901);
or UO_1279 (O_1279,N_9906,N_9935);
nor UO_1280 (O_1280,N_9993,N_9973);
nand UO_1281 (O_1281,N_9905,N_9930);
nor UO_1282 (O_1282,N_9951,N_9977);
or UO_1283 (O_1283,N_9953,N_9986);
nand UO_1284 (O_1284,N_9939,N_9908);
and UO_1285 (O_1285,N_9936,N_9952);
or UO_1286 (O_1286,N_9969,N_9937);
and UO_1287 (O_1287,N_9960,N_9954);
nand UO_1288 (O_1288,N_9993,N_9995);
nor UO_1289 (O_1289,N_9992,N_9901);
nand UO_1290 (O_1290,N_9947,N_9989);
or UO_1291 (O_1291,N_9981,N_9965);
nand UO_1292 (O_1292,N_9941,N_9913);
nand UO_1293 (O_1293,N_9941,N_9984);
nand UO_1294 (O_1294,N_9917,N_9945);
nor UO_1295 (O_1295,N_9977,N_9915);
nand UO_1296 (O_1296,N_9964,N_9912);
nand UO_1297 (O_1297,N_9990,N_9953);
or UO_1298 (O_1298,N_9920,N_9949);
nand UO_1299 (O_1299,N_9982,N_9931);
nor UO_1300 (O_1300,N_9941,N_9903);
and UO_1301 (O_1301,N_9925,N_9953);
or UO_1302 (O_1302,N_9939,N_9977);
and UO_1303 (O_1303,N_9930,N_9981);
and UO_1304 (O_1304,N_9966,N_9910);
and UO_1305 (O_1305,N_9958,N_9946);
and UO_1306 (O_1306,N_9942,N_9906);
or UO_1307 (O_1307,N_9931,N_9961);
nand UO_1308 (O_1308,N_9977,N_9914);
xor UO_1309 (O_1309,N_9977,N_9942);
and UO_1310 (O_1310,N_9999,N_9997);
or UO_1311 (O_1311,N_9911,N_9993);
nor UO_1312 (O_1312,N_9976,N_9957);
and UO_1313 (O_1313,N_9979,N_9943);
and UO_1314 (O_1314,N_9993,N_9931);
and UO_1315 (O_1315,N_9909,N_9993);
nand UO_1316 (O_1316,N_9973,N_9998);
xor UO_1317 (O_1317,N_9902,N_9912);
or UO_1318 (O_1318,N_9907,N_9920);
and UO_1319 (O_1319,N_9975,N_9977);
or UO_1320 (O_1320,N_9968,N_9977);
and UO_1321 (O_1321,N_9957,N_9921);
or UO_1322 (O_1322,N_9970,N_9981);
and UO_1323 (O_1323,N_9912,N_9911);
nor UO_1324 (O_1324,N_9932,N_9900);
nor UO_1325 (O_1325,N_9968,N_9955);
nand UO_1326 (O_1326,N_9904,N_9990);
nor UO_1327 (O_1327,N_9908,N_9912);
and UO_1328 (O_1328,N_9920,N_9913);
nor UO_1329 (O_1329,N_9947,N_9966);
and UO_1330 (O_1330,N_9948,N_9970);
nor UO_1331 (O_1331,N_9915,N_9945);
or UO_1332 (O_1332,N_9949,N_9955);
or UO_1333 (O_1333,N_9929,N_9912);
and UO_1334 (O_1334,N_9969,N_9906);
nand UO_1335 (O_1335,N_9983,N_9932);
or UO_1336 (O_1336,N_9900,N_9912);
or UO_1337 (O_1337,N_9937,N_9925);
and UO_1338 (O_1338,N_9982,N_9945);
and UO_1339 (O_1339,N_9930,N_9903);
or UO_1340 (O_1340,N_9971,N_9956);
and UO_1341 (O_1341,N_9950,N_9921);
or UO_1342 (O_1342,N_9969,N_9919);
and UO_1343 (O_1343,N_9945,N_9954);
nand UO_1344 (O_1344,N_9994,N_9991);
or UO_1345 (O_1345,N_9933,N_9995);
nor UO_1346 (O_1346,N_9987,N_9963);
or UO_1347 (O_1347,N_9979,N_9923);
or UO_1348 (O_1348,N_9953,N_9955);
nor UO_1349 (O_1349,N_9935,N_9970);
nor UO_1350 (O_1350,N_9999,N_9919);
or UO_1351 (O_1351,N_9934,N_9994);
nor UO_1352 (O_1352,N_9936,N_9991);
and UO_1353 (O_1353,N_9997,N_9976);
or UO_1354 (O_1354,N_9920,N_9993);
nor UO_1355 (O_1355,N_9975,N_9919);
nor UO_1356 (O_1356,N_9902,N_9962);
nand UO_1357 (O_1357,N_9965,N_9946);
and UO_1358 (O_1358,N_9913,N_9919);
nor UO_1359 (O_1359,N_9956,N_9928);
or UO_1360 (O_1360,N_9943,N_9939);
xnor UO_1361 (O_1361,N_9956,N_9953);
xor UO_1362 (O_1362,N_9955,N_9916);
nand UO_1363 (O_1363,N_9906,N_9977);
nand UO_1364 (O_1364,N_9987,N_9961);
nand UO_1365 (O_1365,N_9923,N_9942);
and UO_1366 (O_1366,N_9956,N_9998);
nand UO_1367 (O_1367,N_9966,N_9989);
nor UO_1368 (O_1368,N_9902,N_9953);
nor UO_1369 (O_1369,N_9926,N_9939);
or UO_1370 (O_1370,N_9984,N_9998);
and UO_1371 (O_1371,N_9905,N_9944);
and UO_1372 (O_1372,N_9959,N_9914);
or UO_1373 (O_1373,N_9900,N_9931);
or UO_1374 (O_1374,N_9976,N_9964);
or UO_1375 (O_1375,N_9971,N_9988);
xnor UO_1376 (O_1376,N_9983,N_9956);
or UO_1377 (O_1377,N_9989,N_9942);
nor UO_1378 (O_1378,N_9971,N_9901);
nand UO_1379 (O_1379,N_9961,N_9950);
xnor UO_1380 (O_1380,N_9969,N_9902);
nor UO_1381 (O_1381,N_9977,N_9967);
or UO_1382 (O_1382,N_9975,N_9945);
and UO_1383 (O_1383,N_9918,N_9955);
nor UO_1384 (O_1384,N_9977,N_9917);
and UO_1385 (O_1385,N_9924,N_9979);
or UO_1386 (O_1386,N_9938,N_9964);
nand UO_1387 (O_1387,N_9987,N_9965);
and UO_1388 (O_1388,N_9985,N_9945);
nand UO_1389 (O_1389,N_9946,N_9973);
nand UO_1390 (O_1390,N_9907,N_9928);
and UO_1391 (O_1391,N_9927,N_9952);
or UO_1392 (O_1392,N_9978,N_9948);
or UO_1393 (O_1393,N_9928,N_9934);
nor UO_1394 (O_1394,N_9967,N_9939);
nand UO_1395 (O_1395,N_9987,N_9960);
nor UO_1396 (O_1396,N_9994,N_9986);
nand UO_1397 (O_1397,N_9949,N_9954);
nand UO_1398 (O_1398,N_9997,N_9931);
nand UO_1399 (O_1399,N_9935,N_9926);
or UO_1400 (O_1400,N_9995,N_9906);
and UO_1401 (O_1401,N_9971,N_9921);
or UO_1402 (O_1402,N_9947,N_9919);
nor UO_1403 (O_1403,N_9901,N_9953);
nor UO_1404 (O_1404,N_9933,N_9983);
or UO_1405 (O_1405,N_9982,N_9942);
and UO_1406 (O_1406,N_9918,N_9994);
nor UO_1407 (O_1407,N_9966,N_9933);
nand UO_1408 (O_1408,N_9946,N_9918);
and UO_1409 (O_1409,N_9962,N_9933);
or UO_1410 (O_1410,N_9974,N_9978);
and UO_1411 (O_1411,N_9935,N_9917);
or UO_1412 (O_1412,N_9948,N_9969);
and UO_1413 (O_1413,N_9934,N_9929);
and UO_1414 (O_1414,N_9961,N_9949);
nor UO_1415 (O_1415,N_9915,N_9994);
or UO_1416 (O_1416,N_9946,N_9935);
nand UO_1417 (O_1417,N_9919,N_9959);
and UO_1418 (O_1418,N_9949,N_9907);
or UO_1419 (O_1419,N_9964,N_9902);
and UO_1420 (O_1420,N_9919,N_9939);
and UO_1421 (O_1421,N_9956,N_9980);
nor UO_1422 (O_1422,N_9905,N_9921);
or UO_1423 (O_1423,N_9940,N_9935);
nand UO_1424 (O_1424,N_9959,N_9971);
or UO_1425 (O_1425,N_9930,N_9934);
or UO_1426 (O_1426,N_9967,N_9960);
nor UO_1427 (O_1427,N_9992,N_9924);
nor UO_1428 (O_1428,N_9917,N_9944);
and UO_1429 (O_1429,N_9900,N_9989);
nor UO_1430 (O_1430,N_9945,N_9947);
or UO_1431 (O_1431,N_9916,N_9962);
nor UO_1432 (O_1432,N_9947,N_9996);
and UO_1433 (O_1433,N_9991,N_9943);
nor UO_1434 (O_1434,N_9953,N_9936);
nand UO_1435 (O_1435,N_9936,N_9928);
or UO_1436 (O_1436,N_9941,N_9950);
nor UO_1437 (O_1437,N_9991,N_9959);
nor UO_1438 (O_1438,N_9982,N_9919);
or UO_1439 (O_1439,N_9905,N_9935);
nand UO_1440 (O_1440,N_9906,N_9957);
nor UO_1441 (O_1441,N_9972,N_9968);
or UO_1442 (O_1442,N_9918,N_9984);
or UO_1443 (O_1443,N_9992,N_9965);
or UO_1444 (O_1444,N_9953,N_9900);
nor UO_1445 (O_1445,N_9945,N_9987);
nand UO_1446 (O_1446,N_9934,N_9945);
nor UO_1447 (O_1447,N_9930,N_9957);
nand UO_1448 (O_1448,N_9967,N_9993);
or UO_1449 (O_1449,N_9964,N_9979);
nor UO_1450 (O_1450,N_9931,N_9924);
nand UO_1451 (O_1451,N_9987,N_9913);
nor UO_1452 (O_1452,N_9978,N_9971);
and UO_1453 (O_1453,N_9987,N_9920);
nand UO_1454 (O_1454,N_9942,N_9953);
nor UO_1455 (O_1455,N_9983,N_9952);
nand UO_1456 (O_1456,N_9901,N_9925);
nand UO_1457 (O_1457,N_9989,N_9919);
or UO_1458 (O_1458,N_9953,N_9919);
and UO_1459 (O_1459,N_9940,N_9990);
nor UO_1460 (O_1460,N_9999,N_9921);
nor UO_1461 (O_1461,N_9965,N_9933);
or UO_1462 (O_1462,N_9976,N_9952);
nor UO_1463 (O_1463,N_9925,N_9963);
nand UO_1464 (O_1464,N_9960,N_9952);
nor UO_1465 (O_1465,N_9908,N_9921);
and UO_1466 (O_1466,N_9916,N_9981);
and UO_1467 (O_1467,N_9903,N_9987);
nand UO_1468 (O_1468,N_9974,N_9930);
or UO_1469 (O_1469,N_9970,N_9934);
xor UO_1470 (O_1470,N_9916,N_9949);
or UO_1471 (O_1471,N_9916,N_9978);
nand UO_1472 (O_1472,N_9935,N_9967);
nand UO_1473 (O_1473,N_9910,N_9920);
nand UO_1474 (O_1474,N_9977,N_9947);
and UO_1475 (O_1475,N_9933,N_9943);
nand UO_1476 (O_1476,N_9959,N_9982);
nand UO_1477 (O_1477,N_9960,N_9934);
nand UO_1478 (O_1478,N_9909,N_9933);
nand UO_1479 (O_1479,N_9918,N_9993);
nand UO_1480 (O_1480,N_9921,N_9969);
nor UO_1481 (O_1481,N_9933,N_9904);
and UO_1482 (O_1482,N_9928,N_9955);
nor UO_1483 (O_1483,N_9935,N_9998);
nor UO_1484 (O_1484,N_9948,N_9992);
nor UO_1485 (O_1485,N_9950,N_9968);
and UO_1486 (O_1486,N_9929,N_9948);
nor UO_1487 (O_1487,N_9988,N_9949);
nor UO_1488 (O_1488,N_9998,N_9946);
nor UO_1489 (O_1489,N_9972,N_9934);
nand UO_1490 (O_1490,N_9933,N_9901);
nand UO_1491 (O_1491,N_9907,N_9932);
nor UO_1492 (O_1492,N_9906,N_9965);
nand UO_1493 (O_1493,N_9971,N_9920);
nor UO_1494 (O_1494,N_9958,N_9943);
nor UO_1495 (O_1495,N_9994,N_9950);
nor UO_1496 (O_1496,N_9918,N_9962);
nand UO_1497 (O_1497,N_9935,N_9933);
nand UO_1498 (O_1498,N_9931,N_9971);
or UO_1499 (O_1499,N_9998,N_9906);
endmodule