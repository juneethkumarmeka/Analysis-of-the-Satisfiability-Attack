module basic_500_3000_500_6_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_448,In_107);
nand U1 (N_1,In_258,In_296);
or U2 (N_2,In_413,In_10);
or U3 (N_3,In_397,In_377);
nor U4 (N_4,In_109,In_101);
and U5 (N_5,In_52,In_419);
or U6 (N_6,In_149,In_429);
nor U7 (N_7,In_382,In_68);
nor U8 (N_8,In_75,In_61);
or U9 (N_9,In_73,In_454);
or U10 (N_10,In_456,In_79);
nor U11 (N_11,In_476,In_472);
nand U12 (N_12,In_358,In_257);
nor U13 (N_13,In_317,In_351);
xnor U14 (N_14,In_243,In_301);
xnor U15 (N_15,In_404,In_49);
xnor U16 (N_16,In_411,In_232);
or U17 (N_17,In_150,In_279);
and U18 (N_18,In_455,In_241);
xor U19 (N_19,In_447,In_340);
nand U20 (N_20,In_58,In_48);
or U21 (N_21,In_294,In_291);
nand U22 (N_22,In_217,In_99);
xnor U23 (N_23,In_238,In_147);
nand U24 (N_24,In_25,In_188);
nor U25 (N_25,In_189,In_348);
xor U26 (N_26,In_30,In_225);
and U27 (N_27,In_298,In_209);
or U28 (N_28,In_441,In_178);
and U29 (N_29,In_249,In_487);
or U30 (N_30,In_40,In_56);
or U31 (N_31,In_313,In_174);
xor U32 (N_32,In_103,In_67);
nor U33 (N_33,In_104,In_426);
or U34 (N_34,In_204,In_435);
xnor U35 (N_35,In_443,In_256);
or U36 (N_36,In_371,In_323);
or U37 (N_37,In_490,In_2);
nand U38 (N_38,In_423,In_100);
xnor U39 (N_39,In_254,In_231);
or U40 (N_40,In_72,In_37);
nand U41 (N_41,In_60,In_195);
and U42 (N_42,In_197,In_444);
xnor U43 (N_43,In_336,In_108);
and U44 (N_44,In_495,In_213);
nor U45 (N_45,In_437,In_163);
or U46 (N_46,In_143,In_171);
or U47 (N_47,In_221,In_338);
and U48 (N_48,In_57,In_310);
xor U49 (N_49,In_8,In_239);
nand U50 (N_50,In_192,In_123);
nor U51 (N_51,In_216,In_71);
nor U52 (N_52,In_461,In_224);
nand U53 (N_53,In_450,In_115);
xnor U54 (N_54,In_141,In_26);
nor U55 (N_55,In_299,In_18);
nand U56 (N_56,In_428,In_119);
nand U57 (N_57,In_96,In_285);
nand U58 (N_58,In_401,In_168);
nand U59 (N_59,In_392,In_384);
or U60 (N_60,In_233,In_311);
nand U61 (N_61,In_356,In_278);
nand U62 (N_62,In_226,In_474);
xnor U63 (N_63,In_480,In_135);
nand U64 (N_64,In_245,In_110);
xnor U65 (N_65,In_342,In_489);
xor U66 (N_66,In_271,In_334);
xnor U67 (N_67,In_167,In_330);
xor U68 (N_68,In_445,In_191);
nand U69 (N_69,In_128,In_247);
nor U70 (N_70,In_302,In_473);
nor U71 (N_71,In_223,In_66);
nand U72 (N_72,In_148,In_399);
nand U73 (N_73,In_389,In_208);
xor U74 (N_74,In_469,In_388);
and U75 (N_75,In_50,In_46);
xnor U76 (N_76,In_492,In_42);
and U77 (N_77,In_54,In_372);
and U78 (N_78,In_357,In_59);
nor U79 (N_79,In_344,In_74);
nand U80 (N_80,In_433,In_207);
or U81 (N_81,In_360,In_264);
nand U82 (N_82,In_451,In_151);
xnor U83 (N_83,In_331,In_470);
and U84 (N_84,In_333,In_95);
nor U85 (N_85,In_303,In_493);
nand U86 (N_86,In_130,In_464);
nand U87 (N_87,In_438,In_272);
nor U88 (N_88,In_280,In_211);
xnor U89 (N_89,In_332,In_77);
nor U90 (N_90,In_196,In_337);
and U91 (N_91,In_418,In_183);
xnor U92 (N_92,In_321,In_111);
nand U93 (N_93,In_477,In_308);
and U94 (N_94,In_312,In_482);
and U95 (N_95,In_12,In_421);
nor U96 (N_96,In_176,In_431);
nand U97 (N_97,In_146,In_459);
or U98 (N_98,In_97,In_289);
and U99 (N_99,In_362,In_94);
or U100 (N_100,In_432,In_1);
or U101 (N_101,In_341,In_133);
xnor U102 (N_102,In_414,In_80);
nor U103 (N_103,In_138,In_152);
and U104 (N_104,In_304,In_307);
xor U105 (N_105,In_394,In_449);
and U106 (N_106,In_186,In_105);
nand U107 (N_107,In_420,In_267);
xnor U108 (N_108,In_7,In_205);
nor U109 (N_109,In_410,In_374);
nand U110 (N_110,In_265,In_380);
xor U111 (N_111,In_165,In_121);
xnor U112 (N_112,In_467,In_203);
and U113 (N_113,In_38,In_9);
and U114 (N_114,In_499,In_282);
nand U115 (N_115,In_64,In_277);
xor U116 (N_116,In_355,In_306);
nor U117 (N_117,In_354,In_236);
nand U118 (N_118,In_252,In_488);
or U119 (N_119,In_270,In_43);
nor U120 (N_120,In_403,In_453);
or U121 (N_121,In_23,In_92);
and U122 (N_122,In_180,In_63);
and U123 (N_123,In_400,In_475);
nand U124 (N_124,In_367,In_398);
or U125 (N_125,In_136,In_113);
nor U126 (N_126,In_266,In_391);
and U127 (N_127,In_320,In_349);
and U128 (N_128,In_200,In_295);
xor U129 (N_129,In_407,In_98);
nand U130 (N_130,In_466,In_190);
nand U131 (N_131,In_248,In_406);
and U132 (N_132,In_84,In_222);
nand U133 (N_133,In_44,In_315);
and U134 (N_134,In_122,In_0);
xnor U135 (N_135,In_288,In_234);
or U136 (N_136,In_415,In_118);
nand U137 (N_137,In_198,In_202);
nand U138 (N_138,In_373,In_327);
and U139 (N_139,In_405,In_242);
and U140 (N_140,In_172,In_300);
nand U141 (N_141,In_283,In_240);
or U142 (N_142,In_370,In_235);
nor U143 (N_143,In_286,In_255);
xnor U144 (N_144,In_462,In_153);
and U145 (N_145,In_326,In_90);
or U146 (N_146,In_309,In_131);
xor U147 (N_147,In_383,In_325);
or U148 (N_148,In_393,In_352);
nor U149 (N_149,In_164,In_206);
nor U150 (N_150,In_27,In_457);
and U151 (N_151,In_155,In_120);
or U152 (N_152,In_182,In_83);
or U153 (N_153,In_62,In_32);
nand U154 (N_154,In_78,In_35);
or U155 (N_155,In_379,In_436);
or U156 (N_156,In_70,In_250);
nand U157 (N_157,In_484,In_175);
or U158 (N_158,In_368,In_424);
nand U159 (N_159,In_422,In_485);
nor U160 (N_160,In_13,In_408);
and U161 (N_161,In_276,In_114);
or U162 (N_162,In_169,In_160);
xor U163 (N_163,In_434,In_194);
xor U164 (N_164,In_6,In_439);
nand U165 (N_165,In_142,In_416);
and U166 (N_166,In_491,In_14);
or U167 (N_167,In_268,In_220);
nor U168 (N_168,In_45,In_324);
xnor U169 (N_169,In_55,In_361);
xnor U170 (N_170,In_259,In_31);
and U171 (N_171,In_88,In_230);
and U172 (N_172,In_47,In_396);
xor U173 (N_173,In_177,In_126);
nor U174 (N_174,In_134,In_284);
and U175 (N_175,In_184,In_446);
xor U176 (N_176,In_215,In_65);
and U177 (N_177,In_157,In_21);
and U178 (N_178,In_11,In_82);
and U179 (N_179,In_161,In_390);
xor U180 (N_180,In_91,In_166);
nand U181 (N_181,In_181,In_350);
or U182 (N_182,In_427,In_497);
nand U183 (N_183,In_251,In_29);
nand U184 (N_184,In_17,In_417);
nor U185 (N_185,In_3,In_385);
nand U186 (N_186,In_51,In_106);
or U187 (N_187,In_20,In_339);
xnor U188 (N_188,In_218,In_36);
and U189 (N_189,In_112,In_481);
nand U190 (N_190,In_137,In_158);
nor U191 (N_191,In_375,In_93);
or U192 (N_192,In_261,In_102);
xnor U193 (N_193,In_366,In_345);
nand U194 (N_194,In_227,In_19);
nand U195 (N_195,In_395,In_262);
nand U196 (N_196,In_293,In_124);
and U197 (N_197,In_129,In_33);
nand U198 (N_198,In_24,In_214);
nor U199 (N_199,In_201,In_69);
nand U200 (N_200,In_144,In_478);
nor U201 (N_201,In_479,In_76);
and U202 (N_202,In_292,In_170);
nand U203 (N_203,In_41,In_440);
xor U204 (N_204,In_316,In_297);
xor U205 (N_205,In_179,In_364);
or U206 (N_206,In_486,In_305);
xor U207 (N_207,In_228,In_173);
nand U208 (N_208,In_263,In_162);
xor U209 (N_209,In_132,In_229);
nor U210 (N_210,In_287,In_193);
and U211 (N_211,In_329,In_402);
nor U212 (N_212,In_156,In_89);
nand U213 (N_213,In_353,In_494);
or U214 (N_214,In_81,In_381);
nand U215 (N_215,In_127,In_86);
nor U216 (N_216,In_154,In_452);
or U217 (N_217,In_187,In_28);
or U218 (N_218,In_15,In_318);
xor U219 (N_219,In_365,In_53);
nor U220 (N_220,In_319,In_237);
nor U221 (N_221,In_369,In_199);
nor U222 (N_222,In_253,In_260);
xnor U223 (N_223,In_498,In_16);
and U224 (N_224,In_463,In_347);
nand U225 (N_225,In_386,In_281);
nor U226 (N_226,In_387,In_139);
and U227 (N_227,In_269,In_471);
xor U228 (N_228,In_39,In_496);
nand U229 (N_229,In_145,In_376);
or U230 (N_230,In_430,In_468);
nor U231 (N_231,In_378,In_210);
xor U232 (N_232,In_22,In_159);
or U233 (N_233,In_290,In_85);
nand U234 (N_234,In_246,In_185);
nand U235 (N_235,In_273,In_465);
and U236 (N_236,In_363,In_328);
and U237 (N_237,In_274,In_412);
nand U238 (N_238,In_335,In_117);
nor U239 (N_239,In_140,In_346);
nor U240 (N_240,In_460,In_425);
nand U241 (N_241,In_409,In_4);
and U242 (N_242,In_275,In_219);
and U243 (N_243,In_5,In_212);
nand U244 (N_244,In_322,In_483);
or U245 (N_245,In_244,In_34);
xnor U246 (N_246,In_343,In_442);
and U247 (N_247,In_314,In_87);
nand U248 (N_248,In_458,In_359);
nor U249 (N_249,In_125,In_116);
xor U250 (N_250,In_295,In_440);
or U251 (N_251,In_299,In_241);
nor U252 (N_252,In_308,In_370);
nand U253 (N_253,In_202,In_347);
xor U254 (N_254,In_366,In_123);
xor U255 (N_255,In_381,In_405);
nor U256 (N_256,In_127,In_375);
or U257 (N_257,In_86,In_77);
and U258 (N_258,In_20,In_229);
nor U259 (N_259,In_182,In_392);
nand U260 (N_260,In_221,In_106);
xor U261 (N_261,In_429,In_252);
nand U262 (N_262,In_119,In_459);
or U263 (N_263,In_265,In_438);
or U264 (N_264,In_72,In_300);
or U265 (N_265,In_474,In_171);
xnor U266 (N_266,In_91,In_416);
and U267 (N_267,In_452,In_87);
and U268 (N_268,In_334,In_287);
xor U269 (N_269,In_308,In_79);
nand U270 (N_270,In_113,In_261);
xnor U271 (N_271,In_286,In_414);
or U272 (N_272,In_332,In_140);
nor U273 (N_273,In_4,In_482);
or U274 (N_274,In_281,In_265);
nor U275 (N_275,In_83,In_345);
xor U276 (N_276,In_39,In_114);
nand U277 (N_277,In_203,In_309);
nor U278 (N_278,In_294,In_177);
xnor U279 (N_279,In_181,In_90);
nor U280 (N_280,In_365,In_251);
nor U281 (N_281,In_214,In_315);
xor U282 (N_282,In_196,In_352);
and U283 (N_283,In_68,In_466);
nor U284 (N_284,In_421,In_9);
nor U285 (N_285,In_300,In_42);
nand U286 (N_286,In_358,In_381);
xor U287 (N_287,In_151,In_75);
xnor U288 (N_288,In_221,In_303);
nor U289 (N_289,In_9,In_124);
xnor U290 (N_290,In_431,In_146);
xor U291 (N_291,In_205,In_162);
xnor U292 (N_292,In_228,In_211);
and U293 (N_293,In_303,In_349);
and U294 (N_294,In_82,In_51);
or U295 (N_295,In_137,In_196);
and U296 (N_296,In_83,In_327);
and U297 (N_297,In_94,In_192);
xnor U298 (N_298,In_291,In_18);
nor U299 (N_299,In_399,In_152);
and U300 (N_300,In_28,In_424);
and U301 (N_301,In_114,In_440);
xnor U302 (N_302,In_334,In_357);
and U303 (N_303,In_300,In_399);
nand U304 (N_304,In_473,In_193);
and U305 (N_305,In_373,In_124);
or U306 (N_306,In_428,In_142);
and U307 (N_307,In_382,In_421);
and U308 (N_308,In_45,In_106);
and U309 (N_309,In_60,In_89);
xor U310 (N_310,In_212,In_229);
and U311 (N_311,In_484,In_226);
nor U312 (N_312,In_286,In_38);
xor U313 (N_313,In_237,In_322);
nand U314 (N_314,In_414,In_281);
nand U315 (N_315,In_341,In_304);
nor U316 (N_316,In_68,In_387);
xor U317 (N_317,In_275,In_5);
or U318 (N_318,In_212,In_357);
xnor U319 (N_319,In_497,In_436);
or U320 (N_320,In_320,In_177);
xor U321 (N_321,In_420,In_304);
nand U322 (N_322,In_59,In_95);
xor U323 (N_323,In_16,In_168);
or U324 (N_324,In_326,In_191);
nor U325 (N_325,In_186,In_194);
and U326 (N_326,In_445,In_293);
nand U327 (N_327,In_6,In_440);
and U328 (N_328,In_466,In_442);
and U329 (N_329,In_351,In_329);
nor U330 (N_330,In_166,In_137);
xor U331 (N_331,In_442,In_244);
or U332 (N_332,In_107,In_242);
xnor U333 (N_333,In_155,In_429);
xnor U334 (N_334,In_275,In_257);
and U335 (N_335,In_417,In_3);
nand U336 (N_336,In_30,In_391);
nor U337 (N_337,In_364,In_308);
xnor U338 (N_338,In_401,In_63);
nand U339 (N_339,In_117,In_448);
nor U340 (N_340,In_110,In_23);
and U341 (N_341,In_26,In_74);
nand U342 (N_342,In_148,In_305);
and U343 (N_343,In_224,In_440);
xnor U344 (N_344,In_149,In_277);
nor U345 (N_345,In_472,In_15);
and U346 (N_346,In_98,In_270);
and U347 (N_347,In_498,In_131);
nor U348 (N_348,In_49,In_326);
nor U349 (N_349,In_154,In_82);
and U350 (N_350,In_425,In_459);
nor U351 (N_351,In_200,In_348);
xor U352 (N_352,In_279,In_329);
and U353 (N_353,In_431,In_67);
xor U354 (N_354,In_199,In_284);
or U355 (N_355,In_46,In_234);
xnor U356 (N_356,In_216,In_214);
xor U357 (N_357,In_459,In_263);
xor U358 (N_358,In_146,In_317);
nor U359 (N_359,In_296,In_398);
or U360 (N_360,In_151,In_349);
or U361 (N_361,In_143,In_413);
nor U362 (N_362,In_367,In_465);
and U363 (N_363,In_70,In_89);
nand U364 (N_364,In_250,In_194);
nand U365 (N_365,In_45,In_72);
and U366 (N_366,In_367,In_387);
xnor U367 (N_367,In_199,In_20);
nand U368 (N_368,In_57,In_428);
nand U369 (N_369,In_414,In_8);
xor U370 (N_370,In_365,In_103);
xor U371 (N_371,In_348,In_195);
nand U372 (N_372,In_445,In_449);
or U373 (N_373,In_330,In_165);
xor U374 (N_374,In_315,In_472);
xor U375 (N_375,In_166,In_85);
and U376 (N_376,In_490,In_69);
and U377 (N_377,In_127,In_111);
xor U378 (N_378,In_97,In_158);
nand U379 (N_379,In_445,In_342);
or U380 (N_380,In_369,In_415);
xnor U381 (N_381,In_438,In_402);
or U382 (N_382,In_285,In_178);
xor U383 (N_383,In_4,In_394);
nor U384 (N_384,In_10,In_148);
nor U385 (N_385,In_96,In_104);
xor U386 (N_386,In_193,In_151);
and U387 (N_387,In_387,In_328);
nor U388 (N_388,In_359,In_71);
or U389 (N_389,In_259,In_226);
nor U390 (N_390,In_43,In_126);
or U391 (N_391,In_477,In_94);
and U392 (N_392,In_117,In_412);
nand U393 (N_393,In_132,In_136);
nand U394 (N_394,In_450,In_28);
or U395 (N_395,In_66,In_487);
or U396 (N_396,In_330,In_393);
and U397 (N_397,In_347,In_393);
nand U398 (N_398,In_19,In_294);
nor U399 (N_399,In_48,In_266);
and U400 (N_400,In_21,In_87);
nor U401 (N_401,In_146,In_182);
nor U402 (N_402,In_54,In_268);
nor U403 (N_403,In_363,In_280);
and U404 (N_404,In_67,In_157);
nand U405 (N_405,In_8,In_154);
xor U406 (N_406,In_176,In_190);
nand U407 (N_407,In_226,In_456);
xor U408 (N_408,In_94,In_352);
nor U409 (N_409,In_20,In_127);
xnor U410 (N_410,In_425,In_490);
nor U411 (N_411,In_442,In_13);
xor U412 (N_412,In_231,In_171);
xnor U413 (N_413,In_304,In_17);
xnor U414 (N_414,In_338,In_325);
xor U415 (N_415,In_48,In_350);
nand U416 (N_416,In_195,In_409);
and U417 (N_417,In_271,In_198);
nor U418 (N_418,In_349,In_128);
or U419 (N_419,In_80,In_377);
nand U420 (N_420,In_399,In_262);
nand U421 (N_421,In_232,In_480);
nand U422 (N_422,In_221,In_318);
and U423 (N_423,In_210,In_280);
xnor U424 (N_424,In_305,In_244);
nand U425 (N_425,In_412,In_232);
and U426 (N_426,In_21,In_390);
nor U427 (N_427,In_209,In_406);
or U428 (N_428,In_395,In_479);
xor U429 (N_429,In_448,In_275);
or U430 (N_430,In_213,In_179);
xor U431 (N_431,In_437,In_149);
nand U432 (N_432,In_459,In_393);
nand U433 (N_433,In_49,In_485);
nand U434 (N_434,In_114,In_4);
xor U435 (N_435,In_48,In_394);
xnor U436 (N_436,In_78,In_460);
nand U437 (N_437,In_180,In_121);
xnor U438 (N_438,In_98,In_57);
nand U439 (N_439,In_181,In_446);
or U440 (N_440,In_105,In_5);
xnor U441 (N_441,In_138,In_61);
nor U442 (N_442,In_9,In_138);
nand U443 (N_443,In_154,In_319);
nor U444 (N_444,In_405,In_488);
xnor U445 (N_445,In_424,In_146);
xnor U446 (N_446,In_202,In_136);
nor U447 (N_447,In_477,In_485);
xnor U448 (N_448,In_440,In_352);
or U449 (N_449,In_217,In_215);
xnor U450 (N_450,In_363,In_128);
and U451 (N_451,In_158,In_200);
or U452 (N_452,In_67,In_132);
or U453 (N_453,In_425,In_410);
xnor U454 (N_454,In_70,In_305);
nor U455 (N_455,In_478,In_228);
xor U456 (N_456,In_17,In_234);
or U457 (N_457,In_280,In_191);
nand U458 (N_458,In_355,In_15);
nand U459 (N_459,In_397,In_160);
nand U460 (N_460,In_400,In_18);
nor U461 (N_461,In_151,In_153);
and U462 (N_462,In_130,In_123);
xnor U463 (N_463,In_43,In_7);
or U464 (N_464,In_40,In_139);
nor U465 (N_465,In_278,In_268);
and U466 (N_466,In_351,In_188);
nor U467 (N_467,In_308,In_490);
xnor U468 (N_468,In_101,In_434);
or U469 (N_469,In_268,In_485);
or U470 (N_470,In_166,In_156);
or U471 (N_471,In_139,In_110);
xnor U472 (N_472,In_174,In_260);
xnor U473 (N_473,In_273,In_208);
or U474 (N_474,In_8,In_268);
or U475 (N_475,In_221,In_372);
nor U476 (N_476,In_70,In_409);
or U477 (N_477,In_464,In_101);
nor U478 (N_478,In_385,In_298);
or U479 (N_479,In_446,In_470);
and U480 (N_480,In_266,In_109);
nand U481 (N_481,In_405,In_72);
or U482 (N_482,In_161,In_29);
nor U483 (N_483,In_351,In_59);
nor U484 (N_484,In_281,In_399);
nand U485 (N_485,In_486,In_292);
and U486 (N_486,In_55,In_400);
nand U487 (N_487,In_418,In_162);
nand U488 (N_488,In_130,In_20);
nor U489 (N_489,In_283,In_493);
xnor U490 (N_490,In_405,In_457);
nor U491 (N_491,In_248,In_167);
xnor U492 (N_492,In_324,In_7);
xnor U493 (N_493,In_203,In_422);
and U494 (N_494,In_211,In_25);
and U495 (N_495,In_211,In_187);
xor U496 (N_496,In_36,In_154);
xnor U497 (N_497,In_465,In_287);
nand U498 (N_498,In_413,In_363);
nand U499 (N_499,In_340,In_187);
nor U500 (N_500,N_173,N_2);
xor U501 (N_501,N_317,N_129);
and U502 (N_502,N_253,N_373);
xnor U503 (N_503,N_438,N_213);
nor U504 (N_504,N_46,N_483);
xor U505 (N_505,N_305,N_144);
nand U506 (N_506,N_261,N_219);
xnor U507 (N_507,N_248,N_328);
xor U508 (N_508,N_223,N_238);
nor U509 (N_509,N_64,N_444);
xnor U510 (N_510,N_11,N_419);
and U511 (N_511,N_320,N_142);
nand U512 (N_512,N_287,N_364);
or U513 (N_513,N_474,N_288);
nand U514 (N_514,N_323,N_24);
nor U515 (N_515,N_35,N_94);
or U516 (N_516,N_293,N_43);
or U517 (N_517,N_299,N_154);
xnor U518 (N_518,N_376,N_63);
and U519 (N_519,N_339,N_255);
xor U520 (N_520,N_335,N_347);
and U521 (N_521,N_8,N_125);
xnor U522 (N_522,N_297,N_420);
and U523 (N_523,N_31,N_498);
and U524 (N_524,N_188,N_414);
or U525 (N_525,N_389,N_89);
and U526 (N_526,N_4,N_0);
nor U527 (N_527,N_300,N_39);
or U528 (N_528,N_367,N_148);
or U529 (N_529,N_123,N_417);
nand U530 (N_530,N_81,N_80);
nand U531 (N_531,N_492,N_137);
nor U532 (N_532,N_270,N_194);
nand U533 (N_533,N_118,N_156);
xor U534 (N_534,N_357,N_454);
xor U535 (N_535,N_282,N_257);
and U536 (N_536,N_108,N_427);
nand U537 (N_537,N_294,N_177);
and U538 (N_538,N_397,N_400);
or U539 (N_539,N_442,N_258);
nor U540 (N_540,N_425,N_243);
nor U541 (N_541,N_9,N_1);
nand U542 (N_542,N_162,N_394);
and U543 (N_543,N_401,N_269);
nand U544 (N_544,N_134,N_489);
nand U545 (N_545,N_67,N_228);
xor U546 (N_546,N_55,N_239);
nand U547 (N_547,N_246,N_475);
and U548 (N_548,N_435,N_384);
nand U549 (N_549,N_146,N_342);
or U550 (N_550,N_232,N_250);
or U551 (N_551,N_464,N_178);
or U552 (N_552,N_259,N_314);
nor U553 (N_553,N_82,N_109);
and U554 (N_554,N_44,N_168);
xnor U555 (N_555,N_407,N_240);
xor U556 (N_556,N_268,N_132);
or U557 (N_557,N_110,N_71);
nand U558 (N_558,N_159,N_190);
xnor U559 (N_559,N_402,N_387);
xor U560 (N_560,N_151,N_256);
nor U561 (N_561,N_143,N_54);
xnor U562 (N_562,N_318,N_16);
nand U563 (N_563,N_399,N_79);
xor U564 (N_564,N_122,N_493);
or U565 (N_565,N_165,N_176);
nor U566 (N_566,N_385,N_431);
xnor U567 (N_567,N_86,N_117);
and U568 (N_568,N_169,N_390);
nor U569 (N_569,N_370,N_153);
nand U570 (N_570,N_303,N_448);
and U571 (N_571,N_313,N_47);
or U572 (N_572,N_104,N_481);
and U573 (N_573,N_391,N_443);
and U574 (N_574,N_344,N_17);
xnor U575 (N_575,N_141,N_85);
nor U576 (N_576,N_233,N_78);
xnor U577 (N_577,N_216,N_230);
or U578 (N_578,N_484,N_345);
xnor U579 (N_579,N_225,N_201);
nor U580 (N_580,N_480,N_33);
nand U581 (N_581,N_205,N_207);
or U582 (N_582,N_93,N_210);
or U583 (N_583,N_195,N_263);
nand U584 (N_584,N_12,N_349);
nor U585 (N_585,N_495,N_167);
nand U586 (N_586,N_488,N_362);
and U587 (N_587,N_276,N_32);
xor U588 (N_588,N_265,N_234);
or U589 (N_589,N_77,N_432);
nor U590 (N_590,N_158,N_170);
nor U591 (N_591,N_105,N_175);
nand U592 (N_592,N_193,N_26);
or U593 (N_593,N_467,N_236);
or U594 (N_594,N_283,N_436);
and U595 (N_595,N_354,N_308);
xnor U596 (N_596,N_472,N_405);
or U597 (N_597,N_301,N_457);
and U598 (N_598,N_372,N_99);
or U599 (N_599,N_174,N_266);
nand U600 (N_600,N_462,N_66);
nor U601 (N_601,N_56,N_202);
xor U602 (N_602,N_49,N_379);
or U603 (N_603,N_249,N_69);
and U604 (N_604,N_189,N_406);
xnor U605 (N_605,N_138,N_494);
and U606 (N_606,N_57,N_490);
and U607 (N_607,N_237,N_451);
or U608 (N_608,N_471,N_329);
and U609 (N_609,N_281,N_113);
xnor U610 (N_610,N_497,N_477);
nor U611 (N_611,N_386,N_459);
nor U612 (N_612,N_461,N_139);
or U613 (N_613,N_452,N_152);
or U614 (N_614,N_27,N_72);
and U615 (N_615,N_127,N_381);
or U616 (N_616,N_353,N_440);
xnor U617 (N_617,N_197,N_41);
xnor U618 (N_618,N_211,N_412);
or U619 (N_619,N_434,N_59);
and U620 (N_620,N_468,N_332);
nor U621 (N_621,N_382,N_53);
nor U622 (N_622,N_366,N_278);
xnor U623 (N_623,N_476,N_140);
xor U624 (N_624,N_430,N_135);
and U625 (N_625,N_333,N_439);
nor U626 (N_626,N_441,N_242);
nor U627 (N_627,N_87,N_90);
nor U628 (N_628,N_115,N_408);
and U629 (N_629,N_334,N_45);
and U630 (N_630,N_360,N_214);
nor U631 (N_631,N_478,N_446);
and U632 (N_632,N_395,N_286);
and U633 (N_633,N_284,N_198);
or U634 (N_634,N_28,N_97);
or U635 (N_635,N_280,N_319);
or U636 (N_636,N_111,N_217);
nand U637 (N_637,N_295,N_264);
nor U638 (N_638,N_470,N_279);
xnor U639 (N_639,N_5,N_460);
nand U640 (N_640,N_3,N_296);
nor U641 (N_641,N_496,N_365);
nor U642 (N_642,N_380,N_13);
or U643 (N_643,N_316,N_83);
nand U644 (N_644,N_116,N_180);
and U645 (N_645,N_274,N_368);
and U646 (N_646,N_445,N_235);
and U647 (N_647,N_38,N_157);
nand U648 (N_648,N_84,N_164);
and U649 (N_649,N_163,N_453);
or U650 (N_650,N_58,N_273);
xnor U651 (N_651,N_336,N_499);
and U652 (N_652,N_220,N_112);
or U653 (N_653,N_371,N_359);
xnor U654 (N_654,N_324,N_312);
or U655 (N_655,N_473,N_183);
or U656 (N_656,N_252,N_131);
and U657 (N_657,N_458,N_463);
xor U658 (N_658,N_449,N_260);
nor U659 (N_659,N_455,N_469);
nor U660 (N_660,N_215,N_227);
or U661 (N_661,N_466,N_222);
and U662 (N_662,N_369,N_348);
and U663 (N_663,N_120,N_292);
or U664 (N_664,N_290,N_6);
xor U665 (N_665,N_346,N_21);
or U666 (N_666,N_245,N_298);
nand U667 (N_667,N_289,N_275);
nand U668 (N_668,N_374,N_363);
and U669 (N_669,N_231,N_361);
or U670 (N_670,N_199,N_130);
nand U671 (N_671,N_34,N_311);
nand U672 (N_672,N_343,N_331);
xor U673 (N_673,N_491,N_433);
nand U674 (N_674,N_61,N_304);
or U675 (N_675,N_37,N_51);
and U676 (N_676,N_150,N_413);
and U677 (N_677,N_309,N_465);
nor U678 (N_678,N_101,N_106);
xor U679 (N_679,N_52,N_326);
nand U680 (N_680,N_10,N_485);
nor U681 (N_681,N_416,N_325);
nor U682 (N_682,N_241,N_421);
and U683 (N_683,N_96,N_383);
xnor U684 (N_684,N_208,N_187);
or U685 (N_685,N_181,N_418);
nor U686 (N_686,N_212,N_254);
nand U687 (N_687,N_25,N_68);
nor U688 (N_688,N_486,N_36);
nand U689 (N_689,N_447,N_330);
and U690 (N_690,N_307,N_437);
nor U691 (N_691,N_100,N_145);
or U692 (N_692,N_415,N_272);
nor U693 (N_693,N_306,N_429);
xor U694 (N_694,N_166,N_341);
or U695 (N_695,N_126,N_358);
nor U696 (N_696,N_352,N_7);
nand U697 (N_697,N_285,N_487);
xor U698 (N_698,N_92,N_98);
nor U699 (N_699,N_271,N_479);
xor U700 (N_700,N_20,N_321);
nand U701 (N_701,N_124,N_396);
xor U702 (N_702,N_456,N_74);
nor U703 (N_703,N_378,N_40);
nor U704 (N_704,N_262,N_119);
nand U705 (N_705,N_160,N_172);
and U706 (N_706,N_107,N_351);
nand U707 (N_707,N_184,N_91);
nor U708 (N_708,N_73,N_133);
xnor U709 (N_709,N_128,N_15);
nand U710 (N_710,N_209,N_200);
and U711 (N_711,N_48,N_377);
nand U712 (N_712,N_424,N_29);
xor U713 (N_713,N_102,N_192);
or U714 (N_714,N_404,N_62);
xor U715 (N_715,N_95,N_327);
nand U716 (N_716,N_393,N_75);
nand U717 (N_717,N_60,N_19);
nand U718 (N_718,N_30,N_403);
nand U719 (N_719,N_103,N_340);
or U720 (N_720,N_18,N_50);
and U721 (N_721,N_147,N_65);
and U722 (N_722,N_251,N_191);
or U723 (N_723,N_76,N_411);
or U724 (N_724,N_355,N_409);
and U725 (N_725,N_267,N_337);
nor U726 (N_726,N_204,N_203);
nor U727 (N_727,N_42,N_171);
and U728 (N_728,N_350,N_247);
xor U729 (N_729,N_206,N_226);
xor U730 (N_730,N_70,N_426);
nor U731 (N_731,N_88,N_136);
and U732 (N_732,N_182,N_388);
and U733 (N_733,N_322,N_186);
xnor U734 (N_734,N_277,N_423);
nand U735 (N_735,N_196,N_218);
nand U736 (N_736,N_375,N_121);
and U737 (N_737,N_155,N_114);
or U738 (N_738,N_161,N_398);
nand U739 (N_739,N_23,N_338);
or U740 (N_740,N_482,N_224);
nor U741 (N_741,N_315,N_291);
and U742 (N_742,N_221,N_310);
nand U743 (N_743,N_185,N_179);
nand U744 (N_744,N_14,N_428);
nor U745 (N_745,N_244,N_356);
and U746 (N_746,N_450,N_302);
and U747 (N_747,N_392,N_149);
or U748 (N_748,N_410,N_229);
and U749 (N_749,N_422,N_22);
nor U750 (N_750,N_322,N_37);
nor U751 (N_751,N_284,N_55);
or U752 (N_752,N_471,N_495);
nand U753 (N_753,N_268,N_154);
xnor U754 (N_754,N_482,N_94);
and U755 (N_755,N_143,N_93);
or U756 (N_756,N_439,N_74);
or U757 (N_757,N_386,N_315);
xnor U758 (N_758,N_356,N_213);
xnor U759 (N_759,N_111,N_104);
and U760 (N_760,N_320,N_400);
or U761 (N_761,N_358,N_141);
xor U762 (N_762,N_180,N_447);
nor U763 (N_763,N_339,N_301);
and U764 (N_764,N_318,N_372);
or U765 (N_765,N_74,N_62);
xnor U766 (N_766,N_239,N_495);
nor U767 (N_767,N_242,N_268);
and U768 (N_768,N_11,N_266);
or U769 (N_769,N_246,N_370);
xor U770 (N_770,N_275,N_267);
and U771 (N_771,N_182,N_465);
xnor U772 (N_772,N_425,N_466);
nand U773 (N_773,N_101,N_300);
xor U774 (N_774,N_103,N_378);
and U775 (N_775,N_295,N_441);
or U776 (N_776,N_415,N_242);
and U777 (N_777,N_320,N_231);
nor U778 (N_778,N_325,N_197);
and U779 (N_779,N_41,N_229);
nand U780 (N_780,N_496,N_458);
and U781 (N_781,N_8,N_272);
nand U782 (N_782,N_335,N_177);
nor U783 (N_783,N_451,N_191);
xor U784 (N_784,N_412,N_284);
xor U785 (N_785,N_337,N_478);
and U786 (N_786,N_425,N_337);
xor U787 (N_787,N_202,N_41);
nand U788 (N_788,N_240,N_226);
xnor U789 (N_789,N_119,N_452);
or U790 (N_790,N_23,N_5);
or U791 (N_791,N_267,N_147);
nand U792 (N_792,N_375,N_399);
or U793 (N_793,N_104,N_165);
nand U794 (N_794,N_472,N_3);
nor U795 (N_795,N_139,N_285);
and U796 (N_796,N_457,N_171);
xor U797 (N_797,N_418,N_115);
and U798 (N_798,N_74,N_109);
xnor U799 (N_799,N_496,N_14);
or U800 (N_800,N_351,N_424);
or U801 (N_801,N_346,N_474);
nor U802 (N_802,N_27,N_314);
and U803 (N_803,N_361,N_4);
or U804 (N_804,N_446,N_453);
and U805 (N_805,N_267,N_72);
and U806 (N_806,N_355,N_211);
nand U807 (N_807,N_163,N_233);
nor U808 (N_808,N_281,N_66);
nand U809 (N_809,N_213,N_63);
nor U810 (N_810,N_382,N_73);
and U811 (N_811,N_265,N_334);
or U812 (N_812,N_43,N_383);
nand U813 (N_813,N_146,N_393);
nor U814 (N_814,N_6,N_213);
nand U815 (N_815,N_192,N_348);
xor U816 (N_816,N_261,N_425);
nand U817 (N_817,N_331,N_32);
nor U818 (N_818,N_73,N_274);
nor U819 (N_819,N_375,N_268);
and U820 (N_820,N_238,N_20);
nor U821 (N_821,N_61,N_1);
nor U822 (N_822,N_171,N_244);
or U823 (N_823,N_193,N_137);
nor U824 (N_824,N_407,N_239);
xnor U825 (N_825,N_344,N_129);
nand U826 (N_826,N_51,N_140);
and U827 (N_827,N_281,N_413);
or U828 (N_828,N_461,N_175);
nand U829 (N_829,N_41,N_434);
nor U830 (N_830,N_463,N_282);
and U831 (N_831,N_429,N_336);
nand U832 (N_832,N_154,N_255);
xor U833 (N_833,N_156,N_198);
nor U834 (N_834,N_84,N_214);
nor U835 (N_835,N_7,N_168);
or U836 (N_836,N_16,N_65);
nand U837 (N_837,N_445,N_149);
nor U838 (N_838,N_377,N_367);
xnor U839 (N_839,N_272,N_356);
xor U840 (N_840,N_463,N_473);
xnor U841 (N_841,N_238,N_75);
and U842 (N_842,N_382,N_210);
nor U843 (N_843,N_316,N_9);
or U844 (N_844,N_171,N_7);
and U845 (N_845,N_440,N_402);
nand U846 (N_846,N_414,N_162);
xor U847 (N_847,N_26,N_64);
nor U848 (N_848,N_46,N_310);
nor U849 (N_849,N_9,N_22);
nand U850 (N_850,N_306,N_288);
or U851 (N_851,N_270,N_205);
and U852 (N_852,N_426,N_209);
nor U853 (N_853,N_286,N_119);
and U854 (N_854,N_132,N_37);
nand U855 (N_855,N_426,N_85);
xor U856 (N_856,N_66,N_292);
nor U857 (N_857,N_383,N_318);
and U858 (N_858,N_308,N_224);
and U859 (N_859,N_18,N_62);
nand U860 (N_860,N_162,N_190);
and U861 (N_861,N_282,N_414);
and U862 (N_862,N_312,N_255);
nor U863 (N_863,N_226,N_59);
or U864 (N_864,N_430,N_471);
nor U865 (N_865,N_11,N_219);
xor U866 (N_866,N_32,N_246);
xnor U867 (N_867,N_6,N_63);
and U868 (N_868,N_166,N_128);
and U869 (N_869,N_275,N_298);
and U870 (N_870,N_300,N_226);
nor U871 (N_871,N_432,N_135);
xor U872 (N_872,N_39,N_18);
or U873 (N_873,N_488,N_367);
and U874 (N_874,N_327,N_499);
nand U875 (N_875,N_417,N_240);
and U876 (N_876,N_330,N_166);
xnor U877 (N_877,N_467,N_493);
or U878 (N_878,N_312,N_396);
nor U879 (N_879,N_77,N_43);
or U880 (N_880,N_217,N_460);
or U881 (N_881,N_147,N_56);
nand U882 (N_882,N_383,N_336);
xnor U883 (N_883,N_259,N_107);
xor U884 (N_884,N_460,N_426);
xnor U885 (N_885,N_170,N_124);
xnor U886 (N_886,N_366,N_267);
nor U887 (N_887,N_106,N_225);
and U888 (N_888,N_67,N_33);
and U889 (N_889,N_484,N_410);
or U890 (N_890,N_269,N_469);
or U891 (N_891,N_486,N_27);
or U892 (N_892,N_205,N_20);
or U893 (N_893,N_319,N_163);
and U894 (N_894,N_250,N_66);
or U895 (N_895,N_124,N_341);
nand U896 (N_896,N_391,N_375);
or U897 (N_897,N_439,N_387);
or U898 (N_898,N_305,N_12);
nand U899 (N_899,N_468,N_93);
nand U900 (N_900,N_270,N_146);
nor U901 (N_901,N_223,N_131);
nand U902 (N_902,N_453,N_158);
nand U903 (N_903,N_285,N_328);
or U904 (N_904,N_361,N_84);
and U905 (N_905,N_353,N_417);
and U906 (N_906,N_36,N_400);
nor U907 (N_907,N_178,N_311);
nand U908 (N_908,N_192,N_303);
or U909 (N_909,N_109,N_165);
and U910 (N_910,N_278,N_240);
and U911 (N_911,N_219,N_444);
nor U912 (N_912,N_370,N_238);
nand U913 (N_913,N_106,N_385);
xor U914 (N_914,N_7,N_43);
and U915 (N_915,N_398,N_100);
xor U916 (N_916,N_329,N_136);
xor U917 (N_917,N_181,N_150);
nor U918 (N_918,N_273,N_339);
and U919 (N_919,N_455,N_100);
nor U920 (N_920,N_200,N_346);
and U921 (N_921,N_20,N_374);
nor U922 (N_922,N_321,N_331);
xor U923 (N_923,N_252,N_463);
or U924 (N_924,N_12,N_1);
xnor U925 (N_925,N_22,N_221);
or U926 (N_926,N_469,N_320);
and U927 (N_927,N_277,N_466);
or U928 (N_928,N_416,N_8);
nor U929 (N_929,N_381,N_233);
and U930 (N_930,N_36,N_355);
nor U931 (N_931,N_55,N_101);
nor U932 (N_932,N_397,N_375);
nand U933 (N_933,N_426,N_244);
nor U934 (N_934,N_116,N_82);
nor U935 (N_935,N_479,N_171);
nor U936 (N_936,N_405,N_74);
xor U937 (N_937,N_231,N_476);
nand U938 (N_938,N_98,N_24);
nand U939 (N_939,N_178,N_56);
nor U940 (N_940,N_348,N_307);
xnor U941 (N_941,N_499,N_326);
xnor U942 (N_942,N_399,N_192);
xor U943 (N_943,N_175,N_211);
or U944 (N_944,N_273,N_80);
nand U945 (N_945,N_397,N_340);
xnor U946 (N_946,N_327,N_57);
xor U947 (N_947,N_353,N_197);
xor U948 (N_948,N_5,N_176);
xor U949 (N_949,N_333,N_187);
nand U950 (N_950,N_404,N_89);
or U951 (N_951,N_241,N_55);
nand U952 (N_952,N_178,N_382);
nor U953 (N_953,N_41,N_374);
or U954 (N_954,N_359,N_447);
or U955 (N_955,N_360,N_166);
or U956 (N_956,N_324,N_171);
xor U957 (N_957,N_46,N_316);
nor U958 (N_958,N_311,N_26);
nor U959 (N_959,N_334,N_212);
and U960 (N_960,N_370,N_15);
or U961 (N_961,N_300,N_333);
and U962 (N_962,N_338,N_59);
nand U963 (N_963,N_440,N_22);
nor U964 (N_964,N_188,N_458);
nand U965 (N_965,N_375,N_356);
nand U966 (N_966,N_114,N_21);
nor U967 (N_967,N_103,N_285);
and U968 (N_968,N_410,N_479);
and U969 (N_969,N_429,N_473);
nor U970 (N_970,N_192,N_167);
xnor U971 (N_971,N_376,N_290);
nor U972 (N_972,N_217,N_327);
nand U973 (N_973,N_42,N_83);
xnor U974 (N_974,N_465,N_125);
xnor U975 (N_975,N_33,N_445);
and U976 (N_976,N_53,N_259);
nor U977 (N_977,N_266,N_493);
and U978 (N_978,N_269,N_356);
or U979 (N_979,N_248,N_236);
xnor U980 (N_980,N_455,N_10);
nor U981 (N_981,N_26,N_342);
nand U982 (N_982,N_151,N_485);
and U983 (N_983,N_441,N_195);
nand U984 (N_984,N_124,N_490);
nor U985 (N_985,N_457,N_177);
or U986 (N_986,N_177,N_411);
xor U987 (N_987,N_21,N_23);
nand U988 (N_988,N_85,N_306);
or U989 (N_989,N_248,N_45);
and U990 (N_990,N_325,N_82);
and U991 (N_991,N_487,N_401);
and U992 (N_992,N_5,N_417);
nor U993 (N_993,N_351,N_82);
or U994 (N_994,N_237,N_31);
and U995 (N_995,N_480,N_29);
nor U996 (N_996,N_428,N_200);
xnor U997 (N_997,N_247,N_68);
nor U998 (N_998,N_157,N_405);
nor U999 (N_999,N_286,N_337);
and U1000 (N_1000,N_536,N_524);
nand U1001 (N_1001,N_513,N_599);
nand U1002 (N_1002,N_967,N_841);
xnor U1003 (N_1003,N_579,N_801);
nand U1004 (N_1004,N_811,N_635);
and U1005 (N_1005,N_937,N_766);
xor U1006 (N_1006,N_807,N_709);
and U1007 (N_1007,N_794,N_743);
or U1008 (N_1008,N_637,N_974);
nor U1009 (N_1009,N_695,N_726);
or U1010 (N_1010,N_580,N_895);
nor U1011 (N_1011,N_976,N_878);
xnor U1012 (N_1012,N_836,N_804);
xor U1013 (N_1013,N_710,N_916);
nand U1014 (N_1014,N_805,N_894);
nor U1015 (N_1015,N_950,N_938);
or U1016 (N_1016,N_633,N_778);
or U1017 (N_1017,N_500,N_682);
and U1018 (N_1018,N_642,N_997);
xor U1019 (N_1019,N_831,N_686);
or U1020 (N_1020,N_575,N_622);
or U1021 (N_1021,N_936,N_738);
nand U1022 (N_1022,N_854,N_824);
nand U1023 (N_1023,N_578,N_549);
nor U1024 (N_1024,N_702,N_505);
xor U1025 (N_1025,N_888,N_918);
nand U1026 (N_1026,N_872,N_977);
or U1027 (N_1027,N_969,N_657);
or U1028 (N_1028,N_693,N_626);
xor U1029 (N_1029,N_874,N_930);
xor U1030 (N_1030,N_763,N_866);
xnor U1031 (N_1031,N_561,N_896);
nor U1032 (N_1032,N_986,N_511);
nor U1033 (N_1033,N_776,N_679);
and U1034 (N_1034,N_596,N_647);
or U1035 (N_1035,N_760,N_759);
nand U1036 (N_1036,N_809,N_560);
and U1037 (N_1037,N_671,N_761);
nor U1038 (N_1038,N_857,N_884);
nand U1039 (N_1039,N_948,N_779);
nor U1040 (N_1040,N_924,N_912);
and U1041 (N_1041,N_898,N_564);
or U1042 (N_1042,N_654,N_961);
xnor U1043 (N_1043,N_661,N_973);
or U1044 (N_1044,N_822,N_725);
and U1045 (N_1045,N_631,N_586);
or U1046 (N_1046,N_862,N_900);
nand U1047 (N_1047,N_909,N_964);
nand U1048 (N_1048,N_814,N_947);
or U1049 (N_1049,N_920,N_603);
nand U1050 (N_1050,N_750,N_843);
nor U1051 (N_1051,N_864,N_887);
nand U1052 (N_1052,N_672,N_777);
nand U1053 (N_1053,N_565,N_503);
and U1054 (N_1054,N_837,N_845);
nor U1055 (N_1055,N_543,N_528);
and U1056 (N_1056,N_933,N_975);
nor U1057 (N_1057,N_703,N_574);
and U1058 (N_1058,N_704,N_753);
and U1059 (N_1059,N_819,N_717);
or U1060 (N_1060,N_567,N_917);
nor U1061 (N_1061,N_956,N_802);
and U1062 (N_1062,N_606,N_516);
or U1063 (N_1063,N_628,N_501);
and U1064 (N_1064,N_576,N_506);
xnor U1065 (N_1065,N_752,N_651);
or U1066 (N_1066,N_867,N_714);
nand U1067 (N_1067,N_572,N_544);
nor U1068 (N_1068,N_548,N_582);
nor U1069 (N_1069,N_529,N_515);
nor U1070 (N_1070,N_624,N_984);
nand U1071 (N_1071,N_768,N_834);
xor U1072 (N_1072,N_663,N_786);
nand U1073 (N_1073,N_553,N_829);
xor U1074 (N_1074,N_527,N_632);
nand U1075 (N_1075,N_988,N_873);
nor U1076 (N_1076,N_530,N_838);
nor U1077 (N_1077,N_616,N_966);
xor U1078 (N_1078,N_788,N_792);
xor U1079 (N_1079,N_540,N_537);
and U1080 (N_1080,N_615,N_604);
or U1081 (N_1081,N_683,N_817);
nor U1082 (N_1082,N_740,N_625);
nor U1083 (N_1083,N_652,N_711);
and U1084 (N_1084,N_601,N_634);
nor U1085 (N_1085,N_876,N_828);
and U1086 (N_1086,N_668,N_787);
and U1087 (N_1087,N_853,N_655);
nor U1088 (N_1088,N_612,N_932);
or U1089 (N_1089,N_534,N_989);
nor U1090 (N_1090,N_546,N_605);
xnor U1091 (N_1091,N_823,N_629);
xor U1092 (N_1092,N_730,N_520);
nor U1093 (N_1093,N_563,N_600);
nand U1094 (N_1094,N_803,N_734);
nand U1095 (N_1095,N_889,N_774);
xor U1096 (N_1096,N_698,N_861);
and U1097 (N_1097,N_885,N_521);
xor U1098 (N_1098,N_636,N_813);
and U1099 (N_1099,N_638,N_700);
or U1100 (N_1100,N_958,N_992);
xor U1101 (N_1101,N_644,N_670);
and U1102 (N_1102,N_990,N_656);
nand U1103 (N_1103,N_689,N_598);
xor U1104 (N_1104,N_588,N_550);
and U1105 (N_1105,N_554,N_962);
nor U1106 (N_1106,N_852,N_971);
nand U1107 (N_1107,N_535,N_609);
nand U1108 (N_1108,N_662,N_556);
xnor U1109 (N_1109,N_681,N_849);
or U1110 (N_1110,N_945,N_509);
xor U1111 (N_1111,N_733,N_705);
nand U1112 (N_1112,N_562,N_905);
xnor U1113 (N_1113,N_879,N_542);
or U1114 (N_1114,N_739,N_840);
xnor U1115 (N_1115,N_869,N_951);
or U1116 (N_1116,N_558,N_648);
nand U1117 (N_1117,N_999,N_593);
nor U1118 (N_1118,N_890,N_815);
nor U1119 (N_1119,N_970,N_782);
and U1120 (N_1120,N_687,N_927);
xnor U1121 (N_1121,N_968,N_883);
xnor U1122 (N_1122,N_858,N_594);
and U1123 (N_1123,N_627,N_832);
and U1124 (N_1124,N_602,N_863);
nor U1125 (N_1125,N_724,N_676);
nor U1126 (N_1126,N_694,N_965);
nand U1127 (N_1127,N_827,N_772);
nand U1128 (N_1128,N_908,N_780);
nand U1129 (N_1129,N_931,N_796);
or U1130 (N_1130,N_795,N_756);
nand U1131 (N_1131,N_715,N_696);
or U1132 (N_1132,N_621,N_706);
or U1133 (N_1133,N_868,N_899);
and U1134 (N_1134,N_959,N_806);
nand U1135 (N_1135,N_886,N_746);
and U1136 (N_1136,N_762,N_685);
nand U1137 (N_1137,N_764,N_941);
nor U1138 (N_1138,N_793,N_666);
nand U1139 (N_1139,N_699,N_915);
nor U1140 (N_1140,N_691,N_566);
or U1141 (N_1141,N_728,N_820);
and U1142 (N_1142,N_587,N_667);
or U1143 (N_1143,N_773,N_720);
nor U1144 (N_1144,N_789,N_929);
xnor U1145 (N_1145,N_904,N_851);
nor U1146 (N_1146,N_673,N_641);
xnor U1147 (N_1147,N_846,N_590);
xor U1148 (N_1148,N_881,N_640);
or U1149 (N_1149,N_865,N_850);
xor U1150 (N_1150,N_519,N_979);
xor U1151 (N_1151,N_911,N_754);
or U1152 (N_1152,N_713,N_983);
nand U1153 (N_1153,N_906,N_613);
or U1154 (N_1154,N_810,N_901);
or U1155 (N_1155,N_835,N_716);
nor U1156 (N_1156,N_591,N_559);
nor U1157 (N_1157,N_649,N_860);
nor U1158 (N_1158,N_953,N_923);
nor U1159 (N_1159,N_645,N_955);
xnor U1160 (N_1160,N_981,N_741);
xnor U1161 (N_1161,N_531,N_914);
and U1162 (N_1162,N_557,N_934);
nor U1163 (N_1163,N_826,N_848);
and U1164 (N_1164,N_978,N_880);
or U1165 (N_1165,N_607,N_985);
and U1166 (N_1166,N_926,N_551);
or U1167 (N_1167,N_569,N_833);
nor U1168 (N_1168,N_946,N_610);
or U1169 (N_1169,N_620,N_922);
and U1170 (N_1170,N_944,N_508);
or U1171 (N_1171,N_630,N_785);
nor U1172 (N_1172,N_902,N_907);
xnor U1173 (N_1173,N_545,N_690);
xor U1174 (N_1174,N_532,N_585);
xor U1175 (N_1175,N_928,N_856);
nor U1176 (N_1176,N_547,N_943);
nor U1177 (N_1177,N_584,N_993);
and U1178 (N_1178,N_664,N_581);
nor U1179 (N_1179,N_619,N_921);
nor U1180 (N_1180,N_723,N_707);
or U1181 (N_1181,N_758,N_712);
or U1182 (N_1182,N_684,N_816);
nor U1183 (N_1183,N_675,N_942);
or U1184 (N_1184,N_538,N_517);
xor U1185 (N_1185,N_893,N_790);
nand U1186 (N_1186,N_775,N_688);
nor U1187 (N_1187,N_963,N_617);
nand U1188 (N_1188,N_749,N_618);
or U1189 (N_1189,N_994,N_646);
and U1190 (N_1190,N_504,N_589);
nor U1191 (N_1191,N_514,N_897);
xnor U1192 (N_1192,N_882,N_518);
or U1193 (N_1193,N_939,N_744);
nor U1194 (N_1194,N_658,N_952);
or U1195 (N_1195,N_525,N_954);
or U1196 (N_1196,N_697,N_957);
or U1197 (N_1197,N_727,N_680);
and U1198 (N_1198,N_665,N_650);
xor U1199 (N_1199,N_996,N_653);
or U1200 (N_1200,N_757,N_842);
xnor U1201 (N_1201,N_982,N_643);
nor U1202 (N_1202,N_701,N_770);
nor U1203 (N_1203,N_592,N_614);
nand U1204 (N_1204,N_799,N_731);
xor U1205 (N_1205,N_745,N_742);
and U1206 (N_1206,N_597,N_674);
nor U1207 (N_1207,N_783,N_771);
or U1208 (N_1208,N_639,N_608);
or U1209 (N_1209,N_583,N_830);
nor U1210 (N_1210,N_847,N_818);
nand U1211 (N_1211,N_722,N_735);
or U1212 (N_1212,N_972,N_748);
and U1213 (N_1213,N_767,N_747);
nor U1214 (N_1214,N_659,N_555);
or U1215 (N_1215,N_736,N_808);
nor U1216 (N_1216,N_595,N_870);
and U1217 (N_1217,N_791,N_825);
and U1218 (N_1218,N_577,N_755);
nand U1219 (N_1219,N_732,N_510);
nand U1220 (N_1220,N_692,N_903);
xor U1221 (N_1221,N_708,N_910);
nor U1222 (N_1222,N_980,N_839);
nor U1223 (N_1223,N_573,N_539);
nand U1224 (N_1224,N_859,N_512);
nand U1225 (N_1225,N_721,N_960);
xnor U1226 (N_1226,N_797,N_913);
or U1227 (N_1227,N_729,N_678);
nand U1228 (N_1228,N_998,N_892);
and U1229 (N_1229,N_719,N_919);
xnor U1230 (N_1230,N_891,N_781);
and U1231 (N_1231,N_995,N_526);
and U1232 (N_1232,N_935,N_751);
and U1233 (N_1233,N_669,N_844);
or U1234 (N_1234,N_568,N_507);
nor U1235 (N_1235,N_570,N_533);
and U1236 (N_1236,N_677,N_800);
and U1237 (N_1237,N_871,N_737);
or U1238 (N_1238,N_855,N_769);
and U1239 (N_1239,N_660,N_502);
nor U1240 (N_1240,N_522,N_949);
and U1241 (N_1241,N_718,N_940);
nand U1242 (N_1242,N_821,N_541);
or U1243 (N_1243,N_875,N_877);
and U1244 (N_1244,N_925,N_798);
or U1245 (N_1245,N_765,N_812);
nor U1246 (N_1246,N_991,N_571);
or U1247 (N_1247,N_987,N_523);
xor U1248 (N_1248,N_552,N_623);
nand U1249 (N_1249,N_611,N_784);
and U1250 (N_1250,N_771,N_828);
xnor U1251 (N_1251,N_590,N_994);
nor U1252 (N_1252,N_626,N_968);
nor U1253 (N_1253,N_888,N_551);
and U1254 (N_1254,N_879,N_875);
nor U1255 (N_1255,N_907,N_672);
nor U1256 (N_1256,N_881,N_951);
and U1257 (N_1257,N_908,N_685);
or U1258 (N_1258,N_539,N_967);
nand U1259 (N_1259,N_685,N_610);
nand U1260 (N_1260,N_614,N_875);
and U1261 (N_1261,N_595,N_572);
and U1262 (N_1262,N_947,N_506);
and U1263 (N_1263,N_602,N_561);
nand U1264 (N_1264,N_592,N_632);
nor U1265 (N_1265,N_934,N_997);
xnor U1266 (N_1266,N_831,N_960);
xnor U1267 (N_1267,N_719,N_541);
and U1268 (N_1268,N_981,N_857);
nor U1269 (N_1269,N_538,N_533);
xor U1270 (N_1270,N_690,N_920);
nand U1271 (N_1271,N_940,N_652);
xnor U1272 (N_1272,N_982,N_703);
and U1273 (N_1273,N_705,N_662);
and U1274 (N_1274,N_763,N_677);
nor U1275 (N_1275,N_726,N_696);
nor U1276 (N_1276,N_990,N_809);
xnor U1277 (N_1277,N_921,N_856);
and U1278 (N_1278,N_856,N_759);
nand U1279 (N_1279,N_923,N_538);
or U1280 (N_1280,N_624,N_986);
nor U1281 (N_1281,N_562,N_738);
xor U1282 (N_1282,N_893,N_595);
or U1283 (N_1283,N_645,N_519);
and U1284 (N_1284,N_739,N_928);
and U1285 (N_1285,N_919,N_501);
and U1286 (N_1286,N_626,N_738);
or U1287 (N_1287,N_914,N_936);
nor U1288 (N_1288,N_677,N_821);
nor U1289 (N_1289,N_563,N_842);
and U1290 (N_1290,N_501,N_829);
or U1291 (N_1291,N_541,N_793);
xor U1292 (N_1292,N_545,N_791);
and U1293 (N_1293,N_919,N_643);
and U1294 (N_1294,N_888,N_957);
and U1295 (N_1295,N_669,N_990);
xnor U1296 (N_1296,N_608,N_726);
nor U1297 (N_1297,N_841,N_740);
or U1298 (N_1298,N_609,N_852);
xnor U1299 (N_1299,N_841,N_951);
xor U1300 (N_1300,N_724,N_654);
nand U1301 (N_1301,N_708,N_882);
and U1302 (N_1302,N_912,N_802);
nand U1303 (N_1303,N_876,N_517);
or U1304 (N_1304,N_997,N_603);
and U1305 (N_1305,N_509,N_899);
or U1306 (N_1306,N_795,N_535);
or U1307 (N_1307,N_607,N_600);
and U1308 (N_1308,N_767,N_737);
xor U1309 (N_1309,N_575,N_606);
nand U1310 (N_1310,N_788,N_921);
and U1311 (N_1311,N_899,N_752);
or U1312 (N_1312,N_504,N_888);
nor U1313 (N_1313,N_768,N_609);
and U1314 (N_1314,N_809,N_910);
or U1315 (N_1315,N_790,N_954);
and U1316 (N_1316,N_752,N_531);
nor U1317 (N_1317,N_908,N_587);
nand U1318 (N_1318,N_645,N_815);
nor U1319 (N_1319,N_894,N_898);
and U1320 (N_1320,N_502,N_803);
nand U1321 (N_1321,N_847,N_913);
nand U1322 (N_1322,N_628,N_984);
nand U1323 (N_1323,N_749,N_556);
xor U1324 (N_1324,N_738,N_823);
nand U1325 (N_1325,N_523,N_530);
nand U1326 (N_1326,N_866,N_676);
xor U1327 (N_1327,N_597,N_751);
and U1328 (N_1328,N_830,N_846);
or U1329 (N_1329,N_530,N_765);
xnor U1330 (N_1330,N_849,N_971);
or U1331 (N_1331,N_808,N_643);
nand U1332 (N_1332,N_664,N_745);
or U1333 (N_1333,N_973,N_699);
and U1334 (N_1334,N_782,N_723);
or U1335 (N_1335,N_542,N_633);
xnor U1336 (N_1336,N_750,N_504);
nor U1337 (N_1337,N_681,N_879);
and U1338 (N_1338,N_522,N_899);
xor U1339 (N_1339,N_904,N_960);
or U1340 (N_1340,N_774,N_956);
and U1341 (N_1341,N_703,N_828);
nor U1342 (N_1342,N_893,N_622);
xnor U1343 (N_1343,N_718,N_838);
and U1344 (N_1344,N_862,N_863);
and U1345 (N_1345,N_544,N_775);
nand U1346 (N_1346,N_881,N_637);
or U1347 (N_1347,N_669,N_549);
or U1348 (N_1348,N_615,N_992);
xor U1349 (N_1349,N_510,N_665);
or U1350 (N_1350,N_547,N_528);
nand U1351 (N_1351,N_688,N_986);
xor U1352 (N_1352,N_932,N_820);
nor U1353 (N_1353,N_630,N_727);
and U1354 (N_1354,N_989,N_920);
and U1355 (N_1355,N_660,N_624);
xnor U1356 (N_1356,N_957,N_819);
nor U1357 (N_1357,N_609,N_746);
xnor U1358 (N_1358,N_606,N_788);
or U1359 (N_1359,N_829,N_660);
nor U1360 (N_1360,N_786,N_739);
xnor U1361 (N_1361,N_597,N_985);
nor U1362 (N_1362,N_554,N_862);
nand U1363 (N_1363,N_595,N_849);
xnor U1364 (N_1364,N_735,N_852);
nor U1365 (N_1365,N_935,N_609);
nor U1366 (N_1366,N_583,N_724);
xnor U1367 (N_1367,N_776,N_729);
or U1368 (N_1368,N_605,N_809);
or U1369 (N_1369,N_895,N_799);
nor U1370 (N_1370,N_735,N_619);
xnor U1371 (N_1371,N_941,N_551);
nor U1372 (N_1372,N_543,N_870);
nor U1373 (N_1373,N_623,N_530);
nor U1374 (N_1374,N_966,N_981);
and U1375 (N_1375,N_896,N_506);
or U1376 (N_1376,N_911,N_596);
and U1377 (N_1377,N_624,N_800);
or U1378 (N_1378,N_764,N_556);
or U1379 (N_1379,N_943,N_657);
or U1380 (N_1380,N_534,N_821);
nand U1381 (N_1381,N_536,N_679);
or U1382 (N_1382,N_701,N_968);
nand U1383 (N_1383,N_536,N_827);
nand U1384 (N_1384,N_623,N_833);
nor U1385 (N_1385,N_878,N_633);
xnor U1386 (N_1386,N_844,N_629);
and U1387 (N_1387,N_613,N_861);
and U1388 (N_1388,N_843,N_652);
nor U1389 (N_1389,N_791,N_645);
and U1390 (N_1390,N_775,N_769);
nor U1391 (N_1391,N_939,N_655);
and U1392 (N_1392,N_709,N_953);
or U1393 (N_1393,N_920,N_960);
xor U1394 (N_1394,N_890,N_795);
and U1395 (N_1395,N_523,N_656);
or U1396 (N_1396,N_894,N_767);
nand U1397 (N_1397,N_985,N_646);
and U1398 (N_1398,N_522,N_910);
nor U1399 (N_1399,N_821,N_988);
or U1400 (N_1400,N_660,N_961);
and U1401 (N_1401,N_957,N_669);
xor U1402 (N_1402,N_716,N_671);
nand U1403 (N_1403,N_905,N_573);
nand U1404 (N_1404,N_835,N_888);
nand U1405 (N_1405,N_866,N_977);
nand U1406 (N_1406,N_621,N_804);
nand U1407 (N_1407,N_560,N_554);
xor U1408 (N_1408,N_936,N_870);
or U1409 (N_1409,N_776,N_654);
xor U1410 (N_1410,N_993,N_518);
nand U1411 (N_1411,N_891,N_712);
xnor U1412 (N_1412,N_715,N_802);
nor U1413 (N_1413,N_861,N_726);
nor U1414 (N_1414,N_974,N_942);
nand U1415 (N_1415,N_824,N_815);
nand U1416 (N_1416,N_672,N_778);
and U1417 (N_1417,N_509,N_783);
xor U1418 (N_1418,N_929,N_837);
and U1419 (N_1419,N_524,N_982);
nor U1420 (N_1420,N_560,N_730);
or U1421 (N_1421,N_942,N_816);
nor U1422 (N_1422,N_517,N_653);
nor U1423 (N_1423,N_615,N_697);
xnor U1424 (N_1424,N_732,N_599);
nor U1425 (N_1425,N_554,N_755);
nand U1426 (N_1426,N_850,N_785);
nor U1427 (N_1427,N_942,N_622);
nor U1428 (N_1428,N_709,N_955);
nand U1429 (N_1429,N_601,N_970);
or U1430 (N_1430,N_984,N_934);
nor U1431 (N_1431,N_787,N_905);
and U1432 (N_1432,N_954,N_824);
or U1433 (N_1433,N_599,N_706);
nor U1434 (N_1434,N_670,N_529);
and U1435 (N_1435,N_525,N_612);
xor U1436 (N_1436,N_784,N_752);
nor U1437 (N_1437,N_883,N_927);
xor U1438 (N_1438,N_823,N_772);
xnor U1439 (N_1439,N_823,N_508);
xnor U1440 (N_1440,N_791,N_535);
and U1441 (N_1441,N_834,N_612);
nor U1442 (N_1442,N_750,N_534);
nand U1443 (N_1443,N_844,N_548);
or U1444 (N_1444,N_786,N_655);
or U1445 (N_1445,N_849,N_979);
and U1446 (N_1446,N_699,N_953);
nor U1447 (N_1447,N_767,N_521);
xnor U1448 (N_1448,N_691,N_891);
nand U1449 (N_1449,N_604,N_653);
or U1450 (N_1450,N_769,N_947);
nand U1451 (N_1451,N_706,N_798);
and U1452 (N_1452,N_940,N_814);
or U1453 (N_1453,N_741,N_770);
and U1454 (N_1454,N_993,N_722);
nor U1455 (N_1455,N_735,N_710);
nor U1456 (N_1456,N_698,N_824);
and U1457 (N_1457,N_713,N_590);
xor U1458 (N_1458,N_522,N_883);
xor U1459 (N_1459,N_939,N_612);
nand U1460 (N_1460,N_844,N_821);
nand U1461 (N_1461,N_779,N_747);
or U1462 (N_1462,N_545,N_944);
nand U1463 (N_1463,N_962,N_602);
nor U1464 (N_1464,N_969,N_811);
or U1465 (N_1465,N_798,N_612);
and U1466 (N_1466,N_535,N_863);
nor U1467 (N_1467,N_616,N_652);
nand U1468 (N_1468,N_908,N_973);
and U1469 (N_1469,N_843,N_589);
nor U1470 (N_1470,N_557,N_803);
or U1471 (N_1471,N_691,N_780);
nand U1472 (N_1472,N_659,N_704);
or U1473 (N_1473,N_837,N_995);
or U1474 (N_1474,N_640,N_545);
nand U1475 (N_1475,N_925,N_552);
nand U1476 (N_1476,N_537,N_921);
xnor U1477 (N_1477,N_603,N_715);
nor U1478 (N_1478,N_502,N_515);
nor U1479 (N_1479,N_536,N_925);
xor U1480 (N_1480,N_912,N_823);
or U1481 (N_1481,N_696,N_624);
or U1482 (N_1482,N_898,N_822);
and U1483 (N_1483,N_956,N_622);
or U1484 (N_1484,N_571,N_727);
and U1485 (N_1485,N_659,N_566);
nand U1486 (N_1486,N_519,N_708);
nor U1487 (N_1487,N_858,N_874);
and U1488 (N_1488,N_656,N_680);
or U1489 (N_1489,N_512,N_860);
nand U1490 (N_1490,N_974,N_958);
or U1491 (N_1491,N_761,N_932);
xnor U1492 (N_1492,N_618,N_807);
nor U1493 (N_1493,N_592,N_731);
nand U1494 (N_1494,N_765,N_966);
nor U1495 (N_1495,N_682,N_945);
xnor U1496 (N_1496,N_665,N_587);
xor U1497 (N_1497,N_602,N_889);
nand U1498 (N_1498,N_531,N_655);
or U1499 (N_1499,N_752,N_821);
and U1500 (N_1500,N_1008,N_1478);
and U1501 (N_1501,N_1455,N_1291);
or U1502 (N_1502,N_1149,N_1301);
nor U1503 (N_1503,N_1389,N_1207);
and U1504 (N_1504,N_1095,N_1175);
xnor U1505 (N_1505,N_1036,N_1374);
xnor U1506 (N_1506,N_1002,N_1040);
xor U1507 (N_1507,N_1365,N_1385);
nor U1508 (N_1508,N_1080,N_1091);
xor U1509 (N_1509,N_1360,N_1174);
xnor U1510 (N_1510,N_1251,N_1458);
nand U1511 (N_1511,N_1266,N_1220);
or U1512 (N_1512,N_1429,N_1334);
xnor U1513 (N_1513,N_1394,N_1336);
or U1514 (N_1514,N_1416,N_1015);
nor U1515 (N_1515,N_1079,N_1109);
nor U1516 (N_1516,N_1319,N_1123);
nor U1517 (N_1517,N_1019,N_1031);
nand U1518 (N_1518,N_1052,N_1067);
or U1519 (N_1519,N_1342,N_1376);
and U1520 (N_1520,N_1388,N_1130);
nand U1521 (N_1521,N_1364,N_1007);
and U1522 (N_1522,N_1049,N_1053);
nand U1523 (N_1523,N_1221,N_1111);
nand U1524 (N_1524,N_1144,N_1375);
or U1525 (N_1525,N_1258,N_1465);
xor U1526 (N_1526,N_1064,N_1443);
and U1527 (N_1527,N_1487,N_1418);
xor U1528 (N_1528,N_1061,N_1104);
and U1529 (N_1529,N_1114,N_1194);
xnor U1530 (N_1530,N_1297,N_1062);
nor U1531 (N_1531,N_1366,N_1432);
or U1532 (N_1532,N_1345,N_1320);
nand U1533 (N_1533,N_1129,N_1236);
or U1534 (N_1534,N_1338,N_1393);
nor U1535 (N_1535,N_1292,N_1076);
or U1536 (N_1536,N_1094,N_1153);
or U1537 (N_1537,N_1029,N_1060);
or U1538 (N_1538,N_1307,N_1211);
or U1539 (N_1539,N_1284,N_1014);
and U1540 (N_1540,N_1093,N_1037);
nand U1541 (N_1541,N_1038,N_1318);
xnor U1542 (N_1542,N_1026,N_1021);
or U1543 (N_1543,N_1113,N_1169);
nand U1544 (N_1544,N_1158,N_1477);
nor U1545 (N_1545,N_1492,N_1197);
xor U1546 (N_1546,N_1032,N_1483);
xor U1547 (N_1547,N_1448,N_1034);
and U1548 (N_1548,N_1261,N_1030);
nor U1549 (N_1549,N_1472,N_1473);
or U1550 (N_1550,N_1071,N_1354);
xnor U1551 (N_1551,N_1117,N_1102);
nand U1552 (N_1552,N_1103,N_1239);
or U1553 (N_1553,N_1488,N_1431);
xor U1554 (N_1554,N_1145,N_1410);
xor U1555 (N_1555,N_1108,N_1051);
nor U1556 (N_1556,N_1459,N_1274);
nor U1557 (N_1557,N_1229,N_1355);
nand U1558 (N_1558,N_1467,N_1137);
nor U1559 (N_1559,N_1122,N_1457);
xnor U1560 (N_1560,N_1240,N_1138);
and U1561 (N_1561,N_1496,N_1439);
nor U1562 (N_1562,N_1163,N_1142);
nor U1563 (N_1563,N_1460,N_1495);
nand U1564 (N_1564,N_1267,N_1497);
or U1565 (N_1565,N_1063,N_1119);
nand U1566 (N_1566,N_1486,N_1214);
and U1567 (N_1567,N_1012,N_1305);
xor U1568 (N_1568,N_1391,N_1367);
nor U1569 (N_1569,N_1105,N_1296);
and U1570 (N_1570,N_1161,N_1203);
nand U1571 (N_1571,N_1302,N_1313);
and U1572 (N_1572,N_1368,N_1110);
nor U1573 (N_1573,N_1127,N_1423);
nor U1574 (N_1574,N_1081,N_1125);
nand U1575 (N_1575,N_1441,N_1245);
or U1576 (N_1576,N_1310,N_1397);
xor U1577 (N_1577,N_1168,N_1200);
or U1578 (N_1578,N_1152,N_1133);
xnor U1579 (N_1579,N_1401,N_1281);
and U1580 (N_1580,N_1445,N_1215);
or U1581 (N_1581,N_1272,N_1396);
nand U1582 (N_1582,N_1248,N_1089);
or U1583 (N_1583,N_1263,N_1233);
xnor U1584 (N_1584,N_1303,N_1300);
nand U1585 (N_1585,N_1208,N_1069);
nand U1586 (N_1586,N_1121,N_1140);
or U1587 (N_1587,N_1413,N_1450);
or U1588 (N_1588,N_1097,N_1290);
and U1589 (N_1589,N_1086,N_1070);
nand U1590 (N_1590,N_1424,N_1382);
nand U1591 (N_1591,N_1430,N_1484);
or U1592 (N_1592,N_1332,N_1010);
and U1593 (N_1593,N_1143,N_1147);
or U1594 (N_1594,N_1124,N_1198);
xor U1595 (N_1595,N_1224,N_1165);
or U1596 (N_1596,N_1048,N_1417);
nor U1597 (N_1597,N_1427,N_1231);
xor U1598 (N_1598,N_1399,N_1253);
and U1599 (N_1599,N_1449,N_1392);
or U1600 (N_1600,N_1337,N_1403);
nor U1601 (N_1601,N_1335,N_1323);
and U1602 (N_1602,N_1400,N_1218);
nand U1603 (N_1603,N_1156,N_1271);
nor U1604 (N_1604,N_1451,N_1325);
and U1605 (N_1605,N_1379,N_1128);
and U1606 (N_1606,N_1442,N_1370);
nor U1607 (N_1607,N_1244,N_1475);
nor U1608 (N_1608,N_1250,N_1499);
nand U1609 (N_1609,N_1206,N_1286);
and U1610 (N_1610,N_1357,N_1005);
xnor U1611 (N_1611,N_1377,N_1404);
xor U1612 (N_1612,N_1273,N_1234);
and U1613 (N_1613,N_1359,N_1425);
nor U1614 (N_1614,N_1277,N_1016);
nand U1615 (N_1615,N_1433,N_1327);
nor U1616 (N_1616,N_1464,N_1287);
or U1617 (N_1617,N_1264,N_1216);
xor U1618 (N_1618,N_1289,N_1322);
or U1619 (N_1619,N_1098,N_1346);
nor U1620 (N_1620,N_1191,N_1176);
nor U1621 (N_1621,N_1440,N_1462);
nand U1622 (N_1622,N_1210,N_1013);
xor U1623 (N_1623,N_1184,N_1056);
nand U1624 (N_1624,N_1447,N_1057);
nand U1625 (N_1625,N_1150,N_1157);
nand U1626 (N_1626,N_1414,N_1304);
and U1627 (N_1627,N_1421,N_1468);
nor U1628 (N_1628,N_1050,N_1333);
nor U1629 (N_1629,N_1087,N_1330);
xnor U1630 (N_1630,N_1341,N_1285);
nor U1631 (N_1631,N_1306,N_1356);
nand U1632 (N_1632,N_1020,N_1480);
xnor U1633 (N_1633,N_1046,N_1172);
xnor U1634 (N_1634,N_1177,N_1275);
nor U1635 (N_1635,N_1136,N_1426);
nor U1636 (N_1636,N_1280,N_1259);
nand U1637 (N_1637,N_1227,N_1077);
nand U1638 (N_1638,N_1316,N_1249);
nor U1639 (N_1639,N_1419,N_1212);
xnor U1640 (N_1640,N_1242,N_1167);
and U1641 (N_1641,N_1456,N_1331);
or U1642 (N_1642,N_1471,N_1171);
and U1643 (N_1643,N_1420,N_1469);
nand U1644 (N_1644,N_1228,N_1294);
nor U1645 (N_1645,N_1225,N_1226);
or U1646 (N_1646,N_1001,N_1185);
xnor U1647 (N_1647,N_1084,N_1238);
nand U1648 (N_1648,N_1186,N_1075);
xnor U1649 (N_1649,N_1378,N_1118);
and U1650 (N_1650,N_1023,N_1344);
nor U1651 (N_1651,N_1395,N_1193);
or U1652 (N_1652,N_1195,N_1132);
or U1653 (N_1653,N_1315,N_1347);
nor U1654 (N_1654,N_1453,N_1134);
or U1655 (N_1655,N_1115,N_1078);
xor U1656 (N_1656,N_1452,N_1232);
and U1657 (N_1657,N_1348,N_1100);
and U1658 (N_1658,N_1213,N_1470);
and U1659 (N_1659,N_1033,N_1082);
or U1660 (N_1660,N_1055,N_1074);
xnor U1661 (N_1661,N_1498,N_1180);
and U1662 (N_1662,N_1326,N_1265);
xor U1663 (N_1663,N_1428,N_1170);
nor U1664 (N_1664,N_1446,N_1293);
and U1665 (N_1665,N_1199,N_1339);
and U1666 (N_1666,N_1025,N_1243);
and U1667 (N_1667,N_1083,N_1159);
or U1668 (N_1668,N_1408,N_1043);
or U1669 (N_1669,N_1278,N_1298);
xnor U1670 (N_1670,N_1383,N_1178);
or U1671 (N_1671,N_1187,N_1205);
and U1672 (N_1672,N_1476,N_1494);
nor U1673 (N_1673,N_1386,N_1350);
xor U1674 (N_1674,N_1112,N_1351);
and U1675 (N_1675,N_1369,N_1329);
nand U1676 (N_1676,N_1328,N_1358);
nor U1677 (N_1677,N_1308,N_1073);
and U1678 (N_1678,N_1444,N_1435);
nand U1679 (N_1679,N_1343,N_1493);
nand U1680 (N_1680,N_1235,N_1268);
nor U1681 (N_1681,N_1387,N_1256);
xnor U1682 (N_1682,N_1024,N_1044);
or U1683 (N_1683,N_1058,N_1255);
nor U1684 (N_1684,N_1035,N_1047);
and U1685 (N_1685,N_1204,N_1295);
nor U1686 (N_1686,N_1257,N_1092);
xnor U1687 (N_1687,N_1042,N_1402);
nor U1688 (N_1688,N_1381,N_1196);
and U1689 (N_1689,N_1415,N_1006);
nor U1690 (N_1690,N_1003,N_1155);
nor U1691 (N_1691,N_1027,N_1202);
or U1692 (N_1692,N_1088,N_1324);
and U1693 (N_1693,N_1352,N_1160);
nor U1694 (N_1694,N_1485,N_1085);
xor U1695 (N_1695,N_1317,N_1314);
and U1696 (N_1696,N_1131,N_1209);
xnor U1697 (N_1697,N_1361,N_1398);
nand U1698 (N_1698,N_1262,N_1201);
nor U1699 (N_1699,N_1162,N_1482);
xnor U1700 (N_1700,N_1059,N_1276);
or U1701 (N_1701,N_1028,N_1438);
and U1702 (N_1702,N_1309,N_1353);
xnor U1703 (N_1703,N_1481,N_1299);
and U1704 (N_1704,N_1154,N_1372);
nor U1705 (N_1705,N_1422,N_1096);
nand U1706 (N_1706,N_1436,N_1454);
and U1707 (N_1707,N_1252,N_1373);
nand U1708 (N_1708,N_1164,N_1279);
nand U1709 (N_1709,N_1054,N_1116);
and U1710 (N_1710,N_1072,N_1407);
nand U1711 (N_1711,N_1380,N_1463);
and U1712 (N_1712,N_1237,N_1011);
or U1713 (N_1713,N_1018,N_1340);
or U1714 (N_1714,N_1190,N_1223);
nand U1715 (N_1715,N_1288,N_1017);
and U1716 (N_1716,N_1384,N_1166);
and U1717 (N_1717,N_1068,N_1311);
or U1718 (N_1718,N_1254,N_1390);
nor U1719 (N_1719,N_1474,N_1090);
and U1720 (N_1720,N_1041,N_1283);
xor U1721 (N_1721,N_1065,N_1107);
nand U1722 (N_1722,N_1411,N_1000);
nand U1723 (N_1723,N_1349,N_1321);
nand U1724 (N_1724,N_1135,N_1270);
xnor U1725 (N_1725,N_1219,N_1004);
nor U1726 (N_1726,N_1412,N_1182);
or U1727 (N_1727,N_1247,N_1269);
or U1728 (N_1728,N_1466,N_1437);
or U1729 (N_1729,N_1009,N_1222);
xnor U1730 (N_1730,N_1101,N_1489);
nand U1731 (N_1731,N_1192,N_1217);
xor U1732 (N_1732,N_1139,N_1363);
nor U1733 (N_1733,N_1173,N_1066);
nand U1734 (N_1734,N_1406,N_1045);
or U1735 (N_1735,N_1022,N_1146);
nor U1736 (N_1736,N_1181,N_1106);
xnor U1737 (N_1737,N_1371,N_1126);
xnor U1738 (N_1738,N_1039,N_1461);
nand U1739 (N_1739,N_1490,N_1362);
or U1740 (N_1740,N_1183,N_1260);
nand U1741 (N_1741,N_1189,N_1179);
or U1742 (N_1742,N_1148,N_1230);
and U1743 (N_1743,N_1479,N_1151);
and U1744 (N_1744,N_1282,N_1141);
nand U1745 (N_1745,N_1409,N_1241);
xor U1746 (N_1746,N_1405,N_1120);
and U1747 (N_1747,N_1312,N_1491);
xor U1748 (N_1748,N_1246,N_1188);
xnor U1749 (N_1749,N_1099,N_1434);
xor U1750 (N_1750,N_1079,N_1359);
nand U1751 (N_1751,N_1305,N_1075);
or U1752 (N_1752,N_1115,N_1467);
or U1753 (N_1753,N_1228,N_1308);
nor U1754 (N_1754,N_1431,N_1225);
and U1755 (N_1755,N_1416,N_1456);
nand U1756 (N_1756,N_1217,N_1152);
nand U1757 (N_1757,N_1191,N_1209);
or U1758 (N_1758,N_1195,N_1459);
xor U1759 (N_1759,N_1444,N_1388);
or U1760 (N_1760,N_1391,N_1460);
and U1761 (N_1761,N_1227,N_1213);
xor U1762 (N_1762,N_1266,N_1390);
or U1763 (N_1763,N_1315,N_1008);
nand U1764 (N_1764,N_1472,N_1184);
nor U1765 (N_1765,N_1404,N_1315);
or U1766 (N_1766,N_1222,N_1226);
or U1767 (N_1767,N_1121,N_1110);
or U1768 (N_1768,N_1077,N_1332);
or U1769 (N_1769,N_1215,N_1024);
or U1770 (N_1770,N_1433,N_1346);
and U1771 (N_1771,N_1301,N_1489);
or U1772 (N_1772,N_1476,N_1391);
nor U1773 (N_1773,N_1238,N_1283);
xnor U1774 (N_1774,N_1234,N_1431);
xor U1775 (N_1775,N_1207,N_1427);
and U1776 (N_1776,N_1390,N_1158);
and U1777 (N_1777,N_1352,N_1400);
and U1778 (N_1778,N_1103,N_1006);
or U1779 (N_1779,N_1328,N_1392);
nand U1780 (N_1780,N_1268,N_1459);
nand U1781 (N_1781,N_1247,N_1094);
nand U1782 (N_1782,N_1283,N_1476);
nand U1783 (N_1783,N_1162,N_1265);
nor U1784 (N_1784,N_1415,N_1324);
and U1785 (N_1785,N_1255,N_1370);
nor U1786 (N_1786,N_1429,N_1432);
and U1787 (N_1787,N_1460,N_1349);
nand U1788 (N_1788,N_1189,N_1305);
or U1789 (N_1789,N_1030,N_1374);
xnor U1790 (N_1790,N_1175,N_1121);
nor U1791 (N_1791,N_1066,N_1091);
nor U1792 (N_1792,N_1039,N_1053);
nor U1793 (N_1793,N_1430,N_1341);
nand U1794 (N_1794,N_1209,N_1223);
and U1795 (N_1795,N_1309,N_1403);
and U1796 (N_1796,N_1382,N_1125);
and U1797 (N_1797,N_1086,N_1367);
or U1798 (N_1798,N_1242,N_1357);
xnor U1799 (N_1799,N_1279,N_1446);
and U1800 (N_1800,N_1298,N_1095);
or U1801 (N_1801,N_1441,N_1093);
and U1802 (N_1802,N_1311,N_1440);
xor U1803 (N_1803,N_1212,N_1420);
xor U1804 (N_1804,N_1014,N_1040);
and U1805 (N_1805,N_1136,N_1184);
nand U1806 (N_1806,N_1330,N_1436);
xor U1807 (N_1807,N_1236,N_1246);
nor U1808 (N_1808,N_1149,N_1362);
and U1809 (N_1809,N_1094,N_1465);
xnor U1810 (N_1810,N_1145,N_1310);
or U1811 (N_1811,N_1091,N_1397);
nand U1812 (N_1812,N_1387,N_1498);
or U1813 (N_1813,N_1495,N_1030);
nor U1814 (N_1814,N_1094,N_1193);
and U1815 (N_1815,N_1258,N_1206);
nor U1816 (N_1816,N_1352,N_1122);
and U1817 (N_1817,N_1119,N_1490);
or U1818 (N_1818,N_1250,N_1082);
nor U1819 (N_1819,N_1047,N_1124);
and U1820 (N_1820,N_1086,N_1182);
xnor U1821 (N_1821,N_1268,N_1065);
xor U1822 (N_1822,N_1194,N_1437);
or U1823 (N_1823,N_1485,N_1049);
and U1824 (N_1824,N_1041,N_1441);
and U1825 (N_1825,N_1278,N_1071);
or U1826 (N_1826,N_1185,N_1245);
and U1827 (N_1827,N_1317,N_1307);
or U1828 (N_1828,N_1172,N_1419);
xnor U1829 (N_1829,N_1197,N_1337);
or U1830 (N_1830,N_1245,N_1222);
and U1831 (N_1831,N_1264,N_1225);
nand U1832 (N_1832,N_1154,N_1428);
and U1833 (N_1833,N_1160,N_1458);
xor U1834 (N_1834,N_1072,N_1155);
xor U1835 (N_1835,N_1361,N_1299);
nand U1836 (N_1836,N_1309,N_1168);
or U1837 (N_1837,N_1173,N_1196);
or U1838 (N_1838,N_1407,N_1123);
nand U1839 (N_1839,N_1446,N_1233);
nor U1840 (N_1840,N_1090,N_1421);
nand U1841 (N_1841,N_1253,N_1282);
and U1842 (N_1842,N_1056,N_1499);
and U1843 (N_1843,N_1049,N_1055);
and U1844 (N_1844,N_1346,N_1267);
or U1845 (N_1845,N_1154,N_1342);
and U1846 (N_1846,N_1481,N_1074);
xor U1847 (N_1847,N_1362,N_1022);
nor U1848 (N_1848,N_1432,N_1208);
nor U1849 (N_1849,N_1343,N_1263);
nand U1850 (N_1850,N_1055,N_1410);
xnor U1851 (N_1851,N_1295,N_1146);
xor U1852 (N_1852,N_1468,N_1242);
xnor U1853 (N_1853,N_1256,N_1329);
nand U1854 (N_1854,N_1089,N_1311);
nand U1855 (N_1855,N_1223,N_1325);
nand U1856 (N_1856,N_1119,N_1018);
xor U1857 (N_1857,N_1423,N_1188);
nand U1858 (N_1858,N_1477,N_1399);
or U1859 (N_1859,N_1189,N_1002);
or U1860 (N_1860,N_1002,N_1339);
xor U1861 (N_1861,N_1195,N_1069);
and U1862 (N_1862,N_1220,N_1073);
or U1863 (N_1863,N_1213,N_1059);
nand U1864 (N_1864,N_1386,N_1298);
or U1865 (N_1865,N_1111,N_1173);
nand U1866 (N_1866,N_1045,N_1197);
nand U1867 (N_1867,N_1023,N_1405);
nor U1868 (N_1868,N_1466,N_1142);
nand U1869 (N_1869,N_1232,N_1337);
nand U1870 (N_1870,N_1203,N_1069);
and U1871 (N_1871,N_1149,N_1484);
xor U1872 (N_1872,N_1472,N_1115);
and U1873 (N_1873,N_1221,N_1250);
nor U1874 (N_1874,N_1195,N_1004);
nor U1875 (N_1875,N_1382,N_1117);
and U1876 (N_1876,N_1233,N_1161);
or U1877 (N_1877,N_1443,N_1125);
xor U1878 (N_1878,N_1025,N_1296);
nor U1879 (N_1879,N_1449,N_1404);
and U1880 (N_1880,N_1437,N_1088);
nor U1881 (N_1881,N_1280,N_1343);
xor U1882 (N_1882,N_1196,N_1436);
xor U1883 (N_1883,N_1002,N_1471);
nand U1884 (N_1884,N_1481,N_1043);
or U1885 (N_1885,N_1068,N_1057);
and U1886 (N_1886,N_1484,N_1458);
and U1887 (N_1887,N_1015,N_1183);
nand U1888 (N_1888,N_1467,N_1422);
or U1889 (N_1889,N_1155,N_1173);
nor U1890 (N_1890,N_1400,N_1297);
nor U1891 (N_1891,N_1392,N_1111);
and U1892 (N_1892,N_1141,N_1006);
xnor U1893 (N_1893,N_1077,N_1295);
nor U1894 (N_1894,N_1127,N_1483);
xor U1895 (N_1895,N_1173,N_1363);
or U1896 (N_1896,N_1385,N_1327);
xor U1897 (N_1897,N_1461,N_1208);
and U1898 (N_1898,N_1016,N_1240);
or U1899 (N_1899,N_1321,N_1365);
nand U1900 (N_1900,N_1191,N_1069);
xor U1901 (N_1901,N_1157,N_1164);
nand U1902 (N_1902,N_1450,N_1185);
nor U1903 (N_1903,N_1294,N_1400);
nor U1904 (N_1904,N_1177,N_1216);
and U1905 (N_1905,N_1470,N_1252);
nor U1906 (N_1906,N_1115,N_1206);
and U1907 (N_1907,N_1274,N_1416);
nor U1908 (N_1908,N_1295,N_1309);
nand U1909 (N_1909,N_1222,N_1215);
or U1910 (N_1910,N_1212,N_1375);
and U1911 (N_1911,N_1348,N_1419);
nand U1912 (N_1912,N_1010,N_1443);
nand U1913 (N_1913,N_1216,N_1085);
or U1914 (N_1914,N_1350,N_1048);
nor U1915 (N_1915,N_1301,N_1207);
or U1916 (N_1916,N_1171,N_1251);
xnor U1917 (N_1917,N_1355,N_1066);
nand U1918 (N_1918,N_1234,N_1371);
nand U1919 (N_1919,N_1238,N_1479);
nor U1920 (N_1920,N_1279,N_1402);
xnor U1921 (N_1921,N_1260,N_1028);
nor U1922 (N_1922,N_1079,N_1093);
nor U1923 (N_1923,N_1252,N_1270);
xnor U1924 (N_1924,N_1050,N_1083);
and U1925 (N_1925,N_1169,N_1402);
and U1926 (N_1926,N_1459,N_1446);
nor U1927 (N_1927,N_1069,N_1123);
or U1928 (N_1928,N_1206,N_1013);
nand U1929 (N_1929,N_1485,N_1069);
or U1930 (N_1930,N_1361,N_1336);
nor U1931 (N_1931,N_1034,N_1357);
or U1932 (N_1932,N_1333,N_1049);
or U1933 (N_1933,N_1308,N_1295);
nor U1934 (N_1934,N_1393,N_1498);
or U1935 (N_1935,N_1360,N_1076);
and U1936 (N_1936,N_1120,N_1493);
or U1937 (N_1937,N_1484,N_1034);
and U1938 (N_1938,N_1263,N_1058);
xnor U1939 (N_1939,N_1011,N_1417);
and U1940 (N_1940,N_1443,N_1075);
nor U1941 (N_1941,N_1347,N_1367);
and U1942 (N_1942,N_1304,N_1349);
nor U1943 (N_1943,N_1224,N_1476);
or U1944 (N_1944,N_1263,N_1497);
nor U1945 (N_1945,N_1057,N_1406);
or U1946 (N_1946,N_1495,N_1079);
nor U1947 (N_1947,N_1276,N_1302);
nand U1948 (N_1948,N_1465,N_1480);
xor U1949 (N_1949,N_1081,N_1261);
nor U1950 (N_1950,N_1400,N_1125);
nand U1951 (N_1951,N_1416,N_1421);
xor U1952 (N_1952,N_1126,N_1009);
and U1953 (N_1953,N_1069,N_1310);
or U1954 (N_1954,N_1302,N_1223);
or U1955 (N_1955,N_1369,N_1335);
and U1956 (N_1956,N_1099,N_1012);
nand U1957 (N_1957,N_1289,N_1259);
and U1958 (N_1958,N_1255,N_1232);
xnor U1959 (N_1959,N_1088,N_1020);
or U1960 (N_1960,N_1202,N_1087);
or U1961 (N_1961,N_1006,N_1199);
xnor U1962 (N_1962,N_1071,N_1038);
xnor U1963 (N_1963,N_1117,N_1105);
nand U1964 (N_1964,N_1188,N_1249);
nor U1965 (N_1965,N_1051,N_1159);
nor U1966 (N_1966,N_1042,N_1006);
or U1967 (N_1967,N_1126,N_1342);
or U1968 (N_1968,N_1203,N_1301);
nor U1969 (N_1969,N_1014,N_1335);
or U1970 (N_1970,N_1439,N_1306);
nor U1971 (N_1971,N_1055,N_1285);
nor U1972 (N_1972,N_1206,N_1423);
nor U1973 (N_1973,N_1018,N_1495);
xor U1974 (N_1974,N_1224,N_1283);
nand U1975 (N_1975,N_1183,N_1410);
and U1976 (N_1976,N_1297,N_1177);
and U1977 (N_1977,N_1023,N_1138);
or U1978 (N_1978,N_1301,N_1484);
and U1979 (N_1979,N_1372,N_1216);
and U1980 (N_1980,N_1492,N_1030);
or U1981 (N_1981,N_1140,N_1125);
nor U1982 (N_1982,N_1302,N_1357);
nand U1983 (N_1983,N_1171,N_1001);
xor U1984 (N_1984,N_1295,N_1461);
or U1985 (N_1985,N_1284,N_1422);
xor U1986 (N_1986,N_1298,N_1494);
and U1987 (N_1987,N_1305,N_1009);
and U1988 (N_1988,N_1345,N_1051);
nand U1989 (N_1989,N_1370,N_1041);
and U1990 (N_1990,N_1467,N_1244);
nand U1991 (N_1991,N_1355,N_1081);
nand U1992 (N_1992,N_1480,N_1139);
xor U1993 (N_1993,N_1293,N_1432);
nand U1994 (N_1994,N_1107,N_1177);
and U1995 (N_1995,N_1234,N_1445);
nand U1996 (N_1996,N_1368,N_1166);
and U1997 (N_1997,N_1409,N_1054);
or U1998 (N_1998,N_1278,N_1040);
and U1999 (N_1999,N_1449,N_1356);
and U2000 (N_2000,N_1704,N_1503);
xor U2001 (N_2001,N_1521,N_1911);
nand U2002 (N_2002,N_1799,N_1548);
or U2003 (N_2003,N_1507,N_1765);
xnor U2004 (N_2004,N_1692,N_1876);
nor U2005 (N_2005,N_1868,N_1897);
nor U2006 (N_2006,N_1536,N_1739);
or U2007 (N_2007,N_1798,N_1590);
nor U2008 (N_2008,N_1557,N_1509);
nand U2009 (N_2009,N_1754,N_1671);
nand U2010 (N_2010,N_1937,N_1885);
nand U2011 (N_2011,N_1629,N_1500);
xor U2012 (N_2012,N_1510,N_1670);
xor U2013 (N_2013,N_1601,N_1830);
xor U2014 (N_2014,N_1811,N_1931);
xor U2015 (N_2015,N_1686,N_1533);
nor U2016 (N_2016,N_1817,N_1818);
nand U2017 (N_2017,N_1839,N_1961);
nand U2018 (N_2018,N_1709,N_1947);
or U2019 (N_2019,N_1644,N_1814);
nor U2020 (N_2020,N_1723,N_1816);
nor U2021 (N_2021,N_1679,N_1565);
xor U2022 (N_2022,N_1726,N_1537);
nor U2023 (N_2023,N_1838,N_1792);
or U2024 (N_2024,N_1829,N_1942);
or U2025 (N_2025,N_1770,N_1802);
and U2026 (N_2026,N_1621,N_1908);
nand U2027 (N_2027,N_1635,N_1619);
xor U2028 (N_2028,N_1851,N_1895);
or U2029 (N_2029,N_1553,N_1694);
or U2030 (N_2030,N_1740,N_1820);
nor U2031 (N_2031,N_1691,N_1615);
nand U2032 (N_2032,N_1984,N_1512);
nand U2033 (N_2033,N_1840,N_1714);
or U2034 (N_2034,N_1748,N_1648);
xor U2035 (N_2035,N_1989,N_1866);
or U2036 (N_2036,N_1620,N_1513);
or U2037 (N_2037,N_1877,N_1583);
nor U2038 (N_2038,N_1586,N_1742);
nor U2039 (N_2039,N_1801,N_1878);
nor U2040 (N_2040,N_1935,N_1999);
nand U2041 (N_2041,N_1633,N_1940);
or U2042 (N_2042,N_1766,N_1954);
or U2043 (N_2043,N_1734,N_1511);
nand U2044 (N_2044,N_1584,N_1891);
xor U2045 (N_2045,N_1501,N_1985);
and U2046 (N_2046,N_1813,N_1927);
nor U2047 (N_2047,N_1899,N_1592);
nand U2048 (N_2048,N_1920,N_1921);
nand U2049 (N_2049,N_1736,N_1699);
nor U2050 (N_2050,N_1857,N_1753);
or U2051 (N_2051,N_1828,N_1969);
and U2052 (N_2052,N_1737,N_1782);
nor U2053 (N_2053,N_1749,N_1566);
nand U2054 (N_2054,N_1731,N_1534);
nand U2055 (N_2055,N_1647,N_1567);
xnor U2056 (N_2056,N_1756,N_1861);
nand U2057 (N_2057,N_1881,N_1707);
or U2058 (N_2058,N_1977,N_1953);
and U2059 (N_2059,N_1658,N_1973);
nand U2060 (N_2060,N_1535,N_1902);
nor U2061 (N_2061,N_1576,N_1915);
and U2062 (N_2062,N_1549,N_1649);
xor U2063 (N_2063,N_1667,N_1729);
nor U2064 (N_2064,N_1762,N_1972);
and U2065 (N_2065,N_1545,N_1626);
xnor U2066 (N_2066,N_1571,N_1672);
nor U2067 (N_2067,N_1594,N_1531);
and U2068 (N_2068,N_1847,N_1903);
and U2069 (N_2069,N_1913,N_1676);
nor U2070 (N_2070,N_1755,N_1646);
and U2071 (N_2071,N_1611,N_1775);
xnor U2072 (N_2072,N_1668,N_1900);
or U2073 (N_2073,N_1779,N_1751);
xor U2074 (N_2074,N_1730,N_1684);
nand U2075 (N_2075,N_1957,N_1759);
nor U2076 (N_2076,N_1997,N_1522);
nand U2077 (N_2077,N_1515,N_1570);
nand U2078 (N_2078,N_1653,N_1735);
or U2079 (N_2079,N_1794,N_1603);
nand U2080 (N_2080,N_1541,N_1781);
xnor U2081 (N_2081,N_1941,N_1763);
xor U2082 (N_2082,N_1708,N_1883);
nand U2083 (N_2083,N_1832,N_1701);
or U2084 (N_2084,N_1559,N_1527);
nand U2085 (N_2085,N_1666,N_1979);
and U2086 (N_2086,N_1597,N_1821);
or U2087 (N_2087,N_1805,N_1882);
xor U2088 (N_2088,N_1767,N_1656);
xnor U2089 (N_2089,N_1909,N_1693);
nand U2090 (N_2090,N_1724,N_1823);
or U2091 (N_2091,N_1623,N_1809);
or U2092 (N_2092,N_1831,N_1773);
and U2093 (N_2093,N_1544,N_1627);
and U2094 (N_2094,N_1853,N_1848);
and U2095 (N_2095,N_1894,N_1540);
or U2096 (N_2096,N_1638,N_1508);
nand U2097 (N_2097,N_1788,N_1791);
nand U2098 (N_2098,N_1778,N_1988);
nand U2099 (N_2099,N_1886,N_1945);
and U2100 (N_2100,N_1804,N_1543);
and U2101 (N_2101,N_1800,N_1980);
xor U2102 (N_2102,N_1514,N_1844);
and U2103 (N_2103,N_1573,N_1850);
nand U2104 (N_2104,N_1574,N_1971);
or U2105 (N_2105,N_1747,N_1991);
nor U2106 (N_2106,N_1661,N_1519);
xor U2107 (N_2107,N_1625,N_1806);
nor U2108 (N_2108,N_1695,N_1604);
nor U2109 (N_2109,N_1854,N_1569);
or U2110 (N_2110,N_1563,N_1674);
and U2111 (N_2111,N_1650,N_1624);
nand U2112 (N_2112,N_1958,N_1986);
xnor U2113 (N_2113,N_1516,N_1618);
nand U2114 (N_2114,N_1572,N_1777);
or U2115 (N_2115,N_1710,N_1595);
xnor U2116 (N_2116,N_1562,N_1612);
or U2117 (N_2117,N_1696,N_1657);
nand U2118 (N_2118,N_1803,N_1933);
nor U2119 (N_2119,N_1700,N_1640);
nor U2120 (N_2120,N_1764,N_1869);
or U2121 (N_2121,N_1705,N_1506);
nand U2122 (N_2122,N_1702,N_1795);
and U2123 (N_2123,N_1682,N_1889);
or U2124 (N_2124,N_1607,N_1606);
and U2125 (N_2125,N_1930,N_1532);
nand U2126 (N_2126,N_1807,N_1884);
xnor U2127 (N_2127,N_1630,N_1873);
and U2128 (N_2128,N_1936,N_1774);
nand U2129 (N_2129,N_1581,N_1698);
xor U2130 (N_2130,N_1962,N_1966);
nor U2131 (N_2131,N_1722,N_1987);
or U2132 (N_2132,N_1636,N_1556);
xor U2133 (N_2133,N_1520,N_1956);
and U2134 (N_2134,N_1968,N_1706);
nand U2135 (N_2135,N_1918,N_1579);
nand U2136 (N_2136,N_1598,N_1622);
nand U2137 (N_2137,N_1716,N_1560);
and U2138 (N_2138,N_1750,N_1810);
and U2139 (N_2139,N_1896,N_1925);
nand U2140 (N_2140,N_1978,N_1951);
nor U2141 (N_2141,N_1796,N_1906);
nor U2142 (N_2142,N_1659,N_1772);
and U2143 (N_2143,N_1959,N_1518);
nand U2144 (N_2144,N_1654,N_1554);
nand U2145 (N_2145,N_1812,N_1744);
or U2146 (N_2146,N_1599,N_1950);
xnor U2147 (N_2147,N_1645,N_1718);
nor U2148 (N_2148,N_1605,N_1655);
nand U2149 (N_2149,N_1863,N_1790);
and U2150 (N_2150,N_1719,N_1610);
or U2151 (N_2151,N_1926,N_1639);
nor U2152 (N_2152,N_1824,N_1517);
and U2153 (N_2153,N_1711,N_1689);
nor U2154 (N_2154,N_1939,N_1907);
nand U2155 (N_2155,N_1524,N_1964);
and U2156 (N_2156,N_1944,N_1929);
nand U2157 (N_2157,N_1628,N_1901);
and U2158 (N_2158,N_1525,N_1547);
xor U2159 (N_2159,N_1786,N_1660);
xnor U2160 (N_2160,N_1688,N_1928);
nand U2161 (N_2161,N_1609,N_1827);
or U2162 (N_2162,N_1793,N_1943);
nand U2163 (N_2163,N_1600,N_1994);
and U2164 (N_2164,N_1585,N_1712);
xor U2165 (N_2165,N_1643,N_1996);
xor U2166 (N_2166,N_1602,N_1697);
and U2167 (N_2167,N_1552,N_1780);
xnor U2168 (N_2168,N_1502,N_1880);
xnor U2169 (N_2169,N_1564,N_1917);
nor U2170 (N_2170,N_1856,N_1651);
nand U2171 (N_2171,N_1613,N_1787);
nor U2172 (N_2172,N_1616,N_1992);
nor U2173 (N_2173,N_1725,N_1975);
xor U2174 (N_2174,N_1924,N_1995);
xor U2175 (N_2175,N_1990,N_1952);
and U2176 (N_2176,N_1631,N_1677);
or U2177 (N_2177,N_1761,N_1703);
or U2178 (N_2178,N_1596,N_1741);
nor U2179 (N_2179,N_1642,N_1577);
and U2180 (N_2180,N_1825,N_1871);
nand U2181 (N_2181,N_1858,N_1842);
xor U2182 (N_2182,N_1912,N_1752);
nand U2183 (N_2183,N_1808,N_1558);
xor U2184 (N_2184,N_1922,N_1919);
and U2185 (N_2185,N_1837,N_1874);
nand U2186 (N_2186,N_1846,N_1591);
nand U2187 (N_2187,N_1529,N_1617);
and U2188 (N_2188,N_1539,N_1946);
nand U2189 (N_2189,N_1923,N_1784);
and U2190 (N_2190,N_1732,N_1965);
nor U2191 (N_2191,N_1538,N_1758);
or U2192 (N_2192,N_1713,N_1687);
xor U2193 (N_2193,N_1561,N_1998);
nand U2194 (N_2194,N_1578,N_1963);
nand U2195 (N_2195,N_1664,N_1681);
nor U2196 (N_2196,N_1738,N_1743);
and U2197 (N_2197,N_1862,N_1879);
xnor U2198 (N_2198,N_1916,N_1855);
or U2199 (N_2199,N_1551,N_1673);
nand U2200 (N_2200,N_1892,N_1637);
or U2201 (N_2201,N_1721,N_1678);
xor U2202 (N_2202,N_1720,N_1665);
xnor U2203 (N_2203,N_1860,N_1608);
or U2204 (N_2204,N_1938,N_1970);
or U2205 (N_2205,N_1690,N_1680);
nand U2206 (N_2206,N_1523,N_1632);
or U2207 (N_2207,N_1776,N_1768);
nor U2208 (N_2208,N_1949,N_1955);
nor U2209 (N_2209,N_1893,N_1905);
or U2210 (N_2210,N_1822,N_1715);
nand U2211 (N_2211,N_1663,N_1981);
xnor U2212 (N_2212,N_1717,N_1634);
or U2213 (N_2213,N_1542,N_1614);
xor U2214 (N_2214,N_1550,N_1641);
or U2215 (N_2215,N_1826,N_1888);
and U2216 (N_2216,N_1890,N_1833);
and U2217 (N_2217,N_1783,N_1575);
nor U2218 (N_2218,N_1867,N_1745);
nor U2219 (N_2219,N_1669,N_1675);
and U2220 (N_2220,N_1746,N_1593);
and U2221 (N_2221,N_1652,N_1834);
or U2222 (N_2222,N_1662,N_1815);
xnor U2223 (N_2223,N_1904,N_1789);
nor U2224 (N_2224,N_1967,N_1797);
or U2225 (N_2225,N_1769,N_1836);
nand U2226 (N_2226,N_1843,N_1504);
nor U2227 (N_2227,N_1760,N_1568);
xor U2228 (N_2228,N_1898,N_1887);
nand U2229 (N_2229,N_1910,N_1932);
xor U2230 (N_2230,N_1555,N_1771);
or U2231 (N_2231,N_1526,N_1875);
nor U2232 (N_2232,N_1580,N_1872);
nand U2233 (N_2233,N_1859,N_1835);
or U2234 (N_2234,N_1841,N_1948);
and U2235 (N_2235,N_1870,N_1728);
or U2236 (N_2236,N_1976,N_1864);
xor U2237 (N_2237,N_1785,N_1505);
nor U2238 (N_2238,N_1589,N_1528);
and U2239 (N_2239,N_1819,N_1960);
and U2240 (N_2240,N_1849,N_1530);
or U2241 (N_2241,N_1588,N_1983);
and U2242 (N_2242,N_1727,N_1546);
or U2243 (N_2243,N_1865,N_1685);
or U2244 (N_2244,N_1993,N_1845);
and U2245 (N_2245,N_1587,N_1934);
or U2246 (N_2246,N_1982,N_1582);
nor U2247 (N_2247,N_1974,N_1683);
xor U2248 (N_2248,N_1914,N_1852);
or U2249 (N_2249,N_1757,N_1733);
and U2250 (N_2250,N_1981,N_1650);
or U2251 (N_2251,N_1972,N_1546);
and U2252 (N_2252,N_1837,N_1595);
xor U2253 (N_2253,N_1923,N_1919);
or U2254 (N_2254,N_1575,N_1881);
nand U2255 (N_2255,N_1664,N_1790);
and U2256 (N_2256,N_1556,N_1517);
xor U2257 (N_2257,N_1915,N_1715);
or U2258 (N_2258,N_1554,N_1761);
nor U2259 (N_2259,N_1759,N_1536);
nand U2260 (N_2260,N_1634,N_1902);
or U2261 (N_2261,N_1595,N_1836);
nor U2262 (N_2262,N_1667,N_1821);
nor U2263 (N_2263,N_1825,N_1958);
xnor U2264 (N_2264,N_1788,N_1723);
and U2265 (N_2265,N_1781,N_1754);
or U2266 (N_2266,N_1571,N_1560);
nand U2267 (N_2267,N_1960,N_1715);
xnor U2268 (N_2268,N_1884,N_1935);
xnor U2269 (N_2269,N_1799,N_1521);
nand U2270 (N_2270,N_1530,N_1522);
nand U2271 (N_2271,N_1566,N_1773);
xnor U2272 (N_2272,N_1675,N_1865);
and U2273 (N_2273,N_1875,N_1601);
xor U2274 (N_2274,N_1526,N_1653);
nor U2275 (N_2275,N_1858,N_1872);
nor U2276 (N_2276,N_1951,N_1790);
xnor U2277 (N_2277,N_1682,N_1548);
nor U2278 (N_2278,N_1934,N_1645);
nor U2279 (N_2279,N_1901,N_1847);
nand U2280 (N_2280,N_1842,N_1591);
nand U2281 (N_2281,N_1566,N_1644);
nor U2282 (N_2282,N_1893,N_1650);
or U2283 (N_2283,N_1970,N_1869);
nor U2284 (N_2284,N_1734,N_1704);
nand U2285 (N_2285,N_1566,N_1690);
nand U2286 (N_2286,N_1621,N_1519);
nor U2287 (N_2287,N_1542,N_1670);
xnor U2288 (N_2288,N_1845,N_1754);
xor U2289 (N_2289,N_1539,N_1963);
xor U2290 (N_2290,N_1997,N_1573);
xnor U2291 (N_2291,N_1998,N_1728);
and U2292 (N_2292,N_1576,N_1886);
nor U2293 (N_2293,N_1525,N_1915);
nor U2294 (N_2294,N_1830,N_1849);
nor U2295 (N_2295,N_1983,N_1814);
or U2296 (N_2296,N_1654,N_1902);
xnor U2297 (N_2297,N_1763,N_1935);
nor U2298 (N_2298,N_1547,N_1728);
or U2299 (N_2299,N_1611,N_1771);
nand U2300 (N_2300,N_1736,N_1845);
nor U2301 (N_2301,N_1597,N_1886);
xnor U2302 (N_2302,N_1694,N_1979);
nand U2303 (N_2303,N_1693,N_1628);
and U2304 (N_2304,N_1740,N_1574);
xnor U2305 (N_2305,N_1928,N_1656);
nor U2306 (N_2306,N_1853,N_1988);
or U2307 (N_2307,N_1792,N_1668);
and U2308 (N_2308,N_1533,N_1593);
and U2309 (N_2309,N_1510,N_1636);
nand U2310 (N_2310,N_1594,N_1883);
nor U2311 (N_2311,N_1585,N_1539);
nor U2312 (N_2312,N_1526,N_1854);
nor U2313 (N_2313,N_1693,N_1832);
nor U2314 (N_2314,N_1815,N_1989);
xor U2315 (N_2315,N_1710,N_1937);
xor U2316 (N_2316,N_1962,N_1576);
nand U2317 (N_2317,N_1807,N_1574);
or U2318 (N_2318,N_1989,N_1669);
nor U2319 (N_2319,N_1558,N_1935);
nand U2320 (N_2320,N_1615,N_1906);
and U2321 (N_2321,N_1524,N_1699);
or U2322 (N_2322,N_1586,N_1681);
nand U2323 (N_2323,N_1917,N_1756);
nor U2324 (N_2324,N_1733,N_1779);
nand U2325 (N_2325,N_1533,N_1530);
and U2326 (N_2326,N_1927,N_1791);
and U2327 (N_2327,N_1771,N_1644);
xnor U2328 (N_2328,N_1523,N_1904);
nand U2329 (N_2329,N_1583,N_1887);
xnor U2330 (N_2330,N_1554,N_1590);
or U2331 (N_2331,N_1811,N_1701);
nor U2332 (N_2332,N_1501,N_1792);
xor U2333 (N_2333,N_1983,N_1548);
nor U2334 (N_2334,N_1590,N_1537);
nand U2335 (N_2335,N_1833,N_1883);
xnor U2336 (N_2336,N_1641,N_1536);
xor U2337 (N_2337,N_1815,N_1723);
nor U2338 (N_2338,N_1862,N_1624);
xnor U2339 (N_2339,N_1601,N_1692);
and U2340 (N_2340,N_1909,N_1542);
nor U2341 (N_2341,N_1852,N_1988);
nand U2342 (N_2342,N_1764,N_1914);
nand U2343 (N_2343,N_1791,N_1549);
and U2344 (N_2344,N_1773,N_1814);
nor U2345 (N_2345,N_1819,N_1694);
or U2346 (N_2346,N_1654,N_1508);
nor U2347 (N_2347,N_1542,N_1506);
nor U2348 (N_2348,N_1640,N_1936);
nand U2349 (N_2349,N_1952,N_1636);
and U2350 (N_2350,N_1816,N_1832);
nand U2351 (N_2351,N_1656,N_1601);
or U2352 (N_2352,N_1502,N_1860);
nor U2353 (N_2353,N_1629,N_1924);
and U2354 (N_2354,N_1907,N_1501);
nand U2355 (N_2355,N_1868,N_1655);
and U2356 (N_2356,N_1933,N_1761);
nand U2357 (N_2357,N_1577,N_1787);
or U2358 (N_2358,N_1923,N_1615);
and U2359 (N_2359,N_1700,N_1997);
or U2360 (N_2360,N_1982,N_1554);
or U2361 (N_2361,N_1594,N_1540);
or U2362 (N_2362,N_1673,N_1820);
or U2363 (N_2363,N_1985,N_1571);
nand U2364 (N_2364,N_1967,N_1923);
xor U2365 (N_2365,N_1550,N_1837);
and U2366 (N_2366,N_1979,N_1761);
and U2367 (N_2367,N_1886,N_1677);
xnor U2368 (N_2368,N_1858,N_1773);
nor U2369 (N_2369,N_1707,N_1937);
or U2370 (N_2370,N_1509,N_1560);
xor U2371 (N_2371,N_1967,N_1871);
nand U2372 (N_2372,N_1631,N_1619);
xor U2373 (N_2373,N_1664,N_1876);
nand U2374 (N_2374,N_1736,N_1719);
nand U2375 (N_2375,N_1594,N_1662);
and U2376 (N_2376,N_1853,N_1742);
and U2377 (N_2377,N_1663,N_1580);
xnor U2378 (N_2378,N_1922,N_1681);
and U2379 (N_2379,N_1620,N_1940);
and U2380 (N_2380,N_1631,N_1607);
or U2381 (N_2381,N_1879,N_1913);
nor U2382 (N_2382,N_1777,N_1662);
xnor U2383 (N_2383,N_1676,N_1816);
nor U2384 (N_2384,N_1863,N_1869);
nand U2385 (N_2385,N_1973,N_1708);
xor U2386 (N_2386,N_1830,N_1574);
and U2387 (N_2387,N_1774,N_1867);
xor U2388 (N_2388,N_1515,N_1636);
nor U2389 (N_2389,N_1759,N_1850);
or U2390 (N_2390,N_1687,N_1820);
nor U2391 (N_2391,N_1704,N_1582);
or U2392 (N_2392,N_1639,N_1697);
xnor U2393 (N_2393,N_1756,N_1918);
xor U2394 (N_2394,N_1506,N_1693);
or U2395 (N_2395,N_1858,N_1793);
and U2396 (N_2396,N_1799,N_1969);
or U2397 (N_2397,N_1514,N_1871);
and U2398 (N_2398,N_1849,N_1641);
nor U2399 (N_2399,N_1688,N_1654);
or U2400 (N_2400,N_1721,N_1707);
or U2401 (N_2401,N_1948,N_1876);
nor U2402 (N_2402,N_1538,N_1620);
or U2403 (N_2403,N_1637,N_1766);
or U2404 (N_2404,N_1837,N_1711);
or U2405 (N_2405,N_1633,N_1763);
xnor U2406 (N_2406,N_1926,N_1649);
and U2407 (N_2407,N_1948,N_1609);
xor U2408 (N_2408,N_1978,N_1571);
nand U2409 (N_2409,N_1819,N_1522);
and U2410 (N_2410,N_1579,N_1689);
nor U2411 (N_2411,N_1793,N_1884);
xnor U2412 (N_2412,N_1545,N_1973);
or U2413 (N_2413,N_1736,N_1952);
and U2414 (N_2414,N_1973,N_1569);
xor U2415 (N_2415,N_1831,N_1563);
xnor U2416 (N_2416,N_1783,N_1721);
nor U2417 (N_2417,N_1708,N_1831);
xnor U2418 (N_2418,N_1751,N_1715);
or U2419 (N_2419,N_1946,N_1624);
or U2420 (N_2420,N_1689,N_1774);
and U2421 (N_2421,N_1660,N_1753);
nor U2422 (N_2422,N_1814,N_1529);
nor U2423 (N_2423,N_1734,N_1776);
xor U2424 (N_2424,N_1863,N_1662);
nand U2425 (N_2425,N_1965,N_1651);
nor U2426 (N_2426,N_1549,N_1775);
xor U2427 (N_2427,N_1732,N_1630);
nor U2428 (N_2428,N_1554,N_1879);
nand U2429 (N_2429,N_1762,N_1605);
and U2430 (N_2430,N_1580,N_1554);
or U2431 (N_2431,N_1691,N_1663);
nor U2432 (N_2432,N_1976,N_1986);
and U2433 (N_2433,N_1755,N_1670);
nand U2434 (N_2434,N_1809,N_1830);
nand U2435 (N_2435,N_1907,N_1620);
nor U2436 (N_2436,N_1733,N_1537);
xnor U2437 (N_2437,N_1970,N_1879);
and U2438 (N_2438,N_1976,N_1949);
or U2439 (N_2439,N_1629,N_1628);
nor U2440 (N_2440,N_1654,N_1889);
nand U2441 (N_2441,N_1636,N_1852);
nor U2442 (N_2442,N_1912,N_1827);
nand U2443 (N_2443,N_1723,N_1997);
xnor U2444 (N_2444,N_1967,N_1870);
and U2445 (N_2445,N_1909,N_1733);
xor U2446 (N_2446,N_1500,N_1983);
nor U2447 (N_2447,N_1645,N_1871);
or U2448 (N_2448,N_1608,N_1779);
and U2449 (N_2449,N_1910,N_1834);
and U2450 (N_2450,N_1740,N_1873);
or U2451 (N_2451,N_1894,N_1883);
nand U2452 (N_2452,N_1781,N_1918);
or U2453 (N_2453,N_1988,N_1756);
nand U2454 (N_2454,N_1643,N_1606);
nand U2455 (N_2455,N_1796,N_1539);
nand U2456 (N_2456,N_1844,N_1521);
nand U2457 (N_2457,N_1949,N_1668);
xnor U2458 (N_2458,N_1652,N_1535);
xor U2459 (N_2459,N_1936,N_1510);
xor U2460 (N_2460,N_1955,N_1912);
and U2461 (N_2461,N_1903,N_1880);
nand U2462 (N_2462,N_1673,N_1885);
xnor U2463 (N_2463,N_1847,N_1842);
xor U2464 (N_2464,N_1935,N_1882);
or U2465 (N_2465,N_1551,N_1918);
nand U2466 (N_2466,N_1648,N_1527);
xor U2467 (N_2467,N_1624,N_1929);
or U2468 (N_2468,N_1732,N_1738);
nand U2469 (N_2469,N_1896,N_1532);
nand U2470 (N_2470,N_1931,N_1723);
nor U2471 (N_2471,N_1745,N_1537);
nand U2472 (N_2472,N_1768,N_1895);
and U2473 (N_2473,N_1541,N_1552);
xor U2474 (N_2474,N_1988,N_1918);
nor U2475 (N_2475,N_1725,N_1537);
nand U2476 (N_2476,N_1876,N_1564);
xor U2477 (N_2477,N_1787,N_1953);
nand U2478 (N_2478,N_1888,N_1721);
and U2479 (N_2479,N_1703,N_1621);
nor U2480 (N_2480,N_1779,N_1617);
xnor U2481 (N_2481,N_1630,N_1887);
xnor U2482 (N_2482,N_1931,N_1577);
nand U2483 (N_2483,N_1984,N_1954);
nand U2484 (N_2484,N_1915,N_1711);
nand U2485 (N_2485,N_1995,N_1537);
nand U2486 (N_2486,N_1720,N_1779);
nand U2487 (N_2487,N_1751,N_1530);
and U2488 (N_2488,N_1650,N_1772);
and U2489 (N_2489,N_1654,N_1790);
nand U2490 (N_2490,N_1884,N_1969);
and U2491 (N_2491,N_1875,N_1509);
or U2492 (N_2492,N_1975,N_1794);
or U2493 (N_2493,N_1724,N_1847);
nand U2494 (N_2494,N_1599,N_1751);
nand U2495 (N_2495,N_1863,N_1644);
and U2496 (N_2496,N_1504,N_1697);
and U2497 (N_2497,N_1986,N_1979);
or U2498 (N_2498,N_1640,N_1892);
xor U2499 (N_2499,N_1710,N_1668);
or U2500 (N_2500,N_2499,N_2156);
or U2501 (N_2501,N_2294,N_2204);
and U2502 (N_2502,N_2066,N_2118);
or U2503 (N_2503,N_2049,N_2009);
and U2504 (N_2504,N_2478,N_2295);
or U2505 (N_2505,N_2025,N_2189);
xor U2506 (N_2506,N_2007,N_2381);
and U2507 (N_2507,N_2271,N_2325);
xor U2508 (N_2508,N_2101,N_2013);
and U2509 (N_2509,N_2423,N_2020);
nor U2510 (N_2510,N_2053,N_2203);
xor U2511 (N_2511,N_2067,N_2158);
or U2512 (N_2512,N_2397,N_2222);
xnor U2513 (N_2513,N_2105,N_2446);
xor U2514 (N_2514,N_2154,N_2087);
and U2515 (N_2515,N_2200,N_2039);
xnor U2516 (N_2516,N_2250,N_2029);
nor U2517 (N_2517,N_2371,N_2050);
nand U2518 (N_2518,N_2255,N_2035);
nor U2519 (N_2519,N_2473,N_2012);
and U2520 (N_2520,N_2194,N_2424);
xnor U2521 (N_2521,N_2292,N_2491);
xnor U2522 (N_2522,N_2162,N_2305);
nor U2523 (N_2523,N_2430,N_2403);
or U2524 (N_2524,N_2248,N_2246);
or U2525 (N_2525,N_2128,N_2361);
nor U2526 (N_2526,N_2316,N_2445);
nor U2527 (N_2527,N_2169,N_2108);
nand U2528 (N_2528,N_2151,N_2284);
and U2529 (N_2529,N_2330,N_2047);
or U2530 (N_2530,N_2016,N_2187);
nand U2531 (N_2531,N_2133,N_2398);
nand U2532 (N_2532,N_2394,N_2166);
nand U2533 (N_2533,N_2319,N_2464);
xnor U2534 (N_2534,N_2136,N_2280);
nand U2535 (N_2535,N_2211,N_2412);
or U2536 (N_2536,N_2475,N_2161);
or U2537 (N_2537,N_2006,N_2326);
nor U2538 (N_2538,N_2487,N_2389);
xor U2539 (N_2539,N_2438,N_2202);
or U2540 (N_2540,N_2314,N_2405);
nor U2541 (N_2541,N_2086,N_2076);
nand U2542 (N_2542,N_2436,N_2228);
or U2543 (N_2543,N_2437,N_2071);
or U2544 (N_2544,N_2341,N_2180);
nor U2545 (N_2545,N_2213,N_2480);
nand U2546 (N_2546,N_2345,N_2278);
nor U2547 (N_2547,N_2494,N_2269);
nand U2548 (N_2548,N_2093,N_2283);
nand U2549 (N_2549,N_2429,N_2303);
or U2550 (N_2550,N_2090,N_2034);
xor U2551 (N_2551,N_2221,N_2210);
nor U2552 (N_2552,N_2315,N_2380);
xnor U2553 (N_2553,N_2028,N_2056);
or U2554 (N_2554,N_2289,N_2214);
nand U2555 (N_2555,N_2374,N_2163);
xnor U2556 (N_2556,N_2311,N_2324);
and U2557 (N_2557,N_2462,N_2011);
and U2558 (N_2558,N_2068,N_2363);
and U2559 (N_2559,N_2279,N_2425);
xnor U2560 (N_2560,N_2134,N_2103);
xor U2561 (N_2561,N_2415,N_2454);
nor U2562 (N_2562,N_2059,N_2064);
nor U2563 (N_2563,N_2320,N_2342);
xor U2564 (N_2564,N_2336,N_2083);
xor U2565 (N_2565,N_2057,N_2227);
nor U2566 (N_2566,N_2078,N_2252);
nand U2567 (N_2567,N_2061,N_2370);
or U2568 (N_2568,N_2205,N_2178);
nand U2569 (N_2569,N_2416,N_2096);
xor U2570 (N_2570,N_2321,N_2244);
nand U2571 (N_2571,N_2075,N_2104);
or U2572 (N_2572,N_2002,N_2331);
and U2573 (N_2573,N_2275,N_2463);
and U2574 (N_2574,N_2179,N_2355);
nand U2575 (N_2575,N_2447,N_2209);
or U2576 (N_2576,N_2024,N_2120);
nor U2577 (N_2577,N_2082,N_2334);
nand U2578 (N_2578,N_2198,N_2339);
xnor U2579 (N_2579,N_2492,N_2015);
xnor U2580 (N_2580,N_2469,N_2155);
nand U2581 (N_2581,N_2407,N_2377);
and U2582 (N_2582,N_2130,N_2387);
and U2583 (N_2583,N_2411,N_2040);
xnor U2584 (N_2584,N_2185,N_2450);
or U2585 (N_2585,N_2100,N_2441);
or U2586 (N_2586,N_2309,N_2270);
nor U2587 (N_2587,N_2274,N_2175);
nand U2588 (N_2588,N_2106,N_2135);
nand U2589 (N_2589,N_2132,N_2223);
and U2590 (N_2590,N_2063,N_2490);
xor U2591 (N_2591,N_2043,N_2141);
or U2592 (N_2592,N_2125,N_2253);
nand U2593 (N_2593,N_2351,N_2240);
xor U2594 (N_2594,N_2297,N_2408);
nor U2595 (N_2595,N_2052,N_2045);
and U2596 (N_2596,N_2177,N_2033);
nand U2597 (N_2597,N_2460,N_2384);
nor U2598 (N_2598,N_2299,N_2391);
nand U2599 (N_2599,N_2433,N_2428);
or U2600 (N_2600,N_2137,N_2335);
nand U2601 (N_2601,N_2296,N_2207);
or U2602 (N_2602,N_2262,N_2085);
nor U2603 (N_2603,N_2353,N_2367);
and U2604 (N_2604,N_2308,N_2476);
or U2605 (N_2605,N_2212,N_2323);
or U2606 (N_2606,N_2307,N_2030);
nand U2607 (N_2607,N_2281,N_2152);
xor U2608 (N_2608,N_2483,N_2406);
and U2609 (N_2609,N_2109,N_2413);
xor U2610 (N_2610,N_2258,N_2074);
nor U2611 (N_2611,N_2265,N_2467);
xnor U2612 (N_2612,N_2129,N_2392);
xnor U2613 (N_2613,N_2306,N_2461);
nand U2614 (N_2614,N_2036,N_2216);
xor U2615 (N_2615,N_2486,N_2373);
or U2616 (N_2616,N_2218,N_2268);
and U2617 (N_2617,N_2208,N_2466);
nand U2618 (N_2618,N_2038,N_2426);
nor U2619 (N_2619,N_2089,N_2010);
nor U2620 (N_2620,N_2440,N_2195);
xnor U2621 (N_2621,N_2239,N_2354);
nand U2622 (N_2622,N_2375,N_2482);
nor U2623 (N_2623,N_2282,N_2472);
or U2624 (N_2624,N_2004,N_2470);
nand U2625 (N_2625,N_2298,N_2251);
or U2626 (N_2626,N_2001,N_2116);
xnor U2627 (N_2627,N_2399,N_2121);
xor U2628 (N_2628,N_2317,N_2044);
nand U2629 (N_2629,N_2184,N_2113);
nor U2630 (N_2630,N_2419,N_2149);
nor U2631 (N_2631,N_2144,N_2172);
and U2632 (N_2632,N_2287,N_2372);
or U2633 (N_2633,N_2427,N_2322);
nor U2634 (N_2634,N_2414,N_2062);
nor U2635 (N_2635,N_2496,N_2362);
nor U2636 (N_2636,N_2365,N_2358);
or U2637 (N_2637,N_2422,N_2140);
or U2638 (N_2638,N_2349,N_2146);
xnor U2639 (N_2639,N_2174,N_2329);
and U2640 (N_2640,N_2165,N_2219);
and U2641 (N_2641,N_2031,N_2225);
and U2642 (N_2642,N_2410,N_2272);
nand U2643 (N_2643,N_2388,N_2153);
xor U2644 (N_2644,N_2193,N_2400);
xor U2645 (N_2645,N_2098,N_2379);
xor U2646 (N_2646,N_2164,N_2452);
or U2647 (N_2647,N_2254,N_2019);
nand U2648 (N_2648,N_2084,N_2266);
nand U2649 (N_2649,N_2139,N_2160);
nand U2650 (N_2650,N_2267,N_2479);
nand U2651 (N_2651,N_2333,N_2233);
or U2652 (N_2652,N_2097,N_2263);
nor U2653 (N_2653,N_2451,N_2347);
xnor U2654 (N_2654,N_2092,N_2008);
nand U2655 (N_2655,N_2310,N_2366);
nor U2656 (N_2656,N_2245,N_2069);
nand U2657 (N_2657,N_2247,N_2201);
or U2658 (N_2658,N_2455,N_2493);
and U2659 (N_2659,N_2236,N_2286);
nor U2660 (N_2660,N_2114,N_2364);
xnor U2661 (N_2661,N_2359,N_2000);
or U2662 (N_2662,N_2264,N_2256);
or U2663 (N_2663,N_2344,N_2439);
and U2664 (N_2664,N_2032,N_2022);
or U2665 (N_2665,N_2402,N_2386);
nand U2666 (N_2666,N_2396,N_2259);
nand U2667 (N_2667,N_2368,N_2434);
xor U2668 (N_2668,N_2277,N_2348);
xor U2669 (N_2669,N_2220,N_2147);
or U2670 (N_2670,N_2276,N_2291);
or U2671 (N_2671,N_2376,N_2023);
xnor U2672 (N_2672,N_2060,N_2079);
xnor U2673 (N_2673,N_2337,N_2046);
and U2674 (N_2674,N_2126,N_2070);
and U2675 (N_2675,N_2356,N_2188);
and U2676 (N_2676,N_2453,N_2346);
or U2677 (N_2677,N_2058,N_2215);
xor U2678 (N_2678,N_2168,N_2197);
nand U2679 (N_2679,N_2091,N_2350);
xor U2680 (N_2680,N_2054,N_2488);
nand U2681 (N_2681,N_2115,N_2431);
xor U2682 (N_2682,N_2312,N_2042);
nor U2683 (N_2683,N_2393,N_2094);
and U2684 (N_2684,N_2241,N_2099);
and U2685 (N_2685,N_2474,N_2382);
or U2686 (N_2686,N_2173,N_2018);
xor U2687 (N_2687,N_2420,N_2449);
xnor U2688 (N_2688,N_2338,N_2051);
and U2689 (N_2689,N_2229,N_2261);
or U2690 (N_2690,N_2003,N_2107);
nor U2691 (N_2691,N_2465,N_2055);
nor U2692 (N_2692,N_2182,N_2448);
nor U2693 (N_2693,N_2378,N_2235);
and U2694 (N_2694,N_2357,N_2199);
xnor U2695 (N_2695,N_2148,N_2131);
or U2696 (N_2696,N_2484,N_2167);
xnor U2697 (N_2697,N_2112,N_2077);
or U2698 (N_2698,N_2138,N_2159);
nor U2699 (N_2699,N_2192,N_2206);
and U2700 (N_2700,N_2327,N_2457);
or U2701 (N_2701,N_2444,N_2142);
xnor U2702 (N_2702,N_2095,N_2421);
and U2703 (N_2703,N_2468,N_2196);
xor U2704 (N_2704,N_2290,N_2318);
nor U2705 (N_2705,N_2170,N_2226);
or U2706 (N_2706,N_2369,N_2111);
or U2707 (N_2707,N_2065,N_2014);
xnor U2708 (N_2708,N_2285,N_2048);
nor U2709 (N_2709,N_2385,N_2328);
nor U2710 (N_2710,N_2224,N_2217);
or U2711 (N_2711,N_2110,N_2080);
nor U2712 (N_2712,N_2143,N_2238);
nor U2713 (N_2713,N_2237,N_2288);
xor U2714 (N_2714,N_2150,N_2304);
or U2715 (N_2715,N_2234,N_2390);
nor U2716 (N_2716,N_2257,N_2191);
and U2717 (N_2717,N_2021,N_2127);
nor U2718 (N_2718,N_2443,N_2293);
and U2719 (N_2719,N_2026,N_2458);
xor U2720 (N_2720,N_2343,N_2383);
nor U2721 (N_2721,N_2360,N_2401);
or U2722 (N_2722,N_2190,N_2300);
nor U2723 (N_2723,N_2302,N_2489);
and U2724 (N_2724,N_2171,N_2027);
nor U2725 (N_2725,N_2481,N_2242);
and U2726 (N_2726,N_2157,N_2497);
nor U2727 (N_2727,N_2395,N_2005);
nand U2728 (N_2728,N_2230,N_2081);
xor U2729 (N_2729,N_2124,N_2243);
xnor U2730 (N_2730,N_2301,N_2495);
nor U2731 (N_2731,N_2249,N_2260);
and U2732 (N_2732,N_2041,N_2477);
nand U2733 (N_2733,N_2471,N_2037);
nor U2734 (N_2734,N_2119,N_2435);
nand U2735 (N_2735,N_2072,N_2485);
and U2736 (N_2736,N_2352,N_2017);
or U2737 (N_2737,N_2232,N_2183);
nand U2738 (N_2738,N_2088,N_2231);
or U2739 (N_2739,N_2409,N_2404);
nand U2740 (N_2740,N_2418,N_2145);
xnor U2741 (N_2741,N_2117,N_2456);
and U2742 (N_2742,N_2181,N_2122);
xor U2743 (N_2743,N_2442,N_2313);
nand U2744 (N_2744,N_2340,N_2273);
or U2745 (N_2745,N_2459,N_2498);
xnor U2746 (N_2746,N_2186,N_2102);
nor U2747 (N_2747,N_2332,N_2123);
and U2748 (N_2748,N_2176,N_2073);
xor U2749 (N_2749,N_2432,N_2417);
xnor U2750 (N_2750,N_2251,N_2074);
or U2751 (N_2751,N_2278,N_2055);
or U2752 (N_2752,N_2418,N_2077);
and U2753 (N_2753,N_2350,N_2411);
or U2754 (N_2754,N_2415,N_2273);
and U2755 (N_2755,N_2220,N_2475);
xnor U2756 (N_2756,N_2211,N_2342);
nand U2757 (N_2757,N_2098,N_2124);
nor U2758 (N_2758,N_2224,N_2103);
nor U2759 (N_2759,N_2180,N_2351);
nand U2760 (N_2760,N_2274,N_2200);
xor U2761 (N_2761,N_2314,N_2327);
xor U2762 (N_2762,N_2472,N_2076);
nor U2763 (N_2763,N_2027,N_2450);
or U2764 (N_2764,N_2249,N_2221);
xor U2765 (N_2765,N_2081,N_2325);
nor U2766 (N_2766,N_2083,N_2250);
nor U2767 (N_2767,N_2381,N_2483);
nor U2768 (N_2768,N_2289,N_2141);
or U2769 (N_2769,N_2232,N_2468);
or U2770 (N_2770,N_2007,N_2413);
xor U2771 (N_2771,N_2470,N_2220);
nand U2772 (N_2772,N_2103,N_2088);
xnor U2773 (N_2773,N_2223,N_2313);
nand U2774 (N_2774,N_2369,N_2455);
and U2775 (N_2775,N_2129,N_2122);
nand U2776 (N_2776,N_2347,N_2494);
nand U2777 (N_2777,N_2476,N_2067);
nor U2778 (N_2778,N_2069,N_2022);
and U2779 (N_2779,N_2013,N_2386);
nand U2780 (N_2780,N_2123,N_2438);
nor U2781 (N_2781,N_2330,N_2426);
and U2782 (N_2782,N_2302,N_2083);
or U2783 (N_2783,N_2370,N_2109);
xor U2784 (N_2784,N_2356,N_2052);
or U2785 (N_2785,N_2131,N_2142);
or U2786 (N_2786,N_2179,N_2287);
and U2787 (N_2787,N_2405,N_2051);
nor U2788 (N_2788,N_2418,N_2127);
nor U2789 (N_2789,N_2176,N_2121);
xnor U2790 (N_2790,N_2112,N_2025);
and U2791 (N_2791,N_2344,N_2088);
and U2792 (N_2792,N_2436,N_2323);
or U2793 (N_2793,N_2464,N_2106);
or U2794 (N_2794,N_2291,N_2159);
and U2795 (N_2795,N_2494,N_2417);
nand U2796 (N_2796,N_2128,N_2119);
or U2797 (N_2797,N_2137,N_2311);
or U2798 (N_2798,N_2450,N_2133);
nand U2799 (N_2799,N_2337,N_2489);
or U2800 (N_2800,N_2397,N_2152);
xor U2801 (N_2801,N_2193,N_2207);
xor U2802 (N_2802,N_2117,N_2050);
and U2803 (N_2803,N_2138,N_2037);
xnor U2804 (N_2804,N_2446,N_2130);
nand U2805 (N_2805,N_2304,N_2027);
or U2806 (N_2806,N_2177,N_2433);
nand U2807 (N_2807,N_2178,N_2456);
or U2808 (N_2808,N_2262,N_2297);
xnor U2809 (N_2809,N_2491,N_2493);
or U2810 (N_2810,N_2020,N_2056);
and U2811 (N_2811,N_2169,N_2264);
xor U2812 (N_2812,N_2394,N_2345);
nand U2813 (N_2813,N_2124,N_2364);
or U2814 (N_2814,N_2265,N_2020);
nor U2815 (N_2815,N_2059,N_2004);
nor U2816 (N_2816,N_2269,N_2295);
xor U2817 (N_2817,N_2320,N_2003);
and U2818 (N_2818,N_2296,N_2102);
and U2819 (N_2819,N_2135,N_2332);
nand U2820 (N_2820,N_2215,N_2455);
and U2821 (N_2821,N_2153,N_2077);
nand U2822 (N_2822,N_2043,N_2002);
nand U2823 (N_2823,N_2148,N_2132);
nand U2824 (N_2824,N_2115,N_2451);
or U2825 (N_2825,N_2208,N_2356);
nor U2826 (N_2826,N_2222,N_2276);
and U2827 (N_2827,N_2131,N_2481);
xnor U2828 (N_2828,N_2270,N_2047);
nor U2829 (N_2829,N_2387,N_2252);
nand U2830 (N_2830,N_2227,N_2045);
nor U2831 (N_2831,N_2229,N_2365);
nor U2832 (N_2832,N_2215,N_2417);
xor U2833 (N_2833,N_2336,N_2206);
nor U2834 (N_2834,N_2447,N_2173);
xnor U2835 (N_2835,N_2066,N_2374);
and U2836 (N_2836,N_2418,N_2300);
xor U2837 (N_2837,N_2160,N_2341);
or U2838 (N_2838,N_2279,N_2170);
and U2839 (N_2839,N_2416,N_2201);
and U2840 (N_2840,N_2153,N_2066);
xor U2841 (N_2841,N_2055,N_2036);
nand U2842 (N_2842,N_2319,N_2233);
and U2843 (N_2843,N_2378,N_2139);
and U2844 (N_2844,N_2301,N_2170);
and U2845 (N_2845,N_2414,N_2336);
nand U2846 (N_2846,N_2161,N_2006);
or U2847 (N_2847,N_2286,N_2064);
nand U2848 (N_2848,N_2298,N_2389);
xor U2849 (N_2849,N_2287,N_2041);
nand U2850 (N_2850,N_2068,N_2040);
xnor U2851 (N_2851,N_2462,N_2328);
nand U2852 (N_2852,N_2255,N_2361);
or U2853 (N_2853,N_2355,N_2322);
xnor U2854 (N_2854,N_2318,N_2305);
nor U2855 (N_2855,N_2356,N_2207);
nand U2856 (N_2856,N_2038,N_2377);
or U2857 (N_2857,N_2042,N_2010);
nor U2858 (N_2858,N_2161,N_2256);
and U2859 (N_2859,N_2147,N_2241);
and U2860 (N_2860,N_2007,N_2089);
or U2861 (N_2861,N_2070,N_2270);
nand U2862 (N_2862,N_2058,N_2183);
nand U2863 (N_2863,N_2130,N_2102);
nor U2864 (N_2864,N_2343,N_2128);
nor U2865 (N_2865,N_2023,N_2065);
and U2866 (N_2866,N_2375,N_2095);
or U2867 (N_2867,N_2493,N_2371);
xor U2868 (N_2868,N_2179,N_2136);
and U2869 (N_2869,N_2064,N_2303);
xnor U2870 (N_2870,N_2092,N_2005);
or U2871 (N_2871,N_2201,N_2121);
xor U2872 (N_2872,N_2023,N_2113);
nand U2873 (N_2873,N_2250,N_2341);
or U2874 (N_2874,N_2316,N_2336);
and U2875 (N_2875,N_2247,N_2179);
and U2876 (N_2876,N_2370,N_2266);
or U2877 (N_2877,N_2084,N_2481);
nor U2878 (N_2878,N_2081,N_2208);
and U2879 (N_2879,N_2389,N_2054);
nor U2880 (N_2880,N_2492,N_2261);
nor U2881 (N_2881,N_2078,N_2431);
and U2882 (N_2882,N_2272,N_2076);
nor U2883 (N_2883,N_2027,N_2345);
nor U2884 (N_2884,N_2015,N_2105);
nand U2885 (N_2885,N_2213,N_2087);
and U2886 (N_2886,N_2466,N_2128);
xor U2887 (N_2887,N_2472,N_2105);
and U2888 (N_2888,N_2260,N_2198);
nand U2889 (N_2889,N_2209,N_2386);
and U2890 (N_2890,N_2109,N_2152);
and U2891 (N_2891,N_2398,N_2113);
nor U2892 (N_2892,N_2255,N_2167);
or U2893 (N_2893,N_2492,N_2335);
nor U2894 (N_2894,N_2023,N_2421);
and U2895 (N_2895,N_2198,N_2316);
nor U2896 (N_2896,N_2270,N_2297);
or U2897 (N_2897,N_2269,N_2360);
nand U2898 (N_2898,N_2068,N_2212);
nor U2899 (N_2899,N_2190,N_2229);
or U2900 (N_2900,N_2366,N_2111);
and U2901 (N_2901,N_2237,N_2259);
nand U2902 (N_2902,N_2266,N_2143);
and U2903 (N_2903,N_2342,N_2456);
or U2904 (N_2904,N_2153,N_2137);
nor U2905 (N_2905,N_2464,N_2316);
nand U2906 (N_2906,N_2398,N_2496);
nor U2907 (N_2907,N_2482,N_2421);
and U2908 (N_2908,N_2020,N_2222);
nor U2909 (N_2909,N_2405,N_2046);
nor U2910 (N_2910,N_2416,N_2215);
nor U2911 (N_2911,N_2395,N_2238);
or U2912 (N_2912,N_2427,N_2005);
nand U2913 (N_2913,N_2185,N_2238);
or U2914 (N_2914,N_2126,N_2246);
nor U2915 (N_2915,N_2458,N_2323);
nand U2916 (N_2916,N_2357,N_2453);
xnor U2917 (N_2917,N_2382,N_2381);
nand U2918 (N_2918,N_2158,N_2272);
or U2919 (N_2919,N_2306,N_2370);
nor U2920 (N_2920,N_2254,N_2429);
nor U2921 (N_2921,N_2431,N_2311);
nand U2922 (N_2922,N_2378,N_2433);
nor U2923 (N_2923,N_2299,N_2189);
nand U2924 (N_2924,N_2199,N_2475);
xnor U2925 (N_2925,N_2358,N_2319);
and U2926 (N_2926,N_2166,N_2208);
nand U2927 (N_2927,N_2405,N_2422);
nor U2928 (N_2928,N_2299,N_2024);
xor U2929 (N_2929,N_2220,N_2090);
nor U2930 (N_2930,N_2079,N_2061);
xor U2931 (N_2931,N_2246,N_2069);
nand U2932 (N_2932,N_2323,N_2085);
xor U2933 (N_2933,N_2052,N_2197);
or U2934 (N_2934,N_2367,N_2406);
nor U2935 (N_2935,N_2239,N_2018);
nand U2936 (N_2936,N_2004,N_2366);
or U2937 (N_2937,N_2234,N_2320);
xor U2938 (N_2938,N_2277,N_2212);
and U2939 (N_2939,N_2238,N_2357);
or U2940 (N_2940,N_2329,N_2409);
nand U2941 (N_2941,N_2274,N_2167);
nor U2942 (N_2942,N_2201,N_2164);
nor U2943 (N_2943,N_2054,N_2307);
xor U2944 (N_2944,N_2156,N_2402);
and U2945 (N_2945,N_2446,N_2464);
xor U2946 (N_2946,N_2406,N_2177);
nor U2947 (N_2947,N_2291,N_2325);
nand U2948 (N_2948,N_2004,N_2403);
or U2949 (N_2949,N_2208,N_2083);
nor U2950 (N_2950,N_2063,N_2060);
and U2951 (N_2951,N_2249,N_2205);
or U2952 (N_2952,N_2084,N_2030);
xnor U2953 (N_2953,N_2296,N_2481);
xnor U2954 (N_2954,N_2427,N_2308);
nand U2955 (N_2955,N_2135,N_2498);
or U2956 (N_2956,N_2073,N_2399);
xnor U2957 (N_2957,N_2260,N_2153);
and U2958 (N_2958,N_2171,N_2233);
nor U2959 (N_2959,N_2007,N_2203);
and U2960 (N_2960,N_2445,N_2317);
or U2961 (N_2961,N_2285,N_2378);
nand U2962 (N_2962,N_2175,N_2296);
and U2963 (N_2963,N_2279,N_2069);
and U2964 (N_2964,N_2256,N_2276);
xor U2965 (N_2965,N_2227,N_2166);
xnor U2966 (N_2966,N_2477,N_2130);
and U2967 (N_2967,N_2341,N_2351);
nor U2968 (N_2968,N_2013,N_2012);
nand U2969 (N_2969,N_2246,N_2475);
nor U2970 (N_2970,N_2002,N_2182);
or U2971 (N_2971,N_2190,N_2036);
and U2972 (N_2972,N_2450,N_2046);
xnor U2973 (N_2973,N_2416,N_2497);
and U2974 (N_2974,N_2330,N_2279);
nor U2975 (N_2975,N_2126,N_2315);
nand U2976 (N_2976,N_2060,N_2360);
nor U2977 (N_2977,N_2187,N_2297);
and U2978 (N_2978,N_2314,N_2497);
nor U2979 (N_2979,N_2002,N_2314);
xnor U2980 (N_2980,N_2446,N_2173);
or U2981 (N_2981,N_2189,N_2349);
nor U2982 (N_2982,N_2001,N_2488);
nand U2983 (N_2983,N_2028,N_2113);
xor U2984 (N_2984,N_2280,N_2169);
and U2985 (N_2985,N_2138,N_2178);
or U2986 (N_2986,N_2453,N_2088);
xor U2987 (N_2987,N_2016,N_2064);
nor U2988 (N_2988,N_2427,N_2347);
or U2989 (N_2989,N_2350,N_2460);
and U2990 (N_2990,N_2402,N_2397);
nand U2991 (N_2991,N_2157,N_2316);
or U2992 (N_2992,N_2138,N_2094);
and U2993 (N_2993,N_2027,N_2150);
and U2994 (N_2994,N_2103,N_2023);
nand U2995 (N_2995,N_2193,N_2345);
or U2996 (N_2996,N_2455,N_2142);
and U2997 (N_2997,N_2145,N_2361);
and U2998 (N_2998,N_2153,N_2474);
xnor U2999 (N_2999,N_2127,N_2120);
nor UO_0 (O_0,N_2588,N_2820);
and UO_1 (O_1,N_2677,N_2688);
nor UO_2 (O_2,N_2650,N_2888);
nand UO_3 (O_3,N_2609,N_2945);
nand UO_4 (O_4,N_2872,N_2699);
xnor UO_5 (O_5,N_2674,N_2540);
nor UO_6 (O_6,N_2806,N_2840);
or UO_7 (O_7,N_2605,N_2722);
nor UO_8 (O_8,N_2902,N_2816);
nor UO_9 (O_9,N_2793,N_2852);
nand UO_10 (O_10,N_2886,N_2538);
nor UO_11 (O_11,N_2817,N_2660);
nor UO_12 (O_12,N_2864,N_2532);
or UO_13 (O_13,N_2529,N_2685);
or UO_14 (O_14,N_2910,N_2720);
xnor UO_15 (O_15,N_2687,N_2871);
nand UO_16 (O_16,N_2726,N_2638);
xor UO_17 (O_17,N_2512,N_2896);
nor UO_18 (O_18,N_2866,N_2736);
xor UO_19 (O_19,N_2525,N_2510);
nand UO_20 (O_20,N_2616,N_2978);
and UO_21 (O_21,N_2517,N_2653);
nor UO_22 (O_22,N_2671,N_2966);
xor UO_23 (O_23,N_2516,N_2629);
or UO_24 (O_24,N_2577,N_2795);
and UO_25 (O_25,N_2649,N_2785);
and UO_26 (O_26,N_2711,N_2825);
nor UO_27 (O_27,N_2654,N_2701);
nor UO_28 (O_28,N_2933,N_2514);
xnor UO_29 (O_29,N_2704,N_2927);
nand UO_30 (O_30,N_2786,N_2628);
or UO_31 (O_31,N_2734,N_2857);
nor UO_32 (O_32,N_2503,N_2944);
and UO_33 (O_33,N_2752,N_2707);
nand UO_34 (O_34,N_2600,N_2909);
nor UO_35 (O_35,N_2501,N_2784);
xnor UO_36 (O_36,N_2770,N_2964);
nand UO_37 (O_37,N_2782,N_2723);
and UO_38 (O_38,N_2568,N_2606);
nand UO_39 (O_39,N_2700,N_2647);
nand UO_40 (O_40,N_2889,N_2810);
nor UO_41 (O_41,N_2648,N_2682);
or UO_42 (O_42,N_2845,N_2772);
and UO_43 (O_43,N_2839,N_2661);
nand UO_44 (O_44,N_2999,N_2958);
and UO_45 (O_45,N_2504,N_2854);
nand UO_46 (O_46,N_2943,N_2994);
or UO_47 (O_47,N_2565,N_2598);
xor UO_48 (O_48,N_2611,N_2849);
nand UO_49 (O_49,N_2774,N_2899);
or UO_50 (O_50,N_2977,N_2741);
nand UO_51 (O_51,N_2619,N_2923);
nor UO_52 (O_52,N_2878,N_2885);
nor UO_53 (O_53,N_2562,N_2986);
or UO_54 (O_54,N_2823,N_2582);
nor UO_55 (O_55,N_2563,N_2881);
nand UO_56 (O_56,N_2815,N_2744);
nor UO_57 (O_57,N_2993,N_2937);
nand UO_58 (O_58,N_2938,N_2891);
xnor UO_59 (O_59,N_2995,N_2511);
xor UO_60 (O_60,N_2928,N_2608);
nand UO_61 (O_61,N_2718,N_2818);
nor UO_62 (O_62,N_2897,N_2528);
or UO_63 (O_63,N_2560,N_2740);
and UO_64 (O_64,N_2811,N_2610);
and UO_65 (O_65,N_2919,N_2939);
xor UO_66 (O_66,N_2614,N_2860);
and UO_67 (O_67,N_2581,N_2961);
xor UO_68 (O_68,N_2679,N_2951);
xnor UO_69 (O_69,N_2515,N_2513);
or UO_70 (O_70,N_2658,N_2756);
or UO_71 (O_71,N_2584,N_2554);
xor UO_72 (O_72,N_2890,N_2997);
or UO_73 (O_73,N_2953,N_2981);
or UO_74 (O_74,N_2985,N_2791);
xnor UO_75 (O_75,N_2970,N_2796);
xor UO_76 (O_76,N_2874,N_2742);
or UO_77 (O_77,N_2809,N_2631);
nand UO_78 (O_78,N_2830,N_2859);
nor UO_79 (O_79,N_2989,N_2672);
and UO_80 (O_80,N_2753,N_2690);
nand UO_81 (O_81,N_2664,N_2968);
nor UO_82 (O_82,N_2789,N_2666);
or UO_83 (O_83,N_2963,N_2586);
nand UO_84 (O_84,N_2965,N_2644);
or UO_85 (O_85,N_2637,N_2551);
xor UO_86 (O_86,N_2534,N_2662);
xor UO_87 (O_87,N_2773,N_2694);
and UO_88 (O_88,N_2639,N_2876);
nor UO_89 (O_89,N_2522,N_2911);
or UO_90 (O_90,N_2670,N_2659);
and UO_91 (O_91,N_2814,N_2642);
nor UO_92 (O_92,N_2634,N_2903);
xor UO_93 (O_93,N_2549,N_2983);
nor UO_94 (O_94,N_2573,N_2622);
nor UO_95 (O_95,N_2776,N_2717);
nor UO_96 (O_96,N_2617,N_2724);
or UO_97 (O_97,N_2657,N_2526);
xnor UO_98 (O_98,N_2761,N_2775);
nand UO_99 (O_99,N_2802,N_2940);
or UO_100 (O_100,N_2745,N_2680);
or UO_101 (O_101,N_2865,N_2804);
nand UO_102 (O_102,N_2507,N_2675);
and UO_103 (O_103,N_2768,N_2976);
or UO_104 (O_104,N_2844,N_2974);
and UO_105 (O_105,N_2781,N_2751);
and UO_106 (O_106,N_2557,N_2728);
nor UO_107 (O_107,N_2867,N_2641);
nand UO_108 (O_108,N_2797,N_2545);
or UO_109 (O_109,N_2596,N_2835);
or UO_110 (O_110,N_2813,N_2992);
xnor UO_111 (O_111,N_2508,N_2962);
xnor UO_112 (O_112,N_2920,N_2935);
or UO_113 (O_113,N_2851,N_2901);
or UO_114 (O_114,N_2542,N_2640);
xor UO_115 (O_115,N_2807,N_2645);
nor UO_116 (O_116,N_2877,N_2838);
or UO_117 (O_117,N_2843,N_2906);
or UO_118 (O_118,N_2982,N_2550);
nand UO_119 (O_119,N_2623,N_2957);
xnor UO_120 (O_120,N_2754,N_2698);
and UO_121 (O_121,N_2712,N_2873);
nor UO_122 (O_122,N_2692,N_2959);
nor UO_123 (O_123,N_2721,N_2571);
and UO_124 (O_124,N_2651,N_2710);
nor UO_125 (O_125,N_2719,N_2758);
nor UO_126 (O_126,N_2892,N_2521);
xor UO_127 (O_127,N_2912,N_2856);
xor UO_128 (O_128,N_2831,N_2686);
nand UO_129 (O_129,N_2738,N_2618);
xnor UO_130 (O_130,N_2778,N_2926);
and UO_131 (O_131,N_2587,N_2621);
nand UO_132 (O_132,N_2601,N_2597);
and UO_133 (O_133,N_2829,N_2625);
nand UO_134 (O_134,N_2805,N_2533);
nor UO_135 (O_135,N_2669,N_2567);
nor UO_136 (O_136,N_2783,N_2833);
xnor UO_137 (O_137,N_2530,N_2705);
nand UO_138 (O_138,N_2564,N_2907);
and UO_139 (O_139,N_2553,N_2627);
nand UO_140 (O_140,N_2991,N_2547);
or UO_141 (O_141,N_2612,N_2633);
nor UO_142 (O_142,N_2914,N_2603);
and UO_143 (O_143,N_2537,N_2714);
and UO_144 (O_144,N_2769,N_2821);
and UO_145 (O_145,N_2592,N_2599);
xor UO_146 (O_146,N_2760,N_2518);
xnor UO_147 (O_147,N_2570,N_2942);
nand UO_148 (O_148,N_2763,N_2822);
nand UO_149 (O_149,N_2536,N_2980);
nor UO_150 (O_150,N_2737,N_2613);
nand UO_151 (O_151,N_2996,N_2936);
or UO_152 (O_152,N_2904,N_2713);
and UO_153 (O_153,N_2759,N_2556);
or UO_154 (O_154,N_2779,N_2579);
nor UO_155 (O_155,N_2555,N_2652);
xnor UO_156 (O_156,N_2749,N_2743);
nor UO_157 (O_157,N_2764,N_2930);
nor UO_158 (O_158,N_2915,N_2655);
xor UO_159 (O_159,N_2541,N_2590);
xnor UO_160 (O_160,N_2826,N_2837);
nor UO_161 (O_161,N_2561,N_2569);
xor UO_162 (O_162,N_2543,N_2746);
and UO_163 (O_163,N_2841,N_2520);
xnor UO_164 (O_164,N_2762,N_2973);
or UO_165 (O_165,N_2956,N_2635);
nand UO_166 (O_166,N_2998,N_2850);
xor UO_167 (O_167,N_2566,N_2790);
xor UO_168 (O_168,N_2552,N_2729);
xor UO_169 (O_169,N_2620,N_2636);
nand UO_170 (O_170,N_2572,N_2574);
and UO_171 (O_171,N_2895,N_2683);
xnor UO_172 (O_172,N_2934,N_2708);
xor UO_173 (O_173,N_2788,N_2955);
or UO_174 (O_174,N_2893,N_2548);
nor UO_175 (O_175,N_2748,N_2665);
or UO_176 (O_176,N_2656,N_2531);
xor UO_177 (O_177,N_2583,N_2602);
xor UO_178 (O_178,N_2727,N_2663);
and UO_179 (O_179,N_2913,N_2500);
or UO_180 (O_180,N_2787,N_2924);
xor UO_181 (O_181,N_2702,N_2643);
xor UO_182 (O_182,N_2506,N_2546);
and UO_183 (O_183,N_2971,N_2767);
or UO_184 (O_184,N_2931,N_2676);
nand UO_185 (O_185,N_2502,N_2735);
xnor UO_186 (O_186,N_2929,N_2509);
nor UO_187 (O_187,N_2585,N_2979);
xor UO_188 (O_188,N_2731,N_2703);
or UO_189 (O_189,N_2750,N_2969);
or UO_190 (O_190,N_2824,N_2771);
or UO_191 (O_191,N_2594,N_2800);
nor UO_192 (O_192,N_2880,N_2862);
xor UO_193 (O_193,N_2855,N_2696);
xor UO_194 (O_194,N_2960,N_2887);
nand UO_195 (O_195,N_2861,N_2595);
and UO_196 (O_196,N_2803,N_2539);
xor UO_197 (O_197,N_2747,N_2716);
or UO_198 (O_198,N_2626,N_2578);
nor UO_199 (O_199,N_2863,N_2681);
and UO_200 (O_200,N_2917,N_2755);
and UO_201 (O_201,N_2832,N_2990);
xor UO_202 (O_202,N_2527,N_2615);
nor UO_203 (O_203,N_2725,N_2870);
nor UO_204 (O_204,N_2827,N_2535);
xnor UO_205 (O_205,N_2975,N_2524);
or UO_206 (O_206,N_2801,N_2875);
and UO_207 (O_207,N_2766,N_2580);
xnor UO_208 (O_208,N_2836,N_2921);
xnor UO_209 (O_209,N_2646,N_2946);
xnor UO_210 (O_210,N_2544,N_2894);
nor UO_211 (O_211,N_2847,N_2792);
nand UO_212 (O_212,N_2984,N_2689);
nand UO_213 (O_213,N_2591,N_2632);
nor UO_214 (O_214,N_2730,N_2883);
and UO_215 (O_215,N_2794,N_2706);
xor UO_216 (O_216,N_2739,N_2882);
and UO_217 (O_217,N_2954,N_2918);
and UO_218 (O_218,N_2624,N_2678);
nor UO_219 (O_219,N_2828,N_2842);
or UO_220 (O_220,N_2922,N_2673);
nand UO_221 (O_221,N_2905,N_2967);
and UO_222 (O_222,N_2630,N_2898);
nor UO_223 (O_223,N_2575,N_2733);
nor UO_224 (O_224,N_2949,N_2668);
or UO_225 (O_225,N_2916,N_2869);
xor UO_226 (O_226,N_2972,N_2819);
or UO_227 (O_227,N_2848,N_2709);
xor UO_228 (O_228,N_2777,N_2948);
nor UO_229 (O_229,N_2812,N_2559);
xor UO_230 (O_230,N_2941,N_2715);
nor UO_231 (O_231,N_2932,N_2684);
nor UO_232 (O_232,N_2765,N_2523);
nand UO_233 (O_233,N_2693,N_2576);
and UO_234 (O_234,N_2952,N_2519);
xnor UO_235 (O_235,N_2950,N_2604);
or UO_236 (O_236,N_2798,N_2834);
xnor UO_237 (O_237,N_2505,N_2589);
or UO_238 (O_238,N_2947,N_2884);
or UO_239 (O_239,N_2695,N_2853);
nand UO_240 (O_240,N_2868,N_2697);
and UO_241 (O_241,N_2900,N_2732);
and UO_242 (O_242,N_2691,N_2925);
or UO_243 (O_243,N_2593,N_2558);
and UO_244 (O_244,N_2858,N_2988);
nor UO_245 (O_245,N_2846,N_2987);
nor UO_246 (O_246,N_2879,N_2607);
or UO_247 (O_247,N_2780,N_2808);
nor UO_248 (O_248,N_2908,N_2667);
or UO_249 (O_249,N_2799,N_2757);
xnor UO_250 (O_250,N_2808,N_2719);
xnor UO_251 (O_251,N_2581,N_2644);
and UO_252 (O_252,N_2503,N_2802);
or UO_253 (O_253,N_2568,N_2574);
xnor UO_254 (O_254,N_2894,N_2614);
nor UO_255 (O_255,N_2798,N_2973);
nor UO_256 (O_256,N_2779,N_2609);
xnor UO_257 (O_257,N_2745,N_2914);
xor UO_258 (O_258,N_2961,N_2678);
and UO_259 (O_259,N_2675,N_2670);
xor UO_260 (O_260,N_2818,N_2975);
or UO_261 (O_261,N_2932,N_2597);
or UO_262 (O_262,N_2586,N_2569);
and UO_263 (O_263,N_2694,N_2561);
or UO_264 (O_264,N_2692,N_2922);
nor UO_265 (O_265,N_2778,N_2799);
and UO_266 (O_266,N_2911,N_2645);
or UO_267 (O_267,N_2673,N_2536);
or UO_268 (O_268,N_2574,N_2540);
nand UO_269 (O_269,N_2797,N_2808);
nor UO_270 (O_270,N_2782,N_2826);
and UO_271 (O_271,N_2520,N_2665);
or UO_272 (O_272,N_2640,N_2695);
or UO_273 (O_273,N_2879,N_2968);
xor UO_274 (O_274,N_2539,N_2521);
and UO_275 (O_275,N_2807,N_2712);
or UO_276 (O_276,N_2533,N_2784);
xnor UO_277 (O_277,N_2779,N_2887);
nand UO_278 (O_278,N_2849,N_2707);
nor UO_279 (O_279,N_2500,N_2794);
or UO_280 (O_280,N_2674,N_2527);
or UO_281 (O_281,N_2870,N_2679);
nor UO_282 (O_282,N_2976,N_2509);
nand UO_283 (O_283,N_2942,N_2952);
or UO_284 (O_284,N_2834,N_2650);
or UO_285 (O_285,N_2936,N_2645);
or UO_286 (O_286,N_2532,N_2594);
nor UO_287 (O_287,N_2719,N_2644);
or UO_288 (O_288,N_2561,N_2910);
nand UO_289 (O_289,N_2800,N_2850);
nand UO_290 (O_290,N_2896,N_2532);
xor UO_291 (O_291,N_2843,N_2535);
and UO_292 (O_292,N_2778,N_2785);
or UO_293 (O_293,N_2636,N_2768);
xor UO_294 (O_294,N_2566,N_2727);
and UO_295 (O_295,N_2987,N_2556);
xnor UO_296 (O_296,N_2685,N_2509);
and UO_297 (O_297,N_2773,N_2906);
nand UO_298 (O_298,N_2850,N_2848);
xor UO_299 (O_299,N_2709,N_2988);
nand UO_300 (O_300,N_2860,N_2953);
xnor UO_301 (O_301,N_2821,N_2801);
nand UO_302 (O_302,N_2647,N_2744);
xnor UO_303 (O_303,N_2611,N_2544);
nor UO_304 (O_304,N_2939,N_2568);
or UO_305 (O_305,N_2595,N_2838);
xor UO_306 (O_306,N_2659,N_2550);
or UO_307 (O_307,N_2518,N_2575);
and UO_308 (O_308,N_2778,N_2751);
and UO_309 (O_309,N_2966,N_2599);
nor UO_310 (O_310,N_2921,N_2507);
nor UO_311 (O_311,N_2877,N_2611);
or UO_312 (O_312,N_2707,N_2828);
nor UO_313 (O_313,N_2737,N_2797);
nand UO_314 (O_314,N_2686,N_2927);
xor UO_315 (O_315,N_2889,N_2674);
and UO_316 (O_316,N_2551,N_2729);
and UO_317 (O_317,N_2724,N_2894);
or UO_318 (O_318,N_2741,N_2579);
or UO_319 (O_319,N_2570,N_2680);
nor UO_320 (O_320,N_2946,N_2654);
and UO_321 (O_321,N_2896,N_2693);
xnor UO_322 (O_322,N_2996,N_2605);
nor UO_323 (O_323,N_2619,N_2620);
nor UO_324 (O_324,N_2895,N_2794);
nor UO_325 (O_325,N_2700,N_2623);
and UO_326 (O_326,N_2775,N_2963);
nand UO_327 (O_327,N_2559,N_2839);
nor UO_328 (O_328,N_2651,N_2632);
xor UO_329 (O_329,N_2763,N_2839);
xnor UO_330 (O_330,N_2920,N_2577);
nand UO_331 (O_331,N_2964,N_2922);
or UO_332 (O_332,N_2671,N_2924);
and UO_333 (O_333,N_2519,N_2811);
and UO_334 (O_334,N_2781,N_2989);
or UO_335 (O_335,N_2832,N_2859);
xnor UO_336 (O_336,N_2645,N_2561);
or UO_337 (O_337,N_2931,N_2911);
xor UO_338 (O_338,N_2749,N_2702);
nor UO_339 (O_339,N_2624,N_2592);
and UO_340 (O_340,N_2944,N_2568);
nand UO_341 (O_341,N_2797,N_2729);
nor UO_342 (O_342,N_2699,N_2583);
nand UO_343 (O_343,N_2749,N_2645);
xnor UO_344 (O_344,N_2712,N_2931);
xnor UO_345 (O_345,N_2948,N_2577);
and UO_346 (O_346,N_2746,N_2802);
nand UO_347 (O_347,N_2987,N_2829);
and UO_348 (O_348,N_2677,N_2580);
nor UO_349 (O_349,N_2776,N_2587);
or UO_350 (O_350,N_2934,N_2935);
nand UO_351 (O_351,N_2571,N_2958);
and UO_352 (O_352,N_2844,N_2954);
and UO_353 (O_353,N_2965,N_2893);
xnor UO_354 (O_354,N_2666,N_2559);
or UO_355 (O_355,N_2580,N_2813);
or UO_356 (O_356,N_2757,N_2733);
or UO_357 (O_357,N_2652,N_2913);
xor UO_358 (O_358,N_2779,N_2977);
nand UO_359 (O_359,N_2682,N_2840);
nand UO_360 (O_360,N_2556,N_2886);
nor UO_361 (O_361,N_2757,N_2992);
xor UO_362 (O_362,N_2568,N_2931);
xor UO_363 (O_363,N_2596,N_2697);
xnor UO_364 (O_364,N_2556,N_2856);
nor UO_365 (O_365,N_2625,N_2938);
nor UO_366 (O_366,N_2863,N_2674);
xor UO_367 (O_367,N_2830,N_2793);
and UO_368 (O_368,N_2828,N_2503);
nand UO_369 (O_369,N_2763,N_2644);
or UO_370 (O_370,N_2825,N_2627);
and UO_371 (O_371,N_2554,N_2762);
or UO_372 (O_372,N_2541,N_2891);
and UO_373 (O_373,N_2608,N_2916);
nand UO_374 (O_374,N_2637,N_2523);
xnor UO_375 (O_375,N_2852,N_2719);
nor UO_376 (O_376,N_2531,N_2808);
and UO_377 (O_377,N_2725,N_2773);
or UO_378 (O_378,N_2728,N_2544);
or UO_379 (O_379,N_2605,N_2570);
xor UO_380 (O_380,N_2766,N_2891);
and UO_381 (O_381,N_2886,N_2992);
nor UO_382 (O_382,N_2949,N_2974);
xor UO_383 (O_383,N_2740,N_2709);
and UO_384 (O_384,N_2556,N_2619);
and UO_385 (O_385,N_2761,N_2932);
xor UO_386 (O_386,N_2561,N_2725);
or UO_387 (O_387,N_2558,N_2975);
or UO_388 (O_388,N_2866,N_2949);
or UO_389 (O_389,N_2613,N_2780);
or UO_390 (O_390,N_2549,N_2554);
or UO_391 (O_391,N_2629,N_2521);
or UO_392 (O_392,N_2720,N_2533);
nand UO_393 (O_393,N_2845,N_2911);
nand UO_394 (O_394,N_2532,N_2762);
nor UO_395 (O_395,N_2881,N_2917);
and UO_396 (O_396,N_2603,N_2869);
nand UO_397 (O_397,N_2561,N_2935);
nor UO_398 (O_398,N_2805,N_2693);
xnor UO_399 (O_399,N_2908,N_2896);
nor UO_400 (O_400,N_2597,N_2531);
or UO_401 (O_401,N_2869,N_2833);
xor UO_402 (O_402,N_2964,N_2863);
nor UO_403 (O_403,N_2969,N_2634);
or UO_404 (O_404,N_2513,N_2798);
or UO_405 (O_405,N_2966,N_2851);
nor UO_406 (O_406,N_2883,N_2933);
or UO_407 (O_407,N_2786,N_2505);
and UO_408 (O_408,N_2896,N_2878);
nand UO_409 (O_409,N_2901,N_2654);
nor UO_410 (O_410,N_2545,N_2660);
nor UO_411 (O_411,N_2623,N_2515);
nor UO_412 (O_412,N_2525,N_2788);
and UO_413 (O_413,N_2548,N_2837);
and UO_414 (O_414,N_2557,N_2744);
or UO_415 (O_415,N_2788,N_2524);
nand UO_416 (O_416,N_2847,N_2788);
nor UO_417 (O_417,N_2858,N_2910);
or UO_418 (O_418,N_2595,N_2776);
nor UO_419 (O_419,N_2833,N_2562);
xor UO_420 (O_420,N_2741,N_2763);
nor UO_421 (O_421,N_2763,N_2637);
or UO_422 (O_422,N_2817,N_2594);
nand UO_423 (O_423,N_2984,N_2851);
or UO_424 (O_424,N_2939,N_2960);
or UO_425 (O_425,N_2835,N_2582);
nor UO_426 (O_426,N_2606,N_2917);
nor UO_427 (O_427,N_2921,N_2813);
nand UO_428 (O_428,N_2814,N_2904);
nor UO_429 (O_429,N_2685,N_2597);
or UO_430 (O_430,N_2982,N_2806);
xnor UO_431 (O_431,N_2991,N_2669);
nor UO_432 (O_432,N_2848,N_2641);
nand UO_433 (O_433,N_2832,N_2501);
nor UO_434 (O_434,N_2515,N_2747);
nand UO_435 (O_435,N_2568,N_2779);
or UO_436 (O_436,N_2802,N_2978);
xor UO_437 (O_437,N_2825,N_2590);
nand UO_438 (O_438,N_2981,N_2797);
or UO_439 (O_439,N_2904,N_2602);
nand UO_440 (O_440,N_2550,N_2541);
nor UO_441 (O_441,N_2713,N_2850);
and UO_442 (O_442,N_2811,N_2739);
or UO_443 (O_443,N_2683,N_2743);
xnor UO_444 (O_444,N_2622,N_2837);
nand UO_445 (O_445,N_2699,N_2568);
nand UO_446 (O_446,N_2701,N_2950);
and UO_447 (O_447,N_2550,N_2813);
xnor UO_448 (O_448,N_2977,N_2529);
nor UO_449 (O_449,N_2886,N_2626);
xor UO_450 (O_450,N_2553,N_2927);
xor UO_451 (O_451,N_2634,N_2549);
xor UO_452 (O_452,N_2784,N_2825);
nand UO_453 (O_453,N_2636,N_2991);
nor UO_454 (O_454,N_2529,N_2659);
and UO_455 (O_455,N_2833,N_2620);
nor UO_456 (O_456,N_2691,N_2736);
nand UO_457 (O_457,N_2985,N_2780);
or UO_458 (O_458,N_2976,N_2697);
xor UO_459 (O_459,N_2770,N_2807);
nand UO_460 (O_460,N_2894,N_2932);
nand UO_461 (O_461,N_2698,N_2594);
and UO_462 (O_462,N_2843,N_2557);
xnor UO_463 (O_463,N_2987,N_2946);
nand UO_464 (O_464,N_2691,N_2979);
nor UO_465 (O_465,N_2923,N_2875);
or UO_466 (O_466,N_2565,N_2771);
or UO_467 (O_467,N_2803,N_2506);
or UO_468 (O_468,N_2764,N_2894);
xor UO_469 (O_469,N_2688,N_2530);
or UO_470 (O_470,N_2780,N_2870);
or UO_471 (O_471,N_2627,N_2628);
or UO_472 (O_472,N_2806,N_2931);
or UO_473 (O_473,N_2532,N_2578);
and UO_474 (O_474,N_2790,N_2922);
or UO_475 (O_475,N_2864,N_2632);
or UO_476 (O_476,N_2920,N_2618);
xor UO_477 (O_477,N_2609,N_2634);
and UO_478 (O_478,N_2576,N_2773);
nor UO_479 (O_479,N_2588,N_2722);
nand UO_480 (O_480,N_2628,N_2536);
nand UO_481 (O_481,N_2589,N_2753);
nor UO_482 (O_482,N_2807,N_2833);
nand UO_483 (O_483,N_2843,N_2995);
xnor UO_484 (O_484,N_2682,N_2764);
nor UO_485 (O_485,N_2627,N_2885);
nor UO_486 (O_486,N_2636,N_2914);
or UO_487 (O_487,N_2587,N_2763);
and UO_488 (O_488,N_2577,N_2838);
nand UO_489 (O_489,N_2509,N_2560);
nand UO_490 (O_490,N_2853,N_2577);
nand UO_491 (O_491,N_2693,N_2728);
nand UO_492 (O_492,N_2559,N_2528);
nand UO_493 (O_493,N_2667,N_2880);
or UO_494 (O_494,N_2876,N_2724);
or UO_495 (O_495,N_2938,N_2961);
nand UO_496 (O_496,N_2941,N_2582);
or UO_497 (O_497,N_2875,N_2957);
xor UO_498 (O_498,N_2649,N_2679);
and UO_499 (O_499,N_2902,N_2646);
endmodule