module basic_750_5000_1000_10_levels_5xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_611,In_90);
and U1 (N_1,In_368,In_205);
xnor U2 (N_2,In_150,In_407);
nor U3 (N_3,In_248,In_235);
nand U4 (N_4,In_355,In_658);
and U5 (N_5,In_741,In_599);
or U6 (N_6,In_613,In_614);
and U7 (N_7,In_366,In_23);
or U8 (N_8,In_274,In_500);
or U9 (N_9,In_172,In_626);
and U10 (N_10,In_344,In_211);
and U11 (N_11,In_67,In_543);
and U12 (N_12,In_226,In_224);
nor U13 (N_13,In_335,In_582);
or U14 (N_14,In_625,In_578);
or U15 (N_15,In_505,In_53);
and U16 (N_16,In_714,In_487);
nand U17 (N_17,In_256,In_33);
nor U18 (N_18,In_214,In_508);
or U19 (N_19,In_557,In_501);
nor U20 (N_20,In_583,In_587);
or U21 (N_21,In_137,In_301);
and U22 (N_22,In_424,In_432);
or U23 (N_23,In_607,In_526);
or U24 (N_24,In_398,In_523);
nand U25 (N_25,In_437,In_725);
xor U26 (N_26,In_654,In_695);
and U27 (N_27,In_32,In_215);
and U28 (N_28,In_401,In_25);
nand U29 (N_29,In_157,In_151);
nand U30 (N_30,In_118,In_569);
nor U31 (N_31,In_649,In_497);
nor U32 (N_32,In_650,In_732);
or U33 (N_33,In_306,In_704);
or U34 (N_34,In_553,In_676);
nor U35 (N_35,In_309,In_162);
nor U36 (N_36,In_455,In_351);
nor U37 (N_37,In_632,In_46);
nor U38 (N_38,In_721,In_337);
nand U39 (N_39,In_324,In_166);
nand U40 (N_40,In_155,In_488);
and U41 (N_41,In_713,In_209);
or U42 (N_42,In_472,In_646);
or U43 (N_43,In_651,In_185);
or U44 (N_44,In_194,In_122);
nand U45 (N_45,In_100,In_482);
nor U46 (N_46,In_664,In_675);
nand U47 (N_47,In_8,In_636);
nand U48 (N_48,In_656,In_711);
and U49 (N_49,In_669,In_643);
nor U50 (N_50,In_445,In_384);
nor U51 (N_51,In_561,In_492);
and U52 (N_52,In_298,In_255);
nand U53 (N_53,In_580,In_165);
xnor U54 (N_54,In_665,In_623);
xnor U55 (N_55,In_45,In_289);
nor U56 (N_56,In_184,In_189);
nand U57 (N_57,In_173,In_320);
nor U58 (N_58,In_302,In_449);
and U59 (N_59,In_18,In_571);
xnor U60 (N_60,In_710,In_315);
nand U61 (N_61,In_633,In_383);
and U62 (N_62,In_388,In_575);
or U63 (N_63,In_551,In_264);
nand U64 (N_64,In_135,In_360);
nor U65 (N_65,In_400,In_683);
or U66 (N_66,In_498,In_534);
nor U67 (N_67,In_568,In_556);
nor U68 (N_68,In_602,In_250);
xnor U69 (N_69,In_567,In_736);
or U70 (N_70,In_120,In_516);
nand U71 (N_71,In_57,In_719);
and U72 (N_72,In_51,In_177);
xnor U73 (N_73,In_574,In_59);
nand U74 (N_74,In_481,In_409);
nor U75 (N_75,In_300,In_674);
xnor U76 (N_76,In_573,In_346);
nand U77 (N_77,In_510,In_609);
xnor U78 (N_78,In_365,In_478);
nand U79 (N_79,In_86,In_446);
and U80 (N_80,In_180,In_463);
xor U81 (N_81,In_295,In_297);
and U82 (N_82,In_486,In_584);
or U83 (N_83,In_415,In_56);
nand U84 (N_84,In_240,In_630);
or U85 (N_85,In_434,In_413);
and U86 (N_86,In_363,In_386);
or U87 (N_87,In_462,In_700);
xor U88 (N_88,In_164,In_405);
nand U89 (N_89,In_742,In_629);
xor U90 (N_90,In_545,In_410);
and U91 (N_91,In_85,In_483);
nor U92 (N_92,In_603,In_290);
and U93 (N_93,In_475,In_348);
nor U94 (N_94,In_378,In_114);
and U95 (N_95,In_749,In_570);
nand U96 (N_96,In_99,In_506);
and U97 (N_97,In_531,In_287);
nor U98 (N_98,In_361,In_113);
nand U99 (N_99,In_98,In_266);
xnor U100 (N_100,In_682,In_563);
or U101 (N_101,In_436,In_225);
xor U102 (N_102,In_572,In_179);
or U103 (N_103,In_75,In_514);
nand U104 (N_104,In_332,In_52);
nor U105 (N_105,In_369,In_129);
nand U106 (N_106,In_291,In_110);
nand U107 (N_107,In_132,In_202);
nand U108 (N_108,In_727,In_37);
nor U109 (N_109,In_97,In_198);
or U110 (N_110,In_484,In_688);
or U111 (N_111,In_616,In_601);
nand U112 (N_112,In_93,In_222);
or U113 (N_113,In_586,In_538);
nand U114 (N_114,In_62,In_660);
nor U115 (N_115,In_564,In_159);
xnor U116 (N_116,In_303,In_652);
nor U117 (N_117,In_10,In_252);
or U118 (N_118,In_319,In_152);
and U119 (N_119,In_269,In_236);
and U120 (N_120,In_154,In_68);
or U121 (N_121,In_178,In_588);
nor U122 (N_122,In_627,In_589);
xor U123 (N_123,In_524,In_525);
nand U124 (N_124,In_380,In_89);
nor U125 (N_125,In_147,In_49);
and U126 (N_126,In_653,In_304);
and U127 (N_127,In_429,In_82);
and U128 (N_128,In_27,In_36);
and U129 (N_129,In_313,In_206);
and U130 (N_130,In_352,In_188);
or U131 (N_131,In_493,In_321);
nor U132 (N_132,In_680,In_458);
or U133 (N_133,In_343,In_530);
xor U134 (N_134,In_280,In_513);
or U135 (N_135,In_195,In_310);
or U136 (N_136,In_681,In_697);
and U137 (N_137,In_55,In_708);
and U138 (N_138,In_375,In_316);
or U139 (N_139,In_119,In_447);
nand U140 (N_140,In_515,In_464);
nor U141 (N_141,In_167,In_423);
xor U142 (N_142,In_123,In_126);
nand U143 (N_143,In_40,In_376);
nand U144 (N_144,In_43,In_473);
nor U145 (N_145,In_237,In_38);
and U146 (N_146,In_596,In_696);
and U147 (N_147,In_91,In_77);
and U148 (N_148,In_581,In_65);
nor U149 (N_149,In_685,In_29);
xor U150 (N_150,In_456,In_47);
nor U151 (N_151,In_326,In_403);
nand U152 (N_152,In_655,In_428);
nand U153 (N_153,In_707,In_535);
and U154 (N_154,In_311,In_84);
nand U155 (N_155,In_318,In_9);
or U156 (N_156,In_554,In_5);
xor U157 (N_157,In_548,In_372);
and U158 (N_158,In_641,In_171);
nand U159 (N_159,In_334,In_116);
nand U160 (N_160,In_489,In_133);
nor U161 (N_161,In_327,In_537);
nor U162 (N_162,In_495,In_81);
nor U163 (N_163,In_17,In_241);
nor U164 (N_164,In_170,In_693);
or U165 (N_165,In_692,In_420);
or U166 (N_166,In_712,In_267);
nor U167 (N_167,In_738,In_48);
and U168 (N_168,In_592,In_740);
nand U169 (N_169,In_396,In_0);
or U170 (N_170,In_190,In_42);
or U171 (N_171,In_3,In_331);
and U172 (N_172,In_13,In_552);
or U173 (N_173,In_438,In_518);
nor U174 (N_174,In_661,In_591);
nand U175 (N_175,In_71,In_659);
or U176 (N_176,In_540,In_726);
nand U177 (N_177,In_419,In_466);
nor U178 (N_178,In_441,In_109);
or U179 (N_179,In_702,In_296);
nor U180 (N_180,In_148,In_528);
nor U181 (N_181,In_533,In_393);
nor U182 (N_182,In_735,In_325);
nand U183 (N_183,In_207,In_314);
or U184 (N_184,In_21,In_253);
and U185 (N_185,In_465,In_34);
nand U186 (N_186,In_720,In_307);
and U187 (N_187,In_634,In_262);
nand U188 (N_188,In_6,In_229);
nor U189 (N_189,In_662,In_480);
or U190 (N_190,In_520,In_20);
and U191 (N_191,In_156,In_258);
xnor U192 (N_192,In_356,In_16);
or U193 (N_193,In_127,In_699);
and U194 (N_194,In_308,In_729);
and U195 (N_195,In_276,In_340);
nand U196 (N_196,In_427,In_174);
nand U197 (N_197,In_115,In_339);
nor U198 (N_198,In_371,In_451);
and U199 (N_199,In_414,In_670);
and U200 (N_200,In_690,In_312);
nand U201 (N_201,In_233,In_1);
nor U202 (N_202,In_457,In_261);
and U203 (N_203,In_134,In_272);
and U204 (N_204,In_718,In_14);
nand U205 (N_205,In_158,In_370);
or U206 (N_206,In_706,In_559);
and U207 (N_207,In_80,In_349);
nand U208 (N_208,In_391,In_30);
nand U209 (N_209,In_293,In_504);
and U210 (N_210,In_358,In_402);
or U211 (N_211,In_193,In_260);
and U212 (N_212,In_389,In_70);
or U213 (N_213,In_743,In_585);
nand U214 (N_214,In_635,In_353);
nand U215 (N_215,In_620,In_476);
nand U216 (N_216,In_390,In_246);
nand U217 (N_217,In_285,In_657);
nor U218 (N_218,In_183,In_239);
nor U219 (N_219,In_160,In_359);
nand U220 (N_220,In_459,In_92);
nand U221 (N_221,In_558,In_204);
or U222 (N_222,In_357,In_176);
nand U223 (N_223,In_136,In_257);
and U224 (N_224,In_108,In_210);
nand U225 (N_225,In_28,In_31);
nor U226 (N_226,In_731,In_50);
or U227 (N_227,In_496,In_213);
or U228 (N_228,In_672,In_106);
nand U229 (N_229,In_41,In_121);
xnor U230 (N_230,In_4,In_541);
nor U231 (N_231,In_2,In_66);
nand U232 (N_232,In_550,In_679);
nand U233 (N_233,In_329,In_220);
or U234 (N_234,In_141,In_221);
or U235 (N_235,In_734,In_74);
xnor U236 (N_236,In_485,In_689);
and U237 (N_237,In_196,In_527);
xor U238 (N_238,In_460,In_263);
and U239 (N_239,In_364,In_145);
or U240 (N_240,In_644,In_104);
nand U241 (N_241,In_615,In_631);
or U242 (N_242,In_101,In_605);
nand U243 (N_243,In_336,In_439);
and U244 (N_244,In_470,In_238);
nor U245 (N_245,In_593,In_7);
nand U246 (N_246,In_490,In_565);
nand U247 (N_247,In_305,In_219);
or U248 (N_248,In_223,In_547);
xnor U249 (N_249,In_88,In_576);
nand U250 (N_250,In_345,In_181);
xnor U251 (N_251,In_251,In_322);
and U252 (N_252,In_277,In_385);
xor U253 (N_253,In_443,In_83);
and U254 (N_254,In_292,In_430);
nand U255 (N_255,In_283,In_271);
and U256 (N_256,In_507,In_191);
or U257 (N_257,In_595,In_454);
nor U258 (N_258,In_39,In_684);
nand U259 (N_259,In_373,In_694);
nor U260 (N_260,In_395,In_667);
xor U261 (N_261,In_717,In_125);
nor U262 (N_262,In_63,In_622);
or U263 (N_263,In_72,In_124);
nor U264 (N_264,In_19,In_87);
and U265 (N_265,In_218,In_648);
nand U266 (N_266,In_254,In_647);
nand U267 (N_267,In_130,In_15);
nor U268 (N_268,In_617,In_442);
nor U269 (N_269,In_444,In_418);
nor U270 (N_270,In_278,In_733);
nand U271 (N_271,In_330,In_416);
and U272 (N_272,In_161,In_452);
nor U273 (N_273,In_44,In_687);
nor U274 (N_274,In_421,In_79);
and U275 (N_275,In_379,In_73);
or U276 (N_276,In_187,In_76);
nor U277 (N_277,In_200,In_265);
and U278 (N_278,In_666,In_747);
or U279 (N_279,In_317,In_362);
nor U280 (N_280,In_737,In_228);
and U281 (N_281,In_663,In_494);
nand U282 (N_282,In_598,In_408);
and U283 (N_283,In_544,In_399);
nor U284 (N_284,In_431,In_724);
nor U285 (N_285,In_640,In_517);
nand U286 (N_286,In_739,In_612);
and U287 (N_287,In_637,In_342);
or U288 (N_288,In_639,In_60);
and U289 (N_289,In_422,In_64);
xor U290 (N_290,In_281,In_354);
or U291 (N_291,In_243,In_96);
and U292 (N_292,In_227,In_149);
xnor U293 (N_293,In_286,In_536);
nand U294 (N_294,In_404,In_471);
and U295 (N_295,In_678,In_521);
nor U296 (N_296,In_668,In_234);
and U297 (N_297,In_381,In_698);
nand U298 (N_298,In_562,In_102);
xnor U299 (N_299,In_146,In_503);
nor U300 (N_300,In_382,In_279);
nor U301 (N_301,In_11,In_341);
and U302 (N_302,In_701,In_212);
or U303 (N_303,In_268,In_208);
xnor U304 (N_304,In_22,In_705);
nor U305 (N_305,In_140,In_610);
nand U306 (N_306,In_367,In_542);
and U307 (N_307,In_186,In_411);
nor U308 (N_308,In_138,In_294);
xnor U309 (N_309,In_549,In_182);
or U310 (N_310,In_128,In_94);
and U311 (N_311,In_426,In_477);
nand U312 (N_312,In_453,In_673);
nor U313 (N_313,In_144,In_519);
and U314 (N_314,In_577,In_139);
or U315 (N_315,In_412,In_532);
and U316 (N_316,In_450,In_703);
and U317 (N_317,In_288,In_579);
and U318 (N_318,In_539,In_231);
xor U319 (N_319,In_249,In_394);
nand U320 (N_320,In_468,In_745);
or U321 (N_321,In_245,In_645);
or U322 (N_322,In_392,In_716);
and U323 (N_323,In_728,In_35);
nor U324 (N_324,In_107,In_597);
nand U325 (N_325,In_397,In_499);
or U326 (N_326,In_638,In_744);
or U327 (N_327,In_230,In_333);
nor U328 (N_328,In_95,In_105);
nor U329 (N_329,In_555,In_621);
nor U330 (N_330,In_677,In_216);
nand U331 (N_331,In_347,In_203);
or U332 (N_332,In_247,In_479);
nor U333 (N_333,In_299,In_374);
or U334 (N_334,In_512,In_560);
and U335 (N_335,In_270,In_522);
or U336 (N_336,In_604,In_628);
nor U337 (N_337,In_474,In_163);
or U338 (N_338,In_594,In_259);
or U339 (N_339,In_417,In_748);
xnor U340 (N_340,In_529,In_217);
nor U341 (N_341,In_606,In_448);
and U342 (N_342,In_103,In_618);
nand U343 (N_343,In_117,In_282);
nand U344 (N_344,In_467,In_168);
and U345 (N_345,In_600,In_26);
nand U346 (N_346,In_619,In_69);
or U347 (N_347,In_377,In_111);
and U348 (N_348,In_509,In_491);
and U349 (N_349,In_723,In_425);
nor U350 (N_350,In_142,In_566);
or U351 (N_351,In_338,In_61);
nor U352 (N_352,In_275,In_78);
nor U353 (N_353,In_284,In_169);
and U354 (N_354,In_350,In_54);
xnor U355 (N_355,In_590,In_244);
and U356 (N_356,In_131,In_273);
or U357 (N_357,In_709,In_433);
and U358 (N_358,In_624,In_671);
nor U359 (N_359,In_58,In_175);
or U360 (N_360,In_511,In_715);
xor U361 (N_361,In_608,In_387);
nor U362 (N_362,In_199,In_197);
and U363 (N_363,In_201,In_546);
or U364 (N_364,In_24,In_242);
or U365 (N_365,In_406,In_232);
nor U366 (N_366,In_12,In_469);
nand U367 (N_367,In_192,In_691);
nand U368 (N_368,In_440,In_730);
xor U369 (N_369,In_686,In_461);
and U370 (N_370,In_328,In_502);
nor U371 (N_371,In_746,In_153);
and U372 (N_372,In_435,In_143);
nand U373 (N_373,In_112,In_722);
nand U374 (N_374,In_642,In_323);
and U375 (N_375,In_379,In_281);
or U376 (N_376,In_121,In_363);
nand U377 (N_377,In_308,In_164);
nand U378 (N_378,In_69,In_94);
or U379 (N_379,In_391,In_439);
nor U380 (N_380,In_297,In_148);
nand U381 (N_381,In_31,In_63);
and U382 (N_382,In_709,In_708);
and U383 (N_383,In_651,In_80);
nand U384 (N_384,In_153,In_468);
nand U385 (N_385,In_575,In_167);
and U386 (N_386,In_700,In_131);
xnor U387 (N_387,In_211,In_22);
xor U388 (N_388,In_96,In_169);
nor U389 (N_389,In_740,In_318);
nor U390 (N_390,In_706,In_314);
xnor U391 (N_391,In_749,In_635);
xnor U392 (N_392,In_705,In_373);
xor U393 (N_393,In_159,In_130);
and U394 (N_394,In_126,In_734);
nand U395 (N_395,In_335,In_455);
nor U396 (N_396,In_339,In_534);
and U397 (N_397,In_632,In_385);
nor U398 (N_398,In_738,In_275);
nor U399 (N_399,In_594,In_289);
nor U400 (N_400,In_392,In_562);
and U401 (N_401,In_662,In_323);
nand U402 (N_402,In_594,In_553);
or U403 (N_403,In_4,In_1);
or U404 (N_404,In_259,In_375);
nor U405 (N_405,In_703,In_604);
nor U406 (N_406,In_439,In_248);
nor U407 (N_407,In_454,In_561);
nand U408 (N_408,In_202,In_709);
nor U409 (N_409,In_445,In_285);
nor U410 (N_410,In_30,In_161);
nor U411 (N_411,In_608,In_711);
xnor U412 (N_412,In_98,In_691);
nand U413 (N_413,In_254,In_142);
or U414 (N_414,In_392,In_267);
or U415 (N_415,In_113,In_690);
nor U416 (N_416,In_214,In_567);
nor U417 (N_417,In_466,In_567);
or U418 (N_418,In_597,In_9);
and U419 (N_419,In_287,In_332);
xnor U420 (N_420,In_272,In_45);
xor U421 (N_421,In_245,In_117);
nor U422 (N_422,In_418,In_678);
and U423 (N_423,In_562,In_598);
and U424 (N_424,In_713,In_656);
nor U425 (N_425,In_452,In_669);
nand U426 (N_426,In_371,In_338);
nor U427 (N_427,In_362,In_714);
and U428 (N_428,In_467,In_498);
and U429 (N_429,In_583,In_433);
nand U430 (N_430,In_444,In_202);
and U431 (N_431,In_625,In_547);
xor U432 (N_432,In_479,In_213);
nand U433 (N_433,In_273,In_172);
or U434 (N_434,In_7,In_415);
nand U435 (N_435,In_157,In_142);
nand U436 (N_436,In_272,In_675);
or U437 (N_437,In_190,In_28);
nor U438 (N_438,In_46,In_152);
or U439 (N_439,In_210,In_131);
or U440 (N_440,In_339,In_149);
nor U441 (N_441,In_81,In_455);
or U442 (N_442,In_73,In_414);
or U443 (N_443,In_719,In_561);
and U444 (N_444,In_475,In_615);
or U445 (N_445,In_101,In_168);
nand U446 (N_446,In_345,In_455);
nor U447 (N_447,In_132,In_470);
and U448 (N_448,In_104,In_684);
nor U449 (N_449,In_588,In_111);
and U450 (N_450,In_389,In_128);
and U451 (N_451,In_605,In_425);
and U452 (N_452,In_276,In_434);
xnor U453 (N_453,In_494,In_498);
nor U454 (N_454,In_199,In_317);
nor U455 (N_455,In_172,In_702);
and U456 (N_456,In_517,In_568);
xnor U457 (N_457,In_298,In_737);
xor U458 (N_458,In_713,In_134);
nand U459 (N_459,In_235,In_306);
nand U460 (N_460,In_131,In_447);
or U461 (N_461,In_394,In_716);
xor U462 (N_462,In_4,In_60);
nand U463 (N_463,In_138,In_116);
xor U464 (N_464,In_356,In_638);
nor U465 (N_465,In_11,In_499);
and U466 (N_466,In_84,In_690);
nor U467 (N_467,In_356,In_68);
and U468 (N_468,In_601,In_648);
and U469 (N_469,In_489,In_112);
nand U470 (N_470,In_16,In_99);
nand U471 (N_471,In_95,In_534);
nand U472 (N_472,In_232,In_157);
or U473 (N_473,In_26,In_548);
xnor U474 (N_474,In_327,In_267);
and U475 (N_475,In_388,In_390);
nand U476 (N_476,In_696,In_189);
or U477 (N_477,In_647,In_297);
and U478 (N_478,In_569,In_568);
xor U479 (N_479,In_599,In_526);
xor U480 (N_480,In_445,In_642);
xnor U481 (N_481,In_328,In_619);
and U482 (N_482,In_442,In_85);
or U483 (N_483,In_481,In_179);
and U484 (N_484,In_693,In_550);
nor U485 (N_485,In_576,In_748);
nor U486 (N_486,In_226,In_652);
nand U487 (N_487,In_549,In_364);
nand U488 (N_488,In_739,In_706);
and U489 (N_489,In_380,In_164);
nor U490 (N_490,In_411,In_202);
and U491 (N_491,In_109,In_580);
and U492 (N_492,In_678,In_168);
or U493 (N_493,In_78,In_289);
or U494 (N_494,In_231,In_391);
or U495 (N_495,In_389,In_535);
xor U496 (N_496,In_342,In_33);
xor U497 (N_497,In_734,In_158);
nand U498 (N_498,In_68,In_353);
nand U499 (N_499,In_714,In_318);
and U500 (N_500,N_248,N_483);
xnor U501 (N_501,N_310,N_356);
nor U502 (N_502,N_241,N_193);
and U503 (N_503,N_5,N_270);
nand U504 (N_504,N_491,N_405);
and U505 (N_505,N_186,N_52);
and U506 (N_506,N_323,N_219);
xnor U507 (N_507,N_83,N_408);
and U508 (N_508,N_335,N_182);
or U509 (N_509,N_150,N_235);
nand U510 (N_510,N_376,N_226);
and U511 (N_511,N_147,N_80);
and U512 (N_512,N_339,N_149);
xnor U513 (N_513,N_175,N_415);
xnor U514 (N_514,N_343,N_214);
or U515 (N_515,N_199,N_489);
nor U516 (N_516,N_81,N_302);
and U517 (N_517,N_3,N_407);
nand U518 (N_518,N_325,N_113);
nor U519 (N_519,N_69,N_224);
nor U520 (N_520,N_369,N_470);
nor U521 (N_521,N_277,N_90);
nand U522 (N_522,N_11,N_347);
nor U523 (N_523,N_447,N_73);
nor U524 (N_524,N_320,N_333);
nand U525 (N_525,N_265,N_57);
and U526 (N_526,N_422,N_331);
and U527 (N_527,N_161,N_432);
and U528 (N_528,N_173,N_359);
nor U529 (N_529,N_1,N_416);
nand U530 (N_530,N_492,N_151);
and U531 (N_531,N_372,N_401);
xor U532 (N_532,N_109,N_273);
nand U533 (N_533,N_212,N_25);
and U534 (N_534,N_472,N_133);
nor U535 (N_535,N_387,N_388);
nand U536 (N_536,N_227,N_384);
xor U537 (N_537,N_108,N_105);
nor U538 (N_538,N_185,N_46);
nor U539 (N_539,N_378,N_215);
nor U540 (N_540,N_77,N_449);
and U541 (N_541,N_276,N_318);
nor U542 (N_542,N_494,N_375);
nor U543 (N_543,N_423,N_282);
and U544 (N_544,N_36,N_306);
nor U545 (N_545,N_255,N_17);
nor U546 (N_546,N_238,N_464);
or U547 (N_547,N_495,N_354);
and U548 (N_548,N_334,N_294);
xor U549 (N_549,N_385,N_418);
nand U550 (N_550,N_431,N_160);
or U551 (N_551,N_480,N_7);
nand U552 (N_552,N_222,N_9);
and U553 (N_553,N_28,N_18);
nor U554 (N_554,N_350,N_380);
and U555 (N_555,N_330,N_89);
nor U556 (N_556,N_391,N_45);
or U557 (N_557,N_392,N_21);
and U558 (N_558,N_481,N_203);
and U559 (N_559,N_386,N_174);
or U560 (N_560,N_466,N_443);
and U561 (N_561,N_184,N_414);
nand U562 (N_562,N_68,N_194);
nor U563 (N_563,N_413,N_201);
and U564 (N_564,N_338,N_74);
and U565 (N_565,N_435,N_123);
nand U566 (N_566,N_287,N_139);
and U567 (N_567,N_179,N_228);
nand U568 (N_568,N_79,N_128);
and U569 (N_569,N_244,N_279);
or U570 (N_570,N_417,N_8);
and U571 (N_571,N_40,N_22);
nor U572 (N_572,N_498,N_288);
and U573 (N_573,N_313,N_138);
and U574 (N_574,N_180,N_344);
nand U575 (N_575,N_455,N_43);
nor U576 (N_576,N_148,N_2);
nand U577 (N_577,N_75,N_245);
or U578 (N_578,N_252,N_55);
nor U579 (N_579,N_397,N_24);
nor U580 (N_580,N_348,N_462);
and U581 (N_581,N_395,N_463);
nor U582 (N_582,N_256,N_192);
or U583 (N_583,N_58,N_187);
xnor U584 (N_584,N_337,N_322);
or U585 (N_585,N_278,N_188);
or U586 (N_586,N_202,N_299);
or U587 (N_587,N_426,N_357);
nand U588 (N_588,N_353,N_144);
or U589 (N_589,N_86,N_259);
nor U590 (N_590,N_246,N_326);
nand U591 (N_591,N_132,N_439);
xor U592 (N_592,N_368,N_381);
or U593 (N_593,N_66,N_26);
or U594 (N_594,N_383,N_116);
and U595 (N_595,N_84,N_493);
nand U596 (N_596,N_373,N_457);
nor U597 (N_597,N_98,N_140);
and U598 (N_598,N_134,N_200);
and U599 (N_599,N_223,N_284);
and U600 (N_600,N_230,N_307);
or U601 (N_601,N_342,N_289);
or U602 (N_602,N_461,N_217);
nor U603 (N_603,N_154,N_243);
and U604 (N_604,N_196,N_321);
nand U605 (N_605,N_268,N_428);
nor U606 (N_606,N_207,N_400);
nor U607 (N_607,N_379,N_389);
and U608 (N_608,N_233,N_136);
and U609 (N_609,N_363,N_456);
and U610 (N_610,N_459,N_267);
nand U611 (N_611,N_345,N_482);
nand U612 (N_612,N_32,N_314);
or U613 (N_613,N_163,N_117);
or U614 (N_614,N_473,N_42);
nor U615 (N_615,N_239,N_213);
or U616 (N_616,N_390,N_258);
nor U617 (N_617,N_62,N_29);
xor U618 (N_618,N_152,N_118);
or U619 (N_619,N_341,N_290);
nand U620 (N_620,N_436,N_424);
nor U621 (N_621,N_37,N_101);
and U622 (N_622,N_293,N_197);
xnor U623 (N_623,N_155,N_340);
and U624 (N_624,N_41,N_458);
nor U625 (N_625,N_216,N_471);
nor U626 (N_626,N_429,N_178);
nand U627 (N_627,N_153,N_355);
and U628 (N_628,N_486,N_60);
nand U629 (N_629,N_271,N_64);
nor U630 (N_630,N_365,N_70);
and U631 (N_631,N_162,N_169);
nor U632 (N_632,N_309,N_16);
nand U633 (N_633,N_497,N_468);
and U634 (N_634,N_398,N_39);
and U635 (N_635,N_336,N_198);
and U636 (N_636,N_51,N_88);
nor U637 (N_637,N_332,N_304);
or U638 (N_638,N_311,N_121);
and U639 (N_639,N_15,N_351);
or U640 (N_640,N_12,N_484);
nand U641 (N_641,N_76,N_104);
and U642 (N_642,N_263,N_382);
nor U643 (N_643,N_362,N_441);
or U644 (N_644,N_452,N_269);
nand U645 (N_645,N_78,N_240);
nand U646 (N_646,N_301,N_454);
or U647 (N_647,N_20,N_329);
xor U648 (N_648,N_210,N_437);
or U649 (N_649,N_485,N_399);
nor U650 (N_650,N_444,N_63);
and U651 (N_651,N_420,N_448);
or U652 (N_652,N_402,N_396);
nor U653 (N_653,N_442,N_308);
nand U654 (N_654,N_266,N_31);
xor U655 (N_655,N_474,N_445);
nand U656 (N_656,N_167,N_49);
or U657 (N_657,N_54,N_142);
xor U658 (N_658,N_465,N_111);
nand U659 (N_659,N_164,N_158);
or U660 (N_660,N_107,N_124);
nor U661 (N_661,N_170,N_67);
nand U662 (N_662,N_377,N_488);
and U663 (N_663,N_440,N_65);
nor U664 (N_664,N_47,N_253);
nor U665 (N_665,N_23,N_221);
or U666 (N_666,N_126,N_127);
nand U667 (N_667,N_434,N_275);
and U668 (N_668,N_131,N_189);
nand U669 (N_669,N_209,N_319);
or U670 (N_670,N_453,N_92);
nand U671 (N_671,N_499,N_61);
nand U672 (N_672,N_119,N_220);
nand U673 (N_673,N_97,N_291);
and U674 (N_674,N_231,N_249);
nand U675 (N_675,N_349,N_146);
nor U676 (N_676,N_324,N_427);
nor U677 (N_677,N_260,N_394);
nand U678 (N_678,N_300,N_234);
and U679 (N_679,N_410,N_120);
or U680 (N_680,N_10,N_225);
or U681 (N_681,N_176,N_183);
and U682 (N_682,N_430,N_251);
nand U683 (N_683,N_195,N_296);
and U684 (N_684,N_285,N_93);
nand U685 (N_685,N_425,N_177);
nor U686 (N_686,N_460,N_112);
nor U687 (N_687,N_469,N_327);
and U688 (N_688,N_141,N_94);
nor U689 (N_689,N_208,N_19);
and U690 (N_690,N_204,N_206);
or U691 (N_691,N_479,N_451);
xnor U692 (N_692,N_91,N_247);
nand U693 (N_693,N_370,N_286);
nand U694 (N_694,N_237,N_190);
or U695 (N_695,N_145,N_242);
xor U696 (N_696,N_450,N_254);
nor U697 (N_697,N_305,N_371);
and U698 (N_698,N_298,N_53);
nor U699 (N_699,N_44,N_303);
nand U700 (N_700,N_115,N_476);
nand U701 (N_701,N_129,N_110);
or U702 (N_702,N_280,N_143);
and U703 (N_703,N_56,N_85);
and U704 (N_704,N_358,N_157);
nor U705 (N_705,N_487,N_166);
and U706 (N_706,N_114,N_467);
nor U707 (N_707,N_404,N_250);
or U708 (N_708,N_393,N_236);
and U709 (N_709,N_281,N_95);
nand U710 (N_710,N_38,N_364);
or U711 (N_711,N_438,N_419);
and U712 (N_712,N_274,N_317);
and U713 (N_713,N_433,N_211);
or U714 (N_714,N_205,N_6);
and U715 (N_715,N_106,N_159);
or U716 (N_716,N_35,N_374);
xnor U717 (N_717,N_315,N_367);
and U718 (N_718,N_295,N_421);
and U719 (N_719,N_328,N_50);
xnor U720 (N_720,N_100,N_346);
nand U721 (N_721,N_361,N_0);
and U722 (N_722,N_262,N_48);
nand U723 (N_723,N_360,N_27);
or U724 (N_724,N_168,N_292);
or U725 (N_725,N_165,N_130);
nor U726 (N_726,N_272,N_446);
or U727 (N_727,N_103,N_412);
and U728 (N_728,N_30,N_87);
nand U729 (N_729,N_172,N_409);
and U730 (N_730,N_34,N_477);
nand U731 (N_731,N_99,N_4);
or U732 (N_732,N_156,N_283);
nor U733 (N_733,N_403,N_312);
nor U734 (N_734,N_411,N_14);
nor U735 (N_735,N_72,N_478);
and U736 (N_736,N_232,N_137);
nor U737 (N_737,N_125,N_71);
nand U738 (N_738,N_191,N_229);
nand U739 (N_739,N_122,N_33);
nand U740 (N_740,N_490,N_352);
nor U741 (N_741,N_496,N_59);
or U742 (N_742,N_171,N_257);
nand U743 (N_743,N_261,N_316);
nand U744 (N_744,N_82,N_96);
nand U745 (N_745,N_297,N_102);
and U746 (N_746,N_135,N_475);
nand U747 (N_747,N_264,N_181);
nor U748 (N_748,N_218,N_406);
nor U749 (N_749,N_366,N_13);
xnor U750 (N_750,N_178,N_27);
and U751 (N_751,N_347,N_275);
or U752 (N_752,N_206,N_354);
xor U753 (N_753,N_76,N_462);
nand U754 (N_754,N_440,N_57);
nand U755 (N_755,N_230,N_334);
nor U756 (N_756,N_190,N_450);
or U757 (N_757,N_413,N_481);
or U758 (N_758,N_225,N_131);
nor U759 (N_759,N_463,N_459);
and U760 (N_760,N_152,N_219);
nand U761 (N_761,N_284,N_291);
nand U762 (N_762,N_244,N_269);
nand U763 (N_763,N_315,N_145);
and U764 (N_764,N_24,N_42);
xnor U765 (N_765,N_495,N_455);
and U766 (N_766,N_254,N_8);
or U767 (N_767,N_4,N_130);
xor U768 (N_768,N_142,N_430);
or U769 (N_769,N_418,N_119);
or U770 (N_770,N_364,N_84);
nand U771 (N_771,N_38,N_186);
or U772 (N_772,N_190,N_56);
or U773 (N_773,N_225,N_194);
or U774 (N_774,N_388,N_94);
and U775 (N_775,N_460,N_300);
and U776 (N_776,N_474,N_209);
nor U777 (N_777,N_293,N_226);
nand U778 (N_778,N_443,N_347);
or U779 (N_779,N_462,N_403);
and U780 (N_780,N_19,N_443);
nand U781 (N_781,N_64,N_427);
nand U782 (N_782,N_311,N_106);
or U783 (N_783,N_325,N_36);
xnor U784 (N_784,N_28,N_243);
nand U785 (N_785,N_324,N_223);
xor U786 (N_786,N_270,N_365);
nand U787 (N_787,N_193,N_454);
nand U788 (N_788,N_426,N_392);
nor U789 (N_789,N_272,N_86);
or U790 (N_790,N_348,N_359);
and U791 (N_791,N_28,N_440);
nand U792 (N_792,N_13,N_153);
and U793 (N_793,N_207,N_491);
xor U794 (N_794,N_84,N_36);
or U795 (N_795,N_82,N_58);
and U796 (N_796,N_261,N_17);
and U797 (N_797,N_244,N_170);
or U798 (N_798,N_227,N_409);
nor U799 (N_799,N_480,N_309);
and U800 (N_800,N_6,N_35);
nand U801 (N_801,N_414,N_256);
and U802 (N_802,N_237,N_378);
nor U803 (N_803,N_417,N_442);
xnor U804 (N_804,N_322,N_367);
nor U805 (N_805,N_437,N_190);
and U806 (N_806,N_105,N_436);
nor U807 (N_807,N_297,N_284);
or U808 (N_808,N_331,N_385);
nor U809 (N_809,N_286,N_435);
nor U810 (N_810,N_45,N_422);
nor U811 (N_811,N_445,N_84);
or U812 (N_812,N_186,N_161);
and U813 (N_813,N_73,N_213);
and U814 (N_814,N_472,N_48);
nand U815 (N_815,N_452,N_477);
nor U816 (N_816,N_491,N_139);
nor U817 (N_817,N_147,N_420);
xor U818 (N_818,N_320,N_105);
and U819 (N_819,N_216,N_197);
or U820 (N_820,N_106,N_439);
nand U821 (N_821,N_41,N_232);
nand U822 (N_822,N_448,N_357);
or U823 (N_823,N_262,N_344);
xor U824 (N_824,N_300,N_329);
or U825 (N_825,N_335,N_482);
or U826 (N_826,N_472,N_342);
nand U827 (N_827,N_217,N_55);
and U828 (N_828,N_361,N_476);
nand U829 (N_829,N_303,N_64);
nor U830 (N_830,N_465,N_37);
and U831 (N_831,N_224,N_167);
nand U832 (N_832,N_403,N_235);
or U833 (N_833,N_145,N_181);
or U834 (N_834,N_250,N_152);
and U835 (N_835,N_17,N_57);
or U836 (N_836,N_57,N_221);
or U837 (N_837,N_99,N_266);
or U838 (N_838,N_260,N_433);
or U839 (N_839,N_465,N_150);
nand U840 (N_840,N_348,N_326);
or U841 (N_841,N_178,N_211);
nor U842 (N_842,N_212,N_487);
nand U843 (N_843,N_33,N_278);
or U844 (N_844,N_345,N_8);
and U845 (N_845,N_213,N_95);
xor U846 (N_846,N_77,N_478);
or U847 (N_847,N_465,N_263);
nor U848 (N_848,N_427,N_351);
and U849 (N_849,N_165,N_52);
nand U850 (N_850,N_50,N_286);
or U851 (N_851,N_237,N_229);
nand U852 (N_852,N_450,N_320);
or U853 (N_853,N_371,N_178);
nand U854 (N_854,N_397,N_61);
or U855 (N_855,N_136,N_279);
xnor U856 (N_856,N_196,N_249);
xor U857 (N_857,N_157,N_87);
or U858 (N_858,N_317,N_443);
or U859 (N_859,N_272,N_37);
nand U860 (N_860,N_156,N_186);
nand U861 (N_861,N_52,N_276);
and U862 (N_862,N_335,N_110);
or U863 (N_863,N_494,N_366);
and U864 (N_864,N_10,N_494);
nand U865 (N_865,N_358,N_417);
xnor U866 (N_866,N_498,N_105);
nor U867 (N_867,N_335,N_257);
nand U868 (N_868,N_310,N_339);
nand U869 (N_869,N_199,N_486);
or U870 (N_870,N_195,N_406);
nor U871 (N_871,N_120,N_452);
and U872 (N_872,N_283,N_140);
nand U873 (N_873,N_246,N_187);
nor U874 (N_874,N_155,N_466);
xnor U875 (N_875,N_260,N_337);
nand U876 (N_876,N_352,N_233);
or U877 (N_877,N_327,N_47);
nand U878 (N_878,N_125,N_182);
nor U879 (N_879,N_494,N_186);
nand U880 (N_880,N_206,N_247);
nor U881 (N_881,N_295,N_304);
and U882 (N_882,N_130,N_425);
or U883 (N_883,N_425,N_355);
nand U884 (N_884,N_233,N_157);
nor U885 (N_885,N_408,N_152);
nor U886 (N_886,N_178,N_499);
xor U887 (N_887,N_451,N_78);
nand U888 (N_888,N_471,N_425);
or U889 (N_889,N_460,N_38);
xnor U890 (N_890,N_289,N_470);
and U891 (N_891,N_437,N_35);
nand U892 (N_892,N_160,N_137);
or U893 (N_893,N_309,N_259);
and U894 (N_894,N_232,N_141);
nand U895 (N_895,N_486,N_478);
or U896 (N_896,N_315,N_186);
nand U897 (N_897,N_439,N_375);
and U898 (N_898,N_95,N_162);
nor U899 (N_899,N_266,N_235);
nand U900 (N_900,N_73,N_404);
nor U901 (N_901,N_239,N_361);
nor U902 (N_902,N_137,N_384);
nand U903 (N_903,N_140,N_82);
and U904 (N_904,N_208,N_422);
nor U905 (N_905,N_263,N_418);
or U906 (N_906,N_408,N_298);
nor U907 (N_907,N_198,N_488);
nor U908 (N_908,N_50,N_379);
nand U909 (N_909,N_139,N_162);
xnor U910 (N_910,N_1,N_196);
xnor U911 (N_911,N_316,N_179);
nand U912 (N_912,N_21,N_20);
nor U913 (N_913,N_150,N_233);
or U914 (N_914,N_115,N_109);
nor U915 (N_915,N_325,N_217);
or U916 (N_916,N_458,N_129);
and U917 (N_917,N_174,N_51);
and U918 (N_918,N_190,N_486);
or U919 (N_919,N_79,N_203);
or U920 (N_920,N_225,N_8);
xor U921 (N_921,N_433,N_133);
and U922 (N_922,N_159,N_372);
and U923 (N_923,N_180,N_107);
nor U924 (N_924,N_138,N_6);
nor U925 (N_925,N_201,N_457);
and U926 (N_926,N_107,N_424);
xnor U927 (N_927,N_53,N_397);
or U928 (N_928,N_101,N_200);
nand U929 (N_929,N_154,N_296);
nand U930 (N_930,N_228,N_70);
and U931 (N_931,N_35,N_169);
or U932 (N_932,N_133,N_386);
nor U933 (N_933,N_486,N_141);
xnor U934 (N_934,N_488,N_141);
and U935 (N_935,N_146,N_86);
xor U936 (N_936,N_272,N_314);
and U937 (N_937,N_427,N_6);
nor U938 (N_938,N_324,N_185);
or U939 (N_939,N_72,N_359);
nor U940 (N_940,N_50,N_439);
nor U941 (N_941,N_235,N_378);
or U942 (N_942,N_346,N_332);
nor U943 (N_943,N_6,N_470);
nor U944 (N_944,N_468,N_151);
or U945 (N_945,N_390,N_416);
and U946 (N_946,N_162,N_456);
nand U947 (N_947,N_62,N_186);
or U948 (N_948,N_429,N_278);
or U949 (N_949,N_61,N_30);
nand U950 (N_950,N_77,N_185);
nor U951 (N_951,N_448,N_116);
nand U952 (N_952,N_199,N_439);
nand U953 (N_953,N_403,N_283);
nor U954 (N_954,N_26,N_353);
nor U955 (N_955,N_153,N_257);
nor U956 (N_956,N_389,N_162);
nor U957 (N_957,N_393,N_258);
or U958 (N_958,N_312,N_460);
or U959 (N_959,N_393,N_288);
and U960 (N_960,N_181,N_120);
or U961 (N_961,N_352,N_485);
and U962 (N_962,N_88,N_364);
xor U963 (N_963,N_431,N_61);
and U964 (N_964,N_24,N_190);
nand U965 (N_965,N_498,N_164);
and U966 (N_966,N_51,N_232);
nor U967 (N_967,N_350,N_264);
nor U968 (N_968,N_219,N_49);
nand U969 (N_969,N_60,N_349);
or U970 (N_970,N_42,N_460);
nand U971 (N_971,N_448,N_16);
and U972 (N_972,N_220,N_180);
nor U973 (N_973,N_357,N_284);
nor U974 (N_974,N_98,N_244);
and U975 (N_975,N_474,N_391);
nand U976 (N_976,N_75,N_83);
nand U977 (N_977,N_3,N_175);
nor U978 (N_978,N_484,N_14);
or U979 (N_979,N_312,N_412);
nor U980 (N_980,N_289,N_442);
or U981 (N_981,N_268,N_399);
and U982 (N_982,N_158,N_365);
or U983 (N_983,N_229,N_293);
nor U984 (N_984,N_8,N_356);
nand U985 (N_985,N_59,N_61);
or U986 (N_986,N_384,N_373);
nor U987 (N_987,N_332,N_292);
xor U988 (N_988,N_84,N_178);
nor U989 (N_989,N_114,N_182);
and U990 (N_990,N_413,N_131);
nor U991 (N_991,N_434,N_104);
and U992 (N_992,N_396,N_53);
or U993 (N_993,N_27,N_18);
nor U994 (N_994,N_184,N_292);
nand U995 (N_995,N_372,N_260);
xnor U996 (N_996,N_44,N_480);
nand U997 (N_997,N_29,N_143);
or U998 (N_998,N_88,N_141);
nand U999 (N_999,N_437,N_147);
and U1000 (N_1000,N_767,N_789);
nor U1001 (N_1001,N_957,N_748);
and U1002 (N_1002,N_854,N_666);
and U1003 (N_1003,N_723,N_855);
nor U1004 (N_1004,N_742,N_901);
or U1005 (N_1005,N_981,N_583);
or U1006 (N_1006,N_701,N_969);
nand U1007 (N_1007,N_597,N_762);
nor U1008 (N_1008,N_752,N_874);
or U1009 (N_1009,N_770,N_779);
and U1010 (N_1010,N_514,N_962);
and U1011 (N_1011,N_792,N_550);
or U1012 (N_1012,N_986,N_622);
nor U1013 (N_1013,N_538,N_853);
and U1014 (N_1014,N_812,N_655);
nand U1015 (N_1015,N_906,N_523);
and U1016 (N_1016,N_643,N_685);
or U1017 (N_1017,N_988,N_977);
nand U1018 (N_1018,N_927,N_574);
xor U1019 (N_1019,N_949,N_821);
or U1020 (N_1020,N_895,N_995);
nor U1021 (N_1021,N_982,N_570);
nor U1022 (N_1022,N_691,N_890);
or U1023 (N_1023,N_862,N_676);
xnor U1024 (N_1024,N_663,N_684);
nand U1025 (N_1025,N_640,N_781);
and U1026 (N_1026,N_950,N_771);
xor U1027 (N_1027,N_674,N_661);
and U1028 (N_1028,N_599,N_630);
nand U1029 (N_1029,N_780,N_985);
nor U1030 (N_1030,N_823,N_642);
nand U1031 (N_1031,N_860,N_700);
or U1032 (N_1032,N_926,N_559);
xor U1033 (N_1033,N_804,N_932);
and U1034 (N_1034,N_659,N_554);
nor U1035 (N_1035,N_600,N_721);
nand U1036 (N_1036,N_914,N_903);
and U1037 (N_1037,N_882,N_992);
or U1038 (N_1038,N_978,N_956);
nor U1039 (N_1039,N_729,N_990);
or U1040 (N_1040,N_754,N_826);
and U1041 (N_1041,N_980,N_925);
nor U1042 (N_1042,N_612,N_686);
xnor U1043 (N_1043,N_934,N_834);
and U1044 (N_1044,N_790,N_818);
nand U1045 (N_1045,N_501,N_549);
or U1046 (N_1046,N_710,N_552);
xnor U1047 (N_1047,N_530,N_712);
nand U1048 (N_1048,N_811,N_794);
xor U1049 (N_1049,N_989,N_555);
and U1050 (N_1050,N_809,N_731);
nor U1051 (N_1051,N_920,N_594);
or U1052 (N_1052,N_911,N_588);
or U1053 (N_1053,N_706,N_520);
or U1054 (N_1054,N_582,N_595);
nand U1055 (N_1055,N_639,N_966);
and U1056 (N_1056,N_539,N_695);
or U1057 (N_1057,N_959,N_718);
and U1058 (N_1058,N_755,N_858);
and U1059 (N_1059,N_740,N_558);
nor U1060 (N_1060,N_546,N_551);
or U1061 (N_1061,N_732,N_608);
nand U1062 (N_1062,N_556,N_849);
nor U1063 (N_1063,N_527,N_509);
and U1064 (N_1064,N_757,N_696);
or U1065 (N_1065,N_843,N_694);
nor U1066 (N_1066,N_940,N_548);
nor U1067 (N_1067,N_802,N_532);
and U1068 (N_1068,N_873,N_540);
nand U1069 (N_1069,N_524,N_775);
and U1070 (N_1070,N_566,N_879);
nor U1071 (N_1071,N_708,N_777);
nor U1072 (N_1072,N_917,N_773);
and U1073 (N_1073,N_921,N_567);
and U1074 (N_1074,N_954,N_835);
and U1075 (N_1075,N_577,N_991);
xnor U1076 (N_1076,N_942,N_620);
or U1077 (N_1077,N_512,N_625);
nor U1078 (N_1078,N_678,N_711);
xor U1079 (N_1079,N_827,N_653);
nor U1080 (N_1080,N_709,N_614);
nor U1081 (N_1081,N_517,N_650);
xor U1082 (N_1082,N_967,N_519);
nor U1083 (N_1083,N_675,N_788);
nand U1084 (N_1084,N_930,N_671);
xnor U1085 (N_1085,N_610,N_964);
or U1086 (N_1086,N_889,N_943);
or U1087 (N_1087,N_621,N_725);
or U1088 (N_1088,N_869,N_592);
xor U1089 (N_1089,N_960,N_839);
or U1090 (N_1090,N_971,N_803);
xnor U1091 (N_1091,N_598,N_738);
or U1092 (N_1092,N_851,N_918);
nand U1093 (N_1093,N_975,N_601);
or U1094 (N_1094,N_717,N_937);
nand U1095 (N_1095,N_660,N_557);
xor U1096 (N_1096,N_627,N_605);
and U1097 (N_1097,N_502,N_850);
nand U1098 (N_1098,N_783,N_953);
nor U1099 (N_1099,N_840,N_974);
and U1100 (N_1100,N_714,N_507);
nor U1101 (N_1101,N_945,N_547);
and U1102 (N_1102,N_923,N_899);
nand U1103 (N_1103,N_531,N_973);
nor U1104 (N_1104,N_506,N_801);
and U1105 (N_1105,N_907,N_968);
nor U1106 (N_1106,N_813,N_970);
and U1107 (N_1107,N_618,N_946);
nor U1108 (N_1108,N_875,N_939);
or U1109 (N_1109,N_707,N_915);
nand U1110 (N_1110,N_815,N_886);
nor U1111 (N_1111,N_680,N_893);
or U1112 (N_1112,N_513,N_947);
nor U1113 (N_1113,N_822,N_673);
and U1114 (N_1114,N_749,N_584);
nand U1115 (N_1115,N_963,N_838);
and U1116 (N_1116,N_744,N_629);
nor U1117 (N_1117,N_845,N_534);
nor U1118 (N_1118,N_833,N_735);
nor U1119 (N_1119,N_586,N_863);
or U1120 (N_1120,N_760,N_900);
nor U1121 (N_1121,N_615,N_791);
and U1122 (N_1122,N_910,N_753);
and U1123 (N_1123,N_571,N_578);
nand U1124 (N_1124,N_994,N_972);
nor U1125 (N_1125,N_844,N_935);
nand U1126 (N_1126,N_572,N_624);
nor U1127 (N_1127,N_983,N_764);
or U1128 (N_1128,N_856,N_814);
or U1129 (N_1129,N_871,N_933);
nand U1130 (N_1130,N_569,N_737);
nand U1131 (N_1131,N_593,N_585);
and U1132 (N_1132,N_836,N_562);
and U1133 (N_1133,N_948,N_580);
or U1134 (N_1134,N_768,N_500);
nor U1135 (N_1135,N_800,N_529);
or U1136 (N_1136,N_736,N_542);
or U1137 (N_1137,N_928,N_602);
and U1138 (N_1138,N_689,N_656);
nand U1139 (N_1139,N_884,N_719);
xnor U1140 (N_1140,N_996,N_817);
or U1141 (N_1141,N_846,N_784);
or U1142 (N_1142,N_636,N_628);
and U1143 (N_1143,N_604,N_533);
xor U1144 (N_1144,N_976,N_763);
or U1145 (N_1145,N_638,N_961);
and U1146 (N_1146,N_831,N_526);
or U1147 (N_1147,N_797,N_703);
xor U1148 (N_1148,N_672,N_929);
xnor U1149 (N_1149,N_944,N_952);
and U1150 (N_1150,N_758,N_722);
or U1151 (N_1151,N_919,N_924);
nand U1152 (N_1152,N_560,N_544);
nand U1153 (N_1153,N_668,N_778);
or U1154 (N_1154,N_829,N_774);
nor U1155 (N_1155,N_649,N_870);
nand U1156 (N_1156,N_824,N_798);
or U1157 (N_1157,N_581,N_787);
nor U1158 (N_1158,N_859,N_525);
nand U1159 (N_1159,N_922,N_563);
or U1160 (N_1160,N_635,N_739);
xnor U1161 (N_1161,N_698,N_880);
or U1162 (N_1162,N_848,N_759);
and U1163 (N_1163,N_677,N_842);
nor U1164 (N_1164,N_564,N_664);
nor U1165 (N_1165,N_887,N_958);
nand U1166 (N_1166,N_704,N_908);
nor U1167 (N_1167,N_646,N_510);
or U1168 (N_1168,N_662,N_634);
and U1169 (N_1169,N_913,N_561);
and U1170 (N_1170,N_637,N_765);
nor U1171 (N_1171,N_866,N_626);
nand U1172 (N_1172,N_613,N_857);
and U1173 (N_1173,N_515,N_715);
or U1174 (N_1174,N_941,N_693);
and U1175 (N_1175,N_568,N_878);
or U1176 (N_1176,N_657,N_734);
and U1177 (N_1177,N_607,N_619);
nand U1178 (N_1178,N_936,N_796);
nand U1179 (N_1179,N_587,N_508);
xnor U1180 (N_1180,N_617,N_852);
and U1181 (N_1181,N_832,N_955);
and U1182 (N_1182,N_505,N_747);
and U1183 (N_1183,N_772,N_891);
nor U1184 (N_1184,N_511,N_828);
or U1185 (N_1185,N_579,N_820);
and U1186 (N_1186,N_647,N_799);
nand U1187 (N_1187,N_687,N_590);
and U1188 (N_1188,N_733,N_769);
or U1189 (N_1189,N_825,N_576);
or U1190 (N_1190,N_905,N_885);
xnor U1191 (N_1191,N_984,N_720);
or U1192 (N_1192,N_682,N_565);
and U1193 (N_1193,N_741,N_808);
nand U1194 (N_1194,N_805,N_697);
xnor U1195 (N_1195,N_589,N_535);
nand U1196 (N_1196,N_645,N_609);
or U1197 (N_1197,N_745,N_904);
and U1198 (N_1198,N_793,N_541);
nor U1199 (N_1199,N_898,N_841);
nand U1200 (N_1200,N_909,N_536);
or U1201 (N_1201,N_782,N_861);
and U1202 (N_1202,N_690,N_931);
xor U1203 (N_1203,N_545,N_776);
xor U1204 (N_1204,N_553,N_713);
nand U1205 (N_1205,N_993,N_746);
nor U1206 (N_1206,N_716,N_670);
nand U1207 (N_1207,N_631,N_837);
xnor U1208 (N_1208,N_591,N_537);
and U1209 (N_1209,N_730,N_916);
and U1210 (N_1210,N_897,N_688);
xnor U1211 (N_1211,N_503,N_894);
nand U1212 (N_1212,N_810,N_756);
xor U1213 (N_1213,N_902,N_766);
nand U1214 (N_1214,N_816,N_632);
nand U1215 (N_1215,N_606,N_633);
nand U1216 (N_1216,N_864,N_819);
and U1217 (N_1217,N_830,N_641);
nor U1218 (N_1218,N_743,N_965);
nand U1219 (N_1219,N_521,N_726);
and U1220 (N_1220,N_665,N_888);
nand U1221 (N_1221,N_699,N_806);
nand U1222 (N_1222,N_603,N_727);
and U1223 (N_1223,N_648,N_847);
or U1224 (N_1224,N_644,N_807);
nor U1225 (N_1225,N_883,N_795);
and U1226 (N_1226,N_522,N_658);
nor U1227 (N_1227,N_998,N_651);
or U1228 (N_1228,N_912,N_868);
nor U1229 (N_1229,N_623,N_705);
or U1230 (N_1230,N_724,N_667);
or U1231 (N_1231,N_596,N_999);
nand U1232 (N_1232,N_761,N_785);
and U1233 (N_1233,N_652,N_876);
xnor U1234 (N_1234,N_681,N_616);
nand U1235 (N_1235,N_938,N_877);
or U1236 (N_1236,N_528,N_881);
and U1237 (N_1237,N_987,N_669);
nor U1238 (N_1238,N_872,N_865);
or U1239 (N_1239,N_979,N_751);
nor U1240 (N_1240,N_654,N_702);
and U1241 (N_1241,N_683,N_504);
xnor U1242 (N_1242,N_573,N_611);
nand U1243 (N_1243,N_896,N_892);
or U1244 (N_1244,N_728,N_516);
or U1245 (N_1245,N_786,N_692);
or U1246 (N_1246,N_997,N_679);
or U1247 (N_1247,N_867,N_575);
or U1248 (N_1248,N_750,N_951);
xor U1249 (N_1249,N_543,N_518);
xnor U1250 (N_1250,N_760,N_514);
or U1251 (N_1251,N_566,N_939);
and U1252 (N_1252,N_939,N_967);
nor U1253 (N_1253,N_833,N_898);
nand U1254 (N_1254,N_602,N_872);
nand U1255 (N_1255,N_615,N_793);
xor U1256 (N_1256,N_869,N_788);
nand U1257 (N_1257,N_923,N_533);
and U1258 (N_1258,N_595,N_586);
xnor U1259 (N_1259,N_983,N_661);
nor U1260 (N_1260,N_525,N_596);
nand U1261 (N_1261,N_920,N_936);
or U1262 (N_1262,N_868,N_515);
nand U1263 (N_1263,N_835,N_873);
or U1264 (N_1264,N_552,N_598);
nand U1265 (N_1265,N_640,N_709);
nand U1266 (N_1266,N_827,N_591);
and U1267 (N_1267,N_521,N_741);
xnor U1268 (N_1268,N_627,N_690);
nand U1269 (N_1269,N_697,N_940);
and U1270 (N_1270,N_982,N_837);
nand U1271 (N_1271,N_656,N_855);
or U1272 (N_1272,N_590,N_790);
and U1273 (N_1273,N_885,N_730);
or U1274 (N_1274,N_523,N_948);
nand U1275 (N_1275,N_554,N_581);
nor U1276 (N_1276,N_887,N_601);
nor U1277 (N_1277,N_675,N_912);
and U1278 (N_1278,N_503,N_714);
xnor U1279 (N_1279,N_910,N_663);
nand U1280 (N_1280,N_578,N_865);
nor U1281 (N_1281,N_752,N_650);
nand U1282 (N_1282,N_740,N_653);
nand U1283 (N_1283,N_765,N_693);
or U1284 (N_1284,N_711,N_886);
and U1285 (N_1285,N_886,N_882);
nor U1286 (N_1286,N_832,N_924);
and U1287 (N_1287,N_761,N_777);
nand U1288 (N_1288,N_515,N_635);
nor U1289 (N_1289,N_530,N_848);
and U1290 (N_1290,N_853,N_697);
nand U1291 (N_1291,N_873,N_866);
and U1292 (N_1292,N_779,N_522);
and U1293 (N_1293,N_515,N_814);
nor U1294 (N_1294,N_715,N_824);
nor U1295 (N_1295,N_861,N_942);
nand U1296 (N_1296,N_556,N_676);
nand U1297 (N_1297,N_607,N_602);
and U1298 (N_1298,N_722,N_516);
nor U1299 (N_1299,N_808,N_913);
and U1300 (N_1300,N_588,N_797);
and U1301 (N_1301,N_866,N_823);
or U1302 (N_1302,N_886,N_562);
nand U1303 (N_1303,N_796,N_848);
nand U1304 (N_1304,N_654,N_951);
or U1305 (N_1305,N_532,N_514);
and U1306 (N_1306,N_947,N_776);
nand U1307 (N_1307,N_524,N_699);
xor U1308 (N_1308,N_648,N_694);
and U1309 (N_1309,N_793,N_773);
and U1310 (N_1310,N_863,N_669);
and U1311 (N_1311,N_527,N_518);
nand U1312 (N_1312,N_529,N_706);
and U1313 (N_1313,N_838,N_832);
and U1314 (N_1314,N_509,N_952);
nor U1315 (N_1315,N_857,N_633);
xnor U1316 (N_1316,N_771,N_830);
and U1317 (N_1317,N_862,N_573);
nand U1318 (N_1318,N_714,N_727);
nand U1319 (N_1319,N_657,N_707);
and U1320 (N_1320,N_952,N_723);
or U1321 (N_1321,N_519,N_964);
nand U1322 (N_1322,N_572,N_701);
nand U1323 (N_1323,N_824,N_705);
nor U1324 (N_1324,N_578,N_596);
nor U1325 (N_1325,N_548,N_556);
and U1326 (N_1326,N_619,N_739);
or U1327 (N_1327,N_960,N_615);
nor U1328 (N_1328,N_504,N_766);
xor U1329 (N_1329,N_614,N_904);
or U1330 (N_1330,N_839,N_658);
and U1331 (N_1331,N_984,N_741);
nor U1332 (N_1332,N_582,N_807);
and U1333 (N_1333,N_897,N_877);
and U1334 (N_1334,N_564,N_504);
nand U1335 (N_1335,N_948,N_612);
or U1336 (N_1336,N_524,N_756);
and U1337 (N_1337,N_892,N_971);
or U1338 (N_1338,N_668,N_553);
nand U1339 (N_1339,N_892,N_853);
nand U1340 (N_1340,N_784,N_955);
or U1341 (N_1341,N_854,N_989);
or U1342 (N_1342,N_619,N_793);
and U1343 (N_1343,N_586,N_991);
or U1344 (N_1344,N_680,N_854);
and U1345 (N_1345,N_505,N_954);
xor U1346 (N_1346,N_875,N_629);
and U1347 (N_1347,N_611,N_629);
nor U1348 (N_1348,N_866,N_822);
or U1349 (N_1349,N_550,N_723);
or U1350 (N_1350,N_829,N_627);
nor U1351 (N_1351,N_678,N_510);
nor U1352 (N_1352,N_911,N_979);
nor U1353 (N_1353,N_816,N_703);
nand U1354 (N_1354,N_536,N_700);
and U1355 (N_1355,N_716,N_971);
nand U1356 (N_1356,N_835,N_596);
or U1357 (N_1357,N_744,N_704);
or U1358 (N_1358,N_671,N_543);
and U1359 (N_1359,N_686,N_683);
nor U1360 (N_1360,N_684,N_548);
nand U1361 (N_1361,N_730,N_672);
nand U1362 (N_1362,N_616,N_514);
xnor U1363 (N_1363,N_775,N_508);
and U1364 (N_1364,N_594,N_988);
nand U1365 (N_1365,N_938,N_905);
and U1366 (N_1366,N_587,N_817);
nand U1367 (N_1367,N_965,N_603);
or U1368 (N_1368,N_543,N_801);
or U1369 (N_1369,N_659,N_887);
and U1370 (N_1370,N_607,N_659);
and U1371 (N_1371,N_867,N_910);
nand U1372 (N_1372,N_545,N_684);
or U1373 (N_1373,N_774,N_818);
nor U1374 (N_1374,N_549,N_766);
xnor U1375 (N_1375,N_713,N_708);
nand U1376 (N_1376,N_659,N_563);
nand U1377 (N_1377,N_638,N_573);
and U1378 (N_1378,N_707,N_946);
or U1379 (N_1379,N_551,N_836);
and U1380 (N_1380,N_701,N_885);
and U1381 (N_1381,N_873,N_871);
nor U1382 (N_1382,N_528,N_783);
and U1383 (N_1383,N_794,N_928);
nor U1384 (N_1384,N_702,N_766);
nor U1385 (N_1385,N_923,N_888);
or U1386 (N_1386,N_754,N_907);
or U1387 (N_1387,N_621,N_606);
nor U1388 (N_1388,N_576,N_717);
xor U1389 (N_1389,N_672,N_964);
and U1390 (N_1390,N_657,N_726);
or U1391 (N_1391,N_642,N_946);
or U1392 (N_1392,N_617,N_902);
or U1393 (N_1393,N_923,N_790);
or U1394 (N_1394,N_610,N_998);
nand U1395 (N_1395,N_835,N_625);
nor U1396 (N_1396,N_551,N_533);
or U1397 (N_1397,N_561,N_523);
nand U1398 (N_1398,N_714,N_838);
or U1399 (N_1399,N_825,N_651);
xor U1400 (N_1400,N_621,N_539);
nor U1401 (N_1401,N_586,N_701);
nor U1402 (N_1402,N_853,N_855);
nand U1403 (N_1403,N_801,N_807);
nor U1404 (N_1404,N_664,N_972);
nor U1405 (N_1405,N_780,N_576);
or U1406 (N_1406,N_529,N_540);
nand U1407 (N_1407,N_897,N_808);
nor U1408 (N_1408,N_753,N_765);
nand U1409 (N_1409,N_821,N_836);
or U1410 (N_1410,N_945,N_660);
and U1411 (N_1411,N_629,N_556);
or U1412 (N_1412,N_545,N_623);
and U1413 (N_1413,N_640,N_814);
or U1414 (N_1414,N_804,N_511);
xor U1415 (N_1415,N_638,N_618);
and U1416 (N_1416,N_775,N_996);
nand U1417 (N_1417,N_531,N_826);
or U1418 (N_1418,N_528,N_576);
nor U1419 (N_1419,N_664,N_876);
or U1420 (N_1420,N_674,N_613);
nor U1421 (N_1421,N_784,N_622);
nand U1422 (N_1422,N_717,N_951);
and U1423 (N_1423,N_772,N_622);
nand U1424 (N_1424,N_726,N_747);
and U1425 (N_1425,N_786,N_782);
xnor U1426 (N_1426,N_924,N_721);
nor U1427 (N_1427,N_997,N_505);
nand U1428 (N_1428,N_588,N_675);
and U1429 (N_1429,N_763,N_932);
nand U1430 (N_1430,N_857,N_814);
nand U1431 (N_1431,N_615,N_693);
or U1432 (N_1432,N_944,N_644);
nand U1433 (N_1433,N_727,N_586);
nor U1434 (N_1434,N_912,N_983);
nand U1435 (N_1435,N_822,N_639);
and U1436 (N_1436,N_721,N_702);
or U1437 (N_1437,N_984,N_647);
and U1438 (N_1438,N_654,N_603);
nand U1439 (N_1439,N_767,N_770);
and U1440 (N_1440,N_703,N_880);
nand U1441 (N_1441,N_789,N_523);
and U1442 (N_1442,N_826,N_615);
or U1443 (N_1443,N_604,N_677);
or U1444 (N_1444,N_524,N_731);
xnor U1445 (N_1445,N_666,N_897);
and U1446 (N_1446,N_899,N_827);
nand U1447 (N_1447,N_878,N_884);
or U1448 (N_1448,N_670,N_614);
or U1449 (N_1449,N_905,N_775);
nor U1450 (N_1450,N_943,N_660);
and U1451 (N_1451,N_543,N_951);
or U1452 (N_1452,N_794,N_647);
xnor U1453 (N_1453,N_605,N_513);
or U1454 (N_1454,N_950,N_699);
xnor U1455 (N_1455,N_614,N_787);
and U1456 (N_1456,N_945,N_911);
nor U1457 (N_1457,N_642,N_752);
or U1458 (N_1458,N_694,N_509);
and U1459 (N_1459,N_810,N_825);
and U1460 (N_1460,N_832,N_987);
or U1461 (N_1461,N_739,N_751);
nor U1462 (N_1462,N_570,N_505);
nand U1463 (N_1463,N_657,N_751);
nor U1464 (N_1464,N_612,N_559);
and U1465 (N_1465,N_663,N_706);
nand U1466 (N_1466,N_869,N_722);
nand U1467 (N_1467,N_727,N_638);
nand U1468 (N_1468,N_523,N_907);
or U1469 (N_1469,N_548,N_841);
and U1470 (N_1470,N_590,N_845);
and U1471 (N_1471,N_769,N_750);
nand U1472 (N_1472,N_578,N_823);
nand U1473 (N_1473,N_586,N_542);
or U1474 (N_1474,N_930,N_808);
nor U1475 (N_1475,N_513,N_747);
or U1476 (N_1476,N_611,N_795);
nor U1477 (N_1477,N_556,N_534);
nor U1478 (N_1478,N_739,N_631);
or U1479 (N_1479,N_788,N_889);
or U1480 (N_1480,N_707,N_819);
nor U1481 (N_1481,N_830,N_904);
or U1482 (N_1482,N_677,N_596);
nand U1483 (N_1483,N_602,N_936);
and U1484 (N_1484,N_542,N_541);
nand U1485 (N_1485,N_771,N_848);
nand U1486 (N_1486,N_628,N_722);
nor U1487 (N_1487,N_546,N_963);
nand U1488 (N_1488,N_733,N_770);
or U1489 (N_1489,N_919,N_914);
or U1490 (N_1490,N_748,N_525);
nand U1491 (N_1491,N_858,N_988);
and U1492 (N_1492,N_612,N_616);
and U1493 (N_1493,N_724,N_816);
or U1494 (N_1494,N_790,N_707);
and U1495 (N_1495,N_585,N_951);
and U1496 (N_1496,N_512,N_854);
nand U1497 (N_1497,N_780,N_544);
nor U1498 (N_1498,N_566,N_796);
nand U1499 (N_1499,N_904,N_699);
nor U1500 (N_1500,N_1468,N_1160);
or U1501 (N_1501,N_1206,N_1432);
xor U1502 (N_1502,N_1475,N_1163);
or U1503 (N_1503,N_1223,N_1312);
nor U1504 (N_1504,N_1327,N_1042);
nor U1505 (N_1505,N_1283,N_1496);
and U1506 (N_1506,N_1458,N_1473);
or U1507 (N_1507,N_1193,N_1478);
or U1508 (N_1508,N_1032,N_1118);
nor U1509 (N_1509,N_1176,N_1197);
or U1510 (N_1510,N_1221,N_1095);
nand U1511 (N_1511,N_1112,N_1009);
nand U1512 (N_1512,N_1040,N_1460);
or U1513 (N_1513,N_1214,N_1339);
xnor U1514 (N_1514,N_1434,N_1436);
and U1515 (N_1515,N_1486,N_1463);
xor U1516 (N_1516,N_1471,N_1162);
and U1517 (N_1517,N_1018,N_1004);
nor U1518 (N_1518,N_1067,N_1236);
or U1519 (N_1519,N_1405,N_1235);
and U1520 (N_1520,N_1244,N_1003);
nor U1521 (N_1521,N_1282,N_1420);
nand U1522 (N_1522,N_1166,N_1355);
and U1523 (N_1523,N_1170,N_1093);
or U1524 (N_1524,N_1487,N_1179);
or U1525 (N_1525,N_1256,N_1451);
nor U1526 (N_1526,N_1153,N_1185);
or U1527 (N_1527,N_1255,N_1302);
nand U1528 (N_1528,N_1378,N_1398);
nor U1529 (N_1529,N_1292,N_1041);
nor U1530 (N_1530,N_1148,N_1469);
nand U1531 (N_1531,N_1152,N_1479);
nand U1532 (N_1532,N_1109,N_1051);
nand U1533 (N_1533,N_1328,N_1135);
nor U1534 (N_1534,N_1181,N_1280);
and U1535 (N_1535,N_1344,N_1300);
or U1536 (N_1536,N_1326,N_1353);
nor U1537 (N_1537,N_1034,N_1357);
nor U1538 (N_1538,N_1251,N_1400);
nand U1539 (N_1539,N_1417,N_1309);
or U1540 (N_1540,N_1284,N_1060);
or U1541 (N_1541,N_1317,N_1299);
and U1542 (N_1542,N_1015,N_1036);
or U1543 (N_1543,N_1443,N_1472);
and U1544 (N_1544,N_1094,N_1026);
nor U1545 (N_1545,N_1329,N_1159);
or U1546 (N_1546,N_1363,N_1184);
nor U1547 (N_1547,N_1401,N_1037);
nand U1548 (N_1548,N_1202,N_1371);
nand U1549 (N_1549,N_1105,N_1254);
xnor U1550 (N_1550,N_1011,N_1272);
nand U1551 (N_1551,N_1158,N_1424);
and U1552 (N_1552,N_1416,N_1389);
xnor U1553 (N_1553,N_1055,N_1406);
nor U1554 (N_1554,N_1481,N_1117);
or U1555 (N_1555,N_1354,N_1133);
and U1556 (N_1556,N_1440,N_1310);
and U1557 (N_1557,N_1392,N_1273);
nand U1558 (N_1558,N_1279,N_1196);
and U1559 (N_1559,N_1495,N_1446);
nand U1560 (N_1560,N_1183,N_1232);
or U1561 (N_1561,N_1080,N_1258);
nand U1562 (N_1562,N_1488,N_1409);
nor U1563 (N_1563,N_1492,N_1340);
nor U1564 (N_1564,N_1088,N_1275);
nand U1565 (N_1565,N_1228,N_1229);
or U1566 (N_1566,N_1342,N_1019);
nor U1567 (N_1567,N_1367,N_1035);
nand U1568 (N_1568,N_1048,N_1107);
nor U1569 (N_1569,N_1000,N_1386);
and U1570 (N_1570,N_1143,N_1316);
nor U1571 (N_1571,N_1125,N_1351);
nand U1572 (N_1572,N_1347,N_1399);
or U1573 (N_1573,N_1305,N_1429);
nand U1574 (N_1574,N_1233,N_1455);
and U1575 (N_1575,N_1209,N_1084);
and U1576 (N_1576,N_1394,N_1022);
nor U1577 (N_1577,N_1053,N_1174);
nand U1578 (N_1578,N_1127,N_1470);
nor U1579 (N_1579,N_1447,N_1192);
nand U1580 (N_1580,N_1155,N_1203);
nand U1581 (N_1581,N_1027,N_1308);
and U1582 (N_1582,N_1226,N_1418);
or U1583 (N_1583,N_1033,N_1131);
nor U1584 (N_1584,N_1039,N_1016);
nor U1585 (N_1585,N_1121,N_1047);
nor U1586 (N_1586,N_1427,N_1146);
or U1587 (N_1587,N_1006,N_1360);
nand U1588 (N_1588,N_1139,N_1090);
and U1589 (N_1589,N_1380,N_1172);
nand U1590 (N_1590,N_1144,N_1007);
and U1591 (N_1591,N_1274,N_1017);
nand U1592 (N_1592,N_1259,N_1165);
nand U1593 (N_1593,N_1407,N_1207);
or U1594 (N_1594,N_1356,N_1178);
and U1595 (N_1595,N_1384,N_1066);
nor U1596 (N_1596,N_1277,N_1349);
or U1597 (N_1597,N_1412,N_1480);
xnor U1598 (N_1598,N_1129,N_1276);
or U1599 (N_1599,N_1134,N_1397);
or U1600 (N_1600,N_1059,N_1457);
or U1601 (N_1601,N_1387,N_1111);
nand U1602 (N_1602,N_1425,N_1194);
or U1603 (N_1603,N_1257,N_1477);
or U1604 (N_1604,N_1270,N_1157);
or U1605 (N_1605,N_1334,N_1122);
and U1606 (N_1606,N_1456,N_1322);
nand U1607 (N_1607,N_1149,N_1216);
or U1608 (N_1608,N_1402,N_1079);
and U1609 (N_1609,N_1227,N_1439);
or U1610 (N_1610,N_1426,N_1001);
nor U1611 (N_1611,N_1150,N_1438);
xnor U1612 (N_1612,N_1391,N_1023);
nand U1613 (N_1613,N_1494,N_1288);
nor U1614 (N_1614,N_1119,N_1187);
nand U1615 (N_1615,N_1045,N_1190);
xnor U1616 (N_1616,N_1373,N_1199);
nor U1617 (N_1617,N_1430,N_1415);
nand U1618 (N_1618,N_1433,N_1465);
xnor U1619 (N_1619,N_1303,N_1106);
nor U1620 (N_1620,N_1046,N_1365);
and U1621 (N_1621,N_1167,N_1422);
nand U1622 (N_1622,N_1115,N_1361);
nor U1623 (N_1623,N_1195,N_1114);
or U1624 (N_1624,N_1291,N_1466);
nand U1625 (N_1625,N_1382,N_1285);
or U1626 (N_1626,N_1081,N_1078);
or U1627 (N_1627,N_1331,N_1219);
nand U1628 (N_1628,N_1267,N_1151);
and U1629 (N_1629,N_1491,N_1213);
or U1630 (N_1630,N_1497,N_1083);
or U1631 (N_1631,N_1164,N_1301);
nor U1632 (N_1632,N_1250,N_1091);
and U1633 (N_1633,N_1321,N_1028);
nand U1634 (N_1634,N_1385,N_1364);
and U1635 (N_1635,N_1147,N_1177);
xor U1636 (N_1636,N_1225,N_1029);
or U1637 (N_1637,N_1087,N_1012);
or U1638 (N_1638,N_1444,N_1345);
nor U1639 (N_1639,N_1061,N_1021);
or U1640 (N_1640,N_1222,N_1484);
xor U1641 (N_1641,N_1411,N_1493);
and U1642 (N_1642,N_1377,N_1057);
nor U1643 (N_1643,N_1205,N_1390);
nand U1644 (N_1644,N_1348,N_1393);
or U1645 (N_1645,N_1437,N_1315);
or U1646 (N_1646,N_1182,N_1242);
xor U1647 (N_1647,N_1379,N_1008);
nand U1648 (N_1648,N_1108,N_1099);
or U1649 (N_1649,N_1063,N_1375);
nand U1650 (N_1650,N_1352,N_1287);
and U1651 (N_1651,N_1137,N_1245);
nor U1652 (N_1652,N_1188,N_1110);
and U1653 (N_1653,N_1096,N_1086);
nor U1654 (N_1654,N_1335,N_1064);
nand U1655 (N_1655,N_1138,N_1498);
nand U1656 (N_1656,N_1201,N_1189);
nand U1657 (N_1657,N_1230,N_1020);
xnor U1658 (N_1658,N_1089,N_1453);
nand U1659 (N_1659,N_1388,N_1013);
xnor U1660 (N_1660,N_1281,N_1265);
nor U1661 (N_1661,N_1298,N_1333);
and U1662 (N_1662,N_1269,N_1113);
or U1663 (N_1663,N_1218,N_1123);
nor U1664 (N_1664,N_1075,N_1318);
nor U1665 (N_1665,N_1168,N_1474);
nor U1666 (N_1666,N_1266,N_1445);
xor U1667 (N_1667,N_1161,N_1056);
and U1668 (N_1668,N_1031,N_1210);
xnor U1669 (N_1669,N_1467,N_1294);
xnor U1670 (N_1670,N_1296,N_1224);
or U1671 (N_1671,N_1337,N_1459);
or U1672 (N_1672,N_1068,N_1076);
nor U1673 (N_1673,N_1208,N_1376);
and U1674 (N_1674,N_1128,N_1103);
and U1675 (N_1675,N_1180,N_1154);
or U1676 (N_1676,N_1464,N_1005);
or U1677 (N_1677,N_1263,N_1220);
or U1678 (N_1678,N_1449,N_1239);
and U1679 (N_1679,N_1304,N_1419);
and U1680 (N_1680,N_1307,N_1198);
nor U1681 (N_1681,N_1332,N_1359);
nor U1682 (N_1682,N_1290,N_1396);
nand U1683 (N_1683,N_1217,N_1191);
nand U1684 (N_1684,N_1362,N_1383);
nor U1685 (N_1685,N_1071,N_1241);
and U1686 (N_1686,N_1140,N_1014);
nand U1687 (N_1687,N_1408,N_1132);
nand U1688 (N_1688,N_1413,N_1052);
nand U1689 (N_1689,N_1098,N_1104);
and U1690 (N_1690,N_1325,N_1072);
or U1691 (N_1691,N_1142,N_1476);
xnor U1692 (N_1692,N_1136,N_1238);
or U1693 (N_1693,N_1002,N_1025);
or U1694 (N_1694,N_1330,N_1489);
or U1695 (N_1695,N_1435,N_1421);
or U1696 (N_1696,N_1246,N_1243);
or U1697 (N_1697,N_1431,N_1278);
nand U1698 (N_1698,N_1452,N_1441);
or U1699 (N_1699,N_1271,N_1404);
or U1700 (N_1700,N_1204,N_1073);
or U1701 (N_1701,N_1070,N_1065);
nor U1702 (N_1702,N_1249,N_1030);
nor U1703 (N_1703,N_1043,N_1101);
and U1704 (N_1704,N_1346,N_1324);
or U1705 (N_1705,N_1343,N_1314);
nand U1706 (N_1706,N_1252,N_1490);
nor U1707 (N_1707,N_1049,N_1295);
and U1708 (N_1708,N_1499,N_1141);
nand U1709 (N_1709,N_1058,N_1366);
xnor U1710 (N_1710,N_1336,N_1050);
and U1711 (N_1711,N_1323,N_1211);
nor U1712 (N_1712,N_1293,N_1024);
nand U1713 (N_1713,N_1381,N_1403);
and U1714 (N_1714,N_1092,N_1423);
and U1715 (N_1715,N_1320,N_1260);
or U1716 (N_1716,N_1074,N_1173);
nor U1717 (N_1717,N_1261,N_1461);
and U1718 (N_1718,N_1062,N_1253);
nor U1719 (N_1719,N_1169,N_1085);
and U1720 (N_1720,N_1313,N_1448);
nand U1721 (N_1721,N_1462,N_1044);
or U1722 (N_1722,N_1395,N_1454);
or U1723 (N_1723,N_1297,N_1156);
nand U1724 (N_1724,N_1350,N_1097);
and U1725 (N_1725,N_1311,N_1120);
nand U1726 (N_1726,N_1200,N_1186);
nand U1727 (N_1727,N_1240,N_1082);
nor U1728 (N_1728,N_1130,N_1171);
nor U1729 (N_1729,N_1374,N_1102);
nand U1730 (N_1730,N_1450,N_1234);
nor U1731 (N_1731,N_1483,N_1116);
nand U1732 (N_1732,N_1369,N_1077);
nand U1733 (N_1733,N_1126,N_1370);
or U1734 (N_1734,N_1485,N_1124);
or U1735 (N_1735,N_1248,N_1268);
and U1736 (N_1736,N_1231,N_1010);
nor U1737 (N_1737,N_1428,N_1100);
nand U1738 (N_1738,N_1145,N_1368);
or U1739 (N_1739,N_1054,N_1286);
or U1740 (N_1740,N_1069,N_1338);
nand U1741 (N_1741,N_1442,N_1262);
nor U1742 (N_1742,N_1289,N_1414);
nor U1743 (N_1743,N_1319,N_1038);
nor U1744 (N_1744,N_1482,N_1264);
nor U1745 (N_1745,N_1212,N_1358);
nand U1746 (N_1746,N_1410,N_1372);
nor U1747 (N_1747,N_1237,N_1215);
or U1748 (N_1748,N_1175,N_1306);
and U1749 (N_1749,N_1341,N_1247);
nor U1750 (N_1750,N_1403,N_1108);
or U1751 (N_1751,N_1114,N_1120);
nor U1752 (N_1752,N_1448,N_1413);
nor U1753 (N_1753,N_1495,N_1314);
xor U1754 (N_1754,N_1426,N_1283);
and U1755 (N_1755,N_1419,N_1355);
or U1756 (N_1756,N_1471,N_1394);
nand U1757 (N_1757,N_1002,N_1367);
nor U1758 (N_1758,N_1207,N_1402);
nand U1759 (N_1759,N_1082,N_1097);
and U1760 (N_1760,N_1056,N_1163);
xor U1761 (N_1761,N_1382,N_1028);
nand U1762 (N_1762,N_1101,N_1204);
nand U1763 (N_1763,N_1057,N_1347);
nor U1764 (N_1764,N_1298,N_1133);
nand U1765 (N_1765,N_1113,N_1483);
or U1766 (N_1766,N_1024,N_1446);
and U1767 (N_1767,N_1140,N_1020);
xnor U1768 (N_1768,N_1036,N_1214);
nand U1769 (N_1769,N_1352,N_1265);
and U1770 (N_1770,N_1452,N_1386);
or U1771 (N_1771,N_1341,N_1265);
xnor U1772 (N_1772,N_1281,N_1200);
nand U1773 (N_1773,N_1423,N_1348);
nor U1774 (N_1774,N_1151,N_1291);
or U1775 (N_1775,N_1250,N_1338);
nand U1776 (N_1776,N_1261,N_1025);
and U1777 (N_1777,N_1111,N_1409);
and U1778 (N_1778,N_1331,N_1397);
nand U1779 (N_1779,N_1158,N_1369);
and U1780 (N_1780,N_1051,N_1135);
nor U1781 (N_1781,N_1230,N_1420);
nor U1782 (N_1782,N_1096,N_1288);
and U1783 (N_1783,N_1117,N_1428);
or U1784 (N_1784,N_1255,N_1269);
nor U1785 (N_1785,N_1490,N_1173);
xnor U1786 (N_1786,N_1037,N_1219);
nor U1787 (N_1787,N_1071,N_1495);
nor U1788 (N_1788,N_1351,N_1081);
nand U1789 (N_1789,N_1148,N_1307);
nand U1790 (N_1790,N_1291,N_1179);
xnor U1791 (N_1791,N_1004,N_1329);
and U1792 (N_1792,N_1429,N_1498);
nor U1793 (N_1793,N_1455,N_1411);
and U1794 (N_1794,N_1431,N_1399);
nor U1795 (N_1795,N_1043,N_1082);
and U1796 (N_1796,N_1053,N_1238);
nor U1797 (N_1797,N_1367,N_1397);
and U1798 (N_1798,N_1080,N_1306);
and U1799 (N_1799,N_1426,N_1468);
xnor U1800 (N_1800,N_1031,N_1117);
nor U1801 (N_1801,N_1487,N_1399);
and U1802 (N_1802,N_1241,N_1231);
nor U1803 (N_1803,N_1205,N_1129);
and U1804 (N_1804,N_1125,N_1186);
and U1805 (N_1805,N_1218,N_1306);
and U1806 (N_1806,N_1014,N_1419);
nand U1807 (N_1807,N_1187,N_1213);
and U1808 (N_1808,N_1177,N_1197);
nand U1809 (N_1809,N_1435,N_1307);
xor U1810 (N_1810,N_1099,N_1435);
nor U1811 (N_1811,N_1048,N_1457);
nand U1812 (N_1812,N_1135,N_1482);
nor U1813 (N_1813,N_1457,N_1091);
nand U1814 (N_1814,N_1274,N_1420);
or U1815 (N_1815,N_1098,N_1239);
or U1816 (N_1816,N_1291,N_1296);
nor U1817 (N_1817,N_1187,N_1156);
nor U1818 (N_1818,N_1070,N_1268);
or U1819 (N_1819,N_1078,N_1076);
and U1820 (N_1820,N_1428,N_1062);
or U1821 (N_1821,N_1233,N_1169);
nand U1822 (N_1822,N_1166,N_1203);
xnor U1823 (N_1823,N_1282,N_1201);
or U1824 (N_1824,N_1381,N_1308);
and U1825 (N_1825,N_1040,N_1148);
nor U1826 (N_1826,N_1249,N_1148);
or U1827 (N_1827,N_1461,N_1398);
nor U1828 (N_1828,N_1240,N_1122);
nand U1829 (N_1829,N_1040,N_1360);
or U1830 (N_1830,N_1336,N_1339);
nand U1831 (N_1831,N_1316,N_1364);
nand U1832 (N_1832,N_1361,N_1432);
and U1833 (N_1833,N_1427,N_1316);
nor U1834 (N_1834,N_1461,N_1334);
and U1835 (N_1835,N_1220,N_1365);
or U1836 (N_1836,N_1162,N_1354);
xor U1837 (N_1837,N_1307,N_1216);
xnor U1838 (N_1838,N_1036,N_1467);
or U1839 (N_1839,N_1107,N_1133);
and U1840 (N_1840,N_1098,N_1270);
and U1841 (N_1841,N_1467,N_1399);
nor U1842 (N_1842,N_1304,N_1031);
and U1843 (N_1843,N_1205,N_1176);
nand U1844 (N_1844,N_1000,N_1294);
nand U1845 (N_1845,N_1325,N_1429);
xor U1846 (N_1846,N_1411,N_1355);
and U1847 (N_1847,N_1065,N_1019);
or U1848 (N_1848,N_1326,N_1067);
nand U1849 (N_1849,N_1267,N_1287);
or U1850 (N_1850,N_1063,N_1260);
nand U1851 (N_1851,N_1132,N_1167);
or U1852 (N_1852,N_1018,N_1470);
or U1853 (N_1853,N_1030,N_1478);
nand U1854 (N_1854,N_1451,N_1145);
and U1855 (N_1855,N_1483,N_1209);
nor U1856 (N_1856,N_1440,N_1359);
nand U1857 (N_1857,N_1074,N_1491);
and U1858 (N_1858,N_1059,N_1331);
or U1859 (N_1859,N_1283,N_1219);
nor U1860 (N_1860,N_1249,N_1048);
nor U1861 (N_1861,N_1358,N_1241);
nor U1862 (N_1862,N_1050,N_1402);
and U1863 (N_1863,N_1422,N_1169);
nor U1864 (N_1864,N_1402,N_1491);
nand U1865 (N_1865,N_1239,N_1406);
and U1866 (N_1866,N_1203,N_1044);
nor U1867 (N_1867,N_1016,N_1327);
and U1868 (N_1868,N_1301,N_1238);
or U1869 (N_1869,N_1139,N_1362);
xor U1870 (N_1870,N_1172,N_1021);
or U1871 (N_1871,N_1035,N_1235);
or U1872 (N_1872,N_1010,N_1190);
nand U1873 (N_1873,N_1463,N_1250);
nor U1874 (N_1874,N_1034,N_1226);
or U1875 (N_1875,N_1224,N_1246);
or U1876 (N_1876,N_1205,N_1485);
nor U1877 (N_1877,N_1360,N_1289);
nor U1878 (N_1878,N_1391,N_1341);
nor U1879 (N_1879,N_1487,N_1356);
nor U1880 (N_1880,N_1379,N_1482);
xor U1881 (N_1881,N_1233,N_1198);
nor U1882 (N_1882,N_1397,N_1296);
nor U1883 (N_1883,N_1227,N_1006);
nor U1884 (N_1884,N_1458,N_1282);
and U1885 (N_1885,N_1182,N_1479);
and U1886 (N_1886,N_1072,N_1007);
nand U1887 (N_1887,N_1143,N_1016);
and U1888 (N_1888,N_1430,N_1479);
nand U1889 (N_1889,N_1135,N_1151);
and U1890 (N_1890,N_1423,N_1131);
or U1891 (N_1891,N_1173,N_1005);
and U1892 (N_1892,N_1280,N_1009);
or U1893 (N_1893,N_1388,N_1410);
nor U1894 (N_1894,N_1406,N_1259);
nand U1895 (N_1895,N_1406,N_1030);
nor U1896 (N_1896,N_1448,N_1165);
or U1897 (N_1897,N_1208,N_1483);
nand U1898 (N_1898,N_1432,N_1083);
nand U1899 (N_1899,N_1105,N_1115);
or U1900 (N_1900,N_1045,N_1178);
nor U1901 (N_1901,N_1126,N_1030);
nor U1902 (N_1902,N_1139,N_1489);
xor U1903 (N_1903,N_1322,N_1003);
nand U1904 (N_1904,N_1137,N_1405);
and U1905 (N_1905,N_1467,N_1042);
and U1906 (N_1906,N_1415,N_1312);
and U1907 (N_1907,N_1095,N_1017);
nor U1908 (N_1908,N_1258,N_1174);
or U1909 (N_1909,N_1261,N_1154);
or U1910 (N_1910,N_1120,N_1302);
nor U1911 (N_1911,N_1290,N_1441);
nor U1912 (N_1912,N_1296,N_1147);
nand U1913 (N_1913,N_1126,N_1377);
or U1914 (N_1914,N_1220,N_1024);
or U1915 (N_1915,N_1062,N_1225);
or U1916 (N_1916,N_1329,N_1388);
and U1917 (N_1917,N_1350,N_1241);
nand U1918 (N_1918,N_1463,N_1080);
or U1919 (N_1919,N_1402,N_1466);
xor U1920 (N_1920,N_1428,N_1196);
nor U1921 (N_1921,N_1047,N_1052);
nor U1922 (N_1922,N_1156,N_1071);
nand U1923 (N_1923,N_1020,N_1178);
and U1924 (N_1924,N_1215,N_1276);
nand U1925 (N_1925,N_1251,N_1176);
nor U1926 (N_1926,N_1372,N_1306);
nor U1927 (N_1927,N_1486,N_1108);
nand U1928 (N_1928,N_1166,N_1010);
nand U1929 (N_1929,N_1264,N_1307);
or U1930 (N_1930,N_1418,N_1343);
or U1931 (N_1931,N_1383,N_1312);
xnor U1932 (N_1932,N_1218,N_1001);
or U1933 (N_1933,N_1189,N_1403);
nand U1934 (N_1934,N_1204,N_1053);
nand U1935 (N_1935,N_1080,N_1303);
nor U1936 (N_1936,N_1015,N_1450);
or U1937 (N_1937,N_1210,N_1124);
and U1938 (N_1938,N_1322,N_1491);
xnor U1939 (N_1939,N_1160,N_1393);
nand U1940 (N_1940,N_1203,N_1426);
and U1941 (N_1941,N_1487,N_1443);
or U1942 (N_1942,N_1172,N_1243);
or U1943 (N_1943,N_1164,N_1233);
xnor U1944 (N_1944,N_1464,N_1149);
nor U1945 (N_1945,N_1136,N_1080);
nor U1946 (N_1946,N_1316,N_1006);
nor U1947 (N_1947,N_1039,N_1213);
nand U1948 (N_1948,N_1215,N_1415);
and U1949 (N_1949,N_1015,N_1211);
nor U1950 (N_1950,N_1066,N_1085);
and U1951 (N_1951,N_1020,N_1441);
xor U1952 (N_1952,N_1397,N_1352);
nand U1953 (N_1953,N_1012,N_1129);
nor U1954 (N_1954,N_1173,N_1236);
nor U1955 (N_1955,N_1446,N_1278);
nor U1956 (N_1956,N_1167,N_1220);
nor U1957 (N_1957,N_1149,N_1198);
or U1958 (N_1958,N_1414,N_1056);
or U1959 (N_1959,N_1449,N_1296);
and U1960 (N_1960,N_1128,N_1055);
nor U1961 (N_1961,N_1477,N_1157);
nor U1962 (N_1962,N_1283,N_1220);
and U1963 (N_1963,N_1331,N_1322);
xnor U1964 (N_1964,N_1462,N_1445);
nand U1965 (N_1965,N_1344,N_1452);
nand U1966 (N_1966,N_1017,N_1331);
nand U1967 (N_1967,N_1112,N_1463);
nand U1968 (N_1968,N_1351,N_1277);
xnor U1969 (N_1969,N_1314,N_1153);
and U1970 (N_1970,N_1276,N_1319);
nor U1971 (N_1971,N_1209,N_1355);
nand U1972 (N_1972,N_1321,N_1303);
or U1973 (N_1973,N_1230,N_1167);
nor U1974 (N_1974,N_1338,N_1429);
and U1975 (N_1975,N_1203,N_1093);
nand U1976 (N_1976,N_1449,N_1424);
or U1977 (N_1977,N_1332,N_1433);
or U1978 (N_1978,N_1405,N_1208);
and U1979 (N_1979,N_1436,N_1046);
nor U1980 (N_1980,N_1194,N_1003);
nor U1981 (N_1981,N_1249,N_1293);
and U1982 (N_1982,N_1382,N_1116);
nor U1983 (N_1983,N_1049,N_1252);
xor U1984 (N_1984,N_1087,N_1207);
xnor U1985 (N_1985,N_1395,N_1420);
xor U1986 (N_1986,N_1149,N_1471);
and U1987 (N_1987,N_1063,N_1166);
nor U1988 (N_1988,N_1308,N_1341);
nand U1989 (N_1989,N_1194,N_1375);
nor U1990 (N_1990,N_1215,N_1053);
xor U1991 (N_1991,N_1465,N_1283);
nor U1992 (N_1992,N_1159,N_1428);
and U1993 (N_1993,N_1085,N_1298);
or U1994 (N_1994,N_1427,N_1208);
and U1995 (N_1995,N_1039,N_1430);
nand U1996 (N_1996,N_1044,N_1216);
nor U1997 (N_1997,N_1047,N_1281);
and U1998 (N_1998,N_1383,N_1287);
and U1999 (N_1999,N_1262,N_1279);
and U2000 (N_2000,N_1823,N_1846);
and U2001 (N_2001,N_1540,N_1943);
and U2002 (N_2002,N_1580,N_1566);
nor U2003 (N_2003,N_1843,N_1639);
nor U2004 (N_2004,N_1537,N_1791);
or U2005 (N_2005,N_1856,N_1881);
or U2006 (N_2006,N_1552,N_1920);
xnor U2007 (N_2007,N_1502,N_1636);
xnor U2008 (N_2008,N_1896,N_1556);
xnor U2009 (N_2009,N_1780,N_1549);
or U2010 (N_2010,N_1532,N_1572);
and U2011 (N_2011,N_1974,N_1642);
nor U2012 (N_2012,N_1753,N_1965);
nand U2013 (N_2013,N_1782,N_1923);
nand U2014 (N_2014,N_1857,N_1792);
or U2015 (N_2015,N_1977,N_1801);
or U2016 (N_2016,N_1661,N_1520);
and U2017 (N_2017,N_1804,N_1699);
and U2018 (N_2018,N_1908,N_1829);
xnor U2019 (N_2019,N_1830,N_1824);
nor U2020 (N_2020,N_1677,N_1509);
or U2021 (N_2021,N_1669,N_1616);
and U2022 (N_2022,N_1649,N_1820);
nand U2023 (N_2023,N_1695,N_1807);
or U2024 (N_2024,N_1646,N_1783);
or U2025 (N_2025,N_1619,N_1858);
xnor U2026 (N_2026,N_1542,N_1945);
nor U2027 (N_2027,N_1859,N_1679);
and U2028 (N_2028,N_1890,N_1963);
xor U2029 (N_2029,N_1799,N_1573);
xor U2030 (N_2030,N_1655,N_1904);
or U2031 (N_2031,N_1902,N_1676);
nand U2032 (N_2032,N_1962,N_1626);
or U2033 (N_2033,N_1795,N_1605);
nand U2034 (N_2034,N_1511,N_1837);
and U2035 (N_2035,N_1627,N_1982);
nor U2036 (N_2036,N_1659,N_1674);
and U2037 (N_2037,N_1749,N_1884);
nor U2038 (N_2038,N_1867,N_1690);
or U2039 (N_2039,N_1821,N_1777);
or U2040 (N_2040,N_1721,N_1657);
xor U2041 (N_2041,N_1522,N_1852);
nor U2042 (N_2042,N_1535,N_1526);
or U2043 (N_2043,N_1814,N_1746);
nand U2044 (N_2044,N_1806,N_1958);
nand U2045 (N_2045,N_1630,N_1893);
nand U2046 (N_2046,N_1991,N_1747);
and U2047 (N_2047,N_1868,N_1827);
nand U2048 (N_2048,N_1938,N_1629);
nand U2049 (N_2049,N_1771,N_1726);
nor U2050 (N_2050,N_1773,N_1874);
or U2051 (N_2051,N_1697,N_1714);
or U2052 (N_2052,N_1975,N_1643);
nand U2053 (N_2053,N_1812,N_1598);
and U2054 (N_2054,N_1545,N_1905);
xnor U2055 (N_2055,N_1797,N_1850);
xor U2056 (N_2056,N_1767,N_1554);
and U2057 (N_2057,N_1609,N_1722);
or U2058 (N_2058,N_1769,N_1940);
and U2059 (N_2059,N_1912,N_1694);
nor U2060 (N_2060,N_1707,N_1591);
and U2061 (N_2061,N_1524,N_1998);
or U2062 (N_2062,N_1666,N_1577);
nand U2063 (N_2063,N_1851,N_1612);
nor U2064 (N_2064,N_1539,N_1741);
or U2065 (N_2065,N_1597,N_1907);
nor U2066 (N_2066,N_1798,N_1621);
nor U2067 (N_2067,N_1805,N_1922);
nor U2068 (N_2068,N_1543,N_1878);
nor U2069 (N_2069,N_1557,N_1832);
and U2070 (N_2070,N_1686,N_1835);
nor U2071 (N_2071,N_1899,N_1723);
or U2072 (N_2072,N_1574,N_1822);
and U2073 (N_2073,N_1620,N_1715);
and U2074 (N_2074,N_1813,N_1533);
and U2075 (N_2075,N_1882,N_1688);
nand U2076 (N_2076,N_1625,N_1706);
xor U2077 (N_2077,N_1633,N_1531);
and U2078 (N_2078,N_1810,N_1918);
and U2079 (N_2079,N_1941,N_1518);
nor U2080 (N_2080,N_1603,N_1624);
nand U2081 (N_2081,N_1634,N_1724);
xnor U2082 (N_2082,N_1709,N_1955);
or U2083 (N_2083,N_1892,N_1880);
or U2084 (N_2084,N_1565,N_1590);
nand U2085 (N_2085,N_1742,N_1503);
nand U2086 (N_2086,N_1917,N_1710);
or U2087 (N_2087,N_1550,N_1986);
nand U2088 (N_2088,N_1578,N_1834);
nand U2089 (N_2089,N_1928,N_1926);
nand U2090 (N_2090,N_1602,N_1754);
and U2091 (N_2091,N_1936,N_1973);
nand U2092 (N_2092,N_1725,N_1685);
and U2093 (N_2093,N_1934,N_1610);
nand U2094 (N_2094,N_1588,N_1700);
nor U2095 (N_2095,N_1637,N_1972);
nor U2096 (N_2096,N_1732,N_1984);
xnor U2097 (N_2097,N_1519,N_1903);
or U2098 (N_2098,N_1995,N_1601);
nand U2099 (N_2099,N_1582,N_1836);
nand U2100 (N_2100,N_1575,N_1964);
nor U2101 (N_2101,N_1877,N_1750);
nand U2102 (N_2102,N_1887,N_1713);
nand U2103 (N_2103,N_1818,N_1735);
nor U2104 (N_2104,N_1534,N_1794);
nor U2105 (N_2105,N_1895,N_1990);
xor U2106 (N_2106,N_1862,N_1615);
nand U2107 (N_2107,N_1757,N_1500);
xnor U2108 (N_2108,N_1931,N_1981);
nand U2109 (N_2109,N_1651,N_1593);
nand U2110 (N_2110,N_1863,N_1942);
or U2111 (N_2111,N_1983,N_1684);
nor U2112 (N_2112,N_1883,N_1528);
or U2113 (N_2113,N_1994,N_1585);
nand U2114 (N_2114,N_1993,N_1848);
nor U2115 (N_2115,N_1613,N_1910);
nand U2116 (N_2116,N_1513,N_1547);
nor U2117 (N_2117,N_1761,N_1996);
and U2118 (N_2118,N_1891,N_1816);
and U2119 (N_2119,N_1606,N_1898);
or U2120 (N_2120,N_1952,N_1825);
and U2121 (N_2121,N_1702,N_1617);
nand U2122 (N_2122,N_1787,N_1793);
and U2123 (N_2123,N_1507,N_1678);
nor U2124 (N_2124,N_1763,N_1841);
and U2125 (N_2125,N_1839,N_1970);
and U2126 (N_2126,N_1939,N_1774);
nor U2127 (N_2127,N_1758,N_1737);
or U2128 (N_2128,N_1762,N_1648);
and U2129 (N_2129,N_1776,N_1584);
nand U2130 (N_2130,N_1809,N_1592);
or U2131 (N_2131,N_1600,N_1933);
nor U2132 (N_2132,N_1564,N_1764);
nand U2133 (N_2133,N_1765,N_1759);
nand U2134 (N_2134,N_1521,N_1872);
nand U2135 (N_2135,N_1927,N_1949);
nor U2136 (N_2136,N_1683,N_1948);
nand U2137 (N_2137,N_1886,N_1583);
xnor U2138 (N_2138,N_1641,N_1711);
and U2139 (N_2139,N_1558,N_1897);
and U2140 (N_2140,N_1527,N_1504);
nor U2141 (N_2141,N_1561,N_1885);
xnor U2142 (N_2142,N_1819,N_1628);
nand U2143 (N_2143,N_1784,N_1576);
and U2144 (N_2144,N_1512,N_1935);
nor U2145 (N_2145,N_1652,N_1658);
nand U2146 (N_2146,N_1760,N_1718);
nor U2147 (N_2147,N_1719,N_1960);
or U2148 (N_2148,N_1790,N_1623);
or U2149 (N_2149,N_1921,N_1662);
nand U2150 (N_2150,N_1635,N_1570);
or U2151 (N_2151,N_1888,N_1731);
or U2152 (N_2152,N_1779,N_1571);
and U2153 (N_2153,N_1736,N_1866);
nand U2154 (N_2154,N_1889,N_1913);
nor U2155 (N_2155,N_1670,N_1650);
or U2156 (N_2156,N_1687,N_1559);
or U2157 (N_2157,N_1696,N_1607);
nor U2158 (N_2158,N_1525,N_1766);
or U2159 (N_2159,N_1640,N_1729);
or U2160 (N_2160,N_1508,N_1781);
and U2161 (N_2161,N_1869,N_1847);
or U2162 (N_2162,N_1673,N_1739);
or U2163 (N_2163,N_1967,N_1811);
or U2164 (N_2164,N_1900,N_1833);
nand U2165 (N_2165,N_1966,N_1738);
and U2166 (N_2166,N_1505,N_1842);
and U2167 (N_2167,N_1663,N_1555);
nand U2168 (N_2168,N_1567,N_1968);
xor U2169 (N_2169,N_1653,N_1712);
nand U2170 (N_2170,N_1800,N_1845);
nor U2171 (N_2171,N_1529,N_1698);
nand U2172 (N_2172,N_1544,N_1915);
and U2173 (N_2173,N_1755,N_1924);
or U2174 (N_2174,N_1789,N_1876);
and U2175 (N_2175,N_1667,N_1681);
nand U2176 (N_2176,N_1853,N_1595);
nor U2177 (N_2177,N_1815,N_1645);
nand U2178 (N_2178,N_1785,N_1560);
xor U2179 (N_2179,N_1596,N_1672);
xor U2180 (N_2180,N_1808,N_1548);
and U2181 (N_2181,N_1870,N_1997);
and U2182 (N_2182,N_1691,N_1817);
and U2183 (N_2183,N_1937,N_1775);
or U2184 (N_2184,N_1553,N_1728);
nor U2185 (N_2185,N_1614,N_1668);
xnor U2186 (N_2186,N_1906,N_1879);
and U2187 (N_2187,N_1638,N_1930);
nor U2188 (N_2188,N_1768,N_1979);
or U2189 (N_2189,N_1956,N_1957);
nor U2190 (N_2190,N_1756,N_1551);
nor U2191 (N_2191,N_1656,N_1778);
xor U2192 (N_2192,N_1969,N_1727);
or U2193 (N_2193,N_1523,N_1589);
nand U2194 (N_2194,N_1987,N_1631);
or U2195 (N_2195,N_1929,N_1701);
nand U2196 (N_2196,N_1716,N_1546);
nor U2197 (N_2197,N_1730,N_1569);
or U2198 (N_2198,N_1950,N_1786);
nor U2199 (N_2199,N_1506,N_1705);
nor U2200 (N_2200,N_1717,N_1618);
nor U2201 (N_2201,N_1682,N_1586);
or U2202 (N_2202,N_1654,N_1978);
nor U2203 (N_2203,N_1541,N_1611);
or U2204 (N_2204,N_1568,N_1587);
or U2205 (N_2205,N_1752,N_1894);
nor U2206 (N_2206,N_1748,N_1594);
nand U2207 (N_2207,N_1675,N_1849);
or U2208 (N_2208,N_1751,N_1875);
nor U2209 (N_2209,N_1860,N_1988);
xnor U2210 (N_2210,N_1703,N_1932);
nor U2211 (N_2211,N_1692,N_1772);
or U2212 (N_2212,N_1720,N_1992);
and U2213 (N_2213,N_1647,N_1733);
nand U2214 (N_2214,N_1861,N_1871);
and U2215 (N_2215,N_1562,N_1944);
nand U2216 (N_2216,N_1515,N_1581);
or U2217 (N_2217,N_1864,N_1501);
nor U2218 (N_2218,N_1514,N_1976);
xnor U2219 (N_2219,N_1919,N_1671);
or U2220 (N_2220,N_1745,N_1743);
nor U2221 (N_2221,N_1563,N_1622);
or U2222 (N_2222,N_1854,N_1516);
and U2223 (N_2223,N_1599,N_1971);
xnor U2224 (N_2224,N_1873,N_1770);
nor U2225 (N_2225,N_1536,N_1953);
nand U2226 (N_2226,N_1664,N_1961);
or U2227 (N_2227,N_1838,N_1901);
and U2228 (N_2228,N_1660,N_1510);
and U2229 (N_2229,N_1538,N_1828);
nor U2230 (N_2230,N_1947,N_1796);
or U2231 (N_2231,N_1704,N_1803);
nand U2232 (N_2232,N_1959,N_1999);
or U2233 (N_2233,N_1802,N_1989);
nand U2234 (N_2234,N_1608,N_1916);
or U2235 (N_2235,N_1909,N_1680);
and U2236 (N_2236,N_1788,N_1708);
nor U2237 (N_2237,N_1579,N_1734);
nand U2238 (N_2238,N_1517,N_1840);
nor U2239 (N_2239,N_1855,N_1911);
nor U2240 (N_2240,N_1644,N_1865);
and U2241 (N_2241,N_1844,N_1744);
or U2242 (N_2242,N_1946,N_1689);
or U2243 (N_2243,N_1740,N_1632);
and U2244 (N_2244,N_1826,N_1831);
nand U2245 (N_2245,N_1985,N_1954);
nand U2246 (N_2246,N_1925,N_1665);
nor U2247 (N_2247,N_1693,N_1604);
nand U2248 (N_2248,N_1980,N_1530);
and U2249 (N_2249,N_1914,N_1951);
nand U2250 (N_2250,N_1720,N_1727);
nand U2251 (N_2251,N_1958,N_1609);
nor U2252 (N_2252,N_1926,N_1643);
nand U2253 (N_2253,N_1790,N_1864);
or U2254 (N_2254,N_1807,N_1673);
nor U2255 (N_2255,N_1553,N_1958);
or U2256 (N_2256,N_1542,N_1905);
xor U2257 (N_2257,N_1735,N_1983);
nand U2258 (N_2258,N_1783,N_1859);
nor U2259 (N_2259,N_1710,N_1886);
xnor U2260 (N_2260,N_1792,N_1523);
or U2261 (N_2261,N_1868,N_1994);
and U2262 (N_2262,N_1591,N_1521);
xnor U2263 (N_2263,N_1507,N_1855);
nor U2264 (N_2264,N_1557,N_1575);
nand U2265 (N_2265,N_1607,N_1790);
or U2266 (N_2266,N_1558,N_1790);
and U2267 (N_2267,N_1793,N_1921);
nor U2268 (N_2268,N_1679,N_1503);
or U2269 (N_2269,N_1838,N_1622);
nor U2270 (N_2270,N_1862,N_1819);
xnor U2271 (N_2271,N_1972,N_1712);
nor U2272 (N_2272,N_1679,N_1841);
or U2273 (N_2273,N_1965,N_1718);
nand U2274 (N_2274,N_1915,N_1820);
and U2275 (N_2275,N_1621,N_1900);
or U2276 (N_2276,N_1946,N_1553);
or U2277 (N_2277,N_1800,N_1958);
or U2278 (N_2278,N_1587,N_1567);
nand U2279 (N_2279,N_1629,N_1883);
xor U2280 (N_2280,N_1898,N_1674);
and U2281 (N_2281,N_1774,N_1623);
or U2282 (N_2282,N_1662,N_1618);
nand U2283 (N_2283,N_1708,N_1916);
nor U2284 (N_2284,N_1895,N_1790);
nand U2285 (N_2285,N_1919,N_1638);
nand U2286 (N_2286,N_1779,N_1812);
nand U2287 (N_2287,N_1618,N_1899);
nor U2288 (N_2288,N_1872,N_1813);
nor U2289 (N_2289,N_1681,N_1977);
nand U2290 (N_2290,N_1901,N_1948);
nand U2291 (N_2291,N_1842,N_1995);
and U2292 (N_2292,N_1929,N_1580);
nand U2293 (N_2293,N_1871,N_1552);
and U2294 (N_2294,N_1987,N_1559);
and U2295 (N_2295,N_1940,N_1975);
and U2296 (N_2296,N_1736,N_1558);
and U2297 (N_2297,N_1823,N_1782);
nor U2298 (N_2298,N_1916,N_1891);
xnor U2299 (N_2299,N_1804,N_1595);
nor U2300 (N_2300,N_1708,N_1687);
nand U2301 (N_2301,N_1589,N_1549);
xor U2302 (N_2302,N_1963,N_1998);
or U2303 (N_2303,N_1587,N_1633);
or U2304 (N_2304,N_1995,N_1867);
or U2305 (N_2305,N_1781,N_1553);
and U2306 (N_2306,N_1934,N_1820);
and U2307 (N_2307,N_1536,N_1504);
nand U2308 (N_2308,N_1539,N_1732);
nor U2309 (N_2309,N_1966,N_1586);
xnor U2310 (N_2310,N_1613,N_1916);
xnor U2311 (N_2311,N_1811,N_1944);
xnor U2312 (N_2312,N_1858,N_1924);
nor U2313 (N_2313,N_1654,N_1761);
nor U2314 (N_2314,N_1990,N_1663);
nor U2315 (N_2315,N_1966,N_1508);
and U2316 (N_2316,N_1900,N_1772);
or U2317 (N_2317,N_1681,N_1843);
or U2318 (N_2318,N_1996,N_1642);
or U2319 (N_2319,N_1602,N_1980);
nand U2320 (N_2320,N_1790,N_1886);
and U2321 (N_2321,N_1874,N_1578);
xnor U2322 (N_2322,N_1933,N_1500);
and U2323 (N_2323,N_1768,N_1628);
or U2324 (N_2324,N_1821,N_1721);
xnor U2325 (N_2325,N_1543,N_1943);
and U2326 (N_2326,N_1591,N_1853);
xor U2327 (N_2327,N_1566,N_1685);
xor U2328 (N_2328,N_1519,N_1538);
and U2329 (N_2329,N_1774,N_1652);
or U2330 (N_2330,N_1874,N_1875);
nor U2331 (N_2331,N_1846,N_1855);
nor U2332 (N_2332,N_1939,N_1586);
nor U2333 (N_2333,N_1512,N_1666);
or U2334 (N_2334,N_1627,N_1890);
or U2335 (N_2335,N_1667,N_1901);
xor U2336 (N_2336,N_1664,N_1769);
and U2337 (N_2337,N_1827,N_1575);
nor U2338 (N_2338,N_1668,N_1503);
nor U2339 (N_2339,N_1722,N_1563);
nand U2340 (N_2340,N_1749,N_1665);
nand U2341 (N_2341,N_1820,N_1973);
or U2342 (N_2342,N_1772,N_1645);
and U2343 (N_2343,N_1872,N_1852);
and U2344 (N_2344,N_1997,N_1538);
nor U2345 (N_2345,N_1666,N_1678);
nor U2346 (N_2346,N_1974,N_1983);
and U2347 (N_2347,N_1776,N_1981);
nor U2348 (N_2348,N_1988,N_1759);
xor U2349 (N_2349,N_1889,N_1829);
and U2350 (N_2350,N_1689,N_1607);
nand U2351 (N_2351,N_1559,N_1845);
or U2352 (N_2352,N_1810,N_1577);
xor U2353 (N_2353,N_1982,N_1671);
or U2354 (N_2354,N_1739,N_1812);
nand U2355 (N_2355,N_1592,N_1926);
and U2356 (N_2356,N_1547,N_1681);
nand U2357 (N_2357,N_1678,N_1894);
nand U2358 (N_2358,N_1796,N_1747);
and U2359 (N_2359,N_1605,N_1821);
and U2360 (N_2360,N_1669,N_1673);
nor U2361 (N_2361,N_1974,N_1993);
or U2362 (N_2362,N_1564,N_1599);
nand U2363 (N_2363,N_1809,N_1693);
nor U2364 (N_2364,N_1677,N_1678);
or U2365 (N_2365,N_1862,N_1812);
nand U2366 (N_2366,N_1975,N_1987);
xnor U2367 (N_2367,N_1853,N_1964);
nor U2368 (N_2368,N_1851,N_1767);
nand U2369 (N_2369,N_1907,N_1767);
nor U2370 (N_2370,N_1895,N_1513);
and U2371 (N_2371,N_1616,N_1743);
nand U2372 (N_2372,N_1763,N_1869);
xor U2373 (N_2373,N_1980,N_1988);
or U2374 (N_2374,N_1706,N_1558);
xnor U2375 (N_2375,N_1956,N_1747);
and U2376 (N_2376,N_1843,N_1559);
xnor U2377 (N_2377,N_1907,N_1746);
and U2378 (N_2378,N_1947,N_1867);
nand U2379 (N_2379,N_1651,N_1663);
nor U2380 (N_2380,N_1711,N_1913);
or U2381 (N_2381,N_1820,N_1557);
nand U2382 (N_2382,N_1589,N_1672);
or U2383 (N_2383,N_1621,N_1819);
and U2384 (N_2384,N_1539,N_1833);
and U2385 (N_2385,N_1946,N_1683);
or U2386 (N_2386,N_1907,N_1846);
nand U2387 (N_2387,N_1933,N_1627);
nand U2388 (N_2388,N_1896,N_1558);
nor U2389 (N_2389,N_1845,N_1626);
nand U2390 (N_2390,N_1730,N_1531);
and U2391 (N_2391,N_1636,N_1560);
and U2392 (N_2392,N_1843,N_1703);
nand U2393 (N_2393,N_1711,N_1536);
nand U2394 (N_2394,N_1581,N_1692);
nor U2395 (N_2395,N_1759,N_1656);
nand U2396 (N_2396,N_1933,N_1966);
and U2397 (N_2397,N_1753,N_1755);
nor U2398 (N_2398,N_1842,N_1898);
nor U2399 (N_2399,N_1706,N_1844);
nand U2400 (N_2400,N_1535,N_1639);
nor U2401 (N_2401,N_1866,N_1919);
nand U2402 (N_2402,N_1657,N_1776);
or U2403 (N_2403,N_1983,N_1734);
nand U2404 (N_2404,N_1906,N_1593);
nor U2405 (N_2405,N_1952,N_1930);
and U2406 (N_2406,N_1660,N_1981);
and U2407 (N_2407,N_1833,N_1668);
nor U2408 (N_2408,N_1602,N_1917);
nand U2409 (N_2409,N_1555,N_1795);
xor U2410 (N_2410,N_1674,N_1569);
nor U2411 (N_2411,N_1846,N_1827);
or U2412 (N_2412,N_1587,N_1703);
xor U2413 (N_2413,N_1687,N_1563);
xnor U2414 (N_2414,N_1529,N_1748);
and U2415 (N_2415,N_1624,N_1609);
nor U2416 (N_2416,N_1708,N_1989);
nand U2417 (N_2417,N_1545,N_1815);
nand U2418 (N_2418,N_1946,N_1531);
nand U2419 (N_2419,N_1657,N_1529);
nor U2420 (N_2420,N_1634,N_1846);
and U2421 (N_2421,N_1844,N_1688);
xor U2422 (N_2422,N_1868,N_1746);
and U2423 (N_2423,N_1758,N_1658);
or U2424 (N_2424,N_1686,N_1982);
nor U2425 (N_2425,N_1812,N_1654);
nand U2426 (N_2426,N_1548,N_1841);
or U2427 (N_2427,N_1714,N_1923);
nand U2428 (N_2428,N_1781,N_1773);
or U2429 (N_2429,N_1681,N_1776);
xnor U2430 (N_2430,N_1772,N_1998);
or U2431 (N_2431,N_1726,N_1515);
nor U2432 (N_2432,N_1811,N_1787);
nand U2433 (N_2433,N_1788,N_1519);
nor U2434 (N_2434,N_1998,N_1529);
nor U2435 (N_2435,N_1530,N_1965);
and U2436 (N_2436,N_1849,N_1976);
or U2437 (N_2437,N_1805,N_1638);
nor U2438 (N_2438,N_1909,N_1698);
xor U2439 (N_2439,N_1959,N_1560);
or U2440 (N_2440,N_1865,N_1688);
and U2441 (N_2441,N_1995,N_1721);
or U2442 (N_2442,N_1985,N_1731);
nor U2443 (N_2443,N_1969,N_1630);
or U2444 (N_2444,N_1977,N_1633);
xor U2445 (N_2445,N_1637,N_1727);
and U2446 (N_2446,N_1718,N_1570);
and U2447 (N_2447,N_1799,N_1825);
nor U2448 (N_2448,N_1696,N_1706);
xor U2449 (N_2449,N_1557,N_1924);
nor U2450 (N_2450,N_1545,N_1702);
nand U2451 (N_2451,N_1500,N_1611);
nor U2452 (N_2452,N_1539,N_1909);
and U2453 (N_2453,N_1847,N_1597);
and U2454 (N_2454,N_1679,N_1938);
or U2455 (N_2455,N_1635,N_1892);
and U2456 (N_2456,N_1644,N_1511);
and U2457 (N_2457,N_1697,N_1509);
nor U2458 (N_2458,N_1704,N_1534);
nor U2459 (N_2459,N_1508,N_1851);
nor U2460 (N_2460,N_1552,N_1589);
or U2461 (N_2461,N_1992,N_1737);
nor U2462 (N_2462,N_1616,N_1998);
nand U2463 (N_2463,N_1716,N_1533);
and U2464 (N_2464,N_1819,N_1641);
and U2465 (N_2465,N_1929,N_1665);
and U2466 (N_2466,N_1603,N_1551);
nand U2467 (N_2467,N_1859,N_1643);
nor U2468 (N_2468,N_1815,N_1832);
or U2469 (N_2469,N_1871,N_1761);
and U2470 (N_2470,N_1830,N_1630);
nand U2471 (N_2471,N_1834,N_1869);
nor U2472 (N_2472,N_1986,N_1744);
nand U2473 (N_2473,N_1938,N_1545);
xnor U2474 (N_2474,N_1800,N_1586);
and U2475 (N_2475,N_1811,N_1734);
or U2476 (N_2476,N_1656,N_1703);
and U2477 (N_2477,N_1796,N_1607);
nor U2478 (N_2478,N_1882,N_1699);
nand U2479 (N_2479,N_1541,N_1886);
nand U2480 (N_2480,N_1659,N_1731);
nor U2481 (N_2481,N_1922,N_1958);
or U2482 (N_2482,N_1949,N_1783);
nand U2483 (N_2483,N_1934,N_1582);
or U2484 (N_2484,N_1868,N_1869);
or U2485 (N_2485,N_1758,N_1915);
nor U2486 (N_2486,N_1664,N_1726);
nand U2487 (N_2487,N_1849,N_1955);
and U2488 (N_2488,N_1795,N_1763);
nor U2489 (N_2489,N_1903,N_1542);
nand U2490 (N_2490,N_1904,N_1525);
nand U2491 (N_2491,N_1538,N_1816);
nand U2492 (N_2492,N_1581,N_1827);
xnor U2493 (N_2493,N_1869,N_1523);
or U2494 (N_2494,N_1865,N_1630);
and U2495 (N_2495,N_1503,N_1874);
nor U2496 (N_2496,N_1604,N_1698);
nand U2497 (N_2497,N_1878,N_1599);
nor U2498 (N_2498,N_1892,N_1945);
or U2499 (N_2499,N_1636,N_1890);
or U2500 (N_2500,N_2059,N_2246);
and U2501 (N_2501,N_2227,N_2192);
nand U2502 (N_2502,N_2431,N_2354);
nor U2503 (N_2503,N_2197,N_2018);
or U2504 (N_2504,N_2161,N_2170);
nor U2505 (N_2505,N_2331,N_2232);
nand U2506 (N_2506,N_2350,N_2153);
and U2507 (N_2507,N_2374,N_2324);
nor U2508 (N_2508,N_2009,N_2330);
or U2509 (N_2509,N_2029,N_2322);
and U2510 (N_2510,N_2352,N_2455);
xor U2511 (N_2511,N_2258,N_2397);
xnor U2512 (N_2512,N_2128,N_2454);
nand U2513 (N_2513,N_2200,N_2235);
or U2514 (N_2514,N_2301,N_2447);
xor U2515 (N_2515,N_2003,N_2090);
nor U2516 (N_2516,N_2412,N_2440);
nand U2517 (N_2517,N_2098,N_2494);
nor U2518 (N_2518,N_2483,N_2473);
nand U2519 (N_2519,N_2384,N_2433);
or U2520 (N_2520,N_2470,N_2326);
nor U2521 (N_2521,N_2104,N_2225);
or U2522 (N_2522,N_2303,N_2135);
and U2523 (N_2523,N_2188,N_2120);
nand U2524 (N_2524,N_2244,N_2492);
nor U2525 (N_2525,N_2425,N_2351);
and U2526 (N_2526,N_2398,N_2248);
and U2527 (N_2527,N_2268,N_2233);
or U2528 (N_2528,N_2243,N_2103);
nor U2529 (N_2529,N_2189,N_2062);
and U2530 (N_2530,N_2367,N_2224);
or U2531 (N_2531,N_2392,N_2485);
nor U2532 (N_2532,N_2482,N_2162);
nand U2533 (N_2533,N_2343,N_2280);
and U2534 (N_2534,N_2495,N_2156);
or U2535 (N_2535,N_2220,N_2068);
and U2536 (N_2536,N_2286,N_2019);
and U2537 (N_2537,N_2006,N_2209);
and U2538 (N_2538,N_2031,N_2279);
or U2539 (N_2539,N_2176,N_2166);
xnor U2540 (N_2540,N_2057,N_2381);
and U2541 (N_2541,N_2345,N_2370);
nor U2542 (N_2542,N_2278,N_2269);
xnor U2543 (N_2543,N_2105,N_2484);
or U2544 (N_2544,N_2493,N_2038);
or U2545 (N_2545,N_2358,N_2346);
nor U2546 (N_2546,N_2382,N_2335);
xor U2547 (N_2547,N_2052,N_2085);
nand U2548 (N_2548,N_2420,N_2064);
nor U2549 (N_2549,N_2298,N_2297);
nand U2550 (N_2550,N_2388,N_2403);
xor U2551 (N_2551,N_2314,N_2216);
nor U2552 (N_2552,N_2313,N_2304);
or U2553 (N_2553,N_2069,N_2179);
nand U2554 (N_2554,N_2137,N_2284);
or U2555 (N_2555,N_2142,N_2087);
xnor U2556 (N_2556,N_2110,N_2404);
or U2557 (N_2557,N_2445,N_2318);
nand U2558 (N_2558,N_2044,N_2228);
and U2559 (N_2559,N_2212,N_2402);
or U2560 (N_2560,N_2187,N_2174);
nand U2561 (N_2561,N_2373,N_2355);
nand U2562 (N_2562,N_2150,N_2293);
nor U2563 (N_2563,N_2287,N_2289);
or U2564 (N_2564,N_2469,N_2210);
xor U2565 (N_2565,N_2146,N_2480);
or U2566 (N_2566,N_2184,N_2121);
nor U2567 (N_2567,N_2256,N_2117);
xor U2568 (N_2568,N_2111,N_2000);
and U2569 (N_2569,N_2362,N_2109);
xnor U2570 (N_2570,N_2453,N_2035);
and U2571 (N_2571,N_2181,N_2101);
nor U2572 (N_2572,N_2321,N_2472);
nor U2573 (N_2573,N_2229,N_2474);
nor U2574 (N_2574,N_2406,N_2338);
xor U2575 (N_2575,N_2028,N_2134);
or U2576 (N_2576,N_2027,N_2122);
xor U2577 (N_2577,N_2058,N_2329);
nor U2578 (N_2578,N_2283,N_2262);
or U2579 (N_2579,N_2276,N_2475);
and U2580 (N_2580,N_2114,N_2395);
nand U2581 (N_2581,N_2159,N_2095);
nor U2582 (N_2582,N_2088,N_2400);
or U2583 (N_2583,N_2257,N_2372);
nand U2584 (N_2584,N_2306,N_2093);
or U2585 (N_2585,N_2154,N_2172);
nand U2586 (N_2586,N_2488,N_2070);
or U2587 (N_2587,N_2079,N_2049);
or U2588 (N_2588,N_2190,N_2061);
nand U2589 (N_2589,N_2496,N_2045);
nand U2590 (N_2590,N_2436,N_2323);
nand U2591 (N_2591,N_2168,N_2039);
nor U2592 (N_2592,N_2389,N_2130);
nor U2593 (N_2593,N_2077,N_2055);
and U2594 (N_2594,N_2364,N_2042);
xor U2595 (N_2595,N_2083,N_2173);
and U2596 (N_2596,N_2040,N_2332);
or U2597 (N_2597,N_2291,N_2020);
nor U2598 (N_2598,N_2127,N_2378);
or U2599 (N_2599,N_2429,N_2094);
or U2600 (N_2600,N_2336,N_2479);
or U2601 (N_2601,N_2295,N_2437);
and U2602 (N_2602,N_2145,N_2241);
nor U2603 (N_2603,N_2033,N_2065);
nor U2604 (N_2604,N_2334,N_2466);
or U2605 (N_2605,N_2219,N_2308);
nor U2606 (N_2606,N_2066,N_2076);
or U2607 (N_2607,N_2271,N_2203);
nand U2608 (N_2608,N_2277,N_2072);
nor U2609 (N_2609,N_2468,N_2490);
nor U2610 (N_2610,N_2337,N_2463);
nor U2611 (N_2611,N_2113,N_2457);
nand U2612 (N_2612,N_2010,N_2043);
or U2613 (N_2613,N_2254,N_2247);
xor U2614 (N_2614,N_2417,N_2396);
nor U2615 (N_2615,N_2091,N_2405);
or U2616 (N_2616,N_2196,N_2311);
or U2617 (N_2617,N_2408,N_2185);
or U2618 (N_2618,N_2261,N_2422);
nand U2619 (N_2619,N_2459,N_2143);
nor U2620 (N_2620,N_2363,N_2218);
or U2621 (N_2621,N_2414,N_2129);
xnor U2622 (N_2622,N_2021,N_2008);
and U2623 (N_2623,N_2164,N_2296);
and U2624 (N_2624,N_2084,N_2266);
nor U2625 (N_2625,N_2089,N_2202);
and U2626 (N_2626,N_2393,N_2419);
nor U2627 (N_2627,N_2237,N_2163);
nand U2628 (N_2628,N_2407,N_2239);
nor U2629 (N_2629,N_2133,N_2319);
or U2630 (N_2630,N_2001,N_2016);
and U2631 (N_2631,N_2305,N_2242);
or U2632 (N_2632,N_2444,N_2071);
or U2633 (N_2633,N_2399,N_2086);
nor U2634 (N_2634,N_2063,N_2100);
or U2635 (N_2635,N_2245,N_2307);
nor U2636 (N_2636,N_2251,N_2149);
nand U2637 (N_2637,N_2231,N_2158);
nor U2638 (N_2638,N_2365,N_2169);
nor U2639 (N_2639,N_2198,N_2073);
and U2640 (N_2640,N_2223,N_2178);
nand U2641 (N_2641,N_2157,N_2285);
and U2642 (N_2642,N_2361,N_2380);
and U2643 (N_2643,N_2348,N_2141);
nor U2644 (N_2644,N_2394,N_2339);
nand U2645 (N_2645,N_2281,N_2467);
or U2646 (N_2646,N_2344,N_2012);
nor U2647 (N_2647,N_2208,N_2102);
or U2648 (N_2648,N_2160,N_2327);
nor U2649 (N_2649,N_2386,N_2259);
and U2650 (N_2650,N_2477,N_2487);
and U2651 (N_2651,N_2265,N_2030);
nand U2652 (N_2652,N_2053,N_2119);
or U2653 (N_2653,N_2385,N_2152);
or U2654 (N_2654,N_2215,N_2371);
and U2655 (N_2655,N_2004,N_2222);
and U2656 (N_2656,N_2423,N_2186);
nor U2657 (N_2657,N_2250,N_2451);
nor U2658 (N_2658,N_2275,N_2140);
and U2659 (N_2659,N_2424,N_2213);
nand U2660 (N_2660,N_2108,N_2106);
or U2661 (N_2661,N_2011,N_2302);
and U2662 (N_2662,N_2067,N_2464);
nand U2663 (N_2663,N_2236,N_2443);
nand U2664 (N_2664,N_2340,N_2204);
nand U2665 (N_2665,N_2206,N_2341);
nor U2666 (N_2666,N_2461,N_2115);
and U2667 (N_2667,N_2409,N_2015);
and U2668 (N_2668,N_2449,N_2132);
nor U2669 (N_2669,N_2497,N_2240);
nand U2670 (N_2670,N_2353,N_2118);
or U2671 (N_2671,N_2014,N_2290);
and U2672 (N_2672,N_2252,N_2050);
nor U2673 (N_2673,N_2448,N_2144);
xnor U2674 (N_2674,N_2441,N_2498);
or U2675 (N_2675,N_2125,N_2180);
or U2676 (N_2676,N_2342,N_2476);
and U2677 (N_2677,N_2465,N_2249);
and U2678 (N_2678,N_2013,N_2138);
nand U2679 (N_2679,N_2201,N_2272);
and U2680 (N_2680,N_2390,N_2489);
or U2681 (N_2681,N_2312,N_2096);
or U2682 (N_2682,N_2136,N_2270);
and U2683 (N_2683,N_2041,N_2195);
nand U2684 (N_2684,N_2401,N_2460);
nand U2685 (N_2685,N_2375,N_2191);
and U2686 (N_2686,N_2415,N_2491);
or U2687 (N_2687,N_2263,N_2238);
and U2688 (N_2688,N_2325,N_2060);
nor U2689 (N_2689,N_2025,N_2116);
nand U2690 (N_2690,N_2317,N_2081);
nor U2691 (N_2691,N_2048,N_2282);
nor U2692 (N_2692,N_2205,N_2387);
and U2693 (N_2693,N_2383,N_2047);
nor U2694 (N_2694,N_2368,N_2421);
or U2695 (N_2695,N_2328,N_2267);
nor U2696 (N_2696,N_2234,N_2446);
or U2697 (N_2697,N_2131,N_2037);
nand U2698 (N_2698,N_2315,N_2023);
or U2699 (N_2699,N_2349,N_2471);
nor U2700 (N_2700,N_2428,N_2036);
and U2701 (N_2701,N_2430,N_2413);
nand U2702 (N_2702,N_2357,N_2226);
or U2703 (N_2703,N_2299,N_2026);
xor U2704 (N_2704,N_2426,N_2456);
and U2705 (N_2705,N_2310,N_2002);
nand U2706 (N_2706,N_2051,N_2123);
nor U2707 (N_2707,N_2264,N_2171);
nand U2708 (N_2708,N_2221,N_2435);
and U2709 (N_2709,N_2481,N_2366);
or U2710 (N_2710,N_2175,N_2418);
and U2711 (N_2711,N_2182,N_2356);
or U2712 (N_2712,N_2292,N_2126);
xor U2713 (N_2713,N_2450,N_2075);
nand U2714 (N_2714,N_2253,N_2124);
and U2715 (N_2715,N_2177,N_2092);
or U2716 (N_2716,N_2112,N_2165);
or U2717 (N_2717,N_2432,N_2217);
xor U2718 (N_2718,N_2074,N_2017);
nor U2719 (N_2719,N_2139,N_2147);
nand U2720 (N_2720,N_2439,N_2434);
or U2721 (N_2721,N_2300,N_2024);
nor U2722 (N_2722,N_2347,N_2097);
xnor U2723 (N_2723,N_2452,N_2214);
nor U2724 (N_2724,N_2230,N_2056);
nor U2725 (N_2725,N_2391,N_2320);
nand U2726 (N_2726,N_2260,N_2078);
and U2727 (N_2727,N_2309,N_2005);
or U2728 (N_2728,N_2034,N_2273);
or U2729 (N_2729,N_2499,N_2359);
xor U2730 (N_2730,N_2411,N_2458);
nand U2731 (N_2731,N_2462,N_2288);
and U2732 (N_2732,N_2082,N_2046);
xnor U2733 (N_2733,N_2360,N_2294);
and U2734 (N_2734,N_2316,N_2199);
and U2735 (N_2735,N_2032,N_2080);
nand U2736 (N_2736,N_2107,N_2442);
nor U2737 (N_2737,N_2194,N_2410);
nor U2738 (N_2738,N_2151,N_2099);
or U2739 (N_2739,N_2274,N_2379);
or U2740 (N_2740,N_2155,N_2054);
or U2741 (N_2741,N_2416,N_2207);
xnor U2742 (N_2742,N_2148,N_2376);
and U2743 (N_2743,N_2333,N_2438);
and U2744 (N_2744,N_2255,N_2007);
or U2745 (N_2745,N_2369,N_2211);
nand U2746 (N_2746,N_2427,N_2193);
xnor U2747 (N_2747,N_2478,N_2183);
nor U2748 (N_2748,N_2167,N_2022);
or U2749 (N_2749,N_2486,N_2377);
nor U2750 (N_2750,N_2296,N_2047);
xor U2751 (N_2751,N_2239,N_2178);
xor U2752 (N_2752,N_2423,N_2328);
or U2753 (N_2753,N_2296,N_2382);
nor U2754 (N_2754,N_2230,N_2028);
and U2755 (N_2755,N_2112,N_2183);
nand U2756 (N_2756,N_2423,N_2266);
or U2757 (N_2757,N_2477,N_2289);
nand U2758 (N_2758,N_2024,N_2312);
nor U2759 (N_2759,N_2375,N_2460);
or U2760 (N_2760,N_2262,N_2000);
xor U2761 (N_2761,N_2303,N_2010);
nor U2762 (N_2762,N_2182,N_2019);
nor U2763 (N_2763,N_2388,N_2146);
nor U2764 (N_2764,N_2455,N_2133);
and U2765 (N_2765,N_2026,N_2335);
or U2766 (N_2766,N_2331,N_2266);
and U2767 (N_2767,N_2372,N_2103);
nor U2768 (N_2768,N_2172,N_2415);
or U2769 (N_2769,N_2071,N_2082);
and U2770 (N_2770,N_2233,N_2221);
xor U2771 (N_2771,N_2131,N_2056);
and U2772 (N_2772,N_2038,N_2279);
or U2773 (N_2773,N_2211,N_2068);
nor U2774 (N_2774,N_2386,N_2392);
or U2775 (N_2775,N_2165,N_2087);
and U2776 (N_2776,N_2266,N_2132);
nand U2777 (N_2777,N_2237,N_2232);
and U2778 (N_2778,N_2007,N_2285);
nor U2779 (N_2779,N_2428,N_2204);
nor U2780 (N_2780,N_2403,N_2278);
xnor U2781 (N_2781,N_2380,N_2145);
nor U2782 (N_2782,N_2482,N_2414);
nand U2783 (N_2783,N_2400,N_2170);
and U2784 (N_2784,N_2137,N_2109);
nand U2785 (N_2785,N_2051,N_2140);
and U2786 (N_2786,N_2120,N_2155);
and U2787 (N_2787,N_2096,N_2392);
and U2788 (N_2788,N_2488,N_2244);
or U2789 (N_2789,N_2201,N_2424);
and U2790 (N_2790,N_2025,N_2166);
xor U2791 (N_2791,N_2367,N_2127);
nor U2792 (N_2792,N_2369,N_2067);
nand U2793 (N_2793,N_2293,N_2367);
xnor U2794 (N_2794,N_2448,N_2094);
nor U2795 (N_2795,N_2286,N_2128);
and U2796 (N_2796,N_2448,N_2118);
nand U2797 (N_2797,N_2011,N_2377);
and U2798 (N_2798,N_2191,N_2130);
or U2799 (N_2799,N_2377,N_2319);
or U2800 (N_2800,N_2394,N_2261);
nor U2801 (N_2801,N_2430,N_2158);
or U2802 (N_2802,N_2016,N_2008);
or U2803 (N_2803,N_2193,N_2167);
nand U2804 (N_2804,N_2414,N_2033);
nor U2805 (N_2805,N_2364,N_2175);
nor U2806 (N_2806,N_2133,N_2140);
or U2807 (N_2807,N_2375,N_2096);
nor U2808 (N_2808,N_2306,N_2239);
and U2809 (N_2809,N_2076,N_2134);
xnor U2810 (N_2810,N_2466,N_2041);
and U2811 (N_2811,N_2230,N_2429);
and U2812 (N_2812,N_2189,N_2363);
nand U2813 (N_2813,N_2363,N_2051);
or U2814 (N_2814,N_2167,N_2084);
and U2815 (N_2815,N_2192,N_2270);
xor U2816 (N_2816,N_2434,N_2345);
nand U2817 (N_2817,N_2024,N_2081);
nor U2818 (N_2818,N_2398,N_2354);
nand U2819 (N_2819,N_2281,N_2485);
and U2820 (N_2820,N_2465,N_2392);
and U2821 (N_2821,N_2388,N_2179);
or U2822 (N_2822,N_2402,N_2496);
nor U2823 (N_2823,N_2004,N_2276);
nand U2824 (N_2824,N_2499,N_2311);
nor U2825 (N_2825,N_2171,N_2295);
nor U2826 (N_2826,N_2408,N_2423);
or U2827 (N_2827,N_2248,N_2490);
and U2828 (N_2828,N_2176,N_2045);
nor U2829 (N_2829,N_2321,N_2435);
or U2830 (N_2830,N_2444,N_2369);
nand U2831 (N_2831,N_2013,N_2385);
and U2832 (N_2832,N_2151,N_2000);
or U2833 (N_2833,N_2426,N_2408);
and U2834 (N_2834,N_2394,N_2439);
and U2835 (N_2835,N_2045,N_2011);
nand U2836 (N_2836,N_2115,N_2187);
nor U2837 (N_2837,N_2225,N_2061);
or U2838 (N_2838,N_2400,N_2057);
nand U2839 (N_2839,N_2245,N_2383);
nand U2840 (N_2840,N_2234,N_2206);
or U2841 (N_2841,N_2356,N_2412);
and U2842 (N_2842,N_2047,N_2410);
nor U2843 (N_2843,N_2477,N_2209);
nor U2844 (N_2844,N_2443,N_2472);
nor U2845 (N_2845,N_2190,N_2046);
nor U2846 (N_2846,N_2024,N_2281);
xor U2847 (N_2847,N_2008,N_2027);
nor U2848 (N_2848,N_2120,N_2174);
nand U2849 (N_2849,N_2117,N_2179);
xnor U2850 (N_2850,N_2160,N_2111);
nand U2851 (N_2851,N_2123,N_2200);
nand U2852 (N_2852,N_2455,N_2108);
nor U2853 (N_2853,N_2298,N_2245);
xnor U2854 (N_2854,N_2135,N_2251);
nor U2855 (N_2855,N_2280,N_2379);
nand U2856 (N_2856,N_2425,N_2347);
xor U2857 (N_2857,N_2276,N_2265);
nor U2858 (N_2858,N_2174,N_2342);
nor U2859 (N_2859,N_2265,N_2043);
nor U2860 (N_2860,N_2468,N_2287);
nor U2861 (N_2861,N_2193,N_2397);
nand U2862 (N_2862,N_2422,N_2166);
nand U2863 (N_2863,N_2412,N_2014);
and U2864 (N_2864,N_2203,N_2223);
nor U2865 (N_2865,N_2125,N_2020);
nor U2866 (N_2866,N_2217,N_2327);
and U2867 (N_2867,N_2492,N_2414);
nand U2868 (N_2868,N_2466,N_2386);
and U2869 (N_2869,N_2356,N_2167);
or U2870 (N_2870,N_2027,N_2330);
or U2871 (N_2871,N_2034,N_2472);
and U2872 (N_2872,N_2132,N_2408);
nor U2873 (N_2873,N_2461,N_2205);
and U2874 (N_2874,N_2234,N_2259);
and U2875 (N_2875,N_2288,N_2365);
nor U2876 (N_2876,N_2199,N_2393);
xnor U2877 (N_2877,N_2316,N_2070);
nor U2878 (N_2878,N_2213,N_2468);
nor U2879 (N_2879,N_2444,N_2242);
xor U2880 (N_2880,N_2015,N_2062);
nand U2881 (N_2881,N_2268,N_2029);
and U2882 (N_2882,N_2190,N_2460);
and U2883 (N_2883,N_2026,N_2112);
xnor U2884 (N_2884,N_2018,N_2156);
nor U2885 (N_2885,N_2390,N_2329);
nand U2886 (N_2886,N_2087,N_2057);
and U2887 (N_2887,N_2187,N_2227);
nand U2888 (N_2888,N_2066,N_2115);
and U2889 (N_2889,N_2182,N_2136);
or U2890 (N_2890,N_2049,N_2132);
and U2891 (N_2891,N_2438,N_2168);
or U2892 (N_2892,N_2171,N_2192);
nand U2893 (N_2893,N_2290,N_2383);
and U2894 (N_2894,N_2338,N_2070);
xnor U2895 (N_2895,N_2144,N_2057);
and U2896 (N_2896,N_2140,N_2458);
nor U2897 (N_2897,N_2411,N_2322);
or U2898 (N_2898,N_2483,N_2001);
or U2899 (N_2899,N_2371,N_2160);
nand U2900 (N_2900,N_2057,N_2330);
nand U2901 (N_2901,N_2258,N_2398);
nor U2902 (N_2902,N_2253,N_2422);
nor U2903 (N_2903,N_2256,N_2175);
nand U2904 (N_2904,N_2319,N_2320);
and U2905 (N_2905,N_2476,N_2330);
xnor U2906 (N_2906,N_2289,N_2141);
and U2907 (N_2907,N_2368,N_2463);
nand U2908 (N_2908,N_2266,N_2097);
nand U2909 (N_2909,N_2064,N_2303);
and U2910 (N_2910,N_2052,N_2469);
xnor U2911 (N_2911,N_2264,N_2047);
nor U2912 (N_2912,N_2473,N_2016);
nand U2913 (N_2913,N_2159,N_2384);
or U2914 (N_2914,N_2486,N_2271);
nand U2915 (N_2915,N_2308,N_2064);
and U2916 (N_2916,N_2037,N_2141);
and U2917 (N_2917,N_2153,N_2398);
and U2918 (N_2918,N_2031,N_2366);
and U2919 (N_2919,N_2409,N_2075);
nand U2920 (N_2920,N_2368,N_2018);
or U2921 (N_2921,N_2487,N_2202);
nor U2922 (N_2922,N_2314,N_2484);
or U2923 (N_2923,N_2021,N_2028);
nor U2924 (N_2924,N_2059,N_2216);
and U2925 (N_2925,N_2340,N_2194);
and U2926 (N_2926,N_2124,N_2447);
or U2927 (N_2927,N_2231,N_2157);
nor U2928 (N_2928,N_2098,N_2069);
nand U2929 (N_2929,N_2215,N_2180);
or U2930 (N_2930,N_2233,N_2001);
nor U2931 (N_2931,N_2050,N_2299);
and U2932 (N_2932,N_2492,N_2487);
nor U2933 (N_2933,N_2034,N_2399);
nand U2934 (N_2934,N_2290,N_2120);
nor U2935 (N_2935,N_2116,N_2260);
nor U2936 (N_2936,N_2281,N_2437);
nor U2937 (N_2937,N_2265,N_2407);
xnor U2938 (N_2938,N_2384,N_2414);
xnor U2939 (N_2939,N_2245,N_2279);
nand U2940 (N_2940,N_2416,N_2442);
or U2941 (N_2941,N_2071,N_2164);
and U2942 (N_2942,N_2292,N_2127);
or U2943 (N_2943,N_2287,N_2016);
nor U2944 (N_2944,N_2137,N_2071);
nand U2945 (N_2945,N_2459,N_2173);
nand U2946 (N_2946,N_2051,N_2263);
xnor U2947 (N_2947,N_2097,N_2211);
nand U2948 (N_2948,N_2281,N_2225);
or U2949 (N_2949,N_2447,N_2097);
xnor U2950 (N_2950,N_2059,N_2324);
or U2951 (N_2951,N_2197,N_2010);
nand U2952 (N_2952,N_2254,N_2427);
and U2953 (N_2953,N_2341,N_2059);
nor U2954 (N_2954,N_2210,N_2348);
nand U2955 (N_2955,N_2029,N_2488);
or U2956 (N_2956,N_2413,N_2005);
or U2957 (N_2957,N_2023,N_2335);
nor U2958 (N_2958,N_2182,N_2381);
and U2959 (N_2959,N_2203,N_2013);
or U2960 (N_2960,N_2253,N_2304);
or U2961 (N_2961,N_2104,N_2376);
or U2962 (N_2962,N_2222,N_2143);
nor U2963 (N_2963,N_2154,N_2443);
xor U2964 (N_2964,N_2376,N_2459);
nand U2965 (N_2965,N_2212,N_2187);
and U2966 (N_2966,N_2045,N_2476);
and U2967 (N_2967,N_2089,N_2018);
nor U2968 (N_2968,N_2012,N_2400);
or U2969 (N_2969,N_2032,N_2264);
and U2970 (N_2970,N_2390,N_2352);
nor U2971 (N_2971,N_2184,N_2222);
and U2972 (N_2972,N_2214,N_2011);
nor U2973 (N_2973,N_2009,N_2015);
nand U2974 (N_2974,N_2347,N_2416);
or U2975 (N_2975,N_2457,N_2011);
and U2976 (N_2976,N_2009,N_2300);
xnor U2977 (N_2977,N_2240,N_2073);
or U2978 (N_2978,N_2192,N_2220);
or U2979 (N_2979,N_2350,N_2173);
and U2980 (N_2980,N_2382,N_2022);
xnor U2981 (N_2981,N_2395,N_2328);
xnor U2982 (N_2982,N_2108,N_2323);
nor U2983 (N_2983,N_2456,N_2292);
or U2984 (N_2984,N_2078,N_2211);
nor U2985 (N_2985,N_2339,N_2235);
or U2986 (N_2986,N_2154,N_2251);
and U2987 (N_2987,N_2173,N_2043);
and U2988 (N_2988,N_2381,N_2442);
and U2989 (N_2989,N_2115,N_2376);
nor U2990 (N_2990,N_2125,N_2450);
or U2991 (N_2991,N_2131,N_2409);
or U2992 (N_2992,N_2496,N_2385);
or U2993 (N_2993,N_2383,N_2077);
nor U2994 (N_2994,N_2466,N_2430);
and U2995 (N_2995,N_2334,N_2265);
nor U2996 (N_2996,N_2497,N_2322);
and U2997 (N_2997,N_2134,N_2407);
nor U2998 (N_2998,N_2037,N_2221);
nor U2999 (N_2999,N_2471,N_2096);
nor U3000 (N_3000,N_2979,N_2548);
and U3001 (N_3001,N_2938,N_2503);
or U3002 (N_3002,N_2819,N_2595);
or U3003 (N_3003,N_2937,N_2678);
nand U3004 (N_3004,N_2813,N_2874);
xnor U3005 (N_3005,N_2531,N_2856);
xor U3006 (N_3006,N_2952,N_2796);
or U3007 (N_3007,N_2839,N_2618);
nand U3008 (N_3008,N_2835,N_2666);
or U3009 (N_3009,N_2764,N_2768);
nand U3010 (N_3010,N_2515,N_2765);
xor U3011 (N_3011,N_2568,N_2545);
nand U3012 (N_3012,N_2975,N_2941);
nor U3013 (N_3013,N_2645,N_2945);
and U3014 (N_3014,N_2907,N_2668);
xor U3015 (N_3015,N_2906,N_2875);
nor U3016 (N_3016,N_2701,N_2532);
nor U3017 (N_3017,N_2556,N_2752);
and U3018 (N_3018,N_2886,N_2629);
nand U3019 (N_3019,N_2639,N_2505);
xnor U3020 (N_3020,N_2627,N_2546);
nand U3021 (N_3021,N_2584,N_2617);
or U3022 (N_3022,N_2721,N_2892);
or U3023 (N_3023,N_2884,N_2836);
nor U3024 (N_3024,N_2911,N_2877);
nand U3025 (N_3025,N_2602,N_2872);
or U3026 (N_3026,N_2832,N_2606);
nor U3027 (N_3027,N_2654,N_2644);
and U3028 (N_3028,N_2727,N_2715);
xnor U3029 (N_3029,N_2923,N_2983);
nand U3030 (N_3030,N_2706,N_2871);
and U3031 (N_3031,N_2587,N_2795);
nand U3032 (N_3032,N_2554,N_2736);
nand U3033 (N_3033,N_2916,N_2868);
or U3034 (N_3034,N_2821,N_2571);
or U3035 (N_3035,N_2843,N_2558);
or U3036 (N_3036,N_2905,N_2737);
nand U3037 (N_3037,N_2812,N_2805);
nand U3038 (N_3038,N_2598,N_2722);
nand U3039 (N_3039,N_2744,N_2588);
nor U3040 (N_3040,N_2502,N_2538);
or U3041 (N_3041,N_2763,N_2616);
nor U3042 (N_3042,N_2771,N_2985);
xnor U3043 (N_3043,N_2684,N_2864);
nor U3044 (N_3044,N_2717,N_2998);
nand U3045 (N_3045,N_2790,N_2567);
or U3046 (N_3046,N_2777,N_2565);
nand U3047 (N_3047,N_2716,N_2641);
and U3048 (N_3048,N_2728,N_2885);
nor U3049 (N_3049,N_2712,N_2637);
or U3050 (N_3050,N_2773,N_2840);
nor U3051 (N_3051,N_2704,N_2566);
or U3052 (N_3052,N_2756,N_2816);
nand U3053 (N_3053,N_2779,N_2927);
nor U3054 (N_3054,N_2829,N_2543);
nor U3055 (N_3055,N_2512,N_2786);
and U3056 (N_3056,N_2517,N_2977);
and U3057 (N_3057,N_2719,N_2803);
or U3058 (N_3058,N_2534,N_2930);
xor U3059 (N_3059,N_2735,N_2610);
or U3060 (N_3060,N_2563,N_2705);
or U3061 (N_3061,N_2966,N_2524);
nor U3062 (N_3062,N_2994,N_2801);
and U3063 (N_3063,N_2853,N_2878);
and U3064 (N_3064,N_2594,N_2963);
and U3065 (N_3065,N_2890,N_2876);
nand U3066 (N_3066,N_2972,N_2899);
or U3067 (N_3067,N_2753,N_2793);
xor U3068 (N_3068,N_2996,N_2544);
nor U3069 (N_3069,N_2647,N_2861);
and U3070 (N_3070,N_2969,N_2895);
and U3071 (N_3071,N_2957,N_2630);
nand U3072 (N_3072,N_2586,N_2622);
or U3073 (N_3073,N_2526,N_2854);
or U3074 (N_3074,N_2902,N_2549);
nor U3075 (N_3075,N_2749,N_2825);
or U3076 (N_3076,N_2676,N_2696);
and U3077 (N_3077,N_2990,N_2750);
or U3078 (N_3078,N_2655,N_2827);
nand U3079 (N_3079,N_2959,N_2656);
or U3080 (N_3080,N_2931,N_2690);
and U3081 (N_3081,N_2600,N_2673);
nor U3082 (N_3082,N_2891,N_2912);
xor U3083 (N_3083,N_2592,N_2557);
nor U3084 (N_3084,N_2652,N_2889);
nand U3085 (N_3085,N_2626,N_2869);
or U3086 (N_3086,N_2738,N_2525);
nor U3087 (N_3087,N_2733,N_2776);
nand U3088 (N_3088,N_2815,N_2604);
and U3089 (N_3089,N_2579,N_2778);
nor U3090 (N_3090,N_2692,N_2976);
nand U3091 (N_3091,N_2746,N_2634);
nor U3092 (N_3092,N_2882,N_2848);
xor U3093 (N_3093,N_2662,N_2693);
and U3094 (N_3094,N_2980,N_2686);
or U3095 (N_3095,N_2995,N_2667);
nand U3096 (N_3096,N_2883,N_2774);
or U3097 (N_3097,N_2699,N_2862);
nand U3098 (N_3098,N_2814,N_2860);
nand U3099 (N_3099,N_2986,N_2504);
xor U3100 (N_3100,N_2909,N_2709);
xnor U3101 (N_3101,N_2611,N_2648);
nor U3102 (N_3102,N_2946,N_2846);
nor U3103 (N_3103,N_2520,N_2865);
and U3104 (N_3104,N_2694,N_2540);
nand U3105 (N_3105,N_2799,N_2870);
nor U3106 (N_3106,N_2593,N_2700);
nor U3107 (N_3107,N_2747,N_2974);
nor U3108 (N_3108,N_2731,N_2620);
xnor U3109 (N_3109,N_2651,N_2950);
nand U3110 (N_3110,N_2675,N_2826);
nand U3111 (N_3111,N_2984,N_2828);
nor U3112 (N_3112,N_2988,N_2834);
and U3113 (N_3113,N_2555,N_2682);
and U3114 (N_3114,N_2997,N_2798);
and U3115 (N_3115,N_2708,N_2521);
and U3116 (N_3116,N_2741,N_2879);
nor U3117 (N_3117,N_2939,N_2880);
xor U3118 (N_3118,N_2925,N_2784);
and U3119 (N_3119,N_2888,N_2809);
nand U3120 (N_3120,N_2724,N_2609);
and U3121 (N_3121,N_2573,N_2797);
or U3122 (N_3122,N_2987,N_2649);
and U3123 (N_3123,N_2913,N_2810);
or U3124 (N_3124,N_2607,N_2729);
or U3125 (N_3125,N_2850,N_2760);
xor U3126 (N_3126,N_2669,N_2533);
nor U3127 (N_3127,N_2962,N_2551);
nor U3128 (N_3128,N_2761,N_2518);
xor U3129 (N_3129,N_2539,N_2991);
xor U3130 (N_3130,N_2585,N_2726);
and U3131 (N_3131,N_2943,N_2646);
or U3132 (N_3132,N_2887,N_2794);
and U3133 (N_3133,N_2614,N_2817);
and U3134 (N_3134,N_2918,N_2837);
and U3135 (N_3135,N_2624,N_2623);
nor U3136 (N_3136,N_2599,N_2581);
nor U3137 (N_3137,N_2500,N_2893);
nor U3138 (N_3138,N_2919,N_2863);
and U3139 (N_3139,N_2903,N_2742);
xnor U3140 (N_3140,N_2612,N_2781);
nand U3141 (N_3141,N_2688,N_2553);
nor U3142 (N_3142,N_2665,N_2552);
xnor U3143 (N_3143,N_2842,N_2775);
and U3144 (N_3144,N_2759,N_2993);
or U3145 (N_3145,N_2823,N_2920);
or U3146 (N_3146,N_2841,N_2528);
nand U3147 (N_3147,N_2510,N_2537);
nand U3148 (N_3148,N_2942,N_2572);
nand U3149 (N_3149,N_2833,N_2661);
nor U3150 (N_3150,N_2921,N_2664);
nor U3151 (N_3151,N_2772,N_2615);
or U3152 (N_3152,N_2922,N_2811);
nor U3153 (N_3153,N_2758,N_2847);
or U3154 (N_3154,N_2806,N_2767);
and U3155 (N_3155,N_2757,N_2859);
nand U3156 (N_3156,N_2770,N_2663);
nor U3157 (N_3157,N_2947,N_2783);
nor U3158 (N_3158,N_2632,N_2591);
and U3159 (N_3159,N_2713,N_2951);
or U3160 (N_3160,N_2898,N_2808);
or U3161 (N_3161,N_2670,N_2718);
or U3162 (N_3162,N_2564,N_2501);
and U3163 (N_3163,N_2621,N_2695);
nand U3164 (N_3164,N_2901,N_2844);
nand U3165 (N_3165,N_2723,N_2857);
or U3166 (N_3166,N_2653,N_2633);
and U3167 (N_3167,N_2792,N_2820);
nor U3168 (N_3168,N_2574,N_2725);
and U3169 (N_3169,N_2978,N_2542);
nand U3170 (N_3170,N_2560,N_2982);
nand U3171 (N_3171,N_2949,N_2769);
nand U3172 (N_3172,N_2740,N_2513);
and U3173 (N_3173,N_2577,N_2589);
nor U3174 (N_3174,N_2917,N_2576);
nand U3175 (N_3175,N_2523,N_2787);
nand U3176 (N_3176,N_2956,N_2849);
and U3177 (N_3177,N_2910,N_2536);
or U3178 (N_3178,N_2968,N_2782);
nand U3179 (N_3179,N_2788,N_2596);
and U3180 (N_3180,N_2698,N_2785);
or U3181 (N_3181,N_2955,N_2672);
nand U3182 (N_3182,N_2958,N_2597);
or U3183 (N_3183,N_2628,N_2999);
nand U3184 (N_3184,N_2804,N_2831);
nand U3185 (N_3185,N_2605,N_2743);
nor U3186 (N_3186,N_2855,N_2680);
nor U3187 (N_3187,N_2852,N_2685);
or U3188 (N_3188,N_2691,N_2766);
and U3189 (N_3189,N_2940,N_2734);
and U3190 (N_3190,N_2754,N_2822);
nand U3191 (N_3191,N_2948,N_2643);
or U3192 (N_3192,N_2702,N_2657);
and U3193 (N_3193,N_2851,N_2707);
or U3194 (N_3194,N_2789,N_2964);
nor U3195 (N_3195,N_2935,N_2638);
xor U3196 (N_3196,N_2755,N_2703);
nor U3197 (N_3197,N_2751,N_2687);
nor U3198 (N_3198,N_2944,N_2780);
and U3199 (N_3199,N_2845,N_2507);
nand U3200 (N_3200,N_2561,N_2683);
nand U3201 (N_3201,N_2580,N_2904);
nand U3202 (N_3202,N_2745,N_2559);
and U3203 (N_3203,N_2575,N_2881);
nor U3204 (N_3204,N_2971,N_2954);
nand U3205 (N_3205,N_2936,N_2896);
nand U3206 (N_3206,N_2710,N_2677);
nor U3207 (N_3207,N_2527,N_2625);
nand U3208 (N_3208,N_2926,N_2867);
nand U3209 (N_3209,N_2508,N_2908);
or U3210 (N_3210,N_2929,N_2511);
xnor U3211 (N_3211,N_2516,N_2681);
and U3212 (N_3212,N_2578,N_2711);
nand U3213 (N_3213,N_2509,N_2529);
or U3214 (N_3214,N_2635,N_2514);
nor U3215 (N_3215,N_2640,N_2981);
and U3216 (N_3216,N_2679,N_2802);
nor U3217 (N_3217,N_2631,N_2838);
nand U3218 (N_3218,N_2547,N_2541);
and U3219 (N_3219,N_2807,N_2915);
or U3220 (N_3220,N_2659,N_2671);
nor U3221 (N_3221,N_2714,N_2619);
xor U3222 (N_3222,N_2914,N_2992);
or U3223 (N_3223,N_2636,N_2989);
nor U3224 (N_3224,N_2689,N_2924);
or U3225 (N_3225,N_2824,N_2660);
nand U3226 (N_3226,N_2800,N_2960);
nor U3227 (N_3227,N_2658,N_2953);
and U3228 (N_3228,N_2583,N_2732);
or U3229 (N_3229,N_2650,N_2762);
or U3230 (N_3230,N_2928,N_2603);
nand U3231 (N_3231,N_2897,N_2697);
nand U3232 (N_3232,N_2900,N_2608);
nor U3233 (N_3233,N_2961,N_2873);
xor U3234 (N_3234,N_2973,N_2570);
and U3235 (N_3235,N_2674,N_2642);
xor U3236 (N_3236,N_2934,N_2932);
and U3237 (N_3237,N_2720,N_2970);
nor U3238 (N_3238,N_2550,N_2791);
and U3239 (N_3239,N_2519,N_2530);
xor U3240 (N_3240,N_2894,N_2613);
and U3241 (N_3241,N_2562,N_2590);
or U3242 (N_3242,N_2506,N_2818);
or U3243 (N_3243,N_2739,N_2582);
nor U3244 (N_3244,N_2967,N_2522);
and U3245 (N_3245,N_2601,N_2830);
nor U3246 (N_3246,N_2748,N_2933);
nand U3247 (N_3247,N_2965,N_2866);
and U3248 (N_3248,N_2730,N_2858);
nor U3249 (N_3249,N_2569,N_2535);
or U3250 (N_3250,N_2841,N_2997);
nand U3251 (N_3251,N_2779,N_2949);
or U3252 (N_3252,N_2547,N_2627);
xnor U3253 (N_3253,N_2644,N_2727);
or U3254 (N_3254,N_2763,N_2895);
or U3255 (N_3255,N_2858,N_2840);
nand U3256 (N_3256,N_2708,N_2538);
xnor U3257 (N_3257,N_2778,N_2814);
nand U3258 (N_3258,N_2801,N_2512);
and U3259 (N_3259,N_2581,N_2540);
nand U3260 (N_3260,N_2754,N_2777);
xor U3261 (N_3261,N_2733,N_2510);
nand U3262 (N_3262,N_2729,N_2769);
or U3263 (N_3263,N_2615,N_2754);
and U3264 (N_3264,N_2854,N_2959);
xnor U3265 (N_3265,N_2710,N_2964);
or U3266 (N_3266,N_2650,N_2655);
and U3267 (N_3267,N_2558,N_2808);
nor U3268 (N_3268,N_2805,N_2786);
and U3269 (N_3269,N_2932,N_2838);
nand U3270 (N_3270,N_2649,N_2622);
and U3271 (N_3271,N_2694,N_2871);
and U3272 (N_3272,N_2607,N_2945);
xor U3273 (N_3273,N_2626,N_2990);
and U3274 (N_3274,N_2719,N_2529);
nand U3275 (N_3275,N_2776,N_2573);
and U3276 (N_3276,N_2647,N_2520);
nand U3277 (N_3277,N_2525,N_2909);
xor U3278 (N_3278,N_2589,N_2530);
nand U3279 (N_3279,N_2589,N_2799);
nor U3280 (N_3280,N_2997,N_2598);
xor U3281 (N_3281,N_2573,N_2666);
and U3282 (N_3282,N_2925,N_2778);
or U3283 (N_3283,N_2527,N_2771);
or U3284 (N_3284,N_2772,N_2732);
or U3285 (N_3285,N_2775,N_2819);
nor U3286 (N_3286,N_2874,N_2896);
and U3287 (N_3287,N_2852,N_2668);
nand U3288 (N_3288,N_2830,N_2539);
and U3289 (N_3289,N_2836,N_2929);
and U3290 (N_3290,N_2807,N_2874);
and U3291 (N_3291,N_2822,N_2592);
nand U3292 (N_3292,N_2595,N_2893);
or U3293 (N_3293,N_2736,N_2571);
nand U3294 (N_3294,N_2721,N_2698);
xnor U3295 (N_3295,N_2593,N_2681);
and U3296 (N_3296,N_2688,N_2796);
nor U3297 (N_3297,N_2745,N_2930);
nand U3298 (N_3298,N_2503,N_2805);
or U3299 (N_3299,N_2966,N_2999);
nor U3300 (N_3300,N_2605,N_2802);
xnor U3301 (N_3301,N_2855,N_2848);
and U3302 (N_3302,N_2849,N_2648);
or U3303 (N_3303,N_2869,N_2670);
or U3304 (N_3304,N_2651,N_2874);
nor U3305 (N_3305,N_2896,N_2918);
nor U3306 (N_3306,N_2788,N_2730);
nand U3307 (N_3307,N_2918,N_2863);
and U3308 (N_3308,N_2858,N_2742);
nor U3309 (N_3309,N_2975,N_2606);
nor U3310 (N_3310,N_2792,N_2559);
nand U3311 (N_3311,N_2740,N_2924);
nand U3312 (N_3312,N_2859,N_2944);
nand U3313 (N_3313,N_2794,N_2690);
nand U3314 (N_3314,N_2822,N_2949);
and U3315 (N_3315,N_2736,N_2710);
nor U3316 (N_3316,N_2637,N_2881);
and U3317 (N_3317,N_2742,N_2927);
nor U3318 (N_3318,N_2772,N_2814);
xor U3319 (N_3319,N_2520,N_2813);
nand U3320 (N_3320,N_2782,N_2743);
or U3321 (N_3321,N_2564,N_2971);
nor U3322 (N_3322,N_2593,N_2758);
nand U3323 (N_3323,N_2852,N_2581);
nand U3324 (N_3324,N_2662,N_2861);
nor U3325 (N_3325,N_2512,N_2597);
nand U3326 (N_3326,N_2728,N_2625);
nor U3327 (N_3327,N_2602,N_2802);
nand U3328 (N_3328,N_2642,N_2923);
nor U3329 (N_3329,N_2809,N_2685);
nand U3330 (N_3330,N_2601,N_2518);
and U3331 (N_3331,N_2863,N_2984);
and U3332 (N_3332,N_2677,N_2778);
nand U3333 (N_3333,N_2741,N_2582);
xnor U3334 (N_3334,N_2707,N_2881);
and U3335 (N_3335,N_2980,N_2864);
nand U3336 (N_3336,N_2509,N_2625);
and U3337 (N_3337,N_2659,N_2688);
and U3338 (N_3338,N_2974,N_2671);
nand U3339 (N_3339,N_2974,N_2958);
nor U3340 (N_3340,N_2607,N_2834);
nand U3341 (N_3341,N_2596,N_2800);
nand U3342 (N_3342,N_2553,N_2839);
and U3343 (N_3343,N_2632,N_2925);
nand U3344 (N_3344,N_2617,N_2777);
xnor U3345 (N_3345,N_2584,N_2648);
nand U3346 (N_3346,N_2799,N_2611);
xor U3347 (N_3347,N_2935,N_2506);
nor U3348 (N_3348,N_2706,N_2702);
nand U3349 (N_3349,N_2736,N_2735);
or U3350 (N_3350,N_2958,N_2708);
nor U3351 (N_3351,N_2911,N_2919);
nand U3352 (N_3352,N_2822,N_2988);
nor U3353 (N_3353,N_2993,N_2714);
and U3354 (N_3354,N_2580,N_2927);
nand U3355 (N_3355,N_2517,N_2716);
nand U3356 (N_3356,N_2857,N_2955);
and U3357 (N_3357,N_2724,N_2705);
or U3358 (N_3358,N_2504,N_2743);
nor U3359 (N_3359,N_2808,N_2991);
or U3360 (N_3360,N_2591,N_2539);
nand U3361 (N_3361,N_2595,N_2890);
or U3362 (N_3362,N_2674,N_2847);
xor U3363 (N_3363,N_2539,N_2523);
nor U3364 (N_3364,N_2804,N_2799);
nand U3365 (N_3365,N_2611,N_2828);
nor U3366 (N_3366,N_2919,N_2684);
nand U3367 (N_3367,N_2842,N_2777);
and U3368 (N_3368,N_2805,N_2608);
nor U3369 (N_3369,N_2738,N_2827);
or U3370 (N_3370,N_2912,N_2940);
nand U3371 (N_3371,N_2978,N_2706);
nor U3372 (N_3372,N_2935,N_2708);
and U3373 (N_3373,N_2577,N_2738);
nor U3374 (N_3374,N_2840,N_2524);
or U3375 (N_3375,N_2570,N_2957);
nand U3376 (N_3376,N_2535,N_2724);
nand U3377 (N_3377,N_2779,N_2775);
nand U3378 (N_3378,N_2743,N_2935);
nand U3379 (N_3379,N_2750,N_2639);
nor U3380 (N_3380,N_2677,N_2808);
nand U3381 (N_3381,N_2968,N_2636);
or U3382 (N_3382,N_2720,N_2740);
or U3383 (N_3383,N_2779,N_2962);
nor U3384 (N_3384,N_2662,N_2727);
nand U3385 (N_3385,N_2570,N_2869);
or U3386 (N_3386,N_2524,N_2995);
or U3387 (N_3387,N_2500,N_2636);
or U3388 (N_3388,N_2545,N_2531);
nor U3389 (N_3389,N_2884,N_2842);
xnor U3390 (N_3390,N_2776,N_2606);
nand U3391 (N_3391,N_2844,N_2742);
or U3392 (N_3392,N_2821,N_2673);
nor U3393 (N_3393,N_2917,N_2942);
nand U3394 (N_3394,N_2581,N_2668);
or U3395 (N_3395,N_2710,N_2980);
or U3396 (N_3396,N_2715,N_2526);
or U3397 (N_3397,N_2633,N_2776);
or U3398 (N_3398,N_2993,N_2970);
and U3399 (N_3399,N_2801,N_2838);
nor U3400 (N_3400,N_2968,N_2987);
nand U3401 (N_3401,N_2667,N_2616);
xnor U3402 (N_3402,N_2738,N_2691);
nand U3403 (N_3403,N_2859,N_2622);
xor U3404 (N_3404,N_2667,N_2941);
nand U3405 (N_3405,N_2634,N_2961);
and U3406 (N_3406,N_2745,N_2628);
nor U3407 (N_3407,N_2824,N_2538);
or U3408 (N_3408,N_2540,N_2737);
or U3409 (N_3409,N_2634,N_2890);
xor U3410 (N_3410,N_2862,N_2846);
or U3411 (N_3411,N_2702,N_2740);
or U3412 (N_3412,N_2790,N_2794);
nor U3413 (N_3413,N_2739,N_2821);
nor U3414 (N_3414,N_2663,N_2751);
nand U3415 (N_3415,N_2528,N_2609);
and U3416 (N_3416,N_2759,N_2840);
xor U3417 (N_3417,N_2584,N_2892);
nand U3418 (N_3418,N_2824,N_2982);
and U3419 (N_3419,N_2526,N_2563);
nor U3420 (N_3420,N_2525,N_2999);
and U3421 (N_3421,N_2702,N_2687);
xor U3422 (N_3422,N_2640,N_2726);
or U3423 (N_3423,N_2910,N_2683);
nand U3424 (N_3424,N_2923,N_2947);
nor U3425 (N_3425,N_2962,N_2866);
and U3426 (N_3426,N_2560,N_2657);
or U3427 (N_3427,N_2855,N_2743);
nand U3428 (N_3428,N_2561,N_2855);
or U3429 (N_3429,N_2999,N_2520);
and U3430 (N_3430,N_2635,N_2911);
and U3431 (N_3431,N_2667,N_2697);
and U3432 (N_3432,N_2821,N_2900);
xnor U3433 (N_3433,N_2775,N_2669);
and U3434 (N_3434,N_2638,N_2643);
or U3435 (N_3435,N_2900,N_2568);
nand U3436 (N_3436,N_2807,N_2544);
and U3437 (N_3437,N_2736,N_2954);
nor U3438 (N_3438,N_2855,N_2879);
nor U3439 (N_3439,N_2865,N_2747);
xnor U3440 (N_3440,N_2674,N_2912);
nand U3441 (N_3441,N_2963,N_2945);
and U3442 (N_3442,N_2853,N_2881);
or U3443 (N_3443,N_2949,N_2757);
nor U3444 (N_3444,N_2535,N_2517);
nand U3445 (N_3445,N_2890,N_2560);
and U3446 (N_3446,N_2700,N_2907);
nor U3447 (N_3447,N_2898,N_2509);
or U3448 (N_3448,N_2939,N_2758);
and U3449 (N_3449,N_2635,N_2637);
and U3450 (N_3450,N_2767,N_2721);
xor U3451 (N_3451,N_2960,N_2871);
nor U3452 (N_3452,N_2932,N_2623);
and U3453 (N_3453,N_2638,N_2870);
and U3454 (N_3454,N_2525,N_2634);
and U3455 (N_3455,N_2850,N_2943);
nor U3456 (N_3456,N_2989,N_2890);
nor U3457 (N_3457,N_2694,N_2576);
and U3458 (N_3458,N_2770,N_2633);
xnor U3459 (N_3459,N_2994,N_2765);
nand U3460 (N_3460,N_2658,N_2877);
or U3461 (N_3461,N_2713,N_2696);
nand U3462 (N_3462,N_2898,N_2745);
and U3463 (N_3463,N_2946,N_2719);
and U3464 (N_3464,N_2532,N_2505);
or U3465 (N_3465,N_2706,N_2870);
and U3466 (N_3466,N_2903,N_2711);
nor U3467 (N_3467,N_2810,N_2824);
and U3468 (N_3468,N_2671,N_2589);
nand U3469 (N_3469,N_2829,N_2891);
nand U3470 (N_3470,N_2997,N_2635);
xor U3471 (N_3471,N_2904,N_2599);
nand U3472 (N_3472,N_2889,N_2788);
nand U3473 (N_3473,N_2699,N_2735);
or U3474 (N_3474,N_2954,N_2821);
nor U3475 (N_3475,N_2853,N_2827);
and U3476 (N_3476,N_2746,N_2881);
nand U3477 (N_3477,N_2719,N_2874);
nand U3478 (N_3478,N_2994,N_2802);
or U3479 (N_3479,N_2959,N_2635);
nand U3480 (N_3480,N_2793,N_2595);
and U3481 (N_3481,N_2992,N_2713);
and U3482 (N_3482,N_2572,N_2780);
nand U3483 (N_3483,N_2940,N_2744);
or U3484 (N_3484,N_2522,N_2977);
xnor U3485 (N_3485,N_2668,N_2606);
and U3486 (N_3486,N_2984,N_2766);
nor U3487 (N_3487,N_2990,N_2571);
nand U3488 (N_3488,N_2608,N_2911);
nand U3489 (N_3489,N_2516,N_2937);
nand U3490 (N_3490,N_2547,N_2974);
xnor U3491 (N_3491,N_2792,N_2952);
nand U3492 (N_3492,N_2787,N_2593);
or U3493 (N_3493,N_2685,N_2789);
or U3494 (N_3494,N_2576,N_2889);
and U3495 (N_3495,N_2527,N_2870);
nand U3496 (N_3496,N_2509,N_2502);
nand U3497 (N_3497,N_2563,N_2933);
nand U3498 (N_3498,N_2565,N_2985);
nor U3499 (N_3499,N_2857,N_2544);
or U3500 (N_3500,N_3334,N_3149);
nand U3501 (N_3501,N_3241,N_3018);
nand U3502 (N_3502,N_3444,N_3299);
nor U3503 (N_3503,N_3128,N_3374);
nand U3504 (N_3504,N_3431,N_3331);
nor U3505 (N_3505,N_3207,N_3085);
nand U3506 (N_3506,N_3349,N_3252);
or U3507 (N_3507,N_3371,N_3411);
nor U3508 (N_3508,N_3094,N_3142);
nand U3509 (N_3509,N_3441,N_3469);
nand U3510 (N_3510,N_3002,N_3466);
nor U3511 (N_3511,N_3440,N_3226);
and U3512 (N_3512,N_3135,N_3329);
nand U3513 (N_3513,N_3141,N_3393);
or U3514 (N_3514,N_3247,N_3130);
or U3515 (N_3515,N_3193,N_3033);
or U3516 (N_3516,N_3176,N_3109);
and U3517 (N_3517,N_3243,N_3035);
or U3518 (N_3518,N_3306,N_3422);
and U3519 (N_3519,N_3391,N_3173);
nor U3520 (N_3520,N_3407,N_3484);
or U3521 (N_3521,N_3446,N_3447);
nor U3522 (N_3522,N_3489,N_3160);
or U3523 (N_3523,N_3114,N_3303);
or U3524 (N_3524,N_3192,N_3316);
nor U3525 (N_3525,N_3244,N_3063);
and U3526 (N_3526,N_3123,N_3106);
nor U3527 (N_3527,N_3433,N_3011);
and U3528 (N_3528,N_3101,N_3464);
or U3529 (N_3529,N_3381,N_3216);
or U3530 (N_3530,N_3387,N_3335);
and U3531 (N_3531,N_3154,N_3091);
nand U3532 (N_3532,N_3443,N_3185);
nand U3533 (N_3533,N_3165,N_3428);
nor U3534 (N_3534,N_3228,N_3188);
or U3535 (N_3535,N_3147,N_3249);
nor U3536 (N_3536,N_3066,N_3292);
nand U3537 (N_3537,N_3022,N_3320);
or U3538 (N_3538,N_3499,N_3020);
nand U3539 (N_3539,N_3352,N_3268);
xnor U3540 (N_3540,N_3060,N_3157);
xnor U3541 (N_3541,N_3198,N_3289);
or U3542 (N_3542,N_3278,N_3458);
or U3543 (N_3543,N_3168,N_3449);
nor U3544 (N_3544,N_3144,N_3494);
and U3545 (N_3545,N_3223,N_3071);
and U3546 (N_3546,N_3034,N_3090);
nor U3547 (N_3547,N_3166,N_3392);
and U3548 (N_3548,N_3263,N_3336);
xnor U3549 (N_3549,N_3257,N_3108);
nor U3550 (N_3550,N_3369,N_3242);
or U3551 (N_3551,N_3430,N_3283);
or U3552 (N_3552,N_3491,N_3016);
nor U3553 (N_3553,N_3382,N_3227);
and U3554 (N_3554,N_3184,N_3010);
nand U3555 (N_3555,N_3052,N_3478);
xor U3556 (N_3556,N_3155,N_3452);
xnor U3557 (N_3557,N_3080,N_3097);
nor U3558 (N_3558,N_3318,N_3426);
nor U3559 (N_3559,N_3246,N_3325);
and U3560 (N_3560,N_3483,N_3277);
nor U3561 (N_3561,N_3412,N_3432);
or U3562 (N_3562,N_3300,N_3055);
nand U3563 (N_3563,N_3008,N_3049);
nand U3564 (N_3564,N_3279,N_3418);
and U3565 (N_3565,N_3107,N_3161);
xor U3566 (N_3566,N_3459,N_3027);
and U3567 (N_3567,N_3272,N_3420);
nor U3568 (N_3568,N_3138,N_3455);
nand U3569 (N_3569,N_3397,N_3140);
or U3570 (N_3570,N_3180,N_3493);
nand U3571 (N_3571,N_3006,N_3380);
and U3572 (N_3572,N_3041,N_3074);
nor U3573 (N_3573,N_3388,N_3386);
and U3574 (N_3574,N_3231,N_3445);
nand U3575 (N_3575,N_3059,N_3124);
xor U3576 (N_3576,N_3088,N_3248);
nor U3577 (N_3577,N_3222,N_3442);
or U3578 (N_3578,N_3462,N_3048);
or U3579 (N_3579,N_3404,N_3133);
and U3580 (N_3580,N_3347,N_3139);
nor U3581 (N_3581,N_3187,N_3217);
nor U3582 (N_3582,N_3364,N_3245);
or U3583 (N_3583,N_3084,N_3062);
nand U3584 (N_3584,N_3186,N_3396);
nor U3585 (N_3585,N_3164,N_3379);
nor U3586 (N_3586,N_3170,N_3288);
or U3587 (N_3587,N_3307,N_3092);
or U3588 (N_3588,N_3014,N_3051);
and U3589 (N_3589,N_3050,N_3351);
nor U3590 (N_3590,N_3073,N_3212);
nor U3591 (N_3591,N_3367,N_3438);
or U3592 (N_3592,N_3281,N_3363);
nor U3593 (N_3593,N_3079,N_3030);
nand U3594 (N_3594,N_3439,N_3450);
nor U3595 (N_3595,N_3159,N_3390);
or U3596 (N_3596,N_3009,N_3043);
nand U3597 (N_3597,N_3456,N_3251);
nor U3598 (N_3598,N_3415,N_3498);
xor U3599 (N_3599,N_3036,N_3267);
or U3600 (N_3600,N_3471,N_3023);
and U3601 (N_3601,N_3204,N_3312);
nor U3602 (N_3602,N_3409,N_3470);
or U3603 (N_3603,N_3116,N_3271);
or U3604 (N_3604,N_3293,N_3465);
nand U3605 (N_3605,N_3044,N_3136);
or U3606 (N_3606,N_3389,N_3287);
nor U3607 (N_3607,N_3341,N_3476);
or U3608 (N_3608,N_3209,N_3342);
xor U3609 (N_3609,N_3496,N_3308);
nand U3610 (N_3610,N_3121,N_3276);
nor U3611 (N_3611,N_3148,N_3310);
or U3612 (N_3612,N_3239,N_3110);
or U3613 (N_3613,N_3229,N_3261);
and U3614 (N_3614,N_3032,N_3007);
nor U3615 (N_3615,N_3453,N_3067);
and U3616 (N_3616,N_3285,N_3435);
and U3617 (N_3617,N_3169,N_3305);
and U3618 (N_3618,N_3368,N_3201);
and U3619 (N_3619,N_3301,N_3211);
and U3620 (N_3620,N_3179,N_3078);
or U3621 (N_3621,N_3053,N_3240);
or U3622 (N_3622,N_3427,N_3421);
or U3623 (N_3623,N_3146,N_3345);
xnor U3624 (N_3624,N_3189,N_3039);
and U3625 (N_3625,N_3087,N_3061);
and U3626 (N_3626,N_3457,N_3102);
or U3627 (N_3627,N_3359,N_3410);
nor U3628 (N_3628,N_3221,N_3385);
xnor U3629 (N_3629,N_3100,N_3357);
or U3630 (N_3630,N_3025,N_3081);
nor U3631 (N_3631,N_3485,N_3394);
or U3632 (N_3632,N_3089,N_3400);
and U3633 (N_3633,N_3236,N_3330);
or U3634 (N_3634,N_3482,N_3468);
and U3635 (N_3635,N_3042,N_3376);
and U3636 (N_3636,N_3406,N_3467);
or U3637 (N_3637,N_3298,N_3125);
nor U3638 (N_3638,N_3026,N_3197);
nor U3639 (N_3639,N_3355,N_3448);
nand U3640 (N_3640,N_3151,N_3000);
xor U3641 (N_3641,N_3321,N_3181);
nand U3642 (N_3642,N_3233,N_3436);
xor U3643 (N_3643,N_3361,N_3461);
and U3644 (N_3644,N_3224,N_3302);
or U3645 (N_3645,N_3474,N_3183);
xnor U3646 (N_3646,N_3434,N_3132);
and U3647 (N_3647,N_3120,N_3045);
or U3648 (N_3648,N_3405,N_3237);
nand U3649 (N_3649,N_3322,N_3037);
and U3650 (N_3650,N_3378,N_3280);
or U3651 (N_3651,N_3343,N_3333);
nor U3652 (N_3652,N_3323,N_3419);
xor U3653 (N_3653,N_3127,N_3117);
or U3654 (N_3654,N_3486,N_3214);
nor U3655 (N_3655,N_3064,N_3260);
or U3656 (N_3656,N_3480,N_3103);
nand U3657 (N_3657,N_3225,N_3111);
and U3658 (N_3658,N_3253,N_3296);
nand U3659 (N_3659,N_3344,N_3425);
and U3660 (N_3660,N_3354,N_3319);
or U3661 (N_3661,N_3338,N_3024);
nor U3662 (N_3662,N_3038,N_3005);
and U3663 (N_3663,N_3099,N_3372);
nand U3664 (N_3664,N_3265,N_3028);
xnor U3665 (N_3665,N_3399,N_3340);
or U3666 (N_3666,N_3473,N_3058);
nor U3667 (N_3667,N_3295,N_3332);
or U3668 (N_3668,N_3460,N_3315);
xor U3669 (N_3669,N_3294,N_3304);
and U3670 (N_3670,N_3375,N_3273);
nand U3671 (N_3671,N_3373,N_3266);
or U3672 (N_3672,N_3402,N_3238);
xor U3673 (N_3673,N_3076,N_3202);
or U3674 (N_3674,N_3029,N_3213);
nand U3675 (N_3675,N_3270,N_3401);
or U3676 (N_3676,N_3001,N_3414);
nor U3677 (N_3677,N_3054,N_3490);
and U3678 (N_3678,N_3200,N_3119);
nand U3679 (N_3679,N_3398,N_3047);
and U3680 (N_3680,N_3365,N_3370);
nor U3681 (N_3681,N_3255,N_3153);
or U3682 (N_3682,N_3384,N_3454);
xor U3683 (N_3683,N_3488,N_3196);
nand U3684 (N_3684,N_3337,N_3015);
nor U3685 (N_3685,N_3360,N_3264);
nor U3686 (N_3686,N_3070,N_3205);
nand U3687 (N_3687,N_3395,N_3259);
nand U3688 (N_3688,N_3291,N_3178);
and U3689 (N_3689,N_3152,N_3250);
nand U3690 (N_3690,N_3040,N_3069);
nand U3691 (N_3691,N_3122,N_3218);
or U3692 (N_3692,N_3056,N_3230);
or U3693 (N_3693,N_3096,N_3383);
or U3694 (N_3694,N_3477,N_3328);
and U3695 (N_3695,N_3215,N_3065);
or U3696 (N_3696,N_3126,N_3417);
or U3697 (N_3697,N_3235,N_3134);
and U3698 (N_3698,N_3309,N_3115);
nor U3699 (N_3699,N_3451,N_3377);
or U3700 (N_3700,N_3068,N_3077);
or U3701 (N_3701,N_3083,N_3326);
and U3702 (N_3702,N_3346,N_3129);
xor U3703 (N_3703,N_3156,N_3017);
xnor U3704 (N_3704,N_3492,N_3019);
xnor U3705 (N_3705,N_3472,N_3282);
nand U3706 (N_3706,N_3182,N_3137);
nand U3707 (N_3707,N_3093,N_3297);
xnor U3708 (N_3708,N_3172,N_3234);
and U3709 (N_3709,N_3208,N_3075);
nor U3710 (N_3710,N_3175,N_3497);
or U3711 (N_3711,N_3113,N_3269);
nand U3712 (N_3712,N_3275,N_3311);
nand U3713 (N_3713,N_3190,N_3162);
nor U3714 (N_3714,N_3317,N_3284);
nand U3715 (N_3715,N_3313,N_3004);
nor U3716 (N_3716,N_3163,N_3104);
or U3717 (N_3717,N_3286,N_3327);
or U3718 (N_3718,N_3105,N_3424);
or U3719 (N_3719,N_3254,N_3481);
xnor U3720 (N_3720,N_3194,N_3290);
nand U3721 (N_3721,N_3362,N_3082);
and U3722 (N_3722,N_3013,N_3219);
nor U3723 (N_3723,N_3487,N_3206);
nand U3724 (N_3724,N_3031,N_3046);
or U3725 (N_3725,N_3350,N_3437);
and U3726 (N_3726,N_3098,N_3171);
and U3727 (N_3727,N_3158,N_3167);
or U3728 (N_3728,N_3274,N_3210);
nor U3729 (N_3729,N_3324,N_3131);
nand U3730 (N_3730,N_3086,N_3177);
and U3731 (N_3731,N_3003,N_3203);
and U3732 (N_3732,N_3479,N_3150);
xnor U3733 (N_3733,N_3339,N_3429);
xor U3734 (N_3734,N_3358,N_3174);
and U3735 (N_3735,N_3262,N_3258);
or U3736 (N_3736,N_3021,N_3232);
xnor U3737 (N_3737,N_3145,N_3220);
nand U3738 (N_3738,N_3495,N_3195);
nor U3739 (N_3739,N_3356,N_3095);
nand U3740 (N_3740,N_3423,N_3416);
nor U3741 (N_3741,N_3143,N_3463);
xnor U3742 (N_3742,N_3314,N_3348);
and U3743 (N_3743,N_3118,N_3112);
or U3744 (N_3744,N_3413,N_3403);
nor U3745 (N_3745,N_3072,N_3408);
nor U3746 (N_3746,N_3199,N_3191);
or U3747 (N_3747,N_3366,N_3012);
nor U3748 (N_3748,N_3353,N_3057);
nor U3749 (N_3749,N_3256,N_3475);
nand U3750 (N_3750,N_3083,N_3436);
xnor U3751 (N_3751,N_3221,N_3001);
nor U3752 (N_3752,N_3245,N_3227);
xor U3753 (N_3753,N_3085,N_3309);
or U3754 (N_3754,N_3492,N_3367);
xnor U3755 (N_3755,N_3158,N_3094);
nand U3756 (N_3756,N_3137,N_3324);
and U3757 (N_3757,N_3156,N_3351);
nand U3758 (N_3758,N_3014,N_3077);
xnor U3759 (N_3759,N_3013,N_3030);
nand U3760 (N_3760,N_3242,N_3234);
nand U3761 (N_3761,N_3129,N_3005);
nor U3762 (N_3762,N_3252,N_3109);
and U3763 (N_3763,N_3227,N_3021);
or U3764 (N_3764,N_3164,N_3122);
and U3765 (N_3765,N_3484,N_3486);
nand U3766 (N_3766,N_3170,N_3458);
xnor U3767 (N_3767,N_3229,N_3169);
nand U3768 (N_3768,N_3039,N_3377);
nor U3769 (N_3769,N_3286,N_3438);
and U3770 (N_3770,N_3152,N_3236);
xor U3771 (N_3771,N_3237,N_3102);
nand U3772 (N_3772,N_3455,N_3363);
nor U3773 (N_3773,N_3060,N_3024);
and U3774 (N_3774,N_3403,N_3207);
nand U3775 (N_3775,N_3032,N_3146);
nand U3776 (N_3776,N_3341,N_3443);
and U3777 (N_3777,N_3299,N_3324);
nor U3778 (N_3778,N_3301,N_3252);
or U3779 (N_3779,N_3393,N_3411);
xnor U3780 (N_3780,N_3278,N_3357);
nor U3781 (N_3781,N_3037,N_3352);
and U3782 (N_3782,N_3323,N_3047);
nor U3783 (N_3783,N_3077,N_3367);
xnor U3784 (N_3784,N_3169,N_3211);
nand U3785 (N_3785,N_3002,N_3467);
nor U3786 (N_3786,N_3094,N_3481);
nand U3787 (N_3787,N_3059,N_3227);
xnor U3788 (N_3788,N_3226,N_3114);
or U3789 (N_3789,N_3422,N_3349);
nand U3790 (N_3790,N_3238,N_3173);
nor U3791 (N_3791,N_3241,N_3233);
and U3792 (N_3792,N_3293,N_3383);
nor U3793 (N_3793,N_3012,N_3216);
and U3794 (N_3794,N_3444,N_3428);
nand U3795 (N_3795,N_3097,N_3211);
or U3796 (N_3796,N_3338,N_3420);
nor U3797 (N_3797,N_3396,N_3488);
nand U3798 (N_3798,N_3032,N_3448);
or U3799 (N_3799,N_3267,N_3344);
and U3800 (N_3800,N_3298,N_3252);
xor U3801 (N_3801,N_3203,N_3422);
nor U3802 (N_3802,N_3273,N_3382);
or U3803 (N_3803,N_3494,N_3206);
and U3804 (N_3804,N_3240,N_3354);
xor U3805 (N_3805,N_3084,N_3456);
and U3806 (N_3806,N_3086,N_3225);
or U3807 (N_3807,N_3335,N_3378);
nor U3808 (N_3808,N_3081,N_3382);
nor U3809 (N_3809,N_3186,N_3246);
or U3810 (N_3810,N_3162,N_3340);
nand U3811 (N_3811,N_3016,N_3144);
nand U3812 (N_3812,N_3200,N_3463);
nor U3813 (N_3813,N_3076,N_3271);
or U3814 (N_3814,N_3083,N_3401);
nand U3815 (N_3815,N_3422,N_3165);
xnor U3816 (N_3816,N_3051,N_3053);
or U3817 (N_3817,N_3096,N_3000);
and U3818 (N_3818,N_3080,N_3433);
and U3819 (N_3819,N_3092,N_3267);
or U3820 (N_3820,N_3273,N_3431);
xnor U3821 (N_3821,N_3194,N_3226);
and U3822 (N_3822,N_3359,N_3093);
nand U3823 (N_3823,N_3122,N_3284);
nand U3824 (N_3824,N_3169,N_3328);
nand U3825 (N_3825,N_3350,N_3223);
or U3826 (N_3826,N_3385,N_3400);
and U3827 (N_3827,N_3474,N_3487);
and U3828 (N_3828,N_3046,N_3092);
and U3829 (N_3829,N_3458,N_3286);
nand U3830 (N_3830,N_3124,N_3194);
nor U3831 (N_3831,N_3206,N_3470);
or U3832 (N_3832,N_3164,N_3169);
and U3833 (N_3833,N_3350,N_3252);
and U3834 (N_3834,N_3422,N_3360);
nor U3835 (N_3835,N_3101,N_3232);
and U3836 (N_3836,N_3283,N_3271);
nor U3837 (N_3837,N_3432,N_3067);
nand U3838 (N_3838,N_3194,N_3144);
or U3839 (N_3839,N_3359,N_3069);
xor U3840 (N_3840,N_3052,N_3177);
and U3841 (N_3841,N_3232,N_3374);
xnor U3842 (N_3842,N_3478,N_3196);
nor U3843 (N_3843,N_3423,N_3294);
and U3844 (N_3844,N_3076,N_3206);
xor U3845 (N_3845,N_3209,N_3139);
nor U3846 (N_3846,N_3162,N_3208);
nor U3847 (N_3847,N_3352,N_3356);
nand U3848 (N_3848,N_3274,N_3389);
nor U3849 (N_3849,N_3283,N_3083);
nor U3850 (N_3850,N_3211,N_3373);
and U3851 (N_3851,N_3225,N_3424);
or U3852 (N_3852,N_3246,N_3014);
and U3853 (N_3853,N_3445,N_3448);
nand U3854 (N_3854,N_3033,N_3147);
nand U3855 (N_3855,N_3102,N_3085);
nand U3856 (N_3856,N_3263,N_3430);
and U3857 (N_3857,N_3294,N_3213);
or U3858 (N_3858,N_3331,N_3054);
nor U3859 (N_3859,N_3468,N_3405);
nand U3860 (N_3860,N_3097,N_3345);
and U3861 (N_3861,N_3453,N_3207);
and U3862 (N_3862,N_3340,N_3187);
and U3863 (N_3863,N_3274,N_3062);
and U3864 (N_3864,N_3463,N_3079);
or U3865 (N_3865,N_3447,N_3117);
and U3866 (N_3866,N_3202,N_3418);
nand U3867 (N_3867,N_3382,N_3097);
or U3868 (N_3868,N_3105,N_3165);
and U3869 (N_3869,N_3015,N_3246);
nand U3870 (N_3870,N_3192,N_3221);
or U3871 (N_3871,N_3276,N_3042);
nand U3872 (N_3872,N_3487,N_3459);
nor U3873 (N_3873,N_3446,N_3471);
nor U3874 (N_3874,N_3247,N_3234);
and U3875 (N_3875,N_3297,N_3062);
xnor U3876 (N_3876,N_3233,N_3049);
xor U3877 (N_3877,N_3387,N_3005);
or U3878 (N_3878,N_3456,N_3468);
and U3879 (N_3879,N_3403,N_3393);
or U3880 (N_3880,N_3310,N_3173);
nor U3881 (N_3881,N_3149,N_3020);
xor U3882 (N_3882,N_3430,N_3177);
xor U3883 (N_3883,N_3054,N_3454);
xor U3884 (N_3884,N_3232,N_3241);
xor U3885 (N_3885,N_3385,N_3274);
nor U3886 (N_3886,N_3242,N_3472);
nor U3887 (N_3887,N_3104,N_3392);
or U3888 (N_3888,N_3124,N_3356);
xor U3889 (N_3889,N_3466,N_3395);
nor U3890 (N_3890,N_3119,N_3044);
nand U3891 (N_3891,N_3286,N_3401);
or U3892 (N_3892,N_3223,N_3101);
and U3893 (N_3893,N_3029,N_3250);
nor U3894 (N_3894,N_3089,N_3317);
or U3895 (N_3895,N_3050,N_3029);
xnor U3896 (N_3896,N_3133,N_3313);
and U3897 (N_3897,N_3276,N_3154);
and U3898 (N_3898,N_3078,N_3105);
xor U3899 (N_3899,N_3236,N_3313);
nor U3900 (N_3900,N_3072,N_3196);
or U3901 (N_3901,N_3131,N_3434);
and U3902 (N_3902,N_3427,N_3300);
nand U3903 (N_3903,N_3425,N_3113);
nand U3904 (N_3904,N_3456,N_3271);
nor U3905 (N_3905,N_3053,N_3381);
nor U3906 (N_3906,N_3482,N_3370);
and U3907 (N_3907,N_3071,N_3062);
xor U3908 (N_3908,N_3152,N_3470);
or U3909 (N_3909,N_3266,N_3318);
or U3910 (N_3910,N_3491,N_3381);
nand U3911 (N_3911,N_3306,N_3169);
nand U3912 (N_3912,N_3335,N_3314);
nand U3913 (N_3913,N_3050,N_3264);
nor U3914 (N_3914,N_3072,N_3484);
nand U3915 (N_3915,N_3236,N_3178);
and U3916 (N_3916,N_3456,N_3019);
xnor U3917 (N_3917,N_3331,N_3263);
or U3918 (N_3918,N_3272,N_3145);
nand U3919 (N_3919,N_3466,N_3231);
nand U3920 (N_3920,N_3328,N_3178);
or U3921 (N_3921,N_3167,N_3332);
nand U3922 (N_3922,N_3247,N_3391);
nand U3923 (N_3923,N_3498,N_3104);
nand U3924 (N_3924,N_3107,N_3030);
nor U3925 (N_3925,N_3007,N_3349);
nand U3926 (N_3926,N_3484,N_3025);
nor U3927 (N_3927,N_3123,N_3198);
nor U3928 (N_3928,N_3309,N_3397);
nand U3929 (N_3929,N_3434,N_3129);
and U3930 (N_3930,N_3497,N_3498);
or U3931 (N_3931,N_3438,N_3214);
xnor U3932 (N_3932,N_3457,N_3198);
or U3933 (N_3933,N_3340,N_3492);
nand U3934 (N_3934,N_3239,N_3001);
nand U3935 (N_3935,N_3446,N_3494);
nand U3936 (N_3936,N_3420,N_3092);
and U3937 (N_3937,N_3302,N_3365);
and U3938 (N_3938,N_3256,N_3098);
nor U3939 (N_3939,N_3047,N_3044);
nand U3940 (N_3940,N_3403,N_3460);
and U3941 (N_3941,N_3345,N_3041);
and U3942 (N_3942,N_3150,N_3399);
nand U3943 (N_3943,N_3362,N_3097);
nor U3944 (N_3944,N_3377,N_3060);
and U3945 (N_3945,N_3024,N_3459);
or U3946 (N_3946,N_3063,N_3386);
or U3947 (N_3947,N_3471,N_3193);
nor U3948 (N_3948,N_3433,N_3464);
and U3949 (N_3949,N_3481,N_3048);
and U3950 (N_3950,N_3160,N_3137);
and U3951 (N_3951,N_3474,N_3273);
or U3952 (N_3952,N_3281,N_3308);
or U3953 (N_3953,N_3323,N_3166);
nand U3954 (N_3954,N_3202,N_3178);
and U3955 (N_3955,N_3260,N_3206);
nand U3956 (N_3956,N_3287,N_3448);
and U3957 (N_3957,N_3170,N_3441);
nand U3958 (N_3958,N_3349,N_3188);
nor U3959 (N_3959,N_3418,N_3419);
nand U3960 (N_3960,N_3179,N_3403);
nor U3961 (N_3961,N_3269,N_3496);
and U3962 (N_3962,N_3092,N_3408);
or U3963 (N_3963,N_3000,N_3220);
and U3964 (N_3964,N_3326,N_3357);
xor U3965 (N_3965,N_3233,N_3171);
nand U3966 (N_3966,N_3008,N_3467);
or U3967 (N_3967,N_3285,N_3485);
or U3968 (N_3968,N_3367,N_3048);
xnor U3969 (N_3969,N_3462,N_3395);
nor U3970 (N_3970,N_3267,N_3446);
nor U3971 (N_3971,N_3029,N_3401);
or U3972 (N_3972,N_3485,N_3096);
nor U3973 (N_3973,N_3426,N_3254);
or U3974 (N_3974,N_3275,N_3005);
nand U3975 (N_3975,N_3031,N_3491);
and U3976 (N_3976,N_3280,N_3442);
or U3977 (N_3977,N_3444,N_3421);
nand U3978 (N_3978,N_3100,N_3161);
nor U3979 (N_3979,N_3122,N_3309);
xnor U3980 (N_3980,N_3390,N_3162);
or U3981 (N_3981,N_3088,N_3382);
nor U3982 (N_3982,N_3212,N_3122);
nor U3983 (N_3983,N_3199,N_3104);
nand U3984 (N_3984,N_3364,N_3077);
xnor U3985 (N_3985,N_3359,N_3248);
xnor U3986 (N_3986,N_3211,N_3102);
nor U3987 (N_3987,N_3048,N_3363);
and U3988 (N_3988,N_3143,N_3410);
or U3989 (N_3989,N_3000,N_3206);
or U3990 (N_3990,N_3430,N_3409);
nand U3991 (N_3991,N_3223,N_3460);
nor U3992 (N_3992,N_3465,N_3029);
and U3993 (N_3993,N_3365,N_3305);
nor U3994 (N_3994,N_3094,N_3178);
or U3995 (N_3995,N_3333,N_3439);
nor U3996 (N_3996,N_3481,N_3038);
and U3997 (N_3997,N_3434,N_3042);
nor U3998 (N_3998,N_3015,N_3219);
nand U3999 (N_3999,N_3417,N_3390);
nor U4000 (N_4000,N_3828,N_3783);
and U4001 (N_4001,N_3734,N_3677);
nand U4002 (N_4002,N_3672,N_3681);
xnor U4003 (N_4003,N_3740,N_3564);
and U4004 (N_4004,N_3501,N_3788);
and U4005 (N_4005,N_3826,N_3764);
xnor U4006 (N_4006,N_3917,N_3526);
nor U4007 (N_4007,N_3996,N_3638);
nor U4008 (N_4008,N_3611,N_3542);
and U4009 (N_4009,N_3876,N_3646);
or U4010 (N_4010,N_3571,N_3918);
nor U4011 (N_4011,N_3811,N_3804);
nand U4012 (N_4012,N_3931,N_3737);
and U4013 (N_4013,N_3796,N_3517);
or U4014 (N_4014,N_3978,N_3742);
and U4015 (N_4015,N_3799,N_3768);
xor U4016 (N_4016,N_3806,N_3547);
nor U4017 (N_4017,N_3756,N_3817);
and U4018 (N_4018,N_3835,N_3892);
nor U4019 (N_4019,N_3823,N_3626);
nor U4020 (N_4020,N_3589,N_3797);
nand U4021 (N_4021,N_3991,N_3697);
or U4022 (N_4022,N_3537,N_3614);
and U4023 (N_4023,N_3849,N_3691);
and U4024 (N_4024,N_3922,N_3718);
nor U4025 (N_4025,N_3843,N_3727);
xor U4026 (N_4026,N_3552,N_3670);
or U4027 (N_4027,N_3512,N_3722);
nor U4028 (N_4028,N_3506,N_3771);
and U4029 (N_4029,N_3902,N_3824);
nand U4030 (N_4030,N_3732,N_3896);
and U4031 (N_4031,N_3781,N_3770);
nand U4032 (N_4032,N_3985,N_3669);
or U4033 (N_4033,N_3898,N_3527);
nor U4034 (N_4034,N_3710,N_3780);
nor U4035 (N_4035,N_3994,N_3642);
or U4036 (N_4036,N_3841,N_3551);
or U4037 (N_4037,N_3704,N_3906);
xor U4038 (N_4038,N_3921,N_3923);
xor U4039 (N_4039,N_3630,N_3977);
xnor U4040 (N_4040,N_3723,N_3757);
and U4041 (N_4041,N_3594,N_3654);
and U4042 (N_4042,N_3827,N_3919);
nor U4043 (N_4043,N_3590,N_3546);
or U4044 (N_4044,N_3945,N_3500);
nor U4045 (N_4045,N_3556,N_3621);
and U4046 (N_4046,N_3949,N_3524);
or U4047 (N_4047,N_3543,N_3709);
nand U4048 (N_4048,N_3576,N_3809);
and U4049 (N_4049,N_3947,N_3731);
or U4050 (N_4050,N_3836,N_3950);
nand U4051 (N_4051,N_3775,N_3636);
and U4052 (N_4052,N_3961,N_3667);
and U4053 (N_4053,N_3511,N_3510);
or U4054 (N_4054,N_3713,N_3563);
nand U4055 (N_4055,N_3599,N_3692);
and U4056 (N_4056,N_3585,N_3608);
and U4057 (N_4057,N_3533,N_3795);
or U4058 (N_4058,N_3728,N_3936);
and U4059 (N_4059,N_3930,N_3908);
or U4060 (N_4060,N_3929,N_3766);
or U4061 (N_4061,N_3530,N_3741);
nand U4062 (N_4062,N_3598,N_3970);
nor U4063 (N_4063,N_3690,N_3749);
and U4064 (N_4064,N_3767,N_3678);
nand U4065 (N_4065,N_3698,N_3820);
xor U4066 (N_4066,N_3875,N_3569);
and U4067 (N_4067,N_3535,N_3658);
or U4068 (N_4068,N_3659,N_3953);
and U4069 (N_4069,N_3759,N_3905);
nand U4070 (N_4070,N_3974,N_3683);
or U4071 (N_4071,N_3565,N_3503);
and U4072 (N_4072,N_3655,N_3647);
nand U4073 (N_4073,N_3976,N_3668);
or U4074 (N_4074,N_3502,N_3584);
or U4075 (N_4075,N_3833,N_3987);
nand U4076 (N_4076,N_3966,N_3831);
xor U4077 (N_4077,N_3889,N_3873);
xor U4078 (N_4078,N_3582,N_3623);
nor U4079 (N_4079,N_3819,N_3591);
nand U4080 (N_4080,N_3975,N_3763);
or U4081 (N_4081,N_3572,N_3720);
nand U4082 (N_4082,N_3782,N_3958);
nand U4083 (N_4083,N_3689,N_3904);
xor U4084 (N_4084,N_3925,N_3665);
nor U4085 (N_4085,N_3748,N_3661);
nand U4086 (N_4086,N_3864,N_3536);
xor U4087 (N_4087,N_3981,N_3913);
and U4088 (N_4088,N_3911,N_3561);
nor U4089 (N_4089,N_3992,N_3562);
or U4090 (N_4090,N_3733,N_3664);
and U4091 (N_4091,N_3635,N_3967);
nand U4092 (N_4092,N_3838,N_3761);
or U4093 (N_4093,N_3529,N_3739);
or U4094 (N_4094,N_3984,N_3867);
or U4095 (N_4095,N_3525,N_3848);
or U4096 (N_4096,N_3729,N_3604);
or U4097 (N_4097,N_3520,N_3968);
nand U4098 (N_4098,N_3586,N_3993);
or U4099 (N_4099,N_3802,N_3825);
or U4100 (N_4100,N_3818,N_3513);
and U4101 (N_4101,N_3699,N_3810);
and U4102 (N_4102,N_3807,N_3721);
or U4103 (N_4103,N_3952,N_3595);
and U4104 (N_4104,N_3883,N_3730);
nor U4105 (N_4105,N_3842,N_3778);
and U4106 (N_4106,N_3587,N_3938);
and U4107 (N_4107,N_3865,N_3888);
nor U4108 (N_4108,N_3592,N_3701);
nor U4109 (N_4109,N_3869,N_3504);
nor U4110 (N_4110,N_3871,N_3762);
nor U4111 (N_4111,N_3909,N_3680);
nor U4112 (N_4112,N_3774,N_3965);
nor U4113 (N_4113,N_3792,N_3924);
xnor U4114 (N_4114,N_3803,N_3726);
nand U4115 (N_4115,N_3695,N_3559);
or U4116 (N_4116,N_3631,N_3858);
xnor U4117 (N_4117,N_3789,N_3753);
nand U4118 (N_4118,N_3518,N_3995);
or U4119 (N_4119,N_3861,N_3575);
nor U4120 (N_4120,N_3893,N_3989);
xor U4121 (N_4121,N_3894,N_3602);
xor U4122 (N_4122,N_3622,N_3581);
xnor U4123 (N_4123,N_3884,N_3983);
xnor U4124 (N_4124,N_3685,N_3760);
and U4125 (N_4125,N_3596,N_3960);
nand U4126 (N_4126,N_3990,N_3580);
or U4127 (N_4127,N_3853,N_3816);
nor U4128 (N_4128,N_3779,N_3866);
nand U4129 (N_4129,N_3752,N_3777);
nand U4130 (N_4130,N_3744,N_3885);
and U4131 (N_4131,N_3850,N_3573);
nand U4132 (N_4132,N_3605,N_3920);
nor U4133 (N_4133,N_3652,N_3639);
nand U4134 (N_4134,N_3675,N_3972);
xnor U4135 (N_4135,N_3508,N_3671);
nand U4136 (N_4136,N_3579,N_3790);
and U4137 (N_4137,N_3891,N_3684);
nand U4138 (N_4138,N_3868,N_3568);
nor U4139 (N_4139,N_3750,N_3969);
or U4140 (N_4140,N_3588,N_3634);
and U4141 (N_4141,N_3886,N_3830);
or U4142 (N_4142,N_3769,N_3619);
nor U4143 (N_4143,N_3736,N_3791);
nand U4144 (N_4144,N_3673,N_3746);
nand U4145 (N_4145,N_3856,N_3532);
or U4146 (N_4146,N_3872,N_3716);
nor U4147 (N_4147,N_3625,N_3932);
or U4148 (N_4148,N_3544,N_3628);
nor U4149 (N_4149,N_3553,N_3583);
nand U4150 (N_4150,N_3808,N_3735);
nand U4151 (N_4151,N_3674,N_3787);
nor U4152 (N_4152,N_3687,N_3812);
nor U4153 (N_4153,N_3815,N_3613);
nand U4154 (N_4154,N_3743,N_3549);
or U4155 (N_4155,N_3890,N_3956);
and U4156 (N_4156,N_3534,N_3711);
nand U4157 (N_4157,N_3900,N_3627);
and U4158 (N_4158,N_3874,N_3988);
and U4159 (N_4159,N_3879,N_3597);
nand U4160 (N_4160,N_3877,N_3725);
nor U4161 (N_4161,N_3959,N_3612);
nor U4162 (N_4162,N_3521,N_3644);
nand U4163 (N_4163,N_3682,N_3948);
or U4164 (N_4164,N_3963,N_3832);
or U4165 (N_4165,N_3852,N_3857);
nand U4166 (N_4166,N_3629,N_3577);
nand U4167 (N_4167,N_3914,N_3954);
xnor U4168 (N_4168,N_3708,N_3751);
nor U4169 (N_4169,N_3528,N_3717);
or U4170 (N_4170,N_3982,N_3705);
and U4171 (N_4171,N_3863,N_3845);
and U4172 (N_4172,N_3951,N_3615);
or U4173 (N_4173,N_3666,N_3662);
or U4174 (N_4174,N_3793,N_3773);
and U4175 (N_4175,N_3765,N_3632);
nand U4176 (N_4176,N_3798,N_3657);
nand U4177 (N_4177,N_3946,N_3957);
nand U4178 (N_4178,N_3523,N_3860);
or U4179 (N_4179,N_3979,N_3916);
or U4180 (N_4180,N_3747,N_3901);
or U4181 (N_4181,N_3618,N_3620);
and U4182 (N_4182,N_3944,N_3641);
xnor U4183 (N_4183,N_3560,N_3882);
or U4184 (N_4184,N_3505,N_3998);
xnor U4185 (N_4185,N_3617,N_3880);
and U4186 (N_4186,N_3707,N_3897);
nand U4187 (N_4187,N_3928,N_3509);
and U4188 (N_4188,N_3813,N_3964);
nand U4189 (N_4189,N_3507,N_3606);
nor U4190 (N_4190,N_3715,N_3558);
xnor U4191 (N_4191,N_3800,N_3514);
or U4192 (N_4192,N_3962,N_3786);
or U4193 (N_4193,N_3999,N_3609);
xor U4194 (N_4194,N_3714,N_3702);
or U4195 (N_4195,N_3941,N_3519);
and U4196 (N_4196,N_3854,N_3834);
nand U4197 (N_4197,N_3821,N_3942);
nor U4198 (N_4198,N_3794,N_3859);
nor U4199 (N_4199,N_3570,N_3785);
nor U4200 (N_4200,N_3550,N_3676);
nor U4201 (N_4201,N_3937,N_3940);
or U4202 (N_4202,N_3939,N_3567);
nand U4203 (N_4203,N_3700,N_3578);
xor U4204 (N_4204,N_3738,N_3943);
and U4205 (N_4205,N_3693,N_3927);
or U4206 (N_4206,N_3837,N_3540);
and U4207 (N_4207,N_3607,N_3610);
and U4208 (N_4208,N_3633,N_3600);
and U4209 (N_4209,N_3755,N_3541);
nand U4210 (N_4210,N_3719,N_3538);
nor U4211 (N_4211,N_3648,N_3555);
or U4212 (N_4212,N_3887,N_3706);
xnor U4213 (N_4213,N_3851,N_3980);
or U4214 (N_4214,N_3829,N_3955);
and U4215 (N_4215,N_3688,N_3912);
xnor U4216 (N_4216,N_3839,N_3784);
or U4217 (N_4217,N_3566,N_3651);
or U4218 (N_4218,N_3515,N_3881);
nor U4219 (N_4219,N_3653,N_3840);
and U4220 (N_4220,N_3640,N_3724);
and U4221 (N_4221,N_3637,N_3557);
nor U4222 (N_4222,N_3663,N_3776);
nor U4223 (N_4223,N_3971,N_3997);
nor U4224 (N_4224,N_3574,N_3686);
or U4225 (N_4225,N_3973,N_3603);
or U4226 (N_4226,N_3660,N_3645);
or U4227 (N_4227,N_3545,N_3933);
or U4228 (N_4228,N_3754,N_3516);
or U4229 (N_4229,N_3758,N_3593);
nor U4230 (N_4230,N_3903,N_3844);
or U4231 (N_4231,N_3649,N_3935);
nand U4232 (N_4232,N_3696,N_3772);
and U4233 (N_4233,N_3855,N_3814);
and U4234 (N_4234,N_3679,N_3650);
nand U4235 (N_4235,N_3862,N_3895);
or U4236 (N_4236,N_3539,N_3616);
nor U4237 (N_4237,N_3643,N_3624);
or U4238 (N_4238,N_3531,N_3548);
nand U4239 (N_4239,N_3745,N_3907);
or U4240 (N_4240,N_3801,N_3712);
and U4241 (N_4241,N_3601,N_3899);
and U4242 (N_4242,N_3822,N_3910);
and U4243 (N_4243,N_3656,N_3934);
or U4244 (N_4244,N_3703,N_3847);
nand U4245 (N_4245,N_3694,N_3870);
or U4246 (N_4246,N_3846,N_3926);
nor U4247 (N_4247,N_3878,N_3915);
and U4248 (N_4248,N_3554,N_3805);
nor U4249 (N_4249,N_3522,N_3986);
nand U4250 (N_4250,N_3589,N_3710);
nand U4251 (N_4251,N_3868,N_3620);
and U4252 (N_4252,N_3667,N_3744);
nor U4253 (N_4253,N_3977,N_3768);
nand U4254 (N_4254,N_3678,N_3527);
or U4255 (N_4255,N_3840,N_3549);
and U4256 (N_4256,N_3945,N_3709);
nand U4257 (N_4257,N_3898,N_3605);
xor U4258 (N_4258,N_3812,N_3633);
xor U4259 (N_4259,N_3979,N_3776);
or U4260 (N_4260,N_3685,N_3563);
nor U4261 (N_4261,N_3780,N_3636);
nand U4262 (N_4262,N_3771,N_3572);
or U4263 (N_4263,N_3568,N_3991);
nand U4264 (N_4264,N_3647,N_3866);
nor U4265 (N_4265,N_3828,N_3606);
and U4266 (N_4266,N_3914,N_3649);
or U4267 (N_4267,N_3918,N_3512);
or U4268 (N_4268,N_3519,N_3722);
nor U4269 (N_4269,N_3536,N_3626);
or U4270 (N_4270,N_3587,N_3721);
and U4271 (N_4271,N_3849,N_3684);
nand U4272 (N_4272,N_3823,N_3830);
xor U4273 (N_4273,N_3888,N_3856);
or U4274 (N_4274,N_3873,N_3559);
nand U4275 (N_4275,N_3731,N_3592);
or U4276 (N_4276,N_3591,N_3930);
nor U4277 (N_4277,N_3808,N_3757);
or U4278 (N_4278,N_3577,N_3920);
and U4279 (N_4279,N_3518,N_3773);
and U4280 (N_4280,N_3948,N_3746);
nand U4281 (N_4281,N_3674,N_3690);
and U4282 (N_4282,N_3853,N_3985);
and U4283 (N_4283,N_3877,N_3569);
xnor U4284 (N_4284,N_3892,N_3675);
nand U4285 (N_4285,N_3553,N_3754);
and U4286 (N_4286,N_3509,N_3768);
and U4287 (N_4287,N_3653,N_3574);
and U4288 (N_4288,N_3767,N_3505);
and U4289 (N_4289,N_3666,N_3704);
and U4290 (N_4290,N_3989,N_3980);
nand U4291 (N_4291,N_3772,N_3508);
nand U4292 (N_4292,N_3984,N_3868);
nand U4293 (N_4293,N_3632,N_3644);
nand U4294 (N_4294,N_3931,N_3791);
and U4295 (N_4295,N_3941,N_3654);
and U4296 (N_4296,N_3895,N_3620);
and U4297 (N_4297,N_3609,N_3621);
nor U4298 (N_4298,N_3618,N_3694);
or U4299 (N_4299,N_3811,N_3583);
nand U4300 (N_4300,N_3966,N_3624);
and U4301 (N_4301,N_3943,N_3676);
nor U4302 (N_4302,N_3820,N_3861);
xnor U4303 (N_4303,N_3708,N_3773);
or U4304 (N_4304,N_3914,N_3908);
and U4305 (N_4305,N_3687,N_3887);
or U4306 (N_4306,N_3905,N_3684);
or U4307 (N_4307,N_3621,N_3978);
xor U4308 (N_4308,N_3506,N_3731);
nor U4309 (N_4309,N_3852,N_3584);
nand U4310 (N_4310,N_3776,N_3791);
nand U4311 (N_4311,N_3744,N_3752);
xor U4312 (N_4312,N_3746,N_3770);
nor U4313 (N_4313,N_3851,N_3691);
nor U4314 (N_4314,N_3987,N_3892);
nand U4315 (N_4315,N_3898,N_3787);
and U4316 (N_4316,N_3707,N_3697);
and U4317 (N_4317,N_3608,N_3978);
or U4318 (N_4318,N_3592,N_3642);
nor U4319 (N_4319,N_3931,N_3657);
and U4320 (N_4320,N_3844,N_3875);
or U4321 (N_4321,N_3766,N_3932);
and U4322 (N_4322,N_3844,N_3929);
nand U4323 (N_4323,N_3709,N_3718);
xnor U4324 (N_4324,N_3629,N_3856);
and U4325 (N_4325,N_3824,N_3611);
nand U4326 (N_4326,N_3565,N_3961);
nor U4327 (N_4327,N_3815,N_3504);
nand U4328 (N_4328,N_3759,N_3951);
nand U4329 (N_4329,N_3963,N_3606);
or U4330 (N_4330,N_3559,N_3518);
and U4331 (N_4331,N_3719,N_3984);
nor U4332 (N_4332,N_3737,N_3525);
or U4333 (N_4333,N_3534,N_3755);
nor U4334 (N_4334,N_3739,N_3956);
and U4335 (N_4335,N_3518,N_3706);
nor U4336 (N_4336,N_3547,N_3914);
nand U4337 (N_4337,N_3889,N_3691);
nand U4338 (N_4338,N_3638,N_3693);
nand U4339 (N_4339,N_3806,N_3803);
or U4340 (N_4340,N_3612,N_3627);
nor U4341 (N_4341,N_3549,N_3531);
or U4342 (N_4342,N_3555,N_3993);
and U4343 (N_4343,N_3810,N_3706);
nor U4344 (N_4344,N_3523,N_3645);
nor U4345 (N_4345,N_3653,N_3945);
nor U4346 (N_4346,N_3585,N_3955);
or U4347 (N_4347,N_3748,N_3745);
nand U4348 (N_4348,N_3627,N_3886);
xnor U4349 (N_4349,N_3993,N_3969);
and U4350 (N_4350,N_3703,N_3951);
nor U4351 (N_4351,N_3500,N_3663);
or U4352 (N_4352,N_3882,N_3676);
and U4353 (N_4353,N_3613,N_3712);
or U4354 (N_4354,N_3980,N_3587);
and U4355 (N_4355,N_3991,N_3593);
and U4356 (N_4356,N_3820,N_3648);
or U4357 (N_4357,N_3554,N_3765);
or U4358 (N_4358,N_3596,N_3836);
or U4359 (N_4359,N_3775,N_3784);
and U4360 (N_4360,N_3617,N_3635);
and U4361 (N_4361,N_3751,N_3616);
nor U4362 (N_4362,N_3646,N_3913);
or U4363 (N_4363,N_3729,N_3757);
nor U4364 (N_4364,N_3863,N_3968);
and U4365 (N_4365,N_3592,N_3804);
nor U4366 (N_4366,N_3869,N_3587);
or U4367 (N_4367,N_3866,N_3530);
and U4368 (N_4368,N_3789,N_3691);
xnor U4369 (N_4369,N_3714,N_3579);
and U4370 (N_4370,N_3858,N_3539);
nor U4371 (N_4371,N_3670,N_3744);
and U4372 (N_4372,N_3944,N_3578);
nand U4373 (N_4373,N_3957,N_3560);
nand U4374 (N_4374,N_3566,N_3718);
nand U4375 (N_4375,N_3832,N_3572);
nor U4376 (N_4376,N_3931,N_3835);
or U4377 (N_4377,N_3774,N_3693);
or U4378 (N_4378,N_3760,N_3848);
nor U4379 (N_4379,N_3559,N_3685);
xor U4380 (N_4380,N_3682,N_3890);
xor U4381 (N_4381,N_3904,N_3741);
nand U4382 (N_4382,N_3869,N_3506);
xnor U4383 (N_4383,N_3657,N_3945);
nor U4384 (N_4384,N_3691,N_3861);
xnor U4385 (N_4385,N_3893,N_3605);
or U4386 (N_4386,N_3759,N_3947);
or U4387 (N_4387,N_3673,N_3505);
nor U4388 (N_4388,N_3975,N_3921);
and U4389 (N_4389,N_3820,N_3624);
or U4390 (N_4390,N_3903,N_3949);
and U4391 (N_4391,N_3756,N_3623);
or U4392 (N_4392,N_3962,N_3872);
nor U4393 (N_4393,N_3695,N_3850);
and U4394 (N_4394,N_3945,N_3887);
and U4395 (N_4395,N_3841,N_3595);
or U4396 (N_4396,N_3843,N_3697);
nand U4397 (N_4397,N_3939,N_3762);
and U4398 (N_4398,N_3963,N_3917);
and U4399 (N_4399,N_3737,N_3576);
nor U4400 (N_4400,N_3552,N_3677);
or U4401 (N_4401,N_3965,N_3791);
nor U4402 (N_4402,N_3770,N_3572);
nand U4403 (N_4403,N_3913,N_3797);
nor U4404 (N_4404,N_3782,N_3677);
or U4405 (N_4405,N_3720,N_3662);
and U4406 (N_4406,N_3578,N_3697);
and U4407 (N_4407,N_3970,N_3872);
nor U4408 (N_4408,N_3651,N_3867);
or U4409 (N_4409,N_3980,N_3962);
or U4410 (N_4410,N_3785,N_3546);
and U4411 (N_4411,N_3627,N_3608);
nand U4412 (N_4412,N_3987,N_3672);
or U4413 (N_4413,N_3530,N_3509);
xor U4414 (N_4414,N_3850,N_3578);
or U4415 (N_4415,N_3615,N_3779);
nand U4416 (N_4416,N_3891,N_3700);
and U4417 (N_4417,N_3540,N_3795);
nand U4418 (N_4418,N_3579,N_3822);
nand U4419 (N_4419,N_3546,N_3569);
xnor U4420 (N_4420,N_3875,N_3639);
xor U4421 (N_4421,N_3559,N_3669);
nor U4422 (N_4422,N_3683,N_3656);
or U4423 (N_4423,N_3860,N_3868);
nand U4424 (N_4424,N_3959,N_3955);
nand U4425 (N_4425,N_3934,N_3501);
nand U4426 (N_4426,N_3824,N_3516);
nor U4427 (N_4427,N_3522,N_3560);
xnor U4428 (N_4428,N_3895,N_3795);
and U4429 (N_4429,N_3583,N_3693);
nand U4430 (N_4430,N_3938,N_3751);
nor U4431 (N_4431,N_3811,N_3810);
xnor U4432 (N_4432,N_3895,N_3586);
and U4433 (N_4433,N_3821,N_3505);
or U4434 (N_4434,N_3533,N_3920);
nand U4435 (N_4435,N_3582,N_3727);
or U4436 (N_4436,N_3831,N_3541);
nor U4437 (N_4437,N_3935,N_3924);
nand U4438 (N_4438,N_3627,N_3567);
xnor U4439 (N_4439,N_3942,N_3780);
nor U4440 (N_4440,N_3741,N_3764);
nand U4441 (N_4441,N_3910,N_3700);
nor U4442 (N_4442,N_3897,N_3906);
or U4443 (N_4443,N_3816,N_3951);
nand U4444 (N_4444,N_3752,N_3612);
xnor U4445 (N_4445,N_3783,N_3670);
and U4446 (N_4446,N_3789,N_3875);
xor U4447 (N_4447,N_3510,N_3611);
nand U4448 (N_4448,N_3682,N_3543);
or U4449 (N_4449,N_3541,N_3543);
nand U4450 (N_4450,N_3784,N_3849);
or U4451 (N_4451,N_3706,N_3984);
or U4452 (N_4452,N_3544,N_3772);
and U4453 (N_4453,N_3934,N_3546);
or U4454 (N_4454,N_3596,N_3639);
xnor U4455 (N_4455,N_3983,N_3766);
nor U4456 (N_4456,N_3782,N_3865);
nor U4457 (N_4457,N_3540,N_3549);
nor U4458 (N_4458,N_3634,N_3556);
or U4459 (N_4459,N_3920,N_3679);
nand U4460 (N_4460,N_3715,N_3501);
nand U4461 (N_4461,N_3613,N_3917);
or U4462 (N_4462,N_3524,N_3772);
nand U4463 (N_4463,N_3602,N_3997);
nand U4464 (N_4464,N_3547,N_3598);
nand U4465 (N_4465,N_3861,N_3636);
nor U4466 (N_4466,N_3945,N_3883);
nand U4467 (N_4467,N_3787,N_3758);
or U4468 (N_4468,N_3748,N_3543);
nor U4469 (N_4469,N_3803,N_3935);
and U4470 (N_4470,N_3901,N_3983);
nand U4471 (N_4471,N_3972,N_3772);
nand U4472 (N_4472,N_3856,N_3674);
nand U4473 (N_4473,N_3917,N_3525);
or U4474 (N_4474,N_3745,N_3674);
xnor U4475 (N_4475,N_3776,N_3533);
nor U4476 (N_4476,N_3911,N_3889);
or U4477 (N_4477,N_3814,N_3771);
nor U4478 (N_4478,N_3581,N_3959);
nand U4479 (N_4479,N_3808,N_3785);
and U4480 (N_4480,N_3698,N_3679);
nor U4481 (N_4481,N_3738,N_3511);
nand U4482 (N_4482,N_3952,N_3546);
xnor U4483 (N_4483,N_3565,N_3513);
nand U4484 (N_4484,N_3520,N_3717);
xnor U4485 (N_4485,N_3647,N_3649);
xnor U4486 (N_4486,N_3623,N_3569);
nor U4487 (N_4487,N_3946,N_3886);
nand U4488 (N_4488,N_3636,N_3541);
or U4489 (N_4489,N_3796,N_3861);
nor U4490 (N_4490,N_3743,N_3789);
or U4491 (N_4491,N_3632,N_3718);
and U4492 (N_4492,N_3969,N_3559);
and U4493 (N_4493,N_3801,N_3909);
or U4494 (N_4494,N_3871,N_3587);
or U4495 (N_4495,N_3601,N_3992);
and U4496 (N_4496,N_3543,N_3959);
and U4497 (N_4497,N_3871,N_3568);
nor U4498 (N_4498,N_3581,N_3615);
nor U4499 (N_4499,N_3728,N_3536);
nor U4500 (N_4500,N_4391,N_4454);
and U4501 (N_4501,N_4459,N_4435);
nor U4502 (N_4502,N_4000,N_4255);
nor U4503 (N_4503,N_4293,N_4025);
nor U4504 (N_4504,N_4195,N_4415);
and U4505 (N_4505,N_4225,N_4235);
nand U4506 (N_4506,N_4183,N_4281);
nand U4507 (N_4507,N_4018,N_4278);
or U4508 (N_4508,N_4353,N_4011);
and U4509 (N_4509,N_4053,N_4298);
nor U4510 (N_4510,N_4354,N_4147);
or U4511 (N_4511,N_4497,N_4153);
nand U4512 (N_4512,N_4388,N_4165);
nand U4513 (N_4513,N_4070,N_4347);
xnor U4514 (N_4514,N_4456,N_4177);
nor U4515 (N_4515,N_4112,N_4125);
nor U4516 (N_4516,N_4083,N_4409);
nor U4517 (N_4517,N_4472,N_4422);
and U4518 (N_4518,N_4020,N_4023);
nor U4519 (N_4519,N_4038,N_4363);
nand U4520 (N_4520,N_4292,N_4368);
and U4521 (N_4521,N_4243,N_4010);
or U4522 (N_4522,N_4002,N_4107);
nand U4523 (N_4523,N_4431,N_4279);
and U4524 (N_4524,N_4437,N_4263);
and U4525 (N_4525,N_4051,N_4009);
and U4526 (N_4526,N_4175,N_4467);
or U4527 (N_4527,N_4260,N_4270);
and U4528 (N_4528,N_4049,N_4072);
nor U4529 (N_4529,N_4275,N_4021);
nand U4530 (N_4530,N_4158,N_4259);
nand U4531 (N_4531,N_4283,N_4077);
or U4532 (N_4532,N_4372,N_4062);
and U4533 (N_4533,N_4233,N_4328);
xnor U4534 (N_4534,N_4035,N_4358);
nand U4535 (N_4535,N_4184,N_4173);
xor U4536 (N_4536,N_4093,N_4345);
or U4537 (N_4537,N_4485,N_4374);
nor U4538 (N_4538,N_4461,N_4264);
and U4539 (N_4539,N_4357,N_4138);
or U4540 (N_4540,N_4236,N_4284);
xnor U4541 (N_4541,N_4491,N_4222);
nand U4542 (N_4542,N_4385,N_4065);
and U4543 (N_4543,N_4288,N_4311);
xnor U4544 (N_4544,N_4280,N_4108);
nand U4545 (N_4545,N_4064,N_4069);
or U4546 (N_4546,N_4470,N_4132);
nor U4547 (N_4547,N_4364,N_4131);
xnor U4548 (N_4548,N_4355,N_4429);
and U4549 (N_4549,N_4192,N_4239);
or U4550 (N_4550,N_4398,N_4223);
nand U4551 (N_4551,N_4334,N_4127);
and U4552 (N_4552,N_4428,N_4095);
or U4553 (N_4553,N_4446,N_4081);
or U4554 (N_4554,N_4155,N_4277);
nor U4555 (N_4555,N_4430,N_4014);
nor U4556 (N_4556,N_4333,N_4336);
and U4557 (N_4557,N_4142,N_4169);
nor U4558 (N_4558,N_4352,N_4375);
nor U4559 (N_4559,N_4031,N_4097);
nand U4560 (N_4560,N_4059,N_4439);
and U4561 (N_4561,N_4008,N_4122);
nand U4562 (N_4562,N_4346,N_4453);
nor U4563 (N_4563,N_4249,N_4143);
nand U4564 (N_4564,N_4228,N_4204);
xor U4565 (N_4565,N_4359,N_4360);
nor U4566 (N_4566,N_4421,N_4396);
and U4567 (N_4567,N_4427,N_4057);
nor U4568 (N_4568,N_4041,N_4489);
xor U4569 (N_4569,N_4113,N_4494);
and U4570 (N_4570,N_4162,N_4212);
and U4571 (N_4571,N_4136,N_4022);
and U4572 (N_4572,N_4180,N_4244);
or U4573 (N_4573,N_4389,N_4268);
nor U4574 (N_4574,N_4488,N_4118);
nor U4575 (N_4575,N_4078,N_4101);
nor U4576 (N_4576,N_4012,N_4106);
xnor U4577 (N_4577,N_4300,N_4337);
or U4578 (N_4578,N_4201,N_4480);
and U4579 (N_4579,N_4105,N_4048);
nand U4580 (N_4580,N_4499,N_4493);
nor U4581 (N_4581,N_4369,N_4438);
xor U4582 (N_4582,N_4272,N_4432);
nand U4583 (N_4583,N_4013,N_4402);
and U4584 (N_4584,N_4301,N_4046);
nand U4585 (N_4585,N_4080,N_4076);
or U4586 (N_4586,N_4412,N_4130);
and U4587 (N_4587,N_4102,N_4075);
or U4588 (N_4588,N_4410,N_4335);
nor U4589 (N_4589,N_4295,N_4256);
nand U4590 (N_4590,N_4026,N_4045);
nor U4591 (N_4591,N_4447,N_4315);
and U4592 (N_4592,N_4322,N_4308);
nor U4593 (N_4593,N_4492,N_4043);
and U4594 (N_4594,N_4110,N_4167);
or U4595 (N_4595,N_4171,N_4006);
nor U4596 (N_4596,N_4242,N_4227);
nor U4597 (N_4597,N_4193,N_4210);
nand U4598 (N_4598,N_4400,N_4157);
and U4599 (N_4599,N_4119,N_4176);
nand U4600 (N_4600,N_4473,N_4405);
or U4601 (N_4601,N_4111,N_4339);
nand U4602 (N_4602,N_4163,N_4302);
or U4603 (N_4603,N_4403,N_4366);
and U4604 (N_4604,N_4063,N_4338);
nand U4605 (N_4605,N_4139,N_4181);
or U4606 (N_4606,N_4191,N_4028);
or U4607 (N_4607,N_4395,N_4310);
nand U4608 (N_4608,N_4269,N_4015);
and U4609 (N_4609,N_4170,N_4325);
and U4610 (N_4610,N_4090,N_4220);
or U4611 (N_4611,N_4361,N_4319);
and U4612 (N_4612,N_4141,N_4408);
or U4613 (N_4613,N_4234,N_4073);
xor U4614 (N_4614,N_4285,N_4017);
and U4615 (N_4615,N_4323,N_4484);
xnor U4616 (N_4616,N_4426,N_4384);
nor U4617 (N_4617,N_4406,N_4103);
nor U4618 (N_4618,N_4331,N_4237);
nand U4619 (N_4619,N_4367,N_4215);
nor U4620 (N_4620,N_4370,N_4133);
nor U4621 (N_4621,N_4379,N_4450);
nand U4622 (N_4622,N_4267,N_4055);
xnor U4623 (N_4623,N_4282,N_4413);
and U4624 (N_4624,N_4146,N_4085);
and U4625 (N_4625,N_4007,N_4265);
nor U4626 (N_4626,N_4382,N_4109);
and U4627 (N_4627,N_4312,N_4207);
xnor U4628 (N_4628,N_4092,N_4126);
nor U4629 (N_4629,N_4340,N_4034);
nand U4630 (N_4630,N_4116,N_4448);
xor U4631 (N_4631,N_4154,N_4187);
or U4632 (N_4632,N_4185,N_4213);
nand U4633 (N_4633,N_4251,N_4399);
and U4634 (N_4634,N_4123,N_4471);
nand U4635 (N_4635,N_4198,N_4460);
or U4636 (N_4636,N_4469,N_4036);
or U4637 (N_4637,N_4378,N_4387);
nand U4638 (N_4638,N_4208,N_4327);
and U4639 (N_4639,N_4232,N_4054);
or U4640 (N_4640,N_4241,N_4124);
nor U4641 (N_4641,N_4307,N_4253);
xnor U4642 (N_4642,N_4100,N_4117);
xnor U4643 (N_4643,N_4197,N_4150);
nor U4644 (N_4644,N_4386,N_4087);
or U4645 (N_4645,N_4047,N_4052);
and U4646 (N_4646,N_4417,N_4152);
nor U4647 (N_4647,N_4481,N_4455);
nor U4648 (N_4648,N_4343,N_4029);
and U4649 (N_4649,N_4380,N_4060);
nor U4650 (N_4650,N_4088,N_4356);
and U4651 (N_4651,N_4351,N_4238);
nand U4652 (N_4652,N_4320,N_4149);
and U4653 (N_4653,N_4250,N_4140);
nor U4654 (N_4654,N_4121,N_4317);
or U4655 (N_4655,N_4324,N_4290);
nor U4656 (N_4656,N_4129,N_4254);
xnor U4657 (N_4657,N_4420,N_4252);
and U4658 (N_4658,N_4287,N_4321);
and U4659 (N_4659,N_4144,N_4445);
nand U4660 (N_4660,N_4424,N_4273);
nand U4661 (N_4661,N_4094,N_4159);
or U4662 (N_4662,N_4019,N_4341);
and U4663 (N_4663,N_4423,N_4457);
and U4664 (N_4664,N_4286,N_4404);
nor U4665 (N_4665,N_4037,N_4271);
or U4666 (N_4666,N_4482,N_4003);
nor U4667 (N_4667,N_4084,N_4004);
or U4668 (N_4668,N_4443,N_4082);
nor U4669 (N_4669,N_4071,N_4458);
xnor U4670 (N_4670,N_4137,N_4276);
and U4671 (N_4671,N_4394,N_4425);
or U4672 (N_4672,N_4040,N_4050);
nand U4673 (N_4673,N_4135,N_4313);
nor U4674 (N_4674,N_4316,N_4161);
nor U4675 (N_4675,N_4291,N_4202);
nand U4676 (N_4676,N_4058,N_4468);
nand U4677 (N_4677,N_4079,N_4479);
nor U4678 (N_4678,N_4168,N_4487);
or U4679 (N_4679,N_4115,N_4477);
nor U4680 (N_4680,N_4464,N_4309);
xnor U4681 (N_4681,N_4416,N_4200);
and U4682 (N_4682,N_4490,N_4483);
and U4683 (N_4683,N_4433,N_4156);
nand U4684 (N_4684,N_4414,N_4027);
or U4685 (N_4685,N_4257,N_4104);
and U4686 (N_4686,N_4318,N_4475);
nand U4687 (N_4687,N_4373,N_4218);
xor U4688 (N_4688,N_4371,N_4274);
nor U4689 (N_4689,N_4326,N_4074);
and U4690 (N_4690,N_4362,N_4206);
nand U4691 (N_4691,N_4348,N_4294);
nand U4692 (N_4692,N_4042,N_4005);
or U4693 (N_4693,N_4033,N_4392);
and U4694 (N_4694,N_4498,N_4306);
nor U4695 (N_4695,N_4381,N_4436);
nand U4696 (N_4696,N_4296,N_4486);
and U4697 (N_4697,N_4216,N_4332);
and U4698 (N_4698,N_4217,N_4190);
and U4699 (N_4699,N_4226,N_4466);
or U4700 (N_4700,N_4066,N_4452);
or U4701 (N_4701,N_4462,N_4016);
and U4702 (N_4702,N_4496,N_4314);
xnor U4703 (N_4703,N_4160,N_4032);
and U4704 (N_4704,N_4248,N_4258);
nand U4705 (N_4705,N_4240,N_4148);
or U4706 (N_4706,N_4196,N_4478);
or U4707 (N_4707,N_4390,N_4451);
and U4708 (N_4708,N_4262,N_4344);
and U4709 (N_4709,N_4182,N_4189);
and U4710 (N_4710,N_4221,N_4303);
nor U4711 (N_4711,N_4444,N_4030);
or U4712 (N_4712,N_4068,N_4178);
xnor U4713 (N_4713,N_4179,N_4230);
nand U4714 (N_4714,N_4349,N_4186);
and U4715 (N_4715,N_4474,N_4297);
or U4716 (N_4716,N_4120,N_4067);
nand U4717 (N_4717,N_4442,N_4099);
nor U4718 (N_4718,N_4305,N_4098);
or U4719 (N_4719,N_4194,N_4266);
nand U4720 (N_4720,N_4350,N_4393);
or U4721 (N_4721,N_4245,N_4205);
nor U4722 (N_4722,N_4397,N_4114);
nor U4723 (N_4723,N_4039,N_4199);
or U4724 (N_4724,N_4418,N_4128);
or U4725 (N_4725,N_4495,N_4329);
xnor U4726 (N_4726,N_4091,N_4134);
nand U4727 (N_4727,N_4229,N_4164);
xnor U4728 (N_4728,N_4289,N_4024);
and U4729 (N_4729,N_4304,N_4465);
nand U4730 (N_4730,N_4166,N_4401);
or U4731 (N_4731,N_4231,N_4203);
nand U4732 (N_4732,N_4440,N_4434);
nor U4733 (N_4733,N_4441,N_4089);
and U4734 (N_4734,N_4342,N_4172);
nor U4735 (N_4735,N_4419,N_4330);
nand U4736 (N_4736,N_4463,N_4056);
or U4737 (N_4737,N_4247,N_4145);
or U4738 (N_4738,N_4151,N_4061);
or U4739 (N_4739,N_4044,N_4449);
nand U4740 (N_4740,N_4188,N_4299);
or U4741 (N_4741,N_4211,N_4407);
nand U4742 (N_4742,N_4383,N_4411);
or U4743 (N_4743,N_4365,N_4174);
nand U4744 (N_4744,N_4261,N_4224);
nand U4745 (N_4745,N_4214,N_4376);
and U4746 (N_4746,N_4476,N_4086);
or U4747 (N_4747,N_4096,N_4246);
and U4748 (N_4748,N_4377,N_4209);
xnor U4749 (N_4749,N_4001,N_4219);
xor U4750 (N_4750,N_4427,N_4486);
xnor U4751 (N_4751,N_4478,N_4366);
nand U4752 (N_4752,N_4094,N_4082);
nor U4753 (N_4753,N_4269,N_4282);
xnor U4754 (N_4754,N_4062,N_4148);
and U4755 (N_4755,N_4275,N_4262);
xor U4756 (N_4756,N_4457,N_4402);
nor U4757 (N_4757,N_4208,N_4464);
and U4758 (N_4758,N_4045,N_4308);
or U4759 (N_4759,N_4368,N_4331);
nand U4760 (N_4760,N_4367,N_4381);
nor U4761 (N_4761,N_4426,N_4153);
nor U4762 (N_4762,N_4187,N_4103);
and U4763 (N_4763,N_4187,N_4362);
or U4764 (N_4764,N_4067,N_4361);
nand U4765 (N_4765,N_4313,N_4382);
or U4766 (N_4766,N_4421,N_4187);
xor U4767 (N_4767,N_4462,N_4434);
or U4768 (N_4768,N_4098,N_4309);
or U4769 (N_4769,N_4341,N_4069);
and U4770 (N_4770,N_4370,N_4181);
or U4771 (N_4771,N_4307,N_4244);
nor U4772 (N_4772,N_4096,N_4110);
nand U4773 (N_4773,N_4335,N_4237);
nand U4774 (N_4774,N_4320,N_4451);
xor U4775 (N_4775,N_4176,N_4257);
nand U4776 (N_4776,N_4285,N_4235);
nor U4777 (N_4777,N_4303,N_4116);
or U4778 (N_4778,N_4338,N_4314);
and U4779 (N_4779,N_4116,N_4178);
or U4780 (N_4780,N_4029,N_4106);
or U4781 (N_4781,N_4416,N_4122);
or U4782 (N_4782,N_4006,N_4498);
nor U4783 (N_4783,N_4405,N_4417);
nand U4784 (N_4784,N_4319,N_4216);
or U4785 (N_4785,N_4017,N_4037);
nor U4786 (N_4786,N_4496,N_4435);
or U4787 (N_4787,N_4169,N_4403);
nor U4788 (N_4788,N_4310,N_4197);
and U4789 (N_4789,N_4204,N_4148);
nor U4790 (N_4790,N_4421,N_4308);
nor U4791 (N_4791,N_4131,N_4415);
and U4792 (N_4792,N_4152,N_4436);
nand U4793 (N_4793,N_4239,N_4155);
or U4794 (N_4794,N_4449,N_4410);
and U4795 (N_4795,N_4263,N_4405);
nand U4796 (N_4796,N_4015,N_4318);
or U4797 (N_4797,N_4386,N_4296);
nand U4798 (N_4798,N_4228,N_4448);
nand U4799 (N_4799,N_4357,N_4402);
nor U4800 (N_4800,N_4223,N_4222);
xor U4801 (N_4801,N_4116,N_4175);
xnor U4802 (N_4802,N_4464,N_4215);
xnor U4803 (N_4803,N_4104,N_4368);
and U4804 (N_4804,N_4348,N_4459);
and U4805 (N_4805,N_4267,N_4014);
nor U4806 (N_4806,N_4437,N_4498);
and U4807 (N_4807,N_4141,N_4039);
nor U4808 (N_4808,N_4271,N_4320);
nand U4809 (N_4809,N_4449,N_4266);
nand U4810 (N_4810,N_4110,N_4177);
nand U4811 (N_4811,N_4163,N_4020);
or U4812 (N_4812,N_4229,N_4260);
nand U4813 (N_4813,N_4078,N_4478);
nor U4814 (N_4814,N_4179,N_4142);
or U4815 (N_4815,N_4195,N_4291);
nand U4816 (N_4816,N_4383,N_4184);
or U4817 (N_4817,N_4083,N_4369);
nor U4818 (N_4818,N_4273,N_4122);
nand U4819 (N_4819,N_4217,N_4345);
nand U4820 (N_4820,N_4392,N_4183);
nor U4821 (N_4821,N_4005,N_4011);
and U4822 (N_4822,N_4095,N_4016);
and U4823 (N_4823,N_4080,N_4396);
nand U4824 (N_4824,N_4275,N_4437);
xor U4825 (N_4825,N_4266,N_4484);
and U4826 (N_4826,N_4389,N_4109);
and U4827 (N_4827,N_4462,N_4195);
or U4828 (N_4828,N_4435,N_4335);
and U4829 (N_4829,N_4346,N_4426);
nand U4830 (N_4830,N_4405,N_4233);
xor U4831 (N_4831,N_4261,N_4383);
nor U4832 (N_4832,N_4333,N_4391);
nor U4833 (N_4833,N_4417,N_4381);
and U4834 (N_4834,N_4434,N_4244);
nor U4835 (N_4835,N_4186,N_4423);
nor U4836 (N_4836,N_4254,N_4030);
or U4837 (N_4837,N_4231,N_4263);
nor U4838 (N_4838,N_4311,N_4018);
nor U4839 (N_4839,N_4497,N_4106);
xor U4840 (N_4840,N_4118,N_4327);
and U4841 (N_4841,N_4217,N_4493);
nand U4842 (N_4842,N_4278,N_4110);
nand U4843 (N_4843,N_4268,N_4347);
nor U4844 (N_4844,N_4374,N_4175);
or U4845 (N_4845,N_4038,N_4177);
nand U4846 (N_4846,N_4211,N_4173);
nand U4847 (N_4847,N_4062,N_4127);
and U4848 (N_4848,N_4465,N_4137);
and U4849 (N_4849,N_4432,N_4440);
and U4850 (N_4850,N_4435,N_4409);
nor U4851 (N_4851,N_4349,N_4115);
and U4852 (N_4852,N_4049,N_4442);
or U4853 (N_4853,N_4257,N_4083);
and U4854 (N_4854,N_4039,N_4257);
and U4855 (N_4855,N_4032,N_4015);
nor U4856 (N_4856,N_4324,N_4458);
xnor U4857 (N_4857,N_4097,N_4378);
nor U4858 (N_4858,N_4032,N_4423);
or U4859 (N_4859,N_4024,N_4389);
or U4860 (N_4860,N_4042,N_4300);
and U4861 (N_4861,N_4022,N_4318);
or U4862 (N_4862,N_4388,N_4436);
nor U4863 (N_4863,N_4372,N_4184);
nor U4864 (N_4864,N_4282,N_4220);
nand U4865 (N_4865,N_4160,N_4447);
or U4866 (N_4866,N_4232,N_4006);
or U4867 (N_4867,N_4099,N_4027);
and U4868 (N_4868,N_4375,N_4295);
nand U4869 (N_4869,N_4388,N_4102);
xor U4870 (N_4870,N_4103,N_4393);
nor U4871 (N_4871,N_4396,N_4106);
nand U4872 (N_4872,N_4453,N_4039);
xor U4873 (N_4873,N_4026,N_4159);
or U4874 (N_4874,N_4322,N_4430);
or U4875 (N_4875,N_4215,N_4470);
and U4876 (N_4876,N_4001,N_4384);
or U4877 (N_4877,N_4366,N_4094);
and U4878 (N_4878,N_4431,N_4179);
nand U4879 (N_4879,N_4157,N_4433);
or U4880 (N_4880,N_4238,N_4081);
nand U4881 (N_4881,N_4164,N_4221);
nor U4882 (N_4882,N_4044,N_4189);
and U4883 (N_4883,N_4484,N_4260);
and U4884 (N_4884,N_4310,N_4128);
nand U4885 (N_4885,N_4160,N_4468);
nor U4886 (N_4886,N_4223,N_4125);
and U4887 (N_4887,N_4068,N_4152);
nand U4888 (N_4888,N_4442,N_4172);
and U4889 (N_4889,N_4395,N_4355);
nor U4890 (N_4890,N_4267,N_4097);
and U4891 (N_4891,N_4425,N_4173);
or U4892 (N_4892,N_4399,N_4116);
or U4893 (N_4893,N_4050,N_4368);
nor U4894 (N_4894,N_4299,N_4124);
or U4895 (N_4895,N_4262,N_4056);
or U4896 (N_4896,N_4322,N_4366);
nand U4897 (N_4897,N_4240,N_4131);
nand U4898 (N_4898,N_4273,N_4253);
nand U4899 (N_4899,N_4424,N_4337);
nor U4900 (N_4900,N_4328,N_4255);
nand U4901 (N_4901,N_4108,N_4271);
or U4902 (N_4902,N_4495,N_4236);
xnor U4903 (N_4903,N_4085,N_4406);
nor U4904 (N_4904,N_4169,N_4304);
nand U4905 (N_4905,N_4497,N_4362);
and U4906 (N_4906,N_4442,N_4434);
or U4907 (N_4907,N_4270,N_4345);
and U4908 (N_4908,N_4392,N_4080);
nor U4909 (N_4909,N_4424,N_4064);
nor U4910 (N_4910,N_4064,N_4413);
nand U4911 (N_4911,N_4081,N_4294);
or U4912 (N_4912,N_4135,N_4489);
nor U4913 (N_4913,N_4052,N_4282);
nor U4914 (N_4914,N_4198,N_4154);
nor U4915 (N_4915,N_4020,N_4241);
nor U4916 (N_4916,N_4105,N_4463);
nand U4917 (N_4917,N_4278,N_4176);
nor U4918 (N_4918,N_4140,N_4350);
nand U4919 (N_4919,N_4264,N_4338);
nand U4920 (N_4920,N_4446,N_4132);
xor U4921 (N_4921,N_4488,N_4142);
and U4922 (N_4922,N_4050,N_4346);
nor U4923 (N_4923,N_4115,N_4215);
nand U4924 (N_4924,N_4082,N_4178);
nor U4925 (N_4925,N_4118,N_4245);
and U4926 (N_4926,N_4475,N_4031);
nand U4927 (N_4927,N_4412,N_4137);
nand U4928 (N_4928,N_4218,N_4227);
nand U4929 (N_4929,N_4083,N_4134);
nor U4930 (N_4930,N_4310,N_4004);
and U4931 (N_4931,N_4046,N_4144);
xnor U4932 (N_4932,N_4341,N_4282);
nor U4933 (N_4933,N_4288,N_4089);
nor U4934 (N_4934,N_4003,N_4256);
and U4935 (N_4935,N_4283,N_4271);
nand U4936 (N_4936,N_4366,N_4024);
and U4937 (N_4937,N_4207,N_4280);
and U4938 (N_4938,N_4468,N_4320);
nor U4939 (N_4939,N_4243,N_4195);
and U4940 (N_4940,N_4127,N_4000);
nand U4941 (N_4941,N_4004,N_4471);
nand U4942 (N_4942,N_4082,N_4152);
and U4943 (N_4943,N_4234,N_4074);
nor U4944 (N_4944,N_4023,N_4458);
nor U4945 (N_4945,N_4171,N_4344);
and U4946 (N_4946,N_4086,N_4444);
nor U4947 (N_4947,N_4132,N_4471);
xnor U4948 (N_4948,N_4021,N_4241);
nand U4949 (N_4949,N_4095,N_4270);
nand U4950 (N_4950,N_4041,N_4097);
or U4951 (N_4951,N_4147,N_4072);
or U4952 (N_4952,N_4032,N_4165);
or U4953 (N_4953,N_4377,N_4055);
and U4954 (N_4954,N_4343,N_4035);
and U4955 (N_4955,N_4107,N_4151);
and U4956 (N_4956,N_4212,N_4046);
nor U4957 (N_4957,N_4124,N_4148);
nand U4958 (N_4958,N_4185,N_4322);
nor U4959 (N_4959,N_4265,N_4295);
nor U4960 (N_4960,N_4267,N_4469);
and U4961 (N_4961,N_4092,N_4187);
and U4962 (N_4962,N_4071,N_4026);
xor U4963 (N_4963,N_4168,N_4362);
and U4964 (N_4964,N_4282,N_4333);
nor U4965 (N_4965,N_4051,N_4456);
or U4966 (N_4966,N_4357,N_4485);
and U4967 (N_4967,N_4479,N_4102);
nand U4968 (N_4968,N_4332,N_4387);
nand U4969 (N_4969,N_4326,N_4397);
nand U4970 (N_4970,N_4103,N_4345);
nand U4971 (N_4971,N_4447,N_4007);
or U4972 (N_4972,N_4150,N_4306);
or U4973 (N_4973,N_4011,N_4446);
nand U4974 (N_4974,N_4496,N_4211);
nor U4975 (N_4975,N_4063,N_4204);
nor U4976 (N_4976,N_4078,N_4432);
or U4977 (N_4977,N_4014,N_4202);
nand U4978 (N_4978,N_4105,N_4373);
or U4979 (N_4979,N_4103,N_4091);
or U4980 (N_4980,N_4312,N_4261);
nand U4981 (N_4981,N_4389,N_4426);
xor U4982 (N_4982,N_4343,N_4140);
or U4983 (N_4983,N_4225,N_4117);
or U4984 (N_4984,N_4086,N_4153);
xnor U4985 (N_4985,N_4284,N_4361);
nand U4986 (N_4986,N_4065,N_4470);
and U4987 (N_4987,N_4415,N_4482);
or U4988 (N_4988,N_4469,N_4131);
nand U4989 (N_4989,N_4004,N_4244);
or U4990 (N_4990,N_4276,N_4103);
nor U4991 (N_4991,N_4104,N_4086);
or U4992 (N_4992,N_4152,N_4103);
nor U4993 (N_4993,N_4070,N_4425);
nor U4994 (N_4994,N_4193,N_4274);
nor U4995 (N_4995,N_4119,N_4216);
xor U4996 (N_4996,N_4357,N_4455);
nand U4997 (N_4997,N_4483,N_4318);
nand U4998 (N_4998,N_4489,N_4342);
nand U4999 (N_4999,N_4130,N_4445);
nand UO_0 (O_0,N_4643,N_4862);
or UO_1 (O_1,N_4715,N_4562);
and UO_2 (O_2,N_4739,N_4778);
nor UO_3 (O_3,N_4842,N_4579);
nand UO_4 (O_4,N_4960,N_4875);
nor UO_5 (O_5,N_4935,N_4798);
and UO_6 (O_6,N_4867,N_4811);
or UO_7 (O_7,N_4527,N_4561);
or UO_8 (O_8,N_4959,N_4830);
nand UO_9 (O_9,N_4767,N_4815);
or UO_10 (O_10,N_4761,N_4922);
nand UO_11 (O_11,N_4760,N_4841);
nor UO_12 (O_12,N_4729,N_4965);
or UO_13 (O_13,N_4551,N_4619);
nand UO_14 (O_14,N_4907,N_4745);
or UO_15 (O_15,N_4649,N_4824);
xnor UO_16 (O_16,N_4775,N_4637);
nor UO_17 (O_17,N_4972,N_4553);
and UO_18 (O_18,N_4709,N_4532);
xnor UO_19 (O_19,N_4512,N_4791);
nand UO_20 (O_20,N_4829,N_4944);
nand UO_21 (O_21,N_4808,N_4873);
nor UO_22 (O_22,N_4618,N_4956);
or UO_23 (O_23,N_4584,N_4894);
or UO_24 (O_24,N_4810,N_4931);
nor UO_25 (O_25,N_4847,N_4547);
and UO_26 (O_26,N_4889,N_4840);
xor UO_27 (O_27,N_4777,N_4999);
nor UO_28 (O_28,N_4518,N_4945);
or UO_29 (O_29,N_4557,N_4742);
nor UO_30 (O_30,N_4912,N_4689);
and UO_31 (O_31,N_4628,N_4664);
xnor UO_32 (O_32,N_4642,N_4913);
nor UO_33 (O_33,N_4874,N_4770);
or UO_34 (O_34,N_4805,N_4502);
nand UO_35 (O_35,N_4638,N_4757);
or UO_36 (O_36,N_4596,N_4820);
or UO_37 (O_37,N_4536,N_4632);
nand UO_38 (O_38,N_4865,N_4995);
and UO_39 (O_39,N_4702,N_4747);
or UO_40 (O_40,N_4564,N_4860);
xor UO_41 (O_41,N_4634,N_4899);
and UO_42 (O_42,N_4881,N_4656);
or UO_43 (O_43,N_4538,N_4831);
or UO_44 (O_44,N_4968,N_4733);
nand UO_45 (O_45,N_4686,N_4648);
or UO_46 (O_46,N_4546,N_4726);
nand UO_47 (O_47,N_4776,N_4950);
nor UO_48 (O_48,N_4615,N_4629);
nand UO_49 (O_49,N_4684,N_4545);
or UO_50 (O_50,N_4550,N_4580);
nor UO_51 (O_51,N_4660,N_4687);
or UO_52 (O_52,N_4974,N_4571);
nor UO_53 (O_53,N_4923,N_4940);
and UO_54 (O_54,N_4523,N_4773);
or UO_55 (O_55,N_4958,N_4688);
nor UO_56 (O_56,N_4762,N_4574);
nor UO_57 (O_57,N_4713,N_4707);
nor UO_58 (O_58,N_4743,N_4736);
nor UO_59 (O_59,N_4855,N_4951);
nor UO_60 (O_60,N_4758,N_4908);
nor UO_61 (O_61,N_4575,N_4671);
nand UO_62 (O_62,N_4700,N_4966);
nand UO_63 (O_63,N_4802,N_4978);
nand UO_64 (O_64,N_4516,N_4524);
nand UO_65 (O_65,N_4566,N_4568);
nand UO_66 (O_66,N_4756,N_4916);
nor UO_67 (O_67,N_4576,N_4549);
or UO_68 (O_68,N_4941,N_4506);
nor UO_69 (O_69,N_4511,N_4926);
or UO_70 (O_70,N_4719,N_4633);
or UO_71 (O_71,N_4987,N_4787);
and UO_72 (O_72,N_4559,N_4592);
nand UO_73 (O_73,N_4980,N_4533);
nor UO_74 (O_74,N_4990,N_4540);
or UO_75 (O_75,N_4902,N_4765);
or UO_76 (O_76,N_4970,N_4668);
or UO_77 (O_77,N_4590,N_4854);
nor UO_78 (O_78,N_4883,N_4716);
nor UO_79 (O_79,N_4784,N_4803);
or UO_80 (O_80,N_4799,N_4613);
nand UO_81 (O_81,N_4779,N_4896);
xor UO_82 (O_82,N_4657,N_4816);
nor UO_83 (O_83,N_4949,N_4578);
nand UO_84 (O_84,N_4645,N_4911);
xnor UO_85 (O_85,N_4626,N_4586);
nand UO_86 (O_86,N_4714,N_4885);
nand UO_87 (O_87,N_4953,N_4955);
nand UO_88 (O_88,N_4833,N_4611);
nor UO_89 (O_89,N_4988,N_4558);
nand UO_90 (O_90,N_4772,N_4582);
nor UO_91 (O_91,N_4903,N_4543);
or UO_92 (O_92,N_4555,N_4720);
nor UO_93 (O_93,N_4795,N_4676);
nand UO_94 (O_94,N_4727,N_4893);
nor UO_95 (O_95,N_4869,N_4814);
nor UO_96 (O_96,N_4690,N_4917);
nand UO_97 (O_97,N_4663,N_4853);
xor UO_98 (O_98,N_4539,N_4868);
or UO_99 (O_99,N_4588,N_4674);
nand UO_100 (O_100,N_4530,N_4548);
or UO_101 (O_101,N_4598,N_4905);
or UO_102 (O_102,N_4909,N_4969);
and UO_103 (O_103,N_4813,N_4501);
nand UO_104 (O_104,N_4694,N_4669);
or UO_105 (O_105,N_4748,N_4892);
nand UO_106 (O_106,N_4740,N_4781);
nand UO_107 (O_107,N_4871,N_4658);
and UO_108 (O_108,N_4672,N_4839);
or UO_109 (O_109,N_4741,N_4888);
nor UO_110 (O_110,N_4610,N_4886);
nand UO_111 (O_111,N_4946,N_4744);
nand UO_112 (O_112,N_4738,N_4717);
and UO_113 (O_113,N_4534,N_4856);
nor UO_114 (O_114,N_4675,N_4603);
or UO_115 (O_115,N_4753,N_4992);
xnor UO_116 (O_116,N_4783,N_4641);
and UO_117 (O_117,N_4652,N_4529);
or UO_118 (O_118,N_4920,N_4774);
and UO_119 (O_119,N_4622,N_4918);
and UO_120 (O_120,N_4806,N_4947);
xnor UO_121 (O_121,N_4693,N_4754);
nand UO_122 (O_122,N_4796,N_4838);
or UO_123 (O_123,N_4979,N_4595);
or UO_124 (O_124,N_4927,N_4976);
and UO_125 (O_125,N_4639,N_4565);
and UO_126 (O_126,N_4901,N_4679);
xor UO_127 (O_127,N_4967,N_4665);
nor UO_128 (O_128,N_4678,N_4851);
xor UO_129 (O_129,N_4725,N_4769);
xor UO_130 (O_130,N_4997,N_4528);
nand UO_131 (O_131,N_4952,N_4554);
nor UO_132 (O_132,N_4573,N_4877);
nor UO_133 (O_133,N_4597,N_4680);
or UO_134 (O_134,N_4520,N_4957);
nand UO_135 (O_135,N_4500,N_4517);
nor UO_136 (O_136,N_4934,N_4964);
nor UO_137 (O_137,N_4801,N_4925);
and UO_138 (O_138,N_4569,N_4504);
nand UO_139 (O_139,N_4789,N_4560);
and UO_140 (O_140,N_4794,N_4503);
xnor UO_141 (O_141,N_4937,N_4975);
nand UO_142 (O_142,N_4818,N_4939);
nor UO_143 (O_143,N_4887,N_4699);
nand UO_144 (O_144,N_4531,N_4526);
nand UO_145 (O_145,N_4681,N_4915);
nand UO_146 (O_146,N_4698,N_4552);
nand UO_147 (O_147,N_4788,N_4817);
nor UO_148 (O_148,N_4822,N_4973);
nor UO_149 (O_149,N_4910,N_4906);
nand UO_150 (O_150,N_4749,N_4751);
or UO_151 (O_151,N_4836,N_4605);
nand UO_152 (O_152,N_4515,N_4542);
and UO_153 (O_153,N_4832,N_4882);
nor UO_154 (O_154,N_4858,N_4696);
nand UO_155 (O_155,N_4591,N_4601);
or UO_156 (O_156,N_4982,N_4864);
or UO_157 (O_157,N_4895,N_4567);
xnor UO_158 (O_158,N_4544,N_4932);
or UO_159 (O_159,N_4505,N_4857);
nand UO_160 (O_160,N_4606,N_4848);
or UO_161 (O_161,N_4635,N_4650);
or UO_162 (O_162,N_4572,N_4942);
or UO_163 (O_163,N_4695,N_4723);
nand UO_164 (O_164,N_4609,N_4730);
nor UO_165 (O_165,N_4616,N_4933);
xor UO_166 (O_166,N_4786,N_4667);
and UO_167 (O_167,N_4921,N_4846);
nor UO_168 (O_168,N_4627,N_4682);
nor UO_169 (O_169,N_4535,N_4706);
or UO_170 (O_170,N_4697,N_4670);
nand UO_171 (O_171,N_4614,N_4845);
or UO_172 (O_172,N_4989,N_4710);
or UO_173 (O_173,N_4625,N_4624);
nor UO_174 (O_174,N_4800,N_4859);
or UO_175 (O_175,N_4589,N_4993);
or UO_176 (O_176,N_4708,N_4604);
or UO_177 (O_177,N_4938,N_4826);
nand UO_178 (O_178,N_4585,N_4984);
xor UO_179 (O_179,N_4876,N_4711);
or UO_180 (O_180,N_4662,N_4904);
nand UO_181 (O_181,N_4631,N_4837);
and UO_182 (O_182,N_4936,N_4691);
xnor UO_183 (O_183,N_4771,N_4793);
or UO_184 (O_184,N_4666,N_4807);
nand UO_185 (O_185,N_4519,N_4701);
nor UO_186 (O_186,N_4620,N_4866);
nor UO_187 (O_187,N_4985,N_4728);
and UO_188 (O_188,N_4659,N_4850);
or UO_189 (O_189,N_4834,N_4821);
nand UO_190 (O_190,N_4943,N_4705);
and UO_191 (O_191,N_4570,N_4509);
xor UO_192 (O_192,N_4843,N_4792);
nand UO_193 (O_193,N_4928,N_4653);
or UO_194 (O_194,N_4819,N_4891);
nand UO_195 (O_195,N_4704,N_4522);
nor UO_196 (O_196,N_4685,N_4594);
or UO_197 (O_197,N_4825,N_4812);
or UO_198 (O_198,N_4963,N_4924);
and UO_199 (O_199,N_4661,N_4986);
nand UO_200 (O_200,N_4612,N_4655);
or UO_201 (O_201,N_4884,N_4654);
or UO_202 (O_202,N_4673,N_4961);
xnor UO_203 (O_203,N_4581,N_4537);
nor UO_204 (O_204,N_4898,N_4731);
nand UO_205 (O_205,N_4750,N_4804);
nand UO_206 (O_206,N_4577,N_4718);
nor UO_207 (O_207,N_4828,N_4724);
nor UO_208 (O_208,N_4863,N_4879);
nor UO_209 (O_209,N_4737,N_4556);
or UO_210 (O_210,N_4644,N_4890);
and UO_211 (O_211,N_4763,N_4593);
nand UO_212 (O_212,N_4599,N_4563);
nor UO_213 (O_213,N_4617,N_4513);
and UO_214 (O_214,N_4514,N_4994);
nand UO_215 (O_215,N_4991,N_4948);
and UO_216 (O_216,N_4608,N_4823);
or UO_217 (O_217,N_4878,N_4766);
or UO_218 (O_218,N_4630,N_4919);
xor UO_219 (O_219,N_4797,N_4683);
nor UO_220 (O_220,N_4962,N_4755);
or UO_221 (O_221,N_4647,N_4600);
nor UO_222 (O_222,N_4752,N_4983);
and UO_223 (O_223,N_4809,N_4692);
nand UO_224 (O_224,N_4977,N_4677);
xnor UO_225 (O_225,N_4712,N_4722);
or UO_226 (O_226,N_4521,N_4827);
or UO_227 (O_227,N_4930,N_4703);
or UO_228 (O_228,N_4607,N_4525);
nor UO_229 (O_229,N_4785,N_4651);
xor UO_230 (O_230,N_4768,N_4583);
nand UO_231 (O_231,N_4621,N_4861);
nand UO_232 (O_232,N_4849,N_4870);
or UO_233 (O_233,N_4844,N_4880);
nor UO_234 (O_234,N_4587,N_4640);
and UO_235 (O_235,N_4998,N_4636);
or UO_236 (O_236,N_4971,N_4541);
or UO_237 (O_237,N_4900,N_4996);
nand UO_238 (O_238,N_4790,N_4764);
or UO_239 (O_239,N_4508,N_4780);
nand UO_240 (O_240,N_4646,N_4897);
nand UO_241 (O_241,N_4602,N_4835);
xor UO_242 (O_242,N_4981,N_4510);
or UO_243 (O_243,N_4721,N_4735);
and UO_244 (O_244,N_4782,N_4732);
nand UO_245 (O_245,N_4507,N_4852);
and UO_246 (O_246,N_4872,N_4914);
and UO_247 (O_247,N_4734,N_4929);
nand UO_248 (O_248,N_4759,N_4746);
nor UO_249 (O_249,N_4623,N_4954);
xor UO_250 (O_250,N_4860,N_4693);
nand UO_251 (O_251,N_4622,N_4971);
or UO_252 (O_252,N_4963,N_4547);
or UO_253 (O_253,N_4992,N_4613);
and UO_254 (O_254,N_4946,N_4599);
or UO_255 (O_255,N_4703,N_4926);
nor UO_256 (O_256,N_4929,N_4896);
and UO_257 (O_257,N_4933,N_4554);
or UO_258 (O_258,N_4864,N_4655);
or UO_259 (O_259,N_4502,N_4914);
nand UO_260 (O_260,N_4795,N_4606);
nor UO_261 (O_261,N_4508,N_4711);
nor UO_262 (O_262,N_4618,N_4556);
nand UO_263 (O_263,N_4750,N_4807);
or UO_264 (O_264,N_4963,N_4604);
and UO_265 (O_265,N_4769,N_4886);
xor UO_266 (O_266,N_4987,N_4776);
nor UO_267 (O_267,N_4914,N_4879);
or UO_268 (O_268,N_4755,N_4564);
nor UO_269 (O_269,N_4563,N_4576);
and UO_270 (O_270,N_4585,N_4923);
and UO_271 (O_271,N_4662,N_4961);
or UO_272 (O_272,N_4761,N_4763);
nor UO_273 (O_273,N_4855,N_4883);
or UO_274 (O_274,N_4727,N_4873);
and UO_275 (O_275,N_4601,N_4650);
nand UO_276 (O_276,N_4978,N_4581);
nand UO_277 (O_277,N_4872,N_4831);
nor UO_278 (O_278,N_4645,N_4669);
xor UO_279 (O_279,N_4578,N_4731);
nand UO_280 (O_280,N_4830,N_4581);
nand UO_281 (O_281,N_4650,N_4767);
or UO_282 (O_282,N_4977,N_4528);
and UO_283 (O_283,N_4755,N_4965);
xor UO_284 (O_284,N_4980,N_4732);
nand UO_285 (O_285,N_4706,N_4692);
xnor UO_286 (O_286,N_4736,N_4639);
or UO_287 (O_287,N_4657,N_4896);
and UO_288 (O_288,N_4657,N_4633);
or UO_289 (O_289,N_4988,N_4633);
nand UO_290 (O_290,N_4643,N_4749);
or UO_291 (O_291,N_4896,N_4946);
and UO_292 (O_292,N_4884,N_4712);
nand UO_293 (O_293,N_4894,N_4832);
or UO_294 (O_294,N_4759,N_4719);
nor UO_295 (O_295,N_4730,N_4620);
nor UO_296 (O_296,N_4977,N_4739);
nand UO_297 (O_297,N_4929,N_4797);
xnor UO_298 (O_298,N_4952,N_4840);
or UO_299 (O_299,N_4951,N_4680);
nand UO_300 (O_300,N_4924,N_4772);
or UO_301 (O_301,N_4632,N_4644);
or UO_302 (O_302,N_4883,N_4834);
or UO_303 (O_303,N_4748,N_4556);
and UO_304 (O_304,N_4645,N_4627);
and UO_305 (O_305,N_4691,N_4579);
nand UO_306 (O_306,N_4828,N_4501);
nor UO_307 (O_307,N_4532,N_4529);
and UO_308 (O_308,N_4778,N_4566);
or UO_309 (O_309,N_4938,N_4633);
nor UO_310 (O_310,N_4703,N_4932);
nor UO_311 (O_311,N_4753,N_4936);
nand UO_312 (O_312,N_4658,N_4668);
and UO_313 (O_313,N_4924,N_4911);
nand UO_314 (O_314,N_4976,N_4930);
or UO_315 (O_315,N_4707,N_4788);
or UO_316 (O_316,N_4848,N_4815);
nor UO_317 (O_317,N_4930,N_4512);
nand UO_318 (O_318,N_4676,N_4946);
nand UO_319 (O_319,N_4838,N_4946);
and UO_320 (O_320,N_4770,N_4546);
nor UO_321 (O_321,N_4716,N_4673);
nand UO_322 (O_322,N_4710,N_4903);
nand UO_323 (O_323,N_4848,N_4755);
xor UO_324 (O_324,N_4709,N_4909);
or UO_325 (O_325,N_4938,N_4679);
nor UO_326 (O_326,N_4687,N_4859);
nor UO_327 (O_327,N_4549,N_4964);
and UO_328 (O_328,N_4559,N_4823);
nor UO_329 (O_329,N_4862,N_4740);
nand UO_330 (O_330,N_4695,N_4712);
or UO_331 (O_331,N_4608,N_4654);
nor UO_332 (O_332,N_4890,N_4581);
and UO_333 (O_333,N_4557,N_4653);
nand UO_334 (O_334,N_4663,N_4852);
and UO_335 (O_335,N_4755,N_4805);
nand UO_336 (O_336,N_4817,N_4812);
nor UO_337 (O_337,N_4520,N_4738);
nand UO_338 (O_338,N_4891,N_4660);
or UO_339 (O_339,N_4757,N_4721);
and UO_340 (O_340,N_4940,N_4625);
nand UO_341 (O_341,N_4626,N_4608);
nor UO_342 (O_342,N_4813,N_4604);
nor UO_343 (O_343,N_4924,N_4860);
xor UO_344 (O_344,N_4609,N_4781);
nand UO_345 (O_345,N_4618,N_4576);
nand UO_346 (O_346,N_4619,N_4625);
xor UO_347 (O_347,N_4728,N_4616);
and UO_348 (O_348,N_4519,N_4652);
or UO_349 (O_349,N_4899,N_4982);
nand UO_350 (O_350,N_4677,N_4906);
and UO_351 (O_351,N_4500,N_4826);
or UO_352 (O_352,N_4746,N_4626);
or UO_353 (O_353,N_4755,N_4842);
xor UO_354 (O_354,N_4765,N_4534);
nand UO_355 (O_355,N_4741,N_4566);
xor UO_356 (O_356,N_4772,N_4832);
or UO_357 (O_357,N_4961,N_4893);
or UO_358 (O_358,N_4864,N_4524);
and UO_359 (O_359,N_4952,N_4930);
xor UO_360 (O_360,N_4767,N_4718);
nor UO_361 (O_361,N_4927,N_4533);
and UO_362 (O_362,N_4901,N_4993);
nand UO_363 (O_363,N_4869,N_4568);
xor UO_364 (O_364,N_4882,N_4965);
nor UO_365 (O_365,N_4621,N_4692);
and UO_366 (O_366,N_4612,N_4982);
and UO_367 (O_367,N_4929,N_4924);
or UO_368 (O_368,N_4938,N_4800);
nand UO_369 (O_369,N_4542,N_4635);
nor UO_370 (O_370,N_4514,N_4836);
xor UO_371 (O_371,N_4948,N_4573);
xor UO_372 (O_372,N_4752,N_4785);
nor UO_373 (O_373,N_4903,N_4807);
nor UO_374 (O_374,N_4583,N_4955);
or UO_375 (O_375,N_4868,N_4751);
nand UO_376 (O_376,N_4760,N_4738);
or UO_377 (O_377,N_4541,N_4835);
nor UO_378 (O_378,N_4583,N_4764);
or UO_379 (O_379,N_4995,N_4909);
or UO_380 (O_380,N_4715,N_4699);
nand UO_381 (O_381,N_4567,N_4788);
and UO_382 (O_382,N_4612,N_4555);
nor UO_383 (O_383,N_4616,N_4745);
xor UO_384 (O_384,N_4668,N_4768);
nor UO_385 (O_385,N_4980,N_4934);
nor UO_386 (O_386,N_4912,N_4878);
or UO_387 (O_387,N_4777,N_4739);
and UO_388 (O_388,N_4733,N_4757);
nor UO_389 (O_389,N_4590,N_4597);
and UO_390 (O_390,N_4742,N_4501);
and UO_391 (O_391,N_4763,N_4929);
and UO_392 (O_392,N_4921,N_4766);
xnor UO_393 (O_393,N_4796,N_4901);
and UO_394 (O_394,N_4690,N_4884);
xnor UO_395 (O_395,N_4743,N_4531);
and UO_396 (O_396,N_4668,N_4523);
xnor UO_397 (O_397,N_4948,N_4868);
nand UO_398 (O_398,N_4702,N_4708);
nand UO_399 (O_399,N_4693,N_4989);
and UO_400 (O_400,N_4783,N_4824);
xnor UO_401 (O_401,N_4919,N_4642);
or UO_402 (O_402,N_4568,N_4936);
nand UO_403 (O_403,N_4613,N_4565);
nand UO_404 (O_404,N_4989,N_4703);
or UO_405 (O_405,N_4796,N_4565);
or UO_406 (O_406,N_4864,N_4595);
or UO_407 (O_407,N_4640,N_4802);
nor UO_408 (O_408,N_4711,N_4654);
xnor UO_409 (O_409,N_4750,N_4571);
and UO_410 (O_410,N_4712,N_4777);
or UO_411 (O_411,N_4803,N_4975);
nor UO_412 (O_412,N_4592,N_4945);
or UO_413 (O_413,N_4526,N_4987);
nor UO_414 (O_414,N_4532,N_4511);
and UO_415 (O_415,N_4925,N_4605);
nor UO_416 (O_416,N_4933,N_4960);
and UO_417 (O_417,N_4597,N_4586);
nor UO_418 (O_418,N_4759,N_4920);
and UO_419 (O_419,N_4613,N_4820);
nor UO_420 (O_420,N_4831,N_4959);
nand UO_421 (O_421,N_4506,N_4968);
xnor UO_422 (O_422,N_4534,N_4696);
or UO_423 (O_423,N_4940,N_4832);
nand UO_424 (O_424,N_4589,N_4745);
and UO_425 (O_425,N_4674,N_4596);
nor UO_426 (O_426,N_4636,N_4973);
or UO_427 (O_427,N_4619,N_4662);
nor UO_428 (O_428,N_4847,N_4842);
nand UO_429 (O_429,N_4614,N_4991);
nor UO_430 (O_430,N_4554,N_4922);
nand UO_431 (O_431,N_4903,N_4933);
nand UO_432 (O_432,N_4628,N_4729);
xnor UO_433 (O_433,N_4852,N_4994);
xnor UO_434 (O_434,N_4833,N_4594);
nor UO_435 (O_435,N_4589,N_4826);
nand UO_436 (O_436,N_4778,N_4983);
nor UO_437 (O_437,N_4847,N_4777);
nand UO_438 (O_438,N_4832,N_4992);
xor UO_439 (O_439,N_4773,N_4903);
or UO_440 (O_440,N_4928,N_4525);
or UO_441 (O_441,N_4636,N_4535);
and UO_442 (O_442,N_4870,N_4761);
and UO_443 (O_443,N_4838,N_4938);
or UO_444 (O_444,N_4787,N_4716);
xor UO_445 (O_445,N_4629,N_4954);
nand UO_446 (O_446,N_4862,N_4902);
and UO_447 (O_447,N_4576,N_4981);
nor UO_448 (O_448,N_4633,N_4940);
nor UO_449 (O_449,N_4564,N_4741);
nor UO_450 (O_450,N_4559,N_4597);
and UO_451 (O_451,N_4701,N_4518);
nor UO_452 (O_452,N_4832,N_4922);
and UO_453 (O_453,N_4657,N_4983);
nand UO_454 (O_454,N_4743,N_4505);
nor UO_455 (O_455,N_4998,N_4750);
xor UO_456 (O_456,N_4539,N_4874);
xor UO_457 (O_457,N_4516,N_4783);
nor UO_458 (O_458,N_4686,N_4884);
nand UO_459 (O_459,N_4828,N_4536);
xnor UO_460 (O_460,N_4612,N_4724);
nand UO_461 (O_461,N_4632,N_4506);
and UO_462 (O_462,N_4656,N_4798);
or UO_463 (O_463,N_4973,N_4614);
or UO_464 (O_464,N_4586,N_4539);
nor UO_465 (O_465,N_4560,N_4814);
nand UO_466 (O_466,N_4878,N_4859);
nor UO_467 (O_467,N_4725,N_4831);
nor UO_468 (O_468,N_4964,N_4538);
nor UO_469 (O_469,N_4773,N_4676);
and UO_470 (O_470,N_4986,N_4501);
nand UO_471 (O_471,N_4742,N_4706);
or UO_472 (O_472,N_4775,N_4988);
xor UO_473 (O_473,N_4870,N_4787);
nand UO_474 (O_474,N_4572,N_4686);
or UO_475 (O_475,N_4572,N_4749);
nand UO_476 (O_476,N_4987,N_4657);
or UO_477 (O_477,N_4713,N_4932);
nand UO_478 (O_478,N_4750,N_4950);
nor UO_479 (O_479,N_4854,N_4580);
and UO_480 (O_480,N_4980,N_4744);
nor UO_481 (O_481,N_4892,N_4870);
or UO_482 (O_482,N_4717,N_4958);
or UO_483 (O_483,N_4690,N_4786);
nand UO_484 (O_484,N_4837,N_4521);
nand UO_485 (O_485,N_4610,N_4735);
and UO_486 (O_486,N_4839,N_4921);
or UO_487 (O_487,N_4891,N_4525);
nand UO_488 (O_488,N_4759,N_4892);
and UO_489 (O_489,N_4580,N_4605);
and UO_490 (O_490,N_4639,N_4631);
nor UO_491 (O_491,N_4793,N_4898);
nand UO_492 (O_492,N_4523,N_4994);
nand UO_493 (O_493,N_4517,N_4507);
or UO_494 (O_494,N_4873,N_4710);
nand UO_495 (O_495,N_4615,N_4699);
and UO_496 (O_496,N_4906,N_4600);
and UO_497 (O_497,N_4697,N_4900);
nand UO_498 (O_498,N_4917,N_4837);
nor UO_499 (O_499,N_4782,N_4633);
nand UO_500 (O_500,N_4948,N_4565);
nand UO_501 (O_501,N_4548,N_4661);
nand UO_502 (O_502,N_4739,N_4947);
nand UO_503 (O_503,N_4922,N_4856);
and UO_504 (O_504,N_4989,N_4871);
or UO_505 (O_505,N_4548,N_4794);
or UO_506 (O_506,N_4652,N_4635);
nand UO_507 (O_507,N_4563,N_4529);
nand UO_508 (O_508,N_4525,N_4824);
xnor UO_509 (O_509,N_4732,N_4566);
xor UO_510 (O_510,N_4558,N_4589);
nand UO_511 (O_511,N_4547,N_4904);
xor UO_512 (O_512,N_4739,N_4504);
nor UO_513 (O_513,N_4949,N_4779);
nand UO_514 (O_514,N_4891,N_4765);
nor UO_515 (O_515,N_4661,N_4789);
nor UO_516 (O_516,N_4578,N_4711);
xnor UO_517 (O_517,N_4660,N_4992);
xor UO_518 (O_518,N_4801,N_4833);
xor UO_519 (O_519,N_4856,N_4882);
and UO_520 (O_520,N_4649,N_4963);
nor UO_521 (O_521,N_4799,N_4624);
nor UO_522 (O_522,N_4717,N_4669);
nor UO_523 (O_523,N_4751,N_4986);
or UO_524 (O_524,N_4798,N_4941);
and UO_525 (O_525,N_4759,N_4782);
and UO_526 (O_526,N_4717,N_4677);
nand UO_527 (O_527,N_4573,N_4809);
and UO_528 (O_528,N_4923,N_4922);
or UO_529 (O_529,N_4646,N_4537);
nor UO_530 (O_530,N_4675,N_4570);
nand UO_531 (O_531,N_4631,N_4901);
nor UO_532 (O_532,N_4750,N_4845);
nand UO_533 (O_533,N_4900,N_4527);
nand UO_534 (O_534,N_4658,N_4548);
and UO_535 (O_535,N_4734,N_4672);
or UO_536 (O_536,N_4768,N_4667);
and UO_537 (O_537,N_4859,N_4592);
and UO_538 (O_538,N_4586,N_4521);
nand UO_539 (O_539,N_4601,N_4679);
or UO_540 (O_540,N_4709,N_4917);
nand UO_541 (O_541,N_4633,N_4572);
or UO_542 (O_542,N_4655,N_4508);
and UO_543 (O_543,N_4500,N_4752);
nor UO_544 (O_544,N_4959,N_4894);
xnor UO_545 (O_545,N_4867,N_4752);
or UO_546 (O_546,N_4834,N_4940);
and UO_547 (O_547,N_4826,N_4568);
nor UO_548 (O_548,N_4840,N_4612);
nand UO_549 (O_549,N_4536,N_4832);
xor UO_550 (O_550,N_4813,N_4526);
nand UO_551 (O_551,N_4723,N_4530);
nand UO_552 (O_552,N_4988,N_4792);
nand UO_553 (O_553,N_4763,N_4737);
or UO_554 (O_554,N_4582,N_4889);
nor UO_555 (O_555,N_4639,N_4857);
and UO_556 (O_556,N_4916,N_4561);
or UO_557 (O_557,N_4934,N_4700);
nor UO_558 (O_558,N_4872,N_4693);
nor UO_559 (O_559,N_4567,N_4922);
and UO_560 (O_560,N_4666,N_4856);
or UO_561 (O_561,N_4628,N_4991);
xor UO_562 (O_562,N_4931,N_4523);
or UO_563 (O_563,N_4933,N_4799);
nand UO_564 (O_564,N_4820,N_4980);
nor UO_565 (O_565,N_4645,N_4705);
nor UO_566 (O_566,N_4629,N_4723);
nand UO_567 (O_567,N_4630,N_4790);
nor UO_568 (O_568,N_4979,N_4658);
nor UO_569 (O_569,N_4596,N_4918);
or UO_570 (O_570,N_4846,N_4630);
nand UO_571 (O_571,N_4629,N_4503);
nand UO_572 (O_572,N_4697,N_4856);
nand UO_573 (O_573,N_4553,N_4893);
and UO_574 (O_574,N_4970,N_4577);
nand UO_575 (O_575,N_4628,N_4813);
and UO_576 (O_576,N_4508,N_4846);
nor UO_577 (O_577,N_4614,N_4719);
nor UO_578 (O_578,N_4863,N_4824);
nor UO_579 (O_579,N_4874,N_4908);
and UO_580 (O_580,N_4908,N_4918);
and UO_581 (O_581,N_4513,N_4768);
nor UO_582 (O_582,N_4709,N_4963);
or UO_583 (O_583,N_4610,N_4936);
or UO_584 (O_584,N_4836,N_4556);
or UO_585 (O_585,N_4989,N_4829);
or UO_586 (O_586,N_4796,N_4819);
xor UO_587 (O_587,N_4739,N_4992);
and UO_588 (O_588,N_4756,N_4731);
or UO_589 (O_589,N_4623,N_4859);
nand UO_590 (O_590,N_4635,N_4651);
or UO_591 (O_591,N_4693,N_4837);
or UO_592 (O_592,N_4667,N_4802);
nand UO_593 (O_593,N_4896,N_4819);
or UO_594 (O_594,N_4542,N_4649);
nand UO_595 (O_595,N_4692,N_4892);
nor UO_596 (O_596,N_4769,N_4859);
or UO_597 (O_597,N_4821,N_4559);
or UO_598 (O_598,N_4753,N_4879);
or UO_599 (O_599,N_4605,N_4682);
or UO_600 (O_600,N_4932,N_4657);
xnor UO_601 (O_601,N_4775,N_4646);
and UO_602 (O_602,N_4653,N_4919);
or UO_603 (O_603,N_4763,N_4591);
and UO_604 (O_604,N_4512,N_4844);
nor UO_605 (O_605,N_4983,N_4912);
nor UO_606 (O_606,N_4690,N_4588);
nand UO_607 (O_607,N_4780,N_4851);
and UO_608 (O_608,N_4606,N_4828);
xnor UO_609 (O_609,N_4559,N_4848);
nor UO_610 (O_610,N_4922,N_4786);
or UO_611 (O_611,N_4590,N_4631);
nand UO_612 (O_612,N_4957,N_4892);
and UO_613 (O_613,N_4562,N_4911);
nand UO_614 (O_614,N_4929,N_4808);
or UO_615 (O_615,N_4821,N_4956);
nand UO_616 (O_616,N_4900,N_4643);
or UO_617 (O_617,N_4731,N_4515);
nor UO_618 (O_618,N_4701,N_4682);
nor UO_619 (O_619,N_4716,N_4607);
nor UO_620 (O_620,N_4554,N_4631);
xor UO_621 (O_621,N_4602,N_4852);
nor UO_622 (O_622,N_4518,N_4660);
or UO_623 (O_623,N_4639,N_4780);
and UO_624 (O_624,N_4723,N_4521);
or UO_625 (O_625,N_4934,N_4993);
or UO_626 (O_626,N_4539,N_4847);
and UO_627 (O_627,N_4744,N_4846);
nand UO_628 (O_628,N_4835,N_4658);
nand UO_629 (O_629,N_4620,N_4896);
and UO_630 (O_630,N_4891,N_4600);
nand UO_631 (O_631,N_4578,N_4536);
or UO_632 (O_632,N_4728,N_4649);
nand UO_633 (O_633,N_4683,N_4575);
nand UO_634 (O_634,N_4695,N_4877);
nand UO_635 (O_635,N_4779,N_4704);
xor UO_636 (O_636,N_4521,N_4843);
nor UO_637 (O_637,N_4960,N_4649);
nor UO_638 (O_638,N_4631,N_4925);
nor UO_639 (O_639,N_4936,N_4540);
nor UO_640 (O_640,N_4771,N_4669);
or UO_641 (O_641,N_4891,N_4534);
and UO_642 (O_642,N_4906,N_4859);
or UO_643 (O_643,N_4515,N_4958);
and UO_644 (O_644,N_4602,N_4818);
and UO_645 (O_645,N_4577,N_4611);
xnor UO_646 (O_646,N_4830,N_4936);
or UO_647 (O_647,N_4625,N_4990);
and UO_648 (O_648,N_4896,N_4844);
and UO_649 (O_649,N_4537,N_4812);
nor UO_650 (O_650,N_4966,N_4710);
nand UO_651 (O_651,N_4660,N_4809);
or UO_652 (O_652,N_4962,N_4951);
and UO_653 (O_653,N_4740,N_4865);
and UO_654 (O_654,N_4668,N_4959);
nand UO_655 (O_655,N_4526,N_4721);
nor UO_656 (O_656,N_4881,N_4859);
nand UO_657 (O_657,N_4774,N_4897);
or UO_658 (O_658,N_4559,N_4862);
xor UO_659 (O_659,N_4610,N_4585);
nor UO_660 (O_660,N_4579,N_4932);
nor UO_661 (O_661,N_4916,N_4841);
and UO_662 (O_662,N_4883,N_4680);
nand UO_663 (O_663,N_4899,N_4665);
nor UO_664 (O_664,N_4857,N_4660);
and UO_665 (O_665,N_4511,N_4843);
and UO_666 (O_666,N_4820,N_4848);
and UO_667 (O_667,N_4899,N_4605);
and UO_668 (O_668,N_4759,N_4509);
or UO_669 (O_669,N_4613,N_4642);
or UO_670 (O_670,N_4639,N_4761);
and UO_671 (O_671,N_4501,N_4691);
nand UO_672 (O_672,N_4751,N_4821);
or UO_673 (O_673,N_4878,N_4945);
and UO_674 (O_674,N_4551,N_4685);
or UO_675 (O_675,N_4723,N_4651);
and UO_676 (O_676,N_4907,N_4579);
or UO_677 (O_677,N_4999,N_4528);
nor UO_678 (O_678,N_4574,N_4627);
and UO_679 (O_679,N_4527,N_4960);
nor UO_680 (O_680,N_4845,N_4706);
and UO_681 (O_681,N_4602,N_4749);
nand UO_682 (O_682,N_4750,N_4511);
and UO_683 (O_683,N_4904,N_4585);
nand UO_684 (O_684,N_4773,N_4595);
and UO_685 (O_685,N_4801,N_4637);
nand UO_686 (O_686,N_4656,N_4900);
nor UO_687 (O_687,N_4928,N_4710);
xor UO_688 (O_688,N_4852,N_4799);
or UO_689 (O_689,N_4910,N_4994);
and UO_690 (O_690,N_4752,N_4896);
nor UO_691 (O_691,N_4952,N_4642);
nor UO_692 (O_692,N_4753,N_4683);
nor UO_693 (O_693,N_4869,N_4592);
xnor UO_694 (O_694,N_4993,N_4672);
xor UO_695 (O_695,N_4968,N_4579);
or UO_696 (O_696,N_4941,N_4533);
nor UO_697 (O_697,N_4624,N_4906);
nand UO_698 (O_698,N_4788,N_4964);
and UO_699 (O_699,N_4945,N_4593);
and UO_700 (O_700,N_4976,N_4752);
and UO_701 (O_701,N_4625,N_4942);
and UO_702 (O_702,N_4994,N_4991);
and UO_703 (O_703,N_4629,N_4532);
or UO_704 (O_704,N_4554,N_4948);
and UO_705 (O_705,N_4504,N_4537);
nor UO_706 (O_706,N_4770,N_4845);
and UO_707 (O_707,N_4628,N_4931);
nor UO_708 (O_708,N_4897,N_4800);
nor UO_709 (O_709,N_4550,N_4747);
nand UO_710 (O_710,N_4680,N_4916);
or UO_711 (O_711,N_4850,N_4733);
nand UO_712 (O_712,N_4807,N_4815);
and UO_713 (O_713,N_4752,N_4675);
nand UO_714 (O_714,N_4829,N_4586);
nand UO_715 (O_715,N_4806,N_4879);
and UO_716 (O_716,N_4628,N_4976);
and UO_717 (O_717,N_4946,N_4966);
or UO_718 (O_718,N_4575,N_4708);
nor UO_719 (O_719,N_4643,N_4676);
nand UO_720 (O_720,N_4753,N_4898);
xor UO_721 (O_721,N_4600,N_4575);
or UO_722 (O_722,N_4775,N_4654);
nand UO_723 (O_723,N_4571,N_4807);
xnor UO_724 (O_724,N_4546,N_4663);
nor UO_725 (O_725,N_4797,N_4754);
nand UO_726 (O_726,N_4751,N_4851);
nor UO_727 (O_727,N_4830,N_4612);
or UO_728 (O_728,N_4909,N_4708);
nor UO_729 (O_729,N_4513,N_4986);
nand UO_730 (O_730,N_4541,N_4819);
nor UO_731 (O_731,N_4693,N_4727);
or UO_732 (O_732,N_4510,N_4666);
xnor UO_733 (O_733,N_4661,N_4715);
nand UO_734 (O_734,N_4813,N_4663);
xor UO_735 (O_735,N_4836,N_4632);
nor UO_736 (O_736,N_4607,N_4973);
and UO_737 (O_737,N_4529,N_4811);
nand UO_738 (O_738,N_4752,N_4672);
nand UO_739 (O_739,N_4976,N_4584);
or UO_740 (O_740,N_4840,N_4905);
or UO_741 (O_741,N_4963,N_4830);
and UO_742 (O_742,N_4976,N_4660);
or UO_743 (O_743,N_4699,N_4999);
nor UO_744 (O_744,N_4770,N_4611);
nand UO_745 (O_745,N_4674,N_4624);
and UO_746 (O_746,N_4569,N_4693);
or UO_747 (O_747,N_4846,N_4911);
xnor UO_748 (O_748,N_4696,N_4898);
xnor UO_749 (O_749,N_4816,N_4758);
or UO_750 (O_750,N_4750,N_4738);
nor UO_751 (O_751,N_4767,N_4765);
and UO_752 (O_752,N_4612,N_4967);
nor UO_753 (O_753,N_4524,N_4619);
xor UO_754 (O_754,N_4955,N_4958);
or UO_755 (O_755,N_4904,N_4876);
and UO_756 (O_756,N_4514,N_4682);
or UO_757 (O_757,N_4527,N_4611);
and UO_758 (O_758,N_4630,N_4547);
nand UO_759 (O_759,N_4789,N_4714);
nor UO_760 (O_760,N_4643,N_4819);
nand UO_761 (O_761,N_4947,N_4751);
nand UO_762 (O_762,N_4838,N_4657);
or UO_763 (O_763,N_4502,N_4681);
nand UO_764 (O_764,N_4916,N_4688);
nor UO_765 (O_765,N_4663,N_4500);
or UO_766 (O_766,N_4882,N_4875);
and UO_767 (O_767,N_4625,N_4870);
and UO_768 (O_768,N_4603,N_4958);
and UO_769 (O_769,N_4998,N_4708);
and UO_770 (O_770,N_4813,N_4606);
or UO_771 (O_771,N_4533,N_4950);
nor UO_772 (O_772,N_4628,N_4927);
xor UO_773 (O_773,N_4932,N_4653);
and UO_774 (O_774,N_4588,N_4840);
or UO_775 (O_775,N_4709,N_4589);
nor UO_776 (O_776,N_4986,N_4541);
or UO_777 (O_777,N_4716,N_4642);
and UO_778 (O_778,N_4633,N_4653);
nand UO_779 (O_779,N_4613,N_4705);
or UO_780 (O_780,N_4612,N_4780);
nor UO_781 (O_781,N_4896,N_4700);
nor UO_782 (O_782,N_4808,N_4514);
or UO_783 (O_783,N_4874,N_4698);
or UO_784 (O_784,N_4527,N_4573);
nand UO_785 (O_785,N_4710,N_4555);
or UO_786 (O_786,N_4944,N_4613);
or UO_787 (O_787,N_4691,N_4637);
and UO_788 (O_788,N_4574,N_4946);
nand UO_789 (O_789,N_4993,N_4903);
and UO_790 (O_790,N_4771,N_4656);
xor UO_791 (O_791,N_4545,N_4700);
and UO_792 (O_792,N_4963,N_4974);
nand UO_793 (O_793,N_4925,N_4691);
and UO_794 (O_794,N_4747,N_4689);
and UO_795 (O_795,N_4918,N_4746);
nand UO_796 (O_796,N_4916,N_4553);
nor UO_797 (O_797,N_4657,N_4772);
and UO_798 (O_798,N_4622,N_4850);
nor UO_799 (O_799,N_4787,N_4517);
nand UO_800 (O_800,N_4743,N_4591);
or UO_801 (O_801,N_4954,N_4756);
nand UO_802 (O_802,N_4573,N_4707);
or UO_803 (O_803,N_4800,N_4591);
or UO_804 (O_804,N_4759,N_4826);
nor UO_805 (O_805,N_4831,N_4693);
xnor UO_806 (O_806,N_4875,N_4689);
nand UO_807 (O_807,N_4720,N_4630);
nor UO_808 (O_808,N_4520,N_4570);
nor UO_809 (O_809,N_4657,N_4508);
nand UO_810 (O_810,N_4929,N_4585);
nand UO_811 (O_811,N_4634,N_4953);
nand UO_812 (O_812,N_4785,N_4761);
nand UO_813 (O_813,N_4857,N_4853);
nand UO_814 (O_814,N_4877,N_4882);
nand UO_815 (O_815,N_4742,N_4788);
xor UO_816 (O_816,N_4820,N_4701);
nor UO_817 (O_817,N_4813,N_4917);
xnor UO_818 (O_818,N_4642,N_4815);
nand UO_819 (O_819,N_4896,N_4843);
nor UO_820 (O_820,N_4794,N_4893);
and UO_821 (O_821,N_4705,N_4571);
nor UO_822 (O_822,N_4539,N_4640);
nand UO_823 (O_823,N_4623,N_4942);
and UO_824 (O_824,N_4521,N_4987);
xnor UO_825 (O_825,N_4619,N_4655);
nand UO_826 (O_826,N_4744,N_4606);
and UO_827 (O_827,N_4964,N_4978);
nand UO_828 (O_828,N_4611,N_4588);
and UO_829 (O_829,N_4614,N_4869);
or UO_830 (O_830,N_4930,N_4994);
xor UO_831 (O_831,N_4847,N_4616);
nand UO_832 (O_832,N_4528,N_4568);
nand UO_833 (O_833,N_4537,N_4602);
and UO_834 (O_834,N_4619,N_4770);
or UO_835 (O_835,N_4760,N_4622);
or UO_836 (O_836,N_4696,N_4942);
or UO_837 (O_837,N_4739,N_4773);
nor UO_838 (O_838,N_4856,N_4980);
nor UO_839 (O_839,N_4964,N_4725);
and UO_840 (O_840,N_4560,N_4782);
or UO_841 (O_841,N_4632,N_4911);
nand UO_842 (O_842,N_4640,N_4720);
xnor UO_843 (O_843,N_4527,N_4544);
xnor UO_844 (O_844,N_4613,N_4812);
xnor UO_845 (O_845,N_4979,N_4934);
nor UO_846 (O_846,N_4978,N_4977);
xnor UO_847 (O_847,N_4670,N_4522);
or UO_848 (O_848,N_4503,N_4537);
nor UO_849 (O_849,N_4823,N_4937);
nor UO_850 (O_850,N_4635,N_4715);
and UO_851 (O_851,N_4616,N_4830);
or UO_852 (O_852,N_4539,N_4998);
nor UO_853 (O_853,N_4831,N_4503);
or UO_854 (O_854,N_4988,N_4732);
nor UO_855 (O_855,N_4680,N_4990);
or UO_856 (O_856,N_4653,N_4850);
or UO_857 (O_857,N_4648,N_4685);
and UO_858 (O_858,N_4514,N_4697);
nand UO_859 (O_859,N_4819,N_4693);
and UO_860 (O_860,N_4525,N_4835);
xnor UO_861 (O_861,N_4617,N_4610);
and UO_862 (O_862,N_4580,N_4848);
nand UO_863 (O_863,N_4957,N_4675);
or UO_864 (O_864,N_4729,N_4595);
and UO_865 (O_865,N_4874,N_4716);
nand UO_866 (O_866,N_4673,N_4924);
or UO_867 (O_867,N_4633,N_4638);
nand UO_868 (O_868,N_4667,N_4994);
or UO_869 (O_869,N_4567,N_4610);
nor UO_870 (O_870,N_4811,N_4851);
nor UO_871 (O_871,N_4722,N_4520);
or UO_872 (O_872,N_4545,N_4820);
nor UO_873 (O_873,N_4620,N_4527);
and UO_874 (O_874,N_4851,N_4738);
nor UO_875 (O_875,N_4934,N_4745);
xnor UO_876 (O_876,N_4872,N_4815);
nor UO_877 (O_877,N_4917,N_4912);
and UO_878 (O_878,N_4845,N_4565);
and UO_879 (O_879,N_4710,N_4507);
nor UO_880 (O_880,N_4625,N_4502);
nor UO_881 (O_881,N_4930,N_4916);
and UO_882 (O_882,N_4710,N_4687);
nand UO_883 (O_883,N_4942,N_4628);
nor UO_884 (O_884,N_4604,N_4891);
and UO_885 (O_885,N_4963,N_4872);
and UO_886 (O_886,N_4624,N_4800);
and UO_887 (O_887,N_4632,N_4500);
or UO_888 (O_888,N_4684,N_4778);
nand UO_889 (O_889,N_4600,N_4888);
and UO_890 (O_890,N_4863,N_4590);
nand UO_891 (O_891,N_4784,N_4684);
and UO_892 (O_892,N_4693,N_4753);
or UO_893 (O_893,N_4847,N_4686);
nor UO_894 (O_894,N_4914,N_4934);
xor UO_895 (O_895,N_4719,N_4881);
or UO_896 (O_896,N_4632,N_4756);
nor UO_897 (O_897,N_4608,N_4927);
nand UO_898 (O_898,N_4690,N_4768);
xor UO_899 (O_899,N_4744,N_4505);
and UO_900 (O_900,N_4656,N_4696);
and UO_901 (O_901,N_4684,N_4626);
nor UO_902 (O_902,N_4931,N_4917);
nand UO_903 (O_903,N_4929,N_4939);
nor UO_904 (O_904,N_4601,N_4939);
and UO_905 (O_905,N_4697,N_4640);
and UO_906 (O_906,N_4594,N_4750);
or UO_907 (O_907,N_4845,N_4575);
nor UO_908 (O_908,N_4749,N_4502);
nand UO_909 (O_909,N_4537,N_4770);
nand UO_910 (O_910,N_4868,N_4932);
nor UO_911 (O_911,N_4500,N_4512);
and UO_912 (O_912,N_4600,N_4533);
nand UO_913 (O_913,N_4971,N_4708);
or UO_914 (O_914,N_4706,N_4974);
and UO_915 (O_915,N_4599,N_4763);
and UO_916 (O_916,N_4886,N_4808);
nand UO_917 (O_917,N_4681,N_4932);
and UO_918 (O_918,N_4850,N_4675);
or UO_919 (O_919,N_4536,N_4860);
nand UO_920 (O_920,N_4779,N_4913);
nand UO_921 (O_921,N_4617,N_4815);
nand UO_922 (O_922,N_4848,N_4896);
nand UO_923 (O_923,N_4680,N_4842);
xnor UO_924 (O_924,N_4710,N_4980);
nand UO_925 (O_925,N_4858,N_4930);
nand UO_926 (O_926,N_4615,N_4514);
nor UO_927 (O_927,N_4974,N_4720);
nor UO_928 (O_928,N_4981,N_4600);
or UO_929 (O_929,N_4747,N_4761);
nor UO_930 (O_930,N_4940,N_4969);
nand UO_931 (O_931,N_4835,N_4923);
nor UO_932 (O_932,N_4945,N_4900);
and UO_933 (O_933,N_4704,N_4630);
and UO_934 (O_934,N_4573,N_4685);
or UO_935 (O_935,N_4699,N_4798);
or UO_936 (O_936,N_4738,N_4573);
nor UO_937 (O_937,N_4888,N_4842);
nor UO_938 (O_938,N_4545,N_4597);
or UO_939 (O_939,N_4839,N_4892);
and UO_940 (O_940,N_4552,N_4779);
or UO_941 (O_941,N_4842,N_4523);
xor UO_942 (O_942,N_4518,N_4650);
or UO_943 (O_943,N_4662,N_4674);
nor UO_944 (O_944,N_4906,N_4608);
nand UO_945 (O_945,N_4708,N_4814);
and UO_946 (O_946,N_4833,N_4598);
and UO_947 (O_947,N_4941,N_4650);
nand UO_948 (O_948,N_4981,N_4675);
nor UO_949 (O_949,N_4581,N_4580);
and UO_950 (O_950,N_4794,N_4686);
nor UO_951 (O_951,N_4655,N_4932);
or UO_952 (O_952,N_4669,N_4557);
nand UO_953 (O_953,N_4606,N_4750);
xor UO_954 (O_954,N_4897,N_4524);
xor UO_955 (O_955,N_4954,N_4951);
nand UO_956 (O_956,N_4568,N_4999);
or UO_957 (O_957,N_4861,N_4683);
nand UO_958 (O_958,N_4864,N_4989);
or UO_959 (O_959,N_4635,N_4805);
nand UO_960 (O_960,N_4757,N_4534);
xnor UO_961 (O_961,N_4821,N_4547);
and UO_962 (O_962,N_4719,N_4926);
or UO_963 (O_963,N_4939,N_4546);
nand UO_964 (O_964,N_4539,N_4752);
and UO_965 (O_965,N_4970,N_4526);
or UO_966 (O_966,N_4608,N_4651);
nor UO_967 (O_967,N_4733,N_4841);
xnor UO_968 (O_968,N_4612,N_4672);
nand UO_969 (O_969,N_4841,N_4754);
nand UO_970 (O_970,N_4657,N_4788);
nor UO_971 (O_971,N_4764,N_4891);
and UO_972 (O_972,N_4887,N_4827);
nor UO_973 (O_973,N_4857,N_4729);
nor UO_974 (O_974,N_4628,N_4686);
or UO_975 (O_975,N_4847,N_4979);
nand UO_976 (O_976,N_4753,N_4624);
nor UO_977 (O_977,N_4954,N_4596);
nand UO_978 (O_978,N_4511,N_4803);
xnor UO_979 (O_979,N_4783,N_4785);
or UO_980 (O_980,N_4908,N_4992);
nor UO_981 (O_981,N_4953,N_4572);
or UO_982 (O_982,N_4816,N_4602);
nand UO_983 (O_983,N_4777,N_4982);
and UO_984 (O_984,N_4884,N_4757);
nor UO_985 (O_985,N_4553,N_4843);
xnor UO_986 (O_986,N_4961,N_4722);
nor UO_987 (O_987,N_4595,N_4709);
nor UO_988 (O_988,N_4883,N_4930);
nor UO_989 (O_989,N_4732,N_4721);
or UO_990 (O_990,N_4512,N_4710);
xnor UO_991 (O_991,N_4614,N_4860);
nand UO_992 (O_992,N_4682,N_4880);
and UO_993 (O_993,N_4847,N_4825);
nand UO_994 (O_994,N_4651,N_4655);
nor UO_995 (O_995,N_4904,N_4955);
or UO_996 (O_996,N_4755,N_4658);
xnor UO_997 (O_997,N_4956,N_4860);
nor UO_998 (O_998,N_4661,N_4809);
nand UO_999 (O_999,N_4845,N_4804);
endmodule