module basic_1500_15000_2000_10_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_223,In_1360);
nor U1 (N_1,In_238,In_147);
or U2 (N_2,In_1393,In_211);
nor U3 (N_3,In_971,In_794);
or U4 (N_4,In_578,In_1400);
nand U5 (N_5,In_881,In_67);
nor U6 (N_6,In_76,In_250);
nor U7 (N_7,In_1189,In_1415);
and U8 (N_8,In_251,In_576);
and U9 (N_9,In_1052,In_663);
and U10 (N_10,In_438,In_1064);
nor U11 (N_11,In_350,In_778);
or U12 (N_12,In_1275,In_841);
nand U13 (N_13,In_950,In_1386);
or U14 (N_14,In_697,In_98);
nor U15 (N_15,In_1298,In_1350);
and U16 (N_16,In_1412,In_1231);
nand U17 (N_17,In_749,In_1396);
nand U18 (N_18,In_534,In_1176);
or U19 (N_19,In_285,In_1286);
and U20 (N_20,In_1076,In_896);
nor U21 (N_21,In_1319,In_204);
nor U22 (N_22,In_277,In_893);
nor U23 (N_23,In_725,In_133);
nor U24 (N_24,In_1483,In_1365);
or U25 (N_25,In_956,In_1445);
nand U26 (N_26,In_1217,In_1123);
nand U27 (N_27,In_1164,In_248);
nand U28 (N_28,In_221,In_1349);
nand U29 (N_29,In_279,In_68);
nor U30 (N_30,In_1326,In_410);
nor U31 (N_31,In_430,In_474);
and U32 (N_32,In_793,In_637);
xor U33 (N_33,In_263,In_107);
xnor U34 (N_34,In_897,In_737);
and U35 (N_35,In_152,In_89);
or U36 (N_36,In_169,In_610);
and U37 (N_37,In_28,In_1495);
nand U38 (N_38,In_597,In_457);
nand U39 (N_39,In_342,In_1213);
or U40 (N_40,In_1180,In_1318);
xor U41 (N_41,In_764,In_198);
or U42 (N_42,In_641,In_115);
or U43 (N_43,In_472,In_1369);
xnor U44 (N_44,In_325,In_295);
and U45 (N_45,In_1188,In_650);
and U46 (N_46,In_236,In_1478);
and U47 (N_47,In_283,In_1424);
xnor U48 (N_48,In_293,In_414);
or U49 (N_49,In_501,In_1031);
xnor U50 (N_50,In_305,In_813);
nand U51 (N_51,In_599,In_464);
nand U52 (N_52,In_979,In_1082);
nor U53 (N_53,In_291,In_1169);
and U54 (N_54,In_520,In_1035);
nor U55 (N_55,In_196,In_174);
and U56 (N_56,In_1362,In_38);
or U57 (N_57,In_441,In_938);
and U58 (N_58,In_690,In_999);
xor U59 (N_59,In_1114,In_354);
and U60 (N_60,In_1437,In_759);
nand U61 (N_61,In_1351,In_621);
or U62 (N_62,In_815,In_1306);
or U63 (N_63,In_1142,In_1370);
and U64 (N_64,In_1055,In_570);
nand U65 (N_65,In_1156,In_1038);
nor U66 (N_66,In_747,In_985);
nor U67 (N_67,In_255,In_378);
and U68 (N_68,In_131,In_398);
xnor U69 (N_69,In_916,In_762);
xnor U70 (N_70,In_21,In_1135);
nand U71 (N_71,In_524,In_848);
and U72 (N_72,In_149,In_473);
or U73 (N_73,In_1497,In_121);
xnor U74 (N_74,In_1460,In_1472);
and U75 (N_75,In_423,In_447);
xor U76 (N_76,In_1476,In_454);
and U77 (N_77,In_1129,In_1207);
or U78 (N_78,In_1446,In_157);
xor U79 (N_79,In_178,In_240);
nor U80 (N_80,In_845,In_1468);
xnor U81 (N_81,In_924,In_1191);
nand U82 (N_82,In_275,In_862);
or U83 (N_83,In_1032,In_1270);
nor U84 (N_84,In_319,In_307);
nor U85 (N_85,In_1183,In_234);
nand U86 (N_86,In_1072,In_1153);
nand U87 (N_87,In_557,In_939);
or U88 (N_88,In_1008,In_268);
and U89 (N_89,In_646,In_45);
and U90 (N_90,In_1074,In_817);
nor U91 (N_91,In_606,In_311);
nand U92 (N_92,In_1090,In_79);
or U93 (N_93,In_321,In_542);
or U94 (N_94,In_361,In_1378);
nand U95 (N_95,In_1493,In_870);
or U96 (N_96,In_568,In_947);
nand U97 (N_97,In_303,In_19);
nand U98 (N_98,In_1131,In_537);
or U99 (N_99,In_475,In_1078);
xnor U100 (N_100,In_538,In_1414);
or U101 (N_101,In_802,In_1019);
and U102 (N_102,In_23,In_755);
and U103 (N_103,In_717,In_1485);
nand U104 (N_104,In_890,In_918);
xor U105 (N_105,In_1484,In_715);
and U106 (N_106,In_182,In_672);
or U107 (N_107,In_381,In_1068);
nor U108 (N_108,In_433,In_276);
or U109 (N_109,In_784,In_128);
and U110 (N_110,In_907,In_412);
xor U111 (N_111,In_1469,In_1436);
xor U112 (N_112,In_1372,In_510);
or U113 (N_113,In_824,In_281);
and U114 (N_114,In_1366,In_1474);
and U115 (N_115,In_1187,In_1039);
nor U116 (N_116,In_1287,In_445);
or U117 (N_117,In_865,In_587);
or U118 (N_118,In_941,In_804);
and U119 (N_119,In_609,In_18);
nand U120 (N_120,In_921,In_420);
and U121 (N_121,In_109,In_408);
or U122 (N_122,In_145,In_1455);
nand U123 (N_123,In_1274,In_83);
nand U124 (N_124,In_161,In_118);
nand U125 (N_125,In_507,In_847);
or U126 (N_126,In_614,In_108);
nand U127 (N_127,In_505,In_991);
xor U128 (N_128,In_1304,In_316);
xnor U129 (N_129,In_181,In_1079);
nor U130 (N_130,In_436,In_143);
xor U131 (N_131,In_1044,In_87);
or U132 (N_132,In_628,In_1144);
and U133 (N_133,In_852,In_1438);
xnor U134 (N_134,In_1220,In_994);
nor U135 (N_135,In_613,In_684);
xor U136 (N_136,In_839,In_403);
and U137 (N_137,In_1101,In_237);
nand U138 (N_138,In_1246,In_478);
or U139 (N_139,In_990,In_17);
nor U140 (N_140,In_1081,In_323);
nor U141 (N_141,In_7,In_590);
nand U142 (N_142,In_165,In_837);
and U143 (N_143,In_153,In_335);
nor U144 (N_144,In_232,In_1206);
and U145 (N_145,In_243,In_411);
nand U146 (N_146,In_270,In_148);
or U147 (N_147,In_1494,In_992);
nand U148 (N_148,In_910,In_935);
nand U149 (N_149,In_1075,In_1264);
or U150 (N_150,In_961,In_333);
and U151 (N_151,In_1185,In_1441);
nor U152 (N_152,In_351,In_1060);
or U153 (N_153,In_1017,In_200);
nor U154 (N_154,In_517,In_861);
xnor U155 (N_155,In_566,In_1395);
and U156 (N_156,In_915,In_675);
and U157 (N_157,In_1439,In_494);
xor U158 (N_158,In_296,In_1095);
and U159 (N_159,In_487,In_431);
nor U160 (N_160,In_928,In_544);
nor U161 (N_161,In_1151,In_241);
or U162 (N_162,In_787,In_668);
and U163 (N_163,In_953,In_1235);
xor U164 (N_164,In_129,In_170);
xnor U165 (N_165,In_721,In_96);
xnor U166 (N_166,In_1499,In_512);
nand U167 (N_167,In_1084,In_547);
xor U168 (N_168,In_693,In_77);
or U169 (N_169,In_229,In_579);
or U170 (N_170,In_56,In_1233);
nor U171 (N_171,In_1121,In_1173);
xnor U172 (N_172,In_482,In_1146);
nand U173 (N_173,In_466,In_957);
xnor U174 (N_174,In_1302,In_1300);
and U175 (N_175,In_465,In_102);
and U176 (N_176,In_620,In_369);
nor U177 (N_177,In_47,In_1087);
or U178 (N_178,In_419,In_1292);
and U179 (N_179,In_239,In_184);
and U180 (N_180,In_989,In_246);
nand U181 (N_181,In_2,In_61);
nand U182 (N_182,In_1279,In_652);
or U183 (N_183,In_415,In_533);
xnor U184 (N_184,In_1036,In_1152);
and U185 (N_185,In_643,In_1);
or U186 (N_186,In_687,In_85);
xor U187 (N_187,In_126,In_1042);
xor U188 (N_188,In_863,In_780);
nor U189 (N_189,In_514,In_429);
or U190 (N_190,In_84,In_830);
nor U191 (N_191,In_52,In_1265);
xnor U192 (N_192,In_730,In_623);
and U193 (N_193,In_1250,In_97);
and U194 (N_194,In_1015,In_888);
and U195 (N_195,In_337,In_159);
and U196 (N_196,In_1467,In_491);
nand U197 (N_197,In_160,In_691);
xnor U198 (N_198,In_1256,In_1228);
nor U199 (N_199,In_1184,In_326);
and U200 (N_200,In_826,In_965);
or U201 (N_201,In_1065,In_1389);
xnor U202 (N_202,In_653,In_689);
nor U203 (N_203,In_1284,In_1307);
nand U204 (N_204,In_545,In_488);
nor U205 (N_205,In_1174,In_1053);
nor U206 (N_206,In_1092,In_162);
xnor U207 (N_207,In_382,In_591);
nor U208 (N_208,In_1221,In_230);
and U209 (N_209,In_1239,In_288);
or U210 (N_210,In_974,In_69);
and U211 (N_211,In_130,In_55);
or U212 (N_212,In_1463,In_427);
nor U213 (N_213,In_676,In_925);
and U214 (N_214,In_976,In_1477);
and U215 (N_215,In_1148,In_806);
and U216 (N_216,In_771,In_753);
nand U217 (N_217,In_214,In_1251);
and U218 (N_218,In_699,In_387);
and U219 (N_219,In_399,In_572);
nor U220 (N_220,In_1198,In_188);
and U221 (N_221,In_1325,In_484);
or U222 (N_222,In_611,In_404);
nand U223 (N_223,In_1117,In_1259);
nor U224 (N_224,In_158,In_267);
or U225 (N_225,In_249,In_1473);
xor U226 (N_226,In_523,In_449);
nand U227 (N_227,In_919,In_1482);
nand U228 (N_228,In_605,In_338);
or U229 (N_229,In_39,In_213);
or U230 (N_230,In_1481,In_805);
xor U231 (N_231,In_1051,In_777);
nor U232 (N_232,In_1194,In_1491);
nor U233 (N_233,In_718,In_603);
xnor U234 (N_234,In_1179,In_1432);
nor U235 (N_235,In_785,In_1358);
xor U236 (N_236,In_882,In_602);
xnor U237 (N_237,In_1273,In_282);
nor U238 (N_238,In_190,In_139);
xor U239 (N_239,In_775,In_205);
xor U240 (N_240,In_177,In_710);
or U241 (N_241,In_1346,In_336);
xor U242 (N_242,In_840,In_1332);
and U243 (N_243,In_1430,In_530);
nand U244 (N_244,In_1301,In_140);
nand U245 (N_245,In_714,In_1345);
xor U246 (N_246,In_1093,In_1451);
nand U247 (N_247,In_903,In_11);
and U248 (N_248,In_511,In_318);
nand U249 (N_249,In_855,In_1263);
nor U250 (N_250,In_773,In_416);
nor U251 (N_251,In_746,In_1280);
nor U252 (N_252,In_1150,In_171);
or U253 (N_253,In_1227,In_782);
or U254 (N_254,In_20,In_801);
xor U255 (N_255,In_183,In_73);
and U256 (N_256,In_1431,In_114);
and U257 (N_257,In_203,In_1354);
and U258 (N_258,In_527,In_1058);
and U259 (N_259,In_552,In_926);
xor U260 (N_260,In_1294,In_1154);
nand U261 (N_261,In_1255,In_1442);
and U262 (N_262,In_745,In_364);
and U263 (N_263,In_1110,In_1040);
or U264 (N_264,In_439,In_1182);
and U265 (N_265,In_127,In_1067);
and U266 (N_266,In_1106,In_618);
and U267 (N_267,In_821,In_993);
and U268 (N_268,In_1492,In_1003);
xor U269 (N_269,In_360,In_1367);
nand U270 (N_270,In_792,In_908);
or U271 (N_271,In_1373,In_854);
xor U272 (N_272,In_563,In_100);
nand U273 (N_273,In_633,In_479);
or U274 (N_274,In_471,In_297);
and U275 (N_275,In_988,In_424);
nand U276 (N_276,In_53,In_1024);
nor U277 (N_277,In_744,In_1281);
nor U278 (N_278,In_498,In_62);
and U279 (N_279,In_1056,In_324);
nor U280 (N_280,In_1097,In_168);
and U281 (N_281,In_960,In_1475);
and U282 (N_282,In_1462,In_1045);
nor U283 (N_283,In_176,In_413);
and U284 (N_284,In_1104,In_972);
nand U285 (N_285,In_885,In_722);
nand U286 (N_286,In_456,In_1080);
nor U287 (N_287,In_958,In_1242);
and U288 (N_288,In_937,In_1125);
nor U289 (N_289,In_669,In_1449);
xnor U290 (N_290,In_207,In_1426);
nand U291 (N_291,In_341,In_1022);
nor U292 (N_292,In_574,In_667);
nor U293 (N_293,In_776,In_559);
nand U294 (N_294,In_320,In_592);
nor U295 (N_295,In_167,In_731);
and U296 (N_296,In_930,In_141);
or U297 (N_297,In_452,In_37);
and U298 (N_298,In_58,In_1061);
xnor U299 (N_299,In_816,In_796);
nor U300 (N_300,In_708,In_1453);
or U301 (N_301,In_1323,In_1070);
nor U302 (N_302,In_1219,In_265);
or U303 (N_303,In_942,In_1488);
nor U304 (N_304,In_173,In_1459);
nor U305 (N_305,In_1405,In_74);
and U306 (N_306,In_1212,In_70);
nor U307 (N_307,In_15,In_701);
xnor U308 (N_308,In_671,In_1407);
or U309 (N_309,In_1324,In_549);
nor U310 (N_310,In_1163,In_220);
or U311 (N_311,In_273,In_1013);
xnor U312 (N_312,In_1429,In_1200);
or U313 (N_313,In_6,In_1160);
xnor U314 (N_314,In_1138,In_16);
nor U315 (N_315,In_1433,In_720);
or U316 (N_316,In_631,In_694);
and U317 (N_317,In_674,In_1119);
nor U318 (N_318,In_1054,In_1140);
xor U319 (N_319,In_119,In_654);
xnor U320 (N_320,In_664,In_573);
xnor U321 (N_321,In_425,In_385);
or U322 (N_322,In_1359,In_460);
xor U323 (N_323,In_673,In_948);
xnor U324 (N_324,In_998,In_60);
nor U325 (N_325,In_509,In_357);
nor U326 (N_326,In_330,In_222);
nor U327 (N_327,In_407,In_1214);
or U328 (N_328,In_348,In_193);
xnor U329 (N_329,In_340,In_356);
xnor U330 (N_330,In_1375,In_851);
or U331 (N_331,In_546,In_1252);
xnor U332 (N_332,In_967,In_81);
or U333 (N_333,In_905,In_352);
or U334 (N_334,In_476,In_832);
nand U335 (N_335,In_41,In_539);
nand U336 (N_336,In_1157,In_54);
nand U337 (N_337,In_1406,In_394);
or U338 (N_338,In_1126,In_984);
nand U339 (N_339,In_331,In_1411);
xor U340 (N_340,In_789,In_634);
xnor U341 (N_341,In_651,In_540);
xnor U342 (N_342,In_662,In_310);
and U343 (N_343,In_146,In_814);
or U344 (N_344,In_940,In_274);
nor U345 (N_345,In_843,In_876);
nor U346 (N_346,In_156,In_1170);
nand U347 (N_347,In_1001,In_1112);
nand U348 (N_348,In_391,In_1371);
xor U349 (N_349,In_261,In_1293);
nor U350 (N_350,In_493,In_791);
xor U351 (N_351,In_125,In_1381);
and U352 (N_352,In_625,In_685);
nand U353 (N_353,In_943,In_883);
or U354 (N_354,In_909,In_453);
xor U355 (N_355,In_1464,In_677);
nor U356 (N_356,In_1248,In_383);
or U357 (N_357,In_808,In_1288);
xor U358 (N_358,In_828,In_818);
or U359 (N_359,In_877,In_224);
xor U360 (N_360,In_1071,In_535);
or U361 (N_361,In_878,In_1330);
xor U362 (N_362,In_418,In_313);
nand U363 (N_363,In_1425,In_1115);
xnor U364 (N_364,In_269,In_1361);
nor U365 (N_365,In_1006,In_833);
or U366 (N_366,In_911,In_900);
xor U367 (N_367,In_1376,In_1422);
or U368 (N_368,In_192,In_1254);
nor U369 (N_369,In_1315,In_1471);
nand U370 (N_370,In_1276,In_422);
nor U371 (N_371,In_554,In_660);
and U372 (N_372,In_1394,In_1109);
nor U373 (N_373,In_1269,In_43);
xor U374 (N_374,In_384,In_639);
and U375 (N_375,In_1343,In_1458);
nand U376 (N_376,In_1331,In_1454);
or U377 (N_377,In_4,In_1046);
nor U378 (N_378,In_91,In_588);
nand U379 (N_379,In_1158,In_867);
and U380 (N_380,In_1007,In_966);
or U381 (N_381,In_895,In_289);
and U382 (N_382,In_1303,In_823);
nor U383 (N_383,In_1073,In_1452);
or U384 (N_384,In_1335,In_665);
or U385 (N_385,In_1107,In_290);
or U386 (N_386,In_724,In_732);
xor U387 (N_387,In_1479,In_1137);
xor U388 (N_388,In_1247,In_345);
and U389 (N_389,In_202,In_1312);
and U390 (N_390,In_210,In_711);
xor U391 (N_391,In_1161,In_1029);
nor U392 (N_392,In_151,In_1347);
nor U393 (N_393,In_1165,In_1224);
and U394 (N_394,In_1193,In_820);
and U395 (N_395,In_51,In_280);
xnor U396 (N_396,In_894,In_1435);
nor U397 (N_397,In_795,In_750);
and U398 (N_398,In_440,In_741);
xor U399 (N_399,In_951,In_1197);
or U400 (N_400,In_1291,In_1018);
and U401 (N_401,In_103,In_949);
nor U402 (N_402,In_1149,In_287);
and U403 (N_403,In_768,In_1313);
nand U404 (N_404,In_580,In_393);
nor U405 (N_405,In_497,In_679);
and U406 (N_406,In_585,In_1145);
nand U407 (N_407,In_1226,In_349);
or U408 (N_408,In_309,In_936);
nand U409 (N_409,In_231,In_358);
nor U410 (N_410,In_34,In_215);
xor U411 (N_411,In_871,In_963);
xor U412 (N_412,In_709,In_850);
nand U413 (N_413,In_595,In_616);
or U414 (N_414,In_1218,In_260);
nand U415 (N_415,In_421,In_469);
nand U416 (N_416,In_569,In_219);
nand U417 (N_417,In_155,In_589);
xnor U418 (N_418,In_432,In_1205);
nor U419 (N_419,In_1111,In_1271);
xnor U420 (N_420,In_1010,In_1457);
nand U421 (N_421,In_1392,In_467);
xor U422 (N_422,In_395,In_739);
or U423 (N_423,In_1223,In_849);
xor U424 (N_424,In_355,In_132);
nand U425 (N_425,In_1216,In_1364);
xor U426 (N_426,In_1159,In_906);
nor U427 (N_427,In_301,In_1133);
xor U428 (N_428,In_1401,In_1278);
nor U429 (N_429,In_27,In_1262);
and U430 (N_430,In_838,In_1329);
xor U431 (N_431,In_1388,In_864);
nand U432 (N_432,In_922,In_292);
nor U433 (N_433,In_640,In_1456);
nor U434 (N_434,In_233,In_648);
or U435 (N_435,In_719,In_154);
nor U436 (N_436,In_363,In_253);
xor U437 (N_437,In_90,In_272);
xnor U438 (N_438,In_1289,In_1447);
nand U439 (N_439,In_496,In_14);
or U440 (N_440,In_1043,In_973);
nor U441 (N_441,In_1113,In_934);
nor U442 (N_442,In_1342,In_88);
nand U443 (N_443,In_627,In_532);
or U444 (N_444,In_807,In_95);
nor U445 (N_445,In_1382,In_138);
nand U446 (N_446,In_742,In_887);
nand U447 (N_447,In_1066,In_195);
or U448 (N_448,In_1423,In_201);
or U449 (N_449,In_1408,In_298);
and U450 (N_450,In_682,In_1098);
or U451 (N_451,In_1421,In_59);
or U452 (N_452,In_247,In_929);
xnor U453 (N_453,In_31,In_1127);
and U454 (N_454,In_185,In_1103);
nor U455 (N_455,In_619,In_670);
xor U456 (N_456,In_377,In_874);
nor U457 (N_457,In_46,In_1450);
xor U458 (N_458,In_1086,In_1105);
nor U459 (N_459,In_1465,In_485);
or U460 (N_460,In_1260,In_1192);
nand U461 (N_461,In_1249,In_1399);
xnor U462 (N_462,In_1186,In_33);
nor U463 (N_463,In_1320,In_733);
and U464 (N_464,In_811,In_831);
xnor U465 (N_465,In_1311,In_767);
and U466 (N_466,In_244,In_825);
xnor U467 (N_467,In_1178,In_1049);
xor U468 (N_468,In_1232,In_286);
nand U469 (N_469,In_600,In_5);
nor U470 (N_470,In_1363,In_583);
xor U471 (N_471,In_528,In_92);
and U472 (N_472,In_913,In_518);
and U473 (N_473,In_1048,In_702);
or U474 (N_474,In_144,In_1210);
nand U475 (N_475,In_561,In_705);
or U476 (N_476,In_32,In_1050);
or U477 (N_477,In_134,In_373);
or U478 (N_478,In_581,In_123);
or U479 (N_479,In_1096,In_1285);
or U480 (N_480,In_729,In_692);
or U481 (N_481,In_122,In_1005);
nand U482 (N_482,In_968,In_172);
and U483 (N_483,In_1091,In_314);
nand U484 (N_484,In_1166,In_136);
nor U485 (N_485,In_612,In_264);
or U486 (N_486,In_1083,In_1296);
nor U487 (N_487,In_1141,In_751);
or U488 (N_488,In_914,In_1403);
or U489 (N_489,In_252,In_553);
nand U490 (N_490,In_712,In_86);
nand U491 (N_491,In_740,In_401);
nand U492 (N_492,In_1384,In_106);
nand U493 (N_493,In_1241,In_803);
nor U494 (N_494,In_101,In_1317);
and U495 (N_495,In_322,In_734);
xnor U496 (N_496,In_1253,In_981);
or U497 (N_497,In_904,In_111);
xor U498 (N_498,In_359,In_284);
and U499 (N_499,In_226,In_1299);
nor U500 (N_500,In_1177,In_72);
nand U501 (N_501,In_622,In_217);
nor U502 (N_502,In_1120,In_800);
xnor U503 (N_503,In_604,In_1314);
or U504 (N_504,In_842,In_562);
and U505 (N_505,In_372,In_923);
xor U506 (N_506,In_1025,In_262);
nor U507 (N_507,In_607,In_375);
or U508 (N_508,In_308,In_1461);
and U509 (N_509,In_615,In_1327);
xor U510 (N_510,In_1374,In_209);
nor U511 (N_511,In_400,In_506);
nor U512 (N_512,In_504,In_703);
nor U513 (N_513,In_834,In_1328);
nand U514 (N_514,In_256,In_1130);
xor U515 (N_515,In_271,In_443);
nor U516 (N_516,In_728,In_1027);
xnor U517 (N_517,In_112,In_1240);
and U518 (N_518,In_376,In_327);
or U519 (N_519,In_649,In_1195);
nor U520 (N_520,In_463,In_945);
and U521 (N_521,In_586,In_1261);
xor U522 (N_522,In_666,In_529);
xor U523 (N_523,In_696,In_713);
nand U524 (N_524,In_50,In_1047);
or U525 (N_525,In_756,In_1122);
or U526 (N_526,In_1136,In_189);
xor U527 (N_527,In_872,In_658);
nor U528 (N_528,In_822,In_996);
nand U529 (N_529,In_810,In_987);
xnor U530 (N_530,In_344,In_1041);
or U531 (N_531,In_779,In_461);
nand U532 (N_532,In_1236,In_1283);
nand U533 (N_533,In_970,In_110);
or U534 (N_534,In_931,In_596);
or U535 (N_535,In_197,In_1295);
nand U536 (N_536,In_437,In_402);
or U537 (N_537,In_1147,In_716);
and U538 (N_538,In_978,In_986);
nand U539 (N_539,In_955,In_1028);
or U540 (N_540,In_790,In_707);
and U541 (N_541,In_946,In_536);
xnor U542 (N_542,In_1139,In_257);
nor U543 (N_543,In_48,In_706);
xor U544 (N_544,In_799,In_495);
xnor U545 (N_545,In_1490,In_49);
nor U546 (N_546,In_278,In_459);
or U547 (N_547,In_1379,In_827);
nor U548 (N_548,In_444,In_763);
nand U549 (N_549,In_199,In_480);
xor U550 (N_550,In_312,In_1377);
xnor U551 (N_551,In_388,In_944);
xor U552 (N_552,In_1258,In_486);
and U553 (N_553,In_695,In_788);
and U554 (N_554,In_1334,In_24);
or U555 (N_555,In_567,In_636);
or U556 (N_556,In_558,In_550);
nor U557 (N_557,In_1094,In_390);
or U558 (N_558,In_1402,In_113);
nor U559 (N_559,In_99,In_513);
nand U560 (N_560,In_142,In_334);
nor U561 (N_561,In_598,In_521);
or U562 (N_562,In_0,In_769);
nor U563 (N_563,In_477,In_22);
and U564 (N_564,In_1390,In_1202);
xnor U565 (N_565,In_856,In_809);
xor U566 (N_566,In_117,In_608);
or U567 (N_567,In_560,In_1063);
nand U568 (N_568,In_704,In_1208);
xor U569 (N_569,In_1204,In_866);
and U570 (N_570,In_392,In_635);
nor U571 (N_571,In_656,In_29);
and U572 (N_572,In_543,In_899);
or U573 (N_573,In_1222,In_245);
nor U574 (N_574,In_770,In_490);
nor U575 (N_575,In_212,In_1108);
or U576 (N_576,In_1418,In_819);
or U577 (N_577,In_1077,In_1199);
xnor U578 (N_578,In_1268,In_593);
and U579 (N_579,In_1012,In_752);
nor U580 (N_580,In_386,In_75);
xor U581 (N_581,In_451,In_175);
nand U582 (N_582,In_206,In_644);
nor U583 (N_583,In_873,In_179);
and U584 (N_584,In_371,In_332);
and U585 (N_585,In_727,In_57);
or U586 (N_586,In_450,In_1498);
xor U587 (N_587,In_299,In_500);
nand U588 (N_588,In_1444,In_626);
xnor U589 (N_589,In_1026,In_1357);
or U590 (N_590,In_8,In_765);
and U591 (N_591,In_489,In_736);
or U592 (N_592,In_455,In_347);
or U593 (N_593,In_1272,In_1201);
or U594 (N_594,In_1118,In_1244);
xnor U595 (N_595,In_1099,In_686);
nand U596 (N_596,In_389,In_164);
nor U597 (N_597,In_629,In_1059);
or U598 (N_598,In_1225,In_1416);
nor U599 (N_599,In_329,In_1181);
xnor U600 (N_600,In_370,In_869);
or U601 (N_601,In_1011,In_1383);
nor U602 (N_602,In_1132,In_1155);
and U603 (N_603,In_601,In_920);
or U604 (N_604,In_1443,In_1348);
and U605 (N_605,In_835,In_760);
and U606 (N_606,In_738,In_26);
or U607 (N_607,In_186,In_1309);
nor U608 (N_608,In_254,In_194);
xor U609 (N_609,In_362,In_1404);
and U610 (N_610,In_481,In_1355);
nand U611 (N_611,In_1440,In_617);
and U612 (N_612,In_754,In_891);
or U613 (N_613,In_1171,In_582);
or U614 (N_614,In_294,In_1229);
nor U615 (N_615,In_462,In_1338);
nand U616 (N_616,In_1167,In_632);
or U617 (N_617,In_124,In_1486);
or U618 (N_618,In_1290,In_959);
and U619 (N_619,In_645,In_397);
and U620 (N_620,In_901,In_1297);
nand U621 (N_621,In_187,In_783);
nand U622 (N_622,In_1002,In_680);
nor U623 (N_623,In_1337,In_575);
or U624 (N_624,In_975,In_1143);
xor U625 (N_625,In_1100,In_798);
xnor U626 (N_626,In_977,In_1172);
or U627 (N_627,In_225,In_1368);
xor U628 (N_628,In_483,In_889);
nand U629 (N_629,In_1196,In_698);
or U630 (N_630,In_94,In_374);
xnor U631 (N_631,In_927,In_166);
xnor U632 (N_632,In_66,In_137);
xor U633 (N_633,In_502,In_1344);
or U634 (N_634,In_10,In_1385);
nand U635 (N_635,In_1062,In_120);
and U636 (N_636,In_556,In_577);
or U637 (N_637,In_366,In_630);
xnor U638 (N_638,In_409,In_525);
nor U639 (N_639,In_1391,In_1310);
or U640 (N_640,In_836,In_380);
nand U641 (N_641,In_726,In_858);
or U642 (N_642,In_860,In_917);
nand U643 (N_643,In_700,In_208);
or U644 (N_644,In_1470,In_1336);
xor U645 (N_645,In_300,In_135);
and U646 (N_646,In_1000,In_1398);
nand U647 (N_647,In_93,In_969);
nor U648 (N_648,In_499,In_302);
or U649 (N_649,In_1496,In_1353);
xor U650 (N_650,In_1203,In_898);
or U651 (N_651,In_1237,In_63);
xnor U652 (N_652,In_515,In_242);
xor U653 (N_653,In_551,In_723);
nor U654 (N_654,In_884,In_406);
nor U655 (N_655,In_1209,In_1266);
xor U656 (N_656,In_584,In_1387);
or U657 (N_657,In_1057,In_952);
nand U658 (N_658,In_879,In_35);
and U659 (N_659,In_40,In_1245);
and U660 (N_660,In_104,In_995);
and U661 (N_661,In_519,In_548);
and U662 (N_662,In_1316,In_65);
and U663 (N_663,In_857,In_42);
nor U664 (N_664,In_315,In_748);
xor U665 (N_665,In_1321,In_428);
xor U666 (N_666,In_774,In_638);
or U667 (N_667,In_1308,In_688);
xnor U668 (N_668,In_1034,In_235);
nand U669 (N_669,In_859,In_757);
nor U670 (N_670,In_1257,In_594);
nand U671 (N_671,In_657,In_1085);
xor U672 (N_672,In_367,In_1215);
nand U673 (N_673,In_565,In_1128);
nor U674 (N_674,In_82,In_216);
nor U675 (N_675,In_353,In_1397);
and U676 (N_676,In_417,In_868);
and U677 (N_677,In_564,In_1211);
xnor U678 (N_678,In_997,In_1162);
and U679 (N_679,In_902,In_105);
nor U680 (N_680,In_78,In_25);
nand U681 (N_681,In_912,In_71);
xor U682 (N_682,In_1341,In_343);
xor U683 (N_683,In_758,In_1134);
or U684 (N_684,In_227,In_1069);
nor U685 (N_685,In_1466,In_1356);
nor U686 (N_686,In_980,In_442);
or U687 (N_687,In_470,In_80);
nor U688 (N_688,In_1023,In_1102);
nand U689 (N_689,In_541,In_1016);
or U690 (N_690,In_180,In_661);
and U691 (N_691,In_1033,In_30);
nand U692 (N_692,In_368,In_1004);
nand U693 (N_693,In_1234,In_1409);
nand U694 (N_694,In_448,In_458);
and U695 (N_695,In_9,In_516);
and U696 (N_696,In_892,In_522);
or U697 (N_697,In_735,In_844);
nand U698 (N_698,In_304,In_1243);
nand U699 (N_699,In_781,In_1420);
nand U700 (N_700,In_492,In_1448);
nor U701 (N_701,In_761,In_1277);
and U702 (N_702,In_624,In_812);
and U703 (N_703,In_3,In_1322);
nor U704 (N_704,In_571,In_743);
or U705 (N_705,In_853,In_531);
nor U706 (N_706,In_1380,In_797);
nand U707 (N_707,In_44,In_346);
xor U708 (N_708,In_786,In_766);
nand U709 (N_709,In_1175,In_1282);
nand U710 (N_710,In_36,In_1434);
nand U711 (N_711,In_266,In_886);
nor U712 (N_712,In_1305,In_875);
xor U713 (N_713,In_683,In_1088);
nand U714 (N_714,In_1037,In_1333);
or U715 (N_715,In_933,In_396);
xor U716 (N_716,In_328,In_642);
xnor U717 (N_717,In_982,In_1230);
xnor U718 (N_718,In_1190,In_932);
or U719 (N_719,In_116,In_772);
or U720 (N_720,In_964,In_1339);
and U721 (N_721,In_365,In_1340);
and U722 (N_722,In_1417,In_218);
nand U723 (N_723,In_1020,In_503);
or U724 (N_724,In_1410,In_1089);
nor U725 (N_725,In_647,In_12);
nor U726 (N_726,In_1116,In_191);
nor U727 (N_727,In_962,In_163);
and U728 (N_728,In_1489,In_1427);
nor U729 (N_729,In_259,In_339);
nor U730 (N_730,In_1428,In_468);
or U731 (N_731,In_1352,In_880);
or U732 (N_732,In_1014,In_13);
xnor U733 (N_733,In_1021,In_1168);
and U734 (N_734,In_1238,In_829);
and U735 (N_735,In_508,In_526);
or U736 (N_736,In_306,In_1487);
xnor U737 (N_737,In_150,In_446);
xnor U738 (N_738,In_435,In_228);
or U739 (N_739,In_555,In_258);
nor U740 (N_740,In_1267,In_983);
nor U741 (N_741,In_405,In_681);
or U742 (N_742,In_379,In_954);
nor U743 (N_743,In_1030,In_64);
or U744 (N_744,In_1413,In_655);
and U745 (N_745,In_1419,In_659);
nor U746 (N_746,In_1124,In_317);
or U747 (N_747,In_1009,In_678);
xor U748 (N_748,In_434,In_1480);
nand U749 (N_749,In_426,In_846);
nor U750 (N_750,In_920,In_575);
and U751 (N_751,In_692,In_686);
xnor U752 (N_752,In_257,In_336);
and U753 (N_753,In_961,In_422);
nand U754 (N_754,In_160,In_1427);
xor U755 (N_755,In_208,In_540);
or U756 (N_756,In_53,In_593);
nand U757 (N_757,In_166,In_711);
xnor U758 (N_758,In_663,In_616);
nor U759 (N_759,In_1086,In_186);
nand U760 (N_760,In_1304,In_957);
and U761 (N_761,In_217,In_826);
and U762 (N_762,In_1146,In_742);
or U763 (N_763,In_66,In_1301);
xor U764 (N_764,In_658,In_435);
or U765 (N_765,In_920,In_413);
xnor U766 (N_766,In_147,In_1128);
nor U767 (N_767,In_1294,In_341);
or U768 (N_768,In_191,In_635);
and U769 (N_769,In_358,In_1056);
nand U770 (N_770,In_1376,In_883);
or U771 (N_771,In_386,In_231);
and U772 (N_772,In_166,In_801);
nand U773 (N_773,In_1080,In_1060);
xor U774 (N_774,In_735,In_103);
nor U775 (N_775,In_747,In_1104);
xnor U776 (N_776,In_1375,In_993);
or U777 (N_777,In_867,In_777);
and U778 (N_778,In_1268,In_645);
and U779 (N_779,In_566,In_362);
nand U780 (N_780,In_658,In_553);
or U781 (N_781,In_1475,In_401);
or U782 (N_782,In_1477,In_146);
xor U783 (N_783,In_219,In_111);
or U784 (N_784,In_185,In_767);
and U785 (N_785,In_1332,In_174);
nand U786 (N_786,In_28,In_24);
or U787 (N_787,In_1026,In_374);
xnor U788 (N_788,In_864,In_1067);
or U789 (N_789,In_1095,In_835);
nor U790 (N_790,In_1192,In_1190);
nor U791 (N_791,In_683,In_576);
xor U792 (N_792,In_435,In_950);
nand U793 (N_793,In_1157,In_1201);
nand U794 (N_794,In_1404,In_302);
nor U795 (N_795,In_862,In_121);
xor U796 (N_796,In_692,In_116);
nand U797 (N_797,In_1056,In_1040);
nand U798 (N_798,In_631,In_68);
nor U799 (N_799,In_1040,In_862);
nand U800 (N_800,In_1463,In_115);
nand U801 (N_801,In_207,In_1345);
or U802 (N_802,In_256,In_1101);
and U803 (N_803,In_1141,In_386);
xor U804 (N_804,In_1092,In_1373);
nand U805 (N_805,In_1443,In_255);
and U806 (N_806,In_248,In_529);
and U807 (N_807,In_642,In_1211);
nor U808 (N_808,In_13,In_1304);
xor U809 (N_809,In_646,In_1257);
nand U810 (N_810,In_8,In_838);
nor U811 (N_811,In_176,In_969);
or U812 (N_812,In_1248,In_239);
xnor U813 (N_813,In_1365,In_150);
nand U814 (N_814,In_205,In_890);
and U815 (N_815,In_182,In_960);
or U816 (N_816,In_1139,In_630);
nand U817 (N_817,In_936,In_707);
xor U818 (N_818,In_329,In_783);
xnor U819 (N_819,In_73,In_160);
or U820 (N_820,In_729,In_1225);
xnor U821 (N_821,In_674,In_819);
nor U822 (N_822,In_1067,In_692);
nor U823 (N_823,In_1491,In_1257);
nand U824 (N_824,In_19,In_508);
nor U825 (N_825,In_1491,In_505);
nand U826 (N_826,In_950,In_631);
nor U827 (N_827,In_113,In_22);
nand U828 (N_828,In_272,In_1471);
or U829 (N_829,In_1106,In_835);
and U830 (N_830,In_770,In_321);
and U831 (N_831,In_1017,In_456);
nor U832 (N_832,In_456,In_158);
nand U833 (N_833,In_1016,In_73);
and U834 (N_834,In_94,In_424);
nor U835 (N_835,In_1301,In_34);
and U836 (N_836,In_220,In_809);
nand U837 (N_837,In_832,In_984);
and U838 (N_838,In_505,In_609);
nand U839 (N_839,In_597,In_19);
or U840 (N_840,In_1325,In_1105);
nor U841 (N_841,In_373,In_1133);
xnor U842 (N_842,In_900,In_897);
or U843 (N_843,In_763,In_1412);
xnor U844 (N_844,In_1456,In_331);
nand U845 (N_845,In_1091,In_1001);
nor U846 (N_846,In_459,In_514);
nor U847 (N_847,In_859,In_1211);
or U848 (N_848,In_275,In_159);
xnor U849 (N_849,In_101,In_351);
and U850 (N_850,In_560,In_1082);
xor U851 (N_851,In_1344,In_1321);
nand U852 (N_852,In_917,In_873);
nor U853 (N_853,In_345,In_402);
nand U854 (N_854,In_595,In_737);
nand U855 (N_855,In_743,In_937);
and U856 (N_856,In_114,In_605);
xnor U857 (N_857,In_50,In_590);
or U858 (N_858,In_777,In_66);
nor U859 (N_859,In_963,In_1187);
nor U860 (N_860,In_604,In_182);
nand U861 (N_861,In_723,In_718);
and U862 (N_862,In_913,In_1422);
xor U863 (N_863,In_958,In_473);
xnor U864 (N_864,In_1395,In_1311);
xnor U865 (N_865,In_487,In_19);
or U866 (N_866,In_1445,In_1128);
and U867 (N_867,In_846,In_449);
nand U868 (N_868,In_1097,In_175);
nor U869 (N_869,In_544,In_1231);
xor U870 (N_870,In_1209,In_1365);
or U871 (N_871,In_120,In_942);
or U872 (N_872,In_1279,In_856);
xor U873 (N_873,In_1384,In_157);
and U874 (N_874,In_1244,In_1136);
or U875 (N_875,In_1229,In_1057);
nand U876 (N_876,In_28,In_71);
or U877 (N_877,In_958,In_1469);
and U878 (N_878,In_967,In_51);
or U879 (N_879,In_856,In_747);
xnor U880 (N_880,In_1271,In_180);
xnor U881 (N_881,In_827,In_649);
xnor U882 (N_882,In_1174,In_973);
nand U883 (N_883,In_678,In_722);
xnor U884 (N_884,In_180,In_291);
nand U885 (N_885,In_1262,In_408);
and U886 (N_886,In_404,In_742);
nor U887 (N_887,In_756,In_904);
nand U888 (N_888,In_382,In_828);
xnor U889 (N_889,In_1089,In_290);
or U890 (N_890,In_445,In_523);
xnor U891 (N_891,In_350,In_979);
xnor U892 (N_892,In_1146,In_972);
and U893 (N_893,In_525,In_1273);
nor U894 (N_894,In_1355,In_1237);
and U895 (N_895,In_657,In_1351);
xor U896 (N_896,In_1055,In_396);
nor U897 (N_897,In_877,In_84);
nand U898 (N_898,In_767,In_1044);
nor U899 (N_899,In_533,In_438);
xnor U900 (N_900,In_132,In_1444);
nand U901 (N_901,In_414,In_432);
nor U902 (N_902,In_646,In_1134);
nand U903 (N_903,In_127,In_758);
xor U904 (N_904,In_323,In_855);
nand U905 (N_905,In_1001,In_1394);
or U906 (N_906,In_20,In_1103);
and U907 (N_907,In_813,In_267);
nor U908 (N_908,In_486,In_861);
nor U909 (N_909,In_196,In_938);
nor U910 (N_910,In_253,In_1476);
or U911 (N_911,In_1448,In_1072);
xor U912 (N_912,In_1152,In_1043);
nand U913 (N_913,In_128,In_769);
xnor U914 (N_914,In_217,In_527);
and U915 (N_915,In_53,In_1404);
or U916 (N_916,In_529,In_316);
nor U917 (N_917,In_449,In_1059);
nand U918 (N_918,In_1124,In_1054);
nor U919 (N_919,In_432,In_1188);
and U920 (N_920,In_319,In_600);
and U921 (N_921,In_283,In_1164);
and U922 (N_922,In_320,In_1266);
nor U923 (N_923,In_1329,In_1336);
nand U924 (N_924,In_1494,In_530);
xnor U925 (N_925,In_931,In_1363);
nor U926 (N_926,In_162,In_1041);
or U927 (N_927,In_1126,In_1454);
xnor U928 (N_928,In_268,In_486);
nand U929 (N_929,In_614,In_1470);
or U930 (N_930,In_117,In_177);
nor U931 (N_931,In_599,In_1152);
or U932 (N_932,In_835,In_809);
xnor U933 (N_933,In_609,In_773);
nor U934 (N_934,In_342,In_418);
or U935 (N_935,In_1299,In_474);
and U936 (N_936,In_1027,In_288);
or U937 (N_937,In_102,In_1389);
xnor U938 (N_938,In_1021,In_1056);
xnor U939 (N_939,In_120,In_815);
and U940 (N_940,In_1343,In_1067);
and U941 (N_941,In_1430,In_284);
or U942 (N_942,In_927,In_324);
nand U943 (N_943,In_1337,In_859);
nor U944 (N_944,In_664,In_1290);
xor U945 (N_945,In_79,In_303);
and U946 (N_946,In_871,In_1352);
nor U947 (N_947,In_304,In_252);
xnor U948 (N_948,In_44,In_981);
and U949 (N_949,In_550,In_1442);
and U950 (N_950,In_903,In_158);
xnor U951 (N_951,In_822,In_671);
xnor U952 (N_952,In_675,In_1241);
nand U953 (N_953,In_1336,In_340);
nor U954 (N_954,In_73,In_171);
and U955 (N_955,In_780,In_128);
nand U956 (N_956,In_382,In_946);
nand U957 (N_957,In_1405,In_221);
nor U958 (N_958,In_1378,In_739);
and U959 (N_959,In_501,In_126);
nor U960 (N_960,In_508,In_799);
and U961 (N_961,In_1402,In_1131);
nand U962 (N_962,In_1461,In_637);
nor U963 (N_963,In_662,In_474);
and U964 (N_964,In_142,In_600);
or U965 (N_965,In_982,In_377);
nand U966 (N_966,In_1079,In_170);
nand U967 (N_967,In_331,In_1018);
and U968 (N_968,In_371,In_28);
xor U969 (N_969,In_1465,In_947);
or U970 (N_970,In_1404,In_6);
or U971 (N_971,In_687,In_688);
nand U972 (N_972,In_917,In_1075);
or U973 (N_973,In_1371,In_1312);
and U974 (N_974,In_1464,In_33);
and U975 (N_975,In_1459,In_992);
nand U976 (N_976,In_771,In_553);
xor U977 (N_977,In_1461,In_608);
nor U978 (N_978,In_170,In_48);
nor U979 (N_979,In_933,In_104);
nor U980 (N_980,In_965,In_1044);
xnor U981 (N_981,In_1364,In_905);
nor U982 (N_982,In_1133,In_423);
nand U983 (N_983,In_425,In_979);
nand U984 (N_984,In_319,In_798);
and U985 (N_985,In_336,In_98);
xor U986 (N_986,In_1057,In_358);
and U987 (N_987,In_1078,In_972);
nor U988 (N_988,In_1464,In_665);
nor U989 (N_989,In_142,In_405);
and U990 (N_990,In_710,In_402);
or U991 (N_991,In_67,In_329);
nand U992 (N_992,In_39,In_326);
and U993 (N_993,In_193,In_389);
or U994 (N_994,In_478,In_518);
nor U995 (N_995,In_1119,In_656);
or U996 (N_996,In_13,In_1163);
nand U997 (N_997,In_128,In_655);
and U998 (N_998,In_905,In_826);
nor U999 (N_999,In_1028,In_656);
xnor U1000 (N_1000,In_725,In_1036);
and U1001 (N_1001,In_709,In_451);
or U1002 (N_1002,In_798,In_26);
and U1003 (N_1003,In_1125,In_826);
or U1004 (N_1004,In_357,In_896);
nand U1005 (N_1005,In_817,In_917);
or U1006 (N_1006,In_151,In_1202);
nor U1007 (N_1007,In_554,In_130);
or U1008 (N_1008,In_1211,In_261);
xnor U1009 (N_1009,In_1030,In_1465);
nor U1010 (N_1010,In_635,In_1111);
and U1011 (N_1011,In_315,In_1038);
or U1012 (N_1012,In_295,In_352);
xnor U1013 (N_1013,In_129,In_340);
nand U1014 (N_1014,In_1086,In_1225);
xnor U1015 (N_1015,In_422,In_737);
and U1016 (N_1016,In_1452,In_1199);
nand U1017 (N_1017,In_482,In_555);
or U1018 (N_1018,In_440,In_1246);
xnor U1019 (N_1019,In_579,In_146);
and U1020 (N_1020,In_1476,In_89);
or U1021 (N_1021,In_261,In_1030);
and U1022 (N_1022,In_10,In_1054);
and U1023 (N_1023,In_1183,In_1188);
and U1024 (N_1024,In_362,In_734);
nand U1025 (N_1025,In_754,In_818);
and U1026 (N_1026,In_957,In_1281);
nor U1027 (N_1027,In_1301,In_135);
or U1028 (N_1028,In_1422,In_213);
and U1029 (N_1029,In_607,In_1259);
nor U1030 (N_1030,In_1133,In_619);
or U1031 (N_1031,In_18,In_385);
and U1032 (N_1032,In_1398,In_1339);
xnor U1033 (N_1033,In_406,In_19);
xor U1034 (N_1034,In_585,In_316);
xor U1035 (N_1035,In_514,In_1448);
nor U1036 (N_1036,In_710,In_970);
or U1037 (N_1037,In_408,In_1099);
or U1038 (N_1038,In_973,In_703);
and U1039 (N_1039,In_288,In_276);
nor U1040 (N_1040,In_472,In_1353);
or U1041 (N_1041,In_1117,In_598);
nor U1042 (N_1042,In_448,In_581);
or U1043 (N_1043,In_153,In_406);
nor U1044 (N_1044,In_675,In_750);
nand U1045 (N_1045,In_997,In_853);
or U1046 (N_1046,In_710,In_458);
or U1047 (N_1047,In_0,In_426);
nand U1048 (N_1048,In_463,In_1398);
nor U1049 (N_1049,In_254,In_1292);
or U1050 (N_1050,In_202,In_961);
nor U1051 (N_1051,In_181,In_385);
or U1052 (N_1052,In_977,In_1498);
nor U1053 (N_1053,In_169,In_589);
xnor U1054 (N_1054,In_222,In_200);
nor U1055 (N_1055,In_91,In_902);
nor U1056 (N_1056,In_364,In_964);
xor U1057 (N_1057,In_673,In_1283);
nand U1058 (N_1058,In_994,In_716);
or U1059 (N_1059,In_1204,In_906);
or U1060 (N_1060,In_1101,In_112);
or U1061 (N_1061,In_1052,In_1497);
nand U1062 (N_1062,In_194,In_1372);
or U1063 (N_1063,In_258,In_1460);
nand U1064 (N_1064,In_362,In_424);
nand U1065 (N_1065,In_1066,In_869);
nor U1066 (N_1066,In_50,In_1368);
and U1067 (N_1067,In_786,In_1228);
or U1068 (N_1068,In_517,In_1090);
xor U1069 (N_1069,In_895,In_561);
nor U1070 (N_1070,In_1133,In_372);
nor U1071 (N_1071,In_1219,In_995);
nor U1072 (N_1072,In_995,In_201);
and U1073 (N_1073,In_484,In_278);
xnor U1074 (N_1074,In_702,In_34);
xnor U1075 (N_1075,In_1162,In_647);
and U1076 (N_1076,In_171,In_165);
and U1077 (N_1077,In_48,In_1024);
or U1078 (N_1078,In_697,In_807);
or U1079 (N_1079,In_317,In_599);
or U1080 (N_1080,In_865,In_598);
xnor U1081 (N_1081,In_957,In_618);
and U1082 (N_1082,In_805,In_644);
and U1083 (N_1083,In_117,In_713);
and U1084 (N_1084,In_844,In_581);
or U1085 (N_1085,In_554,In_552);
xnor U1086 (N_1086,In_1088,In_395);
nand U1087 (N_1087,In_1428,In_584);
nor U1088 (N_1088,In_184,In_1202);
or U1089 (N_1089,In_605,In_724);
or U1090 (N_1090,In_1225,In_386);
or U1091 (N_1091,In_1124,In_805);
nor U1092 (N_1092,In_646,In_1345);
and U1093 (N_1093,In_657,In_1459);
nand U1094 (N_1094,In_1235,In_1177);
and U1095 (N_1095,In_628,In_1254);
xnor U1096 (N_1096,In_341,In_1002);
xor U1097 (N_1097,In_218,In_376);
and U1098 (N_1098,In_515,In_598);
and U1099 (N_1099,In_781,In_637);
nand U1100 (N_1100,In_1103,In_1192);
xnor U1101 (N_1101,In_1459,In_279);
nand U1102 (N_1102,In_1128,In_829);
or U1103 (N_1103,In_87,In_725);
and U1104 (N_1104,In_326,In_1244);
and U1105 (N_1105,In_1237,In_222);
xnor U1106 (N_1106,In_333,In_479);
nand U1107 (N_1107,In_976,In_1204);
nor U1108 (N_1108,In_1452,In_1413);
or U1109 (N_1109,In_1081,In_704);
and U1110 (N_1110,In_229,In_1347);
and U1111 (N_1111,In_1122,In_1301);
or U1112 (N_1112,In_297,In_1309);
and U1113 (N_1113,In_132,In_91);
nor U1114 (N_1114,In_779,In_326);
xor U1115 (N_1115,In_610,In_1289);
nor U1116 (N_1116,In_1141,In_155);
and U1117 (N_1117,In_21,In_1047);
nor U1118 (N_1118,In_1142,In_875);
or U1119 (N_1119,In_114,In_1242);
or U1120 (N_1120,In_442,In_20);
or U1121 (N_1121,In_344,In_352);
or U1122 (N_1122,In_658,In_1464);
or U1123 (N_1123,In_841,In_1324);
nor U1124 (N_1124,In_1407,In_776);
xor U1125 (N_1125,In_1308,In_371);
xnor U1126 (N_1126,In_500,In_12);
nor U1127 (N_1127,In_440,In_283);
xor U1128 (N_1128,In_700,In_150);
nand U1129 (N_1129,In_802,In_499);
xor U1130 (N_1130,In_905,In_663);
nor U1131 (N_1131,In_866,In_1227);
xor U1132 (N_1132,In_230,In_1200);
nor U1133 (N_1133,In_1204,In_272);
xnor U1134 (N_1134,In_899,In_336);
and U1135 (N_1135,In_306,In_1405);
or U1136 (N_1136,In_1081,In_399);
nand U1137 (N_1137,In_286,In_4);
nor U1138 (N_1138,In_789,In_238);
or U1139 (N_1139,In_1222,In_9);
nor U1140 (N_1140,In_515,In_437);
or U1141 (N_1141,In_102,In_1411);
xor U1142 (N_1142,In_203,In_1109);
xor U1143 (N_1143,In_785,In_188);
nand U1144 (N_1144,In_692,In_219);
nand U1145 (N_1145,In_437,In_1115);
nor U1146 (N_1146,In_355,In_1043);
or U1147 (N_1147,In_915,In_151);
nor U1148 (N_1148,In_749,In_1107);
nor U1149 (N_1149,In_616,In_1216);
nor U1150 (N_1150,In_846,In_232);
or U1151 (N_1151,In_601,In_985);
nand U1152 (N_1152,In_927,In_1353);
or U1153 (N_1153,In_1442,In_409);
and U1154 (N_1154,In_915,In_1344);
nor U1155 (N_1155,In_1157,In_385);
or U1156 (N_1156,In_1445,In_411);
or U1157 (N_1157,In_1433,In_268);
or U1158 (N_1158,In_35,In_938);
and U1159 (N_1159,In_905,In_206);
and U1160 (N_1160,In_299,In_243);
nor U1161 (N_1161,In_1357,In_315);
xor U1162 (N_1162,In_41,In_730);
xor U1163 (N_1163,In_5,In_620);
nor U1164 (N_1164,In_998,In_847);
and U1165 (N_1165,In_220,In_337);
xor U1166 (N_1166,In_734,In_751);
or U1167 (N_1167,In_991,In_1122);
xnor U1168 (N_1168,In_1424,In_52);
xor U1169 (N_1169,In_520,In_764);
and U1170 (N_1170,In_1296,In_1012);
nand U1171 (N_1171,In_119,In_1325);
and U1172 (N_1172,In_130,In_1414);
xor U1173 (N_1173,In_176,In_403);
nor U1174 (N_1174,In_474,In_376);
nand U1175 (N_1175,In_1098,In_722);
nor U1176 (N_1176,In_1078,In_52);
and U1177 (N_1177,In_1350,In_1016);
xnor U1178 (N_1178,In_1393,In_1466);
and U1179 (N_1179,In_954,In_1348);
or U1180 (N_1180,In_464,In_1306);
xnor U1181 (N_1181,In_475,In_995);
and U1182 (N_1182,In_363,In_769);
nand U1183 (N_1183,In_766,In_1104);
xnor U1184 (N_1184,In_1448,In_698);
or U1185 (N_1185,In_1181,In_159);
xor U1186 (N_1186,In_195,In_750);
nor U1187 (N_1187,In_864,In_872);
nor U1188 (N_1188,In_1031,In_1486);
or U1189 (N_1189,In_676,In_1074);
and U1190 (N_1190,In_795,In_898);
xor U1191 (N_1191,In_1247,In_143);
nor U1192 (N_1192,In_313,In_1013);
and U1193 (N_1193,In_729,In_56);
and U1194 (N_1194,In_261,In_1263);
or U1195 (N_1195,In_484,In_705);
nor U1196 (N_1196,In_662,In_870);
or U1197 (N_1197,In_184,In_1387);
nor U1198 (N_1198,In_846,In_1422);
nor U1199 (N_1199,In_948,In_1162);
xor U1200 (N_1200,In_996,In_37);
nor U1201 (N_1201,In_1418,In_65);
or U1202 (N_1202,In_1263,In_978);
nand U1203 (N_1203,In_1177,In_60);
xor U1204 (N_1204,In_1038,In_1263);
nand U1205 (N_1205,In_1263,In_1313);
or U1206 (N_1206,In_496,In_1024);
nor U1207 (N_1207,In_1016,In_1179);
nand U1208 (N_1208,In_437,In_0);
nor U1209 (N_1209,In_1006,In_71);
nor U1210 (N_1210,In_280,In_801);
nand U1211 (N_1211,In_727,In_519);
xor U1212 (N_1212,In_192,In_157);
xor U1213 (N_1213,In_1312,In_772);
nand U1214 (N_1214,In_856,In_318);
nor U1215 (N_1215,In_1047,In_498);
and U1216 (N_1216,In_283,In_665);
nand U1217 (N_1217,In_345,In_561);
or U1218 (N_1218,In_1459,In_162);
nand U1219 (N_1219,In_222,In_264);
or U1220 (N_1220,In_1473,In_698);
xnor U1221 (N_1221,In_1432,In_498);
nor U1222 (N_1222,In_1305,In_605);
xor U1223 (N_1223,In_544,In_620);
and U1224 (N_1224,In_197,In_1104);
nand U1225 (N_1225,In_266,In_979);
nor U1226 (N_1226,In_844,In_1091);
xnor U1227 (N_1227,In_322,In_1163);
xnor U1228 (N_1228,In_389,In_444);
nor U1229 (N_1229,In_906,In_507);
nand U1230 (N_1230,In_1079,In_614);
nand U1231 (N_1231,In_852,In_1376);
xnor U1232 (N_1232,In_963,In_464);
and U1233 (N_1233,In_954,In_526);
xnor U1234 (N_1234,In_88,In_757);
or U1235 (N_1235,In_1408,In_844);
xor U1236 (N_1236,In_171,In_1216);
or U1237 (N_1237,In_348,In_924);
or U1238 (N_1238,In_1290,In_1091);
nand U1239 (N_1239,In_9,In_951);
nor U1240 (N_1240,In_536,In_110);
or U1241 (N_1241,In_1338,In_1267);
and U1242 (N_1242,In_543,In_1185);
nor U1243 (N_1243,In_782,In_1287);
nand U1244 (N_1244,In_1075,In_1291);
nand U1245 (N_1245,In_1466,In_516);
nor U1246 (N_1246,In_1237,In_682);
or U1247 (N_1247,In_1103,In_237);
nor U1248 (N_1248,In_1021,In_541);
and U1249 (N_1249,In_1159,In_440);
nand U1250 (N_1250,In_1321,In_328);
xor U1251 (N_1251,In_567,In_725);
nand U1252 (N_1252,In_310,In_601);
xor U1253 (N_1253,In_1191,In_1115);
nand U1254 (N_1254,In_1415,In_286);
nor U1255 (N_1255,In_590,In_673);
or U1256 (N_1256,In_508,In_697);
nand U1257 (N_1257,In_60,In_1458);
and U1258 (N_1258,In_93,In_1415);
or U1259 (N_1259,In_1188,In_117);
nand U1260 (N_1260,In_358,In_1472);
nor U1261 (N_1261,In_1246,In_480);
or U1262 (N_1262,In_805,In_29);
or U1263 (N_1263,In_500,In_196);
and U1264 (N_1264,In_425,In_90);
xor U1265 (N_1265,In_103,In_642);
xnor U1266 (N_1266,In_641,In_535);
nand U1267 (N_1267,In_933,In_849);
xnor U1268 (N_1268,In_1012,In_447);
nand U1269 (N_1269,In_606,In_106);
nand U1270 (N_1270,In_665,In_694);
nor U1271 (N_1271,In_134,In_1226);
nor U1272 (N_1272,In_1494,In_795);
or U1273 (N_1273,In_966,In_917);
nand U1274 (N_1274,In_1331,In_993);
nor U1275 (N_1275,In_1430,In_257);
nor U1276 (N_1276,In_1198,In_285);
xor U1277 (N_1277,In_1221,In_13);
xor U1278 (N_1278,In_1204,In_1280);
nor U1279 (N_1279,In_1300,In_227);
and U1280 (N_1280,In_698,In_55);
or U1281 (N_1281,In_868,In_1057);
and U1282 (N_1282,In_1332,In_1333);
nand U1283 (N_1283,In_1413,In_336);
or U1284 (N_1284,In_992,In_714);
xor U1285 (N_1285,In_553,In_1378);
nand U1286 (N_1286,In_201,In_1426);
and U1287 (N_1287,In_1298,In_490);
and U1288 (N_1288,In_1006,In_437);
or U1289 (N_1289,In_1291,In_563);
nand U1290 (N_1290,In_1053,In_1169);
or U1291 (N_1291,In_1338,In_1060);
or U1292 (N_1292,In_294,In_1140);
nand U1293 (N_1293,In_40,In_1067);
xnor U1294 (N_1294,In_691,In_552);
and U1295 (N_1295,In_442,In_300);
and U1296 (N_1296,In_378,In_740);
or U1297 (N_1297,In_1455,In_1192);
and U1298 (N_1298,In_1225,In_495);
nand U1299 (N_1299,In_447,In_49);
or U1300 (N_1300,In_101,In_385);
nand U1301 (N_1301,In_826,In_1020);
xnor U1302 (N_1302,In_964,In_1489);
nand U1303 (N_1303,In_255,In_428);
xnor U1304 (N_1304,In_19,In_1252);
or U1305 (N_1305,In_35,In_135);
xnor U1306 (N_1306,In_228,In_1024);
nand U1307 (N_1307,In_774,In_1058);
nor U1308 (N_1308,In_1427,In_1223);
nand U1309 (N_1309,In_683,In_185);
nand U1310 (N_1310,In_298,In_525);
and U1311 (N_1311,In_871,In_620);
nand U1312 (N_1312,In_364,In_570);
nand U1313 (N_1313,In_1030,In_1418);
nand U1314 (N_1314,In_776,In_438);
nand U1315 (N_1315,In_1022,In_1087);
or U1316 (N_1316,In_988,In_12);
or U1317 (N_1317,In_0,In_889);
nand U1318 (N_1318,In_1128,In_7);
nand U1319 (N_1319,In_215,In_60);
or U1320 (N_1320,In_1424,In_36);
nor U1321 (N_1321,In_612,In_1178);
xnor U1322 (N_1322,In_192,In_452);
xnor U1323 (N_1323,In_1116,In_1499);
nor U1324 (N_1324,In_868,In_1212);
and U1325 (N_1325,In_652,In_563);
nor U1326 (N_1326,In_465,In_74);
and U1327 (N_1327,In_50,In_547);
nand U1328 (N_1328,In_1252,In_419);
and U1329 (N_1329,In_110,In_668);
nand U1330 (N_1330,In_541,In_400);
or U1331 (N_1331,In_1146,In_961);
xnor U1332 (N_1332,In_13,In_1146);
and U1333 (N_1333,In_1058,In_269);
nor U1334 (N_1334,In_1044,In_922);
nand U1335 (N_1335,In_1327,In_1356);
xor U1336 (N_1336,In_302,In_210);
or U1337 (N_1337,In_314,In_423);
nor U1338 (N_1338,In_1421,In_1390);
or U1339 (N_1339,In_1225,In_894);
or U1340 (N_1340,In_541,In_1245);
nor U1341 (N_1341,In_1061,In_654);
nand U1342 (N_1342,In_1315,In_876);
and U1343 (N_1343,In_1368,In_943);
or U1344 (N_1344,In_81,In_800);
nor U1345 (N_1345,In_1090,In_1387);
nor U1346 (N_1346,In_100,In_116);
xor U1347 (N_1347,In_1142,In_982);
xor U1348 (N_1348,In_1404,In_951);
nor U1349 (N_1349,In_768,In_372);
and U1350 (N_1350,In_1425,In_143);
nand U1351 (N_1351,In_518,In_793);
and U1352 (N_1352,In_680,In_346);
nand U1353 (N_1353,In_208,In_44);
and U1354 (N_1354,In_309,In_1138);
nor U1355 (N_1355,In_223,In_1461);
and U1356 (N_1356,In_809,In_353);
or U1357 (N_1357,In_1390,In_487);
or U1358 (N_1358,In_72,In_336);
nand U1359 (N_1359,In_770,In_173);
nand U1360 (N_1360,In_615,In_96);
and U1361 (N_1361,In_1379,In_649);
or U1362 (N_1362,In_864,In_1158);
nand U1363 (N_1363,In_866,In_1397);
and U1364 (N_1364,In_1352,In_986);
and U1365 (N_1365,In_1002,In_100);
or U1366 (N_1366,In_850,In_284);
xnor U1367 (N_1367,In_391,In_813);
and U1368 (N_1368,In_1153,In_1434);
and U1369 (N_1369,In_1338,In_1190);
and U1370 (N_1370,In_933,In_1064);
or U1371 (N_1371,In_603,In_555);
xor U1372 (N_1372,In_238,In_1436);
nor U1373 (N_1373,In_1248,In_573);
and U1374 (N_1374,In_411,In_471);
xnor U1375 (N_1375,In_646,In_1414);
nor U1376 (N_1376,In_661,In_235);
nand U1377 (N_1377,In_1074,In_1117);
xnor U1378 (N_1378,In_1440,In_228);
nor U1379 (N_1379,In_565,In_324);
or U1380 (N_1380,In_724,In_210);
nor U1381 (N_1381,In_145,In_749);
xor U1382 (N_1382,In_93,In_838);
xnor U1383 (N_1383,In_755,In_581);
nor U1384 (N_1384,In_261,In_441);
nand U1385 (N_1385,In_511,In_959);
or U1386 (N_1386,In_114,In_512);
nor U1387 (N_1387,In_655,In_832);
nand U1388 (N_1388,In_211,In_1002);
or U1389 (N_1389,In_1478,In_767);
xor U1390 (N_1390,In_1066,In_235);
or U1391 (N_1391,In_1121,In_1463);
xnor U1392 (N_1392,In_702,In_519);
and U1393 (N_1393,In_1100,In_240);
nor U1394 (N_1394,In_481,In_1400);
and U1395 (N_1395,In_880,In_32);
nor U1396 (N_1396,In_420,In_450);
and U1397 (N_1397,In_560,In_1124);
and U1398 (N_1398,In_1487,In_704);
or U1399 (N_1399,In_32,In_464);
and U1400 (N_1400,In_990,In_874);
and U1401 (N_1401,In_543,In_1379);
xor U1402 (N_1402,In_1348,In_897);
nor U1403 (N_1403,In_772,In_722);
and U1404 (N_1404,In_1220,In_918);
or U1405 (N_1405,In_199,In_876);
and U1406 (N_1406,In_62,In_833);
nand U1407 (N_1407,In_165,In_393);
xnor U1408 (N_1408,In_1000,In_880);
or U1409 (N_1409,In_1336,In_680);
xor U1410 (N_1410,In_389,In_834);
nor U1411 (N_1411,In_1414,In_1258);
or U1412 (N_1412,In_917,In_56);
and U1413 (N_1413,In_637,In_533);
nand U1414 (N_1414,In_1456,In_470);
nand U1415 (N_1415,In_148,In_1358);
or U1416 (N_1416,In_147,In_1334);
and U1417 (N_1417,In_1253,In_446);
nand U1418 (N_1418,In_651,In_1023);
and U1419 (N_1419,In_1233,In_758);
xnor U1420 (N_1420,In_498,In_288);
nand U1421 (N_1421,In_406,In_1392);
nor U1422 (N_1422,In_1491,In_758);
or U1423 (N_1423,In_907,In_947);
or U1424 (N_1424,In_496,In_127);
and U1425 (N_1425,In_475,In_153);
and U1426 (N_1426,In_704,In_1490);
xor U1427 (N_1427,In_671,In_133);
and U1428 (N_1428,In_1370,In_383);
nor U1429 (N_1429,In_1021,In_1073);
or U1430 (N_1430,In_401,In_1183);
xor U1431 (N_1431,In_75,In_576);
xor U1432 (N_1432,In_244,In_130);
or U1433 (N_1433,In_701,In_808);
nand U1434 (N_1434,In_176,In_287);
or U1435 (N_1435,In_570,In_927);
xnor U1436 (N_1436,In_539,In_795);
xnor U1437 (N_1437,In_694,In_1086);
nor U1438 (N_1438,In_1136,In_458);
or U1439 (N_1439,In_810,In_1457);
xor U1440 (N_1440,In_1290,In_458);
and U1441 (N_1441,In_1056,In_252);
and U1442 (N_1442,In_671,In_1171);
nor U1443 (N_1443,In_784,In_1339);
and U1444 (N_1444,In_574,In_252);
nor U1445 (N_1445,In_1055,In_902);
or U1446 (N_1446,In_1307,In_914);
and U1447 (N_1447,In_1350,In_618);
nand U1448 (N_1448,In_1132,In_738);
or U1449 (N_1449,In_1430,In_36);
and U1450 (N_1450,In_220,In_1409);
or U1451 (N_1451,In_299,In_657);
xor U1452 (N_1452,In_662,In_698);
xor U1453 (N_1453,In_750,In_68);
or U1454 (N_1454,In_1248,In_1398);
and U1455 (N_1455,In_1060,In_1252);
xor U1456 (N_1456,In_966,In_449);
and U1457 (N_1457,In_329,In_1491);
xor U1458 (N_1458,In_974,In_162);
nand U1459 (N_1459,In_1468,In_87);
or U1460 (N_1460,In_964,In_846);
nand U1461 (N_1461,In_919,In_491);
nand U1462 (N_1462,In_210,In_578);
nand U1463 (N_1463,In_375,In_1359);
and U1464 (N_1464,In_887,In_516);
nor U1465 (N_1465,In_1023,In_1399);
nor U1466 (N_1466,In_938,In_1278);
or U1467 (N_1467,In_650,In_120);
xnor U1468 (N_1468,In_140,In_1297);
or U1469 (N_1469,In_419,In_388);
or U1470 (N_1470,In_435,In_1063);
nand U1471 (N_1471,In_1255,In_486);
nand U1472 (N_1472,In_522,In_1280);
nor U1473 (N_1473,In_1477,In_200);
nor U1474 (N_1474,In_496,In_426);
xor U1475 (N_1475,In_180,In_316);
and U1476 (N_1476,In_1366,In_703);
nor U1477 (N_1477,In_119,In_463);
nand U1478 (N_1478,In_1052,In_31);
nor U1479 (N_1479,In_603,In_1425);
xnor U1480 (N_1480,In_343,In_182);
or U1481 (N_1481,In_323,In_1335);
nand U1482 (N_1482,In_712,In_68);
or U1483 (N_1483,In_1084,In_210);
and U1484 (N_1484,In_686,In_964);
and U1485 (N_1485,In_1343,In_175);
nand U1486 (N_1486,In_1278,In_1321);
and U1487 (N_1487,In_36,In_667);
or U1488 (N_1488,In_1192,In_236);
nand U1489 (N_1489,In_394,In_171);
xnor U1490 (N_1490,In_527,In_549);
nor U1491 (N_1491,In_170,In_1410);
and U1492 (N_1492,In_1376,In_1131);
or U1493 (N_1493,In_1382,In_159);
xnor U1494 (N_1494,In_409,In_88);
nand U1495 (N_1495,In_1068,In_581);
xnor U1496 (N_1496,In_1281,In_1220);
xor U1497 (N_1497,In_445,In_916);
and U1498 (N_1498,In_351,In_1287);
xor U1499 (N_1499,In_161,In_52);
nand U1500 (N_1500,N_1085,N_1495);
xor U1501 (N_1501,N_427,N_1254);
or U1502 (N_1502,N_24,N_1477);
xnor U1503 (N_1503,N_1068,N_97);
nor U1504 (N_1504,N_667,N_239);
nor U1505 (N_1505,N_701,N_598);
nor U1506 (N_1506,N_356,N_259);
nor U1507 (N_1507,N_567,N_108);
or U1508 (N_1508,N_882,N_447);
or U1509 (N_1509,N_1437,N_63);
or U1510 (N_1510,N_330,N_73);
and U1511 (N_1511,N_311,N_1329);
nor U1512 (N_1512,N_1391,N_771);
or U1513 (N_1513,N_1160,N_1222);
or U1514 (N_1514,N_225,N_1136);
and U1515 (N_1515,N_1397,N_364);
nand U1516 (N_1516,N_272,N_552);
or U1517 (N_1517,N_650,N_1383);
or U1518 (N_1518,N_1053,N_1194);
or U1519 (N_1519,N_766,N_1321);
nand U1520 (N_1520,N_827,N_758);
nor U1521 (N_1521,N_959,N_873);
xnor U1522 (N_1522,N_437,N_953);
xor U1523 (N_1523,N_1025,N_997);
xor U1524 (N_1524,N_352,N_1129);
and U1525 (N_1525,N_934,N_210);
and U1526 (N_1526,N_81,N_638);
xnor U1527 (N_1527,N_512,N_1275);
and U1528 (N_1528,N_1484,N_147);
and U1529 (N_1529,N_1086,N_910);
nand U1530 (N_1530,N_819,N_1173);
nand U1531 (N_1531,N_877,N_944);
nor U1532 (N_1532,N_1171,N_991);
nand U1533 (N_1533,N_682,N_1307);
or U1534 (N_1534,N_648,N_490);
or U1535 (N_1535,N_537,N_871);
or U1536 (N_1536,N_1192,N_445);
or U1537 (N_1537,N_266,N_930);
and U1538 (N_1538,N_150,N_1335);
xnor U1539 (N_1539,N_548,N_46);
nor U1540 (N_1540,N_449,N_602);
nor U1541 (N_1541,N_212,N_1107);
or U1542 (N_1542,N_1353,N_105);
nand U1543 (N_1543,N_1088,N_419);
nand U1544 (N_1544,N_1216,N_1390);
nor U1545 (N_1545,N_608,N_1457);
nor U1546 (N_1546,N_220,N_783);
nand U1547 (N_1547,N_1236,N_207);
nor U1548 (N_1548,N_547,N_148);
or U1549 (N_1549,N_1474,N_999);
xnor U1550 (N_1550,N_1319,N_580);
xor U1551 (N_1551,N_494,N_182);
xnor U1552 (N_1552,N_1190,N_78);
or U1553 (N_1553,N_1041,N_410);
nor U1554 (N_1554,N_460,N_304);
and U1555 (N_1555,N_1165,N_965);
and U1556 (N_1556,N_666,N_1366);
and U1557 (N_1557,N_125,N_228);
and U1558 (N_1558,N_249,N_1142);
nor U1559 (N_1559,N_392,N_1073);
nor U1560 (N_1560,N_1003,N_227);
and U1561 (N_1561,N_872,N_1234);
and U1562 (N_1562,N_1151,N_36);
xnor U1563 (N_1563,N_811,N_521);
nor U1564 (N_1564,N_1035,N_735);
nor U1565 (N_1565,N_679,N_727);
and U1566 (N_1566,N_189,N_1130);
nand U1567 (N_1567,N_1471,N_647);
or U1568 (N_1568,N_564,N_80);
nor U1569 (N_1569,N_510,N_1359);
xnor U1570 (N_1570,N_625,N_469);
xnor U1571 (N_1571,N_838,N_1200);
or U1572 (N_1572,N_68,N_1111);
and U1573 (N_1573,N_1405,N_741);
or U1574 (N_1574,N_1380,N_358);
xor U1575 (N_1575,N_1435,N_990);
nand U1576 (N_1576,N_146,N_1009);
nand U1577 (N_1577,N_1418,N_870);
nor U1578 (N_1578,N_1376,N_946);
or U1579 (N_1579,N_926,N_20);
or U1580 (N_1580,N_657,N_1233);
nor U1581 (N_1581,N_372,N_145);
xnor U1582 (N_1582,N_745,N_1467);
xor U1583 (N_1583,N_628,N_699);
or U1584 (N_1584,N_982,N_874);
nand U1585 (N_1585,N_5,N_504);
nand U1586 (N_1586,N_1395,N_730);
xor U1587 (N_1587,N_1120,N_1058);
nand U1588 (N_1588,N_1400,N_893);
or U1589 (N_1589,N_457,N_376);
nor U1590 (N_1590,N_116,N_143);
and U1591 (N_1591,N_1064,N_1038);
and U1592 (N_1592,N_1269,N_1119);
nor U1593 (N_1593,N_1040,N_473);
and U1594 (N_1594,N_1270,N_1011);
or U1595 (N_1595,N_35,N_913);
xnor U1596 (N_1596,N_806,N_496);
nand U1597 (N_1597,N_1350,N_787);
and U1598 (N_1598,N_1166,N_889);
xor U1599 (N_1599,N_61,N_310);
and U1600 (N_1600,N_561,N_1159);
nand U1601 (N_1601,N_1416,N_130);
nand U1602 (N_1602,N_185,N_1488);
nor U1603 (N_1603,N_1230,N_398);
nor U1604 (N_1604,N_1274,N_579);
nor U1605 (N_1605,N_1137,N_560);
xnor U1606 (N_1606,N_917,N_1134);
nand U1607 (N_1607,N_303,N_174);
or U1608 (N_1608,N_698,N_1452);
nor U1609 (N_1609,N_949,N_956);
and U1610 (N_1610,N_428,N_726);
or U1611 (N_1611,N_129,N_1162);
xor U1612 (N_1612,N_1066,N_85);
or U1613 (N_1613,N_271,N_995);
or U1614 (N_1614,N_1407,N_1180);
nand U1615 (N_1615,N_1348,N_1339);
xor U1616 (N_1616,N_477,N_405);
nor U1617 (N_1617,N_171,N_224);
or U1618 (N_1618,N_1243,N_720);
nand U1619 (N_1619,N_115,N_293);
and U1620 (N_1620,N_86,N_403);
or U1621 (N_1621,N_576,N_362);
and U1622 (N_1622,N_850,N_732);
xor U1623 (N_1623,N_696,N_301);
xor U1624 (N_1624,N_1045,N_828);
or U1625 (N_1625,N_1049,N_743);
nand U1626 (N_1626,N_118,N_455);
and U1627 (N_1627,N_281,N_1020);
nand U1628 (N_1628,N_975,N_675);
and U1629 (N_1629,N_752,N_267);
nor U1630 (N_1630,N_961,N_760);
and U1631 (N_1631,N_686,N_695);
nor U1632 (N_1632,N_1331,N_493);
and U1633 (N_1633,N_154,N_1404);
xor U1634 (N_1634,N_1365,N_1317);
or U1635 (N_1635,N_23,N_393);
or U1636 (N_1636,N_1168,N_268);
xnor U1637 (N_1637,N_206,N_1256);
nor U1638 (N_1638,N_756,N_178);
xnor U1639 (N_1639,N_1195,N_825);
xnor U1640 (N_1640,N_160,N_141);
nor U1641 (N_1641,N_248,N_1481);
xnor U1642 (N_1642,N_746,N_313);
nand U1643 (N_1643,N_1033,N_1369);
nor U1644 (N_1644,N_1028,N_41);
or U1645 (N_1645,N_27,N_865);
and U1646 (N_1646,N_110,N_553);
or U1647 (N_1647,N_1202,N_1379);
nand U1648 (N_1648,N_1189,N_1110);
or U1649 (N_1649,N_967,N_823);
or U1650 (N_1650,N_1490,N_137);
or U1651 (N_1651,N_840,N_1204);
xor U1652 (N_1652,N_500,N_739);
nor U1653 (N_1653,N_1109,N_176);
xnor U1654 (N_1654,N_375,N_1393);
or U1655 (N_1655,N_38,N_587);
nor U1656 (N_1656,N_1394,N_1145);
or U1657 (N_1657,N_1060,N_669);
or U1658 (N_1658,N_1268,N_163);
nand U1659 (N_1659,N_593,N_968);
nand U1660 (N_1660,N_592,N_1399);
nor U1661 (N_1661,N_290,N_688);
xor U1662 (N_1662,N_253,N_350);
or U1663 (N_1663,N_438,N_19);
and U1664 (N_1664,N_585,N_801);
or U1665 (N_1665,N_422,N_1310);
and U1666 (N_1666,N_831,N_238);
nand U1667 (N_1667,N_1022,N_911);
xor U1668 (N_1668,N_1021,N_881);
or U1669 (N_1669,N_1357,N_725);
or U1670 (N_1670,N_53,N_1371);
nor U1671 (N_1671,N_621,N_4);
and U1672 (N_1672,N_334,N_1434);
or U1673 (N_1673,N_1079,N_361);
and U1674 (N_1674,N_246,N_1485);
xor U1675 (N_1675,N_192,N_309);
nor U1676 (N_1676,N_179,N_400);
xnor U1677 (N_1677,N_94,N_702);
nor U1678 (N_1678,N_66,N_918);
or U1679 (N_1679,N_1398,N_395);
or U1680 (N_1680,N_1148,N_93);
nand U1681 (N_1681,N_1402,N_514);
xor U1682 (N_1682,N_605,N_700);
nand U1683 (N_1683,N_749,N_1211);
nand U1684 (N_1684,N_1453,N_273);
or U1685 (N_1685,N_211,N_584);
and U1686 (N_1686,N_1157,N_456);
nor U1687 (N_1687,N_404,N_131);
and U1688 (N_1688,N_123,N_339);
nand U1689 (N_1689,N_1247,N_287);
nand U1690 (N_1690,N_908,N_1259);
or U1691 (N_1691,N_574,N_1266);
nand U1692 (N_1692,N_729,N_104);
xor U1693 (N_1693,N_1403,N_254);
nand U1694 (N_1694,N_941,N_1342);
and U1695 (N_1695,N_315,N_1155);
xnor U1696 (N_1696,N_784,N_1262);
nand U1697 (N_1697,N_319,N_581);
nand U1698 (N_1698,N_280,N_1141);
and U1699 (N_1699,N_938,N_651);
nor U1700 (N_1700,N_476,N_181);
nand U1701 (N_1701,N_1065,N_351);
nor U1702 (N_1702,N_627,N_1445);
nand U1703 (N_1703,N_524,N_899);
xnor U1704 (N_1704,N_717,N_216);
xor U1705 (N_1705,N_399,N_662);
nor U1706 (N_1706,N_241,N_1083);
xnor U1707 (N_1707,N_1267,N_935);
and U1708 (N_1708,N_299,N_325);
and U1709 (N_1709,N_785,N_337);
xor U1710 (N_1710,N_1007,N_486);
or U1711 (N_1711,N_55,N_1330);
and U1712 (N_1712,N_417,N_165);
xnor U1713 (N_1713,N_658,N_704);
xnor U1714 (N_1714,N_180,N_1124);
and U1715 (N_1715,N_107,N_895);
and U1716 (N_1716,N_788,N_34);
or U1717 (N_1717,N_1183,N_1448);
nor U1718 (N_1718,N_221,N_1334);
and U1719 (N_1719,N_1252,N_1214);
xor U1720 (N_1720,N_1455,N_1440);
or U1721 (N_1721,N_1279,N_541);
nor U1722 (N_1722,N_1355,N_931);
and U1723 (N_1723,N_1464,N_374);
nor U1724 (N_1724,N_1037,N_639);
or U1725 (N_1725,N_640,N_478);
and U1726 (N_1726,N_925,N_1123);
nand U1727 (N_1727,N_166,N_1298);
and U1728 (N_1728,N_236,N_1131);
nand U1729 (N_1729,N_1430,N_201);
nor U1730 (N_1730,N_942,N_1167);
and U1731 (N_1731,N_183,N_878);
and U1732 (N_1732,N_517,N_862);
and U1733 (N_1733,N_1231,N_1326);
nand U1734 (N_1734,N_962,N_157);
nor U1735 (N_1735,N_1140,N_526);
nand U1736 (N_1736,N_582,N_406);
nand U1737 (N_1737,N_12,N_571);
or U1738 (N_1738,N_1006,N_95);
nand U1739 (N_1739,N_367,N_668);
nand U1740 (N_1740,N_800,N_485);
or U1741 (N_1741,N_1095,N_1122);
xnor U1742 (N_1742,N_421,N_1218);
xnor U1743 (N_1743,N_1062,N_1483);
or U1744 (N_1744,N_134,N_1108);
nor U1745 (N_1745,N_529,N_1116);
nor U1746 (N_1746,N_891,N_62);
or U1747 (N_1747,N_1163,N_243);
nand U1748 (N_1748,N_450,N_484);
nand U1749 (N_1749,N_820,N_462);
or U1750 (N_1750,N_1177,N_533);
nand U1751 (N_1751,N_719,N_572);
xor U1752 (N_1752,N_578,N_349);
xor U1753 (N_1753,N_1302,N_413);
or U1754 (N_1754,N_296,N_412);
nor U1755 (N_1755,N_1293,N_1186);
and U1756 (N_1756,N_366,N_1206);
nand U1757 (N_1757,N_441,N_863);
and U1758 (N_1758,N_282,N_920);
nand U1759 (N_1759,N_1,N_188);
and U1760 (N_1760,N_915,N_527);
nand U1761 (N_1761,N_868,N_834);
nor U1762 (N_1762,N_195,N_1286);
and U1763 (N_1763,N_300,N_1075);
nor U1764 (N_1764,N_1055,N_1389);
nor U1765 (N_1765,N_1422,N_759);
or U1766 (N_1766,N_551,N_25);
nand U1767 (N_1767,N_340,N_847);
or U1768 (N_1768,N_158,N_109);
and U1769 (N_1769,N_1074,N_937);
nand U1770 (N_1770,N_260,N_607);
nor U1771 (N_1771,N_1087,N_14);
and U1772 (N_1772,N_21,N_467);
and U1773 (N_1773,N_794,N_316);
nor U1774 (N_1774,N_1303,N_434);
and U1775 (N_1775,N_1287,N_75);
nor U1776 (N_1776,N_379,N_416);
nand U1777 (N_1777,N_89,N_1248);
or U1778 (N_1778,N_976,N_1375);
xnor U1779 (N_1779,N_851,N_1258);
nor U1780 (N_1780,N_11,N_318);
nor U1781 (N_1781,N_520,N_452);
xor U1782 (N_1782,N_1158,N_397);
or U1783 (N_1783,N_544,N_972);
nor U1784 (N_1784,N_60,N_994);
or U1785 (N_1785,N_1069,N_275);
nand U1786 (N_1786,N_1244,N_1314);
nor U1787 (N_1787,N_278,N_7);
or U1788 (N_1788,N_988,N_693);
xor U1789 (N_1789,N_951,N_928);
xor U1790 (N_1790,N_875,N_654);
or U1791 (N_1791,N_119,N_977);
and U1792 (N_1792,N_807,N_594);
nand U1793 (N_1793,N_663,N_1426);
xor U1794 (N_1794,N_1272,N_223);
nand U1795 (N_1795,N_538,N_957);
or U1796 (N_1796,N_507,N_338);
nor U1797 (N_1797,N_151,N_54);
nand U1798 (N_1798,N_641,N_710);
xor U1799 (N_1799,N_591,N_661);
nand U1800 (N_1800,N_575,N_573);
and U1801 (N_1801,N_217,N_866);
or U1802 (N_1802,N_960,N_1260);
nand U1803 (N_1803,N_390,N_229);
nor U1804 (N_1804,N_43,N_1181);
or U1805 (N_1805,N_1364,N_1133);
nand U1806 (N_1806,N_1304,N_1029);
xnor U1807 (N_1807,N_215,N_1264);
nand U1808 (N_1808,N_389,N_17);
nor U1809 (N_1809,N_565,N_939);
nor U1810 (N_1810,N_479,N_691);
and U1811 (N_1811,N_796,N_499);
and U1812 (N_1812,N_1297,N_1301);
or U1813 (N_1813,N_1128,N_323);
xor U1814 (N_1814,N_1265,N_1325);
nand U1815 (N_1815,N_1447,N_646);
or U1816 (N_1816,N_683,N_48);
xnor U1817 (N_1817,N_1280,N_804);
or U1818 (N_1818,N_1240,N_8);
xor U1819 (N_1819,N_1188,N_444);
nand U1820 (N_1820,N_1284,N_164);
nor U1821 (N_1821,N_363,N_84);
xor U1822 (N_1822,N_630,N_114);
xnor U1823 (N_1823,N_634,N_1410);
nor U1824 (N_1824,N_1449,N_128);
nand U1825 (N_1825,N_502,N_64);
or U1826 (N_1826,N_122,N_262);
xnor U1827 (N_1827,N_1349,N_927);
xor U1828 (N_1828,N_6,N_10);
and U1829 (N_1829,N_1486,N_812);
xor U1830 (N_1830,N_1071,N_1104);
or U1831 (N_1831,N_277,N_234);
xor U1832 (N_1832,N_539,N_1150);
nand U1833 (N_1833,N_274,N_769);
nand U1834 (N_1834,N_175,N_508);
nand U1835 (N_1835,N_355,N_906);
nor U1836 (N_1836,N_1344,N_82);
xnor U1837 (N_1837,N_1493,N_1253);
xor U1838 (N_1838,N_904,N_121);
nand U1839 (N_1839,N_909,N_264);
nand U1840 (N_1840,N_1356,N_761);
nand U1841 (N_1841,N_219,N_989);
or U1842 (N_1842,N_414,N_1438);
and U1843 (N_1843,N_1185,N_849);
nor U1844 (N_1844,N_1296,N_779);
nand U1845 (N_1845,N_1276,N_1368);
xor U1846 (N_1846,N_615,N_149);
and U1847 (N_1847,N_966,N_1067);
or U1848 (N_1848,N_1146,N_633);
and U1849 (N_1849,N_563,N_841);
nand U1850 (N_1850,N_1225,N_102);
nor U1851 (N_1851,N_1179,N_770);
and U1852 (N_1852,N_933,N_609);
or U1853 (N_1853,N_1413,N_550);
xnor U1854 (N_1854,N_855,N_96);
nor U1855 (N_1855,N_136,N_844);
and U1856 (N_1856,N_907,N_1091);
and U1857 (N_1857,N_1468,N_359);
nand U1858 (N_1858,N_1249,N_112);
or U1859 (N_1859,N_173,N_543);
xor U1860 (N_1860,N_606,N_692);
or U1861 (N_1861,N_51,N_568);
or U1862 (N_1862,N_74,N_464);
nand U1863 (N_1863,N_50,N_71);
or U1864 (N_1864,N_1292,N_588);
and U1865 (N_1865,N_1299,N_394);
nor U1866 (N_1866,N_1409,N_1315);
or U1867 (N_1867,N_797,N_629);
or U1868 (N_1868,N_1460,N_624);
nor U1869 (N_1869,N_135,N_49);
or U1870 (N_1870,N_488,N_1360);
nand U1871 (N_1871,N_803,N_1005);
and U1872 (N_1872,N_1333,N_226);
or U1873 (N_1873,N_13,N_706);
nor U1874 (N_1874,N_705,N_475);
or U1875 (N_1875,N_531,N_1139);
nand U1876 (N_1876,N_678,N_570);
nor U1877 (N_1877,N_993,N_368);
and U1878 (N_1878,N_816,N_306);
nor U1879 (N_1879,N_974,N_333);
or U1880 (N_1880,N_829,N_244);
nor U1881 (N_1881,N_777,N_736);
and U1882 (N_1882,N_786,N_1217);
nor U1883 (N_1883,N_291,N_519);
xor U1884 (N_1884,N_193,N_781);
nand U1885 (N_1885,N_1324,N_365);
nor U1886 (N_1886,N_1103,N_1044);
nand U1887 (N_1887,N_83,N_1017);
xnor U1888 (N_1888,N_292,N_963);
and U1889 (N_1889,N_167,N_984);
xnor U1890 (N_1890,N_1309,N_1496);
nand U1891 (N_1891,N_747,N_952);
xor U1892 (N_1892,N_322,N_424);
or U1893 (N_1893,N_635,N_451);
or U1894 (N_1894,N_32,N_853);
xor U1895 (N_1895,N_1487,N_649);
and U1896 (N_1896,N_815,N_1036);
nor U1897 (N_1897,N_1482,N_1229);
or U1898 (N_1898,N_562,N_1050);
nor U1899 (N_1899,N_1018,N_230);
nor U1900 (N_1900,N_100,N_1092);
and U1901 (N_1901,N_1196,N_970);
or U1902 (N_1902,N_1332,N_522);
nand U1903 (N_1903,N_295,N_1323);
or U1904 (N_1904,N_222,N_1370);
nand U1905 (N_1905,N_1377,N_619);
or U1906 (N_1906,N_169,N_724);
and U1907 (N_1907,N_1327,N_768);
xor U1908 (N_1908,N_1238,N_1096);
and U1909 (N_1909,N_1221,N_1070);
nand U1910 (N_1910,N_1176,N_380);
and U1911 (N_1911,N_604,N_90);
and U1912 (N_1912,N_795,N_101);
nor U1913 (N_1913,N_612,N_525);
or U1914 (N_1914,N_832,N_643);
nor U1915 (N_1915,N_1494,N_331);
or U1916 (N_1916,N_329,N_139);
nand U1917 (N_1917,N_425,N_1205);
nor U1918 (N_1918,N_1432,N_645);
xnor U1919 (N_1919,N_709,N_324);
nor U1920 (N_1920,N_1456,N_1282);
xor U1921 (N_1921,N_1382,N_532);
or U1922 (N_1922,N_1076,N_708);
nand U1923 (N_1923,N_1191,N_284);
xor U1924 (N_1924,N_1237,N_1014);
and U1925 (N_1925,N_1425,N_664);
xor U1926 (N_1926,N_814,N_733);
nand U1927 (N_1927,N_1156,N_1089);
xor U1928 (N_1928,N_817,N_320);
and U1929 (N_1929,N_1255,N_401);
nand U1930 (N_1930,N_214,N_1472);
xnor U1931 (N_1931,N_1340,N_1198);
or U1932 (N_1932,N_213,N_1012);
and U1933 (N_1933,N_1479,N_902);
nor U1934 (N_1934,N_1093,N_255);
xor U1935 (N_1935,N_923,N_1439);
nand U1936 (N_1936,N_307,N_936);
or U1937 (N_1937,N_1209,N_799);
and U1938 (N_1938,N_270,N_1153);
xor U1939 (N_1939,N_345,N_1285);
and U1940 (N_1940,N_487,N_597);
and U1941 (N_1941,N_636,N_901);
and U1942 (N_1942,N_660,N_549);
nor U1943 (N_1943,N_716,N_1415);
nor U1944 (N_1944,N_839,N_1213);
xor U1945 (N_1945,N_1039,N_245);
nor U1946 (N_1946,N_595,N_809);
nor U1947 (N_1947,N_1476,N_391);
nor U1948 (N_1948,N_1362,N_1424);
or U1949 (N_1949,N_88,N_72);
or U1950 (N_1950,N_793,N_545);
nor U1951 (N_1951,N_559,N_30);
or U1952 (N_1952,N_892,N_737);
and U1953 (N_1953,N_203,N_1312);
or U1954 (N_1954,N_1197,N_177);
xor U1955 (N_1955,N_914,N_600);
nor U1956 (N_1956,N_1420,N_184);
nand U1957 (N_1957,N_577,N_1105);
and U1958 (N_1958,N_617,N_821);
and U1959 (N_1959,N_958,N_69);
nor U1960 (N_1960,N_481,N_1313);
xor U1961 (N_1961,N_92,N_342);
and U1962 (N_1962,N_555,N_347);
or U1963 (N_1963,N_197,N_463);
nand U1964 (N_1964,N_67,N_586);
or U1965 (N_1965,N_199,N_1212);
xor U1966 (N_1966,N_232,N_894);
or U1967 (N_1967,N_233,N_734);
xnor U1968 (N_1968,N_1419,N_388);
and U1969 (N_1969,N_1164,N_680);
xnor U1970 (N_1970,N_1271,N_858);
xnor U1971 (N_1971,N_269,N_465);
nand U1972 (N_1972,N_1143,N_16);
and U1973 (N_1973,N_656,N_87);
nor U1974 (N_1974,N_386,N_637);
and U1975 (N_1975,N_1113,N_336);
nor U1976 (N_1976,N_187,N_998);
nor U1977 (N_1977,N_900,N_314);
nor U1978 (N_1978,N_1132,N_1126);
or U1979 (N_1979,N_1421,N_681);
or U1980 (N_1980,N_106,N_369);
or U1981 (N_1981,N_156,N_3);
xnor U1982 (N_1982,N_1414,N_1351);
or U1983 (N_1983,N_1475,N_370);
and U1984 (N_1984,N_1345,N_186);
or U1985 (N_1985,N_556,N_558);
and U1986 (N_1986,N_824,N_29);
xnor U1987 (N_1987,N_1170,N_940);
or U1988 (N_1988,N_912,N_190);
and U1989 (N_1989,N_987,N_1388);
and U1990 (N_1990,N_242,N_1466);
nor U1991 (N_1991,N_1316,N_802);
and U1992 (N_1992,N_943,N_509);
or U1993 (N_1993,N_111,N_1199);
or U1994 (N_1994,N_505,N_65);
nand U1995 (N_1995,N_127,N_857);
nor U1996 (N_1996,N_436,N_343);
nand U1997 (N_1997,N_1152,N_429);
nand U1998 (N_1998,N_1227,N_289);
nand U1999 (N_1999,N_610,N_155);
nor U2000 (N_2000,N_1354,N_620);
nand U2001 (N_2001,N_665,N_1363);
and U2002 (N_2002,N_218,N_440);
xnor U2003 (N_2003,N_1463,N_470);
or U2004 (N_2004,N_929,N_945);
and U2005 (N_2005,N_924,N_1401);
xnor U2006 (N_2006,N_335,N_903);
nor U2007 (N_2007,N_91,N_1178);
or U2008 (N_2008,N_653,N_431);
xnor U2009 (N_2009,N_1015,N_905);
nand U2010 (N_2010,N_738,N_1473);
nor U2011 (N_2011,N_778,N_742);
nor U2012 (N_2012,N_2,N_1320);
or U2013 (N_2013,N_762,N_837);
xor U2014 (N_2014,N_1470,N_1373);
nand U2015 (N_2015,N_26,N_466);
and U2016 (N_2016,N_789,N_1013);
nand U2017 (N_2017,N_623,N_480);
nand U2018 (N_2018,N_140,N_1406);
nand U2019 (N_2019,N_1090,N_453);
nand U2020 (N_2020,N_459,N_540);
nor U2021 (N_2021,N_1138,N_1118);
nor U2022 (N_2022,N_0,N_332);
or U2023 (N_2023,N_1056,N_1352);
or U2024 (N_2024,N_546,N_58);
xnor U2025 (N_2025,N_671,N_518);
nand U2026 (N_2026,N_757,N_888);
and U2027 (N_2027,N_1219,N_1024);
nor U2028 (N_2028,N_867,N_744);
nor U2029 (N_2029,N_28,N_1305);
and U2030 (N_2030,N_1174,N_415);
or U2031 (N_2031,N_826,N_120);
nor U2032 (N_2032,N_382,N_305);
nand U2033 (N_2033,N_1101,N_722);
nand U2034 (N_2034,N_357,N_1207);
or U2035 (N_2035,N_842,N_1441);
xor U2036 (N_2036,N_1228,N_1378);
and U2037 (N_2037,N_99,N_1387);
nor U2038 (N_2038,N_1436,N_235);
nand U2039 (N_2039,N_302,N_644);
and U2040 (N_2040,N_1288,N_1239);
xor U2041 (N_2041,N_1061,N_981);
and U2042 (N_2042,N_328,N_344);
xor U2043 (N_2043,N_1054,N_835);
or U2044 (N_2044,N_886,N_1361);
xor U2045 (N_2045,N_1367,N_845);
or U2046 (N_2046,N_47,N_782);
nor U2047 (N_2047,N_124,N_1097);
and U2048 (N_2048,N_1281,N_1290);
and U2049 (N_2049,N_1187,N_1154);
nor U2050 (N_2050,N_198,N_1257);
xnor U2051 (N_2051,N_1346,N_138);
nand U2052 (N_2052,N_1289,N_435);
nor U2053 (N_2053,N_31,N_955);
or U2054 (N_2054,N_1497,N_1492);
xor U2055 (N_2055,N_79,N_1182);
nor U2056 (N_2056,N_1032,N_791);
or U2057 (N_2057,N_448,N_978);
xnor U2058 (N_2058,N_161,N_1004);
nor U2059 (N_2059,N_703,N_250);
and U2060 (N_2060,N_848,N_341);
nand U2061 (N_2061,N_632,N_513);
nand U2062 (N_2062,N_566,N_534);
xnor U2063 (N_2063,N_1149,N_1081);
nand U2064 (N_2064,N_986,N_430);
or U2065 (N_2065,N_1343,N_162);
and U2066 (N_2066,N_590,N_1208);
or U2067 (N_2067,N_1384,N_317);
nand U2068 (N_2068,N_1459,N_1027);
nor U2069 (N_2069,N_1019,N_1094);
and U2070 (N_2070,N_276,N_589);
nor U2071 (N_2071,N_596,N_1458);
nor U2072 (N_2072,N_1223,N_601);
and U2073 (N_2073,N_712,N_1431);
xnor U2074 (N_2074,N_200,N_715);
or U2075 (N_2075,N_18,N_659);
xnor U2076 (N_2076,N_1427,N_674);
nand U2077 (N_2077,N_780,N_1002);
nand U2078 (N_2078,N_286,N_378);
xor U2079 (N_2079,N_418,N_569);
and U2080 (N_2080,N_728,N_346);
nand U2081 (N_2081,N_501,N_247);
or U2082 (N_2082,N_15,N_884);
nor U2083 (N_2083,N_1235,N_879);
and U2084 (N_2084,N_76,N_297);
nor U2085 (N_2085,N_98,N_1428);
nor U2086 (N_2086,N_689,N_792);
or U2087 (N_2087,N_360,N_1023);
nand U2088 (N_2088,N_387,N_42);
xor U2089 (N_2089,N_257,N_1300);
nor U2090 (N_2090,N_194,N_861);
or U2091 (N_2091,N_1077,N_126);
nor U2092 (N_2092,N_1184,N_258);
nor U2093 (N_2093,N_33,N_626);
xnor U2094 (N_2094,N_774,N_642);
nand U2095 (N_2095,N_298,N_1232);
or U2096 (N_2096,N_44,N_1048);
or U2097 (N_2097,N_713,N_1454);
and U2098 (N_2098,N_979,N_535);
and U2099 (N_2099,N_694,N_1294);
nor U2100 (N_2100,N_1308,N_754);
nand U2101 (N_2101,N_377,N_869);
nor U2102 (N_2102,N_511,N_948);
nand U2103 (N_2103,N_1051,N_113);
or U2104 (N_2104,N_231,N_39);
and U2105 (N_2105,N_898,N_1386);
nor U2106 (N_2106,N_1498,N_1030);
nor U2107 (N_2107,N_461,N_1322);
nor U2108 (N_2108,N_132,N_426);
nor U2109 (N_2109,N_1220,N_1480);
nor U2110 (N_2110,N_1026,N_312);
xor U2111 (N_2111,N_1047,N_763);
nor U2112 (N_2112,N_883,N_950);
nand U2113 (N_2113,N_458,N_373);
or U2114 (N_2114,N_1311,N_498);
and U2115 (N_2115,N_808,N_880);
xnor U2116 (N_2116,N_263,N_204);
or U2117 (N_2117,N_718,N_1429);
xor U2118 (N_2118,N_1461,N_265);
nand U2119 (N_2119,N_70,N_1251);
nor U2120 (N_2120,N_1080,N_1411);
and U2121 (N_2121,N_916,N_921);
xor U2122 (N_2122,N_1125,N_836);
nand U2123 (N_2123,N_672,N_1135);
nor U2124 (N_2124,N_103,N_1381);
or U2125 (N_2125,N_483,N_618);
and U2126 (N_2126,N_1396,N_1462);
and U2127 (N_2127,N_613,N_294);
or U2128 (N_2128,N_776,N_1385);
xor U2129 (N_2129,N_983,N_1224);
nand U2130 (N_2130,N_652,N_77);
nor U2131 (N_2131,N_755,N_1193);
nand U2132 (N_2132,N_687,N_1295);
and U2133 (N_2133,N_396,N_170);
or U2134 (N_2134,N_1444,N_616);
or U2135 (N_2135,N_384,N_1278);
nor U2136 (N_2136,N_285,N_1291);
xor U2137 (N_2137,N_859,N_711);
nand U2138 (N_2138,N_153,N_1446);
or U2139 (N_2139,N_446,N_583);
nand U2140 (N_2140,N_1082,N_822);
nor U2141 (N_2141,N_790,N_1169);
and U2142 (N_2142,N_1337,N_954);
and U2143 (N_2143,N_685,N_614);
xor U2144 (N_2144,N_321,N_690);
nand U2145 (N_2145,N_772,N_1112);
nand U2146 (N_2146,N_1491,N_491);
xnor U2147 (N_2147,N_1117,N_751);
xor U2148 (N_2148,N_371,N_468);
nor U2149 (N_2149,N_622,N_208);
and U2150 (N_2150,N_753,N_256);
and U2151 (N_2151,N_1059,N_56);
xor U2152 (N_2152,N_506,N_1100);
nand U2153 (N_2153,N_773,N_1336);
xor U2154 (N_2154,N_1450,N_673);
nor U2155 (N_2155,N_1273,N_1372);
nor U2156 (N_2156,N_516,N_202);
nor U2157 (N_2157,N_1412,N_818);
nor U2158 (N_2158,N_707,N_714);
or U2159 (N_2159,N_1052,N_876);
and U2160 (N_2160,N_775,N_1241);
or U2161 (N_2161,N_843,N_676);
xnor U2162 (N_2162,N_611,N_59);
or U2163 (N_2163,N_764,N_348);
nand U2164 (N_2164,N_1442,N_523);
nand U2165 (N_2165,N_1443,N_947);
nand U2166 (N_2166,N_1099,N_495);
or U2167 (N_2167,N_932,N_57);
nand U2168 (N_2168,N_554,N_454);
and U2169 (N_2169,N_142,N_492);
nor U2170 (N_2170,N_1000,N_1283);
nand U2171 (N_2171,N_237,N_442);
xor U2172 (N_2172,N_599,N_261);
nand U2173 (N_2173,N_1057,N_381);
nand U2174 (N_2174,N_1478,N_172);
xnor U2175 (N_2175,N_283,N_798);
xor U2176 (N_2176,N_1451,N_472);
and U2177 (N_2177,N_1115,N_52);
nor U2178 (N_2178,N_697,N_117);
xnor U2179 (N_2179,N_1203,N_1226);
and U2180 (N_2180,N_196,N_1408);
xor U2181 (N_2181,N_864,N_1042);
and U2182 (N_2182,N_1078,N_964);
nand U2183 (N_2183,N_308,N_432);
or U2184 (N_2184,N_383,N_846);
nor U2185 (N_2185,N_503,N_1417);
xnor U2186 (N_2186,N_252,N_971);
and U2187 (N_2187,N_279,N_439);
xor U2188 (N_2188,N_1010,N_897);
nand U2189 (N_2189,N_1318,N_474);
and U2190 (N_2190,N_1338,N_1261);
nand U2191 (N_2191,N_1161,N_353);
or U2192 (N_2192,N_1469,N_890);
nand U2193 (N_2193,N_1341,N_765);
nor U2194 (N_2194,N_750,N_402);
nand U2195 (N_2195,N_1102,N_1201);
and U2196 (N_2196,N_326,N_251);
xor U2197 (N_2197,N_1001,N_408);
or U2198 (N_2198,N_896,N_973);
nand U2199 (N_2199,N_191,N_168);
nor U2200 (N_2200,N_1358,N_40);
nor U2201 (N_2201,N_1098,N_980);
and U2202 (N_2202,N_1306,N_471);
nor U2203 (N_2203,N_813,N_1465);
or U2204 (N_2204,N_433,N_830);
nor U2205 (N_2205,N_45,N_805);
nand U2206 (N_2206,N_9,N_1374);
or U2207 (N_2207,N_1328,N_655);
and U2208 (N_2208,N_407,N_1008);
and U2209 (N_2209,N_209,N_1277);
nor U2210 (N_2210,N_1215,N_1250);
xor U2211 (N_2211,N_670,N_1499);
and U2212 (N_2212,N_852,N_420);
and U2213 (N_2213,N_854,N_723);
nor U2214 (N_2214,N_985,N_542);
xnor U2215 (N_2215,N_1144,N_530);
and U2216 (N_2216,N_1172,N_205);
xnor U2217 (N_2217,N_767,N_919);
or U2218 (N_2218,N_810,N_1114);
or U2219 (N_2219,N_22,N_1046);
nor U2220 (N_2220,N_1084,N_603);
or U2221 (N_2221,N_833,N_133);
or U2222 (N_2222,N_1433,N_887);
nand U2223 (N_2223,N_885,N_631);
and U2224 (N_2224,N_489,N_1245);
and U2225 (N_2225,N_677,N_288);
xor U2226 (N_2226,N_856,N_536);
or U2227 (N_2227,N_860,N_1031);
nand U2228 (N_2228,N_411,N_969);
and U2229 (N_2229,N_515,N_1263);
xnor U2230 (N_2230,N_497,N_748);
and U2231 (N_2231,N_144,N_1063);
nor U2232 (N_2232,N_684,N_1043);
xor U2233 (N_2233,N_1147,N_721);
xnor U2234 (N_2234,N_996,N_327);
or U2235 (N_2235,N_1072,N_482);
xnor U2236 (N_2236,N_740,N_922);
or U2237 (N_2237,N_240,N_1034);
or U2238 (N_2238,N_1175,N_1347);
nor U2239 (N_2239,N_159,N_1106);
nand U2240 (N_2240,N_409,N_385);
nand U2241 (N_2241,N_992,N_1246);
nand U2242 (N_2242,N_528,N_443);
xnor U2243 (N_2243,N_557,N_1127);
and U2244 (N_2244,N_423,N_1489);
nor U2245 (N_2245,N_37,N_152);
and U2246 (N_2246,N_1121,N_1423);
and U2247 (N_2247,N_1016,N_1392);
or U2248 (N_2248,N_731,N_1210);
nor U2249 (N_2249,N_1242,N_354);
nor U2250 (N_2250,N_1290,N_940);
xor U2251 (N_2251,N_1468,N_1012);
or U2252 (N_2252,N_487,N_886);
xor U2253 (N_2253,N_1334,N_930);
xnor U2254 (N_2254,N_913,N_846);
and U2255 (N_2255,N_654,N_808);
xnor U2256 (N_2256,N_1321,N_347);
xnor U2257 (N_2257,N_943,N_91);
nor U2258 (N_2258,N_1323,N_659);
and U2259 (N_2259,N_610,N_1240);
and U2260 (N_2260,N_512,N_1);
nor U2261 (N_2261,N_1169,N_882);
nand U2262 (N_2262,N_1043,N_378);
or U2263 (N_2263,N_803,N_1149);
xor U2264 (N_2264,N_38,N_1404);
or U2265 (N_2265,N_1243,N_1295);
and U2266 (N_2266,N_860,N_1325);
nand U2267 (N_2267,N_1118,N_461);
and U2268 (N_2268,N_1405,N_790);
xnor U2269 (N_2269,N_537,N_335);
or U2270 (N_2270,N_949,N_1228);
and U2271 (N_2271,N_526,N_1329);
and U2272 (N_2272,N_1292,N_460);
xor U2273 (N_2273,N_991,N_1377);
xor U2274 (N_2274,N_1000,N_1334);
xor U2275 (N_2275,N_1187,N_426);
or U2276 (N_2276,N_894,N_658);
nand U2277 (N_2277,N_1430,N_676);
and U2278 (N_2278,N_322,N_1025);
and U2279 (N_2279,N_1445,N_184);
or U2280 (N_2280,N_547,N_1037);
nand U2281 (N_2281,N_91,N_117);
or U2282 (N_2282,N_127,N_1267);
or U2283 (N_2283,N_882,N_755);
and U2284 (N_2284,N_143,N_1305);
xnor U2285 (N_2285,N_22,N_1169);
nand U2286 (N_2286,N_84,N_1372);
nand U2287 (N_2287,N_503,N_338);
or U2288 (N_2288,N_1486,N_144);
and U2289 (N_2289,N_1164,N_1171);
xor U2290 (N_2290,N_1139,N_814);
nor U2291 (N_2291,N_1267,N_741);
and U2292 (N_2292,N_86,N_60);
nand U2293 (N_2293,N_483,N_1309);
or U2294 (N_2294,N_470,N_613);
nand U2295 (N_2295,N_641,N_575);
nor U2296 (N_2296,N_529,N_787);
and U2297 (N_2297,N_436,N_771);
xor U2298 (N_2298,N_287,N_1375);
nor U2299 (N_2299,N_298,N_758);
and U2300 (N_2300,N_1092,N_58);
xor U2301 (N_2301,N_477,N_728);
xnor U2302 (N_2302,N_1423,N_412);
and U2303 (N_2303,N_952,N_198);
nor U2304 (N_2304,N_1434,N_988);
or U2305 (N_2305,N_892,N_1382);
nand U2306 (N_2306,N_1066,N_686);
xor U2307 (N_2307,N_311,N_644);
and U2308 (N_2308,N_53,N_490);
xnor U2309 (N_2309,N_1241,N_1435);
or U2310 (N_2310,N_522,N_619);
and U2311 (N_2311,N_1495,N_90);
or U2312 (N_2312,N_121,N_1086);
nand U2313 (N_2313,N_621,N_1395);
nor U2314 (N_2314,N_752,N_178);
nand U2315 (N_2315,N_619,N_1301);
nor U2316 (N_2316,N_605,N_629);
nand U2317 (N_2317,N_1077,N_705);
or U2318 (N_2318,N_1163,N_1350);
or U2319 (N_2319,N_276,N_1386);
xnor U2320 (N_2320,N_1171,N_882);
xor U2321 (N_2321,N_585,N_1317);
and U2322 (N_2322,N_46,N_812);
and U2323 (N_2323,N_158,N_386);
xor U2324 (N_2324,N_1114,N_1264);
and U2325 (N_2325,N_142,N_1472);
xor U2326 (N_2326,N_584,N_138);
or U2327 (N_2327,N_1268,N_982);
and U2328 (N_2328,N_234,N_1402);
xnor U2329 (N_2329,N_97,N_67);
xor U2330 (N_2330,N_698,N_241);
or U2331 (N_2331,N_196,N_526);
or U2332 (N_2332,N_1014,N_1280);
xnor U2333 (N_2333,N_1283,N_1189);
nor U2334 (N_2334,N_198,N_1485);
nor U2335 (N_2335,N_862,N_84);
and U2336 (N_2336,N_1084,N_978);
and U2337 (N_2337,N_1043,N_1421);
and U2338 (N_2338,N_989,N_1415);
and U2339 (N_2339,N_50,N_1212);
xnor U2340 (N_2340,N_338,N_367);
nand U2341 (N_2341,N_936,N_620);
xnor U2342 (N_2342,N_366,N_1487);
or U2343 (N_2343,N_1099,N_502);
nor U2344 (N_2344,N_736,N_590);
xnor U2345 (N_2345,N_542,N_1202);
or U2346 (N_2346,N_225,N_148);
and U2347 (N_2347,N_1176,N_2);
or U2348 (N_2348,N_573,N_1194);
and U2349 (N_2349,N_509,N_575);
or U2350 (N_2350,N_1233,N_720);
and U2351 (N_2351,N_253,N_742);
or U2352 (N_2352,N_515,N_1137);
nand U2353 (N_2353,N_1234,N_951);
and U2354 (N_2354,N_1469,N_878);
nor U2355 (N_2355,N_460,N_216);
xnor U2356 (N_2356,N_623,N_335);
nor U2357 (N_2357,N_679,N_180);
or U2358 (N_2358,N_195,N_402);
or U2359 (N_2359,N_1445,N_992);
and U2360 (N_2360,N_409,N_1469);
xnor U2361 (N_2361,N_209,N_122);
or U2362 (N_2362,N_956,N_998);
nand U2363 (N_2363,N_219,N_582);
xnor U2364 (N_2364,N_1025,N_544);
and U2365 (N_2365,N_995,N_1478);
nor U2366 (N_2366,N_214,N_811);
xor U2367 (N_2367,N_1348,N_429);
nor U2368 (N_2368,N_1400,N_494);
nand U2369 (N_2369,N_1086,N_260);
or U2370 (N_2370,N_560,N_1410);
and U2371 (N_2371,N_1436,N_1386);
nor U2372 (N_2372,N_179,N_1088);
or U2373 (N_2373,N_1019,N_462);
nor U2374 (N_2374,N_1412,N_1246);
nand U2375 (N_2375,N_798,N_1377);
nor U2376 (N_2376,N_971,N_1170);
nor U2377 (N_2377,N_1482,N_1041);
xnor U2378 (N_2378,N_667,N_400);
xor U2379 (N_2379,N_1006,N_225);
and U2380 (N_2380,N_323,N_576);
nand U2381 (N_2381,N_1325,N_467);
xor U2382 (N_2382,N_1365,N_88);
and U2383 (N_2383,N_1306,N_453);
nor U2384 (N_2384,N_866,N_1438);
xnor U2385 (N_2385,N_307,N_810);
or U2386 (N_2386,N_1069,N_404);
nor U2387 (N_2387,N_1239,N_126);
nand U2388 (N_2388,N_1221,N_872);
nor U2389 (N_2389,N_905,N_6);
xnor U2390 (N_2390,N_1035,N_312);
and U2391 (N_2391,N_242,N_1451);
nor U2392 (N_2392,N_1404,N_1428);
nor U2393 (N_2393,N_1392,N_138);
or U2394 (N_2394,N_840,N_461);
xnor U2395 (N_2395,N_757,N_738);
nand U2396 (N_2396,N_483,N_706);
or U2397 (N_2397,N_882,N_186);
xnor U2398 (N_2398,N_784,N_230);
nand U2399 (N_2399,N_836,N_1143);
or U2400 (N_2400,N_521,N_1051);
and U2401 (N_2401,N_341,N_273);
nor U2402 (N_2402,N_1171,N_1374);
and U2403 (N_2403,N_163,N_1136);
or U2404 (N_2404,N_612,N_577);
nand U2405 (N_2405,N_397,N_560);
xnor U2406 (N_2406,N_1441,N_445);
and U2407 (N_2407,N_1471,N_883);
and U2408 (N_2408,N_651,N_1321);
and U2409 (N_2409,N_35,N_1430);
nand U2410 (N_2410,N_1258,N_1144);
and U2411 (N_2411,N_664,N_699);
xor U2412 (N_2412,N_31,N_288);
nand U2413 (N_2413,N_1291,N_1181);
nand U2414 (N_2414,N_603,N_1063);
and U2415 (N_2415,N_968,N_913);
nor U2416 (N_2416,N_751,N_634);
xnor U2417 (N_2417,N_56,N_797);
nand U2418 (N_2418,N_1022,N_545);
nor U2419 (N_2419,N_274,N_1387);
nand U2420 (N_2420,N_906,N_291);
and U2421 (N_2421,N_1386,N_451);
nand U2422 (N_2422,N_383,N_454);
nand U2423 (N_2423,N_589,N_973);
or U2424 (N_2424,N_529,N_289);
and U2425 (N_2425,N_73,N_1146);
or U2426 (N_2426,N_768,N_787);
nand U2427 (N_2427,N_1083,N_1097);
nand U2428 (N_2428,N_815,N_1352);
xor U2429 (N_2429,N_326,N_864);
nand U2430 (N_2430,N_990,N_1254);
or U2431 (N_2431,N_876,N_222);
nor U2432 (N_2432,N_664,N_802);
nand U2433 (N_2433,N_313,N_923);
or U2434 (N_2434,N_739,N_650);
or U2435 (N_2435,N_1009,N_1212);
and U2436 (N_2436,N_167,N_1201);
or U2437 (N_2437,N_242,N_534);
or U2438 (N_2438,N_44,N_1302);
xnor U2439 (N_2439,N_700,N_1083);
nand U2440 (N_2440,N_295,N_1443);
xor U2441 (N_2441,N_1382,N_1234);
nand U2442 (N_2442,N_461,N_1425);
xnor U2443 (N_2443,N_1294,N_663);
nor U2444 (N_2444,N_312,N_507);
or U2445 (N_2445,N_175,N_1274);
nor U2446 (N_2446,N_697,N_57);
xor U2447 (N_2447,N_766,N_116);
and U2448 (N_2448,N_1119,N_86);
xnor U2449 (N_2449,N_804,N_1461);
xor U2450 (N_2450,N_973,N_1118);
xnor U2451 (N_2451,N_612,N_629);
nor U2452 (N_2452,N_1074,N_1432);
and U2453 (N_2453,N_1356,N_385);
nor U2454 (N_2454,N_922,N_916);
xnor U2455 (N_2455,N_1301,N_443);
xor U2456 (N_2456,N_458,N_762);
or U2457 (N_2457,N_306,N_526);
nand U2458 (N_2458,N_1372,N_1018);
nor U2459 (N_2459,N_340,N_859);
and U2460 (N_2460,N_1119,N_685);
or U2461 (N_2461,N_95,N_250);
or U2462 (N_2462,N_744,N_1203);
or U2463 (N_2463,N_844,N_2);
nor U2464 (N_2464,N_486,N_72);
nor U2465 (N_2465,N_743,N_945);
or U2466 (N_2466,N_819,N_938);
xnor U2467 (N_2467,N_1263,N_134);
and U2468 (N_2468,N_112,N_1074);
nand U2469 (N_2469,N_418,N_1382);
nand U2470 (N_2470,N_855,N_1152);
xor U2471 (N_2471,N_1295,N_795);
xnor U2472 (N_2472,N_925,N_1126);
or U2473 (N_2473,N_1305,N_60);
xnor U2474 (N_2474,N_531,N_189);
xnor U2475 (N_2475,N_409,N_1035);
xor U2476 (N_2476,N_1445,N_856);
or U2477 (N_2477,N_1171,N_357);
xnor U2478 (N_2478,N_612,N_492);
nand U2479 (N_2479,N_1068,N_815);
xor U2480 (N_2480,N_208,N_363);
xnor U2481 (N_2481,N_1176,N_439);
xor U2482 (N_2482,N_992,N_490);
xor U2483 (N_2483,N_1152,N_1239);
nand U2484 (N_2484,N_767,N_619);
nand U2485 (N_2485,N_556,N_1479);
nor U2486 (N_2486,N_1063,N_527);
or U2487 (N_2487,N_1372,N_1062);
and U2488 (N_2488,N_612,N_751);
nor U2489 (N_2489,N_606,N_661);
or U2490 (N_2490,N_59,N_1366);
nand U2491 (N_2491,N_45,N_19);
and U2492 (N_2492,N_590,N_388);
and U2493 (N_2493,N_106,N_28);
and U2494 (N_2494,N_1069,N_623);
nand U2495 (N_2495,N_603,N_1341);
nand U2496 (N_2496,N_1316,N_534);
nor U2497 (N_2497,N_715,N_794);
and U2498 (N_2498,N_1313,N_1363);
and U2499 (N_2499,N_396,N_1125);
nor U2500 (N_2500,N_29,N_624);
nand U2501 (N_2501,N_1042,N_710);
or U2502 (N_2502,N_1279,N_760);
nand U2503 (N_2503,N_321,N_425);
or U2504 (N_2504,N_957,N_1008);
or U2505 (N_2505,N_182,N_1107);
xnor U2506 (N_2506,N_0,N_508);
xnor U2507 (N_2507,N_1070,N_1271);
and U2508 (N_2508,N_552,N_1420);
and U2509 (N_2509,N_583,N_1041);
xnor U2510 (N_2510,N_1408,N_1017);
and U2511 (N_2511,N_1178,N_1363);
nor U2512 (N_2512,N_1358,N_1310);
xor U2513 (N_2513,N_948,N_193);
nor U2514 (N_2514,N_556,N_318);
nor U2515 (N_2515,N_852,N_1200);
and U2516 (N_2516,N_1481,N_614);
or U2517 (N_2517,N_150,N_381);
nand U2518 (N_2518,N_403,N_983);
nor U2519 (N_2519,N_1404,N_1093);
nor U2520 (N_2520,N_1332,N_808);
nor U2521 (N_2521,N_971,N_344);
nor U2522 (N_2522,N_1140,N_685);
and U2523 (N_2523,N_874,N_606);
xnor U2524 (N_2524,N_1151,N_1222);
and U2525 (N_2525,N_598,N_792);
nand U2526 (N_2526,N_1397,N_830);
xnor U2527 (N_2527,N_190,N_149);
and U2528 (N_2528,N_196,N_1458);
nor U2529 (N_2529,N_1008,N_685);
nor U2530 (N_2530,N_580,N_317);
nor U2531 (N_2531,N_694,N_677);
xnor U2532 (N_2532,N_930,N_717);
or U2533 (N_2533,N_1015,N_805);
xnor U2534 (N_2534,N_1282,N_1296);
or U2535 (N_2535,N_395,N_1145);
nand U2536 (N_2536,N_1017,N_517);
or U2537 (N_2537,N_1403,N_321);
or U2538 (N_2538,N_1315,N_199);
and U2539 (N_2539,N_952,N_1147);
or U2540 (N_2540,N_230,N_675);
nand U2541 (N_2541,N_293,N_211);
xor U2542 (N_2542,N_1114,N_920);
xor U2543 (N_2543,N_1427,N_742);
and U2544 (N_2544,N_1051,N_640);
or U2545 (N_2545,N_923,N_1380);
xnor U2546 (N_2546,N_1050,N_492);
and U2547 (N_2547,N_781,N_576);
xor U2548 (N_2548,N_205,N_187);
nor U2549 (N_2549,N_182,N_226);
nor U2550 (N_2550,N_463,N_816);
or U2551 (N_2551,N_1277,N_1030);
xnor U2552 (N_2552,N_731,N_1118);
xnor U2553 (N_2553,N_280,N_25);
or U2554 (N_2554,N_1122,N_31);
nor U2555 (N_2555,N_7,N_545);
xor U2556 (N_2556,N_251,N_1120);
nand U2557 (N_2557,N_1016,N_1096);
xor U2558 (N_2558,N_1104,N_729);
nor U2559 (N_2559,N_904,N_420);
nand U2560 (N_2560,N_1206,N_755);
nand U2561 (N_2561,N_668,N_393);
and U2562 (N_2562,N_1215,N_301);
or U2563 (N_2563,N_152,N_1035);
or U2564 (N_2564,N_661,N_12);
nand U2565 (N_2565,N_1114,N_821);
and U2566 (N_2566,N_1197,N_767);
xnor U2567 (N_2567,N_1088,N_1171);
xnor U2568 (N_2568,N_764,N_463);
or U2569 (N_2569,N_1133,N_1023);
nor U2570 (N_2570,N_1291,N_214);
nor U2571 (N_2571,N_944,N_1268);
nand U2572 (N_2572,N_1427,N_159);
xnor U2573 (N_2573,N_312,N_431);
and U2574 (N_2574,N_641,N_596);
or U2575 (N_2575,N_650,N_766);
xor U2576 (N_2576,N_157,N_975);
and U2577 (N_2577,N_690,N_590);
and U2578 (N_2578,N_157,N_1184);
nand U2579 (N_2579,N_653,N_815);
nand U2580 (N_2580,N_1131,N_1170);
and U2581 (N_2581,N_105,N_236);
or U2582 (N_2582,N_53,N_454);
and U2583 (N_2583,N_1159,N_1180);
nand U2584 (N_2584,N_1465,N_1182);
or U2585 (N_2585,N_1156,N_816);
nand U2586 (N_2586,N_828,N_1108);
and U2587 (N_2587,N_120,N_722);
nand U2588 (N_2588,N_545,N_1366);
xor U2589 (N_2589,N_428,N_826);
nand U2590 (N_2590,N_989,N_1239);
and U2591 (N_2591,N_511,N_916);
or U2592 (N_2592,N_572,N_1466);
and U2593 (N_2593,N_873,N_259);
nand U2594 (N_2594,N_1099,N_1125);
or U2595 (N_2595,N_279,N_77);
or U2596 (N_2596,N_312,N_166);
xnor U2597 (N_2597,N_42,N_601);
nand U2598 (N_2598,N_489,N_1304);
nand U2599 (N_2599,N_45,N_945);
or U2600 (N_2600,N_372,N_1235);
nor U2601 (N_2601,N_731,N_497);
or U2602 (N_2602,N_356,N_1028);
xor U2603 (N_2603,N_888,N_909);
and U2604 (N_2604,N_963,N_1194);
xnor U2605 (N_2605,N_339,N_1163);
and U2606 (N_2606,N_874,N_1078);
and U2607 (N_2607,N_1494,N_643);
and U2608 (N_2608,N_61,N_104);
xor U2609 (N_2609,N_725,N_615);
or U2610 (N_2610,N_1167,N_1277);
xnor U2611 (N_2611,N_125,N_1086);
xor U2612 (N_2612,N_819,N_114);
xnor U2613 (N_2613,N_1159,N_540);
nor U2614 (N_2614,N_119,N_881);
nor U2615 (N_2615,N_1206,N_1127);
and U2616 (N_2616,N_668,N_120);
nand U2617 (N_2617,N_360,N_1405);
nor U2618 (N_2618,N_822,N_559);
nand U2619 (N_2619,N_960,N_183);
nand U2620 (N_2620,N_140,N_497);
xnor U2621 (N_2621,N_1242,N_1354);
xor U2622 (N_2622,N_311,N_954);
xnor U2623 (N_2623,N_411,N_721);
nand U2624 (N_2624,N_140,N_1160);
nand U2625 (N_2625,N_833,N_516);
nand U2626 (N_2626,N_361,N_444);
nand U2627 (N_2627,N_1020,N_1107);
nor U2628 (N_2628,N_141,N_28);
or U2629 (N_2629,N_1103,N_1417);
and U2630 (N_2630,N_730,N_363);
xnor U2631 (N_2631,N_333,N_1456);
or U2632 (N_2632,N_1035,N_160);
and U2633 (N_2633,N_1047,N_1496);
or U2634 (N_2634,N_1366,N_1244);
and U2635 (N_2635,N_89,N_394);
and U2636 (N_2636,N_1456,N_296);
nand U2637 (N_2637,N_559,N_498);
xnor U2638 (N_2638,N_800,N_687);
or U2639 (N_2639,N_1226,N_514);
xor U2640 (N_2640,N_146,N_644);
and U2641 (N_2641,N_989,N_1193);
xnor U2642 (N_2642,N_970,N_438);
xnor U2643 (N_2643,N_210,N_1244);
or U2644 (N_2644,N_711,N_47);
nand U2645 (N_2645,N_885,N_514);
or U2646 (N_2646,N_38,N_174);
nand U2647 (N_2647,N_116,N_719);
or U2648 (N_2648,N_1228,N_80);
xnor U2649 (N_2649,N_435,N_101);
xnor U2650 (N_2650,N_821,N_401);
nor U2651 (N_2651,N_1463,N_79);
nor U2652 (N_2652,N_200,N_1462);
or U2653 (N_2653,N_1399,N_249);
nand U2654 (N_2654,N_966,N_1083);
nor U2655 (N_2655,N_1380,N_383);
nor U2656 (N_2656,N_49,N_1421);
nor U2657 (N_2657,N_1345,N_1312);
nand U2658 (N_2658,N_1240,N_634);
nor U2659 (N_2659,N_1205,N_698);
and U2660 (N_2660,N_791,N_1221);
xnor U2661 (N_2661,N_1166,N_465);
or U2662 (N_2662,N_1010,N_820);
nor U2663 (N_2663,N_618,N_919);
nand U2664 (N_2664,N_73,N_263);
xor U2665 (N_2665,N_1478,N_802);
and U2666 (N_2666,N_1483,N_1374);
and U2667 (N_2667,N_45,N_1277);
or U2668 (N_2668,N_915,N_1376);
nor U2669 (N_2669,N_822,N_286);
and U2670 (N_2670,N_954,N_261);
nand U2671 (N_2671,N_286,N_55);
or U2672 (N_2672,N_947,N_802);
xnor U2673 (N_2673,N_1037,N_434);
or U2674 (N_2674,N_1385,N_1101);
nor U2675 (N_2675,N_15,N_1241);
nor U2676 (N_2676,N_1319,N_964);
xor U2677 (N_2677,N_190,N_1333);
nor U2678 (N_2678,N_1491,N_223);
and U2679 (N_2679,N_1322,N_66);
or U2680 (N_2680,N_1470,N_446);
xnor U2681 (N_2681,N_604,N_1423);
and U2682 (N_2682,N_493,N_1416);
nor U2683 (N_2683,N_1402,N_430);
nand U2684 (N_2684,N_566,N_245);
nor U2685 (N_2685,N_212,N_131);
nor U2686 (N_2686,N_379,N_1393);
nand U2687 (N_2687,N_1170,N_496);
nand U2688 (N_2688,N_699,N_1466);
or U2689 (N_2689,N_102,N_662);
and U2690 (N_2690,N_586,N_918);
and U2691 (N_2691,N_509,N_979);
nor U2692 (N_2692,N_1459,N_571);
and U2693 (N_2693,N_147,N_122);
and U2694 (N_2694,N_687,N_841);
and U2695 (N_2695,N_78,N_1236);
and U2696 (N_2696,N_1282,N_676);
nand U2697 (N_2697,N_799,N_931);
nand U2698 (N_2698,N_1241,N_311);
nor U2699 (N_2699,N_511,N_387);
xor U2700 (N_2700,N_751,N_152);
or U2701 (N_2701,N_244,N_467);
nor U2702 (N_2702,N_922,N_492);
and U2703 (N_2703,N_909,N_1433);
or U2704 (N_2704,N_1142,N_1167);
or U2705 (N_2705,N_138,N_529);
and U2706 (N_2706,N_85,N_410);
or U2707 (N_2707,N_771,N_105);
nor U2708 (N_2708,N_99,N_818);
nor U2709 (N_2709,N_54,N_786);
and U2710 (N_2710,N_1481,N_918);
and U2711 (N_2711,N_269,N_1386);
and U2712 (N_2712,N_1365,N_404);
and U2713 (N_2713,N_744,N_1257);
nor U2714 (N_2714,N_570,N_468);
nor U2715 (N_2715,N_633,N_1161);
and U2716 (N_2716,N_444,N_638);
nand U2717 (N_2717,N_1307,N_776);
and U2718 (N_2718,N_1258,N_174);
and U2719 (N_2719,N_338,N_949);
nor U2720 (N_2720,N_1123,N_191);
nand U2721 (N_2721,N_187,N_749);
xor U2722 (N_2722,N_916,N_1281);
nor U2723 (N_2723,N_63,N_757);
or U2724 (N_2724,N_1453,N_1461);
or U2725 (N_2725,N_437,N_290);
nand U2726 (N_2726,N_932,N_928);
or U2727 (N_2727,N_1150,N_413);
or U2728 (N_2728,N_1089,N_0);
nor U2729 (N_2729,N_714,N_697);
or U2730 (N_2730,N_1459,N_1012);
or U2731 (N_2731,N_162,N_460);
nand U2732 (N_2732,N_955,N_657);
and U2733 (N_2733,N_573,N_89);
and U2734 (N_2734,N_745,N_837);
nand U2735 (N_2735,N_153,N_660);
nand U2736 (N_2736,N_727,N_1032);
nor U2737 (N_2737,N_1481,N_1222);
xnor U2738 (N_2738,N_1419,N_1422);
and U2739 (N_2739,N_1189,N_1397);
and U2740 (N_2740,N_441,N_1185);
and U2741 (N_2741,N_895,N_1033);
nand U2742 (N_2742,N_758,N_1426);
nor U2743 (N_2743,N_542,N_1255);
xnor U2744 (N_2744,N_69,N_1222);
and U2745 (N_2745,N_974,N_438);
and U2746 (N_2746,N_1191,N_867);
xor U2747 (N_2747,N_1226,N_1398);
nand U2748 (N_2748,N_176,N_996);
nor U2749 (N_2749,N_279,N_404);
or U2750 (N_2750,N_731,N_851);
nand U2751 (N_2751,N_164,N_847);
xnor U2752 (N_2752,N_674,N_672);
nand U2753 (N_2753,N_255,N_48);
and U2754 (N_2754,N_859,N_547);
and U2755 (N_2755,N_1074,N_1218);
nor U2756 (N_2756,N_936,N_765);
or U2757 (N_2757,N_1114,N_517);
or U2758 (N_2758,N_476,N_890);
or U2759 (N_2759,N_1416,N_343);
xor U2760 (N_2760,N_389,N_105);
xnor U2761 (N_2761,N_601,N_836);
and U2762 (N_2762,N_1269,N_649);
xor U2763 (N_2763,N_1123,N_320);
or U2764 (N_2764,N_21,N_1045);
or U2765 (N_2765,N_536,N_259);
nor U2766 (N_2766,N_498,N_1235);
and U2767 (N_2767,N_1,N_197);
and U2768 (N_2768,N_1178,N_69);
nor U2769 (N_2769,N_1323,N_1406);
and U2770 (N_2770,N_1470,N_355);
and U2771 (N_2771,N_812,N_611);
and U2772 (N_2772,N_580,N_1119);
and U2773 (N_2773,N_743,N_9);
nor U2774 (N_2774,N_657,N_428);
and U2775 (N_2775,N_71,N_986);
nor U2776 (N_2776,N_1145,N_308);
and U2777 (N_2777,N_1037,N_1157);
nor U2778 (N_2778,N_1367,N_808);
nor U2779 (N_2779,N_1085,N_1092);
or U2780 (N_2780,N_991,N_1204);
and U2781 (N_2781,N_1096,N_731);
nor U2782 (N_2782,N_42,N_448);
or U2783 (N_2783,N_792,N_478);
xnor U2784 (N_2784,N_375,N_350);
and U2785 (N_2785,N_791,N_1038);
nor U2786 (N_2786,N_1431,N_97);
nor U2787 (N_2787,N_1182,N_181);
xnor U2788 (N_2788,N_1437,N_1159);
or U2789 (N_2789,N_770,N_29);
and U2790 (N_2790,N_1337,N_996);
or U2791 (N_2791,N_1358,N_1186);
or U2792 (N_2792,N_1429,N_163);
xnor U2793 (N_2793,N_790,N_1251);
and U2794 (N_2794,N_599,N_1009);
xnor U2795 (N_2795,N_402,N_613);
xnor U2796 (N_2796,N_1286,N_840);
and U2797 (N_2797,N_1296,N_913);
nor U2798 (N_2798,N_89,N_1413);
nor U2799 (N_2799,N_376,N_968);
nor U2800 (N_2800,N_1394,N_90);
and U2801 (N_2801,N_1212,N_1483);
nand U2802 (N_2802,N_1245,N_276);
xnor U2803 (N_2803,N_328,N_265);
xnor U2804 (N_2804,N_1448,N_1104);
xor U2805 (N_2805,N_1477,N_188);
xor U2806 (N_2806,N_193,N_8);
or U2807 (N_2807,N_1355,N_1215);
or U2808 (N_2808,N_77,N_1150);
nand U2809 (N_2809,N_1109,N_411);
xnor U2810 (N_2810,N_1065,N_1157);
nor U2811 (N_2811,N_575,N_332);
nand U2812 (N_2812,N_1062,N_544);
and U2813 (N_2813,N_1202,N_464);
nor U2814 (N_2814,N_1070,N_1367);
nand U2815 (N_2815,N_1277,N_821);
nor U2816 (N_2816,N_645,N_1299);
or U2817 (N_2817,N_1465,N_749);
or U2818 (N_2818,N_589,N_412);
and U2819 (N_2819,N_177,N_570);
or U2820 (N_2820,N_1097,N_1401);
nor U2821 (N_2821,N_228,N_1495);
nand U2822 (N_2822,N_1171,N_1406);
xnor U2823 (N_2823,N_376,N_549);
xor U2824 (N_2824,N_1432,N_224);
nand U2825 (N_2825,N_1403,N_562);
nor U2826 (N_2826,N_945,N_604);
nand U2827 (N_2827,N_527,N_1144);
nand U2828 (N_2828,N_723,N_1274);
nor U2829 (N_2829,N_385,N_1358);
and U2830 (N_2830,N_1432,N_623);
and U2831 (N_2831,N_1266,N_0);
xor U2832 (N_2832,N_1051,N_1144);
xor U2833 (N_2833,N_440,N_1303);
nor U2834 (N_2834,N_957,N_451);
or U2835 (N_2835,N_1095,N_1043);
nor U2836 (N_2836,N_595,N_949);
xnor U2837 (N_2837,N_570,N_1007);
nand U2838 (N_2838,N_1339,N_1031);
nor U2839 (N_2839,N_472,N_1342);
xnor U2840 (N_2840,N_1245,N_75);
xnor U2841 (N_2841,N_22,N_622);
nor U2842 (N_2842,N_1490,N_288);
nand U2843 (N_2843,N_1097,N_686);
nand U2844 (N_2844,N_399,N_19);
xnor U2845 (N_2845,N_862,N_1379);
xnor U2846 (N_2846,N_718,N_473);
nor U2847 (N_2847,N_635,N_862);
nand U2848 (N_2848,N_1136,N_1406);
and U2849 (N_2849,N_452,N_1437);
nor U2850 (N_2850,N_534,N_179);
or U2851 (N_2851,N_171,N_18);
xnor U2852 (N_2852,N_518,N_185);
nand U2853 (N_2853,N_1122,N_663);
xnor U2854 (N_2854,N_1458,N_305);
and U2855 (N_2855,N_871,N_173);
nor U2856 (N_2856,N_1306,N_1064);
and U2857 (N_2857,N_9,N_491);
nand U2858 (N_2858,N_802,N_129);
or U2859 (N_2859,N_787,N_922);
and U2860 (N_2860,N_163,N_934);
nand U2861 (N_2861,N_1245,N_645);
nor U2862 (N_2862,N_1401,N_566);
and U2863 (N_2863,N_1333,N_841);
nand U2864 (N_2864,N_900,N_1147);
or U2865 (N_2865,N_135,N_938);
nand U2866 (N_2866,N_1464,N_1479);
nor U2867 (N_2867,N_30,N_1280);
or U2868 (N_2868,N_1104,N_1209);
or U2869 (N_2869,N_57,N_472);
or U2870 (N_2870,N_1083,N_426);
and U2871 (N_2871,N_820,N_993);
and U2872 (N_2872,N_108,N_1389);
or U2873 (N_2873,N_666,N_1085);
and U2874 (N_2874,N_1027,N_107);
xnor U2875 (N_2875,N_509,N_1476);
and U2876 (N_2876,N_1010,N_343);
or U2877 (N_2877,N_149,N_308);
nand U2878 (N_2878,N_711,N_1464);
xor U2879 (N_2879,N_1060,N_124);
nor U2880 (N_2880,N_386,N_944);
or U2881 (N_2881,N_929,N_1222);
or U2882 (N_2882,N_901,N_642);
nand U2883 (N_2883,N_584,N_216);
or U2884 (N_2884,N_774,N_417);
and U2885 (N_2885,N_1092,N_1273);
nor U2886 (N_2886,N_263,N_1203);
and U2887 (N_2887,N_353,N_64);
and U2888 (N_2888,N_1335,N_1099);
nor U2889 (N_2889,N_1030,N_790);
nor U2890 (N_2890,N_562,N_50);
and U2891 (N_2891,N_1444,N_294);
xor U2892 (N_2892,N_1353,N_1382);
nand U2893 (N_2893,N_118,N_739);
nand U2894 (N_2894,N_488,N_791);
or U2895 (N_2895,N_1011,N_378);
or U2896 (N_2896,N_1024,N_83);
xnor U2897 (N_2897,N_664,N_374);
or U2898 (N_2898,N_113,N_210);
and U2899 (N_2899,N_1103,N_1147);
nor U2900 (N_2900,N_1471,N_592);
nor U2901 (N_2901,N_1153,N_1089);
or U2902 (N_2902,N_363,N_98);
nor U2903 (N_2903,N_48,N_267);
and U2904 (N_2904,N_256,N_618);
nand U2905 (N_2905,N_450,N_88);
nand U2906 (N_2906,N_124,N_1445);
nand U2907 (N_2907,N_1298,N_297);
or U2908 (N_2908,N_1385,N_330);
xor U2909 (N_2909,N_983,N_1313);
or U2910 (N_2910,N_454,N_78);
and U2911 (N_2911,N_1139,N_720);
or U2912 (N_2912,N_1008,N_230);
and U2913 (N_2913,N_1204,N_1018);
or U2914 (N_2914,N_1498,N_326);
xnor U2915 (N_2915,N_792,N_1254);
and U2916 (N_2916,N_289,N_235);
or U2917 (N_2917,N_1122,N_436);
xor U2918 (N_2918,N_368,N_634);
nand U2919 (N_2919,N_1213,N_544);
xor U2920 (N_2920,N_999,N_287);
xor U2921 (N_2921,N_782,N_1397);
and U2922 (N_2922,N_59,N_1192);
nand U2923 (N_2923,N_5,N_14);
or U2924 (N_2924,N_929,N_1371);
nand U2925 (N_2925,N_994,N_377);
and U2926 (N_2926,N_21,N_1493);
and U2927 (N_2927,N_119,N_1173);
xor U2928 (N_2928,N_1184,N_1160);
or U2929 (N_2929,N_713,N_1104);
or U2930 (N_2930,N_715,N_465);
and U2931 (N_2931,N_1306,N_745);
or U2932 (N_2932,N_1273,N_435);
or U2933 (N_2933,N_1468,N_173);
xor U2934 (N_2934,N_25,N_1001);
nand U2935 (N_2935,N_825,N_848);
nor U2936 (N_2936,N_448,N_845);
or U2937 (N_2937,N_660,N_573);
xnor U2938 (N_2938,N_416,N_227);
nand U2939 (N_2939,N_624,N_604);
nor U2940 (N_2940,N_234,N_1187);
nor U2941 (N_2941,N_294,N_1440);
xor U2942 (N_2942,N_519,N_609);
nor U2943 (N_2943,N_706,N_450);
xnor U2944 (N_2944,N_1148,N_61);
xnor U2945 (N_2945,N_885,N_319);
nand U2946 (N_2946,N_79,N_770);
nand U2947 (N_2947,N_670,N_1387);
nand U2948 (N_2948,N_595,N_115);
nand U2949 (N_2949,N_1287,N_1186);
nor U2950 (N_2950,N_986,N_995);
xnor U2951 (N_2951,N_521,N_963);
nor U2952 (N_2952,N_114,N_401);
nor U2953 (N_2953,N_343,N_1130);
xnor U2954 (N_2954,N_1390,N_567);
xor U2955 (N_2955,N_1013,N_386);
xor U2956 (N_2956,N_444,N_1372);
xnor U2957 (N_2957,N_453,N_621);
nand U2958 (N_2958,N_1305,N_636);
nor U2959 (N_2959,N_1009,N_1400);
or U2960 (N_2960,N_458,N_1300);
nor U2961 (N_2961,N_1497,N_1228);
and U2962 (N_2962,N_734,N_780);
xor U2963 (N_2963,N_826,N_930);
xor U2964 (N_2964,N_309,N_604);
nand U2965 (N_2965,N_1226,N_352);
xnor U2966 (N_2966,N_803,N_114);
or U2967 (N_2967,N_1156,N_667);
xnor U2968 (N_2968,N_156,N_1416);
nor U2969 (N_2969,N_751,N_443);
xor U2970 (N_2970,N_600,N_1275);
xnor U2971 (N_2971,N_75,N_1364);
nand U2972 (N_2972,N_829,N_744);
nand U2973 (N_2973,N_620,N_1363);
and U2974 (N_2974,N_615,N_232);
xor U2975 (N_2975,N_1121,N_42);
xnor U2976 (N_2976,N_1293,N_20);
or U2977 (N_2977,N_365,N_1072);
nand U2978 (N_2978,N_1003,N_57);
or U2979 (N_2979,N_564,N_515);
or U2980 (N_2980,N_142,N_488);
xor U2981 (N_2981,N_1481,N_276);
nand U2982 (N_2982,N_470,N_266);
xnor U2983 (N_2983,N_1398,N_1422);
nor U2984 (N_2984,N_1433,N_363);
and U2985 (N_2985,N_550,N_809);
nor U2986 (N_2986,N_144,N_1342);
xor U2987 (N_2987,N_42,N_1354);
xor U2988 (N_2988,N_275,N_1260);
nand U2989 (N_2989,N_591,N_1202);
xor U2990 (N_2990,N_1449,N_576);
and U2991 (N_2991,N_1284,N_247);
and U2992 (N_2992,N_367,N_219);
or U2993 (N_2993,N_81,N_1134);
and U2994 (N_2994,N_247,N_1048);
xor U2995 (N_2995,N_1067,N_1252);
nand U2996 (N_2996,N_443,N_503);
and U2997 (N_2997,N_608,N_377);
nor U2998 (N_2998,N_768,N_103);
and U2999 (N_2999,N_150,N_1123);
nor U3000 (N_3000,N_2672,N_2012);
xor U3001 (N_3001,N_2310,N_1694);
nor U3002 (N_3002,N_2671,N_2673);
or U3003 (N_3003,N_1809,N_1986);
nor U3004 (N_3004,N_2630,N_2738);
nand U3005 (N_3005,N_2354,N_2072);
or U3006 (N_3006,N_1811,N_2667);
or U3007 (N_3007,N_2773,N_1538);
and U3008 (N_3008,N_2639,N_2790);
nand U3009 (N_3009,N_2538,N_1923);
nand U3010 (N_3010,N_1963,N_2005);
nand U3011 (N_3011,N_2471,N_1934);
xnor U3012 (N_3012,N_1582,N_1855);
and U3013 (N_3013,N_1964,N_1877);
nor U3014 (N_3014,N_2832,N_1559);
nor U3015 (N_3015,N_1971,N_2323);
xor U3016 (N_3016,N_1524,N_2737);
xnor U3017 (N_3017,N_1626,N_2021);
nor U3018 (N_3018,N_2339,N_1565);
xnor U3019 (N_3019,N_2719,N_2970);
or U3020 (N_3020,N_2782,N_2324);
xor U3021 (N_3021,N_2210,N_2933);
nand U3022 (N_3022,N_2155,N_2349);
nand U3023 (N_3023,N_2894,N_2849);
xor U3024 (N_3024,N_2979,N_2247);
xor U3025 (N_3025,N_1662,N_2208);
and U3026 (N_3026,N_1701,N_2263);
and U3027 (N_3027,N_1543,N_2364);
nand U3028 (N_3028,N_2664,N_2862);
and U3029 (N_3029,N_2957,N_2513);
or U3030 (N_3030,N_2212,N_1653);
or U3031 (N_3031,N_1527,N_2746);
and U3032 (N_3032,N_2020,N_2000);
nand U3033 (N_3033,N_1967,N_2176);
or U3034 (N_3034,N_2465,N_1896);
xor U3035 (N_3035,N_2990,N_2512);
or U3036 (N_3036,N_2190,N_2917);
and U3037 (N_3037,N_1925,N_2191);
and U3038 (N_3038,N_1797,N_2615);
and U3039 (N_3039,N_1723,N_1898);
and U3040 (N_3040,N_2199,N_2996);
or U3041 (N_3041,N_1875,N_2861);
nor U3042 (N_3042,N_2087,N_2459);
and U3043 (N_3043,N_1759,N_1608);
or U3044 (N_3044,N_1622,N_2988);
nand U3045 (N_3045,N_2076,N_2825);
nand U3046 (N_3046,N_1750,N_2332);
nor U3047 (N_3047,N_2940,N_2807);
nand U3048 (N_3048,N_1610,N_2198);
nor U3049 (N_3049,N_1516,N_2216);
nor U3050 (N_3050,N_1724,N_2074);
nor U3051 (N_3051,N_1501,N_1748);
xor U3052 (N_3052,N_1767,N_1857);
nor U3053 (N_3053,N_1871,N_1771);
nor U3054 (N_3054,N_1692,N_2706);
and U3055 (N_3055,N_2469,N_2014);
nor U3056 (N_3056,N_1799,N_2860);
xor U3057 (N_3057,N_1769,N_1914);
and U3058 (N_3058,N_1932,N_2575);
nor U3059 (N_3059,N_1534,N_2817);
nor U3060 (N_3060,N_2347,N_2529);
nand U3061 (N_3061,N_2759,N_1677);
xor U3062 (N_3062,N_2740,N_2404);
and U3063 (N_3063,N_1589,N_1900);
and U3064 (N_3064,N_1599,N_1737);
nor U3065 (N_3065,N_1979,N_1879);
or U3066 (N_3066,N_2268,N_2408);
or U3067 (N_3067,N_2246,N_1581);
nand U3068 (N_3068,N_1834,N_1808);
or U3069 (N_3069,N_2526,N_2472);
nand U3070 (N_3070,N_1725,N_1508);
and U3071 (N_3071,N_1937,N_2666);
nand U3072 (N_3072,N_2953,N_2995);
or U3073 (N_3073,N_2889,N_2045);
nor U3074 (N_3074,N_2770,N_1732);
xor U3075 (N_3075,N_2941,N_2421);
nand U3076 (N_3076,N_1933,N_2233);
nand U3077 (N_3077,N_2458,N_1783);
and U3078 (N_3078,N_1598,N_2697);
nand U3079 (N_3079,N_1576,N_2569);
xor U3080 (N_3080,N_2661,N_2333);
or U3081 (N_3081,N_2618,N_2476);
or U3082 (N_3082,N_2031,N_2629);
or U3083 (N_3083,N_2820,N_1616);
or U3084 (N_3084,N_2209,N_2428);
nand U3085 (N_3085,N_2919,N_2822);
xnor U3086 (N_3086,N_2343,N_1786);
nand U3087 (N_3087,N_1736,N_2909);
nor U3088 (N_3088,N_2732,N_2296);
xor U3089 (N_3089,N_2637,N_2857);
xnor U3090 (N_3090,N_1792,N_1890);
and U3091 (N_3091,N_2346,N_1530);
nand U3092 (N_3092,N_2295,N_2393);
or U3093 (N_3093,N_1948,N_2748);
xor U3094 (N_3094,N_2511,N_2287);
nand U3095 (N_3095,N_1968,N_2207);
xor U3096 (N_3096,N_2974,N_2138);
nand U3097 (N_3097,N_2029,N_1632);
nor U3098 (N_3098,N_1717,N_2897);
xnor U3099 (N_3099,N_1515,N_1707);
xnor U3100 (N_3100,N_2419,N_2888);
nor U3101 (N_3101,N_2409,N_2131);
and U3102 (N_3102,N_1615,N_2388);
nor U3103 (N_3103,N_2612,N_2293);
nand U3104 (N_3104,N_2032,N_2997);
and U3105 (N_3105,N_2305,N_2621);
and U3106 (N_3106,N_1838,N_2555);
xor U3107 (N_3107,N_2687,N_2464);
or U3108 (N_3108,N_2470,N_2224);
or U3109 (N_3109,N_2405,N_2378);
and U3110 (N_3110,N_1836,N_2396);
or U3111 (N_3111,N_2248,N_1824);
nor U3112 (N_3112,N_2192,N_2731);
nor U3113 (N_3113,N_2185,N_2656);
xnor U3114 (N_3114,N_2586,N_2973);
or U3115 (N_3115,N_2286,N_2805);
and U3116 (N_3116,N_1863,N_2927);
nand U3117 (N_3117,N_1651,N_2447);
and U3118 (N_3118,N_1931,N_2699);
nand U3119 (N_3119,N_1828,N_2800);
nand U3120 (N_3120,N_2942,N_2379);
or U3121 (N_3121,N_2478,N_2360);
and U3122 (N_3122,N_1664,N_2585);
xor U3123 (N_3123,N_2754,N_2027);
nand U3124 (N_3124,N_2395,N_2509);
nor U3125 (N_3125,N_2826,N_2230);
or U3126 (N_3126,N_2718,N_2382);
nor U3127 (N_3127,N_1944,N_2689);
xor U3128 (N_3128,N_2389,N_1675);
nor U3129 (N_3129,N_2978,N_2406);
xnor U3130 (N_3130,N_1974,N_2607);
or U3131 (N_3131,N_1734,N_1917);
or U3132 (N_3132,N_1669,N_2231);
or U3133 (N_3133,N_2505,N_1636);
xnor U3134 (N_3134,N_2438,N_1595);
nor U3135 (N_3135,N_2819,N_1679);
nor U3136 (N_3136,N_1523,N_1922);
or U3137 (N_3137,N_2847,N_1854);
nand U3138 (N_3138,N_2106,N_2308);
or U3139 (N_3139,N_1689,N_1814);
and U3140 (N_3140,N_1874,N_2911);
nand U3141 (N_3141,N_1887,N_2537);
nand U3142 (N_3142,N_2194,N_1548);
or U3143 (N_3143,N_1529,N_2709);
nor U3144 (N_3144,N_2399,N_2119);
nor U3145 (N_3145,N_1696,N_2864);
xnor U3146 (N_3146,N_2040,N_1577);
nand U3147 (N_3147,N_2550,N_2427);
and U3148 (N_3148,N_2603,N_2884);
or U3149 (N_3149,N_1815,N_2734);
nand U3150 (N_3150,N_2763,N_1729);
nand U3151 (N_3151,N_2402,N_1652);
or U3152 (N_3152,N_2651,N_2275);
nor U3153 (N_3153,N_1590,N_2368);
xor U3154 (N_3154,N_1721,N_2613);
or U3155 (N_3155,N_2180,N_2262);
nor U3156 (N_3156,N_2278,N_1657);
nor U3157 (N_3157,N_2223,N_2253);
or U3158 (N_3158,N_2939,N_1753);
and U3159 (N_3159,N_2831,N_2004);
or U3160 (N_3160,N_2558,N_2760);
and U3161 (N_3161,N_1770,N_1568);
and U3162 (N_3162,N_1884,N_2636);
nand U3163 (N_3163,N_1775,N_2196);
xor U3164 (N_3164,N_2264,N_2442);
nor U3165 (N_3165,N_1605,N_2779);
nor U3166 (N_3166,N_2153,N_2147);
xnor U3167 (N_3167,N_2975,N_2983);
and U3168 (N_3168,N_2808,N_2980);
or U3169 (N_3169,N_2658,N_1682);
nand U3170 (N_3170,N_2869,N_1525);
or U3171 (N_3171,N_2092,N_2755);
nor U3172 (N_3172,N_1902,N_1895);
and U3173 (N_3173,N_2735,N_2705);
nand U3174 (N_3174,N_1904,N_1790);
nor U3175 (N_3175,N_1791,N_2200);
xor U3176 (N_3176,N_2007,N_1969);
xor U3177 (N_3177,N_2814,N_2945);
nor U3178 (N_3178,N_2815,N_2110);
and U3179 (N_3179,N_2767,N_2798);
xor U3180 (N_3180,N_2015,N_1713);
nand U3181 (N_3181,N_1778,N_2976);
or U3182 (N_3182,N_1951,N_2056);
or U3183 (N_3183,N_1620,N_2033);
and U3184 (N_3184,N_2958,N_2670);
nand U3185 (N_3185,N_2843,N_2340);
xor U3186 (N_3186,N_1659,N_1945);
nor U3187 (N_3187,N_2193,N_2619);
nand U3188 (N_3188,N_2236,N_1740);
nor U3189 (N_3189,N_2758,N_2398);
nand U3190 (N_3190,N_2969,N_2749);
nor U3191 (N_3191,N_2502,N_2440);
nor U3192 (N_3192,N_2693,N_2225);
or U3193 (N_3193,N_2016,N_1640);
xnor U3194 (N_3194,N_1924,N_1893);
or U3195 (N_3195,N_1788,N_2606);
or U3196 (N_3196,N_2307,N_2099);
and U3197 (N_3197,N_2806,N_2828);
nor U3198 (N_3198,N_2044,N_1929);
xnor U3199 (N_3199,N_1774,N_1983);
nand U3200 (N_3200,N_1848,N_1935);
nor U3201 (N_3201,N_2149,N_2752);
and U3202 (N_3202,N_2648,N_2517);
nand U3203 (N_3203,N_1830,N_2313);
nand U3204 (N_3204,N_1978,N_1625);
or U3205 (N_3205,N_2736,N_2183);
nor U3206 (N_3206,N_2947,N_1741);
and U3207 (N_3207,N_2314,N_1649);
or U3208 (N_3208,N_2886,N_2152);
xnor U3209 (N_3209,N_2720,N_1995);
nand U3210 (N_3210,N_1596,N_1954);
nor U3211 (N_3211,N_2416,N_1812);
nand U3212 (N_3212,N_1905,N_2563);
and U3213 (N_3213,N_2468,N_2091);
and U3214 (N_3214,N_2453,N_2038);
xnor U3215 (N_3215,N_2053,N_2113);
or U3216 (N_3216,N_1521,N_2877);
xor U3217 (N_3217,N_2120,N_2116);
xor U3218 (N_3218,N_1704,N_1813);
or U3219 (N_3219,N_2257,N_1624);
xnor U3220 (N_3220,N_2226,N_2080);
nor U3221 (N_3221,N_2177,N_2593);
and U3222 (N_3222,N_1678,N_1901);
nand U3223 (N_3223,N_2677,N_1756);
xnor U3224 (N_3224,N_1897,N_2241);
nand U3225 (N_3225,N_2583,N_2083);
nor U3226 (N_3226,N_2187,N_2048);
and U3227 (N_3227,N_1795,N_1899);
or U3228 (N_3228,N_2627,N_2551);
or U3229 (N_3229,N_2809,N_2006);
and U3230 (N_3230,N_2853,N_1735);
or U3231 (N_3231,N_2986,N_2361);
xor U3232 (N_3232,N_2963,N_2559);
xnor U3233 (N_3233,N_2655,N_2436);
xnor U3234 (N_3234,N_2011,N_2829);
or U3235 (N_3235,N_2994,N_2730);
xor U3236 (N_3236,N_1798,N_2154);
and U3237 (N_3237,N_2306,N_1910);
and U3238 (N_3238,N_2552,N_2678);
or U3239 (N_3239,N_2383,N_1613);
nor U3240 (N_3240,N_1670,N_2486);
xnor U3241 (N_3241,N_2240,N_1645);
or U3242 (N_3242,N_1804,N_2365);
xor U3243 (N_3243,N_2878,N_1747);
nor U3244 (N_3244,N_1697,N_2576);
nand U3245 (N_3245,N_1999,N_2542);
nor U3246 (N_3246,N_2483,N_2355);
nand U3247 (N_3247,N_1635,N_2777);
nand U3248 (N_3248,N_1742,N_1558);
or U3249 (N_3249,N_1593,N_1540);
xor U3250 (N_3250,N_2810,N_2665);
or U3251 (N_3251,N_1858,N_2319);
nand U3252 (N_3252,N_2725,N_2686);
xnor U3253 (N_3253,N_2245,N_2218);
xnor U3254 (N_3254,N_2766,N_1843);
nand U3255 (N_3255,N_2858,N_1684);
and U3256 (N_3256,N_2097,N_2114);
and U3257 (N_3257,N_2867,N_2088);
nand U3258 (N_3258,N_1793,N_2950);
xor U3259 (N_3259,N_1578,N_2201);
or U3260 (N_3260,N_1876,N_1965);
nor U3261 (N_3261,N_1668,N_2765);
nand U3262 (N_3262,N_2384,N_1998);
nor U3263 (N_3263,N_1566,N_2567);
and U3264 (N_3264,N_2222,N_1891);
xnor U3265 (N_3265,N_2645,N_1644);
and U3266 (N_3266,N_1604,N_1611);
xor U3267 (N_3267,N_2420,N_1569);
xor U3268 (N_3268,N_2444,N_1617);
or U3269 (N_3269,N_2675,N_1821);
and U3270 (N_3270,N_2217,N_1686);
and U3271 (N_3271,N_1535,N_2273);
or U3272 (N_3272,N_2165,N_2882);
nor U3273 (N_3273,N_2682,N_2516);
nand U3274 (N_3274,N_1502,N_2277);
nand U3275 (N_3275,N_1544,N_2249);
xor U3276 (N_3276,N_1818,N_2497);
xnor U3277 (N_3277,N_1514,N_2414);
nand U3278 (N_3278,N_2663,N_2780);
nand U3279 (N_3279,N_1950,N_2608);
nand U3280 (N_3280,N_2572,N_2587);
nor U3281 (N_3281,N_2424,N_2433);
nor U3282 (N_3282,N_1762,N_2485);
or U3283 (N_3283,N_2244,N_1563);
and U3284 (N_3284,N_1602,N_1648);
and U3285 (N_3285,N_1851,N_2359);
nand U3286 (N_3286,N_2003,N_2842);
nor U3287 (N_3287,N_2900,N_1953);
nor U3288 (N_3288,N_1634,N_2337);
nand U3289 (N_3289,N_1827,N_2523);
or U3290 (N_3290,N_2981,N_2065);
or U3291 (N_3291,N_2134,N_2018);
nand U3292 (N_3292,N_2881,N_1779);
xnor U3293 (N_3293,N_2885,N_2167);
xor U3294 (N_3294,N_1955,N_2142);
nand U3295 (N_3295,N_2646,N_2381);
and U3296 (N_3296,N_2616,N_2727);
nand U3297 (N_3297,N_2600,N_2928);
nor U3298 (N_3298,N_2024,N_1731);
nor U3299 (N_3299,N_2300,N_1641);
nor U3300 (N_3300,N_2772,N_1739);
nor U3301 (N_3301,N_2852,N_2804);
or U3302 (N_3302,N_2172,N_2066);
nand U3303 (N_3303,N_1591,N_2292);
nand U3304 (N_3304,N_2127,N_2220);
or U3305 (N_3305,N_1660,N_2547);
and U3306 (N_3306,N_2188,N_2090);
or U3307 (N_3307,N_2144,N_2951);
and U3308 (N_3308,N_2256,N_1772);
nand U3309 (N_3309,N_2683,N_2078);
and U3310 (N_3310,N_2905,N_2922);
or U3311 (N_3311,N_2660,N_2640);
and U3312 (N_3312,N_2930,N_1532);
nand U3313 (N_3313,N_1962,N_1504);
nand U3314 (N_3314,N_2123,N_2899);
xnor U3315 (N_3315,N_2330,N_1867);
xnor U3316 (N_3316,N_2270,N_2688);
nor U3317 (N_3317,N_2774,N_2653);
nand U3318 (N_3318,N_2624,N_2329);
and U3319 (N_3319,N_2801,N_1958);
and U3320 (N_3320,N_2694,N_2013);
and U3321 (N_3321,N_2258,N_2681);
and U3322 (N_3322,N_1882,N_1961);
xnor U3323 (N_3323,N_2069,N_2622);
or U3324 (N_3324,N_2943,N_2281);
and U3325 (N_3325,N_2499,N_2534);
xor U3326 (N_3326,N_2309,N_1913);
and U3327 (N_3327,N_2617,N_2866);
or U3328 (N_3328,N_2541,N_2136);
or U3329 (N_3329,N_2077,N_2906);
nand U3330 (N_3330,N_2315,N_2489);
or U3331 (N_3331,N_2284,N_1564);
nand U3332 (N_3332,N_1687,N_2034);
nor U3333 (N_3333,N_1623,N_2674);
or U3334 (N_3334,N_1861,N_2680);
nor U3335 (N_3335,N_2265,N_2584);
or U3336 (N_3336,N_1586,N_1702);
nand U3337 (N_3337,N_1561,N_2261);
xor U3338 (N_3338,N_2023,N_2311);
and U3339 (N_3339,N_1722,N_1820);
and U3340 (N_3340,N_2026,N_2903);
or U3341 (N_3341,N_2631,N_1583);
nor U3342 (N_3342,N_1839,N_2601);
nand U3343 (N_3343,N_1650,N_2336);
or U3344 (N_3344,N_2987,N_1763);
nand U3345 (N_3345,N_2375,N_2385);
or U3346 (N_3346,N_2039,N_1878);
nand U3347 (N_3347,N_1628,N_1703);
and U3348 (N_3348,N_1868,N_2321);
and U3349 (N_3349,N_1784,N_2955);
nand U3350 (N_3350,N_2449,N_2043);
and U3351 (N_3351,N_2303,N_2202);
or U3352 (N_3352,N_2566,N_2448);
and U3353 (N_3353,N_1881,N_2064);
nor U3354 (N_3354,N_2374,N_2952);
nor U3355 (N_3355,N_2422,N_2707);
nand U3356 (N_3356,N_2166,N_2999);
xnor U3357 (N_3357,N_1556,N_2966);
xnor U3358 (N_3358,N_2462,N_2904);
nand U3359 (N_3359,N_2451,N_2169);
nor U3360 (N_3360,N_2250,N_2669);
nor U3361 (N_3361,N_2148,N_2086);
xnor U3362 (N_3362,N_2369,N_2984);
and U3363 (N_3363,N_2289,N_2778);
or U3364 (N_3364,N_1567,N_2989);
or U3365 (N_3365,N_2733,N_1614);
or U3366 (N_3366,N_1823,N_1572);
nand U3367 (N_3367,N_1960,N_1700);
nor U3368 (N_3368,N_1849,N_2366);
xnor U3369 (N_3369,N_2691,N_2260);
nor U3370 (N_3370,N_2353,N_1505);
nor U3371 (N_3371,N_1860,N_2662);
nand U3372 (N_3372,N_2873,N_1579);
nor U3373 (N_3373,N_2923,N_1852);
or U3374 (N_3374,N_2839,N_1571);
or U3375 (N_3375,N_2161,N_1959);
or U3376 (N_3376,N_1847,N_1690);
nand U3377 (N_3377,N_2961,N_1536);
xor U3378 (N_3378,N_2920,N_2797);
or U3379 (N_3379,N_1714,N_2386);
xnor U3380 (N_3380,N_2290,N_2418);
or U3381 (N_3381,N_2741,N_2503);
xnor U3382 (N_3382,N_1506,N_2100);
nor U3383 (N_3383,N_1850,N_2628);
and U3384 (N_3384,N_2874,N_2764);
or U3385 (N_3385,N_2341,N_1681);
xor U3386 (N_3386,N_1671,N_2883);
xnor U3387 (N_3387,N_2276,N_2460);
xnor U3388 (N_3388,N_1691,N_2357);
xnor U3389 (N_3389,N_2299,N_1912);
nand U3390 (N_3390,N_2948,N_2178);
and U3391 (N_3391,N_2850,N_1560);
xor U3392 (N_3392,N_1726,N_2577);
and U3393 (N_3393,N_1573,N_2022);
nor U3394 (N_3394,N_1949,N_2791);
or U3395 (N_3395,N_2221,N_2539);
or U3396 (N_3396,N_2750,N_2242);
xor U3397 (N_3397,N_2708,N_1517);
nor U3398 (N_3398,N_2163,N_2528);
nor U3399 (N_3399,N_2568,N_2756);
nand U3400 (N_3400,N_1727,N_1621);
or U3401 (N_3401,N_2322,N_1744);
and U3402 (N_3402,N_2229,N_1637);
xnor U3403 (N_3403,N_2514,N_2959);
or U3404 (N_3404,N_2507,N_2243);
nor U3405 (N_3405,N_1832,N_2157);
or U3406 (N_3406,N_2602,N_1667);
xor U3407 (N_3407,N_2232,N_2742);
nor U3408 (N_3408,N_2103,N_2457);
nand U3409 (N_3409,N_2373,N_1512);
and U3410 (N_3410,N_1764,N_2480);
xor U3411 (N_3411,N_2377,N_2545);
xor U3412 (N_3412,N_2813,N_2796);
nand U3413 (N_3413,N_1992,N_1807);
xor U3414 (N_3414,N_1943,N_2578);
nand U3415 (N_3415,N_1552,N_2685);
nor U3416 (N_3416,N_2895,N_2397);
nor U3417 (N_3417,N_1865,N_2633);
nor U3418 (N_3418,N_1844,N_2085);
nor U3419 (N_3419,N_2964,N_2834);
nand U3420 (N_3420,N_2965,N_2017);
and U3421 (N_3421,N_1688,N_2916);
nand U3422 (N_3422,N_2174,N_2695);
and U3423 (N_3423,N_2345,N_1746);
nor U3424 (N_3424,N_1845,N_1630);
and U3425 (N_3425,N_1862,N_1743);
or U3426 (N_3426,N_2700,N_1580);
nor U3427 (N_3427,N_2151,N_2929);
xnor U3428 (N_3428,N_2274,N_1672);
xnor U3429 (N_3429,N_2946,N_1683);
xnor U3430 (N_3430,N_2871,N_1663);
nor U3431 (N_3431,N_2859,N_2490);
nand U3432 (N_3432,N_2824,N_2252);
nor U3433 (N_3433,N_2267,N_2721);
and U3434 (N_3434,N_1574,N_2073);
nand U3435 (N_3435,N_1647,N_1500);
or U3436 (N_3436,N_1711,N_1547);
or U3437 (N_3437,N_2926,N_1592);
and U3438 (N_3438,N_1705,N_2376);
nand U3439 (N_3439,N_2692,N_2561);
nor U3440 (N_3440,N_2937,N_2219);
or U3441 (N_3441,N_2652,N_1720);
or U3442 (N_3442,N_1507,N_1526);
nor U3443 (N_3443,N_1888,N_1864);
nand U3444 (N_3444,N_2344,N_1835);
nor U3445 (N_3445,N_2008,N_2121);
or U3446 (N_3446,N_2591,N_2908);
or U3447 (N_3447,N_1708,N_2837);
nor U3448 (N_3448,N_1826,N_2704);
or U3449 (N_3449,N_2358,N_2823);
or U3450 (N_3450,N_2280,N_2696);
nor U3451 (N_3451,N_2876,N_1712);
xor U3452 (N_3452,N_2599,N_2326);
and U3453 (N_3453,N_1751,N_2060);
and U3454 (N_3454,N_1886,N_1654);
xor U3455 (N_3455,N_1908,N_2962);
nor U3456 (N_3456,N_1894,N_2811);
or U3457 (N_3457,N_1982,N_2175);
and U3458 (N_3458,N_1991,N_1941);
and U3459 (N_3459,N_2320,N_1819);
nor U3460 (N_3460,N_2082,N_2010);
nor U3461 (N_3461,N_2816,N_2129);
and U3462 (N_3462,N_2715,N_2075);
nor U3463 (N_3463,N_2028,N_2415);
or U3464 (N_3464,N_2195,N_2757);
nand U3465 (N_3465,N_2504,N_2124);
xnor U3466 (N_3466,N_1587,N_1988);
nand U3467 (N_3467,N_2872,N_2743);
nor U3468 (N_3468,N_2605,N_1776);
or U3469 (N_3469,N_2851,N_2794);
or U3470 (N_3470,N_1833,N_2821);
or U3471 (N_3471,N_2972,N_2840);
xor U3472 (N_3472,N_2595,N_2795);
or U3473 (N_3473,N_2977,N_2488);
xnor U3474 (N_3474,N_2215,N_2132);
nor U3475 (N_3475,N_2789,N_2907);
or U3476 (N_3476,N_1817,N_1907);
and U3477 (N_3477,N_2102,N_2213);
or U3478 (N_3478,N_2387,N_1738);
nor U3479 (N_3479,N_1889,N_2186);
nor U3480 (N_3480,N_2392,N_1892);
nor U3481 (N_3481,N_2435,N_1519);
nor U3482 (N_3482,N_1994,N_2592);
or U3483 (N_3483,N_2095,N_1940);
nor U3484 (N_3484,N_2146,N_1869);
nand U3485 (N_3485,N_2351,N_2500);
nor U3486 (N_3486,N_1952,N_1942);
nand U3487 (N_3487,N_2520,N_1509);
or U3488 (N_3488,N_1619,N_1584);
nor U3489 (N_3489,N_2001,N_1977);
and U3490 (N_3490,N_1709,N_2400);
xnor U3491 (N_3491,N_2647,N_1758);
nor U3492 (N_3492,N_2168,N_2835);
and U3493 (N_3493,N_2848,N_2634);
and U3494 (N_3494,N_2938,N_2170);
nor U3495 (N_3495,N_2515,N_2564);
nor U3496 (N_3496,N_1541,N_2527);
or U3497 (N_3497,N_1903,N_2506);
xnor U3498 (N_3498,N_2137,N_2115);
and U3499 (N_3499,N_2162,N_2712);
or U3500 (N_3500,N_2496,N_1699);
and U3501 (N_3501,N_2009,N_2158);
and U3502 (N_3502,N_2203,N_2050);
or U3503 (N_3503,N_2063,N_2912);
nand U3504 (N_3504,N_2423,N_2690);
nor U3505 (N_3505,N_1780,N_2610);
or U3506 (N_3506,N_2025,N_2710);
or U3507 (N_3507,N_2722,N_2474);
nor U3508 (N_3508,N_2312,N_2494);
xnor U3509 (N_3509,N_1752,N_2644);
or U3510 (N_3510,N_1685,N_2540);
nor U3511 (N_3511,N_2784,N_2604);
and U3512 (N_3512,N_2745,N_1926);
or U3513 (N_3513,N_1522,N_1537);
or U3514 (N_3514,N_2944,N_2128);
nor U3515 (N_3515,N_2173,N_2508);
nor U3516 (N_3516,N_2833,N_2543);
or U3517 (N_3517,N_1927,N_1642);
xor U3518 (N_3518,N_2454,N_1656);
nand U3519 (N_3519,N_2108,N_2761);
xor U3520 (N_3520,N_1542,N_1570);
nand U3521 (N_3521,N_2327,N_1825);
nand U3522 (N_3522,N_2184,N_1872);
and U3523 (N_3523,N_1956,N_1531);
and U3524 (N_3524,N_2533,N_1665);
or U3525 (N_3525,N_2067,N_2799);
xor U3526 (N_3526,N_2035,N_1631);
xnor U3527 (N_3527,N_1985,N_2266);
xor U3528 (N_3528,N_1822,N_2298);
nor U3529 (N_3529,N_2519,N_2432);
and U3530 (N_3530,N_1840,N_2051);
and U3531 (N_3531,N_1545,N_1539);
xnor U3532 (N_3532,N_2334,N_1806);
or U3533 (N_3533,N_2614,N_2282);
or U3534 (N_3534,N_2096,N_2046);
or U3535 (N_3535,N_1966,N_2431);
or U3536 (N_3536,N_1607,N_2998);
nor U3537 (N_3537,N_1603,N_1518);
nand U3538 (N_3538,N_2632,N_2181);
nor U3539 (N_3539,N_2856,N_2724);
or U3540 (N_3540,N_2301,N_2679);
xnor U3541 (N_3541,N_2126,N_1760);
nand U3542 (N_3542,N_2531,N_2473);
and U3543 (N_3543,N_2536,N_1710);
xnor U3544 (N_3544,N_2654,N_2921);
xor U3545 (N_3545,N_2788,N_2117);
xor U3546 (N_3546,N_2863,N_2391);
xor U3547 (N_3547,N_2793,N_2211);
xor U3548 (N_3548,N_2501,N_2487);
and U3549 (N_3549,N_2297,N_2620);
nand U3550 (N_3550,N_2914,N_2403);
nor U3551 (N_3551,N_1765,N_2641);
or U3552 (N_3552,N_2288,N_2058);
or U3553 (N_3553,N_2380,N_1639);
nand U3554 (N_3554,N_2141,N_2112);
xnor U3555 (N_3555,N_2093,N_2179);
xnor U3556 (N_3556,N_2122,N_1996);
xor U3557 (N_3557,N_2925,N_1503);
nor U3558 (N_3558,N_1606,N_1754);
nor U3559 (N_3559,N_2104,N_2283);
and U3560 (N_3560,N_1693,N_2739);
nor U3561 (N_3561,N_2036,N_1975);
nand U3562 (N_3562,N_1773,N_2140);
and U3563 (N_3563,N_2827,N_2371);
nand U3564 (N_3564,N_2455,N_2079);
nand U3565 (N_3565,N_2703,N_2484);
nand U3566 (N_3566,N_2237,N_1916);
xor U3567 (N_3567,N_1716,N_1557);
nor U3568 (N_3568,N_1859,N_2803);
nand U3569 (N_3569,N_2560,N_2350);
nand U3570 (N_3570,N_1511,N_2145);
nor U3571 (N_3571,N_2716,N_1918);
xnor U3572 (N_3572,N_2887,N_2896);
nor U3573 (N_3573,N_2934,N_2495);
nand U3574 (N_3574,N_2450,N_1989);
xnor U3575 (N_3575,N_2698,N_2316);
or U3576 (N_3576,N_2626,N_1883);
nor U3577 (N_3577,N_1920,N_2635);
xor U3578 (N_3578,N_1643,N_2935);
or U3579 (N_3579,N_2960,N_2491);
and U3580 (N_3580,N_2783,N_2071);
or U3581 (N_3581,N_2055,N_2352);
xnor U3582 (N_3582,N_2898,N_1749);
or U3583 (N_3583,N_1718,N_2107);
nand U3584 (N_3584,N_1618,N_2331);
and U3585 (N_3585,N_1549,N_2271);
nor U3586 (N_3586,N_1842,N_2325);
or U3587 (N_3587,N_2931,N_2477);
xor U3588 (N_3588,N_2590,N_1629);
or U3589 (N_3589,N_2394,N_2426);
or U3590 (N_3590,N_2294,N_2492);
xnor U3591 (N_3591,N_2135,N_2875);
or U3592 (N_3592,N_2717,N_2956);
nand U3593 (N_3593,N_2781,N_1970);
nor U3594 (N_3594,N_2407,N_1789);
or U3595 (N_3595,N_2052,N_2238);
xnor U3596 (N_3596,N_1655,N_2846);
and U3597 (N_3597,N_2510,N_2818);
nor U3598 (N_3598,N_1676,N_2372);
nor U3599 (N_3599,N_1984,N_2659);
nand U3600 (N_3600,N_2580,N_2753);
xnor U3601 (N_3601,N_1551,N_1785);
nand U3602 (N_3602,N_2150,N_2227);
and U3603 (N_3603,N_2723,N_2481);
xor U3604 (N_3604,N_1866,N_2596);
or U3605 (N_3605,N_2437,N_1936);
nor U3606 (N_3606,N_1782,N_1766);
xnor U3607 (N_3607,N_2910,N_2893);
or U3608 (N_3608,N_2932,N_2643);
and U3609 (N_3609,N_1800,N_2475);
or U3610 (N_3610,N_2776,N_2676);
nor U3611 (N_3611,N_2463,N_2411);
and U3612 (N_3612,N_2164,N_2042);
nand U3613 (N_3613,N_2581,N_2769);
nand U3614 (N_3614,N_2002,N_1698);
or U3615 (N_3615,N_1976,N_2019);
nor U3616 (N_3616,N_2836,N_2668);
xor U3617 (N_3617,N_2802,N_2574);
xor U3618 (N_3618,N_2467,N_1919);
nand U3619 (N_3619,N_2985,N_2768);
nand U3620 (N_3620,N_2684,N_1939);
nand U3621 (N_3621,N_2189,N_2461);
or U3622 (N_3622,N_1921,N_2030);
and U3623 (N_3623,N_1906,N_2439);
and U3624 (N_3624,N_2094,N_1787);
or U3625 (N_3625,N_1885,N_2870);
nand U3626 (N_3626,N_1562,N_2855);
xor U3627 (N_3627,N_1846,N_1550);
xnor U3628 (N_3628,N_2554,N_2061);
nand U3629 (N_3629,N_2589,N_2918);
nor U3630 (N_3630,N_1805,N_2139);
or U3631 (N_3631,N_2650,N_2701);
nor U3632 (N_3632,N_1829,N_2111);
nor U3633 (N_3633,N_2342,N_2070);
xor U3634 (N_3634,N_2390,N_2328);
and U3635 (N_3635,N_2524,N_2098);
or U3636 (N_3636,N_1801,N_2588);
and U3637 (N_3637,N_2452,N_2159);
xnor U3638 (N_3638,N_1673,N_2304);
and U3639 (N_3639,N_2285,N_1594);
xnor U3640 (N_3640,N_1987,N_2785);
nand U3641 (N_3641,N_1554,N_1597);
nand U3642 (N_3642,N_2892,N_2197);
and U3643 (N_3643,N_2992,N_2049);
or U3644 (N_3644,N_2844,N_2556);
nand U3645 (N_3645,N_2054,N_2775);
nor U3646 (N_3646,N_2206,N_2335);
and U3647 (N_3647,N_1761,N_2228);
nor U3648 (N_3648,N_2182,N_2713);
or U3649 (N_3649,N_2714,N_2841);
xnor U3650 (N_3650,N_2982,N_2544);
nand U3651 (N_3651,N_2649,N_2214);
nor U3652 (N_3652,N_1553,N_1930);
xor U3653 (N_3653,N_2562,N_2367);
nand U3654 (N_3654,N_2845,N_2425);
nand U3655 (N_3655,N_2204,N_1781);
nand U3656 (N_3656,N_1973,N_1745);
and U3657 (N_3657,N_1520,N_2711);
or U3658 (N_3658,N_1972,N_2254);
nor U3659 (N_3659,N_1997,N_2251);
or U3660 (N_3660,N_1715,N_2993);
and U3661 (N_3661,N_2412,N_2865);
or U3662 (N_3662,N_2726,N_2417);
xor U3663 (N_3663,N_2272,N_1947);
nand U3664 (N_3664,N_2446,N_1873);
nand U3665 (N_3665,N_2105,N_2548);
xnor U3666 (N_3666,N_2868,N_1796);
xor U3667 (N_3667,N_1880,N_1810);
and U3668 (N_3668,N_2401,N_2239);
or U3669 (N_3669,N_1915,N_1733);
xnor U3670 (N_3670,N_1510,N_2812);
xnor U3671 (N_3671,N_2623,N_1853);
and U3672 (N_3672,N_2830,N_1627);
or U3673 (N_3673,N_2259,N_2109);
and U3674 (N_3674,N_2081,N_1837);
or U3675 (N_3675,N_2786,N_2891);
and U3676 (N_3676,N_2089,N_1658);
nor U3677 (N_3677,N_2879,N_2936);
xnor U3678 (N_3678,N_2047,N_1757);
xnor U3679 (N_3679,N_1728,N_2949);
or U3680 (N_3680,N_1831,N_2570);
nand U3681 (N_3681,N_2302,N_2493);
and U3682 (N_3682,N_2597,N_1674);
nor U3683 (N_3683,N_1609,N_1638);
and U3684 (N_3684,N_2594,N_2611);
xor U3685 (N_3685,N_1980,N_1666);
nor U3686 (N_3686,N_2787,N_2269);
nor U3687 (N_3687,N_2657,N_1981);
nor U3688 (N_3688,N_2041,N_1911);
nor U3689 (N_3689,N_1585,N_1794);
nor U3690 (N_3690,N_2792,N_2901);
nor U3691 (N_3691,N_1588,N_2235);
or U3692 (N_3692,N_2160,N_1528);
nand U3693 (N_3693,N_2413,N_2625);
and U3694 (N_3694,N_2441,N_2902);
nand U3695 (N_3695,N_2445,N_2234);
and U3696 (N_3696,N_2101,N_2522);
and U3697 (N_3697,N_1555,N_2702);
nand U3698 (N_3698,N_1601,N_2370);
or U3699 (N_3699,N_2971,N_2771);
or U3700 (N_3700,N_2546,N_1661);
nor U3701 (N_3701,N_2968,N_2924);
nand U3702 (N_3702,N_2156,N_2443);
xor U3703 (N_3703,N_2525,N_2143);
or U3704 (N_3704,N_1706,N_2171);
and U3705 (N_3705,N_2430,N_2318);
nor U3706 (N_3706,N_1513,N_2890);
and U3707 (N_3707,N_1755,N_2728);
or U3708 (N_3708,N_2518,N_2479);
nor U3709 (N_3709,N_2532,N_2549);
xnor U3710 (N_3710,N_1856,N_1928);
and U3711 (N_3711,N_2609,N_2456);
nand U3712 (N_3712,N_2279,N_1909);
or U3713 (N_3713,N_2363,N_1777);
xnor U3714 (N_3714,N_2466,N_1802);
nor U3715 (N_3715,N_1533,N_2571);
nor U3716 (N_3716,N_2747,N_2744);
and U3717 (N_3717,N_2642,N_2133);
xnor U3718 (N_3718,N_2729,N_2582);
nor U3719 (N_3719,N_1695,N_1841);
and U3720 (N_3720,N_1803,N_2991);
or U3721 (N_3721,N_2967,N_2205);
xnor U3722 (N_3722,N_2762,N_2059);
or U3723 (N_3723,N_1680,N_1768);
xor U3724 (N_3724,N_2557,N_2573);
nor U3725 (N_3725,N_2598,N_2565);
nand U3726 (N_3726,N_2854,N_1600);
nor U3727 (N_3727,N_2084,N_1938);
xnor U3728 (N_3728,N_2255,N_2535);
xnor U3729 (N_3729,N_1990,N_2521);
nand U3730 (N_3730,N_2130,N_2482);
or U3731 (N_3731,N_2579,N_2057);
or U3732 (N_3732,N_1646,N_2062);
nand U3733 (N_3733,N_1816,N_1575);
nand U3734 (N_3734,N_2838,N_1946);
nand U3735 (N_3735,N_2751,N_2434);
nand U3736 (N_3736,N_2338,N_2530);
and U3737 (N_3737,N_2068,N_1612);
nand U3738 (N_3738,N_2037,N_2954);
and U3739 (N_3739,N_2915,N_2317);
and U3740 (N_3740,N_2410,N_2348);
nor U3741 (N_3741,N_1870,N_2638);
xnor U3742 (N_3742,N_2880,N_2291);
xnor U3743 (N_3743,N_1730,N_1633);
and U3744 (N_3744,N_2356,N_2553);
nand U3745 (N_3745,N_1993,N_2125);
nor U3746 (N_3746,N_2429,N_2498);
or U3747 (N_3747,N_1957,N_1546);
nand U3748 (N_3748,N_2118,N_1719);
xor U3749 (N_3749,N_2913,N_2362);
xnor U3750 (N_3750,N_2734,N_2639);
or U3751 (N_3751,N_2166,N_2207);
and U3752 (N_3752,N_1663,N_1549);
nor U3753 (N_3753,N_1707,N_2115);
nand U3754 (N_3754,N_2007,N_2462);
or U3755 (N_3755,N_1637,N_2237);
xnor U3756 (N_3756,N_2663,N_2150);
nor U3757 (N_3757,N_2203,N_2262);
nand U3758 (N_3758,N_2633,N_1733);
and U3759 (N_3759,N_2021,N_1627);
nand U3760 (N_3760,N_1545,N_1810);
and U3761 (N_3761,N_2096,N_2916);
and U3762 (N_3762,N_2789,N_1766);
or U3763 (N_3763,N_1979,N_1953);
nor U3764 (N_3764,N_2527,N_2342);
xnor U3765 (N_3765,N_2110,N_2348);
xnor U3766 (N_3766,N_1676,N_1996);
nor U3767 (N_3767,N_2384,N_2959);
and U3768 (N_3768,N_2611,N_2387);
and U3769 (N_3769,N_2494,N_2874);
xnor U3770 (N_3770,N_2654,N_1790);
nor U3771 (N_3771,N_2994,N_1695);
nand U3772 (N_3772,N_2842,N_2873);
nor U3773 (N_3773,N_2329,N_2049);
nand U3774 (N_3774,N_2235,N_2700);
or U3775 (N_3775,N_2726,N_2525);
xor U3776 (N_3776,N_2336,N_2741);
nand U3777 (N_3777,N_2112,N_2338);
nor U3778 (N_3778,N_2232,N_1663);
nand U3779 (N_3779,N_1517,N_1516);
nor U3780 (N_3780,N_2738,N_1650);
nor U3781 (N_3781,N_1718,N_2763);
or U3782 (N_3782,N_2569,N_2620);
nand U3783 (N_3783,N_1580,N_2928);
xor U3784 (N_3784,N_1733,N_1819);
or U3785 (N_3785,N_1709,N_2198);
and U3786 (N_3786,N_1636,N_2055);
nand U3787 (N_3787,N_1768,N_1519);
nor U3788 (N_3788,N_2673,N_2981);
nand U3789 (N_3789,N_2509,N_1872);
xor U3790 (N_3790,N_2224,N_2328);
xnor U3791 (N_3791,N_2558,N_1751);
or U3792 (N_3792,N_2567,N_1809);
or U3793 (N_3793,N_2599,N_1916);
or U3794 (N_3794,N_1572,N_2967);
xnor U3795 (N_3795,N_2297,N_2065);
or U3796 (N_3796,N_2571,N_2760);
nor U3797 (N_3797,N_2474,N_2017);
and U3798 (N_3798,N_2041,N_2220);
or U3799 (N_3799,N_2431,N_2614);
and U3800 (N_3800,N_2628,N_1933);
nor U3801 (N_3801,N_2633,N_2987);
nor U3802 (N_3802,N_2774,N_1704);
nor U3803 (N_3803,N_2719,N_2173);
or U3804 (N_3804,N_2176,N_2877);
and U3805 (N_3805,N_1778,N_1825);
or U3806 (N_3806,N_2997,N_1500);
nand U3807 (N_3807,N_1951,N_2972);
nor U3808 (N_3808,N_2116,N_1814);
nand U3809 (N_3809,N_1956,N_1959);
xor U3810 (N_3810,N_1557,N_1537);
and U3811 (N_3811,N_2422,N_2639);
xnor U3812 (N_3812,N_2165,N_1517);
xnor U3813 (N_3813,N_2029,N_1825);
and U3814 (N_3814,N_2985,N_2375);
nand U3815 (N_3815,N_2317,N_2924);
nor U3816 (N_3816,N_2383,N_2505);
and U3817 (N_3817,N_2940,N_2580);
or U3818 (N_3818,N_1589,N_2801);
nor U3819 (N_3819,N_2737,N_2586);
or U3820 (N_3820,N_2996,N_1712);
nand U3821 (N_3821,N_2256,N_2144);
nand U3822 (N_3822,N_2718,N_1671);
nor U3823 (N_3823,N_2698,N_1721);
nor U3824 (N_3824,N_1584,N_2717);
or U3825 (N_3825,N_1706,N_1887);
nand U3826 (N_3826,N_2387,N_1565);
and U3827 (N_3827,N_1593,N_2649);
xor U3828 (N_3828,N_2812,N_1886);
and U3829 (N_3829,N_1532,N_1926);
xor U3830 (N_3830,N_2944,N_2320);
xor U3831 (N_3831,N_2926,N_2249);
xnor U3832 (N_3832,N_2056,N_1628);
nor U3833 (N_3833,N_1918,N_1948);
nor U3834 (N_3834,N_1769,N_2892);
and U3835 (N_3835,N_2629,N_2921);
or U3836 (N_3836,N_2873,N_1791);
or U3837 (N_3837,N_1915,N_2921);
xnor U3838 (N_3838,N_1883,N_2045);
or U3839 (N_3839,N_2858,N_2654);
xor U3840 (N_3840,N_2214,N_2047);
or U3841 (N_3841,N_2090,N_2171);
or U3842 (N_3842,N_2764,N_1644);
xnor U3843 (N_3843,N_1689,N_2176);
or U3844 (N_3844,N_2527,N_1812);
and U3845 (N_3845,N_2683,N_2164);
or U3846 (N_3846,N_1697,N_2272);
and U3847 (N_3847,N_2359,N_2881);
and U3848 (N_3848,N_2474,N_1890);
nor U3849 (N_3849,N_2947,N_2959);
nand U3850 (N_3850,N_2221,N_2585);
nor U3851 (N_3851,N_2539,N_1915);
or U3852 (N_3852,N_2452,N_1555);
nor U3853 (N_3853,N_2550,N_1810);
nand U3854 (N_3854,N_2537,N_2411);
or U3855 (N_3855,N_2846,N_2569);
nand U3856 (N_3856,N_2591,N_2174);
nand U3857 (N_3857,N_1818,N_1957);
nor U3858 (N_3858,N_2451,N_1724);
or U3859 (N_3859,N_1505,N_2242);
nand U3860 (N_3860,N_2214,N_2966);
or U3861 (N_3861,N_1738,N_2319);
xor U3862 (N_3862,N_1599,N_2007);
and U3863 (N_3863,N_1617,N_2987);
nand U3864 (N_3864,N_1828,N_2443);
and U3865 (N_3865,N_2303,N_2465);
xor U3866 (N_3866,N_2908,N_2436);
xor U3867 (N_3867,N_1667,N_1701);
or U3868 (N_3868,N_2777,N_2316);
nor U3869 (N_3869,N_1826,N_2537);
xor U3870 (N_3870,N_2722,N_1835);
nor U3871 (N_3871,N_1824,N_2088);
and U3872 (N_3872,N_2911,N_2400);
and U3873 (N_3873,N_1853,N_2292);
or U3874 (N_3874,N_2811,N_2647);
nor U3875 (N_3875,N_2367,N_2542);
and U3876 (N_3876,N_1861,N_2889);
or U3877 (N_3877,N_1629,N_1616);
or U3878 (N_3878,N_2730,N_1734);
xnor U3879 (N_3879,N_1514,N_2506);
nand U3880 (N_3880,N_2446,N_2360);
xor U3881 (N_3881,N_1529,N_1720);
xor U3882 (N_3882,N_1646,N_2118);
or U3883 (N_3883,N_2922,N_2603);
xnor U3884 (N_3884,N_2939,N_2820);
or U3885 (N_3885,N_1555,N_2757);
and U3886 (N_3886,N_1536,N_2451);
or U3887 (N_3887,N_2911,N_2053);
nor U3888 (N_3888,N_1863,N_1532);
or U3889 (N_3889,N_1515,N_2917);
xor U3890 (N_3890,N_1695,N_2607);
nor U3891 (N_3891,N_1613,N_2670);
nor U3892 (N_3892,N_2800,N_2171);
nor U3893 (N_3893,N_2228,N_1971);
nand U3894 (N_3894,N_1809,N_2131);
xnor U3895 (N_3895,N_2775,N_1555);
nand U3896 (N_3896,N_1621,N_2202);
or U3897 (N_3897,N_1878,N_2456);
or U3898 (N_3898,N_2738,N_1616);
xor U3899 (N_3899,N_2873,N_2572);
nand U3900 (N_3900,N_2756,N_2398);
nor U3901 (N_3901,N_2957,N_1824);
nor U3902 (N_3902,N_2612,N_2899);
and U3903 (N_3903,N_2246,N_2319);
and U3904 (N_3904,N_2344,N_2049);
nand U3905 (N_3905,N_1554,N_2198);
xnor U3906 (N_3906,N_2208,N_2247);
and U3907 (N_3907,N_1910,N_1746);
xnor U3908 (N_3908,N_2082,N_2028);
or U3909 (N_3909,N_2249,N_1904);
nand U3910 (N_3910,N_2439,N_1674);
nand U3911 (N_3911,N_1868,N_2056);
and U3912 (N_3912,N_2185,N_2776);
nand U3913 (N_3913,N_2966,N_1722);
xor U3914 (N_3914,N_1955,N_2865);
and U3915 (N_3915,N_1698,N_1687);
and U3916 (N_3916,N_1683,N_2288);
xor U3917 (N_3917,N_2650,N_1747);
nor U3918 (N_3918,N_1871,N_2205);
and U3919 (N_3919,N_2975,N_2752);
or U3920 (N_3920,N_1621,N_2051);
xnor U3921 (N_3921,N_1744,N_2696);
or U3922 (N_3922,N_1565,N_2292);
nand U3923 (N_3923,N_1565,N_2095);
and U3924 (N_3924,N_2749,N_1841);
nor U3925 (N_3925,N_2203,N_2966);
nand U3926 (N_3926,N_1543,N_1820);
and U3927 (N_3927,N_2234,N_2053);
xor U3928 (N_3928,N_1571,N_1514);
nor U3929 (N_3929,N_2800,N_2256);
nand U3930 (N_3930,N_2920,N_1838);
xnor U3931 (N_3931,N_2398,N_1668);
nor U3932 (N_3932,N_2547,N_2962);
nor U3933 (N_3933,N_1998,N_2487);
nor U3934 (N_3934,N_2173,N_2079);
and U3935 (N_3935,N_1536,N_2233);
nand U3936 (N_3936,N_1574,N_1830);
nor U3937 (N_3937,N_2041,N_2067);
or U3938 (N_3938,N_2784,N_2774);
nand U3939 (N_3939,N_2369,N_1894);
or U3940 (N_3940,N_2605,N_2926);
nand U3941 (N_3941,N_2308,N_1982);
and U3942 (N_3942,N_1836,N_2670);
or U3943 (N_3943,N_2622,N_2531);
nor U3944 (N_3944,N_1564,N_2295);
xnor U3945 (N_3945,N_2495,N_1821);
nand U3946 (N_3946,N_2592,N_2937);
and U3947 (N_3947,N_1670,N_2741);
nor U3948 (N_3948,N_1725,N_1918);
nor U3949 (N_3949,N_1703,N_1704);
and U3950 (N_3950,N_2159,N_1787);
xnor U3951 (N_3951,N_2137,N_2338);
xnor U3952 (N_3952,N_1592,N_2008);
xor U3953 (N_3953,N_1800,N_2097);
nand U3954 (N_3954,N_2419,N_2669);
nor U3955 (N_3955,N_2387,N_2077);
or U3956 (N_3956,N_2079,N_1519);
nor U3957 (N_3957,N_2827,N_2998);
xnor U3958 (N_3958,N_2996,N_2399);
or U3959 (N_3959,N_1884,N_2918);
or U3960 (N_3960,N_2353,N_1787);
xor U3961 (N_3961,N_2947,N_2634);
xnor U3962 (N_3962,N_1597,N_2014);
nor U3963 (N_3963,N_2605,N_2577);
nor U3964 (N_3964,N_2717,N_2161);
and U3965 (N_3965,N_2093,N_1617);
xnor U3966 (N_3966,N_2990,N_1640);
and U3967 (N_3967,N_1602,N_2588);
xor U3968 (N_3968,N_2103,N_2482);
or U3969 (N_3969,N_1726,N_1521);
and U3970 (N_3970,N_1681,N_1632);
and U3971 (N_3971,N_1962,N_1963);
xnor U3972 (N_3972,N_2444,N_2473);
nand U3973 (N_3973,N_1681,N_2902);
or U3974 (N_3974,N_2665,N_1773);
or U3975 (N_3975,N_2966,N_1642);
xor U3976 (N_3976,N_1671,N_2181);
or U3977 (N_3977,N_2952,N_2215);
nand U3978 (N_3978,N_2171,N_1802);
and U3979 (N_3979,N_2026,N_1824);
xnor U3980 (N_3980,N_1883,N_2883);
nand U3981 (N_3981,N_2572,N_2859);
and U3982 (N_3982,N_1962,N_2219);
nor U3983 (N_3983,N_1921,N_2913);
xor U3984 (N_3984,N_2653,N_2540);
nand U3985 (N_3985,N_2183,N_2327);
xnor U3986 (N_3986,N_2725,N_2084);
nor U3987 (N_3987,N_1990,N_1526);
or U3988 (N_3988,N_1887,N_2862);
xnor U3989 (N_3989,N_2353,N_2799);
or U3990 (N_3990,N_2101,N_2940);
or U3991 (N_3991,N_2817,N_1632);
or U3992 (N_3992,N_2315,N_1889);
and U3993 (N_3993,N_2632,N_2678);
xor U3994 (N_3994,N_2589,N_1942);
and U3995 (N_3995,N_2862,N_2641);
or U3996 (N_3996,N_2922,N_1688);
and U3997 (N_3997,N_2701,N_2975);
nor U3998 (N_3998,N_2784,N_2595);
xor U3999 (N_3999,N_2695,N_2443);
or U4000 (N_4000,N_2917,N_2418);
or U4001 (N_4001,N_1658,N_2428);
nand U4002 (N_4002,N_2420,N_2276);
nor U4003 (N_4003,N_2419,N_1892);
nand U4004 (N_4004,N_2822,N_1792);
and U4005 (N_4005,N_2927,N_1747);
nor U4006 (N_4006,N_2534,N_1588);
nand U4007 (N_4007,N_1741,N_2691);
xnor U4008 (N_4008,N_2911,N_2943);
nor U4009 (N_4009,N_2232,N_1628);
or U4010 (N_4010,N_2952,N_2357);
nand U4011 (N_4011,N_2313,N_2709);
xnor U4012 (N_4012,N_1944,N_2525);
xnor U4013 (N_4013,N_2860,N_2850);
or U4014 (N_4014,N_2591,N_1656);
xnor U4015 (N_4015,N_2049,N_2652);
nand U4016 (N_4016,N_1610,N_2664);
xor U4017 (N_4017,N_2891,N_1665);
and U4018 (N_4018,N_2690,N_2009);
nor U4019 (N_4019,N_1881,N_1834);
xor U4020 (N_4020,N_1888,N_2251);
nor U4021 (N_4021,N_2531,N_2200);
or U4022 (N_4022,N_1944,N_2920);
nand U4023 (N_4023,N_2887,N_1664);
nand U4024 (N_4024,N_2139,N_2118);
nand U4025 (N_4025,N_1589,N_1837);
nand U4026 (N_4026,N_2496,N_1971);
nor U4027 (N_4027,N_2992,N_2151);
and U4028 (N_4028,N_1571,N_1661);
and U4029 (N_4029,N_2029,N_2615);
or U4030 (N_4030,N_2830,N_2794);
nand U4031 (N_4031,N_2578,N_2436);
and U4032 (N_4032,N_1975,N_2939);
or U4033 (N_4033,N_1923,N_2241);
nand U4034 (N_4034,N_2874,N_2433);
nor U4035 (N_4035,N_2735,N_1915);
and U4036 (N_4036,N_2636,N_2102);
nor U4037 (N_4037,N_2807,N_2907);
nand U4038 (N_4038,N_1850,N_2994);
nand U4039 (N_4039,N_2149,N_2223);
and U4040 (N_4040,N_2714,N_1891);
nand U4041 (N_4041,N_2527,N_1580);
or U4042 (N_4042,N_2246,N_2058);
or U4043 (N_4043,N_1658,N_2640);
nor U4044 (N_4044,N_1595,N_1548);
and U4045 (N_4045,N_2422,N_2282);
nand U4046 (N_4046,N_2820,N_1719);
or U4047 (N_4047,N_2861,N_1534);
and U4048 (N_4048,N_1512,N_1771);
and U4049 (N_4049,N_2476,N_2267);
nor U4050 (N_4050,N_1864,N_2338);
nor U4051 (N_4051,N_2442,N_1750);
nand U4052 (N_4052,N_1942,N_2917);
nand U4053 (N_4053,N_2541,N_2468);
and U4054 (N_4054,N_1551,N_2617);
nand U4055 (N_4055,N_1799,N_2406);
nand U4056 (N_4056,N_2402,N_2200);
nor U4057 (N_4057,N_2101,N_2312);
xor U4058 (N_4058,N_1613,N_1803);
or U4059 (N_4059,N_2548,N_2903);
xor U4060 (N_4060,N_2487,N_1790);
xor U4061 (N_4061,N_2811,N_2766);
and U4062 (N_4062,N_1697,N_1815);
nor U4063 (N_4063,N_2237,N_1874);
xnor U4064 (N_4064,N_2150,N_1897);
or U4065 (N_4065,N_2559,N_1655);
nand U4066 (N_4066,N_2821,N_2465);
xor U4067 (N_4067,N_2125,N_2111);
xnor U4068 (N_4068,N_1611,N_1622);
and U4069 (N_4069,N_2148,N_1686);
or U4070 (N_4070,N_1624,N_2738);
xor U4071 (N_4071,N_2170,N_1960);
xor U4072 (N_4072,N_2501,N_2368);
and U4073 (N_4073,N_2478,N_1520);
or U4074 (N_4074,N_2345,N_2964);
nand U4075 (N_4075,N_2601,N_2063);
or U4076 (N_4076,N_1891,N_1687);
nor U4077 (N_4077,N_2240,N_1514);
and U4078 (N_4078,N_2821,N_2512);
or U4079 (N_4079,N_2863,N_2758);
xor U4080 (N_4080,N_1861,N_2485);
xnor U4081 (N_4081,N_1759,N_2288);
nor U4082 (N_4082,N_2251,N_1707);
xnor U4083 (N_4083,N_2044,N_2148);
xnor U4084 (N_4084,N_2872,N_2982);
xnor U4085 (N_4085,N_2796,N_1731);
nand U4086 (N_4086,N_2746,N_2337);
xor U4087 (N_4087,N_1638,N_1650);
nor U4088 (N_4088,N_2114,N_2564);
and U4089 (N_4089,N_1548,N_2778);
xor U4090 (N_4090,N_2252,N_1932);
nand U4091 (N_4091,N_1642,N_1501);
nand U4092 (N_4092,N_1583,N_2590);
and U4093 (N_4093,N_2096,N_1511);
nand U4094 (N_4094,N_1932,N_2879);
nor U4095 (N_4095,N_2545,N_2618);
or U4096 (N_4096,N_1523,N_2674);
or U4097 (N_4097,N_2650,N_2262);
nor U4098 (N_4098,N_2874,N_1579);
or U4099 (N_4099,N_2347,N_2576);
or U4100 (N_4100,N_2659,N_2331);
nand U4101 (N_4101,N_2042,N_1563);
xor U4102 (N_4102,N_1647,N_2956);
or U4103 (N_4103,N_2882,N_1760);
or U4104 (N_4104,N_2607,N_2536);
xor U4105 (N_4105,N_1701,N_1997);
or U4106 (N_4106,N_1675,N_1902);
and U4107 (N_4107,N_2206,N_2089);
xor U4108 (N_4108,N_2415,N_2485);
xor U4109 (N_4109,N_2442,N_1935);
xor U4110 (N_4110,N_1831,N_1863);
nor U4111 (N_4111,N_1686,N_2033);
and U4112 (N_4112,N_2551,N_2272);
nand U4113 (N_4113,N_1813,N_1672);
xor U4114 (N_4114,N_2945,N_2383);
nor U4115 (N_4115,N_2314,N_2914);
nor U4116 (N_4116,N_2059,N_1811);
nor U4117 (N_4117,N_2964,N_1989);
xnor U4118 (N_4118,N_1703,N_2904);
xor U4119 (N_4119,N_1894,N_1931);
nor U4120 (N_4120,N_2404,N_2516);
nand U4121 (N_4121,N_1866,N_2251);
and U4122 (N_4122,N_1848,N_2256);
and U4123 (N_4123,N_2251,N_2983);
xor U4124 (N_4124,N_2976,N_1796);
and U4125 (N_4125,N_1644,N_1680);
and U4126 (N_4126,N_1573,N_2492);
xnor U4127 (N_4127,N_2653,N_2087);
and U4128 (N_4128,N_2384,N_2693);
or U4129 (N_4129,N_2173,N_1548);
and U4130 (N_4130,N_2201,N_1642);
nand U4131 (N_4131,N_1739,N_2181);
nand U4132 (N_4132,N_2843,N_1751);
or U4133 (N_4133,N_2392,N_2527);
nand U4134 (N_4134,N_1763,N_2759);
xor U4135 (N_4135,N_1798,N_2766);
nand U4136 (N_4136,N_2007,N_1869);
nand U4137 (N_4137,N_2249,N_2426);
and U4138 (N_4138,N_1663,N_1806);
nor U4139 (N_4139,N_2768,N_2227);
or U4140 (N_4140,N_1836,N_2491);
or U4141 (N_4141,N_2432,N_2806);
and U4142 (N_4142,N_1973,N_1658);
nor U4143 (N_4143,N_1738,N_2212);
and U4144 (N_4144,N_1582,N_1668);
xor U4145 (N_4145,N_2832,N_2326);
or U4146 (N_4146,N_1591,N_1578);
and U4147 (N_4147,N_2887,N_2306);
or U4148 (N_4148,N_2751,N_2056);
nor U4149 (N_4149,N_1919,N_2513);
and U4150 (N_4150,N_2807,N_1597);
or U4151 (N_4151,N_2475,N_2415);
or U4152 (N_4152,N_1883,N_1590);
and U4153 (N_4153,N_2134,N_2046);
xnor U4154 (N_4154,N_1586,N_2008);
nand U4155 (N_4155,N_1767,N_2707);
xor U4156 (N_4156,N_2430,N_2690);
xnor U4157 (N_4157,N_1777,N_2088);
nand U4158 (N_4158,N_2699,N_2376);
and U4159 (N_4159,N_1840,N_2863);
xor U4160 (N_4160,N_2798,N_2574);
xor U4161 (N_4161,N_2297,N_2897);
nand U4162 (N_4162,N_1558,N_1607);
xor U4163 (N_4163,N_2715,N_2641);
and U4164 (N_4164,N_2802,N_1817);
nor U4165 (N_4165,N_2470,N_1821);
nand U4166 (N_4166,N_1771,N_2009);
and U4167 (N_4167,N_2370,N_2899);
xor U4168 (N_4168,N_1935,N_1940);
nand U4169 (N_4169,N_2419,N_2790);
xor U4170 (N_4170,N_2626,N_2602);
and U4171 (N_4171,N_1624,N_2130);
or U4172 (N_4172,N_2670,N_1522);
and U4173 (N_4173,N_1772,N_2955);
nand U4174 (N_4174,N_1782,N_2443);
or U4175 (N_4175,N_2908,N_2621);
xnor U4176 (N_4176,N_1720,N_2573);
and U4177 (N_4177,N_2866,N_2939);
xnor U4178 (N_4178,N_2030,N_1637);
or U4179 (N_4179,N_2576,N_1543);
and U4180 (N_4180,N_1808,N_2328);
and U4181 (N_4181,N_2608,N_2746);
and U4182 (N_4182,N_1576,N_1832);
nor U4183 (N_4183,N_1601,N_2494);
xnor U4184 (N_4184,N_1568,N_2169);
nor U4185 (N_4185,N_2617,N_1613);
or U4186 (N_4186,N_2997,N_2947);
nand U4187 (N_4187,N_2057,N_2605);
nand U4188 (N_4188,N_2398,N_1887);
nand U4189 (N_4189,N_1552,N_2806);
nand U4190 (N_4190,N_2068,N_2341);
xor U4191 (N_4191,N_2266,N_1907);
xor U4192 (N_4192,N_1957,N_2900);
or U4193 (N_4193,N_1587,N_1674);
and U4194 (N_4194,N_1743,N_1878);
or U4195 (N_4195,N_2535,N_2813);
nand U4196 (N_4196,N_2031,N_2277);
and U4197 (N_4197,N_2876,N_1957);
xnor U4198 (N_4198,N_2425,N_2115);
xnor U4199 (N_4199,N_2519,N_2640);
and U4200 (N_4200,N_1935,N_1654);
and U4201 (N_4201,N_2981,N_2045);
nor U4202 (N_4202,N_2186,N_2520);
xor U4203 (N_4203,N_1828,N_2714);
or U4204 (N_4204,N_2704,N_1812);
and U4205 (N_4205,N_1911,N_2201);
or U4206 (N_4206,N_2978,N_2794);
nor U4207 (N_4207,N_2447,N_2772);
xnor U4208 (N_4208,N_2415,N_1618);
and U4209 (N_4209,N_2119,N_2232);
xnor U4210 (N_4210,N_1832,N_2742);
xnor U4211 (N_4211,N_1991,N_1612);
nand U4212 (N_4212,N_2385,N_2999);
xor U4213 (N_4213,N_2539,N_2641);
or U4214 (N_4214,N_1878,N_2775);
xor U4215 (N_4215,N_1820,N_2853);
and U4216 (N_4216,N_1531,N_2685);
xnor U4217 (N_4217,N_2175,N_1624);
nor U4218 (N_4218,N_2874,N_2028);
and U4219 (N_4219,N_1539,N_1995);
xnor U4220 (N_4220,N_2289,N_2332);
xnor U4221 (N_4221,N_2955,N_2005);
xor U4222 (N_4222,N_2337,N_2615);
and U4223 (N_4223,N_2809,N_2243);
nand U4224 (N_4224,N_2508,N_2080);
nor U4225 (N_4225,N_1525,N_2672);
nand U4226 (N_4226,N_1707,N_1876);
xnor U4227 (N_4227,N_2411,N_1604);
nand U4228 (N_4228,N_2136,N_2636);
and U4229 (N_4229,N_2922,N_1668);
nand U4230 (N_4230,N_1908,N_1691);
nor U4231 (N_4231,N_1590,N_2218);
nor U4232 (N_4232,N_2627,N_2810);
or U4233 (N_4233,N_1627,N_2784);
and U4234 (N_4234,N_1957,N_2910);
nand U4235 (N_4235,N_2640,N_1621);
and U4236 (N_4236,N_1612,N_2817);
xor U4237 (N_4237,N_2430,N_2501);
xnor U4238 (N_4238,N_2666,N_1705);
nand U4239 (N_4239,N_2846,N_2698);
nand U4240 (N_4240,N_2680,N_2575);
or U4241 (N_4241,N_2786,N_2591);
xnor U4242 (N_4242,N_2635,N_2291);
nand U4243 (N_4243,N_2854,N_2200);
xor U4244 (N_4244,N_1946,N_2575);
and U4245 (N_4245,N_2485,N_2976);
xor U4246 (N_4246,N_2198,N_1603);
and U4247 (N_4247,N_2578,N_1589);
xnor U4248 (N_4248,N_2556,N_2133);
nor U4249 (N_4249,N_1840,N_2437);
nand U4250 (N_4250,N_2919,N_1859);
nor U4251 (N_4251,N_1552,N_1894);
xnor U4252 (N_4252,N_2557,N_2158);
nand U4253 (N_4253,N_2297,N_2399);
or U4254 (N_4254,N_2658,N_2741);
nor U4255 (N_4255,N_2423,N_1616);
xor U4256 (N_4256,N_1737,N_2540);
or U4257 (N_4257,N_2711,N_2022);
and U4258 (N_4258,N_2354,N_2953);
or U4259 (N_4259,N_2935,N_2367);
nor U4260 (N_4260,N_2053,N_2902);
and U4261 (N_4261,N_1852,N_1534);
nor U4262 (N_4262,N_1905,N_2303);
nor U4263 (N_4263,N_1927,N_2786);
and U4264 (N_4264,N_2403,N_1885);
nor U4265 (N_4265,N_2750,N_1676);
nor U4266 (N_4266,N_1997,N_2751);
and U4267 (N_4267,N_1798,N_2433);
or U4268 (N_4268,N_2455,N_1859);
and U4269 (N_4269,N_2429,N_2732);
nand U4270 (N_4270,N_2768,N_2851);
nor U4271 (N_4271,N_2729,N_2606);
and U4272 (N_4272,N_2533,N_2929);
xnor U4273 (N_4273,N_2806,N_1612);
or U4274 (N_4274,N_1928,N_1528);
nand U4275 (N_4275,N_1827,N_2247);
or U4276 (N_4276,N_1517,N_2734);
nand U4277 (N_4277,N_1525,N_2715);
nand U4278 (N_4278,N_2356,N_2914);
and U4279 (N_4279,N_1841,N_1749);
nor U4280 (N_4280,N_1781,N_2115);
nand U4281 (N_4281,N_2462,N_2122);
and U4282 (N_4282,N_2685,N_2637);
and U4283 (N_4283,N_2869,N_1529);
and U4284 (N_4284,N_2377,N_1785);
nor U4285 (N_4285,N_1607,N_2900);
or U4286 (N_4286,N_2093,N_1831);
and U4287 (N_4287,N_2139,N_2781);
and U4288 (N_4288,N_2929,N_2536);
xor U4289 (N_4289,N_2434,N_2745);
and U4290 (N_4290,N_2491,N_2916);
nor U4291 (N_4291,N_2056,N_2404);
or U4292 (N_4292,N_2439,N_1648);
and U4293 (N_4293,N_1763,N_2297);
nor U4294 (N_4294,N_2032,N_2141);
and U4295 (N_4295,N_2227,N_1571);
xnor U4296 (N_4296,N_2045,N_2667);
xor U4297 (N_4297,N_2913,N_2583);
xor U4298 (N_4298,N_1878,N_1608);
or U4299 (N_4299,N_2756,N_2126);
and U4300 (N_4300,N_1588,N_1716);
xnor U4301 (N_4301,N_1849,N_2948);
and U4302 (N_4302,N_2418,N_2213);
and U4303 (N_4303,N_1642,N_2563);
or U4304 (N_4304,N_1601,N_1791);
xnor U4305 (N_4305,N_2698,N_2961);
xnor U4306 (N_4306,N_2585,N_2706);
xor U4307 (N_4307,N_2462,N_2944);
or U4308 (N_4308,N_2582,N_2243);
and U4309 (N_4309,N_2408,N_1745);
nand U4310 (N_4310,N_2061,N_2423);
xor U4311 (N_4311,N_2847,N_2059);
xnor U4312 (N_4312,N_1991,N_1685);
or U4313 (N_4313,N_2607,N_2937);
and U4314 (N_4314,N_1568,N_2089);
and U4315 (N_4315,N_1764,N_2808);
xnor U4316 (N_4316,N_2611,N_1503);
nand U4317 (N_4317,N_1874,N_2677);
or U4318 (N_4318,N_2837,N_2545);
xnor U4319 (N_4319,N_1698,N_2597);
or U4320 (N_4320,N_1533,N_2372);
xor U4321 (N_4321,N_2044,N_2447);
or U4322 (N_4322,N_2568,N_2747);
nor U4323 (N_4323,N_2779,N_2296);
xnor U4324 (N_4324,N_2862,N_2537);
xor U4325 (N_4325,N_2518,N_1567);
nor U4326 (N_4326,N_2543,N_2080);
and U4327 (N_4327,N_2548,N_2012);
and U4328 (N_4328,N_2941,N_1833);
and U4329 (N_4329,N_2496,N_2299);
and U4330 (N_4330,N_1525,N_2882);
nand U4331 (N_4331,N_2678,N_2829);
nand U4332 (N_4332,N_1664,N_2286);
or U4333 (N_4333,N_2663,N_2751);
xor U4334 (N_4334,N_2878,N_2103);
or U4335 (N_4335,N_2981,N_2427);
or U4336 (N_4336,N_1557,N_2867);
nand U4337 (N_4337,N_2488,N_2854);
or U4338 (N_4338,N_2340,N_1736);
nor U4339 (N_4339,N_2550,N_2244);
or U4340 (N_4340,N_1796,N_2384);
and U4341 (N_4341,N_2920,N_2506);
nor U4342 (N_4342,N_2722,N_1721);
or U4343 (N_4343,N_1971,N_1687);
or U4344 (N_4344,N_2991,N_1783);
xnor U4345 (N_4345,N_1531,N_2617);
nor U4346 (N_4346,N_1631,N_2090);
and U4347 (N_4347,N_1742,N_2650);
xor U4348 (N_4348,N_1717,N_2807);
or U4349 (N_4349,N_2282,N_1910);
xor U4350 (N_4350,N_1634,N_2188);
and U4351 (N_4351,N_2412,N_2475);
nand U4352 (N_4352,N_1800,N_1938);
nor U4353 (N_4353,N_2588,N_2392);
nand U4354 (N_4354,N_1927,N_1926);
and U4355 (N_4355,N_2054,N_2358);
nand U4356 (N_4356,N_2134,N_2327);
xor U4357 (N_4357,N_2677,N_2546);
nand U4358 (N_4358,N_2608,N_1534);
nor U4359 (N_4359,N_1608,N_1914);
or U4360 (N_4360,N_2629,N_2239);
and U4361 (N_4361,N_2851,N_1923);
or U4362 (N_4362,N_2166,N_2579);
or U4363 (N_4363,N_2287,N_2047);
nor U4364 (N_4364,N_1749,N_1929);
xor U4365 (N_4365,N_2792,N_2155);
xor U4366 (N_4366,N_2608,N_1815);
nor U4367 (N_4367,N_2106,N_1684);
nor U4368 (N_4368,N_2242,N_2448);
and U4369 (N_4369,N_2639,N_1527);
or U4370 (N_4370,N_2740,N_1591);
or U4371 (N_4371,N_2305,N_1758);
or U4372 (N_4372,N_1633,N_1526);
nand U4373 (N_4373,N_2872,N_1682);
and U4374 (N_4374,N_2108,N_2340);
and U4375 (N_4375,N_2159,N_1826);
nor U4376 (N_4376,N_2594,N_1694);
xor U4377 (N_4377,N_2235,N_1508);
nor U4378 (N_4378,N_2627,N_2080);
and U4379 (N_4379,N_1674,N_1999);
nor U4380 (N_4380,N_2745,N_2144);
or U4381 (N_4381,N_2027,N_2181);
or U4382 (N_4382,N_1827,N_2929);
nor U4383 (N_4383,N_2511,N_1515);
and U4384 (N_4384,N_2028,N_1695);
and U4385 (N_4385,N_1884,N_2429);
and U4386 (N_4386,N_2441,N_2113);
xnor U4387 (N_4387,N_2781,N_2234);
or U4388 (N_4388,N_2674,N_2136);
and U4389 (N_4389,N_2857,N_1638);
or U4390 (N_4390,N_2787,N_2327);
or U4391 (N_4391,N_1825,N_2535);
nor U4392 (N_4392,N_2763,N_2304);
nor U4393 (N_4393,N_1743,N_2503);
and U4394 (N_4394,N_1584,N_2093);
and U4395 (N_4395,N_1620,N_1802);
and U4396 (N_4396,N_2110,N_2848);
xnor U4397 (N_4397,N_2962,N_2649);
xnor U4398 (N_4398,N_2096,N_2663);
nand U4399 (N_4399,N_1722,N_2033);
and U4400 (N_4400,N_2560,N_1567);
xnor U4401 (N_4401,N_1594,N_2371);
or U4402 (N_4402,N_2424,N_1969);
nor U4403 (N_4403,N_2768,N_2696);
nor U4404 (N_4404,N_2452,N_1913);
nand U4405 (N_4405,N_1543,N_1654);
xnor U4406 (N_4406,N_1546,N_2886);
or U4407 (N_4407,N_2481,N_1944);
nor U4408 (N_4408,N_1785,N_1660);
and U4409 (N_4409,N_1914,N_2453);
nand U4410 (N_4410,N_1879,N_2833);
or U4411 (N_4411,N_2710,N_2416);
and U4412 (N_4412,N_1834,N_2375);
nor U4413 (N_4413,N_2988,N_2281);
or U4414 (N_4414,N_2544,N_2666);
xnor U4415 (N_4415,N_2192,N_2357);
nand U4416 (N_4416,N_2784,N_2161);
xnor U4417 (N_4417,N_2975,N_1915);
nor U4418 (N_4418,N_2430,N_1674);
nor U4419 (N_4419,N_2640,N_2244);
or U4420 (N_4420,N_2947,N_1977);
or U4421 (N_4421,N_2910,N_2060);
nor U4422 (N_4422,N_2241,N_1510);
and U4423 (N_4423,N_2774,N_2550);
or U4424 (N_4424,N_2139,N_1776);
and U4425 (N_4425,N_1982,N_2191);
xnor U4426 (N_4426,N_1842,N_2584);
or U4427 (N_4427,N_1860,N_1895);
and U4428 (N_4428,N_2147,N_1754);
and U4429 (N_4429,N_1541,N_2457);
nand U4430 (N_4430,N_2674,N_1749);
nor U4431 (N_4431,N_2966,N_2388);
or U4432 (N_4432,N_2477,N_1775);
or U4433 (N_4433,N_1960,N_2215);
xnor U4434 (N_4434,N_2662,N_1862);
nor U4435 (N_4435,N_2743,N_2702);
nor U4436 (N_4436,N_2242,N_2762);
or U4437 (N_4437,N_2680,N_1698);
and U4438 (N_4438,N_1834,N_2529);
nand U4439 (N_4439,N_1547,N_1605);
xor U4440 (N_4440,N_2610,N_2699);
or U4441 (N_4441,N_2878,N_1520);
xor U4442 (N_4442,N_1912,N_2742);
xor U4443 (N_4443,N_2399,N_2899);
nor U4444 (N_4444,N_1763,N_1560);
nor U4445 (N_4445,N_2784,N_2840);
and U4446 (N_4446,N_2718,N_2400);
nand U4447 (N_4447,N_1525,N_2989);
xnor U4448 (N_4448,N_2132,N_1880);
nor U4449 (N_4449,N_2249,N_2448);
or U4450 (N_4450,N_2578,N_2243);
xor U4451 (N_4451,N_2351,N_2628);
nand U4452 (N_4452,N_2553,N_1811);
nand U4453 (N_4453,N_2815,N_1832);
or U4454 (N_4454,N_2083,N_2600);
and U4455 (N_4455,N_1918,N_2494);
or U4456 (N_4456,N_2630,N_2804);
xnor U4457 (N_4457,N_1821,N_2611);
nand U4458 (N_4458,N_1552,N_2878);
nor U4459 (N_4459,N_2626,N_1673);
nand U4460 (N_4460,N_2065,N_1749);
and U4461 (N_4461,N_1598,N_1503);
and U4462 (N_4462,N_2979,N_2288);
and U4463 (N_4463,N_1766,N_2155);
nand U4464 (N_4464,N_1898,N_2667);
nor U4465 (N_4465,N_2584,N_1916);
and U4466 (N_4466,N_1781,N_1532);
nor U4467 (N_4467,N_2358,N_1506);
xnor U4468 (N_4468,N_2367,N_1956);
xor U4469 (N_4469,N_2573,N_2564);
nand U4470 (N_4470,N_1954,N_2519);
or U4471 (N_4471,N_2277,N_2709);
nor U4472 (N_4472,N_2877,N_1530);
nand U4473 (N_4473,N_1776,N_1981);
xnor U4474 (N_4474,N_1985,N_2771);
or U4475 (N_4475,N_2391,N_2020);
nor U4476 (N_4476,N_2596,N_1743);
xnor U4477 (N_4477,N_1522,N_2052);
nor U4478 (N_4478,N_2709,N_1942);
nand U4479 (N_4479,N_2153,N_2140);
or U4480 (N_4480,N_2495,N_2254);
or U4481 (N_4481,N_2536,N_2055);
or U4482 (N_4482,N_2683,N_2687);
and U4483 (N_4483,N_2956,N_1903);
xor U4484 (N_4484,N_2159,N_1680);
and U4485 (N_4485,N_2750,N_2152);
xnor U4486 (N_4486,N_1881,N_2150);
or U4487 (N_4487,N_2419,N_1720);
or U4488 (N_4488,N_2542,N_1784);
nand U4489 (N_4489,N_1717,N_1656);
nor U4490 (N_4490,N_2236,N_2503);
and U4491 (N_4491,N_2519,N_1543);
xor U4492 (N_4492,N_2565,N_2208);
nand U4493 (N_4493,N_2418,N_2953);
nand U4494 (N_4494,N_2976,N_2637);
xor U4495 (N_4495,N_2664,N_2853);
nor U4496 (N_4496,N_1808,N_2608);
nand U4497 (N_4497,N_2188,N_1917);
nand U4498 (N_4498,N_2125,N_2979);
nand U4499 (N_4499,N_2586,N_2927);
nand U4500 (N_4500,N_3597,N_3053);
xnor U4501 (N_4501,N_4285,N_3767);
or U4502 (N_4502,N_3673,N_3244);
and U4503 (N_4503,N_4087,N_4219);
nor U4504 (N_4504,N_3562,N_3643);
nor U4505 (N_4505,N_3474,N_4128);
or U4506 (N_4506,N_3963,N_4191);
or U4507 (N_4507,N_3095,N_3699);
nor U4508 (N_4508,N_3152,N_4346);
nand U4509 (N_4509,N_3971,N_3674);
or U4510 (N_4510,N_3621,N_4214);
or U4511 (N_4511,N_3873,N_3956);
nor U4512 (N_4512,N_4218,N_3002);
nor U4513 (N_4513,N_3990,N_3602);
nor U4514 (N_4514,N_4321,N_4021);
or U4515 (N_4515,N_3126,N_4386);
or U4516 (N_4516,N_3202,N_3694);
nand U4517 (N_4517,N_3949,N_4116);
xor U4518 (N_4518,N_3294,N_3013);
or U4519 (N_4519,N_3731,N_3450);
or U4520 (N_4520,N_3286,N_4269);
or U4521 (N_4521,N_4223,N_4339);
or U4522 (N_4522,N_4075,N_4041);
or U4523 (N_4523,N_3018,N_3008);
nor U4524 (N_4524,N_3118,N_3044);
xnor U4525 (N_4525,N_4361,N_3498);
nor U4526 (N_4526,N_4394,N_3434);
xnor U4527 (N_4527,N_3556,N_4089);
or U4528 (N_4528,N_4497,N_3872);
xor U4529 (N_4529,N_3338,N_3882);
nor U4530 (N_4530,N_3136,N_3153);
and U4531 (N_4531,N_4084,N_4176);
nor U4532 (N_4532,N_3577,N_3783);
and U4533 (N_4533,N_3506,N_3780);
and U4534 (N_4534,N_4015,N_3850);
xor U4535 (N_4535,N_3930,N_3826);
or U4536 (N_4536,N_3446,N_4138);
nand U4537 (N_4537,N_3677,N_3661);
xnor U4538 (N_4538,N_3750,N_3361);
xnor U4539 (N_4539,N_3906,N_4039);
xor U4540 (N_4540,N_3158,N_3427);
and U4541 (N_4541,N_3140,N_4229);
nand U4542 (N_4542,N_3318,N_4452);
or U4543 (N_4543,N_4080,N_3776);
xor U4544 (N_4544,N_4451,N_3048);
nor U4545 (N_4545,N_4371,N_3966);
nor U4546 (N_4546,N_4294,N_3309);
and U4547 (N_4547,N_3821,N_3521);
nor U4548 (N_4548,N_3486,N_3571);
and U4549 (N_4549,N_3865,N_3142);
nor U4550 (N_4550,N_3638,N_3735);
or U4551 (N_4551,N_3669,N_3021);
xnor U4552 (N_4552,N_3372,N_4301);
nor U4553 (N_4553,N_4335,N_3995);
nand U4554 (N_4554,N_3250,N_3033);
nor U4555 (N_4555,N_3358,N_3066);
nor U4556 (N_4556,N_3631,N_4174);
xnor U4557 (N_4557,N_3998,N_3281);
xnor U4558 (N_4558,N_4184,N_3027);
or U4559 (N_4559,N_3500,N_3799);
xnor U4560 (N_4560,N_4125,N_3070);
xor U4561 (N_4561,N_4145,N_3374);
and U4562 (N_4562,N_4363,N_3404);
nand U4563 (N_4563,N_3005,N_3160);
and U4564 (N_4564,N_3311,N_4070);
and U4565 (N_4565,N_4434,N_4048);
nor U4566 (N_4566,N_3321,N_3977);
and U4567 (N_4567,N_3641,N_4444);
nand U4568 (N_4568,N_3259,N_4029);
nand U4569 (N_4569,N_3478,N_3364);
nor U4570 (N_4570,N_3700,N_3391);
nor U4571 (N_4571,N_4035,N_4281);
nor U4572 (N_4572,N_3415,N_4439);
nand U4573 (N_4573,N_3968,N_4430);
nand U4574 (N_4574,N_3993,N_4162);
xnor U4575 (N_4575,N_4000,N_3078);
xnor U4576 (N_4576,N_3749,N_4284);
and U4577 (N_4577,N_4494,N_4250);
xnor U4578 (N_4578,N_4073,N_4115);
nand U4579 (N_4579,N_3769,N_4256);
nand U4580 (N_4580,N_3130,N_4358);
xor U4581 (N_4581,N_3495,N_4493);
xor U4582 (N_4582,N_3085,N_3093);
nor U4583 (N_4583,N_3941,N_4207);
nand U4584 (N_4584,N_4387,N_4297);
nor U4585 (N_4585,N_3291,N_3802);
nand U4586 (N_4586,N_4094,N_3194);
and U4587 (N_4587,N_4401,N_4320);
or U4588 (N_4588,N_3473,N_3736);
xnor U4589 (N_4589,N_4330,N_4448);
or U4590 (N_4590,N_3649,N_3986);
xnor U4591 (N_4591,N_4283,N_3547);
and U4592 (N_4592,N_3241,N_4109);
nand U4593 (N_4593,N_3572,N_4274);
nor U4594 (N_4594,N_3333,N_4326);
and U4595 (N_4595,N_3324,N_3795);
nand U4596 (N_4596,N_4340,N_3067);
nand U4597 (N_4597,N_3386,N_4093);
or U4598 (N_4598,N_3718,N_3970);
nor U4599 (N_4599,N_3532,N_3658);
nor U4600 (N_4600,N_3617,N_3838);
or U4601 (N_4601,N_4032,N_3603);
xnor U4602 (N_4602,N_3646,N_4064);
nor U4603 (N_4603,N_4117,N_4054);
and U4604 (N_4604,N_3952,N_3740);
or U4605 (N_4605,N_3965,N_3744);
and U4606 (N_4606,N_3665,N_3756);
nand U4607 (N_4607,N_3509,N_3932);
xnor U4608 (N_4608,N_3245,N_3396);
or U4609 (N_4609,N_3787,N_3947);
xnor U4610 (N_4610,N_4423,N_3211);
xnor U4611 (N_4611,N_4013,N_3895);
and U4612 (N_4612,N_3090,N_3055);
xor U4613 (N_4613,N_4262,N_3558);
and U4614 (N_4614,N_4017,N_3465);
xnor U4615 (N_4615,N_3543,N_4275);
nand U4616 (N_4616,N_4183,N_3604);
nand U4617 (N_4617,N_3162,N_4239);
nand U4618 (N_4618,N_3133,N_3430);
nor U4619 (N_4619,N_4113,N_3908);
or U4620 (N_4620,N_3255,N_3796);
xnor U4621 (N_4621,N_3484,N_3851);
or U4622 (N_4622,N_3733,N_4243);
nor U4623 (N_4623,N_3452,N_3525);
or U4624 (N_4624,N_4022,N_4071);
nand U4625 (N_4625,N_3398,N_3269);
nand U4626 (N_4626,N_3809,N_3823);
nand U4627 (N_4627,N_4270,N_3905);
xnor U4628 (N_4628,N_3272,N_4111);
or U4629 (N_4629,N_3943,N_3278);
or U4630 (N_4630,N_4293,N_4486);
or U4631 (N_4631,N_4446,N_3931);
nor U4632 (N_4632,N_3719,N_3569);
or U4633 (N_4633,N_4136,N_3991);
xnor U4634 (N_4634,N_4466,N_3462);
or U4635 (N_4635,N_4004,N_3611);
nor U4636 (N_4636,N_4489,N_3605);
nand U4637 (N_4637,N_4034,N_3068);
xor U4638 (N_4638,N_3356,N_3794);
xnor U4639 (N_4639,N_3367,N_4478);
or U4640 (N_4640,N_3708,N_4171);
nand U4641 (N_4641,N_3504,N_3979);
xnor U4642 (N_4642,N_4158,N_3302);
or U4643 (N_4643,N_3343,N_4026);
nor U4644 (N_4644,N_4266,N_3325);
nand U4645 (N_4645,N_3359,N_3377);
and U4646 (N_4646,N_4336,N_4127);
nand U4647 (N_4647,N_3370,N_3188);
nor U4648 (N_4648,N_3079,N_4414);
and U4649 (N_4649,N_3154,N_4425);
xor U4650 (N_4650,N_3728,N_4043);
and U4651 (N_4651,N_4398,N_3151);
xnor U4652 (N_4652,N_3257,N_4259);
xor U4653 (N_4653,N_4118,N_4051);
nor U4654 (N_4654,N_3698,N_3322);
xnor U4655 (N_4655,N_4210,N_3805);
nand U4656 (N_4656,N_4147,N_4159);
and U4657 (N_4657,N_4213,N_4106);
nor U4658 (N_4658,N_4310,N_4231);
or U4659 (N_4659,N_3529,N_3655);
nand U4660 (N_4660,N_4272,N_3135);
or U4661 (N_4661,N_3179,N_4143);
nor U4662 (N_4662,N_4146,N_4167);
and U4663 (N_4663,N_3123,N_4357);
xor U4664 (N_4664,N_3493,N_3389);
xnor U4665 (N_4665,N_3094,N_3662);
nand U4666 (N_4666,N_3001,N_3014);
or U4667 (N_4667,N_3209,N_3258);
or U4668 (N_4668,N_3644,N_3976);
nor U4669 (N_4669,N_4066,N_3299);
or U4670 (N_4670,N_3582,N_3913);
nor U4671 (N_4671,N_3835,N_3900);
nor U4672 (N_4672,N_3782,N_4324);
or U4673 (N_4673,N_3683,N_3688);
xor U4674 (N_4674,N_4186,N_4194);
and U4675 (N_4675,N_3435,N_3307);
or U4676 (N_4676,N_4247,N_4236);
nand U4677 (N_4677,N_3992,N_4288);
xnor U4678 (N_4678,N_3166,N_4433);
nand U4679 (N_4679,N_3748,N_3693);
nand U4680 (N_4680,N_3394,N_3598);
nor U4681 (N_4681,N_3100,N_3980);
nor U4682 (N_4682,N_3513,N_3867);
xor U4683 (N_4683,N_3354,N_3552);
and U4684 (N_4684,N_4226,N_4488);
or U4685 (N_4685,N_3612,N_3475);
nor U4686 (N_4686,N_3472,N_3401);
nor U4687 (N_4687,N_3113,N_4142);
and U4688 (N_4688,N_4056,N_4251);
nand U4689 (N_4689,N_3149,N_3650);
nor U4690 (N_4690,N_3104,N_4144);
and U4691 (N_4691,N_3029,N_3116);
nand U4692 (N_4692,N_3634,N_4232);
xor U4693 (N_4693,N_4141,N_3304);
or U4694 (N_4694,N_4360,N_4173);
and U4695 (N_4695,N_3248,N_3148);
nor U4696 (N_4696,N_3530,N_3360);
or U4697 (N_4697,N_3606,N_3449);
nand U4698 (N_4698,N_4457,N_4382);
nor U4699 (N_4699,N_3216,N_4437);
xnor U4700 (N_4700,N_4168,N_4291);
nand U4701 (N_4701,N_3228,N_3551);
or U4702 (N_4702,N_3349,N_3168);
xnor U4703 (N_4703,N_3199,N_4241);
nor U4704 (N_4704,N_3645,N_3635);
nand U4705 (N_4705,N_3889,N_4307);
or U4706 (N_4706,N_3408,N_4190);
xor U4707 (N_4707,N_3538,N_4422);
nand U4708 (N_4708,N_3798,N_4295);
and U4709 (N_4709,N_3219,N_3315);
and U4710 (N_4710,N_3494,N_3978);
or U4711 (N_4711,N_3592,N_4216);
or U4712 (N_4712,N_4345,N_3923);
or U4713 (N_4713,N_4028,N_3549);
nand U4714 (N_4714,N_3870,N_4354);
nand U4715 (N_4715,N_3666,N_3576);
nor U4716 (N_4716,N_3040,N_3006);
nor U4717 (N_4717,N_3955,N_3487);
nand U4718 (N_4718,N_4428,N_3758);
and U4719 (N_4719,N_4060,N_3050);
nor U4720 (N_4720,N_3550,N_4476);
xor U4721 (N_4721,N_3935,N_3784);
xor U4722 (N_4722,N_3911,N_3668);
and U4723 (N_4723,N_3839,N_3405);
nor U4724 (N_4724,N_4456,N_3218);
and U4725 (N_4725,N_3157,N_3523);
xor U4726 (N_4726,N_3766,N_3035);
nand U4727 (N_4727,N_4419,N_3418);
or U4728 (N_4728,N_3200,N_4323);
xor U4729 (N_4729,N_3036,N_3887);
nand U4730 (N_4730,N_4040,N_3566);
nor U4731 (N_4731,N_3378,N_3103);
and U4732 (N_4732,N_4472,N_3489);
xnor U4733 (N_4733,N_3178,N_3287);
or U4734 (N_4734,N_3071,N_3579);
nor U4735 (N_4735,N_4140,N_4083);
nand U4736 (N_4736,N_4078,N_3648);
nand U4737 (N_4737,N_3413,N_3351);
nor U4738 (N_4738,N_3402,N_3266);
xor U4739 (N_4739,N_3410,N_3857);
nor U4740 (N_4740,N_3681,N_4192);
xor U4741 (N_4741,N_3928,N_4156);
nand U4742 (N_4742,N_4042,N_3220);
and U4743 (N_4743,N_3777,N_3653);
and U4744 (N_4744,N_3076,N_3455);
xnor U4745 (N_4745,N_3845,N_4067);
nand U4746 (N_4746,N_4495,N_3852);
and U4747 (N_4747,N_3313,N_4068);
or U4748 (N_4748,N_3853,N_3187);
or U4749 (N_4749,N_3144,N_3260);
xor U4750 (N_4750,N_3204,N_3934);
xor U4751 (N_4751,N_3195,N_4459);
xor U4752 (N_4752,N_3056,N_3247);
or U4753 (N_4753,N_3898,N_4009);
xnor U4754 (N_4754,N_4391,N_4396);
xnor U4755 (N_4755,N_3461,N_3974);
or U4756 (N_4756,N_3409,N_3843);
nand U4757 (N_4757,N_4101,N_4408);
xor U4758 (N_4758,N_3442,N_3707);
nand U4759 (N_4759,N_3711,N_3483);
xor U4760 (N_4760,N_4416,N_4133);
nand U4761 (N_4761,N_4081,N_3701);
nand U4762 (N_4762,N_4129,N_4249);
nor U4763 (N_4763,N_3015,N_3920);
nor U4764 (N_4764,N_3964,N_3131);
and U4765 (N_4765,N_3061,N_3832);
or U4766 (N_4766,N_4209,N_4264);
nor U4767 (N_4767,N_3752,N_3855);
and U4768 (N_4768,N_4248,N_3706);
and U4769 (N_4769,N_3680,N_4135);
or U4770 (N_4770,N_4347,N_3412);
nand U4771 (N_4771,N_3371,N_3770);
and U4772 (N_4772,N_3052,N_3159);
nor U4773 (N_4773,N_3833,N_3491);
and U4774 (N_4774,N_4368,N_4329);
nand U4775 (N_4775,N_3233,N_3406);
and U4776 (N_4776,N_3596,N_3860);
or U4777 (N_4777,N_4049,N_3098);
or U4778 (N_4778,N_3994,N_3283);
xor U4779 (N_4779,N_3099,N_4123);
and U4780 (N_4780,N_3205,N_3856);
nor U4781 (N_4781,N_3105,N_3501);
xnor U4782 (N_4782,N_4352,N_3280);
and U4783 (N_4783,N_3512,N_3830);
or U4784 (N_4784,N_3466,N_3252);
or U4785 (N_4785,N_4234,N_3390);
and U4786 (N_4786,N_4204,N_4119);
xor U4787 (N_4787,N_3792,N_3049);
and U4788 (N_4788,N_3137,N_4490);
nor U4789 (N_4789,N_4404,N_3958);
and U4790 (N_4790,N_3768,N_4037);
nor U4791 (N_4791,N_3518,N_3265);
nand U4792 (N_4792,N_4157,N_3346);
nor U4793 (N_4793,N_3164,N_3548);
and U4794 (N_4794,N_3077,N_3112);
or U4795 (N_4795,N_4227,N_3003);
nand U4796 (N_4796,N_3277,N_3428);
or U4797 (N_4797,N_3884,N_3256);
nor U4798 (N_4798,N_3771,N_4011);
xor U4799 (N_4799,N_3894,N_3117);
and U4800 (N_4800,N_4188,N_3540);
or U4801 (N_4801,N_3326,N_4341);
nor U4802 (N_4802,N_4440,N_4046);
xor U4803 (N_4803,N_3037,N_3125);
and U4804 (N_4804,N_3709,N_3660);
nand U4805 (N_4805,N_3625,N_3942);
nor U4806 (N_4806,N_3073,N_3392);
and U4807 (N_4807,N_3224,N_3186);
nand U4808 (N_4808,N_3725,N_3962);
xnor U4809 (N_4809,N_3996,N_3369);
or U4810 (N_4810,N_4364,N_4412);
nand U4811 (N_4811,N_4014,N_4211);
xnor U4812 (N_4812,N_3064,N_3193);
xnor U4813 (N_4813,N_4454,N_4203);
nand U4814 (N_4814,N_3987,N_3937);
and U4815 (N_4815,N_4179,N_3951);
xnor U4816 (N_4816,N_3505,N_3936);
nand U4817 (N_4817,N_3511,N_4383);
and U4818 (N_4818,N_3824,N_3763);
xnor U4819 (N_4819,N_3423,N_3139);
xnor U4820 (N_4820,N_3109,N_3888);
nand U4821 (N_4821,N_3901,N_4074);
and U4822 (N_4822,N_3230,N_3330);
nand U4823 (N_4823,N_4008,N_3000);
or U4824 (N_4824,N_4005,N_3785);
xor U4825 (N_4825,N_4044,N_3613);
nand U4826 (N_4826,N_3414,N_3051);
nor U4827 (N_4827,N_3570,N_4019);
nand U4828 (N_4828,N_4279,N_4189);
nor U4829 (N_4829,N_3614,N_3310);
or U4830 (N_4830,N_3899,N_3088);
xnor U4831 (N_4831,N_3817,N_3022);
xor U4832 (N_4832,N_3276,N_3800);
xnor U4833 (N_4833,N_3883,N_4058);
or U4834 (N_4834,N_3445,N_3528);
nand U4835 (N_4835,N_3636,N_4443);
and U4836 (N_4836,N_3897,N_3557);
and U4837 (N_4837,N_3344,N_4356);
and U4838 (N_4838,N_3023,N_3335);
xnor U4839 (N_4839,N_3946,N_3647);
nor U4840 (N_4840,N_4063,N_4221);
xnor U4841 (N_4841,N_3063,N_4090);
nand U4842 (N_4842,N_4164,N_3510);
nand U4843 (N_4843,N_3329,N_3909);
and U4844 (N_4844,N_3810,N_3834);
nor U4845 (N_4845,N_3469,N_3350);
or U4846 (N_4846,N_3146,N_3268);
nand U4847 (N_4847,N_4491,N_3741);
nor U4848 (N_4848,N_4062,N_3586);
nor U4849 (N_4849,N_4228,N_4470);
nand U4850 (N_4850,N_3290,N_3890);
nand U4851 (N_4851,N_3804,N_3069);
nand U4852 (N_4852,N_3041,N_3594);
and U4853 (N_4853,N_3871,N_4020);
and U4854 (N_4854,N_3689,N_4261);
nand U4855 (N_4855,N_4122,N_3047);
and U4856 (N_4856,N_3365,N_3175);
and U4857 (N_4857,N_3774,N_4379);
and U4858 (N_4858,N_4348,N_3039);
xnor U4859 (N_4859,N_3497,N_4312);
and U4860 (N_4860,N_3261,N_3081);
nand U4861 (N_4861,N_4155,N_3686);
xor U4862 (N_4862,N_4399,N_3734);
nand U4863 (N_4863,N_4018,N_3308);
and U4864 (N_4864,N_3132,N_3411);
nor U4865 (N_4865,N_4327,N_4222);
nand U4866 (N_4866,N_3988,N_3282);
and U4867 (N_4867,N_3587,N_3171);
or U4868 (N_4868,N_3864,N_4055);
or U4869 (N_4869,N_3764,N_4095);
nand U4870 (N_4870,N_4025,N_4469);
and U4871 (N_4871,N_3786,N_4200);
or U4872 (N_4872,N_3183,N_3526);
nand U4873 (N_4873,N_3831,N_3381);
nor U4874 (N_4874,N_4468,N_3999);
nand U4875 (N_4875,N_3240,N_3759);
and U4876 (N_4876,N_3385,N_3246);
and U4877 (N_4877,N_3916,N_3337);
nand U4878 (N_4878,N_3926,N_3448);
and U4879 (N_4879,N_3388,N_4316);
nand U4880 (N_4880,N_3387,N_3122);
or U4881 (N_4881,N_3753,N_3384);
and U4882 (N_4882,N_3622,N_3807);
xnor U4883 (N_4883,N_4132,N_4397);
nor U4884 (N_4884,N_4045,N_3944);
nor U4885 (N_4885,N_4177,N_4303);
or U4886 (N_4886,N_3981,N_4376);
and U4887 (N_4887,N_3896,N_3347);
and U4888 (N_4888,N_3654,N_3184);
nand U4889 (N_4889,N_3182,N_4027);
xnor U4890 (N_4890,N_3189,N_3031);
nand U4891 (N_4891,N_3043,N_3516);
or U4892 (N_4892,N_3479,N_4088);
or U4893 (N_4893,N_3531,N_4367);
nand U4894 (N_4894,N_3989,N_4099);
nor U4895 (N_4895,N_4381,N_3262);
nand U4896 (N_4896,N_3742,N_3751);
and U4897 (N_4897,N_3222,N_3656);
and U4898 (N_4898,N_3637,N_3436);
or U4899 (N_4899,N_4237,N_3957);
or U4900 (N_4900,N_3058,N_3115);
or U4901 (N_4901,N_3443,N_3514);
nor U4902 (N_4902,N_3096,N_4393);
and U4903 (N_4903,N_4036,N_4315);
or U4904 (N_4904,N_4409,N_3924);
xnor U4905 (N_4905,N_3395,N_3585);
and U4906 (N_4906,N_3467,N_4201);
or U4907 (N_4907,N_4322,N_3590);
or U4908 (N_4908,N_3292,N_3581);
and U4909 (N_4909,N_3323,N_3279);
nand U4910 (N_4910,N_3236,N_3659);
and U4911 (N_4911,N_3717,N_3788);
nand U4912 (N_4912,N_3874,N_3515);
xnor U4913 (N_4913,N_4392,N_4332);
and U4914 (N_4914,N_3703,N_4395);
xnor U4915 (N_4915,N_3074,N_3102);
or U4916 (N_4916,N_3985,N_4003);
and U4917 (N_4917,N_4206,N_3327);
xor U4918 (N_4918,N_3716,N_3431);
or U4919 (N_4919,N_3914,N_4001);
or U4920 (N_4920,N_3176,N_3667);
xnor U4921 (N_4921,N_3772,N_4484);
nand U4922 (N_4922,N_3967,N_4350);
nor U4923 (N_4923,N_4377,N_4212);
xnor U4924 (N_4924,N_3714,N_3861);
or U4925 (N_4925,N_3975,N_3458);
nor U4926 (N_4926,N_3174,N_3564);
and U4927 (N_4927,N_4400,N_3803);
xnor U4928 (N_4928,N_4252,N_4344);
and U4929 (N_4929,N_3563,N_4442);
or U4930 (N_4930,N_4137,N_4405);
or U4931 (N_4931,N_3438,N_3600);
and U4932 (N_4932,N_3355,N_4338);
or U4933 (N_4933,N_3470,N_4403);
nand U4934 (N_4934,N_4267,N_3542);
nor U4935 (N_4935,N_3082,N_3948);
and U4936 (N_4936,N_3463,N_4402);
nor U4937 (N_4937,N_4107,N_4012);
or U4938 (N_4938,N_4388,N_4407);
nor U4939 (N_4939,N_3722,N_3320);
nand U4940 (N_4940,N_3440,N_4180);
or U4941 (N_4941,N_3363,N_4096);
nor U4942 (N_4942,N_3016,N_4334);
nor U4943 (N_4943,N_3362,N_4224);
xnor U4944 (N_4944,N_3163,N_4198);
nand U4945 (N_4945,N_3950,N_3567);
and U4946 (N_4946,N_3517,N_4485);
nor U4947 (N_4947,N_3812,N_3198);
and U4948 (N_4948,N_4429,N_3295);
nand U4949 (N_4949,N_4130,N_3982);
nor U4950 (N_4950,N_4260,N_3433);
nand U4951 (N_4951,N_3972,N_4072);
nand U4952 (N_4952,N_3161,N_3177);
nand U4953 (N_4953,N_3822,N_3108);
or U4954 (N_4954,N_3249,N_3004);
and U4955 (N_4955,N_4286,N_3778);
nand U4956 (N_4956,N_3997,N_4421);
and U4957 (N_4957,N_3904,N_4121);
or U4958 (N_4958,N_4304,N_4053);
or U4959 (N_4959,N_3848,N_4187);
xnor U4960 (N_4960,N_4172,N_3691);
nor U4961 (N_4961,N_4426,N_3827);
nand U4962 (N_4962,N_3447,N_4217);
or U4963 (N_4963,N_4479,N_3541);
and U4964 (N_4964,N_3203,N_3185);
nor U4965 (N_4965,N_3403,N_4278);
nor U4966 (N_4966,N_3232,N_4365);
or U4967 (N_4967,N_3573,N_4110);
and U4968 (N_4968,N_4465,N_3042);
and U4969 (N_4969,N_3902,N_3969);
or U4970 (N_4970,N_4410,N_3046);
or U4971 (N_4971,N_3207,N_4010);
and U4972 (N_4972,N_3379,N_3057);
and U4973 (N_4973,N_4165,N_3328);
nor U4974 (N_4974,N_4052,N_3012);
nand U4975 (N_4975,N_3545,N_3813);
xnor U4976 (N_4976,N_4477,N_3945);
nor U4977 (N_4977,N_4319,N_3492);
nand U4978 (N_4978,N_3459,N_3973);
xor U4979 (N_4979,N_3825,N_3574);
or U4980 (N_4980,N_3933,N_3679);
or U4981 (N_4981,N_3560,N_3720);
xor U4982 (N_4982,N_3009,N_4464);
and U4983 (N_4983,N_4215,N_3565);
nand U4984 (N_4984,N_3197,N_3375);
xor U4985 (N_4985,N_3138,N_3017);
or U4986 (N_4986,N_3849,N_4126);
and U4987 (N_4987,N_3929,N_3829);
or U4988 (N_4988,N_3629,N_3651);
nor U4989 (N_4989,N_3524,N_3704);
or U4990 (N_4990,N_3710,N_3601);
nor U4991 (N_4991,N_3721,N_3773);
or U4992 (N_4992,N_3954,N_4235);
nor U4993 (N_4993,N_3555,N_3808);
xnor U4994 (N_4994,N_3312,N_3754);
and U4995 (N_4995,N_3444,N_4333);
xnor U4996 (N_4996,N_3739,N_4205);
xor U4997 (N_4997,N_3862,N_3591);
and U4998 (N_4998,N_3858,N_4417);
nor U4999 (N_4999,N_3007,N_3632);
and U5000 (N_5000,N_3726,N_4242);
nand U5001 (N_5001,N_3271,N_3910);
nand U5002 (N_5002,N_4153,N_3239);
nand U5003 (N_5003,N_4104,N_4082);
and U5004 (N_5004,N_3107,N_4467);
nand U5005 (N_5005,N_3696,N_4098);
nand U5006 (N_5006,N_3713,N_3075);
nand U5007 (N_5007,N_4331,N_3289);
or U5008 (N_5008,N_4355,N_3128);
xnor U5009 (N_5009,N_4366,N_3034);
xor U5010 (N_5010,N_4265,N_4112);
xnor U5011 (N_5011,N_3143,N_3353);
and U5012 (N_5012,N_3623,N_4163);
and U5013 (N_5013,N_3306,N_3877);
or U5014 (N_5014,N_3425,N_3229);
or U5015 (N_5015,N_3471,N_4353);
nor U5016 (N_5016,N_4289,N_3038);
nor U5017 (N_5017,N_3421,N_3419);
or U5018 (N_5018,N_3520,N_4273);
and U5019 (N_5019,N_3456,N_3331);
nor U5020 (N_5020,N_4277,N_3441);
or U5021 (N_5021,N_3296,N_4233);
xnor U5022 (N_5022,N_4449,N_3628);
and U5023 (N_5023,N_3357,N_4475);
or U5024 (N_5024,N_3030,N_3737);
xor U5025 (N_5025,N_3866,N_3797);
nand U5026 (N_5026,N_3336,N_4077);
and U5027 (N_5027,N_4185,N_3083);
xnor U5028 (N_5028,N_3869,N_4375);
and U5029 (N_5029,N_3820,N_3917);
and U5030 (N_5030,N_3464,N_4024);
or U5031 (N_5031,N_4384,N_3254);
and U5032 (N_5032,N_4050,N_4351);
and U5033 (N_5033,N_3251,N_3640);
and U5034 (N_5034,N_3150,N_3242);
and U5035 (N_5035,N_3885,N_4427);
nand U5036 (N_5036,N_4196,N_3213);
nand U5037 (N_5037,N_3121,N_4373);
nand U5038 (N_5038,N_3690,N_4151);
xor U5039 (N_5039,N_3578,N_4287);
nand U5040 (N_5040,N_4002,N_3420);
nor U5041 (N_5041,N_3366,N_3267);
nor U5042 (N_5042,N_3490,N_3319);
and U5043 (N_5043,N_3173,N_3842);
and U5044 (N_5044,N_3671,N_3275);
xor U5045 (N_5045,N_4328,N_3097);
and U5046 (N_5046,N_3912,N_3836);
xor U5047 (N_5047,N_4139,N_4240);
and U5048 (N_5048,N_3383,N_3147);
or U5049 (N_5049,N_4195,N_4079);
and U5050 (N_5050,N_3091,N_4487);
nor U5051 (N_5051,N_3072,N_3089);
nor U5052 (N_5052,N_3729,N_3273);
or U5053 (N_5053,N_4496,N_4065);
xnor U5054 (N_5054,N_3397,N_3960);
xor U5055 (N_5055,N_3429,N_4492);
and U5056 (N_5056,N_4306,N_3903);
xnor U5057 (N_5057,N_3539,N_3298);
and U5058 (N_5058,N_3544,N_3854);
and U5059 (N_5059,N_4076,N_3300);
nand U5060 (N_5060,N_3791,N_3806);
nand U5061 (N_5061,N_3180,N_4435);
nand U5062 (N_5062,N_3607,N_4169);
or U5063 (N_5063,N_3062,N_4482);
xnor U5064 (N_5064,N_3399,N_3106);
or U5065 (N_5065,N_3624,N_4238);
and U5066 (N_5066,N_3881,N_3234);
or U5067 (N_5067,N_4268,N_3846);
xor U5068 (N_5068,N_4438,N_3819);
xor U5069 (N_5069,N_3352,N_3535);
nand U5070 (N_5070,N_3675,N_3476);
and U5071 (N_5071,N_3692,N_3170);
or U5072 (N_5072,N_3407,N_4450);
and U5073 (N_5073,N_4091,N_4370);
or U5074 (N_5074,N_3114,N_3922);
and U5075 (N_5075,N_4471,N_3907);
nand U5076 (N_5076,N_4314,N_3712);
nor U5077 (N_5077,N_3664,N_3891);
nor U5078 (N_5078,N_3382,N_3285);
nand U5079 (N_5079,N_3755,N_3032);
nor U5080 (N_5080,N_4061,N_3685);
or U5081 (N_5081,N_4150,N_3274);
nand U5082 (N_5082,N_4193,N_3223);
nor U5083 (N_5083,N_3789,N_3652);
or U5084 (N_5084,N_3761,N_3380);
and U5085 (N_5085,N_3477,N_3816);
nor U5086 (N_5086,N_3878,N_3025);
and U5087 (N_5087,N_4473,N_4463);
nor U5088 (N_5088,N_4033,N_3765);
nand U5089 (N_5089,N_3024,N_3214);
xor U5090 (N_5090,N_3192,N_3536);
and U5091 (N_5091,N_3297,N_3437);
xor U5092 (N_5092,N_4225,N_3886);
and U5093 (N_5093,N_3695,N_3376);
nand U5094 (N_5094,N_3210,N_3460);
nand U5095 (N_5095,N_3801,N_3663);
nand U5096 (N_5096,N_4499,N_3340);
or U5097 (N_5097,N_3984,N_3270);
or U5098 (N_5098,N_4296,N_4030);
nand U5099 (N_5099,N_3348,N_3422);
xnor U5100 (N_5100,N_4372,N_3317);
xnor U5101 (N_5101,N_3080,N_3828);
nand U5102 (N_5102,N_3264,N_3670);
nor U5103 (N_5103,N_3595,N_3169);
nand U5104 (N_5104,N_3961,N_3314);
xor U5105 (N_5105,N_3011,N_3575);
nand U5106 (N_5106,N_3507,N_3859);
xor U5107 (N_5107,N_4498,N_3844);
nor U5108 (N_5108,N_3568,N_4406);
and U5109 (N_5109,N_4305,N_4300);
nand U5110 (N_5110,N_3527,N_3045);
nand U5111 (N_5111,N_4458,N_4102);
nand U5112 (N_5112,N_4161,N_4181);
xnor U5113 (N_5113,N_3293,N_4311);
or U5114 (N_5114,N_3457,N_4160);
xor U5115 (N_5115,N_3927,N_4148);
nor U5116 (N_5116,N_4245,N_3775);
or U5117 (N_5117,N_3496,N_3599);
nor U5118 (N_5118,N_3468,N_3940);
nand U5119 (N_5119,N_3172,N_3892);
and U5120 (N_5120,N_4166,N_4092);
xor U5121 (N_5121,N_4244,N_4359);
nand U5122 (N_5122,N_4420,N_4202);
xor U5123 (N_5123,N_4378,N_4124);
nand U5124 (N_5124,N_3227,N_4309);
nand U5125 (N_5125,N_4170,N_3837);
nand U5126 (N_5126,N_4481,N_4105);
xnor U5127 (N_5127,N_3747,N_3875);
nor U5128 (N_5128,N_3225,N_3760);
or U5129 (N_5129,N_3156,N_3485);
nor U5130 (N_5130,N_4325,N_3678);
nor U5131 (N_5131,N_4308,N_3615);
nor U5132 (N_5132,N_3841,N_3393);
and U5133 (N_5133,N_3129,N_3705);
nor U5134 (N_5134,N_4343,N_4349);
and U5135 (N_5135,N_4178,N_3453);
and U5136 (N_5136,N_3702,N_4097);
xor U5137 (N_5137,N_3134,N_3793);
xor U5138 (N_5138,N_4038,N_3630);
nor U5139 (N_5139,N_3953,N_3811);
xor U5140 (N_5140,N_4208,N_4292);
or U5141 (N_5141,N_3181,N_4385);
xor U5142 (N_5142,N_4103,N_3779);
xnor U5143 (N_5143,N_4280,N_4154);
or U5144 (N_5144,N_3616,N_3373);
nand U5145 (N_5145,N_3482,N_3983);
nand U5146 (N_5146,N_4152,N_3481);
xnor U5147 (N_5147,N_4453,N_4114);
and U5148 (N_5148,N_3814,N_3730);
and U5149 (N_5149,N_3316,N_4031);
or U5150 (N_5150,N_3110,N_4254);
xor U5151 (N_5151,N_3145,N_4006);
and U5152 (N_5152,N_3790,N_4100);
nand U5153 (N_5153,N_3334,N_3727);
nand U5154 (N_5154,N_3167,N_4016);
or U5155 (N_5155,N_3155,N_3212);
xor U5156 (N_5156,N_3191,N_3303);
nand U5157 (N_5157,N_4134,N_3368);
nand U5158 (N_5158,N_3618,N_3165);
xor U5159 (N_5159,N_4253,N_4276);
nor U5160 (N_5160,N_4337,N_3687);
and U5161 (N_5161,N_3499,N_3215);
nor U5162 (N_5162,N_3559,N_4282);
or U5163 (N_5163,N_3488,N_4255);
xnor U5164 (N_5164,N_4318,N_3339);
xnor U5165 (N_5165,N_3519,N_4197);
or U5166 (N_5166,N_3757,N_3876);
nor U5167 (N_5167,N_3724,N_3231);
or U5168 (N_5168,N_4374,N_3676);
and U5169 (N_5169,N_4131,N_3480);
xor U5170 (N_5170,N_3593,N_3451);
and U5171 (N_5171,N_4120,N_3086);
nand U5172 (N_5172,N_3417,N_3010);
xnor U5173 (N_5173,N_3288,N_3815);
xnor U5174 (N_5174,N_3263,N_3284);
or U5175 (N_5175,N_3684,N_4445);
and U5176 (N_5176,N_4271,N_3208);
nand U5177 (N_5177,N_4220,N_4175);
xor U5178 (N_5178,N_3633,N_3238);
and U5179 (N_5179,N_4461,N_3546);
or U5180 (N_5180,N_3345,N_3400);
or U5181 (N_5181,N_4462,N_4230);
nand U5182 (N_5182,N_3092,N_4057);
nand U5183 (N_5183,N_3639,N_3609);
and U5184 (N_5184,N_4069,N_3508);
and U5185 (N_5185,N_3553,N_3682);
xor U5186 (N_5186,N_3141,N_3627);
xor U5187 (N_5187,N_3584,N_4389);
nand U5188 (N_5188,N_3738,N_3847);
xnor U5189 (N_5189,N_3723,N_4317);
xnor U5190 (N_5190,N_3060,N_3589);
and U5191 (N_5191,N_3054,N_3084);
nor U5192 (N_5192,N_3697,N_3424);
and U5193 (N_5193,N_3868,N_4290);
nand U5194 (N_5194,N_3879,N_3657);
nor U5195 (N_5195,N_3065,N_4302);
nand U5196 (N_5196,N_3206,N_4474);
nor U5197 (N_5197,N_3672,N_4313);
xnor U5198 (N_5198,N_4413,N_3026);
or U5199 (N_5199,N_3939,N_3124);
xnor U5200 (N_5200,N_3119,N_3921);
xnor U5201 (N_5201,N_4483,N_3915);
or U5202 (N_5202,N_3561,N_3190);
and U5203 (N_5203,N_4432,N_3111);
nor U5204 (N_5204,N_3840,N_4362);
nor U5205 (N_5205,N_3715,N_3342);
or U5206 (N_5206,N_3959,N_3938);
xor U5207 (N_5207,N_3028,N_3201);
or U5208 (N_5208,N_4085,N_4447);
or U5209 (N_5209,N_4436,N_3522);
xnor U5210 (N_5210,N_3745,N_4246);
nand U5211 (N_5211,N_3305,N_3893);
nor U5212 (N_5212,N_4299,N_4415);
xnor U5213 (N_5213,N_3781,N_4460);
or U5214 (N_5214,N_3918,N_3880);
xnor U5215 (N_5215,N_3537,N_3059);
xnor U5216 (N_5216,N_3642,N_4263);
xnor U5217 (N_5217,N_3626,N_4149);
and U5218 (N_5218,N_3127,N_4418);
nand U5219 (N_5219,N_3818,N_3588);
nor U5220 (N_5220,N_3253,N_4059);
and U5221 (N_5221,N_4431,N_3301);
nand U5222 (N_5222,N_4298,N_3196);
or U5223 (N_5223,N_3503,N_4199);
or U5224 (N_5224,N_3619,N_3554);
xnor U5225 (N_5225,N_3583,N_4258);
and U5226 (N_5226,N_3087,N_3235);
or U5227 (N_5227,N_4424,N_3743);
or U5228 (N_5228,N_3925,N_3226);
nor U5229 (N_5229,N_3020,N_4455);
nor U5230 (N_5230,N_3341,N_3019);
or U5231 (N_5231,N_3620,N_4411);
nand U5232 (N_5232,N_3580,N_4390);
xor U5233 (N_5233,N_4257,N_3243);
or U5234 (N_5234,N_4047,N_3919);
nand U5235 (N_5235,N_3534,N_3221);
or U5236 (N_5236,N_3762,N_3863);
nand U5237 (N_5237,N_4182,N_3732);
nor U5238 (N_5238,N_3120,N_3432);
or U5239 (N_5239,N_3454,N_4108);
and U5240 (N_5240,N_4441,N_3101);
nor U5241 (N_5241,N_3502,N_3217);
or U5242 (N_5242,N_4023,N_3439);
xor U5243 (N_5243,N_3237,N_3533);
nor U5244 (N_5244,N_3610,N_4369);
or U5245 (N_5245,N_3416,N_4007);
nor U5246 (N_5246,N_4342,N_4380);
or U5247 (N_5247,N_3746,N_4480);
nand U5248 (N_5248,N_3332,N_3608);
and U5249 (N_5249,N_4086,N_3426);
or U5250 (N_5250,N_3268,N_3405);
nand U5251 (N_5251,N_4291,N_4023);
and U5252 (N_5252,N_3560,N_3321);
nand U5253 (N_5253,N_4370,N_3932);
xor U5254 (N_5254,N_3397,N_3931);
xor U5255 (N_5255,N_3700,N_3184);
xor U5256 (N_5256,N_3232,N_3177);
xor U5257 (N_5257,N_3888,N_3601);
xnor U5258 (N_5258,N_3454,N_3202);
xor U5259 (N_5259,N_3440,N_3223);
xnor U5260 (N_5260,N_4206,N_3596);
nand U5261 (N_5261,N_3729,N_4450);
and U5262 (N_5262,N_4446,N_3793);
or U5263 (N_5263,N_4401,N_3019);
nand U5264 (N_5264,N_3396,N_3562);
nand U5265 (N_5265,N_3528,N_4359);
and U5266 (N_5266,N_3155,N_3659);
xor U5267 (N_5267,N_3514,N_3229);
nand U5268 (N_5268,N_4185,N_3809);
xnor U5269 (N_5269,N_3947,N_3244);
nor U5270 (N_5270,N_3464,N_4284);
nor U5271 (N_5271,N_4375,N_4382);
and U5272 (N_5272,N_4202,N_3675);
nor U5273 (N_5273,N_4474,N_3239);
and U5274 (N_5274,N_3619,N_3772);
nor U5275 (N_5275,N_3456,N_3487);
xor U5276 (N_5276,N_3072,N_3311);
nand U5277 (N_5277,N_3740,N_3222);
xnor U5278 (N_5278,N_3573,N_3997);
xor U5279 (N_5279,N_3375,N_4470);
nor U5280 (N_5280,N_3223,N_3282);
and U5281 (N_5281,N_3767,N_3209);
or U5282 (N_5282,N_3520,N_3145);
nand U5283 (N_5283,N_3920,N_3971);
nor U5284 (N_5284,N_3907,N_3928);
xor U5285 (N_5285,N_3486,N_3903);
nand U5286 (N_5286,N_3605,N_3229);
xor U5287 (N_5287,N_4388,N_3443);
or U5288 (N_5288,N_3575,N_3471);
or U5289 (N_5289,N_4198,N_3831);
nor U5290 (N_5290,N_3870,N_4344);
and U5291 (N_5291,N_4225,N_3251);
xor U5292 (N_5292,N_3586,N_3453);
and U5293 (N_5293,N_3497,N_3722);
nor U5294 (N_5294,N_4467,N_3906);
or U5295 (N_5295,N_3789,N_3363);
and U5296 (N_5296,N_4251,N_4467);
and U5297 (N_5297,N_3415,N_3515);
nor U5298 (N_5298,N_4240,N_4355);
nor U5299 (N_5299,N_3655,N_4120);
and U5300 (N_5300,N_3051,N_4019);
or U5301 (N_5301,N_3069,N_3237);
xnor U5302 (N_5302,N_4372,N_3447);
nand U5303 (N_5303,N_3728,N_3114);
and U5304 (N_5304,N_3366,N_4035);
nand U5305 (N_5305,N_4282,N_3831);
and U5306 (N_5306,N_4336,N_3903);
xnor U5307 (N_5307,N_4035,N_3505);
xnor U5308 (N_5308,N_3482,N_3786);
nand U5309 (N_5309,N_3410,N_4457);
nor U5310 (N_5310,N_3475,N_3452);
xnor U5311 (N_5311,N_4014,N_4321);
nor U5312 (N_5312,N_4382,N_3585);
and U5313 (N_5313,N_4461,N_4219);
xor U5314 (N_5314,N_3040,N_4465);
xnor U5315 (N_5315,N_3640,N_3153);
and U5316 (N_5316,N_3822,N_4060);
nor U5317 (N_5317,N_4079,N_3525);
and U5318 (N_5318,N_4090,N_3355);
or U5319 (N_5319,N_3296,N_3067);
and U5320 (N_5320,N_3230,N_3258);
xnor U5321 (N_5321,N_4187,N_3447);
or U5322 (N_5322,N_3552,N_3671);
nand U5323 (N_5323,N_3411,N_3253);
nor U5324 (N_5324,N_4320,N_3058);
or U5325 (N_5325,N_4323,N_4384);
xnor U5326 (N_5326,N_3364,N_4486);
xnor U5327 (N_5327,N_3814,N_3749);
xnor U5328 (N_5328,N_3162,N_3012);
xor U5329 (N_5329,N_3506,N_3000);
or U5330 (N_5330,N_3197,N_4421);
nand U5331 (N_5331,N_4007,N_4056);
nand U5332 (N_5332,N_3999,N_4039);
and U5333 (N_5333,N_3569,N_3902);
or U5334 (N_5334,N_3226,N_3737);
xor U5335 (N_5335,N_3863,N_3205);
nand U5336 (N_5336,N_3324,N_3510);
or U5337 (N_5337,N_4126,N_4275);
or U5338 (N_5338,N_3130,N_3650);
nor U5339 (N_5339,N_3897,N_3322);
nor U5340 (N_5340,N_3861,N_3868);
xnor U5341 (N_5341,N_3996,N_3378);
xor U5342 (N_5342,N_3133,N_3830);
or U5343 (N_5343,N_3813,N_3027);
or U5344 (N_5344,N_4319,N_3303);
xor U5345 (N_5345,N_3461,N_3502);
xor U5346 (N_5346,N_3416,N_3893);
and U5347 (N_5347,N_3371,N_4105);
and U5348 (N_5348,N_3108,N_3099);
nor U5349 (N_5349,N_4207,N_3522);
nand U5350 (N_5350,N_4147,N_3194);
and U5351 (N_5351,N_3913,N_3522);
xor U5352 (N_5352,N_4468,N_3626);
or U5353 (N_5353,N_3318,N_3325);
xor U5354 (N_5354,N_3974,N_4448);
xnor U5355 (N_5355,N_3213,N_4462);
nand U5356 (N_5356,N_4310,N_3561);
or U5357 (N_5357,N_4078,N_3702);
or U5358 (N_5358,N_3931,N_4177);
nor U5359 (N_5359,N_4087,N_4446);
nor U5360 (N_5360,N_3940,N_3579);
nor U5361 (N_5361,N_3180,N_3052);
and U5362 (N_5362,N_4492,N_3712);
and U5363 (N_5363,N_3607,N_3966);
nand U5364 (N_5364,N_3200,N_3965);
nor U5365 (N_5365,N_3230,N_3785);
or U5366 (N_5366,N_3405,N_3383);
nor U5367 (N_5367,N_4172,N_3860);
xor U5368 (N_5368,N_3555,N_3383);
xnor U5369 (N_5369,N_4138,N_3162);
xnor U5370 (N_5370,N_3830,N_3771);
and U5371 (N_5371,N_4066,N_3076);
nand U5372 (N_5372,N_4180,N_4206);
xor U5373 (N_5373,N_4277,N_4455);
nor U5374 (N_5374,N_3655,N_3297);
and U5375 (N_5375,N_3568,N_4357);
nor U5376 (N_5376,N_3607,N_3643);
nand U5377 (N_5377,N_4201,N_3206);
and U5378 (N_5378,N_3957,N_3482);
or U5379 (N_5379,N_3738,N_3304);
xnor U5380 (N_5380,N_4363,N_4063);
xnor U5381 (N_5381,N_3524,N_3791);
nor U5382 (N_5382,N_4090,N_3722);
nand U5383 (N_5383,N_4275,N_3507);
nor U5384 (N_5384,N_3196,N_4306);
nand U5385 (N_5385,N_3546,N_3883);
and U5386 (N_5386,N_3155,N_3651);
and U5387 (N_5387,N_4249,N_3363);
or U5388 (N_5388,N_3109,N_3156);
xnor U5389 (N_5389,N_3062,N_3520);
and U5390 (N_5390,N_4197,N_3543);
and U5391 (N_5391,N_4252,N_4213);
nand U5392 (N_5392,N_3774,N_3849);
and U5393 (N_5393,N_3881,N_3230);
xnor U5394 (N_5394,N_3506,N_3821);
or U5395 (N_5395,N_4266,N_3566);
and U5396 (N_5396,N_3966,N_3199);
and U5397 (N_5397,N_3068,N_3234);
or U5398 (N_5398,N_3959,N_4051);
xnor U5399 (N_5399,N_3104,N_3120);
xnor U5400 (N_5400,N_4126,N_4475);
nand U5401 (N_5401,N_3427,N_3437);
nand U5402 (N_5402,N_3908,N_3163);
nor U5403 (N_5403,N_3826,N_4007);
nand U5404 (N_5404,N_4391,N_4431);
nand U5405 (N_5405,N_4313,N_3877);
nand U5406 (N_5406,N_4124,N_4456);
nand U5407 (N_5407,N_3000,N_3059);
xnor U5408 (N_5408,N_3554,N_3963);
nor U5409 (N_5409,N_3590,N_3892);
or U5410 (N_5410,N_4120,N_3361);
nor U5411 (N_5411,N_4145,N_3232);
and U5412 (N_5412,N_3993,N_3165);
xor U5413 (N_5413,N_4203,N_3305);
nand U5414 (N_5414,N_3681,N_3726);
nand U5415 (N_5415,N_3922,N_3892);
xnor U5416 (N_5416,N_3748,N_4225);
xnor U5417 (N_5417,N_3377,N_3329);
or U5418 (N_5418,N_3357,N_3183);
nor U5419 (N_5419,N_4184,N_3071);
or U5420 (N_5420,N_4449,N_3244);
or U5421 (N_5421,N_3155,N_3907);
nand U5422 (N_5422,N_3228,N_4167);
nand U5423 (N_5423,N_4314,N_3622);
or U5424 (N_5424,N_3628,N_3713);
or U5425 (N_5425,N_3195,N_3732);
and U5426 (N_5426,N_3864,N_4118);
nand U5427 (N_5427,N_3281,N_4111);
xor U5428 (N_5428,N_3996,N_3322);
and U5429 (N_5429,N_3049,N_3362);
and U5430 (N_5430,N_4332,N_3856);
nand U5431 (N_5431,N_3875,N_3237);
nor U5432 (N_5432,N_4146,N_4072);
and U5433 (N_5433,N_4125,N_3612);
nand U5434 (N_5434,N_3882,N_3643);
nor U5435 (N_5435,N_4037,N_4415);
and U5436 (N_5436,N_3532,N_3278);
nor U5437 (N_5437,N_3918,N_3235);
or U5438 (N_5438,N_3687,N_4308);
and U5439 (N_5439,N_3204,N_4263);
nor U5440 (N_5440,N_4462,N_4202);
xnor U5441 (N_5441,N_4133,N_4380);
and U5442 (N_5442,N_3200,N_3714);
xor U5443 (N_5443,N_3137,N_3961);
xnor U5444 (N_5444,N_3102,N_3846);
xor U5445 (N_5445,N_3732,N_3823);
and U5446 (N_5446,N_4436,N_4158);
nor U5447 (N_5447,N_3715,N_4333);
nand U5448 (N_5448,N_4162,N_3018);
xor U5449 (N_5449,N_4326,N_4467);
xor U5450 (N_5450,N_3804,N_3029);
xnor U5451 (N_5451,N_3419,N_3329);
or U5452 (N_5452,N_3598,N_3497);
xnor U5453 (N_5453,N_4048,N_3626);
and U5454 (N_5454,N_3442,N_3808);
or U5455 (N_5455,N_4467,N_3790);
and U5456 (N_5456,N_3462,N_3417);
or U5457 (N_5457,N_3728,N_3651);
xor U5458 (N_5458,N_4224,N_3840);
nor U5459 (N_5459,N_4437,N_3348);
and U5460 (N_5460,N_3906,N_4136);
or U5461 (N_5461,N_3567,N_4343);
or U5462 (N_5462,N_3349,N_3076);
or U5463 (N_5463,N_3545,N_4093);
nand U5464 (N_5464,N_4014,N_3177);
or U5465 (N_5465,N_3922,N_3650);
nand U5466 (N_5466,N_4267,N_4042);
nand U5467 (N_5467,N_3733,N_3074);
xnor U5468 (N_5468,N_3458,N_4489);
and U5469 (N_5469,N_3666,N_4026);
or U5470 (N_5470,N_3851,N_3478);
or U5471 (N_5471,N_4219,N_3724);
or U5472 (N_5472,N_3206,N_4226);
and U5473 (N_5473,N_4030,N_3329);
nand U5474 (N_5474,N_3936,N_3432);
xor U5475 (N_5475,N_3332,N_3373);
xor U5476 (N_5476,N_3705,N_3722);
nand U5477 (N_5477,N_4003,N_3885);
and U5478 (N_5478,N_4115,N_3193);
xor U5479 (N_5479,N_3266,N_4042);
or U5480 (N_5480,N_3033,N_3568);
or U5481 (N_5481,N_3514,N_3769);
or U5482 (N_5482,N_3908,N_3799);
and U5483 (N_5483,N_3531,N_3853);
nor U5484 (N_5484,N_3056,N_4134);
nor U5485 (N_5485,N_4437,N_3032);
nand U5486 (N_5486,N_4002,N_3153);
or U5487 (N_5487,N_4173,N_3482);
or U5488 (N_5488,N_3118,N_4111);
xnor U5489 (N_5489,N_4262,N_3064);
nand U5490 (N_5490,N_4434,N_3062);
nand U5491 (N_5491,N_3598,N_3052);
and U5492 (N_5492,N_4208,N_4374);
nor U5493 (N_5493,N_3089,N_3587);
nand U5494 (N_5494,N_3249,N_4053);
nor U5495 (N_5495,N_4471,N_3218);
nor U5496 (N_5496,N_3626,N_3806);
xor U5497 (N_5497,N_4104,N_3023);
and U5498 (N_5498,N_3243,N_4092);
and U5499 (N_5499,N_3319,N_3082);
or U5500 (N_5500,N_3426,N_4351);
nand U5501 (N_5501,N_4257,N_3473);
nor U5502 (N_5502,N_3673,N_3984);
xnor U5503 (N_5503,N_3557,N_4168);
and U5504 (N_5504,N_4325,N_3361);
and U5505 (N_5505,N_3000,N_4353);
or U5506 (N_5506,N_3582,N_3181);
nor U5507 (N_5507,N_4434,N_3917);
or U5508 (N_5508,N_3003,N_3484);
and U5509 (N_5509,N_4106,N_3272);
nand U5510 (N_5510,N_3141,N_3915);
and U5511 (N_5511,N_3394,N_3327);
or U5512 (N_5512,N_4273,N_3845);
nor U5513 (N_5513,N_3394,N_4108);
and U5514 (N_5514,N_3485,N_3587);
and U5515 (N_5515,N_3697,N_3118);
and U5516 (N_5516,N_3673,N_3994);
and U5517 (N_5517,N_4243,N_3769);
and U5518 (N_5518,N_3797,N_3601);
nand U5519 (N_5519,N_3788,N_3124);
xnor U5520 (N_5520,N_4229,N_3304);
xnor U5521 (N_5521,N_3530,N_3731);
nand U5522 (N_5522,N_3837,N_3609);
and U5523 (N_5523,N_4035,N_3356);
or U5524 (N_5524,N_3811,N_4283);
nor U5525 (N_5525,N_4062,N_3095);
nand U5526 (N_5526,N_4243,N_3319);
or U5527 (N_5527,N_3778,N_3868);
xor U5528 (N_5528,N_3689,N_3844);
nand U5529 (N_5529,N_3383,N_4264);
xnor U5530 (N_5530,N_3108,N_3841);
nand U5531 (N_5531,N_3406,N_4023);
nand U5532 (N_5532,N_4449,N_4052);
nor U5533 (N_5533,N_3727,N_3215);
nor U5534 (N_5534,N_3554,N_3914);
or U5535 (N_5535,N_3854,N_4206);
and U5536 (N_5536,N_3830,N_3839);
and U5537 (N_5537,N_4169,N_3819);
xor U5538 (N_5538,N_4288,N_4111);
nand U5539 (N_5539,N_4188,N_3157);
xnor U5540 (N_5540,N_4232,N_3665);
and U5541 (N_5541,N_4263,N_3316);
xnor U5542 (N_5542,N_3058,N_4149);
xnor U5543 (N_5543,N_3235,N_4152);
or U5544 (N_5544,N_3000,N_3587);
xnor U5545 (N_5545,N_3505,N_4220);
nor U5546 (N_5546,N_3534,N_3907);
xor U5547 (N_5547,N_3694,N_3417);
or U5548 (N_5548,N_4474,N_3715);
and U5549 (N_5549,N_3899,N_3447);
or U5550 (N_5550,N_3285,N_3452);
or U5551 (N_5551,N_3564,N_3371);
nor U5552 (N_5552,N_3165,N_4427);
nor U5553 (N_5553,N_4421,N_4077);
or U5554 (N_5554,N_3498,N_3427);
nor U5555 (N_5555,N_4144,N_4314);
or U5556 (N_5556,N_3850,N_3505);
nor U5557 (N_5557,N_3400,N_4359);
nand U5558 (N_5558,N_3654,N_4240);
xnor U5559 (N_5559,N_3449,N_3764);
xnor U5560 (N_5560,N_3140,N_3145);
nor U5561 (N_5561,N_3326,N_4265);
or U5562 (N_5562,N_4345,N_3420);
nand U5563 (N_5563,N_4393,N_3399);
nor U5564 (N_5564,N_4173,N_3419);
xor U5565 (N_5565,N_4075,N_4499);
xnor U5566 (N_5566,N_3237,N_4034);
xor U5567 (N_5567,N_3706,N_4237);
nor U5568 (N_5568,N_3133,N_4004);
or U5569 (N_5569,N_4125,N_4496);
xnor U5570 (N_5570,N_3505,N_4399);
xnor U5571 (N_5571,N_3881,N_4368);
or U5572 (N_5572,N_3516,N_3007);
xor U5573 (N_5573,N_4055,N_4068);
and U5574 (N_5574,N_3049,N_4431);
or U5575 (N_5575,N_4159,N_3307);
nand U5576 (N_5576,N_4119,N_3341);
nor U5577 (N_5577,N_3546,N_3892);
nor U5578 (N_5578,N_3640,N_3941);
or U5579 (N_5579,N_3770,N_3875);
and U5580 (N_5580,N_3058,N_4421);
or U5581 (N_5581,N_3135,N_4010);
and U5582 (N_5582,N_4326,N_4317);
or U5583 (N_5583,N_3123,N_4007);
nor U5584 (N_5584,N_3896,N_3072);
or U5585 (N_5585,N_4038,N_3760);
nor U5586 (N_5586,N_4255,N_3720);
and U5587 (N_5587,N_4184,N_3418);
xnor U5588 (N_5588,N_3762,N_3475);
and U5589 (N_5589,N_3015,N_4402);
xor U5590 (N_5590,N_3316,N_3670);
nand U5591 (N_5591,N_3698,N_3550);
nor U5592 (N_5592,N_3599,N_4283);
and U5593 (N_5593,N_3790,N_3987);
nor U5594 (N_5594,N_4003,N_3467);
nor U5595 (N_5595,N_3648,N_3025);
and U5596 (N_5596,N_4119,N_3153);
nor U5597 (N_5597,N_4497,N_3111);
nor U5598 (N_5598,N_3808,N_3692);
xnor U5599 (N_5599,N_3809,N_3983);
or U5600 (N_5600,N_4435,N_3138);
nor U5601 (N_5601,N_4060,N_3497);
nand U5602 (N_5602,N_3245,N_4111);
or U5603 (N_5603,N_3727,N_3743);
nor U5604 (N_5604,N_3467,N_3531);
xor U5605 (N_5605,N_4344,N_4266);
nand U5606 (N_5606,N_3550,N_3743);
xor U5607 (N_5607,N_3832,N_4170);
nand U5608 (N_5608,N_4289,N_3816);
xor U5609 (N_5609,N_3018,N_3259);
xor U5610 (N_5610,N_3760,N_3218);
or U5611 (N_5611,N_3376,N_3612);
or U5612 (N_5612,N_3357,N_4099);
or U5613 (N_5613,N_3386,N_3405);
nand U5614 (N_5614,N_3073,N_3214);
nor U5615 (N_5615,N_3569,N_4089);
nand U5616 (N_5616,N_4039,N_3965);
or U5617 (N_5617,N_3834,N_4058);
nor U5618 (N_5618,N_4429,N_3967);
nand U5619 (N_5619,N_3783,N_4034);
nand U5620 (N_5620,N_3854,N_3406);
xor U5621 (N_5621,N_3103,N_4212);
xnor U5622 (N_5622,N_3079,N_3149);
nor U5623 (N_5623,N_3055,N_4249);
nor U5624 (N_5624,N_4251,N_3220);
nor U5625 (N_5625,N_3258,N_3943);
xor U5626 (N_5626,N_3998,N_3018);
nand U5627 (N_5627,N_3191,N_3558);
nand U5628 (N_5628,N_3259,N_3869);
xnor U5629 (N_5629,N_3761,N_3580);
nor U5630 (N_5630,N_3562,N_3285);
xor U5631 (N_5631,N_4326,N_3205);
and U5632 (N_5632,N_4297,N_3557);
or U5633 (N_5633,N_3753,N_4446);
and U5634 (N_5634,N_4209,N_3164);
xor U5635 (N_5635,N_4435,N_3662);
nand U5636 (N_5636,N_3964,N_3694);
xor U5637 (N_5637,N_4377,N_3205);
xnor U5638 (N_5638,N_4027,N_3850);
or U5639 (N_5639,N_3193,N_3173);
or U5640 (N_5640,N_3533,N_3879);
nand U5641 (N_5641,N_3172,N_3460);
or U5642 (N_5642,N_3075,N_4270);
nor U5643 (N_5643,N_3606,N_3117);
and U5644 (N_5644,N_3933,N_4037);
nor U5645 (N_5645,N_4113,N_3287);
xnor U5646 (N_5646,N_4002,N_3468);
or U5647 (N_5647,N_4428,N_4449);
xnor U5648 (N_5648,N_3009,N_3102);
xnor U5649 (N_5649,N_4321,N_3603);
nor U5650 (N_5650,N_4375,N_4394);
and U5651 (N_5651,N_3315,N_3310);
or U5652 (N_5652,N_4095,N_4451);
nor U5653 (N_5653,N_3309,N_3490);
nor U5654 (N_5654,N_3035,N_3738);
or U5655 (N_5655,N_3107,N_3473);
nor U5656 (N_5656,N_4318,N_4297);
nand U5657 (N_5657,N_3555,N_4347);
nand U5658 (N_5658,N_4358,N_4118);
and U5659 (N_5659,N_3222,N_3012);
xor U5660 (N_5660,N_4227,N_3159);
or U5661 (N_5661,N_3022,N_4022);
and U5662 (N_5662,N_3474,N_3491);
nand U5663 (N_5663,N_4156,N_3451);
nor U5664 (N_5664,N_4364,N_3440);
nand U5665 (N_5665,N_3393,N_3028);
nand U5666 (N_5666,N_3520,N_3370);
nor U5667 (N_5667,N_4464,N_4311);
xnor U5668 (N_5668,N_4368,N_3711);
and U5669 (N_5669,N_3595,N_3061);
or U5670 (N_5670,N_3539,N_3338);
and U5671 (N_5671,N_4428,N_3089);
nand U5672 (N_5672,N_3483,N_3375);
nand U5673 (N_5673,N_4379,N_4120);
nand U5674 (N_5674,N_4328,N_4158);
or U5675 (N_5675,N_4009,N_3073);
nand U5676 (N_5676,N_3169,N_3980);
nor U5677 (N_5677,N_3544,N_3065);
and U5678 (N_5678,N_4063,N_3921);
or U5679 (N_5679,N_3356,N_3580);
xnor U5680 (N_5680,N_4217,N_4074);
or U5681 (N_5681,N_3879,N_3449);
nor U5682 (N_5682,N_3857,N_3805);
nand U5683 (N_5683,N_3856,N_3151);
xnor U5684 (N_5684,N_3142,N_4199);
nand U5685 (N_5685,N_3124,N_3658);
xor U5686 (N_5686,N_3249,N_3416);
and U5687 (N_5687,N_4233,N_4458);
nand U5688 (N_5688,N_4459,N_3421);
nor U5689 (N_5689,N_3752,N_3264);
xnor U5690 (N_5690,N_3702,N_3366);
and U5691 (N_5691,N_3427,N_3911);
xor U5692 (N_5692,N_3217,N_3645);
nor U5693 (N_5693,N_3729,N_4171);
nor U5694 (N_5694,N_3398,N_4492);
nand U5695 (N_5695,N_4497,N_4484);
or U5696 (N_5696,N_4351,N_3516);
nand U5697 (N_5697,N_3270,N_3566);
or U5698 (N_5698,N_3946,N_3359);
xnor U5699 (N_5699,N_3550,N_3410);
xnor U5700 (N_5700,N_3917,N_3825);
and U5701 (N_5701,N_3015,N_3259);
or U5702 (N_5702,N_3600,N_3163);
xnor U5703 (N_5703,N_3875,N_3259);
xnor U5704 (N_5704,N_4479,N_4274);
xor U5705 (N_5705,N_3479,N_3555);
nand U5706 (N_5706,N_3946,N_3111);
nand U5707 (N_5707,N_3176,N_3716);
xor U5708 (N_5708,N_4061,N_4045);
or U5709 (N_5709,N_4050,N_3184);
xnor U5710 (N_5710,N_3982,N_4065);
or U5711 (N_5711,N_4404,N_3652);
nor U5712 (N_5712,N_3434,N_3888);
xnor U5713 (N_5713,N_3343,N_4005);
xor U5714 (N_5714,N_4140,N_3095);
xnor U5715 (N_5715,N_4043,N_4391);
nor U5716 (N_5716,N_3639,N_3301);
nand U5717 (N_5717,N_3268,N_3050);
nand U5718 (N_5718,N_4128,N_4317);
nand U5719 (N_5719,N_4400,N_3653);
nor U5720 (N_5720,N_3856,N_3509);
nor U5721 (N_5721,N_3631,N_4073);
or U5722 (N_5722,N_4286,N_3420);
xor U5723 (N_5723,N_4002,N_3144);
or U5724 (N_5724,N_3894,N_3957);
or U5725 (N_5725,N_3220,N_3020);
or U5726 (N_5726,N_3810,N_3877);
xor U5727 (N_5727,N_3700,N_3863);
xor U5728 (N_5728,N_3631,N_4244);
nand U5729 (N_5729,N_4081,N_3482);
nand U5730 (N_5730,N_3374,N_3290);
or U5731 (N_5731,N_3620,N_3944);
xor U5732 (N_5732,N_3220,N_4353);
nand U5733 (N_5733,N_3346,N_3158);
nor U5734 (N_5734,N_3881,N_4164);
and U5735 (N_5735,N_4146,N_3749);
or U5736 (N_5736,N_3886,N_3968);
and U5737 (N_5737,N_3059,N_3791);
xor U5738 (N_5738,N_3438,N_3594);
and U5739 (N_5739,N_3151,N_3082);
nor U5740 (N_5740,N_3411,N_3395);
nor U5741 (N_5741,N_3361,N_3893);
nor U5742 (N_5742,N_4325,N_4178);
nor U5743 (N_5743,N_4067,N_4251);
or U5744 (N_5744,N_4010,N_3792);
or U5745 (N_5745,N_3141,N_3704);
nand U5746 (N_5746,N_4069,N_4180);
nor U5747 (N_5747,N_3879,N_4471);
nand U5748 (N_5748,N_3093,N_3584);
nand U5749 (N_5749,N_3588,N_4051);
nor U5750 (N_5750,N_3453,N_4059);
nor U5751 (N_5751,N_3585,N_3381);
or U5752 (N_5752,N_4235,N_3212);
xnor U5753 (N_5753,N_3400,N_3881);
nand U5754 (N_5754,N_3729,N_3713);
nand U5755 (N_5755,N_4422,N_3263);
or U5756 (N_5756,N_3405,N_3313);
and U5757 (N_5757,N_3646,N_3914);
nor U5758 (N_5758,N_3250,N_4150);
or U5759 (N_5759,N_3734,N_3044);
or U5760 (N_5760,N_3721,N_3842);
or U5761 (N_5761,N_3706,N_3423);
xor U5762 (N_5762,N_4008,N_3516);
or U5763 (N_5763,N_4312,N_4005);
nand U5764 (N_5764,N_3907,N_3444);
xnor U5765 (N_5765,N_4040,N_3875);
nand U5766 (N_5766,N_3031,N_3795);
xor U5767 (N_5767,N_3681,N_4416);
xnor U5768 (N_5768,N_3824,N_4211);
nand U5769 (N_5769,N_3636,N_4282);
or U5770 (N_5770,N_3340,N_3464);
nor U5771 (N_5771,N_3420,N_3910);
and U5772 (N_5772,N_3516,N_3817);
xnor U5773 (N_5773,N_3424,N_3566);
nand U5774 (N_5774,N_4280,N_4396);
and U5775 (N_5775,N_4396,N_3281);
nand U5776 (N_5776,N_3194,N_4035);
nand U5777 (N_5777,N_3244,N_3431);
xor U5778 (N_5778,N_3693,N_3698);
and U5779 (N_5779,N_4229,N_4191);
or U5780 (N_5780,N_4255,N_4187);
nand U5781 (N_5781,N_4218,N_3445);
and U5782 (N_5782,N_3534,N_3543);
or U5783 (N_5783,N_3005,N_4078);
nand U5784 (N_5784,N_4265,N_4171);
or U5785 (N_5785,N_3718,N_3274);
nor U5786 (N_5786,N_3318,N_3089);
and U5787 (N_5787,N_3169,N_3231);
and U5788 (N_5788,N_3797,N_3189);
xnor U5789 (N_5789,N_4132,N_3022);
nor U5790 (N_5790,N_3996,N_3274);
xor U5791 (N_5791,N_3420,N_3237);
nand U5792 (N_5792,N_3694,N_3023);
nand U5793 (N_5793,N_3304,N_3568);
and U5794 (N_5794,N_3621,N_3219);
and U5795 (N_5795,N_3609,N_3465);
or U5796 (N_5796,N_4411,N_3500);
nor U5797 (N_5797,N_3241,N_3088);
xor U5798 (N_5798,N_3922,N_3948);
and U5799 (N_5799,N_3709,N_3963);
or U5800 (N_5800,N_3436,N_4429);
or U5801 (N_5801,N_4302,N_3146);
nor U5802 (N_5802,N_3938,N_3848);
nand U5803 (N_5803,N_3135,N_4174);
nor U5804 (N_5804,N_3463,N_4297);
nor U5805 (N_5805,N_3458,N_3313);
and U5806 (N_5806,N_3006,N_4256);
xnor U5807 (N_5807,N_3231,N_3129);
and U5808 (N_5808,N_3324,N_3157);
nor U5809 (N_5809,N_3562,N_4333);
xnor U5810 (N_5810,N_3996,N_3205);
nand U5811 (N_5811,N_3275,N_4307);
or U5812 (N_5812,N_4177,N_3018);
nand U5813 (N_5813,N_3428,N_3641);
nand U5814 (N_5814,N_4334,N_3592);
or U5815 (N_5815,N_3217,N_3508);
nor U5816 (N_5816,N_3394,N_3406);
and U5817 (N_5817,N_3217,N_4018);
nand U5818 (N_5818,N_3291,N_3568);
or U5819 (N_5819,N_3346,N_4031);
nand U5820 (N_5820,N_4264,N_4412);
xor U5821 (N_5821,N_4182,N_3315);
nand U5822 (N_5822,N_3431,N_3124);
nand U5823 (N_5823,N_4159,N_3637);
nor U5824 (N_5824,N_4114,N_4399);
and U5825 (N_5825,N_3090,N_3696);
and U5826 (N_5826,N_4030,N_4464);
and U5827 (N_5827,N_3331,N_3854);
or U5828 (N_5828,N_4484,N_3012);
and U5829 (N_5829,N_3531,N_4360);
and U5830 (N_5830,N_4053,N_4149);
nand U5831 (N_5831,N_3291,N_3631);
or U5832 (N_5832,N_3343,N_4215);
xor U5833 (N_5833,N_3222,N_3923);
or U5834 (N_5834,N_4450,N_4131);
and U5835 (N_5835,N_3674,N_3704);
xor U5836 (N_5836,N_4035,N_4350);
or U5837 (N_5837,N_3109,N_3487);
nand U5838 (N_5838,N_3772,N_3136);
and U5839 (N_5839,N_4405,N_3081);
nand U5840 (N_5840,N_4436,N_4445);
nand U5841 (N_5841,N_4115,N_3457);
or U5842 (N_5842,N_3529,N_3014);
nand U5843 (N_5843,N_4142,N_3814);
or U5844 (N_5844,N_3035,N_3201);
nor U5845 (N_5845,N_3021,N_3860);
nand U5846 (N_5846,N_3073,N_3885);
nor U5847 (N_5847,N_3772,N_4183);
xor U5848 (N_5848,N_3351,N_3669);
and U5849 (N_5849,N_4499,N_3993);
and U5850 (N_5850,N_4361,N_3377);
xnor U5851 (N_5851,N_3209,N_3640);
xnor U5852 (N_5852,N_4399,N_3252);
nand U5853 (N_5853,N_4351,N_4222);
nand U5854 (N_5854,N_3203,N_3515);
and U5855 (N_5855,N_3651,N_3273);
or U5856 (N_5856,N_3927,N_3949);
nand U5857 (N_5857,N_3136,N_3468);
or U5858 (N_5858,N_4122,N_3364);
and U5859 (N_5859,N_3809,N_3389);
nand U5860 (N_5860,N_3183,N_3982);
nor U5861 (N_5861,N_4073,N_4468);
nand U5862 (N_5862,N_3949,N_3965);
xnor U5863 (N_5863,N_4104,N_3942);
nand U5864 (N_5864,N_4231,N_4296);
nor U5865 (N_5865,N_3566,N_3484);
nand U5866 (N_5866,N_4267,N_3522);
and U5867 (N_5867,N_3121,N_4178);
and U5868 (N_5868,N_4439,N_3040);
and U5869 (N_5869,N_3002,N_3835);
or U5870 (N_5870,N_4398,N_3213);
and U5871 (N_5871,N_3854,N_3950);
xor U5872 (N_5872,N_3357,N_3259);
and U5873 (N_5873,N_3659,N_3486);
or U5874 (N_5874,N_3291,N_4371);
xor U5875 (N_5875,N_4267,N_3818);
xor U5876 (N_5876,N_3494,N_3608);
xor U5877 (N_5877,N_4486,N_4075);
xnor U5878 (N_5878,N_3379,N_3668);
nand U5879 (N_5879,N_3823,N_4195);
or U5880 (N_5880,N_3777,N_3285);
xor U5881 (N_5881,N_3459,N_4197);
nand U5882 (N_5882,N_3348,N_4036);
nor U5883 (N_5883,N_3106,N_3439);
or U5884 (N_5884,N_3298,N_3500);
nand U5885 (N_5885,N_3637,N_3756);
xnor U5886 (N_5886,N_3815,N_4337);
or U5887 (N_5887,N_3948,N_3517);
or U5888 (N_5888,N_4386,N_3591);
or U5889 (N_5889,N_3708,N_3181);
or U5890 (N_5890,N_3678,N_3519);
xor U5891 (N_5891,N_4127,N_4399);
and U5892 (N_5892,N_4397,N_3605);
and U5893 (N_5893,N_3187,N_3532);
and U5894 (N_5894,N_3573,N_4104);
nor U5895 (N_5895,N_4290,N_3536);
or U5896 (N_5896,N_4300,N_3408);
xor U5897 (N_5897,N_3185,N_4320);
or U5898 (N_5898,N_3329,N_3098);
nor U5899 (N_5899,N_3856,N_3162);
nand U5900 (N_5900,N_3180,N_3210);
nor U5901 (N_5901,N_3080,N_3025);
and U5902 (N_5902,N_3620,N_4464);
nand U5903 (N_5903,N_4247,N_4029);
nand U5904 (N_5904,N_3210,N_3762);
and U5905 (N_5905,N_3022,N_3416);
or U5906 (N_5906,N_3453,N_3918);
nor U5907 (N_5907,N_3176,N_4301);
or U5908 (N_5908,N_3433,N_3077);
and U5909 (N_5909,N_3313,N_3026);
xor U5910 (N_5910,N_4274,N_3729);
and U5911 (N_5911,N_4354,N_3235);
and U5912 (N_5912,N_3146,N_3030);
nand U5913 (N_5913,N_4244,N_3802);
or U5914 (N_5914,N_3332,N_3912);
or U5915 (N_5915,N_3714,N_3882);
or U5916 (N_5916,N_3295,N_4008);
nor U5917 (N_5917,N_3169,N_3518);
xor U5918 (N_5918,N_4215,N_3186);
and U5919 (N_5919,N_3846,N_3948);
nand U5920 (N_5920,N_3432,N_4291);
or U5921 (N_5921,N_4257,N_3527);
nand U5922 (N_5922,N_3080,N_3672);
or U5923 (N_5923,N_3661,N_3910);
nor U5924 (N_5924,N_4173,N_3739);
nand U5925 (N_5925,N_3766,N_4044);
nand U5926 (N_5926,N_3090,N_3101);
and U5927 (N_5927,N_3784,N_4488);
xor U5928 (N_5928,N_3685,N_3810);
xor U5929 (N_5929,N_4256,N_3953);
or U5930 (N_5930,N_3066,N_3378);
xor U5931 (N_5931,N_4155,N_3182);
xor U5932 (N_5932,N_3084,N_4380);
xnor U5933 (N_5933,N_3452,N_4324);
or U5934 (N_5934,N_3002,N_3784);
and U5935 (N_5935,N_3935,N_3837);
xor U5936 (N_5936,N_4267,N_4117);
xnor U5937 (N_5937,N_3904,N_4004);
and U5938 (N_5938,N_3625,N_3916);
nand U5939 (N_5939,N_3267,N_3790);
and U5940 (N_5940,N_4459,N_4205);
nand U5941 (N_5941,N_3271,N_3334);
and U5942 (N_5942,N_3927,N_3473);
xnor U5943 (N_5943,N_3044,N_3780);
xor U5944 (N_5944,N_3754,N_3490);
and U5945 (N_5945,N_4139,N_3439);
nand U5946 (N_5946,N_4053,N_3251);
and U5947 (N_5947,N_3406,N_3895);
xor U5948 (N_5948,N_4148,N_4005);
nor U5949 (N_5949,N_3830,N_3858);
and U5950 (N_5950,N_3617,N_4146);
nand U5951 (N_5951,N_3356,N_3299);
nor U5952 (N_5952,N_4275,N_3546);
and U5953 (N_5953,N_3212,N_4162);
nand U5954 (N_5954,N_4053,N_3333);
nand U5955 (N_5955,N_4354,N_4226);
or U5956 (N_5956,N_3936,N_3045);
or U5957 (N_5957,N_4390,N_4466);
nand U5958 (N_5958,N_3919,N_3684);
xnor U5959 (N_5959,N_4490,N_3011);
and U5960 (N_5960,N_3501,N_3091);
nand U5961 (N_5961,N_3556,N_3758);
nor U5962 (N_5962,N_3779,N_4140);
and U5963 (N_5963,N_4259,N_3356);
nand U5964 (N_5964,N_3557,N_4193);
and U5965 (N_5965,N_3205,N_4477);
nand U5966 (N_5966,N_3334,N_3703);
nor U5967 (N_5967,N_3676,N_4220);
nor U5968 (N_5968,N_3709,N_4361);
xnor U5969 (N_5969,N_3577,N_3309);
or U5970 (N_5970,N_3705,N_3868);
or U5971 (N_5971,N_3942,N_4119);
and U5972 (N_5972,N_4159,N_3857);
nor U5973 (N_5973,N_4227,N_3858);
nand U5974 (N_5974,N_3037,N_4171);
nand U5975 (N_5975,N_4016,N_4378);
nand U5976 (N_5976,N_3640,N_3413);
xor U5977 (N_5977,N_3226,N_3833);
xnor U5978 (N_5978,N_3774,N_3234);
nor U5979 (N_5979,N_3464,N_4186);
nor U5980 (N_5980,N_4235,N_3290);
and U5981 (N_5981,N_4253,N_3962);
or U5982 (N_5982,N_4184,N_3356);
and U5983 (N_5983,N_4017,N_3773);
xnor U5984 (N_5984,N_3822,N_3033);
and U5985 (N_5985,N_3737,N_3669);
nand U5986 (N_5986,N_3115,N_3076);
xnor U5987 (N_5987,N_4389,N_3209);
nor U5988 (N_5988,N_3336,N_4245);
and U5989 (N_5989,N_3088,N_3075);
nand U5990 (N_5990,N_3159,N_4235);
nand U5991 (N_5991,N_4256,N_3289);
or U5992 (N_5992,N_3828,N_4306);
xor U5993 (N_5993,N_3698,N_4447);
nand U5994 (N_5994,N_4480,N_3072);
and U5995 (N_5995,N_3329,N_3921);
and U5996 (N_5996,N_3138,N_4183);
nand U5997 (N_5997,N_3175,N_3694);
nand U5998 (N_5998,N_3074,N_3322);
and U5999 (N_5999,N_3709,N_4048);
nand U6000 (N_6000,N_5256,N_5686);
xor U6001 (N_6001,N_4599,N_5721);
or U6002 (N_6002,N_5581,N_4649);
and U6003 (N_6003,N_5364,N_4638);
or U6004 (N_6004,N_5536,N_5767);
nand U6005 (N_6005,N_4914,N_4570);
xnor U6006 (N_6006,N_5317,N_5279);
nor U6007 (N_6007,N_4841,N_4537);
or U6008 (N_6008,N_4620,N_5793);
nand U6009 (N_6009,N_4913,N_4601);
and U6010 (N_6010,N_5494,N_5040);
and U6011 (N_6011,N_5782,N_5458);
and U6012 (N_6012,N_4732,N_5174);
xor U6013 (N_6013,N_4854,N_5672);
xnor U6014 (N_6014,N_4922,N_5950);
nor U6015 (N_6015,N_5539,N_4549);
and U6016 (N_6016,N_4604,N_5342);
nor U6017 (N_6017,N_4832,N_4778);
and U6018 (N_6018,N_5841,N_5169);
nor U6019 (N_6019,N_5923,N_5197);
nor U6020 (N_6020,N_5816,N_4659);
nor U6021 (N_6021,N_4676,N_4925);
and U6022 (N_6022,N_5319,N_4643);
or U6023 (N_6023,N_5257,N_5131);
nor U6024 (N_6024,N_4629,N_4806);
nor U6025 (N_6025,N_5114,N_4651);
or U6026 (N_6026,N_5071,N_5368);
and U6027 (N_6027,N_5199,N_5359);
and U6028 (N_6028,N_5920,N_5451);
nor U6029 (N_6029,N_5490,N_4703);
nor U6030 (N_6030,N_5892,N_5527);
or U6031 (N_6031,N_5992,N_4945);
nor U6032 (N_6032,N_5238,N_5370);
nand U6033 (N_6033,N_4605,N_5618);
and U6034 (N_6034,N_5975,N_5388);
xnor U6035 (N_6035,N_5705,N_4710);
or U6036 (N_6036,N_5086,N_5204);
xnor U6037 (N_6037,N_4892,N_5945);
or U6038 (N_6038,N_4987,N_5965);
nand U6039 (N_6039,N_5399,N_5676);
nor U6040 (N_6040,N_5855,N_5020);
nand U6041 (N_6041,N_5988,N_5980);
xor U6042 (N_6042,N_5015,N_5674);
xnor U6043 (N_6043,N_4609,N_4654);
nand U6044 (N_6044,N_5515,N_4756);
or U6045 (N_6045,N_4689,N_5185);
or U6046 (N_6046,N_5749,N_5208);
nor U6047 (N_6047,N_5847,N_4993);
xnor U6048 (N_6048,N_5813,N_5003);
or U6049 (N_6049,N_5396,N_4837);
nand U6050 (N_6050,N_5982,N_5122);
nand U6051 (N_6051,N_4575,N_5156);
nor U6052 (N_6052,N_4765,N_5507);
nor U6053 (N_6053,N_4800,N_5424);
or U6054 (N_6054,N_5292,N_5972);
xor U6055 (N_6055,N_4717,N_5990);
or U6056 (N_6056,N_5378,N_4555);
nor U6057 (N_6057,N_4773,N_5382);
nor U6058 (N_6058,N_5710,N_5177);
xor U6059 (N_6059,N_4641,N_5836);
xnor U6060 (N_6060,N_5662,N_5597);
or U6061 (N_6061,N_4571,N_4504);
and U6062 (N_6062,N_5949,N_4634);
and U6063 (N_6063,N_5121,N_5734);
and U6064 (N_6064,N_4940,N_4650);
nor U6065 (N_6065,N_5299,N_5790);
nor U6066 (N_6066,N_4866,N_5008);
or U6067 (N_6067,N_4997,N_5777);
and U6068 (N_6068,N_5338,N_5851);
nand U6069 (N_6069,N_5496,N_4934);
xor U6070 (N_6070,N_4972,N_5126);
and U6071 (N_6071,N_5442,N_4506);
or U6072 (N_6072,N_4804,N_5628);
and U6073 (N_6073,N_4895,N_5498);
xnor U6074 (N_6074,N_4858,N_5145);
xor U6075 (N_6075,N_5420,N_5843);
nor U6076 (N_6076,N_5233,N_5077);
nor U6077 (N_6077,N_4781,N_4603);
xor U6078 (N_6078,N_5158,N_4818);
xor U6079 (N_6079,N_5989,N_5026);
nand U6080 (N_6080,N_4885,N_5373);
nor U6081 (N_6081,N_5955,N_5390);
and U6082 (N_6082,N_5694,N_5172);
nand U6083 (N_6083,N_4876,N_5886);
nand U6084 (N_6084,N_5437,N_4730);
and U6085 (N_6085,N_5859,N_4708);
or U6086 (N_6086,N_5544,N_4891);
and U6087 (N_6087,N_4927,N_5203);
nand U6088 (N_6088,N_5309,N_5042);
nor U6089 (N_6089,N_5592,N_4842);
and U6090 (N_6090,N_5247,N_5932);
nand U6091 (N_6091,N_4662,N_5577);
and U6092 (N_6092,N_4748,N_5022);
nand U6093 (N_6093,N_4663,N_5068);
and U6094 (N_6094,N_5792,N_5695);
xor U6095 (N_6095,N_4742,N_4655);
nor U6096 (N_6096,N_4721,N_5845);
or U6097 (N_6097,N_5271,N_5134);
or U6098 (N_6098,N_5983,N_5113);
nand U6099 (N_6099,N_4574,N_4500);
nand U6100 (N_6100,N_5787,N_5838);
or U6101 (N_6101,N_5820,N_5439);
or U6102 (N_6102,N_5291,N_4592);
and U6103 (N_6103,N_4896,N_5282);
nand U6104 (N_6104,N_5229,N_4980);
and U6105 (N_6105,N_5385,N_5994);
xor U6106 (N_6106,N_4660,N_4967);
xor U6107 (N_6107,N_5211,N_5427);
xnor U6108 (N_6108,N_5685,N_5996);
nand U6109 (N_6109,N_5173,N_4633);
or U6110 (N_6110,N_5181,N_4652);
and U6111 (N_6111,N_5105,N_5154);
nand U6112 (N_6112,N_4690,N_5899);
and U6113 (N_6113,N_5314,N_5028);
and U6114 (N_6114,N_5800,N_5088);
or U6115 (N_6115,N_5822,N_5944);
or U6116 (N_6116,N_4734,N_5726);
and U6117 (N_6117,N_5973,N_5339);
nand U6118 (N_6118,N_5664,N_5423);
and U6119 (N_6119,N_5715,N_5522);
nor U6120 (N_6120,N_5725,N_5625);
nand U6121 (N_6121,N_4758,N_4658);
nor U6122 (N_6122,N_5999,N_5153);
xnor U6123 (N_6123,N_5948,N_5605);
and U6124 (N_6124,N_4779,N_5658);
xnor U6125 (N_6125,N_4761,N_4939);
and U6126 (N_6126,N_5106,N_5019);
and U6127 (N_6127,N_5261,N_5642);
nor U6128 (N_6128,N_4751,N_4507);
nor U6129 (N_6129,N_4816,N_5495);
or U6130 (N_6130,N_5554,N_5450);
and U6131 (N_6131,N_5645,N_4801);
nand U6132 (N_6132,N_4681,N_5748);
or U6133 (N_6133,N_5445,N_5723);
and U6134 (N_6134,N_4912,N_4821);
and U6135 (N_6135,N_4520,N_4589);
nand U6136 (N_6136,N_5010,N_4695);
and U6137 (N_6137,N_5497,N_5500);
or U6138 (N_6138,N_5818,N_5283);
or U6139 (N_6139,N_4870,N_5732);
and U6140 (N_6140,N_4796,N_4745);
and U6141 (N_6141,N_4607,N_5051);
nand U6142 (N_6142,N_5140,N_4606);
and U6143 (N_6143,N_4984,N_4992);
xnor U6144 (N_6144,N_5575,N_5417);
and U6145 (N_6145,N_4554,N_5812);
xnor U6146 (N_6146,N_5516,N_4965);
nand U6147 (N_6147,N_5614,N_4840);
nand U6148 (N_6148,N_5655,N_4580);
xor U6149 (N_6149,N_5700,N_5549);
nor U6150 (N_6150,N_5082,N_5954);
xor U6151 (N_6151,N_5183,N_4808);
nand U6152 (N_6152,N_5833,N_5906);
and U6153 (N_6153,N_5743,N_5601);
nor U6154 (N_6154,N_5995,N_5201);
nand U6155 (N_6155,N_5320,N_5104);
and U6156 (N_6156,N_5819,N_5719);
and U6157 (N_6157,N_5831,N_5880);
xor U6158 (N_6158,N_4883,N_5135);
nand U6159 (N_6159,N_4834,N_4583);
and U6160 (N_6160,N_4872,N_5834);
or U6161 (N_6161,N_5136,N_5002);
nand U6162 (N_6162,N_4701,N_4971);
or U6163 (N_6163,N_5746,N_5991);
or U6164 (N_6164,N_4904,N_5771);
xnor U6165 (N_6165,N_5683,N_5877);
nand U6166 (N_6166,N_5421,N_5621);
xnor U6167 (N_6167,N_4964,N_4882);
xnor U6168 (N_6168,N_4849,N_4615);
xnor U6169 (N_6169,N_5084,N_4587);
and U6170 (N_6170,N_5934,N_4924);
xnor U6171 (N_6171,N_5893,N_5479);
nand U6172 (N_6172,N_5325,N_5039);
and U6173 (N_6173,N_5017,N_4713);
and U6174 (N_6174,N_5250,N_4795);
nor U6175 (N_6175,N_5332,N_4665);
or U6176 (N_6176,N_4624,N_5119);
xnor U6177 (N_6177,N_4829,N_5894);
xor U6178 (N_6178,N_5330,N_5901);
or U6179 (N_6179,N_4978,N_5759);
and U6180 (N_6180,N_4722,N_5200);
nor U6181 (N_6181,N_5046,N_5150);
nand U6182 (N_6182,N_5503,N_5272);
nor U6183 (N_6183,N_4811,N_5228);
or U6184 (N_6184,N_5524,N_4657);
xnor U6185 (N_6185,N_5138,N_5363);
nand U6186 (N_6186,N_5722,N_5352);
or U6187 (N_6187,N_4564,N_4548);
or U6188 (N_6188,N_4672,N_5799);
xnor U6189 (N_6189,N_4738,N_4519);
or U6190 (N_6190,N_4505,N_4878);
or U6191 (N_6191,N_5116,N_5778);
and U6192 (N_6192,N_5684,N_5059);
or U6193 (N_6193,N_5141,N_5227);
or U6194 (N_6194,N_5548,N_5085);
and U6195 (N_6195,N_5783,N_5047);
and U6196 (N_6196,N_4792,N_5281);
nor U6197 (N_6197,N_4707,N_5638);
or U6198 (N_6198,N_5191,N_5579);
and U6199 (N_6199,N_4935,N_5323);
or U6200 (N_6200,N_5187,N_5570);
and U6201 (N_6201,N_5933,N_5340);
or U6202 (N_6202,N_5938,N_5049);
and U6203 (N_6203,N_4825,N_5069);
or U6204 (N_6204,N_4611,N_4595);
or U6205 (N_6205,N_4524,N_5418);
nor U6206 (N_6206,N_4529,N_4823);
nand U6207 (N_6207,N_4897,N_4983);
and U6208 (N_6208,N_4942,N_5697);
nor U6209 (N_6209,N_5569,N_5898);
or U6210 (N_6210,N_5699,N_4747);
nand U6211 (N_6211,N_4953,N_5306);
and U6212 (N_6212,N_4588,N_4508);
and U6213 (N_6213,N_4715,N_4780);
nor U6214 (N_6214,N_5875,N_5770);
or U6215 (N_6215,N_4740,N_5907);
nand U6216 (N_6216,N_5160,N_5962);
nor U6217 (N_6217,N_5830,N_5184);
or U6218 (N_6218,N_5728,N_5571);
and U6219 (N_6219,N_4797,N_5667);
nor U6220 (N_6220,N_5629,N_5037);
nor U6221 (N_6221,N_5824,N_5426);
nor U6222 (N_6222,N_4950,N_5061);
or U6223 (N_6223,N_5429,N_5795);
xor U6224 (N_6224,N_5916,N_4704);
and U6225 (N_6225,N_5466,N_5487);
or U6226 (N_6226,N_5506,N_5966);
and U6227 (N_6227,N_4810,N_5375);
or U6228 (N_6228,N_5033,N_5112);
or U6229 (N_6229,N_5448,N_5758);
nand U6230 (N_6230,N_4510,N_5963);
nand U6231 (N_6231,N_4838,N_5313);
and U6232 (N_6232,N_4943,N_5129);
nor U6233 (N_6233,N_4687,N_5666);
nor U6234 (N_6234,N_4711,N_4726);
nand U6235 (N_6235,N_5155,N_4819);
xor U6236 (N_6236,N_5198,N_4626);
xor U6237 (N_6237,N_5351,N_5517);
nand U6238 (N_6238,N_5852,N_4642);
and U6239 (N_6239,N_5882,N_5808);
nor U6240 (N_6240,N_5157,N_5231);
and U6241 (N_6241,N_4608,N_5453);
nand U6242 (N_6242,N_5095,N_4512);
nand U6243 (N_6243,N_5904,N_4824);
and U6244 (N_6244,N_5166,N_5985);
or U6245 (N_6245,N_4528,N_4898);
or U6246 (N_6246,N_5724,N_4817);
or U6247 (N_6247,N_4929,N_4814);
nand U6248 (N_6248,N_5930,N_5005);
and U6249 (N_6249,N_5263,N_4621);
xor U6250 (N_6250,N_5000,N_5066);
and U6251 (N_6251,N_5840,N_5925);
nand U6252 (N_6252,N_5585,N_5692);
and U6253 (N_6253,N_5300,N_4514);
nor U6254 (N_6254,N_4909,N_4550);
and U6255 (N_6255,N_5482,N_5682);
nand U6256 (N_6256,N_5297,N_5997);
nor U6257 (N_6257,N_5584,N_5961);
xor U6258 (N_6258,N_5656,N_5290);
and U6259 (N_6259,N_5897,N_5626);
and U6260 (N_6260,N_5414,N_5805);
nor U6261 (N_6261,N_5083,N_5730);
and U6262 (N_6262,N_5394,N_4557);
nor U6263 (N_6263,N_5092,N_5050);
and U6264 (N_6264,N_4783,N_5600);
nand U6265 (N_6265,N_5243,N_5214);
xor U6266 (N_6266,N_5305,N_5698);
or U6267 (N_6267,N_5251,N_4716);
or U6268 (N_6268,N_5333,N_5718);
or U6269 (N_6269,N_4737,N_5193);
or U6270 (N_6270,N_4576,N_4622);
xnor U6271 (N_6271,N_5736,N_5196);
xnor U6272 (N_6272,N_4600,N_5491);
or U6273 (N_6273,N_5555,N_5087);
xnor U6274 (N_6274,N_5668,N_5964);
nand U6275 (N_6275,N_4631,N_5739);
xor U6276 (N_6276,N_5761,N_5354);
and U6277 (N_6277,N_5557,N_5124);
xnor U6278 (N_6278,N_4692,N_4637);
xor U6279 (N_6279,N_5031,N_4820);
or U6280 (N_6280,N_4614,N_4805);
nor U6281 (N_6281,N_5435,N_5784);
nor U6282 (N_6282,N_5849,N_5977);
nor U6283 (N_6283,N_4705,N_5304);
or U6284 (N_6284,N_4616,N_5910);
nand U6285 (N_6285,N_4563,N_4789);
and U6286 (N_6286,N_4976,N_4851);
xor U6287 (N_6287,N_5559,N_5170);
or U6288 (N_6288,N_4661,N_5096);
xor U6289 (N_6289,N_5641,N_4847);
nand U6290 (N_6290,N_5232,N_4749);
nand U6291 (N_6291,N_5774,N_4848);
nand U6292 (N_6292,N_5034,N_5355);
nand U6293 (N_6293,N_5216,N_5615);
nor U6294 (N_6294,N_5460,N_5318);
nand U6295 (N_6295,N_5461,N_5463);
and U6296 (N_6296,N_5775,N_5312);
nand U6297 (N_6297,N_5884,N_4936);
or U6298 (N_6298,N_5891,N_5689);
nand U6299 (N_6299,N_5081,N_4932);
nand U6300 (N_6300,N_5434,N_4731);
nor U6301 (N_6301,N_5727,N_4602);
or U6302 (N_6302,N_5946,N_5098);
xnor U6303 (N_6303,N_5956,N_4969);
and U6304 (N_6304,N_4910,N_5372);
nor U6305 (N_6305,N_5623,N_5217);
xnor U6306 (N_6306,N_5711,N_4900);
nor U6307 (N_6307,N_4799,N_4996);
nand U6308 (N_6308,N_5935,N_4668);
nand U6309 (N_6309,N_5480,N_4887);
nand U6310 (N_6310,N_5254,N_4618);
nand U6311 (N_6311,N_5888,N_5287);
and U6312 (N_6312,N_5873,N_5235);
nand U6313 (N_6313,N_5869,N_4839);
nand U6314 (N_6314,N_5979,N_5179);
xnor U6315 (N_6315,N_4802,N_5709);
or U6316 (N_6316,N_5298,N_4544);
nor U6317 (N_6317,N_4613,N_5163);
nand U6318 (N_6318,N_5713,N_4509);
and U6319 (N_6319,N_5814,N_5970);
xnor U6320 (N_6320,N_5974,N_5918);
or U6321 (N_6321,N_4886,N_5653);
nor U6322 (N_6322,N_5789,N_4877);
nor U6323 (N_6323,N_5073,N_4868);
xor U6324 (N_6324,N_5596,N_4764);
and U6325 (N_6325,N_5143,N_5681);
nand U6326 (N_6326,N_5921,N_5374);
nand U6327 (N_6327,N_4884,N_5896);
xnor U6328 (N_6328,N_5589,N_5981);
or U6329 (N_6329,N_5574,N_5205);
and U6330 (N_6330,N_4938,N_4541);
nand U6331 (N_6331,N_5563,N_4990);
or U6332 (N_6332,N_4766,N_4906);
xnor U6333 (N_6333,N_5958,N_5769);
nand U6334 (N_6334,N_5070,N_5102);
and U6335 (N_6335,N_4719,N_5405);
or U6336 (N_6336,N_4867,N_5558);
xor U6337 (N_6337,N_5207,N_4919);
and U6338 (N_6338,N_5249,N_5643);
and U6339 (N_6339,N_5613,N_5062);
nand U6340 (N_6340,N_5108,N_5474);
xnor U6341 (N_6341,N_5123,N_5871);
or U6342 (N_6342,N_4966,N_4926);
or U6343 (N_6343,N_4777,N_5195);
nor U6344 (N_6344,N_4908,N_5785);
nand U6345 (N_6345,N_4894,N_5376);
xnor U6346 (N_6346,N_5860,N_5815);
nand U6347 (N_6347,N_4572,N_5438);
or U6348 (N_6348,N_4700,N_4947);
xor U6349 (N_6349,N_4970,N_5294);
nand U6350 (N_6350,N_5139,N_4684);
or U6351 (N_6351,N_5986,N_4573);
nor U6352 (N_6352,N_4937,N_4850);
and U6353 (N_6353,N_5529,N_5079);
nor U6354 (N_6354,N_4803,N_4836);
or U6355 (N_6355,N_4647,N_5941);
xnor U6356 (N_6356,N_5452,N_5056);
nor U6357 (N_6357,N_5707,N_5336);
nand U6358 (N_6358,N_4812,N_5742);
xnor U6359 (N_6359,N_5278,N_5604);
or U6360 (N_6360,N_4561,N_4869);
xor U6361 (N_6361,N_4873,N_5532);
and U6362 (N_6362,N_5366,N_4759);
xnor U6363 (N_6363,N_5118,N_5665);
nand U6364 (N_6364,N_5343,N_4709);
and U6365 (N_6365,N_5895,N_5165);
nor U6366 (N_6366,N_5090,N_5520);
and U6367 (N_6367,N_5928,N_5236);
or U6368 (N_6368,N_5477,N_5013);
nand U6369 (N_6369,N_5391,N_5846);
or U6370 (N_6370,N_5308,N_4678);
or U6371 (N_6371,N_5523,N_5848);
or U6372 (N_6372,N_4941,N_4723);
and U6373 (N_6373,N_5993,N_4623);
xor U6374 (N_6374,N_5543,N_5821);
nor U6375 (N_6375,N_4597,N_5164);
and U6376 (N_6376,N_5350,N_5470);
xnor U6377 (N_6377,N_4833,N_5055);
and U6378 (N_6378,N_5219,N_5075);
nor U6379 (N_6379,N_5768,N_5583);
or U6380 (N_6380,N_5255,N_5624);
and U6381 (N_6381,N_5043,N_4579);
nand U6382 (N_6382,N_5607,N_5392);
nand U6383 (N_6383,N_5735,N_4645);
or U6384 (N_6384,N_5659,N_5978);
and U6385 (N_6385,N_5680,N_5802);
nand U6386 (N_6386,N_5940,N_5663);
nand U6387 (N_6387,N_5001,N_5572);
nor U6388 (N_6388,N_4864,N_5133);
nand U6389 (N_6389,N_5178,N_5631);
and U6390 (N_6390,N_4562,N_5284);
nand U6391 (N_6391,N_4539,N_5765);
xor U6392 (N_6392,N_5107,N_5652);
nand U6393 (N_6393,N_5957,N_5398);
and U6394 (N_6394,N_4920,N_5007);
and U6395 (N_6395,N_5639,N_5349);
nand U6396 (N_6396,N_4899,N_4968);
xor U6397 (N_6397,N_4948,N_4610);
nand U6398 (N_6398,N_5696,N_4809);
or U6399 (N_6399,N_4862,N_4835);
or U6400 (N_6400,N_5514,N_5969);
or U6401 (N_6401,N_4852,N_5717);
and U6402 (N_6402,N_5553,N_4502);
xor U6403 (N_6403,N_5416,N_5541);
xnor U6404 (N_6404,N_5488,N_4793);
nor U6405 (N_6405,N_5415,N_4827);
nand U6406 (N_6406,N_5443,N_4888);
nand U6407 (N_6407,N_4590,N_5436);
xnor U6408 (N_6408,N_4578,N_5212);
nand U6409 (N_6409,N_4857,N_5273);
xor U6410 (N_6410,N_5267,N_4782);
xor U6411 (N_6411,N_5265,N_5125);
nand U6412 (N_6412,N_5644,N_5733);
xor U6413 (N_6413,N_5408,N_5471);
xnor U6414 (N_6414,N_4995,N_5706);
xnor U6415 (N_6415,N_4526,N_4879);
and U6416 (N_6416,N_5384,N_5902);
nand U6417 (N_6417,N_5266,N_5159);
or U6418 (N_6418,N_5738,N_5310);
nand U6419 (N_6419,N_4787,N_5874);
nand U6420 (N_6420,N_5649,N_4959);
nor U6421 (N_6421,N_5701,N_5922);
nor U6422 (N_6422,N_5825,N_5412);
nor U6423 (N_6423,N_5357,N_5027);
or U6424 (N_6424,N_5798,N_5844);
nand U6425 (N_6425,N_5410,N_5111);
nand U6426 (N_6426,N_5720,N_5878);
xnor U6427 (N_6427,N_4917,N_5303);
and U6428 (N_6428,N_5456,N_4930);
or U6429 (N_6429,N_5926,N_5911);
nand U6430 (N_6430,N_5044,N_5741);
or U6431 (N_6431,N_5064,N_5806);
nand U6432 (N_6432,N_4625,N_5402);
and U6433 (N_6433,N_4923,N_5371);
nand U6434 (N_6434,N_4523,N_5327);
or U6435 (N_6435,N_4794,N_4591);
and U6436 (N_6436,N_5610,N_5063);
nor U6437 (N_6437,N_5400,N_4569);
nand U6438 (N_6438,N_4784,N_5637);
and U6439 (N_6439,N_5671,N_5430);
nand U6440 (N_6440,N_5634,N_5862);
and U6441 (N_6441,N_5632,N_5564);
or U6442 (N_6442,N_5100,N_5530);
or U6443 (N_6443,N_5128,N_5057);
xor U6444 (N_6444,N_4585,N_5225);
xor U6445 (N_6445,N_5021,N_5508);
nand U6446 (N_6446,N_5246,N_5237);
xor U6447 (N_6447,N_5478,N_5099);
and U6448 (N_6448,N_5850,N_5616);
or U6449 (N_6449,N_5221,N_4762);
nand U6450 (N_6450,N_5702,N_5485);
or U6451 (N_6451,N_4702,N_4944);
and U6452 (N_6452,N_5486,N_4960);
xnor U6453 (N_6453,N_4915,N_5241);
and U6454 (N_6454,N_5565,N_5080);
xnor U6455 (N_6455,N_4536,N_5344);
xor U6456 (N_6456,N_5296,N_5828);
and U6457 (N_6457,N_4534,N_5275);
nor U6458 (N_6458,N_5675,N_4741);
nor U6459 (N_6459,N_5146,N_5397);
nand U6460 (N_6460,N_4981,N_5752);
xor U6461 (N_6461,N_4517,N_5411);
nor U6462 (N_6462,N_5137,N_5288);
and U6463 (N_6463,N_5381,N_4556);
or U6464 (N_6464,N_4677,N_4669);
and U6465 (N_6465,N_5929,N_5213);
nor U6466 (N_6466,N_5756,N_4515);
nand U6467 (N_6467,N_4712,N_5976);
and U6468 (N_6468,N_5457,N_4513);
nor U6469 (N_6469,N_5867,N_4846);
nor U6470 (N_6470,N_5513,N_4577);
and U6471 (N_6471,N_5927,N_4949);
and U6472 (N_6472,N_5014,N_5714);
nand U6473 (N_6473,N_4753,N_4511);
nand U6474 (N_6474,N_5148,N_5868);
and U6475 (N_6475,N_5377,N_4553);
or U6476 (N_6476,N_4963,N_5640);
nand U6477 (N_6477,N_5931,N_5222);
and U6478 (N_6478,N_4598,N_4828);
or U6479 (N_6479,N_5446,N_5537);
or U6480 (N_6480,N_4593,N_5762);
nor U6481 (N_6481,N_5598,N_5499);
xor U6482 (N_6482,N_4636,N_5234);
nor U6483 (N_6483,N_5244,N_5504);
and U6484 (N_6484,N_4584,N_4640);
or U6485 (N_6485,N_5109,N_5791);
nor U6486 (N_6486,N_4986,N_4786);
nor U6487 (N_6487,N_5811,N_5712);
or U6488 (N_6488,N_5827,N_5431);
nand U6489 (N_6489,N_4646,N_5132);
and U6490 (N_6490,N_5804,N_4648);
or U6491 (N_6491,N_5588,N_4755);
nor U6492 (N_6492,N_4918,N_5704);
and U6493 (N_6493,N_5053,N_5542);
xnor U6494 (N_6494,N_4582,N_5089);
nor U6495 (N_6495,N_5115,N_5839);
or U6496 (N_6496,N_4697,N_5780);
or U6497 (N_6497,N_5489,N_5876);
or U6498 (N_6498,N_5942,N_5276);
or U6499 (N_6499,N_5147,N_5753);
or U6500 (N_6500,N_5295,N_4855);
and U6501 (N_6501,N_5029,N_5369);
nand U6502 (N_6502,N_5023,N_5259);
nand U6503 (N_6503,N_5809,N_5012);
xnor U6504 (N_6504,N_4694,N_5518);
nor U6505 (N_6505,N_5065,N_4683);
xnor U6506 (N_6506,N_5383,N_5647);
or U6507 (N_6507,N_5472,N_4632);
xnor U6508 (N_6508,N_4671,N_4612);
and U6509 (N_6509,N_5379,N_4735);
or U6510 (N_6510,N_5865,N_4727);
xnor U6511 (N_6511,N_4813,N_5142);
and U6512 (N_6512,N_5110,N_4736);
nor U6513 (N_6513,N_4552,N_5286);
and U6514 (N_6514,N_5018,N_4815);
nand U6515 (N_6515,N_4503,N_4865);
and U6516 (N_6516,N_4696,N_4844);
or U6517 (N_6517,N_5097,N_5881);
or U6518 (N_6518,N_5578,N_5751);
or U6519 (N_6519,N_5669,N_5590);
xor U6520 (N_6520,N_5130,N_4501);
and U6521 (N_6521,N_5484,N_4951);
or U6522 (N_6522,N_5546,N_5353);
or U6523 (N_6523,N_5599,N_5226);
or U6524 (N_6524,N_4525,N_4889);
nand U6525 (N_6525,N_4962,N_4985);
xnor U6526 (N_6526,N_5321,N_5740);
or U6527 (N_6527,N_4546,N_5535);
xnor U6528 (N_6528,N_5387,N_4543);
nor U6529 (N_6529,N_5481,N_5863);
xnor U6530 (N_6530,N_5573,N_4558);
nor U6531 (N_6531,N_5716,N_4725);
and U6532 (N_6532,N_5552,N_4890);
nor U6533 (N_6533,N_4977,N_4853);
nor U6534 (N_6534,N_5678,N_5262);
xor U6535 (N_6535,N_5413,N_5492);
nor U6536 (N_6536,N_5252,N_4958);
or U6537 (N_6537,N_4933,N_5464);
and U6538 (N_6538,N_5576,N_4670);
and U6539 (N_6539,N_5952,N_5914);
nor U6540 (N_6540,N_5890,N_4627);
and U6541 (N_6541,N_4724,N_5781);
and U6542 (N_6542,N_5467,N_5857);
and U6543 (N_6543,N_4826,N_5688);
nand U6544 (N_6544,N_5602,N_4656);
or U6545 (N_6545,N_5547,N_5538);
nor U6546 (N_6546,N_5534,N_5889);
or U6547 (N_6547,N_5924,N_4688);
nand U6548 (N_6548,N_4905,N_5315);
nand U6549 (N_6549,N_5776,N_4791);
and U6550 (N_6550,N_5188,N_5186);
or U6551 (N_6551,N_5365,N_4581);
nand U6552 (N_6552,N_4775,N_5817);
nand U6553 (N_6553,N_5016,N_5620);
nand U6554 (N_6554,N_5264,N_5505);
nand U6555 (N_6555,N_5386,N_5519);
and U6556 (N_6556,N_4921,N_5347);
or U6557 (N_6557,N_5866,N_5289);
and U6558 (N_6558,N_4871,N_4785);
or U6559 (N_6559,N_5215,N_4691);
nor U6560 (N_6560,N_5971,N_5052);
and U6561 (N_6561,N_5947,N_5673);
or U6562 (N_6562,N_5594,N_5754);
or U6563 (N_6563,N_5341,N_5937);
nor U6564 (N_6564,N_5091,N_4635);
xor U6565 (N_6565,N_5953,N_4706);
nor U6566 (N_6566,N_4565,N_4679);
or U6567 (N_6567,N_5545,N_5803);
xor U6568 (N_6568,N_5540,N_5210);
nor U6569 (N_6569,N_4863,N_4682);
nand U6570 (N_6570,N_4617,N_5041);
nor U6571 (N_6571,N_5679,N_5617);
nand U6572 (N_6572,N_5277,N_5009);
and U6573 (N_6573,N_4788,N_5409);
and U6574 (N_6574,N_4961,N_5316);
or U6575 (N_6575,N_5428,N_4666);
or U6576 (N_6576,N_5074,N_5960);
and U6577 (N_6577,N_5872,N_4542);
xor U6578 (N_6578,N_5744,N_5915);
nand U6579 (N_6579,N_5404,N_5654);
or U6580 (N_6580,N_4531,N_5531);
nand U6581 (N_6581,N_5025,N_4540);
xor U6582 (N_6582,N_5612,N_4772);
and U6583 (N_6583,N_5912,N_5036);
xor U6584 (N_6584,N_5242,N_5737);
nand U6585 (N_6585,N_5224,N_5483);
xor U6586 (N_6586,N_4644,N_5189);
and U6587 (N_6587,N_5260,N_5447);
or U6588 (N_6588,N_4928,N_5346);
nor U6589 (N_6589,N_5245,N_5525);
xor U6590 (N_6590,N_5936,N_5335);
nor U6591 (N_6591,N_4568,N_4956);
nand U6592 (N_6592,N_5636,N_5651);
or U6593 (N_6593,N_5511,N_5406);
or U6594 (N_6594,N_5968,N_5550);
nor U6595 (N_6595,N_5285,N_5909);
xor U6596 (N_6596,N_5389,N_5885);
nor U6597 (N_6597,N_5832,N_5766);
and U6598 (N_6598,N_4667,N_4916);
or U6599 (N_6599,N_5919,N_5407);
nor U6600 (N_6600,N_4760,N_4776);
or U6601 (N_6601,N_5455,N_5660);
and U6602 (N_6602,N_4988,N_5274);
or U6603 (N_6603,N_5801,N_5206);
nor U6604 (N_6604,N_5773,N_5943);
nand U6605 (N_6605,N_4680,N_5622);
nor U6606 (N_6606,N_4718,N_4974);
nor U6607 (N_6607,N_5441,N_5708);
xnor U6608 (N_6608,N_5324,N_4770);
nand U6609 (N_6609,N_5861,N_4975);
and U6610 (N_6610,N_5329,N_5328);
nand U6611 (N_6611,N_5853,N_5176);
or U6612 (N_6612,N_4881,N_5218);
nand U6613 (N_6613,N_5433,N_5951);
xnor U6614 (N_6614,N_4946,N_4750);
nand U6615 (N_6615,N_5835,N_5842);
or U6616 (N_6616,N_5240,N_5356);
or U6617 (N_6617,N_4685,N_4952);
or U6618 (N_6618,N_5345,N_4521);
and U6619 (N_6619,N_5076,N_5657);
or U6620 (N_6620,N_4551,N_5301);
xnor U6621 (N_6621,N_5887,N_4880);
nor U6622 (N_6622,N_5072,N_5760);
xnor U6623 (N_6623,N_4628,N_5510);
and U6624 (N_6624,N_5796,N_4527);
nor U6625 (N_6625,N_5432,N_4533);
nand U6626 (N_6626,N_5180,N_4798);
nand U6627 (N_6627,N_5648,N_5687);
or U6628 (N_6628,N_5870,N_5619);
nand U6629 (N_6629,N_5587,N_4875);
or U6630 (N_6630,N_5582,N_5512);
or U6631 (N_6631,N_5425,N_4567);
nand U6632 (N_6632,N_5794,N_5331);
nor U6633 (N_6633,N_4586,N_5334);
or U6634 (N_6634,N_4653,N_4743);
nand U6635 (N_6635,N_5311,N_5194);
and U6636 (N_6636,N_5788,N_4566);
nor U6637 (N_6637,N_5182,N_4790);
or U6638 (N_6638,N_5454,N_5502);
nand U6639 (N_6639,N_5120,N_5269);
and U6640 (N_6640,N_5468,N_5058);
nand U6641 (N_6641,N_5608,N_4518);
nand U6642 (N_6642,N_5011,N_5473);
or U6643 (N_6643,N_5462,N_4673);
or U6644 (N_6644,N_5293,N_5360);
xor U6645 (N_6645,N_5152,N_4874);
or U6646 (N_6646,N_4859,N_4860);
nor U6647 (N_6647,N_4955,N_5998);
nor U6648 (N_6648,N_4664,N_4729);
nor U6649 (N_6649,N_5823,N_4739);
or U6650 (N_6650,N_4768,N_5220);
nand U6651 (N_6651,N_5302,N_4999);
and U6652 (N_6652,N_5670,N_5395);
xor U6653 (N_6653,N_4538,N_5054);
xor U6654 (N_6654,N_5268,N_5757);
or U6655 (N_6655,N_5987,N_5103);
nand U6656 (N_6656,N_5646,N_5348);
nand U6657 (N_6657,N_4728,N_5797);
nor U6658 (N_6658,N_4902,N_4845);
xor U6659 (N_6659,N_5528,N_5903);
nor U6660 (N_6660,N_5476,N_4901);
and U6661 (N_6661,N_5959,N_5567);
and U6662 (N_6662,N_5459,N_5449);
nand U6663 (N_6663,N_4763,N_5627);
xor U6664 (N_6664,N_4754,N_4757);
xnor U6665 (N_6665,N_4771,N_5509);
or U6666 (N_6666,N_4843,N_5175);
xor U6667 (N_6667,N_5856,N_4746);
nor U6668 (N_6668,N_5192,N_5444);
or U6669 (N_6669,N_5038,N_5117);
or U6670 (N_6670,N_4744,N_5807);
and U6671 (N_6671,N_5908,N_5763);
nand U6672 (N_6672,N_5560,N_5337);
nor U6673 (N_6673,N_5190,N_5611);
or U6674 (N_6674,N_5521,N_5270);
nor U6675 (N_6675,N_5393,N_5209);
xor U6676 (N_6676,N_5035,N_5703);
nor U6677 (N_6677,N_4994,N_5078);
nor U6678 (N_6678,N_4619,N_5595);
nand U6679 (N_6679,N_5465,N_5045);
nor U6680 (N_6680,N_5501,N_5779);
nor U6681 (N_6681,N_5067,N_5593);
or U6682 (N_6682,N_5151,N_5755);
or U6683 (N_6683,N_4686,N_5786);
nor U6684 (N_6684,N_5322,N_4535);
nor U6685 (N_6685,N_5475,N_5826);
and U6686 (N_6686,N_5401,N_4698);
nor U6687 (N_6687,N_4957,N_5030);
or U6688 (N_6688,N_5248,N_4807);
nand U6689 (N_6689,N_5609,N_4907);
and U6690 (N_6690,N_4532,N_5280);
and U6691 (N_6691,N_4856,N_5362);
nor U6692 (N_6692,N_4954,N_5913);
xnor U6693 (N_6693,N_5419,N_5661);
and U6694 (N_6694,N_5586,N_5060);
or U6695 (N_6695,N_5917,N_5690);
nand U6696 (N_6696,N_4547,N_4774);
or U6697 (N_6697,N_5772,N_5533);
xor U6698 (N_6698,N_5144,N_5879);
or U6699 (N_6699,N_4831,N_5149);
nand U6700 (N_6700,N_4594,N_5326);
or U6701 (N_6701,N_5469,N_5731);
or U6702 (N_6702,N_5750,N_5094);
and U6703 (N_6703,N_4973,N_5171);
nand U6704 (N_6704,N_5745,N_5747);
nand U6705 (N_6705,N_5230,N_5854);
or U6706 (N_6706,N_5606,N_5367);
or U6707 (N_6707,N_5635,N_5258);
xnor U6708 (N_6708,N_5526,N_4560);
or U6709 (N_6709,N_4714,N_5004);
or U6710 (N_6710,N_5403,N_5361);
or U6711 (N_6711,N_4767,N_5422);
xor U6712 (N_6712,N_5161,N_5729);
or U6713 (N_6713,N_5562,N_5380);
xor U6714 (N_6714,N_5048,N_4931);
xnor U6715 (N_6715,N_5127,N_4699);
nand U6716 (N_6716,N_5093,N_5810);
or U6717 (N_6717,N_5764,N_4893);
xnor U6718 (N_6718,N_4720,N_4822);
nor U6719 (N_6719,N_4693,N_5239);
or U6720 (N_6720,N_5677,N_4516);
nor U6721 (N_6721,N_5556,N_4989);
or U6722 (N_6722,N_5493,N_4752);
nor U6723 (N_6723,N_5829,N_4903);
nand U6724 (N_6724,N_5883,N_4674);
xor U6725 (N_6725,N_5568,N_5691);
nand U6726 (N_6726,N_5561,N_5162);
xnor U6727 (N_6727,N_5633,N_4911);
or U6728 (N_6728,N_5900,N_4982);
nor U6729 (N_6729,N_4769,N_5603);
xnor U6730 (N_6730,N_5440,N_5168);
nor U6731 (N_6731,N_4979,N_5358);
or U6732 (N_6732,N_5837,N_5858);
xnor U6733 (N_6733,N_5693,N_4991);
xnor U6734 (N_6734,N_4861,N_4830);
nand U6735 (N_6735,N_4675,N_4630);
nand U6736 (N_6736,N_4596,N_5006);
nor U6737 (N_6737,N_5580,N_5202);
and U6738 (N_6738,N_4998,N_5101);
xor U6739 (N_6739,N_5630,N_5650);
or U6740 (N_6740,N_5864,N_5253);
and U6741 (N_6741,N_4522,N_4530);
nor U6742 (N_6742,N_5223,N_5307);
xor U6743 (N_6743,N_4733,N_4559);
xor U6744 (N_6744,N_5984,N_5167);
xor U6745 (N_6745,N_5591,N_5566);
xnor U6746 (N_6746,N_5024,N_4639);
nand U6747 (N_6747,N_5032,N_5551);
or U6748 (N_6748,N_5967,N_5939);
xnor U6749 (N_6749,N_4545,N_5905);
or U6750 (N_6750,N_4898,N_5314);
or U6751 (N_6751,N_5151,N_5243);
or U6752 (N_6752,N_5067,N_4926);
and U6753 (N_6753,N_4602,N_4724);
or U6754 (N_6754,N_4591,N_5710);
xor U6755 (N_6755,N_4819,N_5993);
xor U6756 (N_6756,N_5621,N_5731);
or U6757 (N_6757,N_5448,N_4973);
and U6758 (N_6758,N_5822,N_5038);
or U6759 (N_6759,N_5025,N_4648);
nor U6760 (N_6760,N_5041,N_4706);
and U6761 (N_6761,N_5901,N_5177);
or U6762 (N_6762,N_5709,N_5263);
or U6763 (N_6763,N_5522,N_4558);
or U6764 (N_6764,N_5236,N_5644);
and U6765 (N_6765,N_5115,N_5821);
or U6766 (N_6766,N_5989,N_5946);
nand U6767 (N_6767,N_5436,N_5811);
and U6768 (N_6768,N_5226,N_5812);
nor U6769 (N_6769,N_5175,N_4641);
nor U6770 (N_6770,N_4692,N_5533);
xor U6771 (N_6771,N_5163,N_5149);
nand U6772 (N_6772,N_5454,N_5351);
or U6773 (N_6773,N_5807,N_4884);
xnor U6774 (N_6774,N_5780,N_5187);
and U6775 (N_6775,N_5776,N_4613);
or U6776 (N_6776,N_5097,N_4862);
nor U6777 (N_6777,N_4860,N_5536);
or U6778 (N_6778,N_5408,N_4957);
nor U6779 (N_6779,N_5866,N_5299);
nand U6780 (N_6780,N_4860,N_4500);
nor U6781 (N_6781,N_5405,N_5258);
nand U6782 (N_6782,N_5851,N_5394);
xnor U6783 (N_6783,N_5053,N_5021);
and U6784 (N_6784,N_5418,N_5895);
nor U6785 (N_6785,N_4639,N_4726);
and U6786 (N_6786,N_4591,N_5910);
nor U6787 (N_6787,N_4978,N_4933);
and U6788 (N_6788,N_5889,N_4798);
or U6789 (N_6789,N_5874,N_4661);
nand U6790 (N_6790,N_5778,N_5314);
and U6791 (N_6791,N_5152,N_5574);
and U6792 (N_6792,N_5515,N_5728);
and U6793 (N_6793,N_4797,N_5345);
or U6794 (N_6794,N_5028,N_5407);
xor U6795 (N_6795,N_4869,N_5890);
and U6796 (N_6796,N_5972,N_4871);
nand U6797 (N_6797,N_5582,N_5432);
and U6798 (N_6798,N_5580,N_4620);
xnor U6799 (N_6799,N_5824,N_5229);
xnor U6800 (N_6800,N_4909,N_4863);
nor U6801 (N_6801,N_5124,N_5566);
xnor U6802 (N_6802,N_5013,N_4701);
nand U6803 (N_6803,N_5787,N_5922);
nor U6804 (N_6804,N_5638,N_4724);
nor U6805 (N_6805,N_5347,N_5999);
and U6806 (N_6806,N_4695,N_5788);
and U6807 (N_6807,N_5233,N_5751);
nor U6808 (N_6808,N_5654,N_4774);
and U6809 (N_6809,N_5501,N_5517);
or U6810 (N_6810,N_5510,N_5395);
xor U6811 (N_6811,N_5752,N_4784);
nand U6812 (N_6812,N_4649,N_4596);
and U6813 (N_6813,N_5043,N_4970);
xnor U6814 (N_6814,N_5555,N_5015);
or U6815 (N_6815,N_5128,N_5929);
or U6816 (N_6816,N_5649,N_4728);
and U6817 (N_6817,N_5425,N_5921);
xnor U6818 (N_6818,N_5930,N_5953);
xor U6819 (N_6819,N_5746,N_4798);
or U6820 (N_6820,N_4616,N_4602);
and U6821 (N_6821,N_5719,N_4546);
xor U6822 (N_6822,N_4957,N_4847);
xor U6823 (N_6823,N_5803,N_4930);
nor U6824 (N_6824,N_4696,N_5518);
nand U6825 (N_6825,N_5554,N_4667);
or U6826 (N_6826,N_4536,N_5647);
or U6827 (N_6827,N_5216,N_5605);
or U6828 (N_6828,N_5811,N_5982);
or U6829 (N_6829,N_4552,N_5017);
nand U6830 (N_6830,N_5958,N_5412);
or U6831 (N_6831,N_5802,N_5033);
and U6832 (N_6832,N_5129,N_5711);
or U6833 (N_6833,N_5147,N_5828);
or U6834 (N_6834,N_4859,N_4746);
xor U6835 (N_6835,N_4625,N_5469);
and U6836 (N_6836,N_4559,N_5482);
or U6837 (N_6837,N_5779,N_5108);
or U6838 (N_6838,N_5312,N_4880);
or U6839 (N_6839,N_4978,N_5335);
xnor U6840 (N_6840,N_5780,N_4754);
nor U6841 (N_6841,N_5623,N_5958);
and U6842 (N_6842,N_5872,N_4531);
xnor U6843 (N_6843,N_5813,N_5049);
xor U6844 (N_6844,N_5929,N_5071);
xor U6845 (N_6845,N_5222,N_5088);
or U6846 (N_6846,N_4575,N_5695);
nor U6847 (N_6847,N_4504,N_4624);
and U6848 (N_6848,N_5499,N_4984);
or U6849 (N_6849,N_4619,N_4743);
and U6850 (N_6850,N_4638,N_4526);
nor U6851 (N_6851,N_5111,N_5571);
xnor U6852 (N_6852,N_4697,N_5869);
and U6853 (N_6853,N_5801,N_5230);
and U6854 (N_6854,N_4913,N_5579);
and U6855 (N_6855,N_4847,N_4921);
and U6856 (N_6856,N_5001,N_5574);
xor U6857 (N_6857,N_5973,N_5199);
nor U6858 (N_6858,N_5417,N_5248);
and U6859 (N_6859,N_4940,N_4913);
nand U6860 (N_6860,N_4990,N_4986);
or U6861 (N_6861,N_5688,N_4626);
or U6862 (N_6862,N_5191,N_5829);
nand U6863 (N_6863,N_5622,N_5423);
and U6864 (N_6864,N_5643,N_5273);
and U6865 (N_6865,N_5043,N_4895);
or U6866 (N_6866,N_5829,N_4741);
nor U6867 (N_6867,N_5903,N_5025);
nand U6868 (N_6868,N_5895,N_5686);
and U6869 (N_6869,N_5121,N_4537);
nor U6870 (N_6870,N_5980,N_5314);
nor U6871 (N_6871,N_5130,N_5449);
or U6872 (N_6872,N_5439,N_5710);
nor U6873 (N_6873,N_4704,N_5818);
nor U6874 (N_6874,N_5922,N_5375);
or U6875 (N_6875,N_4721,N_5049);
xor U6876 (N_6876,N_4744,N_4562);
xnor U6877 (N_6877,N_5325,N_5930);
nand U6878 (N_6878,N_5343,N_4810);
nor U6879 (N_6879,N_5620,N_5657);
nor U6880 (N_6880,N_4762,N_5384);
nor U6881 (N_6881,N_5580,N_4526);
xor U6882 (N_6882,N_5626,N_5111);
and U6883 (N_6883,N_5667,N_5732);
xnor U6884 (N_6884,N_4535,N_5955);
and U6885 (N_6885,N_5480,N_4805);
nand U6886 (N_6886,N_5974,N_5152);
nand U6887 (N_6887,N_5123,N_5551);
and U6888 (N_6888,N_5726,N_5458);
nor U6889 (N_6889,N_4889,N_4537);
nand U6890 (N_6890,N_5324,N_4645);
and U6891 (N_6891,N_5504,N_4810);
or U6892 (N_6892,N_5893,N_5239);
nor U6893 (N_6893,N_5768,N_5816);
or U6894 (N_6894,N_5982,N_5705);
nand U6895 (N_6895,N_5138,N_5044);
and U6896 (N_6896,N_5255,N_4925);
nand U6897 (N_6897,N_4669,N_5379);
nand U6898 (N_6898,N_4920,N_5565);
and U6899 (N_6899,N_4853,N_5635);
and U6900 (N_6900,N_5052,N_5264);
nand U6901 (N_6901,N_4643,N_4548);
xor U6902 (N_6902,N_4592,N_5712);
nand U6903 (N_6903,N_5394,N_5655);
nand U6904 (N_6904,N_5556,N_5828);
or U6905 (N_6905,N_5637,N_4949);
and U6906 (N_6906,N_5374,N_5687);
nor U6907 (N_6907,N_4956,N_5961);
nor U6908 (N_6908,N_5807,N_5748);
or U6909 (N_6909,N_5921,N_5470);
nand U6910 (N_6910,N_4790,N_5388);
or U6911 (N_6911,N_5286,N_5548);
nor U6912 (N_6912,N_5691,N_5150);
nand U6913 (N_6913,N_4506,N_5523);
nand U6914 (N_6914,N_5065,N_5690);
nor U6915 (N_6915,N_4699,N_5803);
nor U6916 (N_6916,N_5040,N_5967);
nand U6917 (N_6917,N_5190,N_5296);
nor U6918 (N_6918,N_5007,N_5475);
or U6919 (N_6919,N_5244,N_5649);
nor U6920 (N_6920,N_5694,N_4828);
and U6921 (N_6921,N_4710,N_5452);
or U6922 (N_6922,N_5702,N_4589);
nor U6923 (N_6923,N_5796,N_4889);
or U6924 (N_6924,N_5804,N_4805);
or U6925 (N_6925,N_5915,N_5633);
nand U6926 (N_6926,N_5869,N_5754);
nor U6927 (N_6927,N_4659,N_5133);
and U6928 (N_6928,N_4533,N_5113);
and U6929 (N_6929,N_5832,N_4762);
nand U6930 (N_6930,N_5463,N_4887);
xnor U6931 (N_6931,N_5668,N_4637);
and U6932 (N_6932,N_5047,N_5158);
and U6933 (N_6933,N_5682,N_5315);
and U6934 (N_6934,N_5149,N_4787);
or U6935 (N_6935,N_4941,N_5493);
xor U6936 (N_6936,N_5541,N_5116);
or U6937 (N_6937,N_5027,N_5399);
or U6938 (N_6938,N_5622,N_5778);
and U6939 (N_6939,N_4743,N_4698);
nor U6940 (N_6940,N_4952,N_5258);
nor U6941 (N_6941,N_4723,N_5359);
and U6942 (N_6942,N_5492,N_5019);
xor U6943 (N_6943,N_5459,N_5318);
nor U6944 (N_6944,N_5731,N_5068);
or U6945 (N_6945,N_5519,N_5339);
and U6946 (N_6946,N_5658,N_5066);
nor U6947 (N_6947,N_5173,N_5839);
nand U6948 (N_6948,N_5562,N_4638);
nand U6949 (N_6949,N_4636,N_4506);
nor U6950 (N_6950,N_5967,N_5881);
nor U6951 (N_6951,N_5026,N_5400);
xnor U6952 (N_6952,N_5941,N_4608);
or U6953 (N_6953,N_5024,N_5066);
or U6954 (N_6954,N_4743,N_5122);
xnor U6955 (N_6955,N_5927,N_4711);
and U6956 (N_6956,N_4758,N_4836);
nand U6957 (N_6957,N_5324,N_5980);
xnor U6958 (N_6958,N_5063,N_4841);
xor U6959 (N_6959,N_4850,N_5761);
nand U6960 (N_6960,N_5803,N_5528);
nor U6961 (N_6961,N_5471,N_5444);
and U6962 (N_6962,N_5022,N_5573);
xor U6963 (N_6963,N_4668,N_4692);
xor U6964 (N_6964,N_4914,N_5973);
nor U6965 (N_6965,N_5138,N_5724);
xnor U6966 (N_6966,N_5480,N_4970);
nor U6967 (N_6967,N_5421,N_5342);
or U6968 (N_6968,N_5358,N_5223);
and U6969 (N_6969,N_5477,N_5347);
and U6970 (N_6970,N_4914,N_4610);
xnor U6971 (N_6971,N_5486,N_5145);
or U6972 (N_6972,N_5030,N_4503);
nor U6973 (N_6973,N_4872,N_5948);
xor U6974 (N_6974,N_5287,N_4828);
nor U6975 (N_6975,N_5549,N_5622);
and U6976 (N_6976,N_5538,N_5980);
nor U6977 (N_6977,N_4542,N_5351);
nor U6978 (N_6978,N_5011,N_4805);
and U6979 (N_6979,N_5396,N_5032);
and U6980 (N_6980,N_5849,N_5699);
nand U6981 (N_6981,N_5229,N_5822);
nor U6982 (N_6982,N_5763,N_5444);
nand U6983 (N_6983,N_4959,N_5594);
nor U6984 (N_6984,N_4825,N_4638);
xor U6985 (N_6985,N_5348,N_5543);
nor U6986 (N_6986,N_5655,N_5466);
or U6987 (N_6987,N_5587,N_4891);
xnor U6988 (N_6988,N_5680,N_4613);
xor U6989 (N_6989,N_4639,N_4649);
xor U6990 (N_6990,N_4871,N_5696);
nor U6991 (N_6991,N_4596,N_5717);
xnor U6992 (N_6992,N_4573,N_4987);
nor U6993 (N_6993,N_5370,N_5122);
nor U6994 (N_6994,N_5792,N_4647);
nor U6995 (N_6995,N_5376,N_4923);
or U6996 (N_6996,N_5458,N_5272);
or U6997 (N_6997,N_5356,N_5806);
nand U6998 (N_6998,N_4871,N_5683);
and U6999 (N_6999,N_5855,N_4505);
xor U7000 (N_7000,N_4627,N_5857);
xnor U7001 (N_7001,N_5783,N_4674);
xor U7002 (N_7002,N_4778,N_5897);
or U7003 (N_7003,N_5080,N_5966);
xnor U7004 (N_7004,N_4676,N_4571);
or U7005 (N_7005,N_5178,N_4922);
nor U7006 (N_7006,N_5188,N_5294);
nor U7007 (N_7007,N_5995,N_5261);
xor U7008 (N_7008,N_4819,N_4799);
nor U7009 (N_7009,N_4831,N_5990);
nand U7010 (N_7010,N_5337,N_5157);
xor U7011 (N_7011,N_5181,N_5867);
xnor U7012 (N_7012,N_4856,N_5478);
or U7013 (N_7013,N_5593,N_5817);
nor U7014 (N_7014,N_5797,N_5997);
xnor U7015 (N_7015,N_4567,N_4976);
and U7016 (N_7016,N_5984,N_5939);
or U7017 (N_7017,N_5817,N_5944);
or U7018 (N_7018,N_4903,N_5737);
or U7019 (N_7019,N_5217,N_4650);
xor U7020 (N_7020,N_5604,N_4941);
and U7021 (N_7021,N_4950,N_4897);
or U7022 (N_7022,N_5045,N_5908);
nand U7023 (N_7023,N_5498,N_5200);
nand U7024 (N_7024,N_5291,N_5341);
or U7025 (N_7025,N_5309,N_5455);
nand U7026 (N_7026,N_5167,N_5964);
and U7027 (N_7027,N_5508,N_5316);
and U7028 (N_7028,N_5326,N_5006);
nor U7029 (N_7029,N_5142,N_4617);
and U7030 (N_7030,N_5960,N_5113);
nand U7031 (N_7031,N_4829,N_4629);
nor U7032 (N_7032,N_5869,N_5494);
or U7033 (N_7033,N_5760,N_4904);
nor U7034 (N_7034,N_5892,N_5610);
and U7035 (N_7035,N_5427,N_4807);
nand U7036 (N_7036,N_5459,N_4773);
xnor U7037 (N_7037,N_4777,N_5715);
nand U7038 (N_7038,N_5221,N_5679);
nand U7039 (N_7039,N_5264,N_4793);
or U7040 (N_7040,N_5804,N_5045);
or U7041 (N_7041,N_5853,N_5064);
nor U7042 (N_7042,N_4886,N_5967);
or U7043 (N_7043,N_5072,N_5410);
and U7044 (N_7044,N_5777,N_4711);
or U7045 (N_7045,N_5849,N_4549);
nor U7046 (N_7046,N_5711,N_4721);
or U7047 (N_7047,N_4518,N_5768);
or U7048 (N_7048,N_5505,N_4960);
and U7049 (N_7049,N_5034,N_4977);
and U7050 (N_7050,N_5346,N_4541);
or U7051 (N_7051,N_4827,N_5305);
xor U7052 (N_7052,N_5629,N_4794);
nor U7053 (N_7053,N_4971,N_5850);
nand U7054 (N_7054,N_5886,N_5261);
nor U7055 (N_7055,N_4622,N_5780);
nor U7056 (N_7056,N_4670,N_5368);
nand U7057 (N_7057,N_5256,N_4948);
nand U7058 (N_7058,N_5938,N_4586);
nand U7059 (N_7059,N_5899,N_5850);
nor U7060 (N_7060,N_4668,N_5057);
nand U7061 (N_7061,N_5268,N_5701);
xnor U7062 (N_7062,N_4987,N_4536);
xor U7063 (N_7063,N_4780,N_5749);
nor U7064 (N_7064,N_4641,N_5378);
and U7065 (N_7065,N_5619,N_5215);
nand U7066 (N_7066,N_5854,N_5196);
nand U7067 (N_7067,N_4928,N_4858);
xnor U7068 (N_7068,N_4554,N_5985);
or U7069 (N_7069,N_4781,N_4962);
or U7070 (N_7070,N_4753,N_4945);
nor U7071 (N_7071,N_5962,N_5598);
nand U7072 (N_7072,N_5552,N_5692);
and U7073 (N_7073,N_5031,N_5029);
or U7074 (N_7074,N_4768,N_5174);
nand U7075 (N_7075,N_5633,N_4979);
xor U7076 (N_7076,N_4818,N_4673);
and U7077 (N_7077,N_5846,N_4613);
xor U7078 (N_7078,N_5860,N_4591);
nor U7079 (N_7079,N_5860,N_5511);
xor U7080 (N_7080,N_4946,N_5141);
or U7081 (N_7081,N_4949,N_5902);
and U7082 (N_7082,N_4747,N_4504);
and U7083 (N_7083,N_4592,N_5046);
or U7084 (N_7084,N_4942,N_5203);
and U7085 (N_7085,N_5702,N_5866);
xor U7086 (N_7086,N_5656,N_5449);
or U7087 (N_7087,N_5583,N_5059);
nor U7088 (N_7088,N_4777,N_5998);
nand U7089 (N_7089,N_5621,N_4530);
or U7090 (N_7090,N_5020,N_5192);
nand U7091 (N_7091,N_5306,N_5760);
nand U7092 (N_7092,N_5113,N_5296);
nand U7093 (N_7093,N_5411,N_5729);
nor U7094 (N_7094,N_5133,N_4845);
and U7095 (N_7095,N_4827,N_5360);
nor U7096 (N_7096,N_5311,N_5839);
nor U7097 (N_7097,N_4873,N_5329);
nor U7098 (N_7098,N_5952,N_5535);
xnor U7099 (N_7099,N_4721,N_5055);
and U7100 (N_7100,N_5025,N_4550);
and U7101 (N_7101,N_4949,N_4933);
nor U7102 (N_7102,N_5738,N_5846);
xor U7103 (N_7103,N_5210,N_5891);
nand U7104 (N_7104,N_5293,N_5398);
and U7105 (N_7105,N_5914,N_5460);
or U7106 (N_7106,N_4686,N_5863);
or U7107 (N_7107,N_5896,N_5228);
nand U7108 (N_7108,N_4788,N_4539);
nor U7109 (N_7109,N_4689,N_4666);
nor U7110 (N_7110,N_5193,N_4824);
xnor U7111 (N_7111,N_4660,N_5286);
nor U7112 (N_7112,N_4995,N_5209);
nor U7113 (N_7113,N_4891,N_5483);
and U7114 (N_7114,N_5249,N_5028);
or U7115 (N_7115,N_5515,N_4630);
xnor U7116 (N_7116,N_5979,N_4837);
nand U7117 (N_7117,N_5818,N_5420);
and U7118 (N_7118,N_5608,N_5986);
nor U7119 (N_7119,N_5785,N_5381);
xnor U7120 (N_7120,N_5764,N_4883);
nor U7121 (N_7121,N_5734,N_5406);
and U7122 (N_7122,N_4874,N_5797);
nand U7123 (N_7123,N_5345,N_4747);
and U7124 (N_7124,N_5099,N_5661);
or U7125 (N_7125,N_5008,N_5342);
nor U7126 (N_7126,N_4755,N_5345);
nand U7127 (N_7127,N_4500,N_4919);
xnor U7128 (N_7128,N_4693,N_5684);
nand U7129 (N_7129,N_5154,N_5698);
nand U7130 (N_7130,N_5716,N_5347);
and U7131 (N_7131,N_5315,N_5320);
xor U7132 (N_7132,N_5118,N_5762);
nand U7133 (N_7133,N_5307,N_5085);
and U7134 (N_7134,N_5022,N_5667);
xnor U7135 (N_7135,N_5876,N_4764);
and U7136 (N_7136,N_5821,N_4950);
nor U7137 (N_7137,N_4790,N_4941);
and U7138 (N_7138,N_4860,N_4745);
nand U7139 (N_7139,N_4884,N_4693);
xnor U7140 (N_7140,N_5879,N_5178);
or U7141 (N_7141,N_4520,N_5867);
nor U7142 (N_7142,N_5580,N_5051);
or U7143 (N_7143,N_5935,N_5922);
nand U7144 (N_7144,N_5886,N_5085);
or U7145 (N_7145,N_5813,N_5374);
nor U7146 (N_7146,N_5109,N_4996);
nand U7147 (N_7147,N_5572,N_5682);
or U7148 (N_7148,N_4917,N_4690);
nand U7149 (N_7149,N_5261,N_5379);
nor U7150 (N_7150,N_4871,N_5866);
nand U7151 (N_7151,N_4942,N_5580);
nand U7152 (N_7152,N_4873,N_5279);
nor U7153 (N_7153,N_5475,N_5512);
xnor U7154 (N_7154,N_5668,N_5976);
nand U7155 (N_7155,N_5793,N_4524);
or U7156 (N_7156,N_4508,N_5867);
nand U7157 (N_7157,N_5615,N_5640);
nand U7158 (N_7158,N_5159,N_5857);
nor U7159 (N_7159,N_5925,N_5551);
nand U7160 (N_7160,N_5616,N_5877);
or U7161 (N_7161,N_5608,N_5303);
xnor U7162 (N_7162,N_4848,N_5640);
nor U7163 (N_7163,N_5138,N_4835);
nand U7164 (N_7164,N_4542,N_5396);
xor U7165 (N_7165,N_5290,N_5438);
and U7166 (N_7166,N_4563,N_4988);
nand U7167 (N_7167,N_5840,N_4640);
nor U7168 (N_7168,N_5629,N_5498);
nor U7169 (N_7169,N_4870,N_4695);
and U7170 (N_7170,N_5399,N_4506);
and U7171 (N_7171,N_4945,N_5237);
xnor U7172 (N_7172,N_5746,N_4942);
xor U7173 (N_7173,N_5872,N_5754);
and U7174 (N_7174,N_5205,N_5372);
or U7175 (N_7175,N_5979,N_4521);
and U7176 (N_7176,N_5385,N_4536);
nor U7177 (N_7177,N_5631,N_4758);
or U7178 (N_7178,N_5503,N_5203);
and U7179 (N_7179,N_4699,N_4804);
nand U7180 (N_7180,N_4910,N_5213);
nor U7181 (N_7181,N_5668,N_4683);
or U7182 (N_7182,N_5176,N_5821);
nor U7183 (N_7183,N_5537,N_5911);
xnor U7184 (N_7184,N_5765,N_5156);
xnor U7185 (N_7185,N_4835,N_4796);
nand U7186 (N_7186,N_4612,N_4505);
xor U7187 (N_7187,N_5719,N_5392);
nor U7188 (N_7188,N_5556,N_5962);
xor U7189 (N_7189,N_5178,N_5372);
and U7190 (N_7190,N_4823,N_5178);
xor U7191 (N_7191,N_4840,N_5188);
nand U7192 (N_7192,N_5793,N_5027);
nor U7193 (N_7193,N_5747,N_5806);
or U7194 (N_7194,N_5838,N_4696);
xnor U7195 (N_7195,N_5171,N_5659);
xnor U7196 (N_7196,N_4572,N_5571);
or U7197 (N_7197,N_4716,N_5450);
nor U7198 (N_7198,N_5583,N_5085);
nor U7199 (N_7199,N_5609,N_5485);
nor U7200 (N_7200,N_5669,N_5966);
nor U7201 (N_7201,N_5519,N_5882);
nand U7202 (N_7202,N_4837,N_5502);
and U7203 (N_7203,N_5313,N_5324);
xor U7204 (N_7204,N_4713,N_4978);
and U7205 (N_7205,N_5802,N_5286);
and U7206 (N_7206,N_4839,N_4877);
and U7207 (N_7207,N_5698,N_4728);
or U7208 (N_7208,N_5998,N_4848);
or U7209 (N_7209,N_5966,N_4831);
or U7210 (N_7210,N_5416,N_5317);
and U7211 (N_7211,N_5730,N_5057);
nor U7212 (N_7212,N_5021,N_5878);
or U7213 (N_7213,N_5158,N_5267);
nand U7214 (N_7214,N_5062,N_5155);
nor U7215 (N_7215,N_5571,N_5291);
and U7216 (N_7216,N_5474,N_5897);
and U7217 (N_7217,N_5904,N_5486);
xor U7218 (N_7218,N_4694,N_5685);
xnor U7219 (N_7219,N_4773,N_5739);
xnor U7220 (N_7220,N_5119,N_5397);
and U7221 (N_7221,N_5670,N_4839);
or U7222 (N_7222,N_5682,N_5073);
xor U7223 (N_7223,N_5303,N_4617);
and U7224 (N_7224,N_5919,N_5867);
or U7225 (N_7225,N_4881,N_5548);
or U7226 (N_7226,N_5457,N_5891);
nand U7227 (N_7227,N_5368,N_5405);
or U7228 (N_7228,N_5747,N_4953);
xor U7229 (N_7229,N_5204,N_5985);
or U7230 (N_7230,N_4571,N_5142);
nand U7231 (N_7231,N_4917,N_5234);
nand U7232 (N_7232,N_5379,N_5145);
and U7233 (N_7233,N_4593,N_4559);
nand U7234 (N_7234,N_5076,N_4722);
nor U7235 (N_7235,N_5730,N_4537);
nand U7236 (N_7236,N_5385,N_5947);
and U7237 (N_7237,N_5616,N_5660);
and U7238 (N_7238,N_5842,N_5951);
nand U7239 (N_7239,N_5853,N_5704);
xnor U7240 (N_7240,N_5051,N_5100);
and U7241 (N_7241,N_5464,N_5183);
nor U7242 (N_7242,N_5435,N_4732);
xnor U7243 (N_7243,N_4752,N_5921);
nor U7244 (N_7244,N_5102,N_5512);
nand U7245 (N_7245,N_5433,N_4619);
nor U7246 (N_7246,N_5008,N_4957);
nor U7247 (N_7247,N_4537,N_4650);
nand U7248 (N_7248,N_4606,N_5765);
nand U7249 (N_7249,N_5602,N_5495);
xor U7250 (N_7250,N_4593,N_5843);
nand U7251 (N_7251,N_5908,N_5269);
or U7252 (N_7252,N_5062,N_4889);
and U7253 (N_7253,N_5598,N_4760);
xnor U7254 (N_7254,N_5056,N_5282);
xor U7255 (N_7255,N_4913,N_5196);
and U7256 (N_7256,N_5909,N_5043);
nor U7257 (N_7257,N_5182,N_4885);
nand U7258 (N_7258,N_4766,N_5921);
nor U7259 (N_7259,N_5561,N_4539);
nand U7260 (N_7260,N_4930,N_5596);
nand U7261 (N_7261,N_5950,N_4524);
or U7262 (N_7262,N_5897,N_5289);
nor U7263 (N_7263,N_5867,N_4893);
nand U7264 (N_7264,N_5969,N_4645);
or U7265 (N_7265,N_5058,N_5258);
nor U7266 (N_7266,N_5710,N_5708);
or U7267 (N_7267,N_5905,N_5276);
or U7268 (N_7268,N_5442,N_5365);
and U7269 (N_7269,N_5868,N_5736);
xnor U7270 (N_7270,N_5398,N_5376);
xor U7271 (N_7271,N_4862,N_5109);
nor U7272 (N_7272,N_4934,N_5497);
nor U7273 (N_7273,N_5867,N_5983);
xor U7274 (N_7274,N_5443,N_5573);
or U7275 (N_7275,N_4550,N_4546);
and U7276 (N_7276,N_5127,N_5295);
and U7277 (N_7277,N_4788,N_5659);
or U7278 (N_7278,N_5566,N_5760);
or U7279 (N_7279,N_4605,N_5428);
nand U7280 (N_7280,N_4642,N_5169);
or U7281 (N_7281,N_5485,N_5085);
and U7282 (N_7282,N_5920,N_5382);
and U7283 (N_7283,N_5677,N_5561);
nor U7284 (N_7284,N_4524,N_5730);
nor U7285 (N_7285,N_5257,N_4800);
nand U7286 (N_7286,N_5092,N_4668);
or U7287 (N_7287,N_4655,N_5868);
and U7288 (N_7288,N_5130,N_4701);
or U7289 (N_7289,N_5603,N_4564);
nor U7290 (N_7290,N_5421,N_5074);
or U7291 (N_7291,N_5499,N_5111);
and U7292 (N_7292,N_4623,N_5578);
nand U7293 (N_7293,N_5986,N_5844);
xor U7294 (N_7294,N_5370,N_5073);
and U7295 (N_7295,N_4897,N_5378);
xor U7296 (N_7296,N_4932,N_5158);
and U7297 (N_7297,N_4841,N_5327);
and U7298 (N_7298,N_5042,N_5197);
nand U7299 (N_7299,N_4513,N_4725);
nand U7300 (N_7300,N_5632,N_4623);
xnor U7301 (N_7301,N_5832,N_5570);
nand U7302 (N_7302,N_5222,N_4661);
and U7303 (N_7303,N_4922,N_4967);
nor U7304 (N_7304,N_5614,N_5978);
nand U7305 (N_7305,N_5232,N_5732);
and U7306 (N_7306,N_5000,N_5146);
or U7307 (N_7307,N_5431,N_4564);
or U7308 (N_7308,N_4818,N_4943);
or U7309 (N_7309,N_5057,N_4754);
nand U7310 (N_7310,N_5052,N_5474);
or U7311 (N_7311,N_5724,N_5860);
nand U7312 (N_7312,N_4559,N_4598);
and U7313 (N_7313,N_4635,N_5321);
nor U7314 (N_7314,N_5130,N_5842);
nand U7315 (N_7315,N_5516,N_4865);
nor U7316 (N_7316,N_5532,N_5083);
or U7317 (N_7317,N_5670,N_5802);
and U7318 (N_7318,N_5789,N_5262);
and U7319 (N_7319,N_4605,N_5563);
nand U7320 (N_7320,N_5423,N_4643);
or U7321 (N_7321,N_5145,N_4914);
nor U7322 (N_7322,N_4940,N_5119);
nor U7323 (N_7323,N_5009,N_4739);
xor U7324 (N_7324,N_4852,N_5485);
nand U7325 (N_7325,N_5126,N_4783);
or U7326 (N_7326,N_5593,N_4853);
and U7327 (N_7327,N_5947,N_5648);
nand U7328 (N_7328,N_5732,N_5617);
or U7329 (N_7329,N_5902,N_4619);
and U7330 (N_7330,N_5914,N_5855);
and U7331 (N_7331,N_5573,N_5807);
and U7332 (N_7332,N_5498,N_4821);
and U7333 (N_7333,N_4728,N_5533);
nand U7334 (N_7334,N_4699,N_5384);
nand U7335 (N_7335,N_5992,N_5276);
nor U7336 (N_7336,N_5077,N_4575);
xor U7337 (N_7337,N_5863,N_4852);
and U7338 (N_7338,N_4771,N_5993);
and U7339 (N_7339,N_5921,N_5670);
and U7340 (N_7340,N_5432,N_5358);
nor U7341 (N_7341,N_5535,N_4684);
xor U7342 (N_7342,N_5552,N_5099);
and U7343 (N_7343,N_5103,N_5390);
or U7344 (N_7344,N_5940,N_5917);
or U7345 (N_7345,N_5021,N_5385);
and U7346 (N_7346,N_4927,N_5467);
xor U7347 (N_7347,N_5037,N_5991);
or U7348 (N_7348,N_4724,N_5712);
xor U7349 (N_7349,N_5074,N_4917);
xor U7350 (N_7350,N_5341,N_5486);
xor U7351 (N_7351,N_4931,N_4544);
or U7352 (N_7352,N_5771,N_4767);
nand U7353 (N_7353,N_5393,N_4625);
xnor U7354 (N_7354,N_5877,N_5788);
nand U7355 (N_7355,N_5837,N_5249);
and U7356 (N_7356,N_4866,N_5542);
nor U7357 (N_7357,N_5853,N_4735);
or U7358 (N_7358,N_5552,N_5667);
xor U7359 (N_7359,N_5312,N_4616);
nor U7360 (N_7360,N_5256,N_5573);
and U7361 (N_7361,N_5691,N_5049);
and U7362 (N_7362,N_5848,N_5092);
and U7363 (N_7363,N_5024,N_5109);
xnor U7364 (N_7364,N_5821,N_5278);
nand U7365 (N_7365,N_5972,N_5273);
xnor U7366 (N_7366,N_5695,N_5885);
xnor U7367 (N_7367,N_5984,N_5828);
or U7368 (N_7368,N_5507,N_4793);
and U7369 (N_7369,N_5831,N_5731);
or U7370 (N_7370,N_4664,N_4842);
nor U7371 (N_7371,N_4692,N_5682);
or U7372 (N_7372,N_4983,N_5252);
or U7373 (N_7373,N_4770,N_5170);
xnor U7374 (N_7374,N_4985,N_5571);
and U7375 (N_7375,N_4734,N_4592);
or U7376 (N_7376,N_5229,N_5324);
or U7377 (N_7377,N_4548,N_4859);
nor U7378 (N_7378,N_5406,N_5887);
nor U7379 (N_7379,N_5198,N_4753);
xor U7380 (N_7380,N_5674,N_5956);
and U7381 (N_7381,N_5247,N_5263);
nand U7382 (N_7382,N_5524,N_4837);
or U7383 (N_7383,N_5082,N_5212);
or U7384 (N_7384,N_4736,N_4877);
xnor U7385 (N_7385,N_5388,N_4780);
nand U7386 (N_7386,N_5471,N_5264);
xor U7387 (N_7387,N_5736,N_5008);
and U7388 (N_7388,N_5825,N_4846);
xor U7389 (N_7389,N_5726,N_5630);
and U7390 (N_7390,N_5404,N_5591);
or U7391 (N_7391,N_5913,N_5706);
xor U7392 (N_7392,N_5914,N_4687);
nor U7393 (N_7393,N_5331,N_4534);
nor U7394 (N_7394,N_5350,N_5816);
xnor U7395 (N_7395,N_5291,N_5603);
xor U7396 (N_7396,N_4768,N_4713);
nand U7397 (N_7397,N_4543,N_5695);
nor U7398 (N_7398,N_5664,N_5820);
and U7399 (N_7399,N_5822,N_5134);
nand U7400 (N_7400,N_5913,N_4832);
and U7401 (N_7401,N_5777,N_5428);
and U7402 (N_7402,N_4512,N_5943);
nor U7403 (N_7403,N_4811,N_4789);
nor U7404 (N_7404,N_5541,N_5654);
xor U7405 (N_7405,N_5852,N_5086);
nand U7406 (N_7406,N_4739,N_5513);
nor U7407 (N_7407,N_5771,N_5438);
and U7408 (N_7408,N_4516,N_5156);
nor U7409 (N_7409,N_5633,N_4892);
and U7410 (N_7410,N_5875,N_5978);
xor U7411 (N_7411,N_5268,N_5563);
and U7412 (N_7412,N_5922,N_5120);
xor U7413 (N_7413,N_5112,N_4748);
and U7414 (N_7414,N_5517,N_4564);
xnor U7415 (N_7415,N_4906,N_5015);
xnor U7416 (N_7416,N_5565,N_5969);
or U7417 (N_7417,N_4873,N_4889);
nand U7418 (N_7418,N_4895,N_5454);
xnor U7419 (N_7419,N_4526,N_5526);
or U7420 (N_7420,N_5125,N_5329);
nand U7421 (N_7421,N_5650,N_5352);
xor U7422 (N_7422,N_4867,N_5902);
xor U7423 (N_7423,N_5569,N_5092);
nand U7424 (N_7424,N_5203,N_5792);
nor U7425 (N_7425,N_5022,N_5064);
and U7426 (N_7426,N_5181,N_5942);
xnor U7427 (N_7427,N_5600,N_5816);
nand U7428 (N_7428,N_5905,N_5472);
or U7429 (N_7429,N_4975,N_5424);
or U7430 (N_7430,N_4877,N_5667);
and U7431 (N_7431,N_5118,N_5115);
and U7432 (N_7432,N_5128,N_4984);
xnor U7433 (N_7433,N_5432,N_5476);
xnor U7434 (N_7434,N_4882,N_5418);
nand U7435 (N_7435,N_5659,N_4576);
nor U7436 (N_7436,N_5999,N_5210);
xnor U7437 (N_7437,N_5486,N_5264);
xor U7438 (N_7438,N_5453,N_5116);
nor U7439 (N_7439,N_5212,N_5582);
or U7440 (N_7440,N_5652,N_5209);
and U7441 (N_7441,N_4612,N_4571);
nand U7442 (N_7442,N_5965,N_4768);
and U7443 (N_7443,N_4751,N_4771);
nand U7444 (N_7444,N_5059,N_5017);
or U7445 (N_7445,N_5275,N_5864);
nand U7446 (N_7446,N_4711,N_5072);
xnor U7447 (N_7447,N_5364,N_5503);
nor U7448 (N_7448,N_5965,N_4730);
xnor U7449 (N_7449,N_5655,N_5736);
nand U7450 (N_7450,N_5277,N_4823);
or U7451 (N_7451,N_4587,N_4945);
nand U7452 (N_7452,N_5872,N_5397);
or U7453 (N_7453,N_5675,N_5755);
nand U7454 (N_7454,N_5395,N_5095);
or U7455 (N_7455,N_5591,N_5260);
xor U7456 (N_7456,N_5092,N_4510);
nor U7457 (N_7457,N_5040,N_5923);
xnor U7458 (N_7458,N_5786,N_5783);
nor U7459 (N_7459,N_5710,N_4601);
nor U7460 (N_7460,N_5658,N_5034);
xnor U7461 (N_7461,N_4842,N_4837);
xor U7462 (N_7462,N_5550,N_5478);
nand U7463 (N_7463,N_5842,N_4709);
or U7464 (N_7464,N_4827,N_4558);
nand U7465 (N_7465,N_4989,N_5548);
xor U7466 (N_7466,N_5987,N_5377);
nor U7467 (N_7467,N_4952,N_5819);
and U7468 (N_7468,N_4697,N_5003);
nand U7469 (N_7469,N_5177,N_5145);
xor U7470 (N_7470,N_4648,N_5611);
and U7471 (N_7471,N_4607,N_5472);
and U7472 (N_7472,N_5342,N_5568);
xor U7473 (N_7473,N_5785,N_5057);
nand U7474 (N_7474,N_5826,N_5064);
nor U7475 (N_7475,N_5607,N_5170);
nand U7476 (N_7476,N_5815,N_4663);
xnor U7477 (N_7477,N_5176,N_4865);
and U7478 (N_7478,N_5261,N_5006);
or U7479 (N_7479,N_4824,N_4725);
nor U7480 (N_7480,N_4914,N_4870);
nand U7481 (N_7481,N_5856,N_4504);
and U7482 (N_7482,N_5425,N_5831);
and U7483 (N_7483,N_4775,N_5227);
xnor U7484 (N_7484,N_5738,N_5350);
nor U7485 (N_7485,N_5158,N_5570);
nor U7486 (N_7486,N_5551,N_5253);
nand U7487 (N_7487,N_5576,N_5338);
nand U7488 (N_7488,N_5428,N_4969);
xnor U7489 (N_7489,N_4787,N_5351);
nand U7490 (N_7490,N_4776,N_5309);
and U7491 (N_7491,N_5445,N_4896);
nand U7492 (N_7492,N_5501,N_5598);
xnor U7493 (N_7493,N_5705,N_5164);
and U7494 (N_7494,N_5787,N_4739);
nor U7495 (N_7495,N_5505,N_5580);
nand U7496 (N_7496,N_5721,N_5645);
and U7497 (N_7497,N_5407,N_5171);
nand U7498 (N_7498,N_5181,N_4908);
nand U7499 (N_7499,N_5855,N_5740);
and U7500 (N_7500,N_6109,N_6348);
and U7501 (N_7501,N_7111,N_6072);
and U7502 (N_7502,N_6576,N_7247);
xor U7503 (N_7503,N_7108,N_6194);
xor U7504 (N_7504,N_6940,N_6448);
nor U7505 (N_7505,N_6938,N_6493);
nand U7506 (N_7506,N_7250,N_6755);
and U7507 (N_7507,N_6705,N_6549);
nor U7508 (N_7508,N_6536,N_6807);
nand U7509 (N_7509,N_7456,N_6308);
nand U7510 (N_7510,N_6313,N_7401);
nand U7511 (N_7511,N_6296,N_6517);
nand U7512 (N_7512,N_7354,N_6502);
xor U7513 (N_7513,N_7136,N_7298);
nor U7514 (N_7514,N_7314,N_7001);
xnor U7515 (N_7515,N_6127,N_7404);
xnor U7516 (N_7516,N_6853,N_6774);
nor U7517 (N_7517,N_7029,N_7253);
nor U7518 (N_7518,N_7408,N_6965);
or U7519 (N_7519,N_7158,N_7074);
and U7520 (N_7520,N_7446,N_7004);
xnor U7521 (N_7521,N_6874,N_6138);
xnor U7522 (N_7522,N_7189,N_6331);
nor U7523 (N_7523,N_7327,N_7166);
nor U7524 (N_7524,N_6144,N_7483);
xor U7525 (N_7525,N_7098,N_6011);
or U7526 (N_7526,N_6663,N_6959);
and U7527 (N_7527,N_6114,N_7142);
xor U7528 (N_7528,N_6652,N_6337);
nor U7529 (N_7529,N_7350,N_7122);
xnor U7530 (N_7530,N_6058,N_6633);
and U7531 (N_7531,N_7195,N_6153);
or U7532 (N_7532,N_6086,N_6364);
and U7533 (N_7533,N_6809,N_7458);
xor U7534 (N_7534,N_6307,N_6232);
or U7535 (N_7535,N_7105,N_6999);
or U7536 (N_7536,N_6883,N_6013);
xnor U7537 (N_7537,N_6944,N_7177);
or U7538 (N_7538,N_7026,N_6150);
and U7539 (N_7539,N_6951,N_7083);
nor U7540 (N_7540,N_6466,N_6597);
nand U7541 (N_7541,N_6410,N_7472);
xnor U7542 (N_7542,N_6686,N_6512);
xor U7543 (N_7543,N_6816,N_6151);
or U7544 (N_7544,N_6146,N_6889);
or U7545 (N_7545,N_6902,N_6192);
and U7546 (N_7546,N_6878,N_6864);
nor U7547 (N_7547,N_7258,N_6321);
xnor U7548 (N_7548,N_7377,N_6112);
xor U7549 (N_7549,N_7190,N_7043);
or U7550 (N_7550,N_6044,N_6798);
or U7551 (N_7551,N_6246,N_6937);
or U7552 (N_7552,N_6697,N_7232);
xnor U7553 (N_7553,N_6757,N_6580);
or U7554 (N_7554,N_6772,N_6462);
xor U7555 (N_7555,N_6645,N_7366);
nor U7556 (N_7556,N_7023,N_7312);
xor U7557 (N_7557,N_7117,N_6780);
or U7558 (N_7558,N_6431,N_6029);
nor U7559 (N_7559,N_6620,N_7019);
and U7560 (N_7560,N_6339,N_6822);
nor U7561 (N_7561,N_6283,N_6602);
nand U7562 (N_7562,N_7181,N_6724);
or U7563 (N_7563,N_6392,N_7073);
or U7564 (N_7564,N_6215,N_6317);
or U7565 (N_7565,N_6273,N_7403);
nor U7566 (N_7566,N_6662,N_7003);
nand U7567 (N_7567,N_7008,N_7447);
nand U7568 (N_7568,N_6183,N_6857);
nor U7569 (N_7569,N_7467,N_7187);
and U7570 (N_7570,N_7249,N_6361);
xor U7571 (N_7571,N_7448,N_6915);
xor U7572 (N_7572,N_6528,N_6116);
xnor U7573 (N_7573,N_6104,N_7347);
or U7574 (N_7574,N_6783,N_6415);
nor U7575 (N_7575,N_6473,N_6209);
xor U7576 (N_7576,N_6142,N_7394);
or U7577 (N_7577,N_6949,N_6129);
nor U7578 (N_7578,N_7342,N_7213);
nor U7579 (N_7579,N_6520,N_6449);
or U7580 (N_7580,N_7490,N_7014);
xor U7581 (N_7581,N_7256,N_6934);
nor U7582 (N_7582,N_6828,N_6794);
xnor U7583 (N_7583,N_6533,N_6530);
or U7584 (N_7584,N_7025,N_6551);
and U7585 (N_7585,N_7222,N_6993);
and U7586 (N_7586,N_6087,N_6992);
or U7587 (N_7587,N_6073,N_7218);
xnor U7588 (N_7588,N_6879,N_6358);
or U7589 (N_7589,N_6529,N_6837);
nand U7590 (N_7590,N_7450,N_6416);
or U7591 (N_7591,N_7307,N_7486);
and U7592 (N_7592,N_7046,N_6744);
and U7593 (N_7593,N_6186,N_6840);
and U7594 (N_7594,N_7297,N_6743);
xnor U7595 (N_7595,N_7086,N_6805);
nand U7596 (N_7596,N_7251,N_7118);
xnor U7597 (N_7597,N_6067,N_6267);
xor U7598 (N_7598,N_7294,N_7234);
and U7599 (N_7599,N_6397,N_6121);
nand U7600 (N_7600,N_6159,N_7487);
xnor U7601 (N_7601,N_7130,N_7388);
nand U7602 (N_7602,N_6801,N_6591);
xor U7603 (N_7603,N_6419,N_6262);
nor U7604 (N_7604,N_7007,N_6737);
xor U7605 (N_7605,N_7402,N_6471);
or U7606 (N_7606,N_6318,N_6522);
and U7607 (N_7607,N_6670,N_6819);
nor U7608 (N_7608,N_7162,N_6479);
nand U7609 (N_7609,N_7042,N_7045);
nor U7610 (N_7610,N_6725,N_6657);
or U7611 (N_7611,N_6438,N_7357);
and U7612 (N_7612,N_6648,N_6120);
nor U7613 (N_7613,N_7422,N_7340);
and U7614 (N_7614,N_7127,N_7259);
nand U7615 (N_7615,N_6792,N_7225);
and U7616 (N_7616,N_7151,N_6031);
xor U7617 (N_7617,N_6342,N_7292);
and U7618 (N_7618,N_7290,N_6735);
nand U7619 (N_7619,N_6835,N_6599);
xor U7620 (N_7620,N_6834,N_6181);
or U7621 (N_7621,N_6156,N_6712);
and U7622 (N_7622,N_7065,N_7468);
or U7623 (N_7623,N_6228,N_6106);
and U7624 (N_7624,N_6688,N_6053);
xnor U7625 (N_7625,N_6326,N_6423);
nor U7626 (N_7626,N_7067,N_6909);
nand U7627 (N_7627,N_6387,N_7305);
xor U7628 (N_7628,N_6564,N_6679);
nand U7629 (N_7629,N_6622,N_6454);
xnor U7630 (N_7630,N_6213,N_6134);
or U7631 (N_7631,N_7433,N_6389);
nor U7632 (N_7632,N_6309,N_7041);
nand U7633 (N_7633,N_7390,N_7245);
nand U7634 (N_7634,N_6420,N_6766);
nand U7635 (N_7635,N_7480,N_6550);
nand U7636 (N_7636,N_6767,N_7119);
and U7637 (N_7637,N_7060,N_6427);
nand U7638 (N_7638,N_6323,N_6340);
xnor U7639 (N_7639,N_7439,N_6226);
or U7640 (N_7640,N_6162,N_6105);
or U7641 (N_7641,N_6941,N_6829);
xnor U7642 (N_7642,N_6861,N_6137);
nor U7643 (N_7643,N_7383,N_6276);
nand U7644 (N_7644,N_6890,N_6925);
or U7645 (N_7645,N_6765,N_7179);
xor U7646 (N_7646,N_6199,N_7457);
xnor U7647 (N_7647,N_7469,N_6238);
or U7648 (N_7648,N_7424,N_6608);
nor U7649 (N_7649,N_6845,N_7360);
or U7650 (N_7650,N_7049,N_6787);
nand U7651 (N_7651,N_6408,N_6220);
xor U7652 (N_7652,N_6268,N_7087);
nor U7653 (N_7653,N_6495,N_7336);
xnor U7654 (N_7654,N_6055,N_6395);
nand U7655 (N_7655,N_6174,N_6758);
nand U7656 (N_7656,N_7077,N_6617);
and U7657 (N_7657,N_7114,N_6019);
and U7658 (N_7658,N_6036,N_7449);
nand U7659 (N_7659,N_6717,N_6923);
nor U7660 (N_7660,N_7129,N_6920);
and U7661 (N_7661,N_7325,N_6190);
xnor U7662 (N_7662,N_6288,N_6726);
or U7663 (N_7663,N_6873,N_6882);
or U7664 (N_7664,N_6930,N_6678);
nor U7665 (N_7665,N_6143,N_6078);
xor U7666 (N_7666,N_7495,N_7202);
and U7667 (N_7667,N_6069,N_7237);
xnor U7668 (N_7668,N_7428,N_6682);
xnor U7669 (N_7669,N_7089,N_7197);
and U7670 (N_7670,N_7092,N_6676);
and U7671 (N_7671,N_6640,N_7126);
xnor U7672 (N_7672,N_6287,N_7462);
xor U7673 (N_7673,N_6931,N_6157);
xor U7674 (N_7674,N_6860,N_6084);
or U7675 (N_7675,N_7267,N_6565);
xor U7676 (N_7676,N_7128,N_6434);
nand U7677 (N_7677,N_6310,N_7319);
or U7678 (N_7678,N_6804,N_6034);
or U7679 (N_7679,N_6642,N_6325);
nor U7680 (N_7680,N_7269,N_6893);
xor U7681 (N_7681,N_6277,N_6535);
nor U7682 (N_7682,N_7382,N_6254);
nor U7683 (N_7683,N_7044,N_7343);
xor U7684 (N_7684,N_7050,N_6612);
nand U7685 (N_7685,N_6002,N_7219);
and U7686 (N_7686,N_6294,N_7134);
nand U7687 (N_7687,N_6411,N_7051);
and U7688 (N_7688,N_6311,N_7315);
xor U7689 (N_7689,N_7465,N_7139);
nor U7690 (N_7690,N_6953,N_6252);
nor U7691 (N_7691,N_6501,N_7263);
xor U7692 (N_7692,N_6338,N_6377);
nor U7693 (N_7693,N_7339,N_6166);
nor U7694 (N_7694,N_6000,N_6082);
and U7695 (N_7695,N_6702,N_6063);
and U7696 (N_7696,N_6349,N_6979);
or U7697 (N_7697,N_6973,N_7420);
or U7698 (N_7698,N_6960,N_6736);
xnor U7699 (N_7699,N_6266,N_6667);
nand U7700 (N_7700,N_6907,N_7123);
xor U7701 (N_7701,N_6230,N_7344);
and U7702 (N_7702,N_7334,N_6083);
and U7703 (N_7703,N_7100,N_6932);
xnor U7704 (N_7704,N_6494,N_6913);
and U7705 (N_7705,N_6750,N_6429);
nor U7706 (N_7706,N_6386,N_6784);
nor U7707 (N_7707,N_6498,N_7082);
and U7708 (N_7708,N_6982,N_7036);
and U7709 (N_7709,N_6871,N_6776);
or U7710 (N_7710,N_6152,N_6527);
and U7711 (N_7711,N_7063,N_6815);
or U7712 (N_7712,N_6826,N_7113);
nand U7713 (N_7713,N_6824,N_7038);
xor U7714 (N_7714,N_6626,N_6426);
nor U7715 (N_7715,N_7188,N_6260);
or U7716 (N_7716,N_6198,N_6988);
and U7717 (N_7717,N_7133,N_6406);
or U7718 (N_7718,N_7176,N_6817);
or U7719 (N_7719,N_6394,N_6546);
xor U7720 (N_7720,N_7296,N_6818);
or U7721 (N_7721,N_7064,N_6672);
and U7722 (N_7722,N_7451,N_6984);
and U7723 (N_7723,N_7248,N_6286);
and U7724 (N_7724,N_6537,N_6996);
and U7725 (N_7725,N_7017,N_7355);
nand U7726 (N_7726,N_6867,N_6135);
xnor U7727 (N_7727,N_7203,N_6762);
and U7728 (N_7728,N_7164,N_7184);
or U7729 (N_7729,N_6500,N_6897);
or U7730 (N_7730,N_6329,N_6716);
xnor U7731 (N_7731,N_7015,N_6887);
and U7732 (N_7732,N_6554,N_6217);
nor U7733 (N_7733,N_6102,N_6666);
or U7734 (N_7734,N_6216,N_6196);
xnor U7735 (N_7735,N_6424,N_7376);
or U7736 (N_7736,N_7473,N_6868);
nand U7737 (N_7737,N_6081,N_6509);
or U7738 (N_7738,N_6435,N_6223);
or U7739 (N_7739,N_6791,N_7024);
and U7740 (N_7740,N_7072,N_6711);
nor U7741 (N_7741,N_6799,N_7069);
xnor U7742 (N_7742,N_6124,N_7299);
and U7743 (N_7743,N_7492,N_6334);
or U7744 (N_7744,N_6698,N_6745);
and U7745 (N_7745,N_7405,N_6171);
nor U7746 (N_7746,N_6202,N_6303);
and U7747 (N_7747,N_7137,N_7321);
or U7748 (N_7748,N_6428,N_6344);
and U7749 (N_7749,N_7317,N_7159);
xor U7750 (N_7750,N_6264,N_7135);
and U7751 (N_7751,N_7191,N_6771);
or U7752 (N_7752,N_6130,N_6467);
or U7753 (N_7753,N_6047,N_7313);
or U7754 (N_7754,N_6110,N_7427);
or U7755 (N_7755,N_6942,N_6123);
nand U7756 (N_7756,N_7095,N_6796);
nand U7757 (N_7757,N_7373,N_6906);
nor U7758 (N_7758,N_6433,N_6604);
or U7759 (N_7759,N_7000,N_6497);
or U7760 (N_7760,N_7423,N_6627);
nand U7761 (N_7761,N_6163,N_6399);
nor U7762 (N_7762,N_6720,N_6594);
nand U7763 (N_7763,N_7417,N_6332);
nor U7764 (N_7764,N_6148,N_6074);
xor U7765 (N_7765,N_6022,N_6628);
and U7766 (N_7766,N_6752,N_6848);
xnor U7767 (N_7767,N_6208,N_6658);
nand U7768 (N_7768,N_6573,N_6369);
nand U7769 (N_7769,N_6919,N_7283);
nand U7770 (N_7770,N_6831,N_7274);
xor U7771 (N_7771,N_7030,N_6506);
nand U7772 (N_7772,N_7198,N_6844);
and U7773 (N_7773,N_6976,N_6849);
xnor U7774 (N_7774,N_6623,N_7378);
nor U7775 (N_7775,N_6224,N_6830);
nand U7776 (N_7776,N_6732,N_6401);
nand U7777 (N_7777,N_6524,N_6231);
nor U7778 (N_7778,N_6068,N_7121);
xor U7779 (N_7779,N_7173,N_7163);
or U7780 (N_7780,N_6299,N_6442);
nand U7781 (N_7781,N_6538,N_6910);
nor U7782 (N_7782,N_6635,N_6929);
xnor U7783 (N_7783,N_6207,N_6723);
and U7784 (N_7784,N_6943,N_7392);
nand U7785 (N_7785,N_6566,N_7395);
and U7786 (N_7786,N_6696,N_6457);
and U7787 (N_7787,N_6885,N_7081);
xor U7788 (N_7788,N_6558,N_7471);
and U7789 (N_7789,N_7300,N_6030);
nand U7790 (N_7790,N_6253,N_6125);
and U7791 (N_7791,N_6681,N_6605);
xnor U7792 (N_7792,N_7115,N_6575);
and U7793 (N_7793,N_6440,N_6490);
nand U7794 (N_7794,N_6584,N_6281);
and U7795 (N_7795,N_6858,N_6094);
and U7796 (N_7796,N_7206,N_6764);
and U7797 (N_7797,N_6997,N_6432);
nand U7798 (N_7798,N_6894,N_6064);
nand U7799 (N_7799,N_6587,N_6598);
and U7800 (N_7800,N_6601,N_6014);
or U7801 (N_7801,N_6655,N_6596);
nor U7802 (N_7802,N_6595,N_6225);
nor U7803 (N_7803,N_7280,N_6091);
nand U7804 (N_7804,N_7367,N_7440);
or U7805 (N_7805,N_7497,N_6324);
or U7806 (N_7806,N_6248,N_6477);
or U7807 (N_7807,N_6131,N_6821);
and U7808 (N_7808,N_7351,N_7287);
and U7809 (N_7809,N_6729,N_6128);
xor U7810 (N_7810,N_6975,N_6214);
nor U7811 (N_7811,N_7398,N_6659);
nand U7812 (N_7812,N_6188,N_6508);
or U7813 (N_7813,N_7443,N_6806);
and U7814 (N_7814,N_6939,N_7271);
nor U7815 (N_7815,N_7146,N_6609);
nor U7816 (N_7816,N_6370,N_6250);
or U7817 (N_7817,N_6483,N_7200);
nor U7818 (N_7818,N_6884,N_6436);
or U7819 (N_7819,N_6354,N_6852);
and U7820 (N_7820,N_6715,N_6734);
or U7821 (N_7821,N_6963,N_6775);
nor U7822 (N_7822,N_6958,N_7037);
nand U7823 (N_7823,N_6024,N_6892);
or U7824 (N_7824,N_6888,N_6185);
or U7825 (N_7825,N_6145,N_6333);
nand U7826 (N_7826,N_6781,N_7012);
and U7827 (N_7827,N_7412,N_6486);
nor U7828 (N_7828,N_6615,N_6341);
or U7829 (N_7829,N_6810,N_7461);
nand U7830 (N_7830,N_6417,N_6272);
or U7831 (N_7831,N_6647,N_7034);
and U7832 (N_7832,N_7236,N_7418);
nor U7833 (N_7833,N_7442,N_6023);
or U7834 (N_7834,N_6895,N_6634);
xor U7835 (N_7835,N_6603,N_6359);
nor U7836 (N_7836,N_7066,N_6704);
or U7837 (N_7837,N_6407,N_6786);
and U7838 (N_7838,N_6139,N_7132);
or U7839 (N_7839,N_6572,N_6859);
nand U7840 (N_7840,N_6691,N_6515);
nor U7841 (N_7841,N_6926,N_6641);
or U7842 (N_7842,N_6970,N_6093);
and U7843 (N_7843,N_6403,N_6579);
or U7844 (N_7844,N_6896,N_7326);
and U7845 (N_7845,N_6210,N_6808);
nor U7846 (N_7846,N_7244,N_7059);
or U7847 (N_7847,N_6684,N_6305);
xor U7848 (N_7848,N_7379,N_6383);
nand U7849 (N_7849,N_7078,N_7363);
nand U7850 (N_7850,N_6050,N_6669);
and U7851 (N_7851,N_7265,N_7454);
and U7852 (N_7852,N_7482,N_7235);
and U7853 (N_7853,N_6274,N_7141);
or U7854 (N_7854,N_6675,N_7459);
nand U7855 (N_7855,N_6221,N_6511);
nor U7856 (N_7856,N_6092,N_6033);
and U7857 (N_7857,N_6051,N_6443);
nand U7858 (N_7858,N_6385,N_6357);
nand U7859 (N_7859,N_6838,N_7138);
or U7860 (N_7860,N_6147,N_7205);
and U7861 (N_7861,N_6170,N_6391);
xnor U7862 (N_7862,N_6079,N_6099);
xor U7863 (N_7863,N_6335,N_7308);
xor U7864 (N_7864,N_6119,N_6983);
and U7865 (N_7865,N_7199,N_7215);
nor U7866 (N_7866,N_6007,N_6785);
nand U7867 (N_7867,N_6870,N_7079);
nand U7868 (N_7868,N_6065,N_6095);
or U7869 (N_7869,N_6090,N_6770);
xnor U7870 (N_7870,N_6905,N_6489);
or U7871 (N_7871,N_6665,N_6468);
and U7872 (N_7872,N_6866,N_7333);
xor U7873 (N_7873,N_7444,N_6330);
or U7874 (N_7874,N_6556,N_7479);
nor U7875 (N_7875,N_6362,N_6351);
and U7876 (N_7876,N_6233,N_6832);
xnor U7877 (N_7877,N_6430,N_6562);
and U7878 (N_7878,N_6204,N_6637);
nor U7879 (N_7879,N_7430,N_7466);
nand U7880 (N_7880,N_6353,N_7431);
and U7881 (N_7881,N_6038,N_7011);
and U7882 (N_7882,N_6010,N_6193);
or U7883 (N_7883,N_7270,N_6492);
or U7884 (N_7884,N_7353,N_6544);
and U7885 (N_7885,N_6160,N_7010);
nor U7886 (N_7886,N_6668,N_6071);
nand U7887 (N_7887,N_6263,N_6977);
nor U7888 (N_7888,N_6460,N_6644);
nor U7889 (N_7889,N_6117,N_6345);
xor U7890 (N_7890,N_6749,N_7053);
and U7891 (N_7891,N_6891,N_6247);
nand U7892 (N_7892,N_6814,N_7346);
xnor U7893 (N_7893,N_6158,N_6021);
xnor U7894 (N_7894,N_6833,N_7494);
or U7895 (N_7895,N_6396,N_6945);
and U7896 (N_7896,N_6740,N_6474);
and U7897 (N_7897,N_6200,N_6446);
xor U7898 (N_7898,N_6346,N_6100);
nand U7899 (N_7899,N_6510,N_6748);
and U7900 (N_7900,N_6012,N_7381);
or U7901 (N_7901,N_7120,N_7436);
xnor U7902 (N_7902,N_7116,N_7056);
or U7903 (N_7903,N_6421,N_6101);
and U7904 (N_7904,N_6096,N_6521);
xor U7905 (N_7905,N_6418,N_6111);
or U7906 (N_7906,N_6936,N_7380);
and U7907 (N_7907,N_6322,N_6673);
and U7908 (N_7908,N_6450,N_6582);
nand U7909 (N_7909,N_6243,N_6412);
or U7910 (N_7910,N_6195,N_7341);
or U7911 (N_7911,N_6719,N_7154);
nand U7912 (N_7912,N_6404,N_7488);
and U7913 (N_7913,N_6149,N_6746);
xor U7914 (N_7914,N_6279,N_6182);
nor U7915 (N_7915,N_6367,N_6865);
xor U7916 (N_7916,N_7039,N_7109);
and U7917 (N_7917,N_6880,N_7358);
or U7918 (N_7918,N_7399,N_6206);
nand U7919 (N_7919,N_7419,N_6178);
nor U7920 (N_7920,N_7107,N_6811);
and U7921 (N_7921,N_6280,N_6855);
nor U7922 (N_7922,N_6827,N_6365);
or U7923 (N_7923,N_6355,N_7145);
nor U7924 (N_7924,N_7091,N_6227);
xnor U7925 (N_7925,N_6189,N_6382);
and U7926 (N_7926,N_6167,N_6126);
and U7927 (N_7927,N_6398,N_6803);
or U7928 (N_7928,N_7273,N_7241);
or U7929 (N_7929,N_6191,N_7435);
and U7930 (N_7930,N_6388,N_6760);
and U7931 (N_7931,N_6018,N_6820);
xnor U7932 (N_7932,N_7359,N_7216);
and U7933 (N_7933,N_6710,N_6306);
nor U7934 (N_7934,N_6847,N_7349);
xor U7935 (N_7935,N_6654,N_7061);
nor U7936 (N_7936,N_6422,N_6585);
or U7937 (N_7937,N_6001,N_6027);
nor U7938 (N_7938,N_6619,N_6289);
nor U7939 (N_7939,N_7304,N_6693);
and U7940 (N_7940,N_6589,N_6249);
or U7941 (N_7941,N_7101,N_6381);
nand U7942 (N_7942,N_7148,N_7210);
xnor U7943 (N_7943,N_7306,N_7481);
and U7944 (N_7944,N_7220,N_7140);
nor U7945 (N_7945,N_7499,N_6759);
xor U7946 (N_7946,N_6995,N_6904);
xor U7947 (N_7947,N_7445,N_7131);
xor U7948 (N_7948,N_6980,N_6779);
xnor U7949 (N_7949,N_6319,N_6451);
nand U7950 (N_7950,N_7028,N_6212);
xor U7951 (N_7951,N_6900,N_7174);
nand U7952 (N_7952,N_7194,N_6463);
nand U7953 (N_7953,N_6561,N_7260);
nor U7954 (N_7954,N_6380,N_7275);
xnor U7955 (N_7955,N_6797,N_6179);
or U7956 (N_7956,N_7452,N_7224);
nor U7957 (N_7957,N_6098,N_7371);
or U7958 (N_7958,N_6085,N_6638);
nor U7959 (N_7959,N_7262,N_6532);
or U7960 (N_7960,N_7476,N_6075);
or U7961 (N_7961,N_7303,N_6708);
xnor U7962 (N_7962,N_7310,N_6015);
nand U7963 (N_7963,N_6251,N_7311);
and U7964 (N_7964,N_6009,N_6269);
nor U7965 (N_7965,N_7183,N_6523);
xor U7966 (N_7966,N_7438,N_7238);
xnor U7967 (N_7967,N_7110,N_6187);
nand U7968 (N_7968,N_6169,N_6695);
nor U7969 (N_7969,N_6742,N_6650);
and U7970 (N_7970,N_7261,N_6846);
nand U7971 (N_7971,N_7209,N_6481);
or U7972 (N_7972,N_7124,N_6020);
nor U7973 (N_7973,N_6025,N_6955);
or U7974 (N_7974,N_6312,N_6842);
xnor U7975 (N_7975,N_7149,N_6707);
xor U7976 (N_7976,N_7147,N_6927);
or U7977 (N_7977,N_6271,N_6136);
nand U7978 (N_7978,N_6548,N_6687);
nand U7979 (N_7979,N_6578,N_6315);
nor U7980 (N_7980,N_6118,N_6470);
xnor U7981 (N_7981,N_6569,N_6588);
and U7982 (N_7982,N_7291,N_6836);
nor U7983 (N_7983,N_6043,N_7040);
or U7984 (N_7984,N_7057,N_7396);
xnor U7985 (N_7985,N_6616,N_7246);
or U7986 (N_7986,N_6229,N_6854);
nand U7987 (N_7987,N_6140,N_7301);
nor U7988 (N_7988,N_6559,N_6950);
nor U7989 (N_7989,N_6076,N_6261);
nor U7990 (N_7990,N_6568,N_7286);
nor U7991 (N_7991,N_6636,N_6851);
xor U7992 (N_7992,N_7293,N_7410);
nor U7993 (N_7993,N_6059,N_6437);
and U7994 (N_7994,N_7182,N_6245);
and U7995 (N_7995,N_7153,N_6244);
or U7996 (N_7996,N_7421,N_7362);
xnor U7997 (N_7997,N_7254,N_6293);
and U7998 (N_7998,N_6184,N_6256);
and U7999 (N_7999,N_7323,N_7088);
or U8000 (N_8000,N_6032,N_6661);
xor U8001 (N_8001,N_6862,N_6475);
xnor U8002 (N_8002,N_6574,N_6553);
nand U8003 (N_8003,N_6685,N_6991);
nand U8004 (N_8004,N_6557,N_6651);
or U8005 (N_8005,N_6378,N_7204);
or U8006 (N_8006,N_6954,N_6802);
nand U8007 (N_8007,N_6618,N_7324);
nor U8008 (N_8008,N_6534,N_7282);
xor U8009 (N_8009,N_7385,N_7397);
xnor U8010 (N_8010,N_6155,N_6747);
nor U8011 (N_8011,N_6692,N_6459);
and U8012 (N_8012,N_6856,N_7309);
nand U8013 (N_8013,N_6543,N_7227);
nand U8014 (N_8014,N_7337,N_6441);
nor U8015 (N_8015,N_6352,N_6778);
and U8016 (N_8016,N_6694,N_6300);
or U8017 (N_8017,N_7242,N_6592);
nor U8018 (N_8018,N_7364,N_6375);
nand U8019 (N_8019,N_6555,N_7231);
or U8020 (N_8020,N_6629,N_6197);
nand U8021 (N_8021,N_6445,N_6593);
or U8022 (N_8022,N_6981,N_7318);
and U8023 (N_8023,N_6291,N_7013);
nor U8024 (N_8024,N_6066,N_6115);
nor U8025 (N_8025,N_7489,N_7085);
nor U8026 (N_8026,N_7230,N_7384);
nand U8027 (N_8027,N_7106,N_6496);
or U8028 (N_8028,N_6518,N_7406);
xor U8029 (N_8029,N_7097,N_6049);
xnor U8030 (N_8030,N_7156,N_7320);
xnor U8031 (N_8031,N_6060,N_6285);
or U8032 (N_8032,N_6630,N_6390);
xor U8033 (N_8033,N_6706,N_7054);
xnor U8034 (N_8034,N_6458,N_6839);
and U8035 (N_8035,N_6132,N_6008);
nor U8036 (N_8036,N_6699,N_6241);
or U8037 (N_8037,N_6173,N_6971);
and U8038 (N_8038,N_6611,N_6606);
nor U8039 (N_8039,N_7062,N_7165);
nor U8040 (N_8040,N_6301,N_6258);
and U8041 (N_8041,N_7170,N_6172);
and U8042 (N_8042,N_6504,N_6823);
and U8043 (N_8043,N_6753,N_6690);
or U8044 (N_8044,N_6639,N_6368);
nand U8045 (N_8045,N_7027,N_7455);
and U8046 (N_8046,N_6653,N_7463);
nand U8047 (N_8047,N_6703,N_6141);
nand U8048 (N_8048,N_7221,N_6994);
nor U8049 (N_8049,N_6077,N_6863);
and U8050 (N_8050,N_7295,N_6218);
nand U8051 (N_8051,N_7322,N_6240);
nor U8052 (N_8052,N_6203,N_6917);
nand U8053 (N_8053,N_7434,N_6107);
or U8054 (N_8054,N_7268,N_7437);
nor U8055 (N_8055,N_6177,N_7103);
and U8056 (N_8056,N_6373,N_6088);
nand U8057 (N_8057,N_6292,N_6825);
xor U8058 (N_8058,N_7208,N_6080);
or U8059 (N_8059,N_6302,N_6769);
nand U8060 (N_8060,N_6540,N_7387);
or U8061 (N_8061,N_6239,N_6164);
xnor U8062 (N_8062,N_6671,N_6877);
or U8063 (N_8063,N_7080,N_6525);
xnor U8064 (N_8064,N_6924,N_7005);
nand U8065 (N_8065,N_7391,N_7018);
nand U8066 (N_8066,N_6026,N_7368);
xnor U8067 (N_8067,N_6800,N_6531);
xnor U8068 (N_8068,N_6374,N_7125);
or U8069 (N_8069,N_6727,N_7161);
nand U8070 (N_8070,N_6986,N_7474);
nor U8071 (N_8071,N_6472,N_7143);
and U8072 (N_8072,N_6414,N_6918);
and U8073 (N_8073,N_6046,N_6133);
and U8074 (N_8074,N_6649,N_7020);
nor U8075 (N_8075,N_6614,N_7369);
nor U8076 (N_8076,N_6176,N_6003);
nor U8077 (N_8077,N_6738,N_7155);
nand U8078 (N_8078,N_7264,N_7196);
and U8079 (N_8079,N_6384,N_6476);
and U8080 (N_8080,N_7460,N_7252);
nor U8081 (N_8081,N_6372,N_6028);
and U8082 (N_8082,N_7257,N_6621);
nand U8083 (N_8083,N_6739,N_7414);
and U8084 (N_8084,N_7058,N_6956);
xnor U8085 (N_8085,N_7052,N_7361);
nand U8086 (N_8086,N_6700,N_6180);
and U8087 (N_8087,N_6974,N_6482);
nand U8088 (N_8088,N_6484,N_6916);
nand U8089 (N_8089,N_7047,N_7084);
nand U8090 (N_8090,N_7160,N_6327);
or U8091 (N_8091,N_6812,N_6777);
nand U8092 (N_8092,N_7285,N_6360);
nor U8093 (N_8093,N_7233,N_7356);
and U8094 (N_8094,N_6061,N_6761);
nor U8095 (N_8095,N_7426,N_7070);
and U8096 (N_8096,N_7207,N_6545);
nor U8097 (N_8097,N_6056,N_6041);
nor U8098 (N_8098,N_7193,N_6656);
xnor U8099 (N_8099,N_6901,N_6488);
nand U8100 (N_8100,N_6947,N_6571);
nand U8101 (N_8101,N_6948,N_7329);
and U8102 (N_8102,N_6040,N_6967);
or U8103 (N_8103,N_6768,N_7400);
xnor U8104 (N_8104,N_6935,N_6843);
nand U8105 (N_8105,N_6205,N_6841);
xnor U8106 (N_8106,N_7002,N_6062);
nand U8107 (N_8107,N_6730,N_7389);
and U8108 (N_8108,N_6567,N_6154);
xor U8109 (N_8109,N_6886,N_7413);
xor U8110 (N_8110,N_6453,N_6017);
or U8111 (N_8111,N_6242,N_7374);
nand U8112 (N_8112,N_6469,N_6298);
or U8113 (N_8113,N_6507,N_6439);
nor U8114 (N_8114,N_6400,N_6563);
and U8115 (N_8115,N_6793,N_7102);
xor U8116 (N_8116,N_6718,N_6570);
nand U8117 (N_8117,N_6499,N_6270);
nand U8118 (N_8118,N_6908,N_7214);
nor U8119 (N_8119,N_7338,N_6456);
and U8120 (N_8120,N_7006,N_7255);
xnor U8121 (N_8121,N_6037,N_7276);
xnor U8122 (N_8122,N_6903,N_6222);
and U8123 (N_8123,N_6985,N_6004);
and U8124 (N_8124,N_6813,N_7068);
nor U8125 (N_8125,N_7345,N_6631);
or U8126 (N_8126,N_7144,N_7175);
and U8127 (N_8127,N_6005,N_6899);
xnor U8128 (N_8128,N_6320,N_7493);
xor U8129 (N_8129,N_7498,N_7093);
nand U8130 (N_8130,N_7112,N_7348);
nor U8131 (N_8131,N_7168,N_6607);
and U8132 (N_8132,N_7228,N_6876);
nor U8133 (N_8133,N_6255,N_6560);
nand U8134 (N_8134,N_7031,N_6175);
xor U8135 (N_8135,N_7186,N_6413);
nand U8136 (N_8136,N_6363,N_6881);
xnor U8137 (N_8137,N_6393,N_6035);
and U8138 (N_8138,N_7243,N_6928);
nand U8139 (N_8139,N_6912,N_6964);
and U8140 (N_8140,N_6505,N_6583);
xor U8141 (N_8141,N_6425,N_6625);
xor U8142 (N_8142,N_6677,N_6600);
nor U8143 (N_8143,N_6048,N_6480);
or U8144 (N_8144,N_6972,N_6683);
xnor U8145 (N_8145,N_7365,N_6850);
and U8146 (N_8146,N_7407,N_6259);
nand U8147 (N_8147,N_7332,N_6284);
and U8148 (N_8148,N_6978,N_6590);
nand U8149 (N_8149,N_7328,N_7009);
xor U8150 (N_8150,N_7432,N_7411);
and U8151 (N_8151,N_6722,N_7032);
and U8152 (N_8152,N_6052,N_7288);
xor U8153 (N_8153,N_7169,N_6356);
and U8154 (N_8154,N_7016,N_6966);
and U8155 (N_8155,N_7352,N_6405);
nand U8156 (N_8156,N_7464,N_6516);
xor U8157 (N_8157,N_7277,N_6444);
nor U8158 (N_8158,N_7441,N_7266);
and U8159 (N_8159,N_6773,N_6968);
and U8160 (N_8160,N_6314,N_6039);
nand U8161 (N_8161,N_6409,N_6042);
or U8162 (N_8162,N_7416,N_6161);
or U8163 (N_8163,N_6343,N_7104);
and U8164 (N_8164,N_6347,N_6613);
and U8165 (N_8165,N_6487,N_6987);
and U8166 (N_8166,N_7171,N_7180);
and U8167 (N_8167,N_6660,N_6016);
nor U8168 (N_8168,N_6045,N_6054);
nor U8169 (N_8169,N_7075,N_6674);
xor U8170 (N_8170,N_6741,N_6552);
nand U8171 (N_8171,N_6234,N_6998);
xor U8172 (N_8172,N_7409,N_7239);
or U8173 (N_8173,N_6872,N_6201);
or U8174 (N_8174,N_6464,N_6278);
nor U8175 (N_8175,N_7485,N_6709);
nor U8176 (N_8176,N_7099,N_6952);
xor U8177 (N_8177,N_6165,N_6455);
or U8178 (N_8178,N_6788,N_6646);
or U8179 (N_8179,N_7331,N_6957);
and U8180 (N_8180,N_7386,N_7055);
and U8181 (N_8181,N_7033,N_7035);
and U8182 (N_8182,N_6782,N_6526);
or U8183 (N_8183,N_7226,N_6282);
and U8184 (N_8184,N_7094,N_6103);
nor U8185 (N_8185,N_6447,N_6006);
xnor U8186 (N_8186,N_6478,N_6946);
and U8187 (N_8187,N_6756,N_6379);
and U8188 (N_8188,N_6057,N_6624);
or U8189 (N_8189,N_7370,N_6689);
xnor U8190 (N_8190,N_6542,N_7415);
or U8191 (N_8191,N_6701,N_6519);
nor U8192 (N_8192,N_6713,N_7212);
and U8193 (N_8193,N_6632,N_6751);
or U8194 (N_8194,N_7201,N_6933);
or U8195 (N_8195,N_6328,N_7278);
nor U8196 (N_8196,N_6721,N_7375);
xor U8197 (N_8197,N_6586,N_6795);
or U8198 (N_8198,N_6581,N_7484);
xor U8199 (N_8199,N_6911,N_7284);
nand U8200 (N_8200,N_6295,N_7470);
nand U8201 (N_8201,N_6990,N_6491);
nor U8202 (N_8202,N_6898,N_7192);
nor U8203 (N_8203,N_6969,N_6168);
or U8204 (N_8204,N_7223,N_7076);
xnor U8205 (N_8205,N_7289,N_7096);
and U8206 (N_8206,N_6366,N_7496);
and U8207 (N_8207,N_6664,N_6113);
xor U8208 (N_8208,N_7157,N_6290);
nand U8209 (N_8209,N_6211,N_7172);
nor U8210 (N_8210,N_6371,N_6731);
nand U8211 (N_8211,N_7477,N_6962);
nor U8212 (N_8212,N_7185,N_7022);
xnor U8213 (N_8213,N_6089,N_6914);
or U8214 (N_8214,N_6921,N_6547);
nand U8215 (N_8215,N_6485,N_7217);
or U8216 (N_8216,N_6236,N_7335);
nand U8217 (N_8217,N_6610,N_7330);
or U8218 (N_8218,N_6763,N_6539);
and U8219 (N_8219,N_6237,N_6070);
and U8220 (N_8220,N_7478,N_7240);
nand U8221 (N_8221,N_6376,N_6336);
or U8222 (N_8222,N_7453,N_6680);
nor U8223 (N_8223,N_6465,N_6257);
xor U8224 (N_8224,N_6922,N_6350);
nor U8225 (N_8225,N_7316,N_7150);
nor U8226 (N_8226,N_7372,N_6265);
and U8227 (N_8227,N_7152,N_6790);
and U8228 (N_8228,N_6961,N_7021);
nor U8229 (N_8229,N_7090,N_6733);
and U8230 (N_8230,N_7167,N_6108);
nand U8231 (N_8231,N_6513,N_7429);
nand U8232 (N_8232,N_6235,N_6503);
xnor U8233 (N_8233,N_6275,N_6643);
or U8234 (N_8234,N_7178,N_6316);
nand U8235 (N_8235,N_7071,N_6989);
or U8236 (N_8236,N_6754,N_6789);
or U8237 (N_8237,N_7491,N_6097);
xnor U8238 (N_8238,N_7279,N_7281);
nor U8239 (N_8239,N_7425,N_7229);
nor U8240 (N_8240,N_6541,N_6461);
or U8241 (N_8241,N_7211,N_6297);
xor U8242 (N_8242,N_6122,N_6577);
nor U8243 (N_8243,N_6304,N_6728);
nand U8244 (N_8244,N_6452,N_7302);
nand U8245 (N_8245,N_6869,N_6402);
nor U8246 (N_8246,N_6219,N_6714);
nor U8247 (N_8247,N_7272,N_7393);
nand U8248 (N_8248,N_6514,N_7475);
and U8249 (N_8249,N_7048,N_6875);
xnor U8250 (N_8250,N_6269,N_6260);
xor U8251 (N_8251,N_7462,N_6363);
and U8252 (N_8252,N_7095,N_6416);
nand U8253 (N_8253,N_6423,N_6466);
nor U8254 (N_8254,N_7148,N_7254);
or U8255 (N_8255,N_6626,N_6483);
nor U8256 (N_8256,N_6023,N_6924);
nand U8257 (N_8257,N_7322,N_7250);
nor U8258 (N_8258,N_7153,N_7379);
nand U8259 (N_8259,N_7075,N_6012);
nor U8260 (N_8260,N_6913,N_6832);
and U8261 (N_8261,N_7210,N_7123);
nand U8262 (N_8262,N_6193,N_6479);
and U8263 (N_8263,N_7390,N_6030);
nor U8264 (N_8264,N_6486,N_6445);
and U8265 (N_8265,N_6373,N_7297);
or U8266 (N_8266,N_6341,N_6153);
xnor U8267 (N_8267,N_6209,N_6461);
nand U8268 (N_8268,N_7085,N_7413);
nor U8269 (N_8269,N_6364,N_7338);
nor U8270 (N_8270,N_6520,N_6206);
or U8271 (N_8271,N_6603,N_6000);
nand U8272 (N_8272,N_6740,N_6917);
nor U8273 (N_8273,N_6934,N_6432);
or U8274 (N_8274,N_7122,N_6973);
nor U8275 (N_8275,N_6095,N_7419);
xnor U8276 (N_8276,N_6672,N_7408);
nand U8277 (N_8277,N_6703,N_6297);
or U8278 (N_8278,N_7325,N_6469);
and U8279 (N_8279,N_6462,N_7196);
and U8280 (N_8280,N_6440,N_6957);
and U8281 (N_8281,N_6985,N_6262);
xor U8282 (N_8282,N_6588,N_6559);
xor U8283 (N_8283,N_6777,N_6804);
or U8284 (N_8284,N_6598,N_6858);
xor U8285 (N_8285,N_7245,N_6171);
xnor U8286 (N_8286,N_7454,N_6895);
and U8287 (N_8287,N_7344,N_6142);
xnor U8288 (N_8288,N_6586,N_7157);
or U8289 (N_8289,N_7165,N_6619);
and U8290 (N_8290,N_6180,N_6388);
and U8291 (N_8291,N_7199,N_6406);
and U8292 (N_8292,N_6217,N_6495);
nand U8293 (N_8293,N_7226,N_6067);
nand U8294 (N_8294,N_6404,N_7005);
or U8295 (N_8295,N_6746,N_6443);
nor U8296 (N_8296,N_6246,N_6136);
or U8297 (N_8297,N_6803,N_7495);
xnor U8298 (N_8298,N_6678,N_6730);
or U8299 (N_8299,N_7132,N_6386);
and U8300 (N_8300,N_6474,N_6944);
or U8301 (N_8301,N_6948,N_6594);
nor U8302 (N_8302,N_6402,N_7471);
nor U8303 (N_8303,N_7120,N_6861);
and U8304 (N_8304,N_6478,N_6824);
and U8305 (N_8305,N_6316,N_6123);
and U8306 (N_8306,N_6772,N_7174);
nor U8307 (N_8307,N_6013,N_6629);
and U8308 (N_8308,N_7127,N_6222);
or U8309 (N_8309,N_6260,N_6592);
and U8310 (N_8310,N_6832,N_6486);
or U8311 (N_8311,N_6164,N_6194);
or U8312 (N_8312,N_6496,N_6548);
nand U8313 (N_8313,N_6529,N_7335);
xnor U8314 (N_8314,N_6762,N_7238);
nand U8315 (N_8315,N_6188,N_6423);
nand U8316 (N_8316,N_6356,N_7442);
nor U8317 (N_8317,N_6762,N_6934);
nand U8318 (N_8318,N_7390,N_6451);
xor U8319 (N_8319,N_6466,N_6168);
xor U8320 (N_8320,N_7171,N_7163);
and U8321 (N_8321,N_6889,N_7032);
nand U8322 (N_8322,N_6930,N_6030);
xor U8323 (N_8323,N_7486,N_6604);
nor U8324 (N_8324,N_6774,N_6905);
nand U8325 (N_8325,N_6976,N_6897);
and U8326 (N_8326,N_7002,N_6558);
nor U8327 (N_8327,N_7326,N_6234);
or U8328 (N_8328,N_6974,N_7353);
or U8329 (N_8329,N_6484,N_6285);
or U8330 (N_8330,N_6066,N_6436);
nand U8331 (N_8331,N_6430,N_7033);
nand U8332 (N_8332,N_7030,N_6814);
nand U8333 (N_8333,N_6183,N_7009);
xor U8334 (N_8334,N_6887,N_6063);
xor U8335 (N_8335,N_6198,N_7003);
nand U8336 (N_8336,N_7095,N_7056);
nor U8337 (N_8337,N_6078,N_6069);
or U8338 (N_8338,N_6392,N_6297);
nor U8339 (N_8339,N_6607,N_6761);
nand U8340 (N_8340,N_7055,N_7118);
nand U8341 (N_8341,N_7474,N_7047);
and U8342 (N_8342,N_7224,N_6666);
xnor U8343 (N_8343,N_6974,N_6087);
nor U8344 (N_8344,N_6518,N_6062);
nor U8345 (N_8345,N_7407,N_7424);
and U8346 (N_8346,N_6047,N_7414);
nand U8347 (N_8347,N_7003,N_6193);
or U8348 (N_8348,N_6427,N_6215);
and U8349 (N_8349,N_7161,N_7160);
nand U8350 (N_8350,N_7148,N_6020);
or U8351 (N_8351,N_7054,N_6894);
nand U8352 (N_8352,N_7272,N_6261);
and U8353 (N_8353,N_6288,N_6908);
nand U8354 (N_8354,N_6453,N_6078);
xor U8355 (N_8355,N_7055,N_7365);
nor U8356 (N_8356,N_7087,N_6979);
xor U8357 (N_8357,N_6894,N_6554);
and U8358 (N_8358,N_6435,N_6065);
and U8359 (N_8359,N_6247,N_6205);
and U8360 (N_8360,N_6312,N_6466);
xnor U8361 (N_8361,N_6585,N_7287);
or U8362 (N_8362,N_6077,N_6476);
and U8363 (N_8363,N_7436,N_7427);
and U8364 (N_8364,N_7243,N_6898);
and U8365 (N_8365,N_6069,N_6318);
nor U8366 (N_8366,N_6559,N_6921);
nor U8367 (N_8367,N_6450,N_7167);
xor U8368 (N_8368,N_6354,N_6067);
nor U8369 (N_8369,N_6973,N_6488);
nor U8370 (N_8370,N_6407,N_7443);
nand U8371 (N_8371,N_6897,N_6664);
or U8372 (N_8372,N_6669,N_6544);
xor U8373 (N_8373,N_7102,N_7125);
xnor U8374 (N_8374,N_6868,N_6360);
nand U8375 (N_8375,N_6767,N_6080);
nor U8376 (N_8376,N_6318,N_6455);
or U8377 (N_8377,N_7072,N_6612);
or U8378 (N_8378,N_7454,N_7133);
or U8379 (N_8379,N_6985,N_6749);
and U8380 (N_8380,N_6845,N_7193);
nor U8381 (N_8381,N_6156,N_7318);
nor U8382 (N_8382,N_7374,N_6972);
nand U8383 (N_8383,N_7090,N_6021);
nor U8384 (N_8384,N_7196,N_7241);
nor U8385 (N_8385,N_6966,N_6495);
nand U8386 (N_8386,N_7143,N_6611);
nor U8387 (N_8387,N_6214,N_7012);
xor U8388 (N_8388,N_7122,N_7270);
nor U8389 (N_8389,N_7012,N_6857);
xor U8390 (N_8390,N_6068,N_7071);
nor U8391 (N_8391,N_7221,N_6600);
or U8392 (N_8392,N_6947,N_7159);
nand U8393 (N_8393,N_7412,N_6634);
or U8394 (N_8394,N_6637,N_7251);
or U8395 (N_8395,N_6050,N_6674);
nand U8396 (N_8396,N_6539,N_6100);
xnor U8397 (N_8397,N_7235,N_7016);
xnor U8398 (N_8398,N_6131,N_6108);
and U8399 (N_8399,N_7116,N_6899);
xnor U8400 (N_8400,N_6360,N_6659);
nor U8401 (N_8401,N_7303,N_6875);
nor U8402 (N_8402,N_6836,N_6564);
xnor U8403 (N_8403,N_7416,N_6493);
xor U8404 (N_8404,N_7139,N_6957);
or U8405 (N_8405,N_7199,N_6348);
or U8406 (N_8406,N_6689,N_6978);
xnor U8407 (N_8407,N_6552,N_7085);
xor U8408 (N_8408,N_6666,N_7304);
xnor U8409 (N_8409,N_6570,N_7176);
xor U8410 (N_8410,N_7314,N_7035);
nor U8411 (N_8411,N_7086,N_6581);
nand U8412 (N_8412,N_7086,N_7175);
xnor U8413 (N_8413,N_6398,N_7225);
or U8414 (N_8414,N_7027,N_6248);
xnor U8415 (N_8415,N_7417,N_6419);
nor U8416 (N_8416,N_6194,N_7318);
xor U8417 (N_8417,N_6746,N_7385);
nor U8418 (N_8418,N_6199,N_6246);
nor U8419 (N_8419,N_7315,N_6117);
xnor U8420 (N_8420,N_6460,N_6361);
nor U8421 (N_8421,N_6232,N_7216);
nand U8422 (N_8422,N_6332,N_6221);
nor U8423 (N_8423,N_7183,N_7247);
nand U8424 (N_8424,N_7133,N_6822);
and U8425 (N_8425,N_6072,N_6805);
xor U8426 (N_8426,N_6802,N_6846);
nand U8427 (N_8427,N_6588,N_6978);
xor U8428 (N_8428,N_7226,N_7369);
and U8429 (N_8429,N_6309,N_7187);
xnor U8430 (N_8430,N_7461,N_6996);
nor U8431 (N_8431,N_6139,N_7366);
xor U8432 (N_8432,N_7429,N_7236);
nor U8433 (N_8433,N_7460,N_6369);
nand U8434 (N_8434,N_6716,N_7433);
and U8435 (N_8435,N_7398,N_6309);
nor U8436 (N_8436,N_6735,N_6449);
and U8437 (N_8437,N_7122,N_6077);
or U8438 (N_8438,N_7391,N_6052);
and U8439 (N_8439,N_6706,N_7184);
and U8440 (N_8440,N_6278,N_6080);
and U8441 (N_8441,N_7471,N_7137);
and U8442 (N_8442,N_7474,N_6685);
xor U8443 (N_8443,N_7377,N_6041);
or U8444 (N_8444,N_6665,N_6884);
or U8445 (N_8445,N_6330,N_7431);
xnor U8446 (N_8446,N_6686,N_7367);
xnor U8447 (N_8447,N_6303,N_7254);
nor U8448 (N_8448,N_7021,N_7383);
xnor U8449 (N_8449,N_7007,N_6094);
nand U8450 (N_8450,N_6895,N_7261);
and U8451 (N_8451,N_6206,N_7011);
xor U8452 (N_8452,N_6012,N_7004);
nand U8453 (N_8453,N_6380,N_6318);
and U8454 (N_8454,N_6719,N_6615);
nand U8455 (N_8455,N_6277,N_6001);
nand U8456 (N_8456,N_7123,N_6601);
xor U8457 (N_8457,N_6168,N_6543);
xor U8458 (N_8458,N_6030,N_6103);
or U8459 (N_8459,N_6459,N_7363);
nor U8460 (N_8460,N_6103,N_6469);
nor U8461 (N_8461,N_7090,N_6731);
and U8462 (N_8462,N_6474,N_6637);
nor U8463 (N_8463,N_7190,N_7399);
or U8464 (N_8464,N_7467,N_6530);
nor U8465 (N_8465,N_6169,N_6957);
nor U8466 (N_8466,N_6186,N_7460);
xnor U8467 (N_8467,N_6482,N_7204);
or U8468 (N_8468,N_7172,N_7056);
nor U8469 (N_8469,N_6962,N_6515);
and U8470 (N_8470,N_6551,N_7327);
or U8471 (N_8471,N_7016,N_7403);
or U8472 (N_8472,N_7382,N_6523);
xnor U8473 (N_8473,N_6475,N_6818);
or U8474 (N_8474,N_6523,N_6215);
nand U8475 (N_8475,N_6070,N_6728);
nor U8476 (N_8476,N_6967,N_7024);
nand U8477 (N_8477,N_6721,N_6469);
or U8478 (N_8478,N_6829,N_7206);
or U8479 (N_8479,N_6309,N_6514);
xnor U8480 (N_8480,N_6949,N_7216);
or U8481 (N_8481,N_6978,N_6057);
nand U8482 (N_8482,N_6629,N_6399);
nand U8483 (N_8483,N_6695,N_6627);
nand U8484 (N_8484,N_6124,N_7461);
and U8485 (N_8485,N_7030,N_7493);
xnor U8486 (N_8486,N_6757,N_7163);
xor U8487 (N_8487,N_7363,N_7382);
or U8488 (N_8488,N_6088,N_7335);
xor U8489 (N_8489,N_6625,N_7240);
or U8490 (N_8490,N_6442,N_6274);
and U8491 (N_8491,N_6374,N_6033);
and U8492 (N_8492,N_7125,N_7184);
or U8493 (N_8493,N_6820,N_6720);
and U8494 (N_8494,N_6188,N_6999);
nor U8495 (N_8495,N_6226,N_6872);
xnor U8496 (N_8496,N_6906,N_6506);
xnor U8497 (N_8497,N_7180,N_6125);
nand U8498 (N_8498,N_7353,N_6451);
nand U8499 (N_8499,N_6368,N_7452);
nand U8500 (N_8500,N_6092,N_6142);
and U8501 (N_8501,N_6964,N_7457);
nand U8502 (N_8502,N_6196,N_6210);
xnor U8503 (N_8503,N_6180,N_6809);
or U8504 (N_8504,N_6052,N_6775);
and U8505 (N_8505,N_6536,N_7236);
nand U8506 (N_8506,N_6157,N_6118);
and U8507 (N_8507,N_6358,N_6632);
nor U8508 (N_8508,N_7348,N_7335);
xnor U8509 (N_8509,N_7348,N_6777);
nor U8510 (N_8510,N_6756,N_6853);
nor U8511 (N_8511,N_7319,N_6093);
xnor U8512 (N_8512,N_6085,N_6886);
xor U8513 (N_8513,N_7312,N_6379);
xnor U8514 (N_8514,N_7295,N_6357);
nor U8515 (N_8515,N_7223,N_6199);
xor U8516 (N_8516,N_6746,N_7042);
and U8517 (N_8517,N_6062,N_7388);
nor U8518 (N_8518,N_6613,N_7369);
or U8519 (N_8519,N_7316,N_6689);
and U8520 (N_8520,N_6086,N_6554);
xor U8521 (N_8521,N_6741,N_7334);
nand U8522 (N_8522,N_6028,N_6076);
and U8523 (N_8523,N_6558,N_6309);
or U8524 (N_8524,N_6465,N_7295);
or U8525 (N_8525,N_6303,N_6338);
and U8526 (N_8526,N_6634,N_6842);
and U8527 (N_8527,N_6950,N_6812);
nor U8528 (N_8528,N_7362,N_7320);
or U8529 (N_8529,N_6617,N_7302);
or U8530 (N_8530,N_7300,N_7299);
xor U8531 (N_8531,N_6468,N_6421);
nor U8532 (N_8532,N_6726,N_7227);
xnor U8533 (N_8533,N_6052,N_6531);
and U8534 (N_8534,N_7447,N_7201);
and U8535 (N_8535,N_7026,N_7330);
nor U8536 (N_8536,N_6797,N_6587);
nor U8537 (N_8537,N_6667,N_7238);
xnor U8538 (N_8538,N_6926,N_7297);
and U8539 (N_8539,N_6552,N_6362);
and U8540 (N_8540,N_6287,N_7333);
nand U8541 (N_8541,N_7235,N_6480);
nand U8542 (N_8542,N_7469,N_6208);
nor U8543 (N_8543,N_7363,N_6030);
nand U8544 (N_8544,N_6816,N_6971);
xor U8545 (N_8545,N_6499,N_7473);
nand U8546 (N_8546,N_7188,N_6638);
or U8547 (N_8547,N_6444,N_6178);
xor U8548 (N_8548,N_7333,N_7109);
nand U8549 (N_8549,N_6930,N_7174);
and U8550 (N_8550,N_6109,N_7136);
and U8551 (N_8551,N_7045,N_7414);
and U8552 (N_8552,N_6685,N_6781);
xor U8553 (N_8553,N_6185,N_7231);
nor U8554 (N_8554,N_7217,N_7143);
nor U8555 (N_8555,N_6348,N_6266);
and U8556 (N_8556,N_6309,N_6587);
nand U8557 (N_8557,N_6835,N_7005);
nor U8558 (N_8558,N_6933,N_6860);
nand U8559 (N_8559,N_6719,N_6789);
nor U8560 (N_8560,N_7301,N_6664);
or U8561 (N_8561,N_6662,N_6534);
or U8562 (N_8562,N_7138,N_6082);
nor U8563 (N_8563,N_6356,N_6884);
nor U8564 (N_8564,N_6194,N_7176);
nand U8565 (N_8565,N_6515,N_6154);
nand U8566 (N_8566,N_6470,N_6012);
or U8567 (N_8567,N_6561,N_6226);
and U8568 (N_8568,N_6431,N_6756);
nor U8569 (N_8569,N_7446,N_6194);
or U8570 (N_8570,N_7434,N_6945);
nor U8571 (N_8571,N_6288,N_6684);
nor U8572 (N_8572,N_7110,N_6758);
xor U8573 (N_8573,N_6497,N_7099);
xor U8574 (N_8574,N_6723,N_6466);
or U8575 (N_8575,N_7262,N_6580);
xor U8576 (N_8576,N_7194,N_6487);
and U8577 (N_8577,N_7338,N_6078);
nand U8578 (N_8578,N_7087,N_7295);
xor U8579 (N_8579,N_6856,N_6027);
or U8580 (N_8580,N_6283,N_6214);
and U8581 (N_8581,N_6793,N_6744);
xnor U8582 (N_8582,N_6358,N_7383);
nor U8583 (N_8583,N_6360,N_7247);
xnor U8584 (N_8584,N_6850,N_7421);
and U8585 (N_8585,N_6134,N_6016);
xnor U8586 (N_8586,N_6906,N_6792);
or U8587 (N_8587,N_6911,N_6818);
nand U8588 (N_8588,N_6657,N_6465);
and U8589 (N_8589,N_6556,N_6587);
and U8590 (N_8590,N_6290,N_7176);
and U8591 (N_8591,N_6716,N_6938);
nand U8592 (N_8592,N_6581,N_7037);
xor U8593 (N_8593,N_7228,N_6040);
nand U8594 (N_8594,N_6899,N_6272);
or U8595 (N_8595,N_6715,N_6356);
and U8596 (N_8596,N_7345,N_6794);
or U8597 (N_8597,N_6858,N_7232);
xor U8598 (N_8598,N_6778,N_6781);
or U8599 (N_8599,N_6309,N_7100);
nand U8600 (N_8600,N_6268,N_7485);
xnor U8601 (N_8601,N_7470,N_7278);
or U8602 (N_8602,N_7471,N_6804);
xnor U8603 (N_8603,N_6723,N_6147);
xor U8604 (N_8604,N_6455,N_7425);
and U8605 (N_8605,N_6621,N_6573);
xnor U8606 (N_8606,N_6772,N_6500);
xor U8607 (N_8607,N_7199,N_7127);
nand U8608 (N_8608,N_7296,N_6242);
and U8609 (N_8609,N_6040,N_6845);
xor U8610 (N_8610,N_6452,N_7078);
nand U8611 (N_8611,N_7198,N_6037);
nand U8612 (N_8612,N_6935,N_6933);
nor U8613 (N_8613,N_7320,N_7397);
nor U8614 (N_8614,N_6314,N_6497);
and U8615 (N_8615,N_7469,N_6956);
nand U8616 (N_8616,N_6946,N_6553);
nand U8617 (N_8617,N_6386,N_6244);
or U8618 (N_8618,N_6265,N_7448);
xor U8619 (N_8619,N_6386,N_6804);
or U8620 (N_8620,N_6088,N_6089);
xor U8621 (N_8621,N_6259,N_7432);
xnor U8622 (N_8622,N_7219,N_6299);
xor U8623 (N_8623,N_6991,N_6832);
nor U8624 (N_8624,N_7307,N_7055);
xor U8625 (N_8625,N_6083,N_6871);
nand U8626 (N_8626,N_6269,N_7270);
and U8627 (N_8627,N_6104,N_7419);
or U8628 (N_8628,N_6055,N_6385);
nor U8629 (N_8629,N_7368,N_7026);
and U8630 (N_8630,N_7404,N_7487);
xnor U8631 (N_8631,N_6787,N_6183);
nor U8632 (N_8632,N_6135,N_6031);
or U8633 (N_8633,N_6316,N_6086);
and U8634 (N_8634,N_6380,N_7181);
and U8635 (N_8635,N_7305,N_6071);
nor U8636 (N_8636,N_6366,N_6793);
nor U8637 (N_8637,N_6695,N_6711);
xor U8638 (N_8638,N_7413,N_6767);
xnor U8639 (N_8639,N_7066,N_6694);
nor U8640 (N_8640,N_6661,N_7247);
xor U8641 (N_8641,N_6332,N_6409);
or U8642 (N_8642,N_6604,N_7215);
nor U8643 (N_8643,N_7440,N_6254);
xnor U8644 (N_8644,N_7468,N_6081);
and U8645 (N_8645,N_7283,N_6670);
and U8646 (N_8646,N_6761,N_6595);
or U8647 (N_8647,N_6514,N_6155);
or U8648 (N_8648,N_6115,N_6449);
or U8649 (N_8649,N_7227,N_6546);
and U8650 (N_8650,N_6795,N_6548);
and U8651 (N_8651,N_6882,N_6092);
nand U8652 (N_8652,N_7121,N_6667);
xor U8653 (N_8653,N_7479,N_6569);
or U8654 (N_8654,N_6404,N_6610);
xnor U8655 (N_8655,N_6398,N_7288);
and U8656 (N_8656,N_7453,N_6215);
nor U8657 (N_8657,N_6113,N_6534);
nor U8658 (N_8658,N_6350,N_7009);
nor U8659 (N_8659,N_7390,N_6771);
and U8660 (N_8660,N_6946,N_6423);
xnor U8661 (N_8661,N_7349,N_7247);
and U8662 (N_8662,N_7206,N_7337);
nor U8663 (N_8663,N_6230,N_7159);
nand U8664 (N_8664,N_7413,N_6223);
and U8665 (N_8665,N_6534,N_7357);
nand U8666 (N_8666,N_7130,N_7381);
xnor U8667 (N_8667,N_6754,N_6882);
nor U8668 (N_8668,N_7042,N_7122);
nand U8669 (N_8669,N_6204,N_6769);
xor U8670 (N_8670,N_6277,N_6655);
xnor U8671 (N_8671,N_7449,N_6670);
nand U8672 (N_8672,N_7345,N_7472);
and U8673 (N_8673,N_6105,N_6428);
xor U8674 (N_8674,N_6542,N_6487);
xnor U8675 (N_8675,N_6148,N_6066);
or U8676 (N_8676,N_7227,N_6265);
and U8677 (N_8677,N_6334,N_6952);
nor U8678 (N_8678,N_7020,N_6995);
nor U8679 (N_8679,N_6654,N_7249);
nor U8680 (N_8680,N_7388,N_7415);
nand U8681 (N_8681,N_7406,N_6328);
nor U8682 (N_8682,N_7146,N_6527);
nor U8683 (N_8683,N_6830,N_7497);
nand U8684 (N_8684,N_7169,N_6749);
nand U8685 (N_8685,N_7311,N_6278);
xor U8686 (N_8686,N_7108,N_6482);
or U8687 (N_8687,N_7391,N_7285);
xor U8688 (N_8688,N_7170,N_6042);
and U8689 (N_8689,N_6477,N_6181);
or U8690 (N_8690,N_6867,N_6326);
and U8691 (N_8691,N_6331,N_6514);
xnor U8692 (N_8692,N_6359,N_6694);
nor U8693 (N_8693,N_6653,N_6071);
and U8694 (N_8694,N_6587,N_6755);
and U8695 (N_8695,N_7185,N_6511);
nor U8696 (N_8696,N_7491,N_6466);
nor U8697 (N_8697,N_6448,N_6168);
nand U8698 (N_8698,N_6672,N_6361);
or U8699 (N_8699,N_7097,N_7291);
nand U8700 (N_8700,N_6933,N_7481);
nand U8701 (N_8701,N_6398,N_6711);
or U8702 (N_8702,N_7167,N_6502);
or U8703 (N_8703,N_7339,N_7095);
and U8704 (N_8704,N_6940,N_6159);
xor U8705 (N_8705,N_7200,N_6896);
xor U8706 (N_8706,N_6663,N_6738);
and U8707 (N_8707,N_6115,N_6546);
xnor U8708 (N_8708,N_7096,N_6063);
nor U8709 (N_8709,N_6179,N_6607);
nand U8710 (N_8710,N_7147,N_6223);
nor U8711 (N_8711,N_6801,N_6300);
nor U8712 (N_8712,N_6337,N_6474);
nor U8713 (N_8713,N_6602,N_7003);
nand U8714 (N_8714,N_6640,N_6000);
and U8715 (N_8715,N_6738,N_6761);
nor U8716 (N_8716,N_7241,N_7242);
nand U8717 (N_8717,N_7056,N_6758);
nand U8718 (N_8718,N_6831,N_6929);
xnor U8719 (N_8719,N_6306,N_6045);
xor U8720 (N_8720,N_6874,N_6249);
xnor U8721 (N_8721,N_6398,N_6515);
and U8722 (N_8722,N_6688,N_7397);
nor U8723 (N_8723,N_6488,N_6401);
or U8724 (N_8724,N_6362,N_7174);
nand U8725 (N_8725,N_6916,N_7275);
nor U8726 (N_8726,N_6358,N_6693);
nand U8727 (N_8727,N_6488,N_6036);
xor U8728 (N_8728,N_7131,N_6104);
nor U8729 (N_8729,N_6864,N_6693);
nor U8730 (N_8730,N_6121,N_6665);
or U8731 (N_8731,N_6146,N_6223);
and U8732 (N_8732,N_6497,N_6175);
xor U8733 (N_8733,N_7185,N_6351);
nand U8734 (N_8734,N_6360,N_6738);
or U8735 (N_8735,N_6995,N_7310);
or U8736 (N_8736,N_7439,N_7378);
nand U8737 (N_8737,N_6892,N_6808);
nor U8738 (N_8738,N_6757,N_7391);
or U8739 (N_8739,N_6138,N_6790);
or U8740 (N_8740,N_6607,N_7201);
xor U8741 (N_8741,N_7243,N_6536);
and U8742 (N_8742,N_6007,N_7180);
or U8743 (N_8743,N_6005,N_7105);
nor U8744 (N_8744,N_6362,N_6835);
and U8745 (N_8745,N_6431,N_6167);
or U8746 (N_8746,N_6569,N_6370);
or U8747 (N_8747,N_6483,N_6233);
xor U8748 (N_8748,N_7103,N_7490);
nand U8749 (N_8749,N_6533,N_7224);
nor U8750 (N_8750,N_6299,N_6175);
nand U8751 (N_8751,N_7298,N_6009);
nor U8752 (N_8752,N_7371,N_6076);
or U8753 (N_8753,N_6102,N_6916);
xnor U8754 (N_8754,N_6852,N_7161);
nand U8755 (N_8755,N_6546,N_6474);
xor U8756 (N_8756,N_6922,N_6686);
and U8757 (N_8757,N_7213,N_6238);
nor U8758 (N_8758,N_7468,N_6142);
or U8759 (N_8759,N_6962,N_7208);
nor U8760 (N_8760,N_7306,N_6432);
xnor U8761 (N_8761,N_6632,N_6912);
nand U8762 (N_8762,N_7430,N_6174);
and U8763 (N_8763,N_7374,N_6310);
xnor U8764 (N_8764,N_6835,N_7335);
nor U8765 (N_8765,N_6361,N_6445);
nand U8766 (N_8766,N_6111,N_7382);
or U8767 (N_8767,N_6395,N_6767);
xnor U8768 (N_8768,N_6753,N_6360);
nand U8769 (N_8769,N_6082,N_6677);
or U8770 (N_8770,N_6313,N_6503);
xnor U8771 (N_8771,N_7112,N_6861);
xor U8772 (N_8772,N_6250,N_6389);
nand U8773 (N_8773,N_6199,N_6229);
and U8774 (N_8774,N_7242,N_7223);
nand U8775 (N_8775,N_7479,N_7069);
or U8776 (N_8776,N_7433,N_6841);
nand U8777 (N_8777,N_6105,N_7207);
xnor U8778 (N_8778,N_7072,N_7011);
nor U8779 (N_8779,N_6410,N_6531);
xnor U8780 (N_8780,N_6914,N_7360);
or U8781 (N_8781,N_6655,N_6116);
xnor U8782 (N_8782,N_6096,N_6783);
xor U8783 (N_8783,N_7342,N_6238);
xor U8784 (N_8784,N_6053,N_6238);
xor U8785 (N_8785,N_6371,N_6924);
xnor U8786 (N_8786,N_6612,N_6149);
xor U8787 (N_8787,N_6001,N_6945);
or U8788 (N_8788,N_6614,N_6184);
nand U8789 (N_8789,N_6654,N_6355);
xor U8790 (N_8790,N_6747,N_6900);
and U8791 (N_8791,N_7023,N_6635);
or U8792 (N_8792,N_6325,N_7173);
nand U8793 (N_8793,N_7388,N_6728);
xnor U8794 (N_8794,N_6676,N_7159);
and U8795 (N_8795,N_6969,N_7306);
or U8796 (N_8796,N_7329,N_6833);
xnor U8797 (N_8797,N_7350,N_6443);
nor U8798 (N_8798,N_7003,N_6718);
nand U8799 (N_8799,N_6474,N_7339);
or U8800 (N_8800,N_6220,N_6802);
or U8801 (N_8801,N_7221,N_7283);
nor U8802 (N_8802,N_7078,N_6592);
or U8803 (N_8803,N_6380,N_6005);
nand U8804 (N_8804,N_7090,N_6130);
nand U8805 (N_8805,N_6037,N_7277);
nor U8806 (N_8806,N_6509,N_6862);
nor U8807 (N_8807,N_7322,N_6836);
and U8808 (N_8808,N_6979,N_7056);
xnor U8809 (N_8809,N_7016,N_6372);
nor U8810 (N_8810,N_6787,N_6619);
nor U8811 (N_8811,N_6937,N_6173);
or U8812 (N_8812,N_7216,N_6394);
or U8813 (N_8813,N_6700,N_6048);
or U8814 (N_8814,N_6127,N_6568);
nand U8815 (N_8815,N_7121,N_6136);
and U8816 (N_8816,N_7011,N_6210);
nor U8817 (N_8817,N_6174,N_7209);
xnor U8818 (N_8818,N_6517,N_7237);
nand U8819 (N_8819,N_6127,N_6242);
or U8820 (N_8820,N_7087,N_7342);
nor U8821 (N_8821,N_6511,N_6478);
xor U8822 (N_8822,N_6037,N_7336);
nand U8823 (N_8823,N_6295,N_6119);
xnor U8824 (N_8824,N_7230,N_6944);
and U8825 (N_8825,N_7444,N_6097);
or U8826 (N_8826,N_7180,N_7395);
nand U8827 (N_8827,N_7438,N_7295);
nand U8828 (N_8828,N_7011,N_6763);
xor U8829 (N_8829,N_6759,N_7059);
xnor U8830 (N_8830,N_6269,N_7413);
or U8831 (N_8831,N_7363,N_6542);
xor U8832 (N_8832,N_7334,N_6690);
and U8833 (N_8833,N_7401,N_7368);
and U8834 (N_8834,N_7177,N_6070);
nor U8835 (N_8835,N_6151,N_7223);
nand U8836 (N_8836,N_7324,N_6795);
xor U8837 (N_8837,N_7496,N_6035);
nor U8838 (N_8838,N_6506,N_6837);
or U8839 (N_8839,N_7174,N_7391);
xnor U8840 (N_8840,N_7022,N_6883);
or U8841 (N_8841,N_7116,N_7179);
xnor U8842 (N_8842,N_6765,N_6503);
nor U8843 (N_8843,N_6204,N_6139);
nand U8844 (N_8844,N_7444,N_6478);
xor U8845 (N_8845,N_7157,N_6165);
nand U8846 (N_8846,N_6095,N_6774);
xor U8847 (N_8847,N_6009,N_7051);
or U8848 (N_8848,N_6976,N_6800);
and U8849 (N_8849,N_7172,N_7367);
nor U8850 (N_8850,N_6897,N_7112);
xnor U8851 (N_8851,N_6512,N_6209);
xnor U8852 (N_8852,N_6287,N_6929);
nor U8853 (N_8853,N_7440,N_6290);
and U8854 (N_8854,N_6895,N_6246);
xor U8855 (N_8855,N_6458,N_6996);
or U8856 (N_8856,N_6193,N_6509);
nand U8857 (N_8857,N_6162,N_6952);
nor U8858 (N_8858,N_7371,N_6411);
and U8859 (N_8859,N_6880,N_6274);
nand U8860 (N_8860,N_6305,N_7260);
nor U8861 (N_8861,N_6893,N_6231);
or U8862 (N_8862,N_6480,N_6830);
nor U8863 (N_8863,N_6665,N_6868);
nand U8864 (N_8864,N_6247,N_6501);
nand U8865 (N_8865,N_7470,N_6223);
xnor U8866 (N_8866,N_6318,N_6641);
xnor U8867 (N_8867,N_7364,N_6942);
nor U8868 (N_8868,N_7296,N_6428);
or U8869 (N_8869,N_7054,N_6680);
nor U8870 (N_8870,N_6848,N_6073);
or U8871 (N_8871,N_6763,N_6729);
xor U8872 (N_8872,N_7270,N_7197);
nor U8873 (N_8873,N_6317,N_7316);
and U8874 (N_8874,N_6183,N_6561);
xor U8875 (N_8875,N_6153,N_6987);
or U8876 (N_8876,N_6641,N_6291);
nand U8877 (N_8877,N_7025,N_6491);
nand U8878 (N_8878,N_6101,N_6927);
nor U8879 (N_8879,N_6335,N_6551);
nand U8880 (N_8880,N_6682,N_7075);
xnor U8881 (N_8881,N_6400,N_7179);
xor U8882 (N_8882,N_6682,N_6794);
nor U8883 (N_8883,N_6582,N_7403);
or U8884 (N_8884,N_6555,N_7116);
and U8885 (N_8885,N_6075,N_6965);
nor U8886 (N_8886,N_6324,N_7408);
nor U8887 (N_8887,N_6761,N_7364);
or U8888 (N_8888,N_7427,N_7224);
nor U8889 (N_8889,N_6889,N_7395);
and U8890 (N_8890,N_6333,N_6517);
xnor U8891 (N_8891,N_6807,N_7300);
xnor U8892 (N_8892,N_6394,N_6730);
and U8893 (N_8893,N_6597,N_6298);
xor U8894 (N_8894,N_7434,N_7417);
nand U8895 (N_8895,N_6866,N_7008);
xor U8896 (N_8896,N_7376,N_6293);
nand U8897 (N_8897,N_7323,N_6921);
or U8898 (N_8898,N_6634,N_6287);
nor U8899 (N_8899,N_6056,N_6449);
nand U8900 (N_8900,N_6431,N_6020);
nor U8901 (N_8901,N_6621,N_6480);
and U8902 (N_8902,N_6230,N_6716);
or U8903 (N_8903,N_6913,N_6352);
xnor U8904 (N_8904,N_7228,N_6092);
or U8905 (N_8905,N_6067,N_7468);
nand U8906 (N_8906,N_6824,N_6117);
xor U8907 (N_8907,N_6569,N_6950);
xnor U8908 (N_8908,N_6278,N_7231);
nor U8909 (N_8909,N_6781,N_6206);
nand U8910 (N_8910,N_7028,N_7099);
nor U8911 (N_8911,N_6293,N_6748);
or U8912 (N_8912,N_6295,N_6331);
nand U8913 (N_8913,N_7317,N_7460);
and U8914 (N_8914,N_6533,N_7358);
nor U8915 (N_8915,N_7249,N_7452);
xnor U8916 (N_8916,N_6474,N_6517);
or U8917 (N_8917,N_6989,N_7037);
and U8918 (N_8918,N_7060,N_6578);
nor U8919 (N_8919,N_7399,N_6060);
and U8920 (N_8920,N_6132,N_6449);
xor U8921 (N_8921,N_6671,N_6464);
nor U8922 (N_8922,N_7314,N_6417);
and U8923 (N_8923,N_7145,N_6748);
nand U8924 (N_8924,N_7382,N_7022);
xor U8925 (N_8925,N_6735,N_6607);
nand U8926 (N_8926,N_6085,N_6612);
nand U8927 (N_8927,N_7306,N_6531);
nor U8928 (N_8928,N_7339,N_7229);
nand U8929 (N_8929,N_6763,N_6405);
and U8930 (N_8930,N_7241,N_6839);
or U8931 (N_8931,N_6052,N_6078);
or U8932 (N_8932,N_6885,N_7070);
xor U8933 (N_8933,N_6372,N_7371);
nand U8934 (N_8934,N_6688,N_6521);
and U8935 (N_8935,N_6832,N_6150);
nor U8936 (N_8936,N_6208,N_6046);
or U8937 (N_8937,N_6893,N_6839);
xor U8938 (N_8938,N_7495,N_6951);
or U8939 (N_8939,N_6014,N_7190);
or U8940 (N_8940,N_6593,N_6470);
xnor U8941 (N_8941,N_6504,N_7443);
and U8942 (N_8942,N_6910,N_7235);
xnor U8943 (N_8943,N_7422,N_6219);
xor U8944 (N_8944,N_6440,N_7305);
and U8945 (N_8945,N_6978,N_7045);
xnor U8946 (N_8946,N_7388,N_6015);
xor U8947 (N_8947,N_7261,N_6863);
nor U8948 (N_8948,N_6211,N_7375);
xor U8949 (N_8949,N_6629,N_6077);
nor U8950 (N_8950,N_6456,N_7261);
nor U8951 (N_8951,N_6452,N_6983);
nor U8952 (N_8952,N_7114,N_7280);
and U8953 (N_8953,N_7053,N_6940);
nand U8954 (N_8954,N_7389,N_6350);
nand U8955 (N_8955,N_6087,N_7280);
xnor U8956 (N_8956,N_7363,N_7438);
nand U8957 (N_8957,N_7062,N_6847);
nor U8958 (N_8958,N_7463,N_7294);
nor U8959 (N_8959,N_6937,N_7193);
xor U8960 (N_8960,N_6048,N_7020);
or U8961 (N_8961,N_6568,N_7011);
xnor U8962 (N_8962,N_7203,N_6506);
nand U8963 (N_8963,N_6684,N_6730);
nand U8964 (N_8964,N_6748,N_6964);
and U8965 (N_8965,N_6529,N_7494);
nor U8966 (N_8966,N_6391,N_6215);
nand U8967 (N_8967,N_6960,N_7013);
nor U8968 (N_8968,N_7055,N_7065);
nor U8969 (N_8969,N_6370,N_6695);
xor U8970 (N_8970,N_7310,N_6100);
and U8971 (N_8971,N_6999,N_7376);
or U8972 (N_8972,N_7160,N_6155);
and U8973 (N_8973,N_7270,N_6031);
xnor U8974 (N_8974,N_7453,N_6449);
nand U8975 (N_8975,N_7189,N_7499);
xor U8976 (N_8976,N_6544,N_6867);
xor U8977 (N_8977,N_6422,N_6702);
xnor U8978 (N_8978,N_6114,N_6626);
nand U8979 (N_8979,N_6698,N_6122);
nand U8980 (N_8980,N_6185,N_7003);
or U8981 (N_8981,N_6772,N_6148);
nor U8982 (N_8982,N_7422,N_6642);
nor U8983 (N_8983,N_6377,N_6259);
nor U8984 (N_8984,N_6542,N_6675);
nand U8985 (N_8985,N_7328,N_6989);
or U8986 (N_8986,N_6886,N_6972);
nand U8987 (N_8987,N_7445,N_7152);
nor U8988 (N_8988,N_7140,N_6370);
or U8989 (N_8989,N_7451,N_7395);
and U8990 (N_8990,N_7081,N_6906);
nand U8991 (N_8991,N_6026,N_6137);
nand U8992 (N_8992,N_6470,N_7327);
nand U8993 (N_8993,N_6645,N_6769);
or U8994 (N_8994,N_6436,N_6113);
nor U8995 (N_8995,N_6640,N_6337);
nor U8996 (N_8996,N_6336,N_7003);
nor U8997 (N_8997,N_7154,N_7394);
nor U8998 (N_8998,N_6765,N_6451);
nand U8999 (N_8999,N_6226,N_7297);
nand U9000 (N_9000,N_7868,N_8500);
nor U9001 (N_9001,N_7738,N_7861);
nor U9002 (N_9002,N_7545,N_8470);
or U9003 (N_9003,N_8450,N_8186);
or U9004 (N_9004,N_8385,N_8201);
xnor U9005 (N_9005,N_8709,N_8603);
nor U9006 (N_9006,N_8409,N_7790);
nand U9007 (N_9007,N_7663,N_7961);
and U9008 (N_9008,N_7804,N_7743);
nor U9009 (N_9009,N_8633,N_8661);
and U9010 (N_9010,N_8260,N_8862);
and U9011 (N_9011,N_8258,N_7864);
nand U9012 (N_9012,N_8317,N_8087);
or U9013 (N_9013,N_8054,N_8442);
nor U9014 (N_9014,N_8535,N_8886);
and U9015 (N_9015,N_8895,N_8935);
xnor U9016 (N_9016,N_8553,N_8524);
nor U9017 (N_9017,N_8520,N_8991);
or U9018 (N_9018,N_8198,N_8729);
nand U9019 (N_9019,N_8602,N_8584);
xor U9020 (N_9020,N_8074,N_8383);
nand U9021 (N_9021,N_8312,N_8680);
and U9022 (N_9022,N_8872,N_7635);
or U9023 (N_9023,N_8767,N_8339);
xnor U9024 (N_9024,N_7816,N_8654);
xor U9025 (N_9025,N_7955,N_7833);
or U9026 (N_9026,N_8301,N_7562);
or U9027 (N_9027,N_8333,N_7681);
or U9028 (N_9028,N_8364,N_8504);
or U9029 (N_9029,N_8901,N_8989);
or U9030 (N_9030,N_8629,N_8229);
and U9031 (N_9031,N_7968,N_7696);
xnor U9032 (N_9032,N_8119,N_8016);
xnor U9033 (N_9033,N_7846,N_7615);
nor U9034 (N_9034,N_7617,N_7783);
and U9035 (N_9035,N_8243,N_8627);
xor U9036 (N_9036,N_8411,N_8847);
nor U9037 (N_9037,N_8340,N_7737);
and U9038 (N_9038,N_8248,N_8064);
nor U9039 (N_9039,N_7597,N_8141);
and U9040 (N_9040,N_8879,N_8306);
nand U9041 (N_9041,N_8816,N_8281);
and U9042 (N_9042,N_8583,N_7902);
xor U9043 (N_9043,N_8342,N_8365);
xnor U9044 (N_9044,N_7767,N_7975);
and U9045 (N_9045,N_8381,N_8022);
and U9046 (N_9046,N_7660,N_8939);
nor U9047 (N_9047,N_8369,N_8486);
nand U9048 (N_9048,N_8880,N_7556);
or U9049 (N_9049,N_7578,N_8776);
nand U9050 (N_9050,N_8058,N_8720);
nor U9051 (N_9051,N_8687,N_8060);
nor U9052 (N_9052,N_8110,N_7772);
nand U9053 (N_9053,N_8810,N_8589);
nand U9054 (N_9054,N_8518,N_7752);
nor U9055 (N_9055,N_7732,N_7634);
nand U9056 (N_9056,N_7843,N_7745);
and U9057 (N_9057,N_7700,N_8594);
xnor U9058 (N_9058,N_7755,N_7910);
xnor U9059 (N_9059,N_7870,N_8351);
or U9060 (N_9060,N_8362,N_8797);
or U9061 (N_9061,N_8322,N_8097);
xnor U9062 (N_9062,N_7820,N_8835);
nor U9063 (N_9063,N_8725,N_8346);
xor U9064 (N_9064,N_8618,N_7609);
and U9065 (N_9065,N_8600,N_8354);
nor U9066 (N_9066,N_8465,N_8832);
xnor U9067 (N_9067,N_8984,N_7920);
nor U9068 (N_9068,N_8021,N_7805);
or U9069 (N_9069,N_8719,N_7942);
nor U9070 (N_9070,N_8491,N_8531);
xnor U9071 (N_9071,N_8757,N_7728);
or U9072 (N_9072,N_8082,N_8636);
or U9073 (N_9073,N_8386,N_8161);
and U9074 (N_9074,N_8623,N_8724);
xnor U9075 (N_9075,N_8887,N_8614);
and U9076 (N_9076,N_8891,N_7701);
xor U9077 (N_9077,N_8608,N_8349);
nand U9078 (N_9078,N_8184,N_8360);
and U9079 (N_9079,N_8404,N_7649);
nor U9080 (N_9080,N_7631,N_7644);
or U9081 (N_9081,N_7552,N_7559);
nor U9082 (N_9082,N_8328,N_7903);
nand U9083 (N_9083,N_8995,N_8451);
or U9084 (N_9084,N_8726,N_7795);
nor U9085 (N_9085,N_8838,N_8239);
nor U9086 (N_9086,N_8131,N_7717);
and U9087 (N_9087,N_8631,N_8336);
and U9088 (N_9088,N_8663,N_8662);
xor U9089 (N_9089,N_8809,N_7827);
xor U9090 (N_9090,N_8867,N_8568);
nor U9091 (N_9091,N_8669,N_8721);
nand U9092 (N_9092,N_8965,N_8051);
and U9093 (N_9093,N_8917,N_7886);
xor U9094 (N_9094,N_8447,N_8743);
xnor U9095 (N_9095,N_8197,N_8413);
xor U9096 (N_9096,N_8483,N_8941);
nand U9097 (N_9097,N_8124,N_8424);
or U9098 (N_9098,N_8780,N_8151);
or U9099 (N_9099,N_8521,N_8812);
or U9100 (N_9100,N_8616,N_7654);
and U9101 (N_9101,N_8546,N_8391);
or U9102 (N_9102,N_8166,N_8502);
xor U9103 (N_9103,N_7514,N_7564);
nand U9104 (N_9104,N_8659,N_8731);
or U9105 (N_9105,N_8821,N_7584);
nor U9106 (N_9106,N_8773,N_8240);
nor U9107 (N_9107,N_7831,N_8918);
nand U9108 (N_9108,N_7930,N_8893);
xor U9109 (N_9109,N_8270,N_8796);
nand U9110 (N_9110,N_8304,N_8075);
and U9111 (N_9111,N_8655,N_7582);
nand U9112 (N_9112,N_7711,N_7802);
xor U9113 (N_9113,N_7810,N_7506);
nor U9114 (N_9114,N_7665,N_8287);
and U9115 (N_9115,N_7759,N_8121);
or U9116 (N_9116,N_8758,N_8059);
nand U9117 (N_9117,N_8220,N_8990);
nor U9118 (N_9118,N_7744,N_7554);
xor U9119 (N_9119,N_8096,N_7957);
xnor U9120 (N_9120,N_7595,N_7551);
or U9121 (N_9121,N_8018,N_8421);
nand U9122 (N_9122,N_8851,N_8238);
xor U9123 (N_9123,N_8936,N_8547);
nor U9124 (N_9124,N_8418,N_8679);
xor U9125 (N_9125,N_8739,N_8505);
xnor U9126 (N_9126,N_7918,N_8723);
nand U9127 (N_9127,N_8045,N_8537);
and U9128 (N_9128,N_8250,N_7958);
or U9129 (N_9129,N_8690,N_7619);
and U9130 (N_9130,N_8760,N_8974);
nor U9131 (N_9131,N_7898,N_8705);
or U9132 (N_9132,N_7651,N_7658);
nor U9133 (N_9133,N_8698,N_7799);
and U9134 (N_9134,N_8696,N_8980);
or U9135 (N_9135,N_8044,N_8792);
xnor U9136 (N_9136,N_8030,N_8653);
and U9137 (N_9137,N_8476,N_8327);
or U9138 (N_9138,N_8083,N_8367);
or U9139 (N_9139,N_8009,N_8912);
nand U9140 (N_9140,N_8909,N_7897);
or U9141 (N_9141,N_8802,N_8630);
xor U9142 (N_9142,N_8542,N_7912);
and U9143 (N_9143,N_8474,N_8291);
nor U9144 (N_9144,N_7726,N_7785);
and U9145 (N_9145,N_8677,N_8707);
and U9146 (N_9146,N_7927,N_8228);
xnor U9147 (N_9147,N_8192,N_8975);
nor U9148 (N_9148,N_8410,N_8251);
or U9149 (N_9149,N_8130,N_8766);
nand U9150 (N_9150,N_7934,N_8566);
and U9151 (N_9151,N_8337,N_8484);
nand U9152 (N_9152,N_8350,N_8013);
nor U9153 (N_9153,N_7685,N_8038);
xnor U9154 (N_9154,N_7760,N_8899);
xnor U9155 (N_9155,N_7561,N_8755);
xor U9156 (N_9156,N_8420,N_8273);
nor U9157 (N_9157,N_8208,N_7567);
and U9158 (N_9158,N_8193,N_7707);
nor U9159 (N_9159,N_7781,N_7867);
xnor U9160 (N_9160,N_8034,N_7842);
xnor U9161 (N_9161,N_8882,N_8138);
nor U9162 (N_9162,N_8977,N_8530);
and U9163 (N_9163,N_8092,N_8162);
nor U9164 (N_9164,N_8836,N_8923);
and U9165 (N_9165,N_8508,N_8276);
or U9166 (N_9166,N_8751,N_7756);
or U9167 (N_9167,N_8914,N_7940);
xor U9168 (N_9168,N_7991,N_7812);
or U9169 (N_9169,N_7819,N_8469);
nor U9170 (N_9170,N_8014,N_8501);
nand U9171 (N_9171,N_8519,N_8468);
nor U9172 (N_9172,N_8570,N_8005);
xnor U9173 (N_9173,N_8595,N_8642);
nand U9174 (N_9174,N_7546,N_7608);
and U9175 (N_9175,N_8405,N_8300);
nand U9176 (N_9176,N_8157,N_8310);
nor U9177 (N_9177,N_8299,N_8894);
and U9178 (N_9178,N_8324,N_8916);
nor U9179 (N_9179,N_8461,N_7645);
and U9180 (N_9180,N_8403,N_8429);
nand U9181 (N_9181,N_8645,N_7880);
and U9182 (N_9182,N_8940,N_8194);
or U9183 (N_9183,N_8428,N_8154);
xnor U9184 (N_9184,N_7593,N_8952);
and U9185 (N_9185,N_7600,N_8219);
xnor U9186 (N_9186,N_7893,N_7703);
and U9187 (N_9187,N_7577,N_7951);
xor U9188 (N_9188,N_8670,N_8311);
and U9189 (N_9189,N_8889,N_8998);
xnor U9190 (N_9190,N_8826,N_8433);
nor U9191 (N_9191,N_8741,N_7549);
or U9192 (N_9192,N_7950,N_8041);
or U9193 (N_9193,N_8233,N_7656);
nand U9194 (N_9194,N_8249,N_7750);
or U9195 (N_9195,N_8230,N_8778);
and U9196 (N_9196,N_8155,N_7859);
xnor U9197 (N_9197,N_8949,N_8804);
nor U9198 (N_9198,N_8791,N_8254);
nor U9199 (N_9199,N_8906,N_7922);
xor U9200 (N_9200,N_8763,N_8609);
and U9201 (N_9201,N_7693,N_8844);
xnor U9202 (N_9202,N_8575,N_8691);
nor U9203 (N_9203,N_8319,N_7691);
nor U9204 (N_9204,N_8070,N_7543);
xnor U9205 (N_9205,N_7839,N_8189);
and U9206 (N_9206,N_8203,N_8762);
xor U9207 (N_9207,N_8928,N_8168);
nor U9208 (N_9208,N_8375,N_8591);
nand U9209 (N_9209,N_8540,N_7550);
and U9210 (N_9210,N_7835,N_7736);
xor U9211 (N_9211,N_8577,N_8167);
xor U9212 (N_9212,N_8264,N_7882);
xor U9213 (N_9213,N_7581,N_8649);
or U9214 (N_9214,N_7747,N_7618);
xor U9215 (N_9215,N_7894,N_7673);
and U9216 (N_9216,N_8997,N_7964);
nor U9217 (N_9217,N_8139,N_8487);
nand U9218 (N_9218,N_7959,N_8266);
or U9219 (N_9219,N_8068,N_8937);
xnor U9220 (N_9220,N_8771,N_8958);
nand U9221 (N_9221,N_8149,N_8527);
nor U9222 (N_9222,N_8283,N_8973);
nor U9223 (N_9223,N_8047,N_8067);
and U9224 (N_9224,N_8927,N_8626);
nand U9225 (N_9225,N_7938,N_8303);
nor U9226 (N_9226,N_7509,N_7683);
xor U9227 (N_9227,N_8695,N_8113);
nor U9228 (N_9228,N_8561,N_7899);
xnor U9229 (N_9229,N_8744,N_7505);
and U9230 (N_9230,N_8789,N_7758);
xnor U9231 (N_9231,N_8828,N_8948);
xor U9232 (N_9232,N_8062,N_8875);
nor U9233 (N_9233,N_7587,N_8427);
nor U9234 (N_9234,N_8190,N_8267);
nand U9235 (N_9235,N_7563,N_7974);
or U9236 (N_9236,N_8775,N_7840);
nand U9237 (N_9237,N_8482,N_7972);
nor U9238 (N_9238,N_7762,N_8255);
nor U9239 (N_9239,N_8379,N_8883);
nor U9240 (N_9240,N_8971,N_8643);
or U9241 (N_9241,N_8782,N_7935);
or U9242 (N_9242,N_8722,N_7829);
nand U9243 (N_9243,N_8459,N_8235);
xnor U9244 (N_9244,N_8993,N_8492);
and U9245 (N_9245,N_7932,N_8770);
nor U9246 (N_9246,N_8332,N_7697);
and U9247 (N_9247,N_8573,N_8697);
or U9248 (N_9248,N_8236,N_8206);
xor U9249 (N_9249,N_8903,N_8942);
nand U9250 (N_9250,N_8033,N_8232);
nor U9251 (N_9251,N_7792,N_8684);
nand U9252 (N_9252,N_7800,N_7858);
and U9253 (N_9253,N_8640,N_8628);
nand U9254 (N_9254,N_8839,N_7716);
xnor U9255 (N_9255,N_8999,N_7588);
nor U9256 (N_9256,N_8037,N_7692);
xor U9257 (N_9257,N_7905,N_8372);
nor U9258 (N_9258,N_8026,N_7598);
or U9259 (N_9259,N_7798,N_8109);
nor U9260 (N_9260,N_8558,N_8529);
nand U9261 (N_9261,N_8079,N_7768);
nor U9262 (N_9262,N_8921,N_8930);
nand U9263 (N_9263,N_7636,N_8713);
nor U9264 (N_9264,N_7949,N_7818);
nand U9265 (N_9265,N_7530,N_8646);
nand U9266 (N_9266,N_8377,N_7647);
nand U9267 (N_9267,N_7945,N_8550);
nor U9268 (N_9268,N_8185,N_7560);
or U9269 (N_9269,N_8737,N_7969);
nor U9270 (N_9270,N_8897,N_8904);
or U9271 (N_9271,N_7933,N_8822);
nand U9272 (N_9272,N_8860,N_8742);
xnor U9273 (N_9273,N_7527,N_8178);
and U9274 (N_9274,N_7815,N_8960);
xnor U9275 (N_9275,N_8036,N_7766);
or U9276 (N_9276,N_8100,N_8514);
and U9277 (N_9277,N_8020,N_8225);
xnor U9278 (N_9278,N_8134,N_7834);
nand U9279 (N_9279,N_8331,N_7718);
or U9280 (N_9280,N_7796,N_7881);
and U9281 (N_9281,N_8783,N_7915);
or U9282 (N_9282,N_7583,N_7540);
nor U9283 (N_9283,N_7962,N_8158);
and U9284 (N_9284,N_7695,N_8601);
xnor U9285 (N_9285,N_8445,N_7601);
and U9286 (N_9286,N_8682,N_8479);
xnor U9287 (N_9287,N_8024,N_8806);
or U9288 (N_9288,N_7978,N_8978);
xnor U9289 (N_9289,N_8132,N_7607);
nor U9290 (N_9290,N_8922,N_7811);
and U9291 (N_9291,N_7592,N_8523);
and U9292 (N_9292,N_7642,N_8261);
xnor U9293 (N_9293,N_8147,N_8126);
nor U9294 (N_9294,N_8736,N_8881);
nand U9295 (N_9295,N_8869,N_7973);
nand U9296 (N_9296,N_7669,N_8086);
nor U9297 (N_9297,N_8006,N_7960);
nand U9298 (N_9298,N_8408,N_7746);
xor U9299 (N_9299,N_8069,N_8543);
xnor U9300 (N_9300,N_8344,N_7875);
nand U9301 (N_9301,N_8257,N_8039);
nand U9302 (N_9302,N_7591,N_8785);
xnor U9303 (N_9303,N_8188,N_8081);
nor U9304 (N_9304,N_8979,N_8911);
nand U9305 (N_9305,N_8905,N_7926);
and U9306 (N_9306,N_8104,N_8735);
or U9307 (N_9307,N_7566,N_8422);
and U9308 (N_9308,N_8888,N_7944);
nand U9309 (N_9309,N_7794,N_8323);
nand U9310 (N_9310,N_8624,N_8610);
or U9311 (N_9311,N_8683,N_7866);
nand U9312 (N_9312,N_8604,N_7638);
and U9313 (N_9313,N_8309,N_8226);
nor U9314 (N_9314,N_8795,N_8416);
and U9315 (N_9315,N_8641,N_7510);
nand U9316 (N_9316,N_8046,N_8652);
or U9317 (N_9317,N_8900,N_8085);
nor U9318 (N_9318,N_8938,N_8480);
nand U9319 (N_9319,N_7605,N_7965);
xnor U9320 (N_9320,N_7535,N_7518);
nand U9321 (N_9321,N_8032,N_7911);
nand U9322 (N_9322,N_7719,N_7573);
nor U9323 (N_9323,N_7906,N_8140);
nor U9324 (N_9324,N_8135,N_8846);
or U9325 (N_9325,N_8932,N_7900);
nand U9326 (N_9326,N_8571,N_7849);
xnor U9327 (N_9327,N_8988,N_7873);
xor U9328 (N_9328,N_8015,N_7572);
or U9329 (N_9329,N_8439,N_7712);
xor U9330 (N_9330,N_8842,N_7739);
nand U9331 (N_9331,N_8008,N_8943);
nor U9332 (N_9332,N_7702,N_7925);
xor U9333 (N_9333,N_8237,N_8982);
xnor U9334 (N_9334,N_8892,N_8656);
xnor U9335 (N_9335,N_8803,N_8195);
or U9336 (N_9336,N_7603,N_7721);
nor U9337 (N_9337,N_8554,N_8288);
nor U9338 (N_9338,N_7836,N_8638);
nand U9339 (N_9339,N_8823,N_8865);
or U9340 (N_9340,N_7513,N_7780);
nand U9341 (N_9341,N_7534,N_8749);
nor U9342 (N_9342,N_8738,N_8830);
or U9343 (N_9343,N_8455,N_8644);
nor U9344 (N_9344,N_8613,N_8790);
or U9345 (N_9345,N_8137,N_8578);
nand U9346 (N_9346,N_8448,N_7878);
nor U9347 (N_9347,N_8902,N_7801);
nand U9348 (N_9348,N_7565,N_8868);
or U9349 (N_9349,N_7710,N_8878);
and U9350 (N_9350,N_7909,N_8473);
nand U9351 (N_9351,N_8710,N_7708);
nand U9352 (N_9352,N_8740,N_8817);
nand U9353 (N_9353,N_8370,N_8080);
xnor U9354 (N_9354,N_7919,N_7659);
xnor U9355 (N_9355,N_7524,N_8551);
or U9356 (N_9356,N_8443,N_8389);
xor U9357 (N_9357,N_7948,N_7981);
nor U9358 (N_9358,N_8384,N_7853);
nand U9359 (N_9359,N_8689,N_8423);
nand U9360 (N_9360,N_8481,N_7825);
nor U9361 (N_9361,N_8477,N_8378);
or U9362 (N_9362,N_8338,N_8102);
xor U9363 (N_9363,N_7672,N_7734);
xnor U9364 (N_9364,N_8211,N_8456);
nor U9365 (N_9365,N_8127,N_8048);
xor U9366 (N_9366,N_7625,N_8286);
xor U9367 (N_9367,N_7862,N_8588);
nand U9368 (N_9368,N_8392,N_7500);
xnor U9369 (N_9369,N_8325,N_8976);
and U9370 (N_9370,N_8136,N_8801);
or U9371 (N_9371,N_8647,N_7520);
xnor U9372 (N_9372,N_8981,N_8268);
nand U9373 (N_9373,N_8125,N_7684);
nand U9374 (N_9374,N_8296,N_8221);
xor U9375 (N_9375,N_7620,N_8387);
nor U9376 (N_9376,N_8056,N_8269);
nand U9377 (N_9377,N_7889,N_8066);
xnor U9378 (N_9378,N_7943,N_8253);
and U9379 (N_9379,N_8884,N_8498);
nand U9380 (N_9380,N_8329,N_7727);
nor U9381 (N_9381,N_7860,N_7763);
nand U9382 (N_9382,N_8569,N_7773);
or U9383 (N_9383,N_8825,N_8307);
xor U9384 (N_9384,N_7516,N_7775);
nor U9385 (N_9385,N_7511,N_8970);
nand U9386 (N_9386,N_8664,N_8494);
xnor U9387 (N_9387,N_7694,N_7674);
xnor U9388 (N_9388,N_8295,N_8478);
nor U9389 (N_9389,N_8793,N_8335);
nand U9390 (N_9390,N_7686,N_8284);
xnor U9391 (N_9391,N_7952,N_7533);
nor U9392 (N_9392,N_7996,N_7753);
or U9393 (N_9393,N_7640,N_8040);
or U9394 (N_9394,N_7709,N_7503);
nand U9395 (N_9395,N_8660,N_8095);
nor U9396 (N_9396,N_8371,N_8896);
and U9397 (N_9397,N_8212,N_7980);
nand U9398 (N_9398,N_8358,N_8497);
nand U9399 (N_9399,N_7725,N_8813);
xnor U9400 (N_9400,N_8272,N_8599);
nor U9401 (N_9401,N_8262,N_7998);
xor U9402 (N_9402,N_8774,N_8637);
or U9403 (N_9403,N_7629,N_7537);
and U9404 (N_9404,N_8858,N_8648);
nor U9405 (N_9405,N_8597,N_7985);
nor U9406 (N_9406,N_7913,N_8992);
or U9407 (N_9407,N_8945,N_7690);
or U9408 (N_9408,N_7544,N_8907);
nor U9409 (N_9409,N_7512,N_7914);
xnor U9410 (N_9410,N_8674,N_8532);
and U9411 (N_9411,N_8460,N_7664);
and U9412 (N_9412,N_8398,N_7541);
nor U9413 (N_9413,N_7786,N_7515);
nand U9414 (N_9414,N_8947,N_7602);
nor U9415 (N_9415,N_8007,N_8968);
nor U9416 (N_9416,N_8853,N_8929);
and U9417 (N_9417,N_8877,N_8012);
nand U9418 (N_9418,N_8073,N_8576);
xnor U9419 (N_9419,N_7992,N_8366);
or U9420 (N_9420,N_7813,N_7953);
xor U9421 (N_9421,N_7988,N_8171);
or U9422 (N_9422,N_8787,N_8934);
xnor U9423 (N_9423,N_8150,N_7883);
or U9424 (N_9424,N_8142,N_8815);
xnor U9425 (N_9425,N_8890,N_8091);
or U9426 (N_9426,N_8466,N_7863);
or U9427 (N_9427,N_8784,N_8105);
and U9428 (N_9428,N_8632,N_8293);
and U9429 (N_9429,N_7528,N_8053);
or U9430 (N_9430,N_8557,N_8457);
nor U9431 (N_9431,N_8088,N_7806);
nor U9432 (N_9432,N_7977,N_8635);
and U9433 (N_9433,N_8857,N_8042);
nand U9434 (N_9434,N_8885,N_8128);
nor U9435 (N_9435,N_8756,N_7838);
nand U9436 (N_9436,N_7966,N_8170);
or U9437 (N_9437,N_7754,N_8926);
and U9438 (N_9438,N_8152,N_8217);
nor U9439 (N_9439,N_7699,N_7999);
and U9440 (N_9440,N_8357,N_8084);
nor U9441 (N_9441,N_8944,N_8620);
nand U9442 (N_9442,N_8446,N_7847);
and U9443 (N_9443,N_8715,N_7793);
nor U9444 (N_9444,N_7621,N_8049);
xnor U9445 (N_9445,N_7823,N_8814);
nor U9446 (N_9446,N_7904,N_8376);
or U9447 (N_9447,N_8436,N_8593);
xor U9448 (N_9448,N_8380,N_7713);
nand U9449 (N_9449,N_8290,N_7655);
nand U9450 (N_9450,N_7797,N_8625);
nand U9451 (N_9451,N_7937,N_7715);
nand U9452 (N_9452,N_8464,N_8967);
and U9453 (N_9453,N_8545,N_8223);
and U9454 (N_9454,N_8396,N_8256);
nor U9455 (N_9455,N_7890,N_7887);
nor U9456 (N_9456,N_7924,N_8651);
and U9457 (N_9457,N_8607,N_7507);
or U9458 (N_9458,N_8750,N_7888);
xnor U9459 (N_9459,N_8702,N_8908);
xnor U9460 (N_9460,N_8298,N_8122);
and U9461 (N_9461,N_7956,N_8289);
or U9462 (N_9462,N_7908,N_7984);
nor U9463 (N_9463,N_7733,N_8712);
and U9464 (N_9464,N_8315,N_7523);
or U9465 (N_9465,N_7627,N_8898);
xnor U9466 (N_9466,N_8834,N_8177);
or U9467 (N_9467,N_7570,N_8764);
nand U9468 (N_9468,N_7947,N_8592);
nand U9469 (N_9469,N_7994,N_8913);
nor U9470 (N_9470,N_8503,N_7782);
or U9471 (N_9471,N_8820,N_8094);
or U9472 (N_9472,N_8347,N_8247);
nand U9473 (N_9473,N_8169,N_8866);
or U9474 (N_9474,N_8129,N_7871);
xor U9475 (N_9475,N_7865,N_8285);
nor U9476 (N_9476,N_8849,N_8556);
and U9477 (N_9477,N_7874,N_8686);
and U9478 (N_9478,N_8574,N_7705);
xnor U9479 (N_9479,N_8522,N_7643);
nand U9480 (N_9480,N_8055,N_8876);
nor U9481 (N_9481,N_7730,N_8539);
nand U9482 (N_9482,N_8533,N_7675);
xor U9483 (N_9483,N_8987,N_8271);
or U9484 (N_9484,N_7923,N_8390);
nand U9485 (N_9485,N_7826,N_7661);
xnor U9486 (N_9486,N_8297,N_8964);
nor U9487 (N_9487,N_8515,N_8714);
or U9488 (N_9488,N_8181,N_8187);
and U9489 (N_9489,N_7650,N_8565);
and U9490 (N_9490,N_8579,N_8116);
nand U9491 (N_9491,N_7854,N_8244);
nor U9492 (N_9492,N_8259,N_8330);
nor U9493 (N_9493,N_8493,N_8402);
nand U9494 (N_9494,N_8246,N_8164);
or U9495 (N_9495,N_8078,N_8856);
nand U9496 (N_9496,N_7677,N_7742);
nor U9497 (N_9497,N_8510,N_7706);
nand U9498 (N_9498,N_7639,N_7616);
xor U9499 (N_9499,N_7828,N_8061);
xor U9500 (N_9500,N_7907,N_7731);
and U9501 (N_9501,N_8214,N_7596);
and U9502 (N_9502,N_8076,N_8855);
nand U9503 (N_9503,N_8560,N_8117);
and U9504 (N_9504,N_7626,N_8210);
or U9505 (N_9505,N_7821,N_8000);
xor U9506 (N_9506,N_8798,N_8475);
and U9507 (N_9507,N_8861,N_8231);
nand U9508 (N_9508,N_7749,N_7832);
nor U9509 (N_9509,N_8174,N_8222);
and U9510 (N_9510,N_8768,N_8202);
and U9511 (N_9511,N_8996,N_7680);
nor U9512 (N_9512,N_8444,N_7856);
nor U9513 (N_9513,N_8148,N_8685);
xor U9514 (N_9514,N_8434,N_7921);
or U9515 (N_9515,N_8753,N_8598);
and U9516 (N_9516,N_7594,N_8419);
or U9517 (N_9517,N_8748,N_8057);
nor U9518 (N_9518,N_8777,N_7579);
or U9519 (N_9519,N_8292,N_8745);
or U9520 (N_9520,N_8345,N_8986);
or U9521 (N_9521,N_8302,N_8837);
nor U9522 (N_9522,N_7982,N_8526);
nand U9523 (N_9523,N_7613,N_8808);
or U9524 (N_9524,N_7536,N_8772);
and U9525 (N_9525,N_8536,N_7771);
nand U9526 (N_9526,N_8692,N_8512);
nand U9527 (N_9527,N_8567,N_7641);
xnor U9528 (N_9528,N_8314,N_8694);
xor U9529 (N_9529,N_8093,N_8728);
nor U9530 (N_9530,N_7611,N_8506);
and U9531 (N_9531,N_8454,N_8280);
or U9532 (N_9532,N_8972,N_8108);
nand U9533 (N_9533,N_8919,N_7539);
xnor U9534 (N_9534,N_8035,N_7789);
xnor U9535 (N_9535,N_8432,N_8352);
nand U9536 (N_9536,N_8827,N_8462);
xnor U9537 (N_9537,N_8933,N_7590);
nor U9538 (N_9538,N_8534,N_7764);
xnor U9539 (N_9539,N_8752,N_8852);
nor U9540 (N_9540,N_8870,N_8871);
nor U9541 (N_9541,N_7993,N_7769);
nor U9542 (N_9542,N_7936,N_7622);
or U9543 (N_9543,N_8549,N_8165);
or U9544 (N_9544,N_8580,N_8509);
nor U9545 (N_9545,N_8089,N_8874);
or U9546 (N_9546,N_8294,N_8417);
or U9547 (N_9547,N_8017,N_8688);
nor U9548 (N_9548,N_7954,N_8572);
and U9549 (N_9549,N_7970,N_8438);
nor U9550 (N_9550,N_8800,N_7928);
xnor U9551 (N_9551,N_7885,N_8356);
or U9552 (N_9552,N_8955,N_8393);
and U9553 (N_9553,N_8316,N_7896);
nor U9554 (N_9554,N_8490,N_8586);
nor U9555 (N_9555,N_7877,N_8397);
xor U9556 (N_9556,N_7585,N_8488);
and U9557 (N_9557,N_8564,N_7735);
xor U9558 (N_9558,N_7501,N_8043);
or U9559 (N_9559,N_8489,N_7990);
nor U9560 (N_9560,N_8472,N_8180);
nor U9561 (N_9561,N_8458,N_8209);
and U9562 (N_9562,N_8156,N_8234);
nor U9563 (N_9563,N_8845,N_8394);
nor U9564 (N_9564,N_8191,N_8708);
xor U9565 (N_9565,N_8452,N_7869);
nor U9566 (N_9566,N_8098,N_7668);
nand U9567 (N_9567,N_8023,N_8824);
nand U9568 (N_9568,N_7704,N_7963);
or U9569 (N_9569,N_7748,N_8496);
nand U9570 (N_9570,N_8650,N_8587);
xnor U9571 (N_9571,N_7698,N_8681);
xnor U9572 (N_9572,N_8555,N_8175);
or U9573 (N_9573,N_7648,N_8924);
nand U9574 (N_9574,N_8673,N_7729);
or U9575 (N_9575,N_7822,N_8538);
nor U9576 (N_9576,N_8807,N_8200);
nand U9577 (N_9577,N_8308,N_7995);
nand U9578 (N_9578,N_8811,N_8562);
and U9579 (N_9579,N_8111,N_8407);
nor U9580 (N_9580,N_8954,N_8961);
nor U9581 (N_9581,N_7722,N_8265);
and U9582 (N_9582,N_8263,N_7687);
and U9583 (N_9583,N_8359,N_8153);
and U9584 (N_9584,N_7844,N_8548);
and U9585 (N_9585,N_8010,N_8011);
and U9586 (N_9586,N_7971,N_8415);
nand U9587 (N_9587,N_8956,N_7547);
nand U9588 (N_9588,N_7845,N_8321);
and U9589 (N_9589,N_7946,N_8326);
and U9590 (N_9590,N_7612,N_8511);
or U9591 (N_9591,N_8090,N_7809);
nor U9592 (N_9592,N_8985,N_7803);
xor U9593 (N_9593,N_8318,N_7610);
nand U9594 (N_9594,N_8507,N_7569);
or U9595 (N_9595,N_8279,N_8133);
and U9596 (N_9596,N_8112,N_8700);
nand U9597 (N_9597,N_7628,N_8590);
nor U9598 (N_9598,N_8946,N_7557);
or U9599 (N_9599,N_8794,N_7895);
and U9600 (N_9600,N_7624,N_8781);
nand U9601 (N_9601,N_7542,N_8950);
xnor U9602 (N_9602,N_8829,N_8163);
nor U9603 (N_9603,N_8395,N_8959);
xor U9604 (N_9604,N_7667,N_8027);
or U9605 (N_9605,N_7967,N_8453);
nor U9606 (N_9606,N_7941,N_7671);
nor U9607 (N_9607,N_7633,N_8274);
or U9608 (N_9608,N_7580,N_7526);
or U9609 (N_9609,N_8159,N_7939);
nand U9610 (N_9610,N_7679,N_7774);
nand U9611 (N_9611,N_8320,N_7519);
and U9612 (N_9612,N_7855,N_8144);
or U9613 (N_9613,N_8622,N_7987);
or U9614 (N_9614,N_7851,N_8788);
nand U9615 (N_9615,N_7632,N_8833);
xor U9616 (N_9616,N_8205,N_8106);
xnor U9617 (N_9617,N_8596,N_8401);
or U9618 (N_9618,N_7777,N_8703);
xnor U9619 (N_9619,N_8848,N_8431);
and U9620 (N_9620,N_8699,N_7857);
and U9621 (N_9621,N_8746,N_8218);
xnor U9622 (N_9622,N_7917,N_7770);
and U9623 (N_9623,N_8204,N_8173);
nor U9624 (N_9624,N_8275,N_7720);
nor U9625 (N_9625,N_7553,N_7646);
xnor U9626 (N_9626,N_8701,N_7614);
xor U9627 (N_9627,N_8541,N_8414);
nand U9628 (N_9628,N_8241,N_8029);
or U9629 (N_9629,N_8818,N_8348);
nor U9630 (N_9630,N_8467,N_8052);
xnor U9631 (N_9631,N_8437,N_8951);
or U9632 (N_9632,N_7751,N_8050);
and U9633 (N_9633,N_8963,N_7521);
nor U9634 (N_9634,N_8841,N_8115);
nand U9635 (N_9635,N_7652,N_8242);
and U9636 (N_9636,N_7637,N_7979);
and U9637 (N_9637,N_8004,N_8585);
or U9638 (N_9638,N_8761,N_8779);
nor U9639 (N_9639,N_7891,N_7986);
and U9640 (N_9640,N_7571,N_7784);
or U9641 (N_9641,N_8957,N_7670);
nand U9642 (N_9642,N_7787,N_8361);
or U9643 (N_9643,N_8305,N_7522);
or U9644 (N_9644,N_8717,N_7558);
nor U9645 (N_9645,N_8611,N_7604);
nand U9646 (N_9646,N_8341,N_8759);
nor U9647 (N_9647,N_8605,N_8671);
and U9648 (N_9648,N_8499,N_8634);
or U9649 (N_9649,N_8374,N_7848);
xnor U9650 (N_9650,N_8382,N_7724);
or U9651 (N_9651,N_7678,N_7723);
xor U9652 (N_9652,N_7630,N_8179);
nor U9653 (N_9653,N_7606,N_7788);
and U9654 (N_9654,N_8843,N_7892);
nand U9655 (N_9655,N_7808,N_8910);
xnor U9656 (N_9656,N_8399,N_8915);
nand U9657 (N_9657,N_8658,N_7901);
nand U9658 (N_9658,N_7599,N_7525);
or U9659 (N_9659,N_8003,N_8864);
nand U9660 (N_9660,N_8966,N_8615);
nor U9661 (N_9661,N_8819,N_8559);
nand U9662 (N_9662,N_7532,N_7548);
xor U9663 (N_9663,N_8730,N_8621);
or U9664 (N_9664,N_8463,N_8612);
and U9665 (N_9665,N_7623,N_7688);
xor U9666 (N_9666,N_8146,N_8435);
or U9667 (N_9667,N_7837,N_8920);
nand U9668 (N_9668,N_7517,N_8859);
and U9669 (N_9669,N_8704,N_8747);
xor U9670 (N_9670,N_8581,N_7576);
or U9671 (N_9671,N_8667,N_8953);
and U9672 (N_9672,N_7574,N_7841);
xnor U9673 (N_9673,N_8400,N_8123);
or U9674 (N_9674,N_7714,N_8831);
xor U9675 (N_9675,N_8118,N_8176);
and U9676 (N_9676,N_8799,N_8207);
and U9677 (N_9677,N_8072,N_7666);
and U9678 (N_9678,N_8019,N_8440);
xor U9679 (N_9679,N_8028,N_8517);
and U9680 (N_9680,N_8353,N_8343);
nor U9681 (N_9681,N_7682,N_8245);
or U9682 (N_9682,N_8199,N_8114);
xnor U9683 (N_9683,N_8716,N_8099);
nor U9684 (N_9684,N_8213,N_8678);
or U9685 (N_9685,N_8665,N_7778);
or U9686 (N_9686,N_8412,N_8182);
nand U9687 (N_9687,N_8754,N_7884);
nand U9688 (N_9688,N_7761,N_8693);
xor U9689 (N_9689,N_8277,N_8227);
and U9690 (N_9690,N_8840,N_8552);
or U9691 (N_9691,N_7791,N_8025);
xor U9692 (N_9692,N_8063,N_8676);
xor U9693 (N_9693,N_8983,N_8363);
or U9694 (N_9694,N_7929,N_8406);
nand U9695 (N_9695,N_7538,N_8582);
nor U9696 (N_9696,N_8513,N_8077);
or U9697 (N_9697,N_8994,N_8001);
nor U9698 (N_9698,N_7830,N_8873);
or U9699 (N_9699,N_8931,N_7817);
or U9700 (N_9700,N_8733,N_8672);
xor U9701 (N_9701,N_8388,N_8160);
and U9702 (N_9702,N_8925,N_8854);
nand U9703 (N_9703,N_8706,N_7568);
nand U9704 (N_9704,N_7740,N_8516);
nor U9705 (N_9705,N_8216,N_8143);
nor U9706 (N_9706,N_8734,N_8765);
nor U9707 (N_9707,N_8334,N_8355);
and U9708 (N_9708,N_7983,N_8368);
nand U9709 (N_9709,N_7586,N_7824);
xnor U9710 (N_9710,N_7850,N_8495);
nand U9711 (N_9711,N_7931,N_7575);
xnor U9712 (N_9712,N_8373,N_7765);
nor U9713 (N_9713,N_8805,N_8425);
or U9714 (N_9714,N_8485,N_8769);
xor U9715 (N_9715,N_7876,N_8101);
and U9716 (N_9716,N_8675,N_8962);
nor U9717 (N_9717,N_7689,N_8426);
nor U9718 (N_9718,N_8619,N_8718);
and U9719 (N_9719,N_8065,N_8031);
nand U9720 (N_9720,N_7589,N_8544);
nand U9721 (N_9721,N_7814,N_7776);
nand U9722 (N_9722,N_8471,N_7989);
or U9723 (N_9723,N_7852,N_8657);
or U9724 (N_9724,N_8666,N_8145);
or U9725 (N_9725,N_8727,N_8224);
nand U9726 (N_9726,N_8430,N_8103);
xnor U9727 (N_9727,N_7976,N_8668);
or U9728 (N_9728,N_7502,N_8732);
or U9729 (N_9729,N_8120,N_8617);
and U9730 (N_9730,N_7997,N_8863);
xnor U9731 (N_9731,N_8252,N_7653);
nor U9732 (N_9732,N_8711,N_7662);
and U9733 (N_9733,N_8278,N_7779);
nand U9734 (N_9734,N_8639,N_8441);
nand U9735 (N_9735,N_7757,N_7657);
xnor U9736 (N_9736,N_8215,N_8002);
and U9737 (N_9737,N_7807,N_8563);
or U9738 (N_9738,N_7504,N_8850);
nor U9739 (N_9739,N_8071,N_7872);
nor U9740 (N_9740,N_7531,N_7555);
nor U9741 (N_9741,N_7676,N_8313);
and U9742 (N_9742,N_8525,N_8196);
nand U9743 (N_9743,N_7879,N_8606);
or U9744 (N_9744,N_8969,N_7508);
xor U9745 (N_9745,N_7741,N_8183);
nor U9746 (N_9746,N_8528,N_7916);
xnor U9747 (N_9747,N_8172,N_8786);
nor U9748 (N_9748,N_8107,N_8449);
and U9749 (N_9749,N_7529,N_8282);
nand U9750 (N_9750,N_7954,N_7737);
nor U9751 (N_9751,N_8667,N_8754);
xor U9752 (N_9752,N_8258,N_8851);
nand U9753 (N_9753,N_8563,N_8660);
or U9754 (N_9754,N_7884,N_8126);
xor U9755 (N_9755,N_8626,N_8226);
and U9756 (N_9756,N_8139,N_7588);
or U9757 (N_9757,N_8787,N_8630);
and U9758 (N_9758,N_8479,N_7567);
nor U9759 (N_9759,N_7550,N_8316);
and U9760 (N_9760,N_8635,N_8722);
nor U9761 (N_9761,N_8295,N_7631);
and U9762 (N_9762,N_8525,N_8860);
and U9763 (N_9763,N_8349,N_7871);
and U9764 (N_9764,N_8323,N_8968);
or U9765 (N_9765,N_8233,N_8258);
nor U9766 (N_9766,N_8420,N_8342);
nand U9767 (N_9767,N_8216,N_8507);
nand U9768 (N_9768,N_8871,N_8928);
and U9769 (N_9769,N_7858,N_7828);
xor U9770 (N_9770,N_8065,N_7666);
xor U9771 (N_9771,N_8676,N_7913);
nand U9772 (N_9772,N_8191,N_7932);
xnor U9773 (N_9773,N_8215,N_7778);
or U9774 (N_9774,N_8326,N_7904);
or U9775 (N_9775,N_7716,N_7918);
and U9776 (N_9776,N_8996,N_8431);
xnor U9777 (N_9777,N_7925,N_7981);
or U9778 (N_9778,N_7974,N_7855);
nand U9779 (N_9779,N_8131,N_7625);
and U9780 (N_9780,N_8390,N_7894);
and U9781 (N_9781,N_7939,N_7508);
nor U9782 (N_9782,N_7627,N_8089);
nor U9783 (N_9783,N_7892,N_8731);
xnor U9784 (N_9784,N_8014,N_7668);
or U9785 (N_9785,N_8159,N_8466);
nand U9786 (N_9786,N_8930,N_8907);
xnor U9787 (N_9787,N_8465,N_7821);
nor U9788 (N_9788,N_8112,N_7714);
nor U9789 (N_9789,N_8099,N_8039);
or U9790 (N_9790,N_8132,N_8128);
xnor U9791 (N_9791,N_8630,N_8881);
nand U9792 (N_9792,N_8439,N_8981);
xnor U9793 (N_9793,N_7752,N_7715);
and U9794 (N_9794,N_8993,N_8948);
nor U9795 (N_9795,N_8215,N_8206);
and U9796 (N_9796,N_7947,N_7699);
nand U9797 (N_9797,N_8823,N_8586);
nand U9798 (N_9798,N_8884,N_8501);
nor U9799 (N_9799,N_8245,N_8022);
xnor U9800 (N_9800,N_7760,N_8924);
nand U9801 (N_9801,N_8599,N_8551);
xor U9802 (N_9802,N_8352,N_8982);
nand U9803 (N_9803,N_7612,N_8871);
nor U9804 (N_9804,N_7751,N_8228);
nor U9805 (N_9805,N_7596,N_8755);
nor U9806 (N_9806,N_7869,N_8844);
or U9807 (N_9807,N_8178,N_8084);
and U9808 (N_9808,N_7924,N_8322);
nand U9809 (N_9809,N_7761,N_8090);
or U9810 (N_9810,N_8928,N_7901);
xnor U9811 (N_9811,N_7614,N_7906);
or U9812 (N_9812,N_8032,N_8484);
nand U9813 (N_9813,N_8211,N_8598);
nand U9814 (N_9814,N_7581,N_7953);
nor U9815 (N_9815,N_8435,N_8736);
xor U9816 (N_9816,N_8221,N_8381);
nor U9817 (N_9817,N_8800,N_7785);
and U9818 (N_9818,N_7643,N_7600);
nand U9819 (N_9819,N_7522,N_8426);
or U9820 (N_9820,N_7683,N_7851);
nand U9821 (N_9821,N_7829,N_7824);
xor U9822 (N_9822,N_8405,N_7780);
xnor U9823 (N_9823,N_7720,N_7904);
nand U9824 (N_9824,N_8132,N_7568);
or U9825 (N_9825,N_8123,N_7929);
nand U9826 (N_9826,N_8658,N_8036);
and U9827 (N_9827,N_7519,N_7549);
nand U9828 (N_9828,N_7518,N_8927);
xor U9829 (N_9829,N_7887,N_8576);
or U9830 (N_9830,N_8685,N_7865);
xnor U9831 (N_9831,N_8461,N_7579);
nand U9832 (N_9832,N_8154,N_8753);
or U9833 (N_9833,N_8701,N_7537);
nand U9834 (N_9834,N_8916,N_8929);
nand U9835 (N_9835,N_7699,N_8270);
and U9836 (N_9836,N_8302,N_7857);
or U9837 (N_9837,N_8138,N_7747);
xor U9838 (N_9838,N_8804,N_7596);
and U9839 (N_9839,N_8777,N_8379);
or U9840 (N_9840,N_8674,N_8172);
nor U9841 (N_9841,N_8403,N_8646);
nand U9842 (N_9842,N_7621,N_8886);
or U9843 (N_9843,N_8502,N_8382);
nand U9844 (N_9844,N_7968,N_8769);
nor U9845 (N_9845,N_8202,N_7906);
nand U9846 (N_9846,N_8811,N_8402);
and U9847 (N_9847,N_8768,N_8114);
and U9848 (N_9848,N_7742,N_7592);
nor U9849 (N_9849,N_8294,N_8827);
nand U9850 (N_9850,N_7832,N_8160);
xnor U9851 (N_9851,N_8426,N_8197);
or U9852 (N_9852,N_8741,N_7645);
xor U9853 (N_9853,N_8350,N_7962);
or U9854 (N_9854,N_7570,N_8854);
nor U9855 (N_9855,N_8712,N_8745);
xor U9856 (N_9856,N_8389,N_8310);
xor U9857 (N_9857,N_8625,N_7532);
and U9858 (N_9858,N_7866,N_7867);
nand U9859 (N_9859,N_8486,N_7868);
or U9860 (N_9860,N_8774,N_7672);
xnor U9861 (N_9861,N_7747,N_7649);
xor U9862 (N_9862,N_8799,N_8098);
nand U9863 (N_9863,N_7791,N_7808);
nand U9864 (N_9864,N_8097,N_8627);
nand U9865 (N_9865,N_8386,N_8461);
nor U9866 (N_9866,N_7950,N_8540);
or U9867 (N_9867,N_7689,N_7593);
and U9868 (N_9868,N_8903,N_8404);
nand U9869 (N_9869,N_8747,N_7666);
nor U9870 (N_9870,N_8582,N_7828);
xor U9871 (N_9871,N_8968,N_8830);
nand U9872 (N_9872,N_7659,N_7700);
xor U9873 (N_9873,N_8097,N_8384);
nand U9874 (N_9874,N_8400,N_7939);
nand U9875 (N_9875,N_7758,N_7854);
nand U9876 (N_9876,N_7565,N_8937);
nor U9877 (N_9877,N_8557,N_8294);
xnor U9878 (N_9878,N_7537,N_7509);
xnor U9879 (N_9879,N_7802,N_8191);
nand U9880 (N_9880,N_8656,N_8056);
and U9881 (N_9881,N_7681,N_8111);
xnor U9882 (N_9882,N_8871,N_7723);
nand U9883 (N_9883,N_7990,N_8209);
nor U9884 (N_9884,N_8688,N_8670);
or U9885 (N_9885,N_8822,N_8161);
or U9886 (N_9886,N_8952,N_8287);
and U9887 (N_9887,N_8993,N_7533);
xor U9888 (N_9888,N_8745,N_8949);
or U9889 (N_9889,N_7602,N_7608);
nor U9890 (N_9890,N_7634,N_7591);
nand U9891 (N_9891,N_8805,N_8053);
nor U9892 (N_9892,N_7897,N_8384);
and U9893 (N_9893,N_7583,N_8294);
and U9894 (N_9894,N_7740,N_7927);
nor U9895 (N_9895,N_8022,N_7653);
and U9896 (N_9896,N_7897,N_7950);
xor U9897 (N_9897,N_8447,N_7857);
or U9898 (N_9898,N_8385,N_8564);
nand U9899 (N_9899,N_8182,N_8074);
and U9900 (N_9900,N_7768,N_7562);
xnor U9901 (N_9901,N_7804,N_7619);
nand U9902 (N_9902,N_8892,N_8527);
nor U9903 (N_9903,N_8585,N_7640);
or U9904 (N_9904,N_8418,N_7761);
nand U9905 (N_9905,N_8996,N_8467);
or U9906 (N_9906,N_7988,N_8931);
or U9907 (N_9907,N_8851,N_8325);
nand U9908 (N_9908,N_8805,N_7532);
nand U9909 (N_9909,N_7558,N_8450);
or U9910 (N_9910,N_8214,N_7956);
nor U9911 (N_9911,N_7559,N_8384);
nand U9912 (N_9912,N_8242,N_8582);
xnor U9913 (N_9913,N_7720,N_7559);
or U9914 (N_9914,N_7841,N_8883);
xnor U9915 (N_9915,N_7996,N_7750);
nor U9916 (N_9916,N_7502,N_7854);
or U9917 (N_9917,N_8977,N_7680);
or U9918 (N_9918,N_7578,N_7916);
and U9919 (N_9919,N_8743,N_8975);
xnor U9920 (N_9920,N_8046,N_8260);
xor U9921 (N_9921,N_8797,N_8592);
xnor U9922 (N_9922,N_8137,N_8781);
nor U9923 (N_9923,N_8656,N_8101);
nand U9924 (N_9924,N_8778,N_8992);
nor U9925 (N_9925,N_8862,N_8196);
xnor U9926 (N_9926,N_8126,N_8647);
nand U9927 (N_9927,N_8035,N_8037);
and U9928 (N_9928,N_8692,N_8617);
and U9929 (N_9929,N_7899,N_8224);
nor U9930 (N_9930,N_8942,N_7645);
and U9931 (N_9931,N_8526,N_8377);
nor U9932 (N_9932,N_8666,N_8814);
xor U9933 (N_9933,N_8137,N_8315);
nor U9934 (N_9934,N_8842,N_7980);
nor U9935 (N_9935,N_8666,N_7732);
xnor U9936 (N_9936,N_8131,N_8098);
nand U9937 (N_9937,N_8223,N_8843);
nand U9938 (N_9938,N_8441,N_8752);
xor U9939 (N_9939,N_8204,N_7868);
and U9940 (N_9940,N_7793,N_7726);
nand U9941 (N_9941,N_7555,N_7696);
and U9942 (N_9942,N_8374,N_8705);
and U9943 (N_9943,N_8750,N_8887);
xor U9944 (N_9944,N_8187,N_8221);
nor U9945 (N_9945,N_7846,N_8989);
and U9946 (N_9946,N_8082,N_8727);
xnor U9947 (N_9947,N_8024,N_8637);
xnor U9948 (N_9948,N_8310,N_8025);
nor U9949 (N_9949,N_8047,N_8739);
nor U9950 (N_9950,N_8039,N_7889);
nor U9951 (N_9951,N_7737,N_8621);
nor U9952 (N_9952,N_7946,N_8046);
nand U9953 (N_9953,N_8230,N_7564);
or U9954 (N_9954,N_8911,N_8375);
or U9955 (N_9955,N_8617,N_7863);
or U9956 (N_9956,N_8002,N_8526);
xnor U9957 (N_9957,N_8515,N_8709);
xnor U9958 (N_9958,N_8590,N_8811);
or U9959 (N_9959,N_8992,N_7956);
xnor U9960 (N_9960,N_8270,N_8432);
nor U9961 (N_9961,N_7615,N_7796);
or U9962 (N_9962,N_7907,N_8408);
and U9963 (N_9963,N_8440,N_7663);
or U9964 (N_9964,N_7513,N_8627);
nand U9965 (N_9965,N_8766,N_8934);
nor U9966 (N_9966,N_8791,N_8977);
nor U9967 (N_9967,N_8555,N_7786);
xnor U9968 (N_9968,N_7871,N_8057);
nor U9969 (N_9969,N_7939,N_7953);
nor U9970 (N_9970,N_8287,N_8326);
nor U9971 (N_9971,N_8378,N_8433);
xor U9972 (N_9972,N_8236,N_8576);
nor U9973 (N_9973,N_7660,N_7922);
or U9974 (N_9974,N_8344,N_7606);
nand U9975 (N_9975,N_7930,N_7939);
nor U9976 (N_9976,N_8377,N_7658);
nor U9977 (N_9977,N_8467,N_8423);
or U9978 (N_9978,N_8862,N_8345);
or U9979 (N_9979,N_8604,N_8306);
xnor U9980 (N_9980,N_8316,N_8843);
xnor U9981 (N_9981,N_8170,N_8930);
xor U9982 (N_9982,N_7946,N_7928);
nor U9983 (N_9983,N_7636,N_8262);
nand U9984 (N_9984,N_8832,N_7678);
nand U9985 (N_9985,N_8388,N_8285);
nor U9986 (N_9986,N_8935,N_7989);
and U9987 (N_9987,N_7863,N_8917);
nand U9988 (N_9988,N_7681,N_7779);
nand U9989 (N_9989,N_7564,N_7727);
or U9990 (N_9990,N_8062,N_8381);
nand U9991 (N_9991,N_7843,N_7957);
and U9992 (N_9992,N_8369,N_8058);
nor U9993 (N_9993,N_8152,N_8448);
nor U9994 (N_9994,N_8469,N_7874);
nand U9995 (N_9995,N_8142,N_8517);
nand U9996 (N_9996,N_7649,N_8525);
nand U9997 (N_9997,N_8708,N_8827);
xnor U9998 (N_9998,N_8323,N_8495);
xnor U9999 (N_9999,N_7724,N_8151);
or U10000 (N_10000,N_8615,N_8023);
xnor U10001 (N_10001,N_8529,N_8684);
and U10002 (N_10002,N_7872,N_8542);
or U10003 (N_10003,N_8183,N_8964);
nor U10004 (N_10004,N_7863,N_7991);
nor U10005 (N_10005,N_7805,N_7575);
and U10006 (N_10006,N_8764,N_7960);
and U10007 (N_10007,N_8354,N_7879);
nand U10008 (N_10008,N_8898,N_8476);
nor U10009 (N_10009,N_7654,N_8294);
nand U10010 (N_10010,N_7521,N_8783);
nand U10011 (N_10011,N_8194,N_8273);
nand U10012 (N_10012,N_7515,N_8647);
nand U10013 (N_10013,N_7829,N_8694);
nand U10014 (N_10014,N_7506,N_8795);
and U10015 (N_10015,N_7808,N_7816);
nor U10016 (N_10016,N_8596,N_8299);
and U10017 (N_10017,N_8595,N_8058);
nand U10018 (N_10018,N_8332,N_7911);
xnor U10019 (N_10019,N_7861,N_7956);
nor U10020 (N_10020,N_8721,N_8525);
nand U10021 (N_10021,N_7776,N_7790);
or U10022 (N_10022,N_8323,N_8515);
and U10023 (N_10023,N_8112,N_8933);
nand U10024 (N_10024,N_8922,N_8758);
xnor U10025 (N_10025,N_8544,N_7505);
xnor U10026 (N_10026,N_7862,N_7572);
nor U10027 (N_10027,N_8004,N_7524);
and U10028 (N_10028,N_7682,N_7799);
and U10029 (N_10029,N_7722,N_7696);
nor U10030 (N_10030,N_8002,N_8753);
nand U10031 (N_10031,N_8701,N_7503);
and U10032 (N_10032,N_8676,N_8644);
nand U10033 (N_10033,N_8555,N_7523);
and U10034 (N_10034,N_7839,N_7723);
nor U10035 (N_10035,N_8177,N_8270);
xor U10036 (N_10036,N_8652,N_8808);
or U10037 (N_10037,N_8638,N_8427);
and U10038 (N_10038,N_8068,N_8493);
nor U10039 (N_10039,N_7849,N_8350);
and U10040 (N_10040,N_8137,N_8149);
or U10041 (N_10041,N_8474,N_8880);
nand U10042 (N_10042,N_8624,N_8595);
or U10043 (N_10043,N_8026,N_8483);
and U10044 (N_10044,N_8900,N_7532);
and U10045 (N_10045,N_8889,N_8477);
xor U10046 (N_10046,N_8893,N_8547);
or U10047 (N_10047,N_7875,N_8522);
nand U10048 (N_10048,N_7885,N_8326);
xnor U10049 (N_10049,N_7743,N_8949);
or U10050 (N_10050,N_7786,N_8883);
nor U10051 (N_10051,N_8254,N_7515);
or U10052 (N_10052,N_7658,N_7537);
xor U10053 (N_10053,N_8317,N_8708);
and U10054 (N_10054,N_8772,N_8638);
nor U10055 (N_10055,N_8155,N_7920);
nor U10056 (N_10056,N_8987,N_7832);
nand U10057 (N_10057,N_7714,N_8900);
and U10058 (N_10058,N_8056,N_8362);
and U10059 (N_10059,N_8548,N_8319);
nand U10060 (N_10060,N_8471,N_8984);
nand U10061 (N_10061,N_8180,N_8853);
or U10062 (N_10062,N_7731,N_8605);
xor U10063 (N_10063,N_7704,N_8922);
and U10064 (N_10064,N_8307,N_8545);
xor U10065 (N_10065,N_8714,N_7591);
nor U10066 (N_10066,N_8643,N_7908);
or U10067 (N_10067,N_7571,N_8502);
and U10068 (N_10068,N_8627,N_8866);
xor U10069 (N_10069,N_8765,N_8714);
xor U10070 (N_10070,N_8732,N_7779);
nand U10071 (N_10071,N_8239,N_7748);
xor U10072 (N_10072,N_8194,N_8816);
nand U10073 (N_10073,N_7860,N_8403);
nand U10074 (N_10074,N_8979,N_8307);
or U10075 (N_10075,N_8262,N_8471);
nor U10076 (N_10076,N_8192,N_8950);
or U10077 (N_10077,N_8524,N_8985);
nand U10078 (N_10078,N_7758,N_8581);
nor U10079 (N_10079,N_8707,N_7862);
xnor U10080 (N_10080,N_8427,N_8721);
xor U10081 (N_10081,N_8974,N_8429);
and U10082 (N_10082,N_7765,N_8787);
nand U10083 (N_10083,N_7935,N_8511);
xnor U10084 (N_10084,N_8120,N_7545);
nand U10085 (N_10085,N_7604,N_8488);
xor U10086 (N_10086,N_8263,N_8069);
or U10087 (N_10087,N_7696,N_7589);
xor U10088 (N_10088,N_8341,N_8004);
nor U10089 (N_10089,N_7765,N_7697);
nor U10090 (N_10090,N_7829,N_7848);
or U10091 (N_10091,N_7963,N_7599);
xor U10092 (N_10092,N_8110,N_7665);
nor U10093 (N_10093,N_8475,N_8051);
nor U10094 (N_10094,N_7889,N_8967);
nor U10095 (N_10095,N_8458,N_7873);
xor U10096 (N_10096,N_8659,N_7836);
nor U10097 (N_10097,N_8012,N_7822);
or U10098 (N_10098,N_8466,N_8915);
nand U10099 (N_10099,N_7753,N_8617);
nand U10100 (N_10100,N_7762,N_8997);
and U10101 (N_10101,N_8761,N_8702);
or U10102 (N_10102,N_8033,N_8456);
and U10103 (N_10103,N_7917,N_7569);
xnor U10104 (N_10104,N_8673,N_8360);
xnor U10105 (N_10105,N_7855,N_7646);
nand U10106 (N_10106,N_7744,N_8486);
or U10107 (N_10107,N_8290,N_7728);
nand U10108 (N_10108,N_8132,N_8067);
nand U10109 (N_10109,N_8335,N_7658);
nor U10110 (N_10110,N_8644,N_8080);
and U10111 (N_10111,N_8999,N_8475);
or U10112 (N_10112,N_8241,N_8051);
nand U10113 (N_10113,N_8919,N_7977);
or U10114 (N_10114,N_7970,N_7620);
xor U10115 (N_10115,N_7879,N_8722);
or U10116 (N_10116,N_7875,N_8816);
nand U10117 (N_10117,N_8941,N_7729);
xor U10118 (N_10118,N_8332,N_7557);
nand U10119 (N_10119,N_8175,N_7974);
nor U10120 (N_10120,N_8341,N_7915);
and U10121 (N_10121,N_7603,N_8362);
nor U10122 (N_10122,N_8508,N_8724);
xor U10123 (N_10123,N_7900,N_8584);
nand U10124 (N_10124,N_7726,N_8070);
and U10125 (N_10125,N_7790,N_8715);
nor U10126 (N_10126,N_8217,N_8196);
nand U10127 (N_10127,N_8672,N_8937);
and U10128 (N_10128,N_7634,N_7987);
nor U10129 (N_10129,N_8046,N_7927);
nand U10130 (N_10130,N_8344,N_7789);
and U10131 (N_10131,N_8034,N_8557);
and U10132 (N_10132,N_8203,N_7958);
nand U10133 (N_10133,N_8275,N_8012);
nor U10134 (N_10134,N_8175,N_7887);
or U10135 (N_10135,N_7891,N_7670);
nand U10136 (N_10136,N_8300,N_8694);
nor U10137 (N_10137,N_7957,N_7868);
or U10138 (N_10138,N_8319,N_8175);
nand U10139 (N_10139,N_8673,N_8825);
and U10140 (N_10140,N_8339,N_8617);
or U10141 (N_10141,N_7708,N_7802);
xnor U10142 (N_10142,N_8558,N_8779);
and U10143 (N_10143,N_8032,N_8797);
xor U10144 (N_10144,N_8919,N_8792);
xnor U10145 (N_10145,N_8478,N_8963);
nand U10146 (N_10146,N_8233,N_8738);
and U10147 (N_10147,N_7602,N_8468);
xor U10148 (N_10148,N_8801,N_8106);
nor U10149 (N_10149,N_8223,N_8784);
xor U10150 (N_10150,N_8643,N_8387);
xnor U10151 (N_10151,N_8608,N_7743);
and U10152 (N_10152,N_7564,N_7781);
or U10153 (N_10153,N_8241,N_7969);
or U10154 (N_10154,N_8338,N_7996);
xnor U10155 (N_10155,N_8894,N_7945);
nor U10156 (N_10156,N_8945,N_8824);
nand U10157 (N_10157,N_7618,N_7568);
and U10158 (N_10158,N_8853,N_8185);
and U10159 (N_10159,N_7659,N_7620);
or U10160 (N_10160,N_8265,N_8682);
and U10161 (N_10161,N_8914,N_7984);
nor U10162 (N_10162,N_8296,N_8945);
or U10163 (N_10163,N_8904,N_8386);
nor U10164 (N_10164,N_7954,N_8574);
or U10165 (N_10165,N_8792,N_7900);
xor U10166 (N_10166,N_8899,N_8295);
or U10167 (N_10167,N_8254,N_7696);
and U10168 (N_10168,N_7991,N_7738);
nor U10169 (N_10169,N_8264,N_7535);
and U10170 (N_10170,N_8959,N_7546);
xnor U10171 (N_10171,N_7968,N_8326);
and U10172 (N_10172,N_8344,N_8704);
xnor U10173 (N_10173,N_7717,N_8759);
nor U10174 (N_10174,N_7754,N_8786);
nor U10175 (N_10175,N_8789,N_8644);
nand U10176 (N_10176,N_8145,N_8937);
and U10177 (N_10177,N_8942,N_8078);
nand U10178 (N_10178,N_8192,N_7534);
and U10179 (N_10179,N_7551,N_7913);
nor U10180 (N_10180,N_8716,N_8573);
nor U10181 (N_10181,N_8895,N_8061);
or U10182 (N_10182,N_7906,N_8057);
nor U10183 (N_10183,N_8496,N_8642);
nand U10184 (N_10184,N_7870,N_8787);
nand U10185 (N_10185,N_8022,N_8393);
nor U10186 (N_10186,N_8372,N_8005);
nor U10187 (N_10187,N_8670,N_8567);
and U10188 (N_10188,N_7924,N_8222);
or U10189 (N_10189,N_7562,N_8677);
xnor U10190 (N_10190,N_8560,N_8266);
or U10191 (N_10191,N_8866,N_7598);
or U10192 (N_10192,N_7629,N_7627);
or U10193 (N_10193,N_7782,N_8374);
xor U10194 (N_10194,N_8757,N_8201);
nand U10195 (N_10195,N_8913,N_7524);
nand U10196 (N_10196,N_8968,N_8207);
xor U10197 (N_10197,N_8887,N_7947);
xor U10198 (N_10198,N_8198,N_8869);
and U10199 (N_10199,N_7910,N_8417);
nor U10200 (N_10200,N_8690,N_7718);
or U10201 (N_10201,N_8996,N_7973);
or U10202 (N_10202,N_8604,N_7573);
xor U10203 (N_10203,N_8716,N_8551);
nor U10204 (N_10204,N_8370,N_8463);
and U10205 (N_10205,N_8460,N_8651);
nor U10206 (N_10206,N_7533,N_7905);
and U10207 (N_10207,N_7860,N_8292);
xor U10208 (N_10208,N_8047,N_8461);
nor U10209 (N_10209,N_7517,N_8117);
or U10210 (N_10210,N_8726,N_8010);
or U10211 (N_10211,N_8027,N_8352);
nor U10212 (N_10212,N_8900,N_7863);
and U10213 (N_10213,N_8097,N_8631);
nand U10214 (N_10214,N_8121,N_8177);
and U10215 (N_10215,N_8638,N_8085);
nor U10216 (N_10216,N_7576,N_7983);
or U10217 (N_10217,N_8583,N_8274);
or U10218 (N_10218,N_7562,N_7622);
or U10219 (N_10219,N_8371,N_8516);
and U10220 (N_10220,N_7749,N_7981);
nor U10221 (N_10221,N_8591,N_7601);
nand U10222 (N_10222,N_8126,N_8380);
xor U10223 (N_10223,N_7602,N_7504);
or U10224 (N_10224,N_8466,N_7517);
nand U10225 (N_10225,N_8079,N_8946);
nand U10226 (N_10226,N_8967,N_8925);
nor U10227 (N_10227,N_8282,N_8945);
nand U10228 (N_10228,N_7806,N_8269);
nand U10229 (N_10229,N_8947,N_7542);
nand U10230 (N_10230,N_8010,N_7893);
nand U10231 (N_10231,N_8792,N_7830);
or U10232 (N_10232,N_8167,N_7606);
nand U10233 (N_10233,N_8089,N_8892);
or U10234 (N_10234,N_8190,N_7616);
xnor U10235 (N_10235,N_8343,N_7995);
xor U10236 (N_10236,N_8762,N_8497);
xnor U10237 (N_10237,N_8296,N_8899);
or U10238 (N_10238,N_8057,N_8050);
or U10239 (N_10239,N_8247,N_7783);
xnor U10240 (N_10240,N_8532,N_8410);
nor U10241 (N_10241,N_7615,N_7527);
xor U10242 (N_10242,N_8347,N_7929);
nor U10243 (N_10243,N_8799,N_8737);
xor U10244 (N_10244,N_8863,N_8247);
nor U10245 (N_10245,N_8964,N_8825);
and U10246 (N_10246,N_7703,N_7808);
xnor U10247 (N_10247,N_8510,N_7672);
and U10248 (N_10248,N_8006,N_7899);
nand U10249 (N_10249,N_8318,N_8190);
nor U10250 (N_10250,N_8279,N_8830);
or U10251 (N_10251,N_7723,N_8843);
xnor U10252 (N_10252,N_7581,N_7958);
and U10253 (N_10253,N_8263,N_8640);
xnor U10254 (N_10254,N_7648,N_7719);
nor U10255 (N_10255,N_8349,N_8123);
xor U10256 (N_10256,N_8038,N_8911);
xor U10257 (N_10257,N_7919,N_8058);
xor U10258 (N_10258,N_8621,N_8830);
nor U10259 (N_10259,N_8890,N_8841);
nor U10260 (N_10260,N_7829,N_8620);
nand U10261 (N_10261,N_8646,N_8413);
and U10262 (N_10262,N_7787,N_8525);
nand U10263 (N_10263,N_8409,N_8159);
nand U10264 (N_10264,N_7633,N_7533);
nor U10265 (N_10265,N_7915,N_8854);
nor U10266 (N_10266,N_8043,N_8982);
and U10267 (N_10267,N_8208,N_8364);
nor U10268 (N_10268,N_8306,N_8456);
nand U10269 (N_10269,N_7817,N_7891);
and U10270 (N_10270,N_8249,N_7826);
nor U10271 (N_10271,N_8545,N_7945);
and U10272 (N_10272,N_7901,N_8870);
or U10273 (N_10273,N_7816,N_8209);
nor U10274 (N_10274,N_8211,N_8265);
nand U10275 (N_10275,N_8207,N_8750);
nand U10276 (N_10276,N_7910,N_7644);
or U10277 (N_10277,N_7750,N_8352);
nor U10278 (N_10278,N_8292,N_7551);
nand U10279 (N_10279,N_8617,N_7870);
xnor U10280 (N_10280,N_8131,N_8528);
nor U10281 (N_10281,N_8208,N_8660);
or U10282 (N_10282,N_8235,N_8833);
nand U10283 (N_10283,N_8791,N_8937);
xor U10284 (N_10284,N_8052,N_8995);
nand U10285 (N_10285,N_8037,N_8890);
or U10286 (N_10286,N_8484,N_8622);
xor U10287 (N_10287,N_8734,N_8367);
and U10288 (N_10288,N_8226,N_7752);
nand U10289 (N_10289,N_8410,N_8909);
xnor U10290 (N_10290,N_8632,N_7994);
xor U10291 (N_10291,N_7989,N_8427);
nor U10292 (N_10292,N_8891,N_8069);
and U10293 (N_10293,N_8864,N_8286);
nand U10294 (N_10294,N_7899,N_8007);
or U10295 (N_10295,N_7681,N_8253);
xnor U10296 (N_10296,N_7861,N_8173);
or U10297 (N_10297,N_8497,N_8625);
nor U10298 (N_10298,N_8715,N_8829);
and U10299 (N_10299,N_8413,N_8777);
xnor U10300 (N_10300,N_8974,N_7758);
nand U10301 (N_10301,N_8870,N_8866);
or U10302 (N_10302,N_8167,N_8063);
nand U10303 (N_10303,N_8681,N_8902);
or U10304 (N_10304,N_7987,N_8857);
nand U10305 (N_10305,N_8395,N_8922);
and U10306 (N_10306,N_8340,N_8555);
and U10307 (N_10307,N_8169,N_8589);
xor U10308 (N_10308,N_8768,N_7558);
or U10309 (N_10309,N_8451,N_8221);
or U10310 (N_10310,N_8259,N_8728);
nand U10311 (N_10311,N_7854,N_8800);
nand U10312 (N_10312,N_8468,N_8494);
xor U10313 (N_10313,N_8719,N_8231);
nand U10314 (N_10314,N_8165,N_8010);
xor U10315 (N_10315,N_8229,N_7725);
nand U10316 (N_10316,N_8780,N_7816);
and U10317 (N_10317,N_8458,N_8054);
xor U10318 (N_10318,N_8377,N_8008);
nor U10319 (N_10319,N_7761,N_7555);
xnor U10320 (N_10320,N_7782,N_8302);
or U10321 (N_10321,N_7749,N_8941);
nor U10322 (N_10322,N_7915,N_8033);
nand U10323 (N_10323,N_8165,N_7907);
and U10324 (N_10324,N_8811,N_8947);
and U10325 (N_10325,N_7658,N_7614);
xor U10326 (N_10326,N_8463,N_8390);
nor U10327 (N_10327,N_7661,N_7514);
nand U10328 (N_10328,N_8302,N_8135);
and U10329 (N_10329,N_8891,N_7742);
nor U10330 (N_10330,N_8507,N_7558);
and U10331 (N_10331,N_8239,N_8638);
nand U10332 (N_10332,N_8990,N_8651);
or U10333 (N_10333,N_8296,N_8739);
and U10334 (N_10334,N_8859,N_8871);
nor U10335 (N_10335,N_7574,N_7640);
nand U10336 (N_10336,N_8661,N_8526);
and U10337 (N_10337,N_8525,N_8296);
xor U10338 (N_10338,N_7867,N_8271);
nand U10339 (N_10339,N_7827,N_8153);
nand U10340 (N_10340,N_8747,N_7540);
or U10341 (N_10341,N_8960,N_8217);
and U10342 (N_10342,N_8445,N_7614);
nor U10343 (N_10343,N_8528,N_8486);
nor U10344 (N_10344,N_7945,N_8929);
and U10345 (N_10345,N_7642,N_8630);
and U10346 (N_10346,N_8237,N_8391);
xor U10347 (N_10347,N_8931,N_8575);
nand U10348 (N_10348,N_7708,N_8504);
and U10349 (N_10349,N_8773,N_7998);
and U10350 (N_10350,N_8900,N_8764);
or U10351 (N_10351,N_7569,N_8875);
or U10352 (N_10352,N_8593,N_8644);
or U10353 (N_10353,N_8248,N_8581);
nand U10354 (N_10354,N_7502,N_7957);
nand U10355 (N_10355,N_8591,N_8968);
or U10356 (N_10356,N_8733,N_8148);
nand U10357 (N_10357,N_8263,N_8569);
or U10358 (N_10358,N_8859,N_8459);
and U10359 (N_10359,N_8718,N_8351);
xnor U10360 (N_10360,N_8158,N_7581);
or U10361 (N_10361,N_8176,N_8036);
nor U10362 (N_10362,N_7545,N_7749);
nor U10363 (N_10363,N_8717,N_7532);
nor U10364 (N_10364,N_7559,N_7836);
or U10365 (N_10365,N_8748,N_8411);
xnor U10366 (N_10366,N_7920,N_8818);
nor U10367 (N_10367,N_8789,N_8844);
nand U10368 (N_10368,N_8061,N_8065);
nand U10369 (N_10369,N_7892,N_7711);
and U10370 (N_10370,N_8444,N_8950);
or U10371 (N_10371,N_8208,N_8501);
nor U10372 (N_10372,N_8864,N_8803);
nand U10373 (N_10373,N_7532,N_8314);
nor U10374 (N_10374,N_8336,N_8574);
or U10375 (N_10375,N_8379,N_8176);
nor U10376 (N_10376,N_8243,N_7625);
nor U10377 (N_10377,N_7567,N_8618);
nand U10378 (N_10378,N_8285,N_8555);
nand U10379 (N_10379,N_8045,N_7608);
nor U10380 (N_10380,N_7831,N_7568);
nor U10381 (N_10381,N_8430,N_8592);
nor U10382 (N_10382,N_7804,N_8811);
and U10383 (N_10383,N_8980,N_8828);
and U10384 (N_10384,N_8588,N_8374);
xor U10385 (N_10385,N_7730,N_7963);
nand U10386 (N_10386,N_8515,N_8729);
xor U10387 (N_10387,N_8289,N_7914);
nand U10388 (N_10388,N_7922,N_7748);
nor U10389 (N_10389,N_8188,N_8628);
or U10390 (N_10390,N_8165,N_7506);
and U10391 (N_10391,N_7731,N_8815);
and U10392 (N_10392,N_8404,N_7536);
or U10393 (N_10393,N_7693,N_7573);
xnor U10394 (N_10394,N_8771,N_8345);
or U10395 (N_10395,N_8513,N_8159);
nor U10396 (N_10396,N_8173,N_8237);
xnor U10397 (N_10397,N_8594,N_7998);
nor U10398 (N_10398,N_7961,N_7829);
nor U10399 (N_10399,N_8222,N_8588);
nor U10400 (N_10400,N_8665,N_7904);
or U10401 (N_10401,N_8506,N_8001);
or U10402 (N_10402,N_7994,N_8262);
and U10403 (N_10403,N_8061,N_7896);
or U10404 (N_10404,N_8857,N_8561);
nand U10405 (N_10405,N_8559,N_7938);
nand U10406 (N_10406,N_7711,N_8338);
nand U10407 (N_10407,N_8678,N_8980);
xor U10408 (N_10408,N_7834,N_7770);
nor U10409 (N_10409,N_8626,N_8091);
nor U10410 (N_10410,N_8681,N_7960);
and U10411 (N_10411,N_7593,N_7517);
xor U10412 (N_10412,N_7852,N_7527);
xor U10413 (N_10413,N_7792,N_8536);
nor U10414 (N_10414,N_8758,N_7983);
nand U10415 (N_10415,N_8224,N_8893);
and U10416 (N_10416,N_8672,N_8842);
xor U10417 (N_10417,N_8665,N_7576);
or U10418 (N_10418,N_8763,N_8186);
or U10419 (N_10419,N_8987,N_7614);
xor U10420 (N_10420,N_7563,N_8444);
or U10421 (N_10421,N_7846,N_8515);
xor U10422 (N_10422,N_8580,N_8317);
xor U10423 (N_10423,N_8402,N_8019);
or U10424 (N_10424,N_7887,N_8121);
and U10425 (N_10425,N_8218,N_8098);
nand U10426 (N_10426,N_8075,N_8613);
and U10427 (N_10427,N_8261,N_7723);
xor U10428 (N_10428,N_8170,N_8660);
and U10429 (N_10429,N_8795,N_7609);
nor U10430 (N_10430,N_8663,N_7923);
nand U10431 (N_10431,N_7820,N_8194);
xor U10432 (N_10432,N_8042,N_8206);
nand U10433 (N_10433,N_8450,N_7760);
and U10434 (N_10434,N_8339,N_7808);
nand U10435 (N_10435,N_8546,N_8563);
xor U10436 (N_10436,N_7681,N_7740);
xnor U10437 (N_10437,N_8111,N_8597);
nand U10438 (N_10438,N_8406,N_8842);
or U10439 (N_10439,N_7766,N_8614);
or U10440 (N_10440,N_8606,N_8408);
nor U10441 (N_10441,N_8911,N_8305);
nand U10442 (N_10442,N_8861,N_7669);
nand U10443 (N_10443,N_8931,N_8219);
xnor U10444 (N_10444,N_8038,N_8369);
and U10445 (N_10445,N_7629,N_8899);
xnor U10446 (N_10446,N_7778,N_8254);
and U10447 (N_10447,N_8413,N_8662);
and U10448 (N_10448,N_8407,N_8654);
xnor U10449 (N_10449,N_8522,N_8466);
or U10450 (N_10450,N_7564,N_7690);
nor U10451 (N_10451,N_7904,N_8432);
xor U10452 (N_10452,N_8015,N_7863);
nand U10453 (N_10453,N_7990,N_8145);
or U10454 (N_10454,N_8210,N_8534);
nor U10455 (N_10455,N_8935,N_8894);
nor U10456 (N_10456,N_8701,N_7857);
nor U10457 (N_10457,N_7505,N_7657);
xnor U10458 (N_10458,N_7609,N_7703);
nand U10459 (N_10459,N_8685,N_8055);
nor U10460 (N_10460,N_7727,N_8205);
nand U10461 (N_10461,N_8942,N_8132);
xor U10462 (N_10462,N_8159,N_8657);
nand U10463 (N_10463,N_7803,N_8395);
xor U10464 (N_10464,N_8229,N_8004);
xor U10465 (N_10465,N_8082,N_7950);
and U10466 (N_10466,N_8113,N_8999);
nand U10467 (N_10467,N_7544,N_8158);
nand U10468 (N_10468,N_8638,N_8353);
and U10469 (N_10469,N_7542,N_8019);
xor U10470 (N_10470,N_8064,N_8916);
or U10471 (N_10471,N_7851,N_8415);
or U10472 (N_10472,N_8175,N_8129);
xor U10473 (N_10473,N_8716,N_8116);
nor U10474 (N_10474,N_8321,N_8895);
nand U10475 (N_10475,N_8812,N_7850);
xnor U10476 (N_10476,N_8529,N_7782);
and U10477 (N_10477,N_8920,N_7564);
nand U10478 (N_10478,N_7676,N_7914);
nor U10479 (N_10479,N_8810,N_8667);
nor U10480 (N_10480,N_8191,N_8274);
nor U10481 (N_10481,N_7794,N_8799);
or U10482 (N_10482,N_7973,N_8192);
and U10483 (N_10483,N_7825,N_8617);
and U10484 (N_10484,N_8213,N_8612);
or U10485 (N_10485,N_7633,N_7899);
xor U10486 (N_10486,N_8199,N_8670);
nor U10487 (N_10487,N_8002,N_7684);
or U10488 (N_10488,N_8807,N_8560);
and U10489 (N_10489,N_7801,N_7585);
nand U10490 (N_10490,N_7522,N_7843);
and U10491 (N_10491,N_8239,N_8498);
or U10492 (N_10492,N_7656,N_8806);
nor U10493 (N_10493,N_8425,N_8510);
or U10494 (N_10494,N_8535,N_8972);
or U10495 (N_10495,N_8014,N_7778);
or U10496 (N_10496,N_8698,N_8239);
or U10497 (N_10497,N_8478,N_8141);
nor U10498 (N_10498,N_7660,N_8235);
nor U10499 (N_10499,N_8663,N_8888);
or U10500 (N_10500,N_9441,N_9682);
xnor U10501 (N_10501,N_9364,N_10207);
and U10502 (N_10502,N_10034,N_9825);
and U10503 (N_10503,N_9181,N_9108);
xnor U10504 (N_10504,N_9871,N_10294);
xnor U10505 (N_10505,N_10360,N_9018);
nor U10506 (N_10506,N_9733,N_10496);
xor U10507 (N_10507,N_9227,N_10334);
or U10508 (N_10508,N_10464,N_9347);
nor U10509 (N_10509,N_10139,N_10470);
nand U10510 (N_10510,N_9664,N_9567);
xor U10511 (N_10511,N_9530,N_9829);
or U10512 (N_10512,N_9639,N_9184);
and U10513 (N_10513,N_9717,N_10367);
or U10514 (N_10514,N_10238,N_10119);
and U10515 (N_10515,N_9028,N_9286);
or U10516 (N_10516,N_9542,N_10146);
nand U10517 (N_10517,N_10155,N_9898);
nor U10518 (N_10518,N_10126,N_10276);
nor U10519 (N_10519,N_9578,N_9708);
nor U10520 (N_10520,N_10018,N_9575);
xnor U10521 (N_10521,N_9662,N_10184);
nand U10522 (N_10522,N_10359,N_10278);
and U10523 (N_10523,N_9237,N_10167);
and U10524 (N_10524,N_9372,N_10208);
xnor U10525 (N_10525,N_10280,N_9460);
nor U10526 (N_10526,N_9442,N_9055);
or U10527 (N_10527,N_9385,N_9369);
xor U10528 (N_10528,N_9930,N_9233);
nor U10529 (N_10529,N_10033,N_9454);
or U10530 (N_10530,N_10240,N_9983);
and U10531 (N_10531,N_10116,N_10447);
xor U10532 (N_10532,N_9675,N_10301);
nor U10533 (N_10533,N_9977,N_9179);
nand U10534 (N_10534,N_9386,N_10486);
nor U10535 (N_10535,N_9025,N_9073);
or U10536 (N_10536,N_10473,N_10308);
nand U10537 (N_10537,N_9243,N_10386);
nor U10538 (N_10538,N_9050,N_9075);
or U10539 (N_10539,N_10160,N_10071);
and U10540 (N_10540,N_9239,N_9023);
nor U10541 (N_10541,N_10299,N_9048);
nor U10542 (N_10542,N_9269,N_9312);
xnor U10543 (N_10543,N_10144,N_9396);
xnor U10544 (N_10544,N_9336,N_9543);
nor U10545 (N_10545,N_9861,N_10279);
or U10546 (N_10546,N_9362,N_10478);
xor U10547 (N_10547,N_9554,N_9735);
xor U10548 (N_10548,N_9823,N_9481);
nand U10549 (N_10549,N_9995,N_9081);
and U10550 (N_10550,N_9057,N_9666);
nor U10551 (N_10551,N_10021,N_10433);
xnor U10552 (N_10552,N_9982,N_9642);
and U10553 (N_10553,N_10472,N_10057);
or U10554 (N_10554,N_9934,N_10412);
nor U10555 (N_10555,N_9496,N_10451);
nand U10556 (N_10556,N_9840,N_10142);
xnor U10557 (N_10557,N_9146,N_9000);
or U10558 (N_10558,N_9244,N_10066);
nand U10559 (N_10559,N_9730,N_9812);
nand U10560 (N_10560,N_9749,N_9498);
and U10561 (N_10561,N_9775,N_10157);
xnor U10562 (N_10562,N_10419,N_9351);
and U10563 (N_10563,N_10064,N_9596);
or U10564 (N_10564,N_9923,N_9301);
xnor U10565 (N_10565,N_9358,N_9981);
xnor U10566 (N_10566,N_10312,N_9284);
nor U10567 (N_10567,N_9070,N_10340);
nand U10568 (N_10568,N_9217,N_9204);
and U10569 (N_10569,N_9990,N_9695);
and U10570 (N_10570,N_9796,N_9544);
or U10571 (N_10571,N_9563,N_9742);
or U10572 (N_10572,N_9870,N_10354);
or U10573 (N_10573,N_9319,N_9451);
xor U10574 (N_10574,N_10007,N_10277);
or U10575 (N_10575,N_9082,N_10151);
nor U10576 (N_10576,N_9446,N_9024);
or U10577 (N_10577,N_9201,N_10356);
nand U10578 (N_10578,N_9277,N_9449);
and U10579 (N_10579,N_10328,N_9719);
xnor U10580 (N_10580,N_9497,N_10118);
or U10581 (N_10581,N_10471,N_10036);
or U10582 (N_10582,N_9091,N_10317);
or U10583 (N_10583,N_9998,N_10257);
nor U10584 (N_10584,N_9152,N_9132);
xnor U10585 (N_10585,N_10095,N_9445);
nor U10586 (N_10586,N_9458,N_9888);
nor U10587 (N_10587,N_9086,N_9387);
or U10588 (N_10588,N_9189,N_9072);
nor U10589 (N_10589,N_9869,N_9203);
xor U10590 (N_10590,N_10313,N_9683);
xnor U10591 (N_10591,N_10015,N_9709);
nor U10592 (N_10592,N_9125,N_9685);
xor U10593 (N_10593,N_10044,N_10474);
nor U10594 (N_10594,N_9536,N_10408);
nor U10595 (N_10595,N_9142,N_10050);
xor U10596 (N_10596,N_10008,N_9216);
nor U10597 (N_10597,N_9459,N_10004);
nand U10598 (N_10598,N_10324,N_9684);
nor U10599 (N_10599,N_9550,N_9852);
or U10600 (N_10600,N_9855,N_9097);
nand U10601 (N_10601,N_9897,N_9137);
and U10602 (N_10602,N_9979,N_9880);
and U10603 (N_10603,N_9323,N_9994);
or U10604 (N_10604,N_10389,N_9223);
or U10605 (N_10605,N_9180,N_9595);
nor U10606 (N_10606,N_9404,N_9661);
or U10607 (N_10607,N_9699,N_10053);
nand U10608 (N_10608,N_10088,N_9740);
nand U10609 (N_10609,N_9365,N_9085);
nand U10610 (N_10610,N_10251,N_9159);
nand U10611 (N_10611,N_10176,N_9980);
nor U10612 (N_10612,N_9197,N_9262);
and U10613 (N_10613,N_9927,N_10393);
xor U10614 (N_10614,N_9105,N_9267);
nor U10615 (N_10615,N_9326,N_9946);
and U10616 (N_10616,N_9864,N_9242);
nor U10617 (N_10617,N_9917,N_9997);
nand U10618 (N_10618,N_9436,N_9729);
and U10619 (N_10619,N_9030,N_10350);
or U10620 (N_10620,N_10010,N_9160);
xnor U10621 (N_10621,N_9753,N_9517);
nand U10622 (N_10622,N_10259,N_9153);
nor U10623 (N_10623,N_9261,N_9360);
and U10624 (N_10624,N_9592,N_9701);
or U10625 (N_10625,N_10410,N_9437);
nor U10626 (N_10626,N_10481,N_10012);
nor U10627 (N_10627,N_10329,N_9165);
nand U10628 (N_10628,N_9193,N_10398);
xor U10629 (N_10629,N_10256,N_9989);
xnor U10630 (N_10630,N_10222,N_9036);
xnor U10631 (N_10631,N_9453,N_10456);
nor U10632 (N_10632,N_9007,N_9327);
and U10633 (N_10633,N_9939,N_10365);
xnor U10634 (N_10634,N_9565,N_9743);
xnor U10635 (N_10635,N_10423,N_9035);
or U10636 (N_10636,N_9405,N_10242);
nor U10637 (N_10637,N_9349,N_10352);
xnor U10638 (N_10638,N_10479,N_9883);
or U10639 (N_10639,N_9031,N_10031);
nor U10640 (N_10640,N_9508,N_10055);
and U10641 (N_10641,N_9417,N_9282);
or U10642 (N_10642,N_10411,N_9915);
and U10643 (N_10643,N_9961,N_9813);
nand U10644 (N_10644,N_10099,N_9808);
or U10645 (N_10645,N_9366,N_10183);
nand U10646 (N_10646,N_9773,N_9856);
nor U10647 (N_10647,N_9175,N_10452);
or U10648 (N_10648,N_9100,N_9561);
and U10649 (N_10649,N_10404,N_10136);
xnor U10650 (N_10650,N_10081,N_9901);
or U10651 (N_10651,N_9389,N_9300);
nand U10652 (N_10652,N_10403,N_9718);
xor U10653 (N_10653,N_9558,N_9359);
nand U10654 (N_10654,N_10069,N_9688);
nor U10655 (N_10655,N_9291,N_10090);
nand U10656 (N_10656,N_9345,N_10191);
nor U10657 (N_10657,N_10011,N_9363);
and U10658 (N_10658,N_9290,N_9134);
nor U10659 (N_10659,N_9511,N_9002);
or U10660 (N_10660,N_10093,N_9967);
xnor U10661 (N_10661,N_9576,N_9435);
nor U10662 (N_10662,N_9212,N_9406);
or U10663 (N_10663,N_9245,N_10371);
and U10664 (N_10664,N_9609,N_9158);
nand U10665 (N_10665,N_10065,N_9540);
and U10666 (N_10666,N_9618,N_10429);
and U10667 (N_10667,N_10235,N_9084);
nand U10668 (N_10668,N_9214,N_10373);
and U10669 (N_10669,N_9518,N_9588);
and U10670 (N_10670,N_9568,N_9424);
and U10671 (N_10671,N_9838,N_9750);
nor U10672 (N_10672,N_9440,N_10296);
and U10673 (N_10673,N_9724,N_9426);
or U10674 (N_10674,N_9628,N_9804);
or U10675 (N_10675,N_9381,N_9090);
or U10676 (N_10676,N_9012,N_9623);
and U10677 (N_10677,N_10427,N_10111);
or U10678 (N_10678,N_9881,N_9877);
or U10679 (N_10679,N_9526,N_10122);
or U10680 (N_10680,N_10458,N_9538);
nand U10681 (N_10681,N_10453,N_9114);
or U10682 (N_10682,N_10089,N_10232);
nor U10683 (N_10683,N_9492,N_9782);
and U10684 (N_10684,N_9288,N_9604);
nand U10685 (N_10685,N_9375,N_9572);
and U10686 (N_10686,N_9110,N_9106);
or U10687 (N_10687,N_10422,N_9045);
nor U10688 (N_10688,N_9064,N_9976);
nand U10689 (N_10689,N_9455,N_10103);
or U10690 (N_10690,N_9135,N_9991);
and U10691 (N_10691,N_9253,N_9936);
xor U10692 (N_10692,N_9850,N_9325);
xnor U10693 (N_10693,N_9736,N_9827);
xor U10694 (N_10694,N_10000,N_10344);
xnor U10695 (N_10695,N_10109,N_10148);
or U10696 (N_10696,N_9419,N_9725);
or U10697 (N_10697,N_9894,N_9238);
nand U10698 (N_10698,N_10337,N_9702);
nor U10699 (N_10699,N_10275,N_10450);
nand U10700 (N_10700,N_10227,N_9904);
or U10701 (N_10701,N_9208,N_10417);
and U10702 (N_10702,N_9001,N_9505);
nor U10703 (N_10703,N_9858,N_10060);
nand U10704 (N_10704,N_9433,N_9042);
or U10705 (N_10705,N_9545,N_9241);
nand U10706 (N_10706,N_9960,N_10061);
and U10707 (N_10707,N_9298,N_9760);
or U10708 (N_10708,N_10223,N_10325);
xor U10709 (N_10709,N_9629,N_10180);
and U10710 (N_10710,N_10288,N_9694);
nor U10711 (N_10711,N_9232,N_10127);
and U10712 (N_10712,N_10174,N_9130);
or U10713 (N_10713,N_9196,N_9633);
or U10714 (N_10714,N_10432,N_10005);
xor U10715 (N_10715,N_9602,N_9993);
or U10716 (N_10716,N_9950,N_10305);
nand U10717 (N_10717,N_9186,N_9015);
and U10718 (N_10718,N_10224,N_10405);
nand U10719 (N_10719,N_10149,N_10290);
nand U10720 (N_10720,N_10024,N_9485);
or U10721 (N_10721,N_9964,N_9150);
nor U10722 (N_10722,N_9329,N_9867);
and U10723 (N_10723,N_9169,N_9706);
nor U10724 (N_10724,N_9376,N_10152);
xnor U10725 (N_10725,N_10048,N_10385);
nand U10726 (N_10726,N_9903,N_10041);
nor U10727 (N_10727,N_9620,N_10233);
or U10728 (N_10728,N_10264,N_9109);
nor U10729 (N_10729,N_10039,N_9972);
and U10730 (N_10730,N_10273,N_10497);
xnor U10731 (N_10731,N_9553,N_10120);
nand U10732 (N_10732,N_9911,N_9136);
xnor U10733 (N_10733,N_9907,N_9800);
xnor U10734 (N_10734,N_9818,N_9373);
nand U10735 (N_10735,N_9198,N_10335);
nor U10736 (N_10736,N_10209,N_9819);
nor U10737 (N_10737,N_9589,N_9305);
xnor U10738 (N_10738,N_10347,N_10401);
xnor U10739 (N_10739,N_9056,N_9738);
xnor U10740 (N_10740,N_10387,N_9182);
or U10741 (N_10741,N_10019,N_9403);
or U10742 (N_10742,N_10032,N_10345);
nand U10743 (N_10743,N_10017,N_9258);
or U10744 (N_10744,N_10049,N_10212);
nor U10745 (N_10745,N_9029,N_9330);
or U10746 (N_10746,N_10391,N_9127);
nor U10747 (N_10747,N_9734,N_9956);
nand U10748 (N_10748,N_9676,N_10321);
xor U10749 (N_10749,N_9693,N_9848);
xor U10750 (N_10750,N_10006,N_10316);
nor U10751 (N_10751,N_10098,N_9077);
xor U10752 (N_10752,N_10020,N_10075);
and U10753 (N_10753,N_9014,N_9475);
nand U10754 (N_10754,N_10203,N_9479);
and U10755 (N_10755,N_10446,N_9026);
nand U10756 (N_10756,N_10477,N_9790);
nor U10757 (N_10757,N_9546,N_9006);
nor U10758 (N_10758,N_10409,N_9107);
nand U10759 (N_10759,N_9087,N_9889);
nor U10760 (N_10760,N_9247,N_9846);
nand U10761 (N_10761,N_9102,N_10488);
or U10762 (N_10762,N_10141,N_10097);
nor U10763 (N_10763,N_9969,N_10192);
and U10764 (N_10764,N_10382,N_10361);
and U10765 (N_10765,N_9635,N_10366);
and U10766 (N_10766,N_10112,N_10295);
or U10767 (N_10767,N_9696,N_9332);
and U10768 (N_10768,N_9401,N_10326);
nor U10769 (N_10769,N_10133,N_10186);
nor U10770 (N_10770,N_9645,N_9421);
nand U10771 (N_10771,N_9624,N_10476);
xor U10772 (N_10772,N_9402,N_9866);
xnor U10773 (N_10773,N_9874,N_10003);
and U10774 (N_10774,N_9133,N_9534);
xor U10775 (N_10775,N_9593,N_10171);
or U10776 (N_10776,N_9672,N_9474);
and U10777 (N_10777,N_9557,N_10498);
xnor U10778 (N_10778,N_9266,N_10253);
nand U10779 (N_10779,N_9104,N_10388);
nor U10780 (N_10780,N_9817,N_9868);
or U10781 (N_10781,N_9257,N_9383);
and U10782 (N_10782,N_10138,N_10384);
xnor U10783 (N_10783,N_9937,N_9842);
xnor U10784 (N_10784,N_10378,N_10267);
xnor U10785 (N_10785,N_9962,N_9586);
or U10786 (N_10786,N_9251,N_9884);
and U10787 (N_10787,N_9154,N_10073);
and U10788 (N_10788,N_9340,N_9723);
nand U10789 (N_10789,N_9078,N_9703);
or U10790 (N_10790,N_9507,N_9318);
and U10791 (N_10791,N_9849,N_10218);
or U10792 (N_10792,N_9556,N_9625);
or U10793 (N_10793,N_10158,N_9971);
or U10794 (N_10794,N_9627,N_9632);
and U10795 (N_10795,N_9611,N_10038);
or U10796 (N_10796,N_9535,N_9339);
nor U10797 (N_10797,N_10499,N_10495);
or U10798 (N_10798,N_10485,N_10414);
and U10799 (N_10799,N_9034,N_9791);
nor U10800 (N_10800,N_9958,N_10102);
nand U10801 (N_10801,N_9178,N_9764);
and U10802 (N_10802,N_10219,N_9619);
nand U10803 (N_10803,N_9605,N_10241);
nand U10804 (N_10804,N_9249,N_10254);
xnor U10805 (N_10805,N_9830,N_10087);
or U10806 (N_10806,N_9415,N_9529);
or U10807 (N_10807,N_9882,N_9940);
nor U10808 (N_10808,N_9959,N_9533);
nor U10809 (N_10809,N_9295,N_10121);
and U10810 (N_10810,N_9255,N_10247);
and U10811 (N_10811,N_10465,N_9681);
xnor U10812 (N_10812,N_9429,N_9952);
or U10813 (N_10813,N_9431,N_10179);
nand U10814 (N_10814,N_9698,N_9103);
or U10815 (N_10815,N_9192,N_9126);
and U10816 (N_10816,N_9809,N_9095);
xor U10817 (N_10817,N_9833,N_9646);
nand U10818 (N_10818,N_9276,N_9795);
xor U10819 (N_10819,N_9256,N_9659);
and U10820 (N_10820,N_10062,N_10287);
xor U10821 (N_10821,N_9263,N_9836);
or U10822 (N_10822,N_9462,N_9674);
nor U10823 (N_10823,N_9384,N_9129);
or U10824 (N_10824,N_9900,N_9422);
xnor U10825 (N_10825,N_10231,N_10094);
nand U10826 (N_10826,N_10194,N_10370);
nor U10827 (N_10827,N_9640,N_9467);
nand U10828 (N_10828,N_10270,N_9948);
or U10829 (N_10829,N_10113,N_10096);
nand U10830 (N_10830,N_10128,N_10397);
xnor U10831 (N_10831,N_10394,N_9116);
and U10832 (N_10832,N_9516,N_9287);
nand U10833 (N_10833,N_10077,N_9494);
nand U10834 (N_10834,N_9834,N_9504);
or U10835 (N_10835,N_9613,N_9626);
and U10836 (N_10836,N_9941,N_9778);
nand U10837 (N_10837,N_10195,N_9416);
xnor U10838 (N_10838,N_10318,N_10029);
nand U10839 (N_10839,N_9054,N_9427);
nand U10840 (N_10840,N_9076,N_9194);
or U10841 (N_10841,N_9788,N_9476);
nor U10842 (N_10842,N_9471,N_9713);
xnor U10843 (N_10843,N_10289,N_10407);
and U10844 (N_10844,N_10045,N_10236);
xor U10845 (N_10845,N_9720,N_9811);
xnor U10846 (N_10846,N_10444,N_9068);
or U10847 (N_10847,N_9726,N_9739);
or U10848 (N_10848,N_9637,N_10091);
and U10849 (N_10849,N_9487,N_9928);
nor U10850 (N_10850,N_10368,N_9816);
or U10851 (N_10851,N_9118,N_9831);
nand U10852 (N_10852,N_10042,N_10322);
nand U10853 (N_10853,N_9652,N_9004);
or U10854 (N_10854,N_9879,N_9168);
nor U10855 (N_10855,N_9308,N_10467);
nand U10856 (N_10856,N_9918,N_9310);
nand U10857 (N_10857,N_9591,N_9786);
nand U10858 (N_10858,N_10415,N_10362);
nand U10859 (N_10859,N_9224,N_9616);
or U10860 (N_10860,N_10177,N_10210);
nand U10861 (N_10861,N_9038,N_9878);
xor U10862 (N_10862,N_9537,N_9931);
and U10863 (N_10863,N_10436,N_9667);
and U10864 (N_10864,N_10035,N_9443);
xor U10865 (N_10865,N_9355,N_9438);
or U10866 (N_10866,N_10249,N_9274);
nor U10867 (N_10867,N_9549,N_10163);
nor U10868 (N_10868,N_9027,N_9480);
nor U10869 (N_10869,N_9752,N_9228);
xnor U10870 (N_10870,N_9264,N_9121);
xnor U10871 (N_10871,N_9170,N_9722);
and U10872 (N_10872,N_9945,N_9774);
nand U10873 (N_10873,N_9714,N_9891);
nand U10874 (N_10874,N_9354,N_9032);
xnor U10875 (N_10875,N_9606,N_9910);
xor U10876 (N_10876,N_10245,N_9469);
nand U10877 (N_10877,N_9630,N_9280);
nor U10878 (N_10878,N_9377,N_9985);
and U10879 (N_10879,N_9079,N_9317);
xor U10880 (N_10880,N_9638,N_9074);
and U10881 (N_10881,N_10100,N_10114);
xor U10882 (N_10882,N_10416,N_9984);
and U10883 (N_10883,N_9872,N_10395);
xnor U10884 (N_10884,N_10248,N_10108);
or U10885 (N_10885,N_9017,N_10330);
and U10886 (N_10886,N_9221,N_10379);
nand U10887 (N_10887,N_10030,N_10262);
and U10888 (N_10888,N_10107,N_9019);
or U10889 (N_10889,N_10482,N_9527);
or U10890 (N_10890,N_9122,N_9350);
and U10891 (N_10891,N_10229,N_9607);
xor U10892 (N_10892,N_9250,N_10320);
or U10893 (N_10893,N_9677,N_9391);
or U10894 (N_10894,N_9631,N_9758);
xnor U10895 (N_10895,N_9761,N_9902);
and U10896 (N_10896,N_10263,N_10376);
xnor U10897 (N_10897,N_9559,N_9409);
nor U10898 (N_10898,N_9689,N_10123);
nor U10899 (N_10899,N_10197,N_10341);
nand U10900 (N_10900,N_9908,N_9707);
or U10901 (N_10901,N_9678,N_9515);
or U10902 (N_10902,N_9430,N_9851);
nand U10903 (N_10903,N_9215,N_9320);
xnor U10904 (N_10904,N_10413,N_9805);
xnor U10905 (N_10905,N_9065,N_10383);
and U10906 (N_10906,N_10309,N_9975);
or U10907 (N_10907,N_9914,N_10175);
and U10908 (N_10908,N_10092,N_9727);
nor U10909 (N_10909,N_9651,N_9163);
nand U10910 (N_10910,N_9577,N_10492);
or U10911 (N_10911,N_10441,N_9873);
nor U10912 (N_10912,N_9293,N_9314);
or U10913 (N_10913,N_9951,N_9597);
and U10914 (N_10914,N_10085,N_9828);
nor U10915 (N_10915,N_9783,N_10201);
xnor U10916 (N_10916,N_9574,N_10292);
or U10917 (N_10917,N_9803,N_9357);
nor U10918 (N_10918,N_10469,N_10137);
xor U10919 (N_10919,N_9202,N_10147);
and U10920 (N_10920,N_10353,N_10214);
nand U10921 (N_10921,N_9794,N_10002);
xnor U10922 (N_10922,N_10494,N_9745);
xor U10923 (N_10923,N_9139,N_10156);
nand U10924 (N_10924,N_9715,N_9209);
xor U10925 (N_10925,N_9470,N_9590);
nor U10926 (N_10926,N_9751,N_9539);
nand U10927 (N_10927,N_9041,N_9776);
or U10928 (N_10928,N_10272,N_9005);
or U10929 (N_10929,N_9060,N_10230);
nor U10930 (N_10930,N_10418,N_9650);
and U10931 (N_10931,N_9226,N_9514);
and U10932 (N_10932,N_10153,N_9283);
xor U10933 (N_10933,N_9862,N_9395);
and U10934 (N_10934,N_9408,N_9051);
nand U10935 (N_10935,N_9352,N_10129);
and U10936 (N_10936,N_9254,N_9929);
or U10937 (N_10937,N_10009,N_10493);
and U10938 (N_10938,N_9564,N_9987);
xor U10939 (N_10939,N_9599,N_9039);
xor U10940 (N_10940,N_9338,N_9731);
xnor U10941 (N_10941,N_9414,N_9865);
and U10942 (N_10942,N_10487,N_10342);
xor U10943 (N_10943,N_10438,N_9140);
or U10944 (N_10944,N_9093,N_9482);
xnor U10945 (N_10945,N_9965,N_10078);
nand U10946 (N_10946,N_9353,N_9787);
and U10947 (N_10947,N_9802,N_9665);
nand U10948 (N_10948,N_10076,N_9887);
xnor U10949 (N_10949,N_9762,N_10448);
and U10950 (N_10950,N_9143,N_10348);
xnor U10951 (N_10951,N_9847,N_10058);
or U10952 (N_10952,N_9636,N_9067);
or U10953 (N_10953,N_9769,N_10014);
and U10954 (N_10954,N_9814,N_10351);
nor U10955 (N_10955,N_9328,N_9399);
xor U10956 (N_10956,N_9615,N_9617);
xor U10957 (N_10957,N_9303,N_9712);
nor U10958 (N_10958,N_10110,N_9839);
xor U10959 (N_10959,N_9837,N_10323);
nor U10960 (N_10960,N_10311,N_10130);
xor U10961 (N_10961,N_9099,N_10182);
nor U10962 (N_10962,N_9423,N_9147);
nand U10963 (N_10963,N_9657,N_9071);
or U10964 (N_10964,N_10215,N_9785);
xnor U10965 (N_10965,N_10285,N_9123);
nand U10966 (N_10966,N_10284,N_10258);
or U10967 (N_10967,N_10083,N_9926);
nand U10968 (N_10968,N_9367,N_9489);
nor U10969 (N_10969,N_10402,N_9111);
nand U10970 (N_10970,N_10023,N_9306);
nand U10971 (N_10971,N_9439,N_10016);
and U10972 (N_10972,N_9601,N_9230);
and U10973 (N_10973,N_10300,N_9716);
and U10974 (N_10974,N_9020,N_9955);
nand U10975 (N_10975,N_10293,N_10054);
nor U10976 (N_10976,N_9711,N_10390);
nor U10977 (N_10977,N_9273,N_9053);
nand U10978 (N_10978,N_9176,N_10443);
nor U10979 (N_10979,N_10134,N_9647);
or U10980 (N_10980,N_9016,N_10420);
and U10981 (N_10981,N_9863,N_10483);
or U10982 (N_10982,N_9010,N_9634);
and U10983 (N_10983,N_9875,N_9853);
and U10984 (N_10984,N_9525,N_10178);
nand U10985 (N_10985,N_9022,N_10297);
nor U10986 (N_10986,N_9011,N_10043);
or U10987 (N_10987,N_9660,N_9473);
and U10988 (N_10988,N_9893,N_10237);
or U10989 (N_10989,N_9673,N_10462);
xnor U10990 (N_10990,N_9046,N_9268);
and U10991 (N_10991,N_9968,N_9947);
xor U10992 (N_10992,N_9779,N_9420);
xnor U10993 (N_10993,N_9755,N_9648);
and U10994 (N_10994,N_10169,N_9608);
and U10995 (N_10995,N_10125,N_10339);
or U10996 (N_10996,N_9149,N_9252);
or U10997 (N_10997,N_10421,N_9299);
nand U10998 (N_10998,N_10220,N_9583);
nand U10999 (N_10999,N_9801,N_9754);
xnor U11000 (N_11000,N_10181,N_9141);
and U11001 (N_11001,N_10302,N_9896);
nor U11002 (N_11002,N_9279,N_9380);
nand U11003 (N_11003,N_9271,N_9986);
nand U11004 (N_11004,N_9653,N_9052);
nand U11005 (N_11005,N_9999,N_9656);
or U11006 (N_11006,N_10027,N_9260);
nand U11007 (N_11007,N_10455,N_9040);
xor U11008 (N_11008,N_9766,N_10440);
xnor U11009 (N_11009,N_10435,N_10298);
nor U11010 (N_11010,N_10271,N_10228);
nor U11011 (N_11011,N_9157,N_9521);
nor U11012 (N_11012,N_9502,N_9705);
xnor U11013 (N_11013,N_9500,N_9285);
nor U11014 (N_11014,N_9321,N_9343);
and U11015 (N_11015,N_10143,N_9043);
or U11016 (N_11016,N_9037,N_10079);
nor U11017 (N_11017,N_10185,N_9499);
xor U11018 (N_11018,N_10468,N_9322);
and U11019 (N_11019,N_10068,N_10307);
and U11020 (N_11020,N_9164,N_10131);
or U11021 (N_11021,N_10430,N_10046);
xor U11022 (N_11022,N_10154,N_10283);
nand U11023 (N_11023,N_10439,N_9465);
xnor U11024 (N_11024,N_9996,N_9822);
xor U11025 (N_11025,N_9680,N_9275);
xor U11026 (N_11026,N_9205,N_10234);
and U11027 (N_11027,N_10211,N_9428);
xnor U11028 (N_11028,N_9368,N_9658);
nor U11029 (N_11029,N_9806,N_9155);
nand U11030 (N_11030,N_10115,N_9207);
xnor U11031 (N_11031,N_10445,N_9770);
nand U11032 (N_11032,N_9522,N_9235);
or U11033 (N_11033,N_9161,N_9225);
xor U11034 (N_11034,N_10037,N_9069);
or U11035 (N_11035,N_9117,N_10052);
nand U11036 (N_11036,N_9570,N_9407);
nand U11037 (N_11037,N_9501,N_9784);
xor U11038 (N_11038,N_9876,N_9344);
nor U11039 (N_11039,N_10056,N_10327);
nor U11040 (N_11040,N_9710,N_9957);
or U11041 (N_11041,N_10150,N_9144);
and U11042 (N_11042,N_9236,N_10086);
nand U11043 (N_11043,N_9062,N_9388);
nand U11044 (N_11044,N_10243,N_9096);
xor U11045 (N_11045,N_9191,N_9584);
or U11046 (N_11046,N_9581,N_10187);
nand U11047 (N_11047,N_9924,N_10104);
xor U11048 (N_11048,N_9411,N_9119);
and U11049 (N_11049,N_10490,N_10489);
nand U11050 (N_11050,N_10442,N_9490);
nor U11051 (N_11051,N_9768,N_9131);
or U11052 (N_11052,N_9434,N_10454);
xnor U11053 (N_11053,N_9356,N_9331);
or U11054 (N_11054,N_9992,N_9748);
nor U11055 (N_11055,N_9145,N_9187);
xor U11056 (N_11056,N_10193,N_9183);
or U11057 (N_11057,N_10315,N_9488);
and U11058 (N_11058,N_10170,N_9741);
xnor U11059 (N_11059,N_10434,N_9483);
nand U11060 (N_11060,N_9560,N_10372);
or U11061 (N_11061,N_10332,N_9777);
xor U11062 (N_11062,N_9151,N_9452);
and U11063 (N_11063,N_9461,N_9337);
and U11064 (N_11064,N_9859,N_9598);
and U11065 (N_11065,N_9447,N_9857);
nand U11066 (N_11066,N_9270,N_9824);
or U11067 (N_11067,N_9562,N_10199);
xor U11068 (N_11068,N_9418,N_9641);
xnor U11069 (N_11069,N_9477,N_9974);
and U11070 (N_11070,N_9379,N_10225);
xor U11071 (N_11071,N_9512,N_9912);
nor U11072 (N_11072,N_10173,N_10082);
or U11073 (N_11073,N_9013,N_9913);
nand U11074 (N_11074,N_9890,N_9061);
nand U11075 (N_11075,N_10291,N_9670);
or U11076 (N_11076,N_9763,N_9219);
nand U11077 (N_11077,N_10304,N_10059);
xnor U11078 (N_11078,N_10190,N_9361);
nand U11079 (N_11079,N_9767,N_9493);
nor U11080 (N_11080,N_9789,N_10025);
or U11081 (N_11081,N_10425,N_9679);
xnor U11082 (N_11082,N_9425,N_9370);
or U11083 (N_11083,N_10047,N_9311);
nor U11084 (N_11084,N_9094,N_9844);
nand U11085 (N_11085,N_9519,N_9200);
nor U11086 (N_11086,N_10466,N_10268);
and U11087 (N_11087,N_10162,N_10449);
or U11088 (N_11088,N_9098,N_9621);
nand U11089 (N_11089,N_10377,N_9973);
or U11090 (N_11090,N_9663,N_10484);
or U11091 (N_11091,N_9885,N_10303);
or U11092 (N_11092,N_9138,N_9622);
xor U11093 (N_11093,N_9832,N_9188);
xnor U11094 (N_11094,N_9008,N_9668);
nand U11095 (N_11095,N_9495,N_9304);
and U11096 (N_11096,N_9772,N_9324);
nor U11097 (N_11097,N_9394,N_9464);
xnor U11098 (N_11098,N_9393,N_9757);
and U11099 (N_11099,N_9371,N_10261);
and U11100 (N_11100,N_10204,N_9297);
and U11101 (N_11101,N_10196,N_10072);
nand U11102 (N_11102,N_9307,N_9174);
nor U11103 (N_11103,N_9821,N_10437);
xnor U11104 (N_11104,N_9547,N_10269);
nor U11105 (N_11105,N_9551,N_9700);
nor U11106 (N_11106,N_10067,N_9166);
nand U11107 (N_11107,N_10117,N_9569);
or U11108 (N_11108,N_9088,N_10244);
or U11109 (N_11109,N_10265,N_10260);
nand U11110 (N_11110,N_10428,N_9506);
and U11111 (N_11111,N_9744,N_10198);
or U11112 (N_11112,N_10381,N_10349);
xor U11113 (N_11113,N_10135,N_9835);
and U11114 (N_11114,N_10431,N_9692);
nand U11115 (N_11115,N_9222,N_9296);
xnor U11116 (N_11116,N_9966,N_10172);
or U11117 (N_11117,N_9797,N_10246);
nand U11118 (N_11118,N_9765,N_9737);
and U11119 (N_11119,N_9649,N_9644);
or U11120 (N_11120,N_9206,N_9571);
nand U11121 (N_11121,N_9240,N_9503);
xor U11122 (N_11122,N_9704,N_9112);
nor U11123 (N_11123,N_10028,N_9059);
or U11124 (N_11124,N_9410,N_10338);
xor U11125 (N_11125,N_9728,N_9793);
nor U11126 (N_11126,N_10255,N_10363);
xor U11127 (N_11127,N_9115,N_9643);
or U11128 (N_11128,N_10206,N_9397);
and U11129 (N_11129,N_10188,N_9400);
or U11130 (N_11130,N_9248,N_9080);
nand U11131 (N_11131,N_9899,N_9342);
or U11132 (N_11132,N_9063,N_9162);
or U11133 (N_11133,N_9472,N_9199);
or U11134 (N_11134,N_10314,N_9654);
nand U11135 (N_11135,N_10266,N_10202);
and U11136 (N_11136,N_9582,N_9392);
nor U11137 (N_11137,N_9292,N_9346);
or U11138 (N_11138,N_10457,N_10166);
xor U11139 (N_11139,N_10013,N_9049);
nor U11140 (N_11140,N_9921,N_9799);
nand U11141 (N_11141,N_9218,N_10040);
and U11142 (N_11142,N_9532,N_9450);
or U11143 (N_11143,N_9732,N_10475);
nand U11144 (N_11144,N_9810,N_9843);
or U11145 (N_11145,N_9905,N_9759);
and U11146 (N_11146,N_9523,N_10164);
nand U11147 (N_11147,N_9463,N_9128);
or U11148 (N_11148,N_10216,N_9780);
nor U11149 (N_11149,N_9920,N_9978);
nand U11150 (N_11150,N_9083,N_10221);
or U11151 (N_11151,N_9348,N_9009);
nor U11152 (N_11152,N_10480,N_10252);
nor U11153 (N_11153,N_9671,N_10331);
xnor U11154 (N_11154,N_9747,N_10392);
nand U11155 (N_11155,N_10426,N_9909);
nor U11156 (N_11156,N_10369,N_9003);
nor U11157 (N_11157,N_9148,N_9234);
or U11158 (N_11158,N_10346,N_9278);
xnor U11159 (N_11159,N_10380,N_9860);
xor U11160 (N_11160,N_10217,N_10070);
nor U11161 (N_11161,N_9229,N_9092);
and U11162 (N_11162,N_9771,N_9478);
or U11163 (N_11163,N_10140,N_9792);
nand U11164 (N_11164,N_9398,N_9089);
or U11165 (N_11165,N_10333,N_9566);
nand U11166 (N_11166,N_10051,N_10250);
or U11167 (N_11167,N_10145,N_9820);
or U11168 (N_11168,N_9841,N_9935);
xnor U11169 (N_11169,N_10357,N_9603);
or U11170 (N_11170,N_10374,N_9826);
and U11171 (N_11171,N_10101,N_10200);
or U11172 (N_11172,N_9854,N_9895);
or U11173 (N_11173,N_9892,N_9378);
and U11174 (N_11174,N_9690,N_9922);
xor U11175 (N_11175,N_9513,N_9669);
nor U11176 (N_11176,N_9721,N_10106);
nand U11177 (N_11177,N_9552,N_10132);
nor U11178 (N_11178,N_9963,N_9906);
or U11179 (N_11179,N_9954,N_10161);
nand U11180 (N_11180,N_9220,N_9541);
xor U11181 (N_11181,N_9815,N_9309);
nor U11182 (N_11182,N_9528,N_10286);
or U11183 (N_11183,N_10400,N_9315);
xnor U11184 (N_11184,N_9687,N_9374);
or U11185 (N_11185,N_9944,N_9456);
xor U11186 (N_11186,N_9173,N_9520);
xor U11187 (N_11187,N_9746,N_9167);
and U11188 (N_11188,N_9211,N_9390);
nand U11189 (N_11189,N_9925,N_9444);
or U11190 (N_11190,N_10168,N_10205);
or U11191 (N_11191,N_9302,N_9341);
xor U11192 (N_11192,N_10063,N_10491);
and U11193 (N_11193,N_9486,N_9886);
nand U11194 (N_11194,N_9066,N_10084);
nor U11195 (N_11195,N_10281,N_9466);
nand U11196 (N_11196,N_9259,N_10336);
and U11197 (N_11197,N_9316,N_9807);
and U11198 (N_11198,N_9047,N_9156);
or U11199 (N_11199,N_10213,N_9113);
or U11200 (N_11200,N_10310,N_9919);
and U11201 (N_11201,N_9412,N_9953);
nand U11202 (N_11202,N_9044,N_9988);
xnor U11203 (N_11203,N_9579,N_9484);
nor U11204 (N_11204,N_10306,N_10105);
nor U11205 (N_11205,N_10463,N_9555);
xnor U11206 (N_11206,N_9798,N_9177);
and U11207 (N_11207,N_10461,N_9058);
nor U11208 (N_11208,N_9120,N_10343);
nor U11209 (N_11209,N_9190,N_9970);
and U11210 (N_11210,N_10239,N_10424);
and U11211 (N_11211,N_10165,N_9531);
or U11212 (N_11212,N_9949,N_9033);
or U11213 (N_11213,N_9172,N_10074);
xnor U11214 (N_11214,N_10406,N_10460);
nor U11215 (N_11215,N_10189,N_9756);
xnor U11216 (N_11216,N_9294,N_9942);
and U11217 (N_11217,N_9448,N_9943);
nand U11218 (N_11218,N_9468,N_9585);
nand U11219 (N_11219,N_9432,N_9213);
and U11220 (N_11220,N_9457,N_9265);
nor U11221 (N_11221,N_9686,N_9781);
and U11222 (N_11222,N_9612,N_9246);
nand U11223 (N_11223,N_9335,N_9610);
xor U11224 (N_11224,N_9614,N_9600);
nor U11225 (N_11225,N_9587,N_10159);
or U11226 (N_11226,N_10226,N_9697);
or U11227 (N_11227,N_10026,N_9334);
nor U11228 (N_11228,N_9195,N_9021);
or U11229 (N_11229,N_9573,N_9281);
nor U11230 (N_11230,N_10399,N_9932);
xnor U11231 (N_11231,N_9655,N_9510);
nand U11232 (N_11232,N_9231,N_9333);
xnor U11233 (N_11233,N_10080,N_9594);
or U11234 (N_11234,N_9171,N_9933);
or U11235 (N_11235,N_9413,N_10001);
or U11236 (N_11236,N_9509,N_10355);
or U11237 (N_11237,N_10124,N_10358);
xnor U11238 (N_11238,N_10282,N_9524);
nor U11239 (N_11239,N_9691,N_9491);
xnor U11240 (N_11240,N_10396,N_10022);
and U11241 (N_11241,N_10375,N_10364);
nor U11242 (N_11242,N_10459,N_9382);
xnor U11243 (N_11243,N_9272,N_9289);
xnor U11244 (N_11244,N_9185,N_10319);
xor U11245 (N_11245,N_9548,N_9210);
or U11246 (N_11246,N_9845,N_9313);
xnor U11247 (N_11247,N_9124,N_9938);
or U11248 (N_11248,N_10274,N_9101);
and U11249 (N_11249,N_9580,N_9916);
nor U11250 (N_11250,N_9449,N_10042);
nand U11251 (N_11251,N_10201,N_10276);
xnor U11252 (N_11252,N_9017,N_9711);
or U11253 (N_11253,N_10082,N_10042);
xor U11254 (N_11254,N_9873,N_9011);
and U11255 (N_11255,N_10020,N_9330);
nand U11256 (N_11256,N_10181,N_10208);
or U11257 (N_11257,N_9833,N_9529);
and U11258 (N_11258,N_9019,N_10119);
or U11259 (N_11259,N_10492,N_9659);
or U11260 (N_11260,N_9311,N_9442);
xor U11261 (N_11261,N_9793,N_10142);
and U11262 (N_11262,N_9514,N_9535);
or U11263 (N_11263,N_10418,N_9932);
and U11264 (N_11264,N_10147,N_9849);
nor U11265 (N_11265,N_9655,N_9268);
and U11266 (N_11266,N_10177,N_9536);
xnor U11267 (N_11267,N_9166,N_9196);
nand U11268 (N_11268,N_9946,N_10252);
or U11269 (N_11269,N_9325,N_9026);
or U11270 (N_11270,N_10462,N_9743);
and U11271 (N_11271,N_9174,N_10308);
or U11272 (N_11272,N_10085,N_9158);
and U11273 (N_11273,N_10129,N_10035);
or U11274 (N_11274,N_9388,N_9123);
nor U11275 (N_11275,N_10322,N_9868);
nor U11276 (N_11276,N_9555,N_9283);
nand U11277 (N_11277,N_9793,N_10165);
nor U11278 (N_11278,N_10226,N_9660);
nor U11279 (N_11279,N_9767,N_9843);
or U11280 (N_11280,N_9647,N_9391);
nor U11281 (N_11281,N_9546,N_10439);
nand U11282 (N_11282,N_9164,N_10274);
or U11283 (N_11283,N_9602,N_10489);
nand U11284 (N_11284,N_10282,N_9452);
nand U11285 (N_11285,N_9262,N_9984);
and U11286 (N_11286,N_9141,N_9339);
xnor U11287 (N_11287,N_9982,N_9343);
nand U11288 (N_11288,N_10195,N_9159);
nand U11289 (N_11289,N_9146,N_9133);
or U11290 (N_11290,N_9623,N_9371);
and U11291 (N_11291,N_9229,N_10298);
and U11292 (N_11292,N_10053,N_9371);
and U11293 (N_11293,N_9907,N_9103);
and U11294 (N_11294,N_10160,N_10359);
nor U11295 (N_11295,N_10250,N_9143);
nand U11296 (N_11296,N_9008,N_10447);
nand U11297 (N_11297,N_10442,N_9603);
nor U11298 (N_11298,N_9168,N_9144);
nand U11299 (N_11299,N_10325,N_10085);
nand U11300 (N_11300,N_10383,N_9027);
nor U11301 (N_11301,N_10094,N_10194);
or U11302 (N_11302,N_9109,N_9446);
nand U11303 (N_11303,N_9173,N_10492);
nand U11304 (N_11304,N_10186,N_9643);
and U11305 (N_11305,N_9031,N_9416);
or U11306 (N_11306,N_9773,N_9368);
or U11307 (N_11307,N_9891,N_9387);
or U11308 (N_11308,N_10316,N_9711);
nand U11309 (N_11309,N_9280,N_9465);
xnor U11310 (N_11310,N_10279,N_10368);
nor U11311 (N_11311,N_9934,N_9096);
nand U11312 (N_11312,N_9984,N_10477);
or U11313 (N_11313,N_9180,N_10363);
nand U11314 (N_11314,N_9091,N_9293);
nand U11315 (N_11315,N_10075,N_10350);
xor U11316 (N_11316,N_10361,N_10051);
nand U11317 (N_11317,N_9972,N_10488);
and U11318 (N_11318,N_10188,N_10230);
or U11319 (N_11319,N_10008,N_9809);
and U11320 (N_11320,N_10337,N_9378);
nand U11321 (N_11321,N_9202,N_9648);
xnor U11322 (N_11322,N_9668,N_9538);
nand U11323 (N_11323,N_9347,N_9801);
or U11324 (N_11324,N_9757,N_9436);
or U11325 (N_11325,N_10344,N_9764);
xnor U11326 (N_11326,N_9677,N_10398);
nor U11327 (N_11327,N_9528,N_10070);
and U11328 (N_11328,N_9747,N_10213);
and U11329 (N_11329,N_10081,N_9708);
nand U11330 (N_11330,N_10037,N_9642);
xnor U11331 (N_11331,N_10473,N_9595);
or U11332 (N_11332,N_9508,N_9769);
nand U11333 (N_11333,N_9433,N_10286);
and U11334 (N_11334,N_9188,N_9357);
nand U11335 (N_11335,N_10202,N_10248);
xor U11336 (N_11336,N_9755,N_9100);
nand U11337 (N_11337,N_9753,N_9041);
nor U11338 (N_11338,N_9639,N_9748);
nor U11339 (N_11339,N_10472,N_10270);
nand U11340 (N_11340,N_9841,N_9928);
or U11341 (N_11341,N_9721,N_10028);
or U11342 (N_11342,N_10334,N_9983);
nand U11343 (N_11343,N_9569,N_9946);
nor U11344 (N_11344,N_9641,N_9468);
xor U11345 (N_11345,N_9368,N_9363);
and U11346 (N_11346,N_10097,N_10087);
nand U11347 (N_11347,N_9824,N_9711);
nor U11348 (N_11348,N_9645,N_9273);
or U11349 (N_11349,N_9600,N_10487);
xnor U11350 (N_11350,N_9626,N_9510);
and U11351 (N_11351,N_9512,N_9549);
or U11352 (N_11352,N_9837,N_9674);
nand U11353 (N_11353,N_9238,N_10313);
xnor U11354 (N_11354,N_9941,N_9186);
nand U11355 (N_11355,N_10450,N_10235);
nand U11356 (N_11356,N_9310,N_9789);
nor U11357 (N_11357,N_10022,N_9260);
and U11358 (N_11358,N_10447,N_9123);
and U11359 (N_11359,N_9908,N_9652);
nand U11360 (N_11360,N_9407,N_10251);
nand U11361 (N_11361,N_9734,N_10332);
xor U11362 (N_11362,N_9263,N_9765);
xnor U11363 (N_11363,N_9397,N_9050);
nor U11364 (N_11364,N_9981,N_10084);
nor U11365 (N_11365,N_10114,N_9595);
nand U11366 (N_11366,N_10359,N_9037);
or U11367 (N_11367,N_9993,N_9424);
nor U11368 (N_11368,N_9071,N_10360);
nor U11369 (N_11369,N_10021,N_9992);
or U11370 (N_11370,N_10475,N_9669);
xor U11371 (N_11371,N_9596,N_10037);
or U11372 (N_11372,N_9308,N_9845);
xor U11373 (N_11373,N_9976,N_10113);
nand U11374 (N_11374,N_9911,N_9375);
nand U11375 (N_11375,N_9856,N_9398);
xnor U11376 (N_11376,N_9414,N_9172);
or U11377 (N_11377,N_9242,N_10034);
nor U11378 (N_11378,N_9380,N_9862);
nor U11379 (N_11379,N_9889,N_10115);
xor U11380 (N_11380,N_9798,N_9294);
nand U11381 (N_11381,N_10020,N_10003);
nand U11382 (N_11382,N_9109,N_9049);
nor U11383 (N_11383,N_9070,N_9074);
or U11384 (N_11384,N_10020,N_9406);
xor U11385 (N_11385,N_9472,N_10310);
nand U11386 (N_11386,N_9573,N_10185);
and U11387 (N_11387,N_9622,N_9177);
nand U11388 (N_11388,N_9801,N_10345);
and U11389 (N_11389,N_9438,N_9471);
or U11390 (N_11390,N_10134,N_10190);
and U11391 (N_11391,N_10300,N_9516);
and U11392 (N_11392,N_9460,N_9456);
xnor U11393 (N_11393,N_10297,N_9781);
xnor U11394 (N_11394,N_10261,N_9925);
and U11395 (N_11395,N_9015,N_9366);
and U11396 (N_11396,N_9359,N_9043);
nor U11397 (N_11397,N_10498,N_10121);
and U11398 (N_11398,N_10371,N_10133);
or U11399 (N_11399,N_9534,N_10155);
or U11400 (N_11400,N_10017,N_9183);
and U11401 (N_11401,N_10405,N_9286);
nand U11402 (N_11402,N_10333,N_9451);
and U11403 (N_11403,N_9176,N_10484);
and U11404 (N_11404,N_10329,N_9450);
xor U11405 (N_11405,N_9660,N_9356);
or U11406 (N_11406,N_9143,N_9366);
nor U11407 (N_11407,N_9637,N_10250);
and U11408 (N_11408,N_9956,N_10294);
or U11409 (N_11409,N_10271,N_9379);
or U11410 (N_11410,N_9852,N_9767);
nand U11411 (N_11411,N_9313,N_10236);
xnor U11412 (N_11412,N_9219,N_9549);
and U11413 (N_11413,N_9733,N_10174);
or U11414 (N_11414,N_9216,N_9856);
nand U11415 (N_11415,N_9668,N_9807);
nor U11416 (N_11416,N_10221,N_9659);
nand U11417 (N_11417,N_9487,N_9142);
and U11418 (N_11418,N_9813,N_9337);
and U11419 (N_11419,N_9814,N_9197);
and U11420 (N_11420,N_10252,N_10460);
or U11421 (N_11421,N_9336,N_9055);
and U11422 (N_11422,N_10381,N_9271);
nand U11423 (N_11423,N_9522,N_9495);
nor U11424 (N_11424,N_9601,N_9661);
nand U11425 (N_11425,N_9323,N_9956);
or U11426 (N_11426,N_9383,N_9653);
nor U11427 (N_11427,N_10367,N_9729);
nor U11428 (N_11428,N_9951,N_10036);
xnor U11429 (N_11429,N_9896,N_9744);
nand U11430 (N_11430,N_10424,N_9759);
and U11431 (N_11431,N_9930,N_9754);
and U11432 (N_11432,N_9454,N_9398);
xnor U11433 (N_11433,N_9865,N_10146);
nor U11434 (N_11434,N_9302,N_9202);
xor U11435 (N_11435,N_9509,N_9448);
xnor U11436 (N_11436,N_9966,N_10015);
and U11437 (N_11437,N_9893,N_9489);
nand U11438 (N_11438,N_10179,N_10487);
or U11439 (N_11439,N_10263,N_9889);
nand U11440 (N_11440,N_10173,N_9418);
and U11441 (N_11441,N_10303,N_9814);
nand U11442 (N_11442,N_10421,N_9020);
xnor U11443 (N_11443,N_9195,N_10231);
nand U11444 (N_11444,N_9558,N_10477);
nand U11445 (N_11445,N_9714,N_9475);
nand U11446 (N_11446,N_10478,N_9345);
nand U11447 (N_11447,N_10244,N_9704);
or U11448 (N_11448,N_9602,N_9564);
nand U11449 (N_11449,N_9235,N_10354);
nor U11450 (N_11450,N_9115,N_10240);
and U11451 (N_11451,N_9215,N_10109);
or U11452 (N_11452,N_9667,N_9813);
nand U11453 (N_11453,N_10215,N_10458);
or U11454 (N_11454,N_10433,N_9703);
or U11455 (N_11455,N_10396,N_9045);
xor U11456 (N_11456,N_10409,N_10462);
nor U11457 (N_11457,N_9420,N_10360);
nand U11458 (N_11458,N_9790,N_9272);
nor U11459 (N_11459,N_9448,N_10202);
nor U11460 (N_11460,N_10128,N_10110);
xor U11461 (N_11461,N_9287,N_10043);
nor U11462 (N_11462,N_10061,N_9860);
nand U11463 (N_11463,N_9414,N_9868);
and U11464 (N_11464,N_10420,N_9441);
or U11465 (N_11465,N_9075,N_9234);
or U11466 (N_11466,N_9845,N_9554);
or U11467 (N_11467,N_9486,N_10112);
nor U11468 (N_11468,N_9088,N_9149);
or U11469 (N_11469,N_9461,N_9181);
xor U11470 (N_11470,N_9678,N_10237);
or U11471 (N_11471,N_9468,N_10076);
or U11472 (N_11472,N_9822,N_9587);
nor U11473 (N_11473,N_9562,N_9535);
and U11474 (N_11474,N_9155,N_9274);
nand U11475 (N_11475,N_10260,N_9019);
and U11476 (N_11476,N_9828,N_9622);
nand U11477 (N_11477,N_10102,N_10269);
and U11478 (N_11478,N_10025,N_10398);
and U11479 (N_11479,N_9997,N_9808);
xor U11480 (N_11480,N_9388,N_9892);
and U11481 (N_11481,N_9716,N_9814);
xnor U11482 (N_11482,N_10368,N_10329);
and U11483 (N_11483,N_9253,N_9063);
xor U11484 (N_11484,N_10239,N_10285);
xor U11485 (N_11485,N_9536,N_9991);
and U11486 (N_11486,N_10089,N_9174);
and U11487 (N_11487,N_10051,N_9020);
nand U11488 (N_11488,N_10175,N_10420);
nor U11489 (N_11489,N_9954,N_10282);
and U11490 (N_11490,N_10323,N_9445);
xor U11491 (N_11491,N_10347,N_10197);
nor U11492 (N_11492,N_9604,N_9402);
xor U11493 (N_11493,N_9389,N_9026);
or U11494 (N_11494,N_9360,N_9422);
nand U11495 (N_11495,N_10268,N_10462);
nor U11496 (N_11496,N_9995,N_9141);
nand U11497 (N_11497,N_9662,N_9910);
or U11498 (N_11498,N_9321,N_9750);
or U11499 (N_11499,N_10034,N_10195);
nor U11500 (N_11500,N_9545,N_9135);
and U11501 (N_11501,N_9624,N_10103);
nand U11502 (N_11502,N_10322,N_10464);
and U11503 (N_11503,N_10428,N_10233);
xor U11504 (N_11504,N_9954,N_9148);
xor U11505 (N_11505,N_10489,N_9282);
nor U11506 (N_11506,N_9516,N_9886);
xor U11507 (N_11507,N_10041,N_10361);
nand U11508 (N_11508,N_10222,N_9481);
and U11509 (N_11509,N_9207,N_9790);
nand U11510 (N_11510,N_9413,N_9754);
nand U11511 (N_11511,N_9348,N_10422);
nor U11512 (N_11512,N_9043,N_9645);
or U11513 (N_11513,N_10136,N_9712);
or U11514 (N_11514,N_9799,N_10046);
and U11515 (N_11515,N_9036,N_9332);
nor U11516 (N_11516,N_9405,N_9323);
xor U11517 (N_11517,N_9723,N_10139);
nor U11518 (N_11518,N_9889,N_10111);
nor U11519 (N_11519,N_9589,N_9127);
nand U11520 (N_11520,N_9458,N_10368);
nand U11521 (N_11521,N_9921,N_9430);
or U11522 (N_11522,N_9371,N_9101);
and U11523 (N_11523,N_10125,N_10132);
and U11524 (N_11524,N_9095,N_10341);
nand U11525 (N_11525,N_9094,N_9027);
and U11526 (N_11526,N_10440,N_9593);
nor U11527 (N_11527,N_10497,N_9016);
and U11528 (N_11528,N_9875,N_10064);
and U11529 (N_11529,N_10135,N_9074);
nor U11530 (N_11530,N_10227,N_9542);
nor U11531 (N_11531,N_10390,N_9069);
nand U11532 (N_11532,N_10295,N_10161);
or U11533 (N_11533,N_10328,N_10315);
or U11534 (N_11534,N_10428,N_9504);
nor U11535 (N_11535,N_10397,N_9923);
xor U11536 (N_11536,N_9557,N_9000);
or U11537 (N_11537,N_9529,N_9032);
nand U11538 (N_11538,N_10227,N_9594);
or U11539 (N_11539,N_10070,N_9320);
xor U11540 (N_11540,N_9566,N_9292);
and U11541 (N_11541,N_10246,N_9500);
nand U11542 (N_11542,N_9944,N_9887);
or U11543 (N_11543,N_9417,N_9782);
xor U11544 (N_11544,N_9384,N_9877);
or U11545 (N_11545,N_9056,N_9396);
nand U11546 (N_11546,N_9959,N_9683);
nand U11547 (N_11547,N_9151,N_10061);
or U11548 (N_11548,N_9604,N_10175);
or U11549 (N_11549,N_10119,N_10420);
nor U11550 (N_11550,N_9131,N_10247);
xnor U11551 (N_11551,N_10098,N_10242);
nand U11552 (N_11552,N_9253,N_10327);
and U11553 (N_11553,N_9699,N_9950);
nor U11554 (N_11554,N_9192,N_10358);
nand U11555 (N_11555,N_10432,N_9930);
nor U11556 (N_11556,N_10344,N_9059);
and U11557 (N_11557,N_10027,N_9008);
nor U11558 (N_11558,N_9850,N_9936);
and U11559 (N_11559,N_10443,N_9804);
nand U11560 (N_11560,N_10031,N_9070);
and U11561 (N_11561,N_9418,N_9753);
nand U11562 (N_11562,N_9138,N_9642);
or U11563 (N_11563,N_9308,N_9544);
nand U11564 (N_11564,N_9699,N_10471);
and U11565 (N_11565,N_9088,N_10412);
and U11566 (N_11566,N_9507,N_10202);
nor U11567 (N_11567,N_10383,N_9698);
xor U11568 (N_11568,N_9316,N_9617);
nor U11569 (N_11569,N_9470,N_9623);
and U11570 (N_11570,N_9966,N_9811);
and U11571 (N_11571,N_9302,N_9947);
xor U11572 (N_11572,N_9789,N_10234);
nand U11573 (N_11573,N_9880,N_9139);
xor U11574 (N_11574,N_9321,N_9176);
nor U11575 (N_11575,N_10439,N_9369);
or U11576 (N_11576,N_9339,N_9154);
and U11577 (N_11577,N_9701,N_9803);
nor U11578 (N_11578,N_9668,N_9909);
xor U11579 (N_11579,N_9712,N_9989);
and U11580 (N_11580,N_9407,N_9576);
nand U11581 (N_11581,N_9020,N_10092);
xnor U11582 (N_11582,N_9404,N_9035);
nand U11583 (N_11583,N_10443,N_10072);
xnor U11584 (N_11584,N_10235,N_10292);
or U11585 (N_11585,N_9560,N_9931);
or U11586 (N_11586,N_9817,N_9637);
and U11587 (N_11587,N_9414,N_10047);
and U11588 (N_11588,N_9928,N_10074);
xnor U11589 (N_11589,N_9700,N_10257);
xor U11590 (N_11590,N_9226,N_9804);
and U11591 (N_11591,N_9628,N_9398);
or U11592 (N_11592,N_10083,N_9551);
nor U11593 (N_11593,N_9617,N_10069);
and U11594 (N_11594,N_9583,N_9836);
and U11595 (N_11595,N_9748,N_10192);
nor U11596 (N_11596,N_9063,N_9840);
xnor U11597 (N_11597,N_9759,N_9261);
nor U11598 (N_11598,N_9551,N_10092);
nand U11599 (N_11599,N_9235,N_10478);
nor U11600 (N_11600,N_9171,N_10069);
nor U11601 (N_11601,N_10498,N_9311);
nor U11602 (N_11602,N_9765,N_9785);
or U11603 (N_11603,N_9228,N_9368);
or U11604 (N_11604,N_9801,N_10452);
nor U11605 (N_11605,N_9675,N_9269);
or U11606 (N_11606,N_9797,N_9697);
nor U11607 (N_11607,N_9123,N_9488);
nor U11608 (N_11608,N_9367,N_9339);
or U11609 (N_11609,N_9255,N_9458);
nand U11610 (N_11610,N_9427,N_10375);
or U11611 (N_11611,N_10247,N_9196);
and U11612 (N_11612,N_10454,N_9977);
nor U11613 (N_11613,N_9664,N_10188);
or U11614 (N_11614,N_10065,N_10177);
xor U11615 (N_11615,N_9274,N_10199);
or U11616 (N_11616,N_9301,N_9329);
nand U11617 (N_11617,N_9834,N_9311);
and U11618 (N_11618,N_10094,N_9690);
and U11619 (N_11619,N_10403,N_10432);
xor U11620 (N_11620,N_10137,N_9497);
nor U11621 (N_11621,N_10278,N_9451);
and U11622 (N_11622,N_9607,N_9740);
and U11623 (N_11623,N_10373,N_9352);
xnor U11624 (N_11624,N_9822,N_9826);
xnor U11625 (N_11625,N_10229,N_9961);
xnor U11626 (N_11626,N_9126,N_9473);
xnor U11627 (N_11627,N_9081,N_9439);
xnor U11628 (N_11628,N_9401,N_9839);
nand U11629 (N_11629,N_9290,N_10254);
and U11630 (N_11630,N_10229,N_9512);
xnor U11631 (N_11631,N_9639,N_9588);
and U11632 (N_11632,N_10155,N_10199);
xor U11633 (N_11633,N_9062,N_9320);
nand U11634 (N_11634,N_9913,N_9276);
nor U11635 (N_11635,N_10467,N_10399);
xor U11636 (N_11636,N_9233,N_9745);
nand U11637 (N_11637,N_10171,N_10052);
xor U11638 (N_11638,N_10297,N_9878);
and U11639 (N_11639,N_9442,N_9412);
and U11640 (N_11640,N_9670,N_9687);
or U11641 (N_11641,N_9946,N_9848);
or U11642 (N_11642,N_10093,N_10011);
xor U11643 (N_11643,N_9988,N_10213);
and U11644 (N_11644,N_10311,N_9704);
and U11645 (N_11645,N_10063,N_9252);
nor U11646 (N_11646,N_10295,N_9384);
nor U11647 (N_11647,N_9727,N_9477);
or U11648 (N_11648,N_9992,N_10436);
and U11649 (N_11649,N_9776,N_9977);
xnor U11650 (N_11650,N_9302,N_9397);
xnor U11651 (N_11651,N_9295,N_9225);
xor U11652 (N_11652,N_9678,N_9861);
nand U11653 (N_11653,N_9695,N_10405);
or U11654 (N_11654,N_10440,N_9873);
and U11655 (N_11655,N_9413,N_10120);
xor U11656 (N_11656,N_9140,N_10344);
xor U11657 (N_11657,N_9381,N_9780);
nand U11658 (N_11658,N_10058,N_9340);
xor U11659 (N_11659,N_10226,N_9920);
nand U11660 (N_11660,N_10485,N_9263);
and U11661 (N_11661,N_9782,N_10440);
nor U11662 (N_11662,N_10243,N_9770);
nand U11663 (N_11663,N_10151,N_9908);
xor U11664 (N_11664,N_10241,N_9524);
and U11665 (N_11665,N_9547,N_10240);
xor U11666 (N_11666,N_9927,N_10145);
xor U11667 (N_11667,N_10005,N_9979);
and U11668 (N_11668,N_10487,N_9405);
or U11669 (N_11669,N_9499,N_10391);
or U11670 (N_11670,N_9397,N_9857);
and U11671 (N_11671,N_9767,N_9373);
and U11672 (N_11672,N_10344,N_9987);
nand U11673 (N_11673,N_10133,N_9671);
and U11674 (N_11674,N_9952,N_9650);
and U11675 (N_11675,N_9843,N_9073);
or U11676 (N_11676,N_9126,N_10407);
and U11677 (N_11677,N_9084,N_9379);
nand U11678 (N_11678,N_9941,N_9661);
or U11679 (N_11679,N_9415,N_10401);
xor U11680 (N_11680,N_9174,N_9298);
xor U11681 (N_11681,N_9842,N_10092);
nand U11682 (N_11682,N_10236,N_9473);
nor U11683 (N_11683,N_9831,N_9712);
xnor U11684 (N_11684,N_9079,N_9151);
xor U11685 (N_11685,N_9781,N_10081);
and U11686 (N_11686,N_9233,N_9863);
nor U11687 (N_11687,N_9863,N_10414);
or U11688 (N_11688,N_10386,N_10485);
nor U11689 (N_11689,N_9222,N_9075);
and U11690 (N_11690,N_10371,N_9648);
nor U11691 (N_11691,N_9074,N_9791);
nor U11692 (N_11692,N_9834,N_10227);
xnor U11693 (N_11693,N_9710,N_9511);
nand U11694 (N_11694,N_10060,N_9879);
or U11695 (N_11695,N_9476,N_10145);
or U11696 (N_11696,N_9412,N_9908);
nor U11697 (N_11697,N_10172,N_9290);
nor U11698 (N_11698,N_10472,N_10277);
and U11699 (N_11699,N_9957,N_9952);
nor U11700 (N_11700,N_9355,N_9911);
nor U11701 (N_11701,N_10157,N_9582);
or U11702 (N_11702,N_9242,N_9863);
xnor U11703 (N_11703,N_10268,N_10235);
and U11704 (N_11704,N_9826,N_10491);
xnor U11705 (N_11705,N_9319,N_9996);
and U11706 (N_11706,N_9418,N_10486);
and U11707 (N_11707,N_9890,N_10031);
nand U11708 (N_11708,N_10481,N_9295);
xnor U11709 (N_11709,N_9398,N_9509);
nor U11710 (N_11710,N_10122,N_9569);
and U11711 (N_11711,N_9165,N_9827);
or U11712 (N_11712,N_9529,N_10460);
nor U11713 (N_11713,N_9128,N_10444);
or U11714 (N_11714,N_9870,N_9568);
and U11715 (N_11715,N_9504,N_9992);
nand U11716 (N_11716,N_9277,N_9979);
xnor U11717 (N_11717,N_9178,N_9771);
xor U11718 (N_11718,N_9457,N_10122);
nor U11719 (N_11719,N_10289,N_9985);
nand U11720 (N_11720,N_9562,N_10236);
xor U11721 (N_11721,N_9900,N_9073);
and U11722 (N_11722,N_10263,N_10323);
and U11723 (N_11723,N_9964,N_10016);
and U11724 (N_11724,N_9573,N_9773);
or U11725 (N_11725,N_9818,N_10231);
or U11726 (N_11726,N_9852,N_9762);
xnor U11727 (N_11727,N_10431,N_9995);
and U11728 (N_11728,N_10413,N_9706);
nor U11729 (N_11729,N_10286,N_9218);
nor U11730 (N_11730,N_10016,N_9366);
xor U11731 (N_11731,N_9272,N_9077);
xor U11732 (N_11732,N_9691,N_9063);
and U11733 (N_11733,N_9350,N_10297);
and U11734 (N_11734,N_10461,N_10226);
and U11735 (N_11735,N_9652,N_9834);
or U11736 (N_11736,N_9092,N_9687);
and U11737 (N_11737,N_10266,N_10420);
and U11738 (N_11738,N_9792,N_10202);
or U11739 (N_11739,N_9410,N_9757);
xor U11740 (N_11740,N_10206,N_9025);
and U11741 (N_11741,N_10390,N_9500);
xnor U11742 (N_11742,N_9305,N_9446);
nand U11743 (N_11743,N_9091,N_9592);
xnor U11744 (N_11744,N_9390,N_9417);
nand U11745 (N_11745,N_9431,N_9424);
xnor U11746 (N_11746,N_10064,N_10427);
xor U11747 (N_11747,N_10449,N_9125);
nand U11748 (N_11748,N_9992,N_10312);
xor U11749 (N_11749,N_9512,N_9727);
nand U11750 (N_11750,N_9650,N_9168);
nor U11751 (N_11751,N_9702,N_9663);
nor U11752 (N_11752,N_10303,N_9464);
or U11753 (N_11753,N_10425,N_9667);
xnor U11754 (N_11754,N_10435,N_9780);
xnor U11755 (N_11755,N_9707,N_9053);
xnor U11756 (N_11756,N_9414,N_9045);
or U11757 (N_11757,N_10443,N_9263);
xnor U11758 (N_11758,N_9450,N_9294);
or U11759 (N_11759,N_9605,N_9907);
nand U11760 (N_11760,N_10215,N_9031);
xor U11761 (N_11761,N_9395,N_9090);
nand U11762 (N_11762,N_10183,N_9751);
nor U11763 (N_11763,N_9029,N_9581);
nor U11764 (N_11764,N_9425,N_9853);
or U11765 (N_11765,N_10203,N_10288);
and U11766 (N_11766,N_9995,N_9404);
nand U11767 (N_11767,N_10347,N_10118);
xnor U11768 (N_11768,N_10084,N_9340);
nor U11769 (N_11769,N_9961,N_9789);
or U11770 (N_11770,N_9064,N_9505);
nand U11771 (N_11771,N_9433,N_9722);
nor U11772 (N_11772,N_9344,N_9147);
nand U11773 (N_11773,N_9964,N_9046);
and U11774 (N_11774,N_9836,N_10132);
xor U11775 (N_11775,N_9477,N_10126);
and U11776 (N_11776,N_10059,N_10331);
xnor U11777 (N_11777,N_9093,N_9746);
or U11778 (N_11778,N_9170,N_10404);
or U11779 (N_11779,N_10304,N_9809);
xnor U11780 (N_11780,N_9203,N_9324);
and U11781 (N_11781,N_9011,N_10378);
nor U11782 (N_11782,N_9500,N_9794);
and U11783 (N_11783,N_9081,N_9564);
and U11784 (N_11784,N_10017,N_9831);
and U11785 (N_11785,N_10224,N_9468);
xor U11786 (N_11786,N_9329,N_9945);
or U11787 (N_11787,N_10370,N_9425);
and U11788 (N_11788,N_9612,N_9243);
xnor U11789 (N_11789,N_9670,N_9581);
nor U11790 (N_11790,N_9144,N_9729);
nand U11791 (N_11791,N_10436,N_9214);
or U11792 (N_11792,N_10172,N_9814);
xor U11793 (N_11793,N_10281,N_9797);
or U11794 (N_11794,N_9311,N_10108);
nor U11795 (N_11795,N_10278,N_10134);
or U11796 (N_11796,N_9761,N_10090);
nand U11797 (N_11797,N_10242,N_10410);
and U11798 (N_11798,N_9426,N_10032);
and U11799 (N_11799,N_9293,N_9681);
xor U11800 (N_11800,N_9020,N_9048);
nand U11801 (N_11801,N_9094,N_9959);
and U11802 (N_11802,N_9775,N_9699);
nand U11803 (N_11803,N_10327,N_10068);
nor U11804 (N_11804,N_9567,N_9347);
or U11805 (N_11805,N_9002,N_9946);
or U11806 (N_11806,N_9504,N_9875);
xnor U11807 (N_11807,N_10397,N_9881);
or U11808 (N_11808,N_10229,N_9632);
xor U11809 (N_11809,N_10042,N_10169);
and U11810 (N_11810,N_9542,N_9923);
nor U11811 (N_11811,N_9900,N_10318);
nor U11812 (N_11812,N_9666,N_10388);
and U11813 (N_11813,N_9385,N_9980);
nor U11814 (N_11814,N_10281,N_10194);
xnor U11815 (N_11815,N_9120,N_9762);
nor U11816 (N_11816,N_9785,N_9975);
nand U11817 (N_11817,N_9993,N_9387);
or U11818 (N_11818,N_9922,N_10262);
nand U11819 (N_11819,N_10077,N_10209);
nand U11820 (N_11820,N_10119,N_9197);
or U11821 (N_11821,N_10120,N_9571);
nand U11822 (N_11822,N_9393,N_9401);
and U11823 (N_11823,N_9944,N_10203);
nand U11824 (N_11824,N_9477,N_9761);
xor U11825 (N_11825,N_9105,N_9634);
or U11826 (N_11826,N_9818,N_9940);
nor U11827 (N_11827,N_9419,N_9627);
xnor U11828 (N_11828,N_9297,N_9349);
nor U11829 (N_11829,N_10301,N_9338);
and U11830 (N_11830,N_9516,N_9632);
nand U11831 (N_11831,N_9724,N_9739);
nor U11832 (N_11832,N_9030,N_10346);
nand U11833 (N_11833,N_9115,N_9648);
xor U11834 (N_11834,N_10048,N_9335);
xor U11835 (N_11835,N_9725,N_9442);
xnor U11836 (N_11836,N_9064,N_9988);
nand U11837 (N_11837,N_10165,N_10390);
or U11838 (N_11838,N_10252,N_9032);
xnor U11839 (N_11839,N_9586,N_9077);
and U11840 (N_11840,N_10330,N_9034);
and U11841 (N_11841,N_9831,N_9901);
nor U11842 (N_11842,N_9896,N_9783);
and U11843 (N_11843,N_10075,N_10145);
and U11844 (N_11844,N_10438,N_9617);
nor U11845 (N_11845,N_10209,N_9075);
and U11846 (N_11846,N_10409,N_9842);
xnor U11847 (N_11847,N_10464,N_9246);
xor U11848 (N_11848,N_9794,N_10298);
or U11849 (N_11849,N_9685,N_10103);
nor U11850 (N_11850,N_9135,N_10378);
nor U11851 (N_11851,N_10020,N_10308);
or U11852 (N_11852,N_9483,N_9491);
or U11853 (N_11853,N_9005,N_10043);
and U11854 (N_11854,N_10336,N_10227);
nand U11855 (N_11855,N_10104,N_10430);
nor U11856 (N_11856,N_10036,N_9521);
nand U11857 (N_11857,N_10381,N_9193);
and U11858 (N_11858,N_10359,N_10223);
xnor U11859 (N_11859,N_9778,N_10121);
and U11860 (N_11860,N_9479,N_9766);
or U11861 (N_11861,N_10492,N_9165);
nand U11862 (N_11862,N_9805,N_9469);
xor U11863 (N_11863,N_9916,N_9739);
or U11864 (N_11864,N_9530,N_9657);
nor U11865 (N_11865,N_9780,N_10067);
xnor U11866 (N_11866,N_9037,N_10322);
nor U11867 (N_11867,N_9246,N_9371);
nor U11868 (N_11868,N_9300,N_10078);
xor U11869 (N_11869,N_9641,N_9077);
nor U11870 (N_11870,N_10436,N_9567);
nor U11871 (N_11871,N_10347,N_9764);
and U11872 (N_11872,N_9397,N_10159);
or U11873 (N_11873,N_9512,N_9602);
nor U11874 (N_11874,N_10169,N_9593);
nand U11875 (N_11875,N_9896,N_10415);
nor U11876 (N_11876,N_10130,N_9719);
or U11877 (N_11877,N_9908,N_9247);
or U11878 (N_11878,N_10278,N_9419);
xnor U11879 (N_11879,N_9955,N_9465);
or U11880 (N_11880,N_10493,N_9955);
nand U11881 (N_11881,N_9771,N_9222);
and U11882 (N_11882,N_10102,N_9434);
or U11883 (N_11883,N_9237,N_9359);
xnor U11884 (N_11884,N_9683,N_10403);
xor U11885 (N_11885,N_9457,N_9449);
xnor U11886 (N_11886,N_9391,N_10107);
xor U11887 (N_11887,N_10289,N_10031);
and U11888 (N_11888,N_9743,N_10351);
xor U11889 (N_11889,N_9721,N_9521);
and U11890 (N_11890,N_9357,N_9906);
and U11891 (N_11891,N_9333,N_10204);
xnor U11892 (N_11892,N_9804,N_9712);
and U11893 (N_11893,N_9191,N_9530);
nor U11894 (N_11894,N_10315,N_10014);
nand U11895 (N_11895,N_10249,N_9732);
or U11896 (N_11896,N_9318,N_9863);
nor U11897 (N_11897,N_10431,N_10015);
or U11898 (N_11898,N_9849,N_9750);
or U11899 (N_11899,N_9046,N_10208);
nand U11900 (N_11900,N_9236,N_9831);
or U11901 (N_11901,N_10204,N_9415);
nor U11902 (N_11902,N_9373,N_9394);
nand U11903 (N_11903,N_10192,N_9663);
or U11904 (N_11904,N_10135,N_9507);
or U11905 (N_11905,N_9065,N_9459);
nand U11906 (N_11906,N_10048,N_9227);
nor U11907 (N_11907,N_9320,N_9221);
nand U11908 (N_11908,N_9837,N_9578);
xnor U11909 (N_11909,N_9846,N_9001);
and U11910 (N_11910,N_9684,N_9436);
or U11911 (N_11911,N_9959,N_9063);
nand U11912 (N_11912,N_9484,N_9031);
xnor U11913 (N_11913,N_10079,N_10190);
or U11914 (N_11914,N_10175,N_9133);
or U11915 (N_11915,N_9506,N_9959);
nand U11916 (N_11916,N_9023,N_10467);
nor U11917 (N_11917,N_10428,N_10260);
xor U11918 (N_11918,N_10201,N_10044);
nand U11919 (N_11919,N_10317,N_10121);
nand U11920 (N_11920,N_9613,N_9542);
nand U11921 (N_11921,N_9011,N_10249);
xor U11922 (N_11922,N_9384,N_10376);
and U11923 (N_11923,N_10308,N_9014);
nor U11924 (N_11924,N_10381,N_9049);
nand U11925 (N_11925,N_9072,N_9777);
and U11926 (N_11926,N_10162,N_9339);
and U11927 (N_11927,N_9342,N_9111);
nand U11928 (N_11928,N_10326,N_9931);
and U11929 (N_11929,N_9632,N_10337);
or U11930 (N_11930,N_9837,N_10084);
nor U11931 (N_11931,N_9243,N_9889);
or U11932 (N_11932,N_10417,N_9448);
or U11933 (N_11933,N_9087,N_9011);
and U11934 (N_11934,N_10318,N_10072);
and U11935 (N_11935,N_9298,N_9384);
nor U11936 (N_11936,N_9108,N_9327);
xor U11937 (N_11937,N_9178,N_10058);
and U11938 (N_11938,N_10149,N_9062);
nor U11939 (N_11939,N_9978,N_9367);
nor U11940 (N_11940,N_9536,N_10375);
xnor U11941 (N_11941,N_10490,N_9533);
nand U11942 (N_11942,N_10071,N_10047);
nor U11943 (N_11943,N_9605,N_9442);
or U11944 (N_11944,N_10342,N_10471);
and U11945 (N_11945,N_9121,N_9675);
nand U11946 (N_11946,N_9738,N_10488);
nor U11947 (N_11947,N_9331,N_9239);
xnor U11948 (N_11948,N_9509,N_9959);
nor U11949 (N_11949,N_9399,N_9103);
or U11950 (N_11950,N_10218,N_10281);
xor U11951 (N_11951,N_9154,N_10285);
and U11952 (N_11952,N_9663,N_9996);
and U11953 (N_11953,N_10271,N_9425);
nor U11954 (N_11954,N_10486,N_9766);
xnor U11955 (N_11955,N_9522,N_9617);
or U11956 (N_11956,N_9162,N_10131);
nor U11957 (N_11957,N_10472,N_9517);
nor U11958 (N_11958,N_9594,N_9976);
and U11959 (N_11959,N_9522,N_9196);
or U11960 (N_11960,N_9431,N_9505);
and U11961 (N_11961,N_10425,N_10373);
nand U11962 (N_11962,N_10366,N_9200);
xnor U11963 (N_11963,N_9253,N_10343);
nand U11964 (N_11964,N_9419,N_9304);
and U11965 (N_11965,N_9533,N_9721);
or U11966 (N_11966,N_9684,N_9547);
and U11967 (N_11967,N_10320,N_10220);
xor U11968 (N_11968,N_10354,N_9996);
xor U11969 (N_11969,N_10358,N_10297);
nand U11970 (N_11970,N_9115,N_10192);
xnor U11971 (N_11971,N_10329,N_9994);
nand U11972 (N_11972,N_9663,N_10457);
nand U11973 (N_11973,N_9991,N_10196);
and U11974 (N_11974,N_9457,N_9193);
nand U11975 (N_11975,N_9518,N_10355);
nor U11976 (N_11976,N_9087,N_10449);
and U11977 (N_11977,N_10130,N_9267);
nand U11978 (N_11978,N_9281,N_9842);
and U11979 (N_11979,N_10403,N_10496);
nand U11980 (N_11980,N_9170,N_9914);
xor U11981 (N_11981,N_9313,N_10294);
and U11982 (N_11982,N_9432,N_9071);
nor U11983 (N_11983,N_10492,N_9526);
and U11984 (N_11984,N_9932,N_9460);
nor U11985 (N_11985,N_9302,N_9190);
nor U11986 (N_11986,N_10324,N_10074);
xnor U11987 (N_11987,N_9348,N_9099);
nor U11988 (N_11988,N_10051,N_10157);
and U11989 (N_11989,N_9201,N_10354);
or U11990 (N_11990,N_9628,N_9141);
nor U11991 (N_11991,N_9998,N_9472);
nor U11992 (N_11992,N_10147,N_9661);
or U11993 (N_11993,N_10390,N_10331);
nand U11994 (N_11994,N_10185,N_10307);
nor U11995 (N_11995,N_10068,N_9121);
nand U11996 (N_11996,N_9533,N_9321);
nor U11997 (N_11997,N_9518,N_9096);
nand U11998 (N_11998,N_10238,N_10225);
xor U11999 (N_11999,N_9658,N_9850);
nand U12000 (N_12000,N_11450,N_11701);
xor U12001 (N_12001,N_11359,N_11861);
nor U12002 (N_12002,N_11950,N_10611);
or U12003 (N_12003,N_11099,N_11700);
xnor U12004 (N_12004,N_11420,N_11839);
nor U12005 (N_12005,N_11334,N_11158);
or U12006 (N_12006,N_11460,N_11092);
and U12007 (N_12007,N_10889,N_11921);
xor U12008 (N_12008,N_10822,N_10801);
or U12009 (N_12009,N_10583,N_11833);
nor U12010 (N_12010,N_11090,N_11976);
xor U12011 (N_12011,N_11271,N_11198);
nand U12012 (N_12012,N_10917,N_11834);
nor U12013 (N_12013,N_11777,N_11414);
nand U12014 (N_12014,N_11072,N_10883);
or U12015 (N_12015,N_11836,N_11370);
nand U12016 (N_12016,N_10531,N_10735);
nand U12017 (N_12017,N_11905,N_11632);
and U12018 (N_12018,N_11298,N_11034);
xor U12019 (N_12019,N_10767,N_11446);
nor U12020 (N_12020,N_11115,N_10699);
or U12021 (N_12021,N_11727,N_10871);
or U12022 (N_12022,N_10588,N_10922);
nand U12023 (N_12023,N_11219,N_11728);
nor U12024 (N_12024,N_11664,N_11780);
or U12025 (N_12025,N_10865,N_11285);
xnor U12026 (N_12026,N_11979,N_10771);
nor U12027 (N_12027,N_11267,N_11181);
nand U12028 (N_12028,N_11653,N_11544);
and U12029 (N_12029,N_11984,N_11637);
nor U12030 (N_12030,N_11476,N_10915);
nor U12031 (N_12031,N_11110,N_11479);
or U12032 (N_12032,N_10624,N_11082);
xor U12033 (N_12033,N_11511,N_11699);
and U12034 (N_12034,N_11445,N_11026);
and U12035 (N_12035,N_11713,N_11991);
or U12036 (N_12036,N_11603,N_10598);
or U12037 (N_12037,N_10843,N_10813);
or U12038 (N_12038,N_11067,N_11430);
xnor U12039 (N_12039,N_11642,N_11711);
xnor U12040 (N_12040,N_11361,N_11744);
nor U12041 (N_12041,N_11855,N_11633);
nand U12042 (N_12042,N_10730,N_10600);
nand U12043 (N_12043,N_10538,N_10511);
xor U12044 (N_12044,N_11341,N_11114);
xor U12045 (N_12045,N_11073,N_10920);
xor U12046 (N_12046,N_11521,N_11952);
or U12047 (N_12047,N_10667,N_11561);
nand U12048 (N_12048,N_11883,N_11537);
xor U12049 (N_12049,N_11529,N_11309);
nor U12050 (N_12050,N_10779,N_11308);
xor U12051 (N_12051,N_11762,N_11214);
and U12052 (N_12052,N_11423,N_10565);
nor U12053 (N_12053,N_11685,N_11721);
nand U12054 (N_12054,N_10552,N_11595);
nand U12055 (N_12055,N_10919,N_11573);
xnor U12056 (N_12056,N_11571,N_11449);
nor U12057 (N_12057,N_11464,N_11550);
nor U12058 (N_12058,N_11586,N_10714);
and U12059 (N_12059,N_11525,N_10683);
xnor U12060 (N_12060,N_10693,N_10826);
nand U12061 (N_12061,N_11129,N_11391);
or U12062 (N_12062,N_11155,N_11208);
xor U12063 (N_12063,N_11792,N_11963);
nand U12064 (N_12064,N_10564,N_10949);
xor U12065 (N_12065,N_11353,N_11469);
or U12066 (N_12066,N_11184,N_11980);
nor U12067 (N_12067,N_11404,N_11927);
or U12068 (N_12068,N_11346,N_11256);
xor U12069 (N_12069,N_11212,N_11327);
nand U12070 (N_12070,N_11615,N_11585);
nand U12071 (N_12071,N_11070,N_11534);
or U12072 (N_12072,N_11645,N_11288);
nor U12073 (N_12073,N_11797,N_10869);
or U12074 (N_12074,N_11580,N_11514);
and U12075 (N_12075,N_11413,N_11251);
xnor U12076 (N_12076,N_11835,N_11107);
and U12077 (N_12077,N_11382,N_11003);
xor U12078 (N_12078,N_11336,N_10757);
nor U12079 (N_12079,N_11668,N_11331);
or U12080 (N_12080,N_11594,N_11007);
nand U12081 (N_12081,N_11051,N_10631);
xor U12082 (N_12082,N_10514,N_11558);
and U12083 (N_12083,N_10759,N_11605);
xnor U12084 (N_12084,N_10815,N_11253);
nor U12085 (N_12085,N_11022,N_11712);
nor U12086 (N_12086,N_11362,N_10851);
and U12087 (N_12087,N_10880,N_10689);
nand U12088 (N_12088,N_11720,N_10633);
nor U12089 (N_12089,N_11305,N_11737);
and U12090 (N_12090,N_11200,N_11406);
and U12091 (N_12091,N_11020,N_11857);
xor U12092 (N_12092,N_10517,N_11671);
and U12093 (N_12093,N_11674,N_11326);
nor U12094 (N_12094,N_11915,N_10964);
or U12095 (N_12095,N_11475,N_11614);
and U12096 (N_12096,N_11439,N_11260);
and U12097 (N_12097,N_10793,N_11820);
nor U12098 (N_12098,N_11386,N_10839);
and U12099 (N_12099,N_10620,N_10977);
nor U12100 (N_12100,N_11023,N_10602);
and U12101 (N_12101,N_11895,N_10664);
xor U12102 (N_12102,N_11799,N_11320);
or U12103 (N_12103,N_11667,N_11095);
and U12104 (N_12104,N_10874,N_11598);
xnor U12105 (N_12105,N_10818,N_10630);
nor U12106 (N_12106,N_11681,N_10934);
nor U12107 (N_12107,N_11228,N_11005);
xor U12108 (N_12108,N_11519,N_10824);
xnor U12109 (N_12109,N_10817,N_11376);
and U12110 (N_12110,N_11093,N_11638);
nand U12111 (N_12111,N_10705,N_11330);
or U12112 (N_12112,N_10594,N_10632);
and U12113 (N_12113,N_11501,N_10581);
nor U12114 (N_12114,N_11455,N_11488);
nor U12115 (N_12115,N_10559,N_10674);
or U12116 (N_12116,N_11788,N_11974);
xnor U12117 (N_12117,N_11136,N_11462);
nor U12118 (N_12118,N_11873,N_11496);
and U12119 (N_12119,N_10729,N_10854);
or U12120 (N_12120,N_11526,N_11069);
and U12121 (N_12121,N_11171,N_11520);
nor U12122 (N_12122,N_11793,N_11492);
xor U12123 (N_12123,N_11821,N_11772);
xor U12124 (N_12124,N_10692,N_10905);
nor U12125 (N_12125,N_11930,N_10606);
or U12126 (N_12126,N_10930,N_10884);
and U12127 (N_12127,N_10503,N_11276);
or U12128 (N_12128,N_11164,N_10777);
xor U12129 (N_12129,N_10673,N_10504);
xor U12130 (N_12130,N_11323,N_11893);
nand U12131 (N_12131,N_11452,N_11695);
and U12132 (N_12132,N_11033,N_11856);
or U12133 (N_12133,N_11961,N_11579);
nand U12134 (N_12134,N_11736,N_11495);
nor U12135 (N_12135,N_11936,N_11485);
and U12136 (N_12136,N_10876,N_10829);
or U12137 (N_12137,N_11163,N_11986);
xor U12138 (N_12138,N_11421,N_10765);
or U12139 (N_12139,N_11207,N_11890);
or U12140 (N_12140,N_10525,N_11043);
and U12141 (N_12141,N_10814,N_11075);
nor U12142 (N_12142,N_11363,N_10838);
nand U12143 (N_12143,N_11670,N_10941);
nor U12144 (N_12144,N_11871,N_10762);
nand U12145 (N_12145,N_11847,N_11328);
or U12146 (N_12146,N_11994,N_11876);
xnor U12147 (N_12147,N_10936,N_11510);
nand U12148 (N_12148,N_10660,N_10867);
nand U12149 (N_12149,N_11289,N_11397);
nor U12150 (N_12150,N_10834,N_11923);
or U12151 (N_12151,N_11045,N_10907);
or U12152 (N_12152,N_11547,N_11787);
nor U12153 (N_12153,N_11217,N_11819);
nor U12154 (N_12154,N_10805,N_11827);
nand U12155 (N_12155,N_10873,N_11731);
or U12156 (N_12156,N_11059,N_11229);
and U12157 (N_12157,N_11355,N_11745);
nor U12158 (N_12158,N_11539,N_11132);
or U12159 (N_12159,N_11942,N_11541);
nand U12160 (N_12160,N_11128,N_11621);
and U12161 (N_12161,N_11196,N_11880);
xnor U12162 (N_12162,N_10519,N_11622);
or U12163 (N_12163,N_10597,N_11896);
nor U12164 (N_12164,N_11407,N_11528);
nand U12165 (N_12165,N_10591,N_11756);
nor U12166 (N_12166,N_11350,N_11802);
nor U12167 (N_12167,N_11428,N_11553);
or U12168 (N_12168,N_11435,N_11805);
xnor U12169 (N_12169,N_10769,N_11778);
and U12170 (N_12170,N_11002,N_11182);
or U12171 (N_12171,N_10760,N_11691);
and U12172 (N_12172,N_10906,N_11723);
nand U12173 (N_12173,N_11818,N_10890);
and U12174 (N_12174,N_11945,N_10790);
nor U12175 (N_12175,N_11249,N_10956);
nand U12176 (N_12176,N_11226,N_11596);
or U12177 (N_12177,N_11148,N_11167);
or U12178 (N_12178,N_10856,N_10555);
or U12179 (N_12179,N_10654,N_11672);
xnor U12180 (N_12180,N_11892,N_10775);
and U12181 (N_12181,N_11054,N_11434);
nor U12182 (N_12182,N_11216,N_10968);
and U12183 (N_12183,N_11879,N_11813);
and U12184 (N_12184,N_10662,N_10537);
xnor U12185 (N_12185,N_11150,N_10811);
nor U12186 (N_12186,N_11565,N_10847);
xnor U12187 (N_12187,N_11848,N_11013);
nand U12188 (N_12188,N_11636,N_11383);
nand U12189 (N_12189,N_10726,N_11490);
nand U12190 (N_12190,N_11201,N_11796);
xor U12191 (N_12191,N_11272,N_11567);
nor U12192 (N_12192,N_11983,N_11969);
nor U12193 (N_12193,N_10960,N_11126);
nor U12194 (N_12194,N_10684,N_11546);
nand U12195 (N_12195,N_10807,N_11004);
nor U12196 (N_12196,N_11960,N_11845);
xnor U12197 (N_12197,N_10959,N_11509);
xor U12198 (N_12198,N_10528,N_10576);
nor U12199 (N_12199,N_10893,N_11590);
nand U12200 (N_12200,N_11837,N_11169);
or U12201 (N_12201,N_10566,N_11889);
and U12202 (N_12202,N_11968,N_10665);
and U12203 (N_12203,N_10535,N_10727);
and U12204 (N_12204,N_10802,N_10663);
or U12205 (N_12205,N_11097,N_10728);
or U12206 (N_12206,N_11442,N_10866);
nand U12207 (N_12207,N_10773,N_11325);
nor U12208 (N_12208,N_10522,N_11888);
and U12209 (N_12209,N_10864,N_10669);
nor U12210 (N_12210,N_11422,N_11849);
and U12211 (N_12211,N_11312,N_10998);
nor U12212 (N_12212,N_11195,N_11763);
or U12213 (N_12213,N_11686,N_11822);
nor U12214 (N_12214,N_11424,N_11478);
nor U12215 (N_12215,N_10637,N_11252);
nand U12216 (N_12216,N_11380,N_11016);
or U12217 (N_12217,N_10652,N_10643);
nand U12218 (N_12218,N_10737,N_10942);
xnor U12219 (N_12219,N_11874,N_11730);
nand U12220 (N_12220,N_11524,N_11116);
nand U12221 (N_12221,N_10912,N_11467);
and U12222 (N_12222,N_11704,N_10512);
or U12223 (N_12223,N_10816,N_11693);
nor U12224 (N_12224,N_11053,N_10534);
and U12225 (N_12225,N_10982,N_10585);
xor U12226 (N_12226,N_11790,N_10544);
xor U12227 (N_12227,N_11178,N_11299);
or U12228 (N_12228,N_10592,N_11953);
or U12229 (N_12229,N_10804,N_11365);
nor U12230 (N_12230,N_10657,N_11610);
nand U12231 (N_12231,N_10943,N_10753);
xor U12232 (N_12232,N_11374,N_10806);
and U12233 (N_12233,N_11076,N_10937);
nand U12234 (N_12234,N_11538,N_11307);
nor U12235 (N_12235,N_11502,N_11808);
and U12236 (N_12236,N_11554,N_11760);
or U12237 (N_12237,N_10543,N_10783);
xor U12238 (N_12238,N_10999,N_11617);
and U12239 (N_12239,N_10885,N_11507);
nor U12240 (N_12240,N_11371,N_11505);
nor U12241 (N_12241,N_11512,N_10572);
and U12242 (N_12242,N_11771,N_11300);
or U12243 (N_12243,N_11191,N_11175);
nand U12244 (N_12244,N_10900,N_11401);
xor U12245 (N_12245,N_10724,N_11940);
nand U12246 (N_12246,N_11078,N_11917);
and U12247 (N_12247,N_10651,N_11747);
or U12248 (N_12248,N_10836,N_10945);
or U12249 (N_12249,N_10896,N_11572);
or U12250 (N_12250,N_10701,N_10635);
or U12251 (N_12251,N_11035,N_10629);
nand U12252 (N_12252,N_11753,N_11902);
and U12253 (N_12253,N_11444,N_11278);
or U12254 (N_12254,N_11911,N_11998);
xnor U12255 (N_12255,N_10579,N_11064);
or U12256 (N_12256,N_11347,N_10723);
nor U12257 (N_12257,N_10653,N_11402);
or U12258 (N_12258,N_11800,N_10800);
or U12259 (N_12259,N_10719,N_10827);
xor U12260 (N_12260,N_10803,N_10764);
or U12261 (N_12261,N_11472,N_10870);
nor U12262 (N_12262,N_10608,N_11448);
nand U12263 (N_12263,N_11678,N_11454);
nor U12264 (N_12264,N_11729,N_11877);
xor U12265 (N_12265,N_11222,N_10888);
or U12266 (N_12266,N_11270,N_11992);
or U12267 (N_12267,N_11243,N_10696);
xor U12268 (N_12268,N_10715,N_11337);
nand U12269 (N_12269,N_10621,N_10939);
xor U12270 (N_12270,N_10685,N_11117);
and U12271 (N_12271,N_11732,N_11801);
xnor U12272 (N_12272,N_11803,N_11342);
or U12273 (N_12273,N_11749,N_11684);
nand U12274 (N_12274,N_11388,N_11863);
nor U12275 (N_12275,N_10704,N_11345);
nor U12276 (N_12276,N_11851,N_11591);
nor U12277 (N_12277,N_10521,N_10840);
and U12278 (N_12278,N_11535,N_10527);
or U12279 (N_12279,N_11060,N_10695);
nand U12280 (N_12280,N_11480,N_11240);
and U12281 (N_12281,N_10823,N_10545);
nor U12282 (N_12282,N_11934,N_11578);
xnor U12283 (N_12283,N_10569,N_11931);
and U12284 (N_12284,N_11247,N_11623);
nand U12285 (N_12285,N_11313,N_11066);
nor U12286 (N_12286,N_10613,N_10754);
nor U12287 (N_12287,N_10553,N_11458);
nor U12288 (N_12288,N_11533,N_10897);
nor U12289 (N_12289,N_11329,N_11844);
and U12290 (N_12290,N_11850,N_11009);
xor U12291 (N_12291,N_11823,N_11018);
or U12292 (N_12292,N_11552,N_11384);
or U12293 (N_12293,N_11599,N_11296);
or U12294 (N_12294,N_11608,N_11532);
and U12295 (N_12295,N_11894,N_11486);
nand U12296 (N_12296,N_10639,N_11971);
xnor U12297 (N_12297,N_11146,N_11755);
xnor U12298 (N_12298,N_11156,N_10722);
and U12299 (N_12299,N_11042,N_11557);
or U12300 (N_12300,N_11716,N_11555);
or U12301 (N_12301,N_11318,N_11959);
or U12302 (N_12302,N_10946,N_11841);
or U12303 (N_12303,N_11708,N_11843);
nand U12304 (N_12304,N_11031,N_10933);
or U12305 (N_12305,N_10821,N_11735);
and U12306 (N_12306,N_10913,N_11881);
nor U12307 (N_12307,N_11666,N_11269);
and U12308 (N_12308,N_11032,N_11926);
nand U12309 (N_12309,N_11068,N_11946);
and U12310 (N_12310,N_11504,N_11138);
nor U12311 (N_12311,N_11812,N_11862);
or U12312 (N_12312,N_10992,N_11981);
nor U12313 (N_12313,N_11688,N_11935);
nand U12314 (N_12314,N_10604,N_11702);
or U12315 (N_12315,N_10970,N_11262);
nor U12316 (N_12316,N_11125,N_11694);
or U12317 (N_12317,N_11280,N_11773);
and U12318 (N_12318,N_10648,N_11611);
nand U12319 (N_12319,N_11202,N_11692);
xor U12320 (N_12320,N_10832,N_10857);
and U12321 (N_12321,N_11542,N_11246);
nand U12322 (N_12322,N_10707,N_10772);
and U12323 (N_12323,N_10666,N_11606);
or U12324 (N_12324,N_11906,N_10603);
and U12325 (N_12325,N_11241,N_10556);
xnor U12326 (N_12326,N_11867,N_10837);
or U12327 (N_12327,N_11754,N_10718);
nor U12328 (N_12328,N_10618,N_11348);
nor U12329 (N_12329,N_10647,N_11127);
and U12330 (N_12330,N_10758,N_10690);
xnor U12331 (N_12331,N_11776,N_11515);
or U12332 (N_12332,N_11814,N_10561);
or U12333 (N_12333,N_10688,N_10577);
and U12334 (N_12334,N_11989,N_11639);
xor U12335 (N_12335,N_11909,N_10686);
and U12336 (N_12336,N_11123,N_11273);
nor U12337 (N_12337,N_11235,N_11140);
or U12338 (N_12338,N_10786,N_11717);
nand U12339 (N_12339,N_10928,N_11183);
nand U12340 (N_12340,N_11643,N_10744);
and U12341 (N_12341,N_11709,N_10776);
or U12342 (N_12342,N_11029,N_11767);
nand U12343 (N_12343,N_11508,N_11338);
nand U12344 (N_12344,N_10770,N_11679);
and U12345 (N_12345,N_11310,N_11830);
or U12346 (N_12346,N_11758,N_11775);
nand U12347 (N_12347,N_10619,N_11624);
nand U12348 (N_12348,N_11914,N_11733);
nor U12349 (N_12349,N_10642,N_10972);
xnor U12350 (N_12350,N_11236,N_11918);
or U12351 (N_12351,N_11696,N_11661);
and U12352 (N_12352,N_10680,N_11768);
xor U12353 (N_12353,N_11030,N_11683);
nand U12354 (N_12354,N_11965,N_11357);
xor U12355 (N_12355,N_10996,N_10710);
nor U12356 (N_12356,N_11098,N_11972);
or U12357 (N_12357,N_11901,N_11274);
and U12358 (N_12358,N_10833,N_11447);
and U12359 (N_12359,N_10574,N_10902);
or U12360 (N_12360,N_11011,N_10971);
nand U12361 (N_12361,N_10986,N_11144);
xor U12362 (N_12362,N_11427,N_11494);
nor U12363 (N_12363,N_11811,N_10713);
nor U12364 (N_12364,N_10988,N_10925);
or U12365 (N_12365,N_11842,N_10991);
or U12366 (N_12366,N_11868,N_10974);
or U12367 (N_12367,N_11807,N_10712);
xor U12368 (N_12368,N_11019,N_10984);
nand U12369 (N_12369,N_11199,N_11369);
nand U12370 (N_12370,N_11872,N_10766);
or U12371 (N_12371,N_11321,N_10761);
and U12372 (N_12372,N_10855,N_11170);
xor U12373 (N_12373,N_11143,N_11366);
and U12374 (N_12374,N_11142,N_10539);
nor U12375 (N_12375,N_11618,N_11319);
or U12376 (N_12376,N_10625,N_10862);
nor U12377 (N_12377,N_10734,N_11131);
nor U12378 (N_12378,N_11197,N_10835);
nand U12379 (N_12379,N_10748,N_11517);
and U12380 (N_12380,N_11231,N_10646);
nand U12381 (N_12381,N_10848,N_11766);
and U12382 (N_12382,N_11609,N_11387);
or U12383 (N_12383,N_11121,N_11451);
nand U12384 (N_12384,N_11025,N_11057);
and U12385 (N_12385,N_10830,N_11548);
xnor U12386 (N_12386,N_11676,N_11049);
nor U12387 (N_12387,N_11001,N_11589);
nor U12388 (N_12388,N_11364,N_11663);
nand U12389 (N_12389,N_10575,N_11266);
nor U12390 (N_12390,N_10557,N_11339);
or U12391 (N_12391,N_11297,N_11860);
nand U12392 (N_12392,N_11764,N_10841);
xor U12393 (N_12393,N_10668,N_11562);
and U12394 (N_12394,N_11726,N_10796);
xnor U12395 (N_12395,N_11491,N_11124);
and U12396 (N_12396,N_10973,N_11828);
or U12397 (N_12397,N_10584,N_11174);
nor U12398 (N_12398,N_11284,N_11597);
xor U12399 (N_12399,N_11660,N_10780);
nor U12400 (N_12400,N_11795,N_11545);
and U12401 (N_12401,N_10911,N_10703);
nor U12402 (N_12402,N_11354,N_11211);
or U12403 (N_12403,N_11024,N_10736);
nand U12404 (N_12404,N_10898,N_11477);
or U12405 (N_12405,N_11159,N_10849);
or U12406 (N_12406,N_10508,N_10781);
nor U12407 (N_12407,N_11224,N_11411);
and U12408 (N_12408,N_10593,N_11089);
nor U12409 (N_12409,N_10809,N_11227);
nand U12410 (N_12410,N_11997,N_10743);
nand U12411 (N_12411,N_11878,N_11283);
xnor U12412 (N_12412,N_11543,N_11405);
nor U12413 (N_12413,N_11014,N_11152);
or U12414 (N_12414,N_11870,N_11705);
or U12415 (N_12415,N_11379,N_11592);
or U12416 (N_12416,N_11286,N_10670);
xnor U12417 (N_12417,N_11306,N_10923);
nand U12418 (N_12418,N_11415,N_11527);
nand U12419 (N_12419,N_11056,N_11218);
nor U12420 (N_12420,N_10975,N_11356);
and U12421 (N_12421,N_11765,N_11503);
nor U12422 (N_12422,N_11628,N_10532);
or U12423 (N_12423,N_10768,N_11722);
xnor U12424 (N_12424,N_10554,N_11094);
and U12425 (N_12425,N_11463,N_10903);
xor U12426 (N_12426,N_11866,N_10716);
xnor U12427 (N_12427,N_11239,N_10978);
xnor U12428 (N_12428,N_10910,N_11457);
nand U12429 (N_12429,N_10799,N_10794);
and U12430 (N_12430,N_10947,N_10706);
and U12431 (N_12431,N_10573,N_11403);
nand U12432 (N_12432,N_11087,N_11186);
xor U12433 (N_12433,N_11203,N_11000);
and U12434 (N_12434,N_11654,N_11255);
or U12435 (N_12435,N_11682,N_10721);
or U12436 (N_12436,N_10810,N_11441);
nor U12437 (N_12437,N_10697,N_10623);
and U12438 (N_12438,N_11122,N_11194);
xor U12439 (N_12439,N_11882,N_10626);
nor U12440 (N_12440,N_10808,N_10795);
nor U12441 (N_12441,N_11938,N_11220);
or U12442 (N_12442,N_11230,N_11738);
xor U12443 (N_12443,N_10877,N_11530);
nor U12444 (N_12444,N_10622,N_10931);
xor U12445 (N_12445,N_11119,N_11644);
nor U12446 (N_12446,N_10587,N_11687);
and U12447 (N_12447,N_10788,N_11052);
and U12448 (N_12448,N_11080,N_11593);
and U12449 (N_12449,N_11245,N_11292);
and U12450 (N_12450,N_11482,N_11264);
xor U12451 (N_12451,N_11038,N_10676);
and U12452 (N_12452,N_10526,N_11824);
nand U12453 (N_12453,N_10739,N_11995);
and U12454 (N_12454,N_10546,N_11697);
nand U12455 (N_12455,N_11794,N_11416);
and U12456 (N_12456,N_11988,N_11440);
nand U12457 (N_12457,N_11962,N_10562);
or U12458 (N_12458,N_10507,N_10506);
nor U12459 (N_12459,N_11392,N_11426);
xor U12460 (N_12460,N_10700,N_10656);
or U12461 (N_12461,N_11396,N_10831);
and U12462 (N_12462,N_11852,N_11061);
nor U12463 (N_12463,N_10568,N_11832);
or U12464 (N_12464,N_10571,N_10580);
nand U12465 (N_12465,N_10709,N_11581);
nor U12466 (N_12466,N_11389,N_10778);
and U12467 (N_12467,N_11349,N_11012);
nand U12468 (N_12468,N_10891,N_10541);
and U12469 (N_12469,N_10963,N_11884);
and U12470 (N_12470,N_11244,N_11027);
xnor U12471 (N_12471,N_10845,N_10958);
nor U12472 (N_12472,N_11784,N_11690);
nand U12473 (N_12473,N_11650,N_11577);
nor U12474 (N_12474,N_11437,N_10976);
and U12475 (N_12475,N_10596,N_11190);
or U12476 (N_12476,N_10746,N_10784);
nor U12477 (N_12477,N_11826,N_10792);
and U12478 (N_12478,N_11903,N_10505);
and U12479 (N_12479,N_11761,N_11919);
or U12480 (N_12480,N_11947,N_11465);
and U12481 (N_12481,N_10549,N_10523);
or U12482 (N_12482,N_11662,N_11804);
or U12483 (N_12483,N_11084,N_11523);
nor U12484 (N_12484,N_11652,N_10895);
and U12485 (N_12485,N_11928,N_11293);
or U12486 (N_12486,N_11655,N_10985);
nor U12487 (N_12487,N_11810,N_11759);
nor U12488 (N_12488,N_10691,N_11205);
and U12489 (N_12489,N_11008,N_11785);
nand U12490 (N_12490,N_10518,N_11659);
nand U12491 (N_12491,N_10542,N_10717);
or U12492 (N_12492,N_11277,N_10560);
nor U12493 (N_12493,N_11139,N_11096);
nor U12494 (N_12494,N_10567,N_11433);
xor U12495 (N_12495,N_11781,N_11335);
nor U12496 (N_12496,N_11176,N_11317);
nand U12497 (N_12497,N_11556,N_10901);
nor U12498 (N_12498,N_10698,N_11036);
nand U12499 (N_12499,N_11091,N_11956);
xor U12500 (N_12500,N_11332,N_10738);
nor U12501 (N_12501,N_10607,N_10842);
and U12502 (N_12502,N_11021,N_11481);
nor U12503 (N_12503,N_10605,N_11620);
nand U12504 (N_12504,N_11301,N_11551);
nand U12505 (N_12505,N_11311,N_11951);
nand U12506 (N_12506,N_11083,N_11303);
or U12507 (N_12507,N_10513,N_11265);
and U12508 (N_12508,N_11470,N_11304);
and U12509 (N_12509,N_10540,N_11887);
nand U12510 (N_12510,N_11275,N_10797);
and U12511 (N_12511,N_11104,N_11041);
nor U12512 (N_12512,N_10500,N_11875);
or U12513 (N_12513,N_11518,N_11993);
xor U12514 (N_12514,N_11160,N_11898);
or U12515 (N_12515,N_11157,N_11063);
nor U12516 (N_12516,N_10732,N_11966);
and U12517 (N_12517,N_11375,N_11314);
xor U12518 (N_12518,N_11734,N_10747);
nand U12519 (N_12519,N_10750,N_11103);
and U12520 (N_12520,N_11215,N_10529);
and U12521 (N_12521,N_10524,N_10601);
or U12522 (N_12522,N_10672,N_11399);
xnor U12523 (N_12523,N_10589,N_10708);
xnor U12524 (N_12524,N_10617,N_11908);
nor U12525 (N_12525,N_11600,N_11315);
xnor U12526 (N_12526,N_11924,N_11932);
xor U12527 (N_12527,N_10872,N_11471);
nor U12528 (N_12528,N_11825,N_10953);
or U12529 (N_12529,N_10957,N_11582);
nand U12530 (N_12530,N_11489,N_11646);
or U12531 (N_12531,N_11757,N_11724);
nand U12532 (N_12532,N_11865,N_10725);
nor U12533 (N_12533,N_10820,N_11268);
nand U12534 (N_12534,N_11419,N_11343);
nor U12535 (N_12535,N_10742,N_11322);
nand U12536 (N_12536,N_11015,N_11640);
xor U12537 (N_12537,N_11566,N_11913);
and U12538 (N_12538,N_10740,N_10774);
nor U12539 (N_12539,N_11789,N_11673);
or U12540 (N_12540,N_10882,N_10550);
nor U12541 (N_12541,N_11185,N_11500);
nand U12542 (N_12542,N_11294,N_11113);
nand U12543 (N_12543,N_11291,N_10645);
nand U12544 (N_12544,N_11740,N_10791);
nor U12545 (N_12545,N_10520,N_11665);
and U12546 (N_12546,N_11718,N_10995);
and U12547 (N_12547,N_10659,N_10952);
and U12548 (N_12548,N_11109,N_10899);
nand U12549 (N_12549,N_11137,N_10515);
nor U12550 (N_12550,N_11147,N_10904);
nor U12551 (N_12551,N_10615,N_11978);
nor U12552 (N_12552,N_11531,N_10547);
nor U12553 (N_12553,N_10983,N_11223);
xnor U12554 (N_12554,N_11151,N_11635);
nand U12555 (N_12555,N_10628,N_11498);
and U12556 (N_12556,N_11575,N_10859);
or U12557 (N_12557,N_10711,N_10745);
xor U12558 (N_12558,N_11111,N_11429);
nand U12559 (N_12559,N_10570,N_11891);
nor U12560 (N_12560,N_11750,N_10614);
and U12561 (N_12561,N_11806,N_11381);
or U12562 (N_12562,N_10918,N_10940);
nor U12563 (N_12563,N_11958,N_11006);
nor U12564 (N_12564,N_11669,N_10861);
xnor U12565 (N_12565,N_11626,N_11910);
or U12566 (N_12566,N_10965,N_11588);
xor U12567 (N_12567,N_11809,N_10661);
or U12568 (N_12568,N_11077,N_11487);
and U12569 (N_12569,N_10682,N_11714);
nor U12570 (N_12570,N_10610,N_11853);
or U12571 (N_12571,N_10927,N_11017);
or U12572 (N_12572,N_11570,N_11050);
xor U12573 (N_12573,N_11385,N_11725);
nor U12574 (N_12574,N_10634,N_11954);
nor U12575 (N_12575,N_11177,N_11497);
nor U12576 (N_12576,N_11680,N_11601);
xnor U12577 (N_12577,N_10756,N_11739);
or U12578 (N_12578,N_11358,N_10997);
or U12579 (N_12579,N_11916,N_11393);
and U12580 (N_12580,N_11563,N_11290);
nand U12581 (N_12581,N_11250,N_10858);
and U12582 (N_12582,N_11333,N_11172);
and U12583 (N_12583,N_11922,N_11037);
nor U12584 (N_12584,N_11612,N_11907);
and U12585 (N_12585,N_11779,N_11657);
and U12586 (N_12586,N_11232,N_11658);
xnor U12587 (N_12587,N_11869,N_11483);
nor U12588 (N_12588,N_11028,N_11135);
and U12589 (N_12589,N_11641,N_11631);
xor U12590 (N_12590,N_10741,N_11436);
nor U12591 (N_12591,N_11840,N_10679);
or U12592 (N_12592,N_11074,N_10879);
xnor U12593 (N_12593,N_10916,N_10502);
or U12594 (N_12594,N_11782,N_10929);
and U12595 (N_12595,N_11368,N_11933);
nand U12596 (N_12596,N_10954,N_11929);
or U12597 (N_12597,N_10558,N_11949);
or U12598 (N_12598,N_10944,N_11257);
and U12599 (N_12599,N_11513,N_10798);
nand U12600 (N_12600,N_11602,N_11540);
and U12601 (N_12601,N_11957,N_11770);
xor U12602 (N_12602,N_11039,N_11937);
and U12603 (N_12603,N_10677,N_11468);
nand U12604 (N_12604,N_10655,N_11786);
or U12605 (N_12605,N_11204,N_11944);
nand U12606 (N_12606,N_11395,N_11912);
nor U12607 (N_12607,N_10812,N_10894);
xor U12608 (N_12608,N_11970,N_11838);
or U12609 (N_12609,N_11677,N_11400);
xor U12610 (N_12610,N_11281,N_11130);
xnor U12611 (N_12611,N_11086,N_11234);
and U12612 (N_12612,N_11817,N_10609);
and U12613 (N_12613,N_10951,N_11999);
nor U12614 (N_12614,N_11259,N_11576);
nor U12615 (N_12615,N_10860,N_11180);
xor U12616 (N_12616,N_10914,N_10678);
and U12617 (N_12617,N_10649,N_11569);
and U12618 (N_12618,N_10852,N_11071);
and U12619 (N_12619,N_11154,N_11048);
nand U12620 (N_12620,N_11619,N_10720);
and U12621 (N_12621,N_11746,N_11560);
or U12622 (N_12622,N_11248,N_11516);
nor U12623 (N_12623,N_11344,N_10509);
nand U12624 (N_12624,N_11188,N_10687);
nand U12625 (N_12625,N_11973,N_10694);
xor U12626 (N_12626,N_11221,N_10878);
nand U12627 (N_12627,N_11258,N_11316);
and U12628 (N_12628,N_10702,N_11706);
xor U12629 (N_12629,N_10681,N_11324);
or U12630 (N_12630,N_11079,N_10536);
nand U12631 (N_12631,N_11102,N_11118);
nor U12632 (N_12632,N_11996,N_11065);
nand U12633 (N_12633,N_10510,N_11864);
or U12634 (N_12634,N_10749,N_10892);
or U12635 (N_12635,N_10501,N_11629);
xor U12636 (N_12636,N_10990,N_11242);
xor U12637 (N_12637,N_11955,N_11584);
xor U12638 (N_12638,N_11261,N_11948);
or U12639 (N_12639,N_10819,N_11967);
xnor U12640 (N_12640,N_11173,N_10961);
and U12641 (N_12641,N_11846,N_11941);
nand U12642 (N_12642,N_11651,N_11453);
nor U12643 (N_12643,N_11040,N_11367);
or U12644 (N_12644,N_11506,N_11703);
nor U12645 (N_12645,N_10881,N_11583);
xor U12646 (N_12646,N_11943,N_10731);
or U12647 (N_12647,N_11990,N_11791);
xor U12648 (N_12648,N_11925,N_11398);
or U12649 (N_12649,N_11886,N_11179);
nand U12650 (N_12650,N_11815,N_11613);
nand U12651 (N_12651,N_10590,N_11568);
nor U12652 (N_12652,N_11373,N_11145);
or U12653 (N_12653,N_11752,N_10787);
nor U12654 (N_12654,N_11340,N_11719);
nor U12655 (N_12655,N_11831,N_11648);
xor U12656 (N_12656,N_11536,N_11484);
xor U12657 (N_12657,N_10932,N_10938);
nor U12658 (N_12658,N_10924,N_11047);
and U12659 (N_12659,N_11168,N_10789);
nor U12660 (N_12660,N_11964,N_11649);
or U12661 (N_12661,N_11431,N_10636);
xnor U12662 (N_12662,N_11743,N_11748);
xor U12663 (N_12663,N_11372,N_10595);
or U12664 (N_12664,N_11522,N_11206);
or U12665 (N_12665,N_10887,N_11210);
xor U12666 (N_12666,N_11153,N_11282);
nand U12667 (N_12667,N_10994,N_11081);
and U12668 (N_12668,N_10886,N_11473);
nand U12669 (N_12669,N_10675,N_11493);
and U12670 (N_12670,N_11377,N_11100);
and U12671 (N_12671,N_10671,N_11408);
or U12672 (N_12672,N_10981,N_11287);
and U12673 (N_12673,N_10979,N_11939);
or U12674 (N_12674,N_10950,N_11412);
or U12675 (N_12675,N_10578,N_10908);
and U12676 (N_12676,N_11162,N_11106);
nand U12677 (N_12677,N_11675,N_11233);
xnor U12678 (N_12678,N_11263,N_10926);
and U12679 (N_12679,N_10844,N_10627);
nor U12680 (N_12680,N_11689,N_11783);
xnor U12681 (N_12681,N_11295,N_11352);
and U12682 (N_12682,N_10551,N_11141);
xnor U12683 (N_12683,N_11459,N_11417);
xor U12684 (N_12684,N_11438,N_11904);
and U12685 (N_12685,N_11607,N_11165);
nor U12686 (N_12686,N_11209,N_10935);
or U12687 (N_12687,N_10863,N_11410);
nor U12688 (N_12688,N_11044,N_11559);
nor U12689 (N_12689,N_10599,N_10955);
nand U12690 (N_12690,N_11751,N_11390);
and U12691 (N_12691,N_11225,N_11432);
xor U12692 (N_12692,N_11213,N_11741);
xor U12693 (N_12693,N_11394,N_10875);
nand U12694 (N_12694,N_10969,N_10966);
or U12695 (N_12695,N_11987,N_11161);
and U12696 (N_12696,N_11647,N_11466);
nor U12697 (N_12697,N_10868,N_11616);
or U12698 (N_12698,N_11187,N_11088);
xnor U12699 (N_12699,N_10563,N_10853);
or U12700 (N_12700,N_11046,N_10921);
and U12701 (N_12701,N_10752,N_11816);
nand U12702 (N_12702,N_11062,N_11166);
and U12703 (N_12703,N_11189,N_10658);
nor U12704 (N_12704,N_11854,N_10989);
nor U12705 (N_12705,N_10980,N_10616);
nand U12706 (N_12706,N_11985,N_11627);
xor U12707 (N_12707,N_10582,N_10586);
nor U12708 (N_12708,N_11105,N_11900);
xor U12709 (N_12709,N_10909,N_10644);
or U12710 (N_12710,N_10967,N_11587);
nor U12711 (N_12711,N_10962,N_11254);
or U12712 (N_12712,N_11378,N_11085);
and U12713 (N_12713,N_11710,N_11698);
and U12714 (N_12714,N_10846,N_10533);
xnor U12715 (N_12715,N_11461,N_10733);
or U12716 (N_12716,N_11133,N_10612);
or U12717 (N_12717,N_11634,N_11982);
or U12718 (N_12718,N_11899,N_11360);
or U12719 (N_12719,N_10825,N_11858);
nor U12720 (N_12720,N_11859,N_10751);
or U12721 (N_12721,N_10850,N_10755);
and U12722 (N_12722,N_11193,N_10828);
nand U12723 (N_12723,N_11897,N_11975);
and U12724 (N_12724,N_11769,N_10987);
and U12725 (N_12725,N_10650,N_11798);
nand U12726 (N_12726,N_11774,N_11742);
nand U12727 (N_12727,N_11149,N_11549);
xnor U12728 (N_12728,N_11474,N_10641);
nand U12729 (N_12729,N_11108,N_11120);
xnor U12730 (N_12730,N_10993,N_10948);
xor U12731 (N_12731,N_11715,N_11058);
and U12732 (N_12732,N_11977,N_11656);
and U12733 (N_12733,N_11010,N_10785);
nor U12734 (N_12734,N_10782,N_11829);
or U12735 (N_12735,N_11707,N_11237);
or U12736 (N_12736,N_11920,N_11418);
and U12737 (N_12737,N_10548,N_10638);
nand U12738 (N_12738,N_10640,N_11302);
or U12739 (N_12739,N_11101,N_10530);
and U12740 (N_12740,N_11192,N_10763);
xnor U12741 (N_12741,N_11630,N_11112);
nand U12742 (N_12742,N_11055,N_11885);
nor U12743 (N_12743,N_11443,N_11279);
and U12744 (N_12744,N_11425,N_11351);
xnor U12745 (N_12745,N_11604,N_11625);
or U12746 (N_12746,N_11238,N_11456);
or U12747 (N_12747,N_11574,N_11564);
xnor U12748 (N_12748,N_11499,N_10516);
xnor U12749 (N_12749,N_11134,N_11409);
nand U12750 (N_12750,N_11633,N_11911);
xor U12751 (N_12751,N_11981,N_11635);
and U12752 (N_12752,N_11491,N_10825);
or U12753 (N_12753,N_10957,N_11197);
xor U12754 (N_12754,N_10987,N_11300);
xnor U12755 (N_12755,N_10937,N_11584);
nand U12756 (N_12756,N_11917,N_11169);
nor U12757 (N_12757,N_11743,N_11333);
nand U12758 (N_12758,N_11352,N_11798);
xor U12759 (N_12759,N_11948,N_11725);
nand U12760 (N_12760,N_10649,N_11763);
nor U12761 (N_12761,N_11512,N_11157);
nor U12762 (N_12762,N_11348,N_11825);
nor U12763 (N_12763,N_11371,N_11231);
nor U12764 (N_12764,N_11894,N_10713);
or U12765 (N_12765,N_10642,N_10980);
nor U12766 (N_12766,N_11713,N_11144);
nand U12767 (N_12767,N_10700,N_11789);
nor U12768 (N_12768,N_11375,N_10883);
and U12769 (N_12769,N_10523,N_11747);
nor U12770 (N_12770,N_10749,N_10509);
and U12771 (N_12771,N_10979,N_11005);
and U12772 (N_12772,N_11855,N_11885);
or U12773 (N_12773,N_10845,N_11723);
xor U12774 (N_12774,N_11457,N_11922);
nand U12775 (N_12775,N_11790,N_10831);
and U12776 (N_12776,N_11530,N_11918);
nor U12777 (N_12777,N_10796,N_11192);
xnor U12778 (N_12778,N_10668,N_10854);
nor U12779 (N_12779,N_11966,N_11253);
nor U12780 (N_12780,N_11089,N_11267);
xor U12781 (N_12781,N_11276,N_11988);
or U12782 (N_12782,N_11265,N_11836);
nand U12783 (N_12783,N_11743,N_11118);
nand U12784 (N_12784,N_11991,N_11483);
and U12785 (N_12785,N_11205,N_11007);
nor U12786 (N_12786,N_11031,N_10676);
xor U12787 (N_12787,N_11070,N_11587);
xnor U12788 (N_12788,N_11086,N_11639);
nor U12789 (N_12789,N_11409,N_10543);
nor U12790 (N_12790,N_11745,N_10546);
nand U12791 (N_12791,N_10579,N_11544);
or U12792 (N_12792,N_11941,N_10905);
and U12793 (N_12793,N_11204,N_11842);
and U12794 (N_12794,N_11158,N_11922);
nand U12795 (N_12795,N_10970,N_11129);
xnor U12796 (N_12796,N_11767,N_11243);
and U12797 (N_12797,N_10941,N_11176);
nor U12798 (N_12798,N_11026,N_11728);
xor U12799 (N_12799,N_10816,N_11482);
nand U12800 (N_12800,N_11363,N_11721);
nor U12801 (N_12801,N_11249,N_10659);
nand U12802 (N_12802,N_10742,N_11528);
or U12803 (N_12803,N_10863,N_10677);
xor U12804 (N_12804,N_11438,N_11391);
nor U12805 (N_12805,N_11135,N_10578);
and U12806 (N_12806,N_11593,N_11009);
nand U12807 (N_12807,N_11548,N_10534);
or U12808 (N_12808,N_10699,N_10918);
and U12809 (N_12809,N_11065,N_11219);
nand U12810 (N_12810,N_11413,N_11683);
or U12811 (N_12811,N_11704,N_10646);
xor U12812 (N_12812,N_11952,N_10671);
or U12813 (N_12813,N_11838,N_11507);
or U12814 (N_12814,N_11112,N_11828);
nor U12815 (N_12815,N_11852,N_11977);
and U12816 (N_12816,N_11612,N_11453);
nor U12817 (N_12817,N_11779,N_11182);
nor U12818 (N_12818,N_10869,N_10949);
xor U12819 (N_12819,N_11742,N_10861);
nor U12820 (N_12820,N_10814,N_10727);
xor U12821 (N_12821,N_10619,N_11894);
or U12822 (N_12822,N_10604,N_11205);
nor U12823 (N_12823,N_10581,N_11148);
nand U12824 (N_12824,N_11029,N_10606);
nand U12825 (N_12825,N_11658,N_11681);
nor U12826 (N_12826,N_11133,N_11565);
or U12827 (N_12827,N_11389,N_11757);
and U12828 (N_12828,N_11273,N_11488);
and U12829 (N_12829,N_11219,N_10900);
xnor U12830 (N_12830,N_11121,N_10921);
xnor U12831 (N_12831,N_11729,N_11854);
and U12832 (N_12832,N_11493,N_11944);
nand U12833 (N_12833,N_10757,N_11436);
and U12834 (N_12834,N_11421,N_10945);
or U12835 (N_12835,N_11351,N_11977);
or U12836 (N_12836,N_11838,N_11082);
or U12837 (N_12837,N_11545,N_11247);
nand U12838 (N_12838,N_11228,N_11726);
or U12839 (N_12839,N_10876,N_11505);
or U12840 (N_12840,N_11832,N_11582);
xor U12841 (N_12841,N_10835,N_11131);
nor U12842 (N_12842,N_11852,N_11578);
or U12843 (N_12843,N_11492,N_11809);
nor U12844 (N_12844,N_11842,N_11872);
and U12845 (N_12845,N_11726,N_11981);
nor U12846 (N_12846,N_11700,N_11813);
xnor U12847 (N_12847,N_11091,N_10595);
xnor U12848 (N_12848,N_10838,N_11404);
or U12849 (N_12849,N_11160,N_11678);
xor U12850 (N_12850,N_11855,N_11589);
and U12851 (N_12851,N_11423,N_11240);
nand U12852 (N_12852,N_10587,N_11163);
and U12853 (N_12853,N_11093,N_10851);
and U12854 (N_12854,N_10565,N_10648);
or U12855 (N_12855,N_10857,N_10542);
nand U12856 (N_12856,N_11506,N_10854);
nor U12857 (N_12857,N_11631,N_11208);
and U12858 (N_12858,N_11460,N_11200);
nor U12859 (N_12859,N_11170,N_11652);
or U12860 (N_12860,N_11405,N_10733);
nor U12861 (N_12861,N_11923,N_10885);
nor U12862 (N_12862,N_11313,N_11341);
xnor U12863 (N_12863,N_11538,N_10890);
nor U12864 (N_12864,N_11669,N_10530);
xnor U12865 (N_12865,N_11283,N_11111);
nand U12866 (N_12866,N_10906,N_11859);
and U12867 (N_12867,N_10741,N_11075);
and U12868 (N_12868,N_11595,N_11615);
and U12869 (N_12869,N_10687,N_10979);
nor U12870 (N_12870,N_11954,N_10604);
or U12871 (N_12871,N_11775,N_11301);
or U12872 (N_12872,N_10583,N_10776);
or U12873 (N_12873,N_11767,N_10803);
nand U12874 (N_12874,N_11540,N_11229);
nand U12875 (N_12875,N_11079,N_11518);
xor U12876 (N_12876,N_11884,N_11787);
nor U12877 (N_12877,N_11124,N_11600);
xnor U12878 (N_12878,N_11174,N_10675);
or U12879 (N_12879,N_11774,N_11757);
nor U12880 (N_12880,N_11793,N_10983);
and U12881 (N_12881,N_10580,N_11367);
nor U12882 (N_12882,N_11714,N_10591);
or U12883 (N_12883,N_10651,N_11608);
nor U12884 (N_12884,N_11580,N_10620);
nand U12885 (N_12885,N_11454,N_11235);
nor U12886 (N_12886,N_11108,N_10724);
nor U12887 (N_12887,N_10585,N_11985);
nor U12888 (N_12888,N_11799,N_11797);
xor U12889 (N_12889,N_11760,N_11067);
and U12890 (N_12890,N_11378,N_11811);
or U12891 (N_12891,N_11257,N_11122);
xnor U12892 (N_12892,N_11490,N_11809);
xnor U12893 (N_12893,N_11374,N_11996);
nand U12894 (N_12894,N_11460,N_11382);
and U12895 (N_12895,N_11217,N_10830);
nor U12896 (N_12896,N_10777,N_11967);
nand U12897 (N_12897,N_11730,N_10511);
or U12898 (N_12898,N_11584,N_11918);
nor U12899 (N_12899,N_10869,N_11320);
and U12900 (N_12900,N_10554,N_11482);
and U12901 (N_12901,N_10933,N_10759);
and U12902 (N_12902,N_10754,N_11092);
xor U12903 (N_12903,N_11293,N_11349);
xor U12904 (N_12904,N_10521,N_11637);
xor U12905 (N_12905,N_11409,N_10605);
nor U12906 (N_12906,N_11961,N_11600);
nand U12907 (N_12907,N_11552,N_10696);
and U12908 (N_12908,N_11886,N_11935);
and U12909 (N_12909,N_11508,N_10735);
and U12910 (N_12910,N_11564,N_11939);
and U12911 (N_12911,N_10585,N_10978);
nor U12912 (N_12912,N_11369,N_11964);
nor U12913 (N_12913,N_10674,N_11085);
and U12914 (N_12914,N_10985,N_11709);
or U12915 (N_12915,N_11072,N_11009);
nor U12916 (N_12916,N_11272,N_10524);
nand U12917 (N_12917,N_11140,N_11980);
nor U12918 (N_12918,N_11078,N_11451);
and U12919 (N_12919,N_11736,N_11279);
nand U12920 (N_12920,N_11907,N_11866);
and U12921 (N_12921,N_11066,N_10988);
and U12922 (N_12922,N_11013,N_11019);
nand U12923 (N_12923,N_11824,N_10583);
xnor U12924 (N_12924,N_10767,N_11653);
and U12925 (N_12925,N_11384,N_10649);
and U12926 (N_12926,N_11537,N_11620);
nand U12927 (N_12927,N_11117,N_10579);
or U12928 (N_12928,N_11343,N_10657);
or U12929 (N_12929,N_10906,N_10738);
nand U12930 (N_12930,N_10719,N_11714);
nand U12931 (N_12931,N_11984,N_11406);
nor U12932 (N_12932,N_10861,N_10982);
or U12933 (N_12933,N_11154,N_10978);
xor U12934 (N_12934,N_11692,N_11182);
nor U12935 (N_12935,N_11419,N_11944);
and U12936 (N_12936,N_11331,N_10894);
xnor U12937 (N_12937,N_10732,N_11951);
and U12938 (N_12938,N_10622,N_11337);
and U12939 (N_12939,N_11250,N_11130);
nand U12940 (N_12940,N_10699,N_11498);
and U12941 (N_12941,N_11732,N_11542);
nand U12942 (N_12942,N_10558,N_11101);
or U12943 (N_12943,N_10726,N_11516);
and U12944 (N_12944,N_11838,N_10842);
and U12945 (N_12945,N_10697,N_10607);
nor U12946 (N_12946,N_11576,N_10877);
or U12947 (N_12947,N_10699,N_11378);
nand U12948 (N_12948,N_11650,N_10590);
xnor U12949 (N_12949,N_11302,N_11610);
and U12950 (N_12950,N_11857,N_11015);
nor U12951 (N_12951,N_10986,N_10946);
and U12952 (N_12952,N_10543,N_11154);
xor U12953 (N_12953,N_11618,N_11742);
nand U12954 (N_12954,N_11586,N_11376);
and U12955 (N_12955,N_10673,N_11639);
or U12956 (N_12956,N_11040,N_11088);
xnor U12957 (N_12957,N_11724,N_10626);
xnor U12958 (N_12958,N_11745,N_11484);
and U12959 (N_12959,N_11837,N_11566);
nand U12960 (N_12960,N_10531,N_11297);
and U12961 (N_12961,N_10996,N_11891);
or U12962 (N_12962,N_11223,N_10859);
nor U12963 (N_12963,N_11444,N_11035);
nor U12964 (N_12964,N_11316,N_10971);
or U12965 (N_12965,N_11586,N_11258);
or U12966 (N_12966,N_11192,N_10797);
nand U12967 (N_12967,N_11105,N_11512);
or U12968 (N_12968,N_11038,N_10977);
xor U12969 (N_12969,N_11855,N_10775);
nor U12970 (N_12970,N_11172,N_10583);
and U12971 (N_12971,N_11620,N_10754);
nor U12972 (N_12972,N_10785,N_10770);
xnor U12973 (N_12973,N_10531,N_11890);
nor U12974 (N_12974,N_11070,N_11885);
nand U12975 (N_12975,N_10625,N_11784);
nand U12976 (N_12976,N_10933,N_10717);
and U12977 (N_12977,N_11754,N_11155);
nand U12978 (N_12978,N_11937,N_11357);
and U12979 (N_12979,N_11216,N_11922);
or U12980 (N_12980,N_10902,N_11045);
xor U12981 (N_12981,N_10763,N_11639);
and U12982 (N_12982,N_11469,N_10508);
xor U12983 (N_12983,N_11920,N_11189);
and U12984 (N_12984,N_10752,N_11441);
or U12985 (N_12985,N_11755,N_10913);
xnor U12986 (N_12986,N_11704,N_11239);
xor U12987 (N_12987,N_11282,N_10954);
and U12988 (N_12988,N_11601,N_11154);
nor U12989 (N_12989,N_11613,N_11088);
nand U12990 (N_12990,N_11850,N_11600);
and U12991 (N_12991,N_11132,N_10961);
xnor U12992 (N_12992,N_11607,N_10814);
nor U12993 (N_12993,N_11866,N_11574);
nand U12994 (N_12994,N_11025,N_10978);
or U12995 (N_12995,N_10606,N_11359);
or U12996 (N_12996,N_10631,N_11220);
nor U12997 (N_12997,N_11346,N_11015);
nand U12998 (N_12998,N_11999,N_10582);
xor U12999 (N_12999,N_11457,N_11565);
or U13000 (N_13000,N_10885,N_11560);
xnor U13001 (N_13001,N_11861,N_11997);
xnor U13002 (N_13002,N_10822,N_11989);
nand U13003 (N_13003,N_11379,N_10822);
and U13004 (N_13004,N_10937,N_11212);
xor U13005 (N_13005,N_10734,N_11242);
and U13006 (N_13006,N_11957,N_11594);
nand U13007 (N_13007,N_11777,N_11873);
xnor U13008 (N_13008,N_11224,N_10916);
nor U13009 (N_13009,N_11020,N_11808);
nor U13010 (N_13010,N_11744,N_11756);
or U13011 (N_13011,N_10697,N_11355);
or U13012 (N_13012,N_11963,N_11245);
and U13013 (N_13013,N_11857,N_10853);
nand U13014 (N_13014,N_10953,N_11269);
nand U13015 (N_13015,N_10661,N_11468);
xnor U13016 (N_13016,N_10938,N_11885);
nor U13017 (N_13017,N_10794,N_11404);
xor U13018 (N_13018,N_11433,N_10973);
nand U13019 (N_13019,N_11383,N_10896);
and U13020 (N_13020,N_11937,N_11233);
xor U13021 (N_13021,N_11566,N_11286);
nand U13022 (N_13022,N_10974,N_11083);
nor U13023 (N_13023,N_11640,N_11432);
xor U13024 (N_13024,N_11196,N_11282);
and U13025 (N_13025,N_11461,N_11062);
xor U13026 (N_13026,N_10827,N_11357);
nand U13027 (N_13027,N_11505,N_10849);
nor U13028 (N_13028,N_11656,N_11408);
or U13029 (N_13029,N_10814,N_11304);
and U13030 (N_13030,N_11204,N_11081);
nor U13031 (N_13031,N_10558,N_11489);
or U13032 (N_13032,N_11391,N_11005);
and U13033 (N_13033,N_11618,N_10881);
and U13034 (N_13034,N_11149,N_10652);
or U13035 (N_13035,N_10582,N_10903);
xnor U13036 (N_13036,N_10831,N_11065);
xnor U13037 (N_13037,N_11359,N_11218);
xor U13038 (N_13038,N_10887,N_11585);
nor U13039 (N_13039,N_10990,N_11305);
xor U13040 (N_13040,N_10912,N_11223);
or U13041 (N_13041,N_10936,N_11872);
and U13042 (N_13042,N_11384,N_10756);
or U13043 (N_13043,N_11907,N_11310);
nor U13044 (N_13044,N_11440,N_10661);
nor U13045 (N_13045,N_11748,N_11363);
nor U13046 (N_13046,N_10931,N_11759);
xnor U13047 (N_13047,N_11983,N_10688);
nand U13048 (N_13048,N_11441,N_10790);
nor U13049 (N_13049,N_11276,N_11938);
nor U13050 (N_13050,N_10589,N_10646);
xor U13051 (N_13051,N_11764,N_10607);
nor U13052 (N_13052,N_10532,N_11410);
and U13053 (N_13053,N_11825,N_11419);
nor U13054 (N_13054,N_10891,N_11596);
or U13055 (N_13055,N_11698,N_11441);
nor U13056 (N_13056,N_10739,N_11013);
nor U13057 (N_13057,N_10819,N_10939);
or U13058 (N_13058,N_10802,N_10961);
xor U13059 (N_13059,N_11956,N_11628);
nor U13060 (N_13060,N_11760,N_11996);
and U13061 (N_13061,N_11997,N_11687);
nand U13062 (N_13062,N_11748,N_11848);
and U13063 (N_13063,N_11815,N_10975);
nand U13064 (N_13064,N_10530,N_11952);
or U13065 (N_13065,N_11673,N_11227);
and U13066 (N_13066,N_11269,N_10984);
nand U13067 (N_13067,N_10687,N_10500);
nor U13068 (N_13068,N_11208,N_10538);
and U13069 (N_13069,N_10995,N_10710);
and U13070 (N_13070,N_11628,N_10716);
and U13071 (N_13071,N_11222,N_10803);
nor U13072 (N_13072,N_11041,N_11704);
or U13073 (N_13073,N_11904,N_11606);
and U13074 (N_13074,N_11416,N_11735);
or U13075 (N_13075,N_11395,N_10578);
and U13076 (N_13076,N_11744,N_11205);
nor U13077 (N_13077,N_11506,N_10599);
or U13078 (N_13078,N_11206,N_11373);
and U13079 (N_13079,N_11140,N_10586);
xnor U13080 (N_13080,N_11158,N_11736);
nor U13081 (N_13081,N_11963,N_10532);
nand U13082 (N_13082,N_11762,N_11777);
nor U13083 (N_13083,N_11144,N_11599);
nand U13084 (N_13084,N_11281,N_11144);
nor U13085 (N_13085,N_10831,N_10564);
and U13086 (N_13086,N_11637,N_10775);
or U13087 (N_13087,N_10851,N_11207);
nand U13088 (N_13088,N_10933,N_11093);
xor U13089 (N_13089,N_10945,N_11663);
or U13090 (N_13090,N_11214,N_11426);
xor U13091 (N_13091,N_11904,N_11537);
or U13092 (N_13092,N_10955,N_11619);
xor U13093 (N_13093,N_11066,N_11925);
xor U13094 (N_13094,N_11878,N_10985);
and U13095 (N_13095,N_11864,N_10829);
or U13096 (N_13096,N_10710,N_11056);
xor U13097 (N_13097,N_10677,N_11353);
nand U13098 (N_13098,N_11806,N_10662);
nand U13099 (N_13099,N_11322,N_11188);
nor U13100 (N_13100,N_11763,N_10551);
or U13101 (N_13101,N_11356,N_11233);
and U13102 (N_13102,N_11369,N_10748);
or U13103 (N_13103,N_11767,N_11120);
nand U13104 (N_13104,N_11768,N_11175);
and U13105 (N_13105,N_11213,N_10522);
or U13106 (N_13106,N_11830,N_11775);
or U13107 (N_13107,N_10853,N_11257);
nand U13108 (N_13108,N_11699,N_11742);
nand U13109 (N_13109,N_11238,N_11617);
or U13110 (N_13110,N_11565,N_11021);
xor U13111 (N_13111,N_10766,N_10941);
nand U13112 (N_13112,N_11470,N_10983);
xnor U13113 (N_13113,N_10673,N_10953);
nand U13114 (N_13114,N_10787,N_11044);
and U13115 (N_13115,N_11477,N_11060);
nor U13116 (N_13116,N_10887,N_10659);
or U13117 (N_13117,N_10595,N_11154);
nor U13118 (N_13118,N_10852,N_10780);
and U13119 (N_13119,N_10968,N_11222);
nand U13120 (N_13120,N_11499,N_11312);
nand U13121 (N_13121,N_11726,N_11899);
or U13122 (N_13122,N_10507,N_11548);
and U13123 (N_13123,N_10716,N_11123);
nand U13124 (N_13124,N_10804,N_11164);
or U13125 (N_13125,N_11765,N_10835);
and U13126 (N_13126,N_10924,N_11877);
or U13127 (N_13127,N_11946,N_10844);
xnor U13128 (N_13128,N_11777,N_11962);
and U13129 (N_13129,N_11924,N_10774);
and U13130 (N_13130,N_11306,N_11877);
nand U13131 (N_13131,N_10699,N_11004);
nand U13132 (N_13132,N_11275,N_11519);
xnor U13133 (N_13133,N_11258,N_11965);
or U13134 (N_13134,N_11951,N_11930);
xor U13135 (N_13135,N_11955,N_10744);
xor U13136 (N_13136,N_11765,N_11994);
xor U13137 (N_13137,N_11886,N_11013);
nand U13138 (N_13138,N_11698,N_11069);
nand U13139 (N_13139,N_11596,N_11704);
or U13140 (N_13140,N_10642,N_11793);
and U13141 (N_13141,N_11260,N_10654);
and U13142 (N_13142,N_10815,N_10698);
nor U13143 (N_13143,N_11169,N_10869);
nand U13144 (N_13144,N_11714,N_11407);
nor U13145 (N_13145,N_11069,N_10660);
or U13146 (N_13146,N_11840,N_11279);
and U13147 (N_13147,N_11813,N_10824);
xor U13148 (N_13148,N_11080,N_11619);
xor U13149 (N_13149,N_11245,N_10977);
xor U13150 (N_13150,N_11580,N_11933);
nor U13151 (N_13151,N_10930,N_10775);
nor U13152 (N_13152,N_11664,N_11408);
nor U13153 (N_13153,N_11932,N_11533);
xor U13154 (N_13154,N_11595,N_11523);
or U13155 (N_13155,N_11855,N_11666);
and U13156 (N_13156,N_10896,N_10846);
nand U13157 (N_13157,N_10657,N_10817);
and U13158 (N_13158,N_11795,N_11499);
and U13159 (N_13159,N_11733,N_11629);
xor U13160 (N_13160,N_11254,N_10580);
nand U13161 (N_13161,N_10686,N_10677);
nand U13162 (N_13162,N_11047,N_11125);
nand U13163 (N_13163,N_11087,N_11532);
nor U13164 (N_13164,N_10980,N_11563);
and U13165 (N_13165,N_11717,N_10873);
nor U13166 (N_13166,N_10506,N_11328);
nand U13167 (N_13167,N_10874,N_11984);
nand U13168 (N_13168,N_10916,N_11672);
or U13169 (N_13169,N_11511,N_11994);
and U13170 (N_13170,N_11230,N_11025);
or U13171 (N_13171,N_11917,N_10718);
and U13172 (N_13172,N_11851,N_11438);
and U13173 (N_13173,N_10896,N_10604);
nor U13174 (N_13174,N_11117,N_11986);
or U13175 (N_13175,N_11939,N_11282);
or U13176 (N_13176,N_10959,N_11789);
nor U13177 (N_13177,N_10539,N_11852);
xnor U13178 (N_13178,N_11974,N_11534);
nand U13179 (N_13179,N_11911,N_11475);
and U13180 (N_13180,N_10879,N_11854);
or U13181 (N_13181,N_11830,N_11988);
nor U13182 (N_13182,N_11386,N_11943);
nor U13183 (N_13183,N_11442,N_11630);
nor U13184 (N_13184,N_11388,N_11479);
nor U13185 (N_13185,N_11369,N_10755);
or U13186 (N_13186,N_11370,N_10542);
nand U13187 (N_13187,N_11233,N_11595);
xor U13188 (N_13188,N_11487,N_11483);
xnor U13189 (N_13189,N_10596,N_11170);
and U13190 (N_13190,N_10521,N_11436);
or U13191 (N_13191,N_10603,N_11656);
nand U13192 (N_13192,N_10919,N_10774);
or U13193 (N_13193,N_10614,N_11358);
nor U13194 (N_13194,N_10857,N_11415);
and U13195 (N_13195,N_10963,N_10718);
nand U13196 (N_13196,N_11923,N_11181);
xor U13197 (N_13197,N_11264,N_10849);
nor U13198 (N_13198,N_11702,N_10777);
nand U13199 (N_13199,N_10595,N_11861);
nand U13200 (N_13200,N_10679,N_11076);
nand U13201 (N_13201,N_11943,N_11967);
or U13202 (N_13202,N_11306,N_10907);
nor U13203 (N_13203,N_11905,N_10918);
or U13204 (N_13204,N_11734,N_11250);
xnor U13205 (N_13205,N_11691,N_10532);
or U13206 (N_13206,N_11076,N_10608);
or U13207 (N_13207,N_11313,N_11135);
xnor U13208 (N_13208,N_10515,N_11653);
and U13209 (N_13209,N_11001,N_11193);
xor U13210 (N_13210,N_11831,N_11445);
or U13211 (N_13211,N_11963,N_10954);
nand U13212 (N_13212,N_11566,N_11585);
nand U13213 (N_13213,N_11681,N_11092);
nor U13214 (N_13214,N_11560,N_10642);
nor U13215 (N_13215,N_11947,N_11566);
nand U13216 (N_13216,N_11657,N_11245);
and U13217 (N_13217,N_11126,N_11898);
and U13218 (N_13218,N_11316,N_11963);
and U13219 (N_13219,N_10943,N_11160);
nand U13220 (N_13220,N_11481,N_11946);
xor U13221 (N_13221,N_11114,N_11566);
or U13222 (N_13222,N_11057,N_11845);
nor U13223 (N_13223,N_11129,N_11794);
xnor U13224 (N_13224,N_11140,N_10691);
nand U13225 (N_13225,N_10805,N_11902);
or U13226 (N_13226,N_10512,N_11292);
or U13227 (N_13227,N_11299,N_11471);
or U13228 (N_13228,N_11792,N_10829);
nand U13229 (N_13229,N_11753,N_10580);
nand U13230 (N_13230,N_10948,N_11522);
xnor U13231 (N_13231,N_10996,N_10503);
xor U13232 (N_13232,N_10845,N_10814);
and U13233 (N_13233,N_10942,N_10988);
xor U13234 (N_13234,N_11751,N_10699);
nor U13235 (N_13235,N_11998,N_10561);
or U13236 (N_13236,N_10753,N_10670);
nor U13237 (N_13237,N_11044,N_11552);
nand U13238 (N_13238,N_11696,N_11948);
or U13239 (N_13239,N_10724,N_11284);
or U13240 (N_13240,N_11870,N_11560);
nand U13241 (N_13241,N_11690,N_10748);
and U13242 (N_13242,N_11289,N_11989);
xor U13243 (N_13243,N_11721,N_11063);
nand U13244 (N_13244,N_11452,N_11334);
nor U13245 (N_13245,N_10866,N_11948);
nand U13246 (N_13246,N_10662,N_11361);
and U13247 (N_13247,N_10676,N_11272);
xnor U13248 (N_13248,N_10863,N_11413);
nand U13249 (N_13249,N_11085,N_10976);
and U13250 (N_13250,N_11970,N_11281);
xnor U13251 (N_13251,N_11855,N_10700);
and U13252 (N_13252,N_10694,N_11558);
xnor U13253 (N_13253,N_10521,N_10713);
nor U13254 (N_13254,N_10616,N_10546);
xor U13255 (N_13255,N_11681,N_11439);
xnor U13256 (N_13256,N_11449,N_11514);
and U13257 (N_13257,N_11439,N_10865);
xor U13258 (N_13258,N_11116,N_11614);
and U13259 (N_13259,N_11723,N_11348);
nand U13260 (N_13260,N_11689,N_11740);
nand U13261 (N_13261,N_10943,N_11438);
or U13262 (N_13262,N_11544,N_11478);
nand U13263 (N_13263,N_10900,N_11134);
nor U13264 (N_13264,N_11240,N_11444);
nor U13265 (N_13265,N_11438,N_11931);
xnor U13266 (N_13266,N_11863,N_11587);
and U13267 (N_13267,N_11523,N_10571);
xor U13268 (N_13268,N_11346,N_11757);
and U13269 (N_13269,N_10991,N_10577);
nor U13270 (N_13270,N_11089,N_10595);
nor U13271 (N_13271,N_10888,N_11661);
nand U13272 (N_13272,N_10830,N_11103);
xnor U13273 (N_13273,N_11493,N_11350);
nand U13274 (N_13274,N_11312,N_10822);
nand U13275 (N_13275,N_11778,N_10713);
or U13276 (N_13276,N_10857,N_10917);
nand U13277 (N_13277,N_11451,N_11148);
nor U13278 (N_13278,N_11172,N_11339);
nor U13279 (N_13279,N_11585,N_11883);
nand U13280 (N_13280,N_11136,N_11156);
xnor U13281 (N_13281,N_11883,N_10865);
xor U13282 (N_13282,N_11056,N_10869);
nor U13283 (N_13283,N_10896,N_11471);
or U13284 (N_13284,N_10770,N_11745);
and U13285 (N_13285,N_11775,N_10799);
and U13286 (N_13286,N_11022,N_10874);
and U13287 (N_13287,N_11733,N_11283);
xor U13288 (N_13288,N_11879,N_11391);
xnor U13289 (N_13289,N_10518,N_10933);
and U13290 (N_13290,N_11958,N_11964);
xnor U13291 (N_13291,N_11164,N_10542);
nand U13292 (N_13292,N_11989,N_11999);
nand U13293 (N_13293,N_11444,N_11265);
nand U13294 (N_13294,N_11393,N_10847);
xnor U13295 (N_13295,N_11620,N_11446);
nand U13296 (N_13296,N_11091,N_11009);
nor U13297 (N_13297,N_11130,N_11033);
and U13298 (N_13298,N_11809,N_10944);
nand U13299 (N_13299,N_11070,N_10836);
and U13300 (N_13300,N_11105,N_11813);
xor U13301 (N_13301,N_11145,N_10913);
and U13302 (N_13302,N_10789,N_11375);
xnor U13303 (N_13303,N_11874,N_11062);
and U13304 (N_13304,N_11594,N_11712);
nor U13305 (N_13305,N_10569,N_11334);
and U13306 (N_13306,N_11558,N_10715);
xnor U13307 (N_13307,N_10719,N_11026);
and U13308 (N_13308,N_10511,N_11141);
nor U13309 (N_13309,N_11629,N_10806);
xor U13310 (N_13310,N_11520,N_11288);
nand U13311 (N_13311,N_11361,N_10712);
nand U13312 (N_13312,N_11872,N_11689);
nand U13313 (N_13313,N_10892,N_11000);
or U13314 (N_13314,N_11268,N_11496);
or U13315 (N_13315,N_10838,N_10609);
nand U13316 (N_13316,N_11669,N_11731);
and U13317 (N_13317,N_10518,N_11661);
xor U13318 (N_13318,N_11350,N_11816);
xor U13319 (N_13319,N_10886,N_11235);
nand U13320 (N_13320,N_10845,N_10650);
nor U13321 (N_13321,N_10692,N_11009);
xor U13322 (N_13322,N_11493,N_11337);
or U13323 (N_13323,N_10916,N_11164);
nand U13324 (N_13324,N_11835,N_11597);
xor U13325 (N_13325,N_11565,N_10881);
and U13326 (N_13326,N_11662,N_10861);
xor U13327 (N_13327,N_10590,N_11316);
nand U13328 (N_13328,N_10532,N_11342);
or U13329 (N_13329,N_11863,N_10538);
nor U13330 (N_13330,N_11557,N_11188);
and U13331 (N_13331,N_11952,N_11791);
xnor U13332 (N_13332,N_10516,N_11955);
nand U13333 (N_13333,N_10948,N_10849);
xor U13334 (N_13334,N_11880,N_11199);
xor U13335 (N_13335,N_10884,N_10684);
or U13336 (N_13336,N_10974,N_11881);
xnor U13337 (N_13337,N_11830,N_11578);
nand U13338 (N_13338,N_11375,N_11929);
nand U13339 (N_13339,N_10536,N_10572);
nand U13340 (N_13340,N_11892,N_11023);
xnor U13341 (N_13341,N_10748,N_10968);
nand U13342 (N_13342,N_11450,N_11064);
or U13343 (N_13343,N_10876,N_10705);
xnor U13344 (N_13344,N_11248,N_11656);
or U13345 (N_13345,N_11838,N_11810);
xnor U13346 (N_13346,N_11113,N_10629);
or U13347 (N_13347,N_10674,N_10771);
nor U13348 (N_13348,N_11286,N_11384);
nand U13349 (N_13349,N_10758,N_11153);
or U13350 (N_13350,N_11707,N_10829);
and U13351 (N_13351,N_11711,N_11956);
nand U13352 (N_13352,N_11004,N_10729);
nand U13353 (N_13353,N_10721,N_11384);
and U13354 (N_13354,N_11070,N_11493);
nand U13355 (N_13355,N_11219,N_11419);
and U13356 (N_13356,N_11460,N_11431);
or U13357 (N_13357,N_11123,N_11865);
xnor U13358 (N_13358,N_10548,N_11115);
and U13359 (N_13359,N_10522,N_10619);
and U13360 (N_13360,N_10767,N_11333);
nand U13361 (N_13361,N_10982,N_10707);
or U13362 (N_13362,N_11268,N_11876);
xnor U13363 (N_13363,N_11004,N_10668);
xor U13364 (N_13364,N_11346,N_11549);
nor U13365 (N_13365,N_10630,N_11527);
nor U13366 (N_13366,N_11759,N_11774);
nor U13367 (N_13367,N_11718,N_11770);
nand U13368 (N_13368,N_11604,N_11337);
nand U13369 (N_13369,N_11408,N_10542);
nand U13370 (N_13370,N_11080,N_11527);
or U13371 (N_13371,N_11060,N_10773);
or U13372 (N_13372,N_11402,N_11796);
nand U13373 (N_13373,N_11682,N_11579);
or U13374 (N_13374,N_11870,N_10727);
and U13375 (N_13375,N_10800,N_10966);
nor U13376 (N_13376,N_11392,N_10770);
or U13377 (N_13377,N_11164,N_11009);
or U13378 (N_13378,N_11315,N_11281);
nor U13379 (N_13379,N_11716,N_10925);
nor U13380 (N_13380,N_11188,N_11176);
or U13381 (N_13381,N_11455,N_11658);
nand U13382 (N_13382,N_11790,N_10846);
or U13383 (N_13383,N_11585,N_11652);
xor U13384 (N_13384,N_10925,N_11606);
xor U13385 (N_13385,N_10665,N_11394);
nor U13386 (N_13386,N_11324,N_11102);
and U13387 (N_13387,N_10863,N_11441);
xor U13388 (N_13388,N_10544,N_11114);
xor U13389 (N_13389,N_11736,N_11545);
nor U13390 (N_13390,N_10862,N_11033);
nor U13391 (N_13391,N_10798,N_10531);
nor U13392 (N_13392,N_11229,N_11087);
and U13393 (N_13393,N_11385,N_11593);
nand U13394 (N_13394,N_11927,N_11909);
and U13395 (N_13395,N_10982,N_11279);
and U13396 (N_13396,N_11301,N_11892);
or U13397 (N_13397,N_11976,N_11810);
nand U13398 (N_13398,N_11468,N_11951);
nand U13399 (N_13399,N_11497,N_11689);
xor U13400 (N_13400,N_10548,N_10788);
nand U13401 (N_13401,N_11661,N_11087);
xor U13402 (N_13402,N_11969,N_10878);
nor U13403 (N_13403,N_11431,N_10529);
and U13404 (N_13404,N_10670,N_11237);
and U13405 (N_13405,N_11710,N_11841);
nor U13406 (N_13406,N_11302,N_11366);
and U13407 (N_13407,N_11812,N_10942);
nor U13408 (N_13408,N_10811,N_11528);
nor U13409 (N_13409,N_11572,N_10516);
xor U13410 (N_13410,N_11334,N_10956);
xor U13411 (N_13411,N_11856,N_10796);
and U13412 (N_13412,N_11733,N_11668);
and U13413 (N_13413,N_10500,N_10679);
nand U13414 (N_13414,N_11284,N_11604);
nand U13415 (N_13415,N_11232,N_11298);
xnor U13416 (N_13416,N_11477,N_10538);
nor U13417 (N_13417,N_10686,N_11594);
and U13418 (N_13418,N_11206,N_11129);
xnor U13419 (N_13419,N_11896,N_11375);
xnor U13420 (N_13420,N_11653,N_11416);
and U13421 (N_13421,N_11443,N_11412);
xor U13422 (N_13422,N_11674,N_10733);
xnor U13423 (N_13423,N_11539,N_10665);
xor U13424 (N_13424,N_11840,N_11610);
or U13425 (N_13425,N_10580,N_11510);
xnor U13426 (N_13426,N_11094,N_11355);
and U13427 (N_13427,N_11708,N_11328);
and U13428 (N_13428,N_11821,N_10705);
xnor U13429 (N_13429,N_10863,N_11327);
nor U13430 (N_13430,N_11270,N_10930);
and U13431 (N_13431,N_11249,N_10984);
nand U13432 (N_13432,N_10755,N_11723);
nor U13433 (N_13433,N_11726,N_10518);
nor U13434 (N_13434,N_11793,N_11737);
or U13435 (N_13435,N_11591,N_10551);
nand U13436 (N_13436,N_11558,N_11573);
nor U13437 (N_13437,N_11084,N_10877);
and U13438 (N_13438,N_10800,N_10997);
nand U13439 (N_13439,N_10595,N_11353);
nand U13440 (N_13440,N_10773,N_11858);
and U13441 (N_13441,N_11736,N_11346);
xor U13442 (N_13442,N_10685,N_11421);
or U13443 (N_13443,N_10748,N_11521);
or U13444 (N_13444,N_11177,N_10666);
xor U13445 (N_13445,N_11629,N_11153);
or U13446 (N_13446,N_10788,N_10865);
xor U13447 (N_13447,N_11698,N_11430);
xor U13448 (N_13448,N_11790,N_11391);
and U13449 (N_13449,N_11651,N_11416);
nor U13450 (N_13450,N_10653,N_11793);
nand U13451 (N_13451,N_11353,N_10600);
or U13452 (N_13452,N_10788,N_11997);
xnor U13453 (N_13453,N_11737,N_11625);
nor U13454 (N_13454,N_11230,N_10554);
and U13455 (N_13455,N_11815,N_11211);
nand U13456 (N_13456,N_11858,N_11388);
or U13457 (N_13457,N_11047,N_11203);
nand U13458 (N_13458,N_11910,N_11149);
and U13459 (N_13459,N_10701,N_11852);
nor U13460 (N_13460,N_11993,N_11758);
or U13461 (N_13461,N_10935,N_10611);
nor U13462 (N_13462,N_11269,N_11586);
xor U13463 (N_13463,N_11515,N_11788);
nor U13464 (N_13464,N_11545,N_11463);
xnor U13465 (N_13465,N_11871,N_11602);
nand U13466 (N_13466,N_11341,N_11688);
or U13467 (N_13467,N_10578,N_11232);
and U13468 (N_13468,N_11829,N_11495);
nand U13469 (N_13469,N_11766,N_11103);
and U13470 (N_13470,N_11177,N_10779);
and U13471 (N_13471,N_11606,N_10756);
xnor U13472 (N_13472,N_11883,N_11017);
or U13473 (N_13473,N_11180,N_11738);
xnor U13474 (N_13474,N_10719,N_11015);
nor U13475 (N_13475,N_10879,N_11114);
xor U13476 (N_13476,N_11674,N_10957);
and U13477 (N_13477,N_11486,N_11860);
and U13478 (N_13478,N_11581,N_10781);
nor U13479 (N_13479,N_11869,N_11625);
xor U13480 (N_13480,N_11322,N_10977);
or U13481 (N_13481,N_10842,N_11327);
nand U13482 (N_13482,N_11474,N_11525);
nand U13483 (N_13483,N_10570,N_11364);
xor U13484 (N_13484,N_11995,N_10765);
and U13485 (N_13485,N_11348,N_10996);
nor U13486 (N_13486,N_10919,N_11608);
xor U13487 (N_13487,N_11440,N_11478);
or U13488 (N_13488,N_11445,N_11345);
nor U13489 (N_13489,N_11743,N_10725);
or U13490 (N_13490,N_10511,N_11183);
xor U13491 (N_13491,N_10999,N_11649);
or U13492 (N_13492,N_11076,N_11201);
nor U13493 (N_13493,N_10728,N_10659);
nand U13494 (N_13494,N_11327,N_11607);
nor U13495 (N_13495,N_11186,N_11395);
nor U13496 (N_13496,N_11032,N_11303);
and U13497 (N_13497,N_10822,N_11550);
and U13498 (N_13498,N_11330,N_11942);
and U13499 (N_13499,N_11785,N_10845);
xor U13500 (N_13500,N_12760,N_12205);
nor U13501 (N_13501,N_13411,N_12624);
or U13502 (N_13502,N_12730,N_13402);
nand U13503 (N_13503,N_12503,N_13368);
nor U13504 (N_13504,N_12831,N_12709);
nand U13505 (N_13505,N_12726,N_12448);
nor U13506 (N_13506,N_13341,N_12969);
xnor U13507 (N_13507,N_13254,N_13346);
nor U13508 (N_13508,N_12770,N_12317);
or U13509 (N_13509,N_12963,N_12718);
nor U13510 (N_13510,N_13059,N_13219);
nand U13511 (N_13511,N_12595,N_12204);
nor U13512 (N_13512,N_12288,N_12540);
nor U13513 (N_13513,N_12435,N_13350);
and U13514 (N_13514,N_12162,N_13279);
nor U13515 (N_13515,N_12738,N_12722);
xnor U13516 (N_13516,N_13386,N_12826);
xnor U13517 (N_13517,N_12386,N_13239);
nand U13518 (N_13518,N_13248,N_13268);
or U13519 (N_13519,N_12615,N_12515);
and U13520 (N_13520,N_12387,N_12130);
and U13521 (N_13521,N_12388,N_13366);
and U13522 (N_13522,N_13029,N_13423);
nand U13523 (N_13523,N_13357,N_13178);
and U13524 (N_13524,N_12869,N_12511);
and U13525 (N_13525,N_12028,N_13300);
nor U13526 (N_13526,N_12566,N_13175);
or U13527 (N_13527,N_12078,N_12497);
nor U13528 (N_13528,N_13427,N_12279);
xor U13529 (N_13529,N_12412,N_13023);
xor U13530 (N_13530,N_12460,N_12899);
nand U13531 (N_13531,N_12865,N_13359);
xor U13532 (N_13532,N_13024,N_13018);
nand U13533 (N_13533,N_12225,N_12104);
xnor U13534 (N_13534,N_13429,N_13140);
or U13535 (N_13535,N_13474,N_13276);
xor U13536 (N_13536,N_12827,N_13403);
and U13537 (N_13537,N_12939,N_13398);
and U13538 (N_13538,N_12820,N_13456);
xor U13539 (N_13539,N_12587,N_12254);
nand U13540 (N_13540,N_12828,N_12608);
and U13541 (N_13541,N_12416,N_12764);
nor U13542 (N_13542,N_13484,N_12466);
or U13543 (N_13543,N_12716,N_13339);
or U13544 (N_13544,N_12598,N_12297);
nor U13545 (N_13545,N_12147,N_12834);
nor U13546 (N_13546,N_13347,N_12055);
nor U13547 (N_13547,N_13183,N_13278);
and U13548 (N_13548,N_12610,N_13288);
nor U13549 (N_13549,N_12380,N_12090);
xnor U13550 (N_13550,N_12282,N_13395);
or U13551 (N_13551,N_12065,N_12061);
or U13552 (N_13552,N_13056,N_12246);
nand U13553 (N_13553,N_12512,N_12656);
nor U13554 (N_13554,N_12620,N_12371);
nor U13555 (N_13555,N_12680,N_12488);
nand U13556 (N_13556,N_12783,N_12189);
and U13557 (N_13557,N_13244,N_12342);
nand U13558 (N_13558,N_13007,N_12493);
xor U13559 (N_13559,N_13103,N_12842);
xnor U13560 (N_13560,N_13010,N_13358);
xor U13561 (N_13561,N_12069,N_13048);
nand U13562 (N_13562,N_13466,N_12663);
xor U13563 (N_13563,N_13038,N_12005);
xor U13564 (N_13564,N_13327,N_13488);
and U13565 (N_13565,N_13040,N_12904);
nand U13566 (N_13566,N_12073,N_12075);
or U13567 (N_13567,N_12588,N_12034);
or U13568 (N_13568,N_13206,N_12607);
nor U13569 (N_13569,N_12965,N_12191);
and U13570 (N_13570,N_13209,N_12487);
or U13571 (N_13571,N_12143,N_12099);
nor U13572 (N_13572,N_12907,N_13397);
nand U13573 (N_13573,N_12547,N_13230);
or U13574 (N_13574,N_12799,N_12704);
nor U13575 (N_13575,N_12968,N_12165);
nand U13576 (N_13576,N_13174,N_13080);
nand U13577 (N_13577,N_13381,N_13044);
and U13578 (N_13578,N_12436,N_13153);
nand U13579 (N_13579,N_12936,N_13246);
and U13580 (N_13580,N_13430,N_12955);
nand U13581 (N_13581,N_12214,N_13160);
nand U13582 (N_13582,N_13476,N_12149);
nor U13583 (N_13583,N_12271,N_13422);
nor U13584 (N_13584,N_12128,N_13020);
or U13585 (N_13585,N_13270,N_12402);
and U13586 (N_13586,N_12697,N_12173);
or U13587 (N_13587,N_13120,N_12888);
xnor U13588 (N_13588,N_12894,N_13022);
and U13589 (N_13589,N_12043,N_12242);
or U13590 (N_13590,N_13417,N_13063);
nor U13591 (N_13591,N_12184,N_12954);
nor U13592 (N_13592,N_12372,N_13033);
xor U13593 (N_13593,N_12791,N_12066);
nand U13594 (N_13594,N_13035,N_13407);
nor U13595 (N_13595,N_12864,N_12074);
or U13596 (N_13596,N_12657,N_12776);
xnor U13597 (N_13597,N_12672,N_13252);
nand U13598 (N_13598,N_13194,N_12685);
or U13599 (N_13599,N_12689,N_13091);
and U13600 (N_13600,N_12578,N_12159);
nand U13601 (N_13601,N_13060,N_12688);
nand U13602 (N_13602,N_12998,N_13337);
nand U13603 (N_13603,N_13169,N_12743);
nor U13604 (N_13604,N_13172,N_12059);
nor U13605 (N_13605,N_12118,N_12352);
nor U13606 (N_13606,N_12422,N_13089);
nor U13607 (N_13607,N_12115,N_13371);
nand U13608 (N_13608,N_12396,N_12261);
and U13609 (N_13609,N_12604,N_12027);
or U13610 (N_13610,N_12433,N_12108);
nand U13611 (N_13611,N_12035,N_12506);
xnor U13612 (N_13612,N_13222,N_13070);
or U13613 (N_13613,N_12878,N_12077);
nand U13614 (N_13614,N_12852,N_12366);
nand U13615 (N_13615,N_12498,N_12980);
and U13616 (N_13616,N_13168,N_12082);
and U13617 (N_13617,N_12221,N_12177);
nor U13618 (N_13618,N_13037,N_12219);
and U13619 (N_13619,N_13264,N_13491);
and U13620 (N_13620,N_13287,N_12345);
and U13621 (N_13621,N_12470,N_12895);
and U13622 (N_13622,N_12986,N_13331);
or U13623 (N_13623,N_13237,N_13375);
nor U13624 (N_13624,N_12974,N_12331);
and U13625 (N_13625,N_12109,N_12772);
xor U13626 (N_13626,N_13134,N_12010);
or U13627 (N_13627,N_13437,N_12196);
nor U13628 (N_13628,N_12464,N_12335);
xor U13629 (N_13629,N_12300,N_12721);
or U13630 (N_13630,N_12792,N_12186);
nand U13631 (N_13631,N_12922,N_13154);
nor U13632 (N_13632,N_12605,N_13139);
and U13633 (N_13633,N_12340,N_13101);
nand U13634 (N_13634,N_13187,N_12307);
nand U13635 (N_13635,N_12921,N_12941);
nand U13636 (N_13636,N_12398,N_12855);
and U13637 (N_13637,N_12731,N_12589);
nor U13638 (N_13638,N_13281,N_12400);
and U13639 (N_13639,N_12253,N_13293);
xor U13640 (N_13640,N_13426,N_12911);
or U13641 (N_13641,N_12138,N_12702);
xnor U13642 (N_13642,N_12033,N_12861);
nand U13643 (N_13643,N_13225,N_12736);
nor U13644 (N_13644,N_12677,N_12741);
nor U13645 (N_13645,N_12517,N_12514);
and U13646 (N_13646,N_13275,N_13431);
and U13647 (N_13647,N_12603,N_13390);
xnor U13648 (N_13648,N_13317,N_13072);
and U13649 (N_13649,N_12083,N_12286);
nor U13650 (N_13650,N_12089,N_12107);
nor U13651 (N_13651,N_12343,N_12364);
or U13652 (N_13652,N_13164,N_12347);
and U13653 (N_13653,N_12612,N_12832);
or U13654 (N_13654,N_12447,N_12454);
or U13655 (N_13655,N_12889,N_13394);
nand U13656 (N_13656,N_13079,N_12209);
and U13657 (N_13657,N_12616,N_13321);
and U13658 (N_13658,N_12215,N_13498);
xnor U13659 (N_13659,N_12560,N_12964);
xor U13660 (N_13660,N_12038,N_12113);
xor U13661 (N_13661,N_13138,N_12009);
or U13662 (N_13662,N_12479,N_13255);
nand U13663 (N_13663,N_13050,N_12505);
nor U13664 (N_13664,N_12759,N_13282);
nand U13665 (N_13665,N_13088,N_12442);
nor U13666 (N_13666,N_12040,N_13235);
and U13667 (N_13667,N_12427,N_12379);
and U13668 (N_13668,N_12644,N_13214);
and U13669 (N_13669,N_12863,N_12139);
nor U13670 (N_13670,N_13298,N_12236);
and U13671 (N_13671,N_12859,N_12407);
nor U13672 (N_13672,N_12749,N_12683);
or U13673 (N_13673,N_12896,N_12893);
xor U13674 (N_13674,N_13418,N_12174);
or U13675 (N_13675,N_12593,N_12885);
xnor U13676 (N_13676,N_13142,N_12182);
nor U13677 (N_13677,N_12080,N_12315);
and U13678 (N_13678,N_12927,N_12081);
nand U13679 (N_13679,N_12449,N_13156);
nand U13680 (N_13680,N_12134,N_12539);
or U13681 (N_13681,N_12240,N_12650);
or U13682 (N_13682,N_13444,N_13081);
and U13683 (N_13683,N_13095,N_13047);
and U13684 (N_13684,N_12789,N_13267);
nand U13685 (N_13685,N_12956,N_12100);
or U13686 (N_13686,N_12959,N_13221);
nor U13687 (N_13687,N_13408,N_12244);
nor U13688 (N_13688,N_13083,N_12361);
or U13689 (N_13689,N_12193,N_12359);
and U13690 (N_13690,N_13285,N_12390);
xnor U13691 (N_13691,N_12092,N_13338);
nand U13692 (N_13692,N_13475,N_12745);
or U13693 (N_13693,N_12735,N_12022);
nor U13694 (N_13694,N_12883,N_12044);
and U13695 (N_13695,N_12687,N_13478);
and U13696 (N_13696,N_12678,N_12846);
nor U13697 (N_13697,N_12706,N_13141);
xnor U13698 (N_13698,N_13041,N_12543);
xnor U13699 (N_13699,N_13376,N_12004);
and U13700 (N_13700,N_13189,N_12144);
nand U13701 (N_13701,N_13470,N_12490);
xor U13702 (N_13702,N_12348,N_13036);
nand U13703 (N_13703,N_13208,N_12001);
nand U13704 (N_13704,N_12131,N_12628);
or U13705 (N_13705,N_12739,N_12141);
xor U13706 (N_13706,N_12525,N_12935);
or U13707 (N_13707,N_12949,N_12905);
nor U13708 (N_13708,N_13343,N_12046);
or U13709 (N_13709,N_13245,N_12919);
or U13710 (N_13710,N_12406,N_13494);
nor U13711 (N_13711,N_13192,N_13211);
nor U13712 (N_13712,N_13111,N_13319);
or U13713 (N_13713,N_12171,N_13008);
or U13714 (N_13714,N_12192,N_12983);
nor U13715 (N_13715,N_13453,N_13305);
nand U13716 (N_13716,N_12692,N_12985);
and U13717 (N_13717,N_13492,N_12877);
and U13718 (N_13718,N_13021,N_13240);
nor U13719 (N_13719,N_13412,N_12041);
and U13720 (N_13720,N_12093,N_12195);
nand U13721 (N_13721,N_12676,N_12950);
xnor U13722 (N_13722,N_12232,N_13065);
xor U13723 (N_13723,N_12328,N_12291);
and U13724 (N_13724,N_13146,N_13441);
and U13725 (N_13725,N_12211,N_12385);
nor U13726 (N_13726,N_13284,N_12946);
nand U13727 (N_13727,N_13457,N_13128);
or U13728 (N_13728,N_12779,N_13017);
nor U13729 (N_13729,N_12336,N_12733);
or U13730 (N_13730,N_12876,N_13039);
nor U13731 (N_13731,N_12853,N_12439);
or U13732 (N_13732,N_12640,N_12701);
and U13733 (N_13733,N_13075,N_12984);
and U13734 (N_13734,N_13271,N_12357);
or U13735 (N_13735,N_13042,N_12966);
or U13736 (N_13736,N_12294,N_12684);
or U13737 (N_13737,N_12953,N_13224);
nor U13738 (N_13738,N_13419,N_12555);
and U13739 (N_13739,N_12837,N_12884);
or U13740 (N_13740,N_13087,N_13265);
and U13741 (N_13741,N_12085,N_12573);
nand U13742 (N_13742,N_13485,N_12520);
and U13743 (N_13743,N_12708,N_12565);
nand U13744 (N_13744,N_12368,N_12169);
xor U13745 (N_13745,N_13262,N_13213);
nand U13746 (N_13746,N_12661,N_12848);
xnor U13747 (N_13747,N_13452,N_13295);
or U13748 (N_13748,N_12961,N_12032);
and U13749 (N_13749,N_13260,N_12463);
nand U13750 (N_13750,N_12017,N_13269);
nor U13751 (N_13751,N_12638,N_13217);
nor U13752 (N_13752,N_12830,N_12582);
or U13753 (N_13753,N_12529,N_13414);
and U13754 (N_13754,N_12474,N_13011);
nand U13755 (N_13755,N_12952,N_12334);
and U13756 (N_13756,N_12409,N_12301);
xnor U13757 (N_13757,N_13000,N_13405);
xnor U13758 (N_13758,N_13393,N_12179);
nand U13759 (N_13759,N_13132,N_12947);
nor U13760 (N_13760,N_12707,N_12531);
xnor U13761 (N_13761,N_13205,N_13105);
xnor U13762 (N_13762,N_13186,N_12989);
nand U13763 (N_13763,N_13344,N_12472);
nor U13764 (N_13764,N_12821,N_13228);
and U13765 (N_13765,N_12519,N_12110);
or U13766 (N_13766,N_13181,N_12781);
nor U13767 (N_13767,N_13071,N_13349);
or U13768 (N_13768,N_12462,N_13152);
nor U13769 (N_13769,N_12012,N_12931);
xnor U13770 (N_13770,N_13045,N_13477);
and U13771 (N_13771,N_13185,N_12908);
nand U13772 (N_13772,N_12356,N_13448);
nor U13773 (N_13773,N_12123,N_12223);
nand U13774 (N_13774,N_12750,N_12914);
xor U13775 (N_13775,N_12339,N_12670);
nor U13776 (N_13776,N_12153,N_12910);
and U13777 (N_13777,N_13336,N_12801);
or U13778 (N_13778,N_12190,N_13299);
and U13779 (N_13779,N_13197,N_12793);
xor U13780 (N_13780,N_13435,N_12805);
nand U13781 (N_13781,N_12039,N_12874);
or U13782 (N_13782,N_12287,N_12623);
and U13783 (N_13783,N_12924,N_12932);
xnor U13784 (N_13784,N_12618,N_12972);
nor U13785 (N_13785,N_13487,N_12606);
or U13786 (N_13786,N_12602,N_12483);
nor U13787 (N_13787,N_13472,N_12554);
nand U13788 (N_13788,N_12424,N_13073);
nor U13789 (N_13789,N_12967,N_12370);
nand U13790 (N_13790,N_13297,N_12091);
nor U13791 (N_13791,N_12243,N_13133);
or U13792 (N_13792,N_12290,N_12634);
and U13793 (N_13793,N_12392,N_12729);
nand U13794 (N_13794,N_12748,N_12930);
nand U13795 (N_13795,N_12137,N_13200);
nand U13796 (N_13796,N_13306,N_13450);
nor U13797 (N_13797,N_12381,N_12228);
nand U13798 (N_13798,N_12203,N_12633);
xnor U13799 (N_13799,N_12358,N_12806);
or U13800 (N_13800,N_12129,N_12576);
and U13801 (N_13801,N_12570,N_13084);
or U13802 (N_13802,N_12744,N_13410);
nor U13803 (N_13803,N_12898,N_12194);
nand U13804 (N_13804,N_12673,N_13232);
nor U13805 (N_13805,N_12599,N_12403);
or U13806 (N_13806,N_13380,N_12662);
or U13807 (N_13807,N_12751,N_12161);
and U13808 (N_13808,N_13135,N_13436);
and U13809 (N_13809,N_12596,N_13363);
or U13810 (N_13810,N_12087,N_12377);
nand U13811 (N_13811,N_13369,N_12306);
and U13812 (N_13812,N_13361,N_13165);
nor U13813 (N_13813,N_13451,N_12882);
nor U13814 (N_13814,N_13340,N_12262);
xnor U13815 (N_13815,N_13307,N_12648);
xnor U13816 (N_13816,N_12333,N_12245);
nand U13817 (N_13817,N_12715,N_13283);
nor U13818 (N_13818,N_12063,N_12785);
nor U13819 (N_13819,N_12250,N_12296);
and U13820 (N_13820,N_13166,N_12816);
or U13821 (N_13821,N_12553,N_12230);
and U13822 (N_13822,N_12248,N_12795);
and U13823 (N_13823,N_12272,N_13462);
xnor U13824 (N_13824,N_12023,N_13207);
nor U13825 (N_13825,N_12982,N_13233);
xnor U13826 (N_13826,N_13467,N_12574);
xnor U13827 (N_13827,N_12796,N_13420);
nor U13828 (N_13828,N_12641,N_13392);
xor U13829 (N_13829,N_12235,N_12923);
nor U13830 (N_13830,N_12142,N_12917);
and U13831 (N_13831,N_12548,N_12480);
xnor U13832 (N_13832,N_12774,N_12766);
or U13833 (N_13833,N_12754,N_13465);
xnor U13834 (N_13834,N_12095,N_12283);
nand U13835 (N_13835,N_13389,N_12056);
and U13836 (N_13836,N_12705,N_13318);
nand U13837 (N_13837,N_13031,N_12494);
and U13838 (N_13838,N_12330,N_12824);
and U13839 (N_13839,N_12536,N_12912);
nor U13840 (N_13840,N_12829,N_12501);
nor U13841 (N_13841,N_12742,N_12549);
nor U13842 (N_13842,N_12929,N_12740);
nand U13843 (N_13843,N_12376,N_12870);
nand U13844 (N_13844,N_12018,N_12029);
nor U13845 (N_13845,N_12489,N_13241);
xor U13846 (N_13846,N_13379,N_12468);
or U13847 (N_13847,N_12613,N_12621);
or U13848 (N_13848,N_12410,N_13226);
nor U13849 (N_13849,N_13328,N_12451);
or U13850 (N_13850,N_12126,N_13312);
or U13851 (N_13851,N_12281,N_12054);
xor U13852 (N_13852,N_12755,N_12378);
nand U13853 (N_13853,N_12327,N_13438);
and U13854 (N_13854,N_12668,N_12355);
or U13855 (N_13855,N_12404,N_12305);
or U13856 (N_13856,N_12627,N_12446);
or U13857 (N_13857,N_13385,N_13176);
or U13858 (N_13858,N_12280,N_12133);
xor U13859 (N_13859,N_12132,N_12158);
nor U13860 (N_13860,N_12713,N_12076);
and U13861 (N_13861,N_13067,N_12854);
and U13862 (N_13862,N_12807,N_12943);
and U13863 (N_13863,N_12401,N_12309);
nor U13864 (N_13864,N_12103,N_12524);
nor U13865 (N_13865,N_12784,N_12900);
xnor U13866 (N_13866,N_13433,N_12875);
nor U13867 (N_13867,N_12362,N_13116);
nor U13868 (N_13868,N_13496,N_12586);
nand U13869 (N_13869,N_12491,N_12654);
or U13870 (N_13870,N_12421,N_13188);
or U13871 (N_13871,N_12259,N_12324);
or U13872 (N_13872,N_12866,N_13325);
or U13873 (N_13873,N_13352,N_13333);
or U13874 (N_13874,N_12238,N_12399);
or U13875 (N_13875,N_13499,N_13308);
nand U13876 (N_13876,N_12310,N_12960);
nand U13877 (N_13877,N_12045,N_13370);
nand U13878 (N_13878,N_13387,N_12275);
xor U13879 (N_13879,N_12011,N_13447);
xor U13880 (N_13880,N_12024,N_12535);
nand U13881 (N_13881,N_12594,N_12559);
nor U13882 (N_13882,N_12106,N_13231);
nor U13883 (N_13883,N_13016,N_12550);
or U13884 (N_13884,N_12881,N_12526);
nor U13885 (N_13885,N_12326,N_13061);
nor U13886 (N_13886,N_12415,N_13330);
or U13887 (N_13887,N_12609,N_12234);
nor U13888 (N_13888,N_12732,N_12318);
or U13889 (N_13889,N_12945,N_12533);
nand U13890 (N_13890,N_12665,N_13212);
xor U13891 (N_13891,N_13471,N_12452);
nor U13892 (N_13892,N_12504,N_12206);
or U13893 (N_13893,N_13074,N_12933);
or U13894 (N_13894,N_13147,N_13449);
and U13895 (N_13895,N_12030,N_12860);
or U13896 (N_13896,N_13202,N_12227);
nand U13897 (N_13897,N_13258,N_12769);
or U13898 (N_13898,N_12712,N_12181);
nor U13899 (N_13899,N_13184,N_12050);
nand U13900 (N_13900,N_12457,N_13002);
xnor U13901 (N_13901,N_12902,N_13401);
nand U13902 (N_13902,N_12581,N_13104);
nand U13903 (N_13903,N_12019,N_12441);
and U13904 (N_13904,N_12437,N_12728);
xor U13905 (N_13905,N_12674,N_13198);
or U13906 (N_13906,N_13109,N_12629);
and U13907 (N_13907,N_13455,N_12431);
and U13908 (N_13908,N_13013,N_13043);
nand U13909 (N_13909,N_13329,N_13323);
or U13910 (N_13910,N_12916,N_13082);
and U13911 (N_13911,N_13253,N_13218);
or U13912 (N_13912,N_12176,N_12101);
nor U13913 (N_13913,N_12995,N_13163);
nor U13914 (N_13914,N_12970,N_13309);
and U13915 (N_13915,N_12341,N_12295);
xnor U13916 (N_13916,N_13173,N_12762);
xnor U13917 (N_13917,N_12237,N_12768);
and U13918 (N_13918,N_12218,N_12389);
xnor U13919 (N_13919,N_12053,N_12714);
and U13920 (N_13920,N_12818,N_12405);
nor U13921 (N_13921,N_12383,N_13144);
and U13922 (N_13922,N_12450,N_12417);
xnor U13923 (N_13923,N_13360,N_13054);
nor U13924 (N_13924,N_12973,N_12298);
nor U13925 (N_13925,N_12188,N_13052);
nand U13926 (N_13926,N_13442,N_12630);
nand U13927 (N_13927,N_12591,N_12098);
or U13928 (N_13928,N_13250,N_12485);
xor U13929 (N_13929,N_12850,N_13122);
nor U13930 (N_13930,N_13236,N_13301);
nand U13931 (N_13931,N_13388,N_13196);
and U13932 (N_13932,N_12200,N_13434);
or U13933 (N_13933,N_12256,N_12021);
or U13934 (N_13934,N_12042,N_13157);
nand U13935 (N_13935,N_13148,N_13171);
nand U13936 (N_13936,N_13257,N_13201);
xor U13937 (N_13937,N_12500,N_13396);
xnor U13938 (N_13938,N_12997,N_12516);
nand U13939 (N_13939,N_12199,N_12551);
xnor U13940 (N_13940,N_12096,N_12432);
nand U13941 (N_13941,N_12469,N_13483);
nand U13942 (N_13942,N_13162,N_13334);
and U13943 (N_13943,N_12977,N_12167);
nor U13944 (N_13944,N_12338,N_12163);
and U13945 (N_13945,N_12459,N_12523);
xnor U13946 (N_13946,N_12567,N_12014);
nor U13947 (N_13947,N_12428,N_13425);
and U13948 (N_13948,N_12871,N_13473);
or U13949 (N_13949,N_12815,N_12572);
or U13950 (N_13950,N_12145,N_12892);
and U13951 (N_13951,N_13351,N_13119);
and U13952 (N_13952,N_12787,N_12325);
and U13953 (N_13953,N_12845,N_12094);
and U13954 (N_13954,N_13234,N_12148);
xor U13955 (N_13955,N_13353,N_12268);
nand U13956 (N_13956,N_13445,N_13497);
xor U13957 (N_13957,N_12047,N_12700);
and U13958 (N_13958,N_12639,N_12651);
or U13959 (N_13959,N_13102,N_12015);
nand U13960 (N_13960,N_13458,N_13372);
nor U13961 (N_13961,N_13409,N_12026);
and U13962 (N_13962,N_12086,N_12937);
nor U13963 (N_13963,N_13332,N_12664);
and U13964 (N_13964,N_12391,N_12563);
xor U13965 (N_13965,N_13159,N_12311);
and U13966 (N_13966,N_12157,N_12693);
xor U13967 (N_13967,N_12564,N_12187);
nor U13968 (N_13968,N_12767,N_13129);
and U13969 (N_13969,N_12292,N_12856);
nor U13970 (N_13970,N_12495,N_12150);
nor U13971 (N_13971,N_12263,N_13019);
xnor U13972 (N_13972,N_12322,N_12507);
or U13973 (N_13973,N_12119,N_13100);
xor U13974 (N_13974,N_12626,N_13415);
nor U13975 (N_13975,N_13005,N_12579);
xor U13976 (N_13976,N_12114,N_12284);
nand U13977 (N_13977,N_12957,N_12467);
or U13978 (N_13978,N_12696,N_12841);
nor U13979 (N_13979,N_13014,N_12675);
xnor U13980 (N_13980,N_12267,N_13106);
xor U13981 (N_13981,N_12168,N_12753);
nor U13982 (N_13982,N_13123,N_12915);
and U13983 (N_13983,N_12988,N_12719);
and U13984 (N_13984,N_12140,N_12455);
nor U13985 (N_13985,N_13364,N_12658);
nand U13986 (N_13986,N_12690,N_12723);
and U13987 (N_13987,N_13290,N_12562);
nor U13988 (N_13988,N_12231,N_12360);
or U13989 (N_13989,N_13404,N_12940);
xor U13990 (N_13990,N_12851,N_13155);
xnor U13991 (N_13991,N_13460,N_12052);
xnor U13992 (N_13992,N_12681,N_13243);
nor U13993 (N_13993,N_12475,N_13463);
nand U13994 (N_13994,N_12659,N_12901);
or U13995 (N_13995,N_12071,N_12951);
nor U13996 (N_13996,N_12546,N_13092);
nand U13997 (N_13997,N_12036,N_12411);
nor U13998 (N_13998,N_13459,N_12773);
and U13999 (N_13999,N_12691,N_12369);
or U14000 (N_14000,N_12367,N_12172);
and U14001 (N_14001,N_13032,N_12590);
nand U14002 (N_14002,N_13377,N_12344);
nand U14003 (N_14003,N_12484,N_12111);
nor U14004 (N_14004,N_12285,N_13313);
and U14005 (N_14005,N_12146,N_13158);
xnor U14006 (N_14006,N_13432,N_12302);
or U14007 (N_14007,N_13464,N_12185);
or U14008 (N_14008,N_12720,N_12365);
or U14009 (N_14009,N_12763,N_12064);
nor U14010 (N_14010,N_12224,N_12928);
nand U14011 (N_14011,N_12575,N_12048);
nand U14012 (N_14012,N_12804,N_13294);
nand U14013 (N_14013,N_12482,N_12652);
nor U14014 (N_14014,N_12070,N_12313);
nand U14015 (N_14015,N_12461,N_13322);
nor U14016 (N_14016,N_12008,N_13454);
nand U14017 (N_14017,N_12320,N_12926);
and U14018 (N_14018,N_13439,N_13383);
nor U14019 (N_14019,N_12207,N_12079);
or U14020 (N_14020,N_12007,N_12703);
and U14021 (N_14021,N_13362,N_12393);
or U14022 (N_14022,N_12948,N_12667);
and U14023 (N_14023,N_13373,N_12031);
xnor U14024 (N_14024,N_12269,N_13127);
or U14025 (N_14025,N_12920,N_13136);
or U14026 (N_14026,N_12552,N_13131);
nor U14027 (N_14027,N_13280,N_13034);
or U14028 (N_14028,N_12260,N_12857);
or U14029 (N_14029,N_13068,N_13469);
and U14030 (N_14030,N_12425,N_12999);
nand U14031 (N_14031,N_12020,N_12180);
and U14032 (N_14032,N_12849,N_13266);
nor U14033 (N_14033,N_12813,N_13272);
nor U14034 (N_14034,N_12558,N_12771);
and U14035 (N_14035,N_13025,N_12303);
xor U14036 (N_14036,N_12121,N_12068);
or U14037 (N_14037,N_13161,N_12758);
and U14038 (N_14038,N_13051,N_12440);
and U14039 (N_14039,N_12653,N_12521);
xor U14040 (N_14040,N_12154,N_13170);
nand U14041 (N_14041,N_13015,N_12135);
and U14042 (N_14042,N_12276,N_13367);
xor U14043 (N_14043,N_12887,N_12847);
xnor U14044 (N_14044,N_12597,N_12698);
nor U14045 (N_14045,N_13193,N_12477);
xnor U14046 (N_14046,N_12934,N_13112);
xnor U14047 (N_14047,N_12112,N_13382);
nand U14048 (N_14048,N_12938,N_13115);
nand U14049 (N_14049,N_12125,N_12277);
nand U14050 (N_14050,N_13216,N_12643);
nand U14051 (N_14051,N_13251,N_12136);
or U14052 (N_14052,N_12962,N_12226);
nor U14053 (N_14053,N_13261,N_13291);
nand U14054 (N_14054,N_12522,N_12016);
xor U14055 (N_14055,N_13098,N_12002);
xor U14056 (N_14056,N_13110,N_13107);
nand U14057 (N_14057,N_13097,N_13446);
nand U14058 (N_14058,N_13391,N_12925);
nand U14059 (N_14059,N_12600,N_12170);
or U14060 (N_14060,N_13296,N_12867);
nor U14061 (N_14061,N_12051,N_13259);
nand U14062 (N_14062,N_12419,N_13324);
nand U14063 (N_14063,N_12067,N_12122);
nand U14064 (N_14064,N_13481,N_13495);
nand U14065 (N_14065,N_13263,N_13093);
nor U14066 (N_14066,N_12373,N_12201);
xor U14067 (N_14067,N_13238,N_12217);
nor U14068 (N_14068,N_13489,N_13304);
and U14069 (N_14069,N_13416,N_12264);
xnor U14070 (N_14070,N_13113,N_13480);
nand U14071 (N_14071,N_12886,N_12838);
or U14072 (N_14072,N_12890,N_12571);
and U14073 (N_14073,N_13374,N_12534);
or U14074 (N_14074,N_12987,N_13076);
and U14075 (N_14075,N_12508,N_12976);
xnor U14076 (N_14076,N_12155,N_13326);
or U14077 (N_14077,N_13108,N_12151);
nor U14078 (N_14078,N_13195,N_12375);
and U14079 (N_14079,N_13302,N_12353);
nor U14080 (N_14080,N_13126,N_12646);
nand U14081 (N_14081,N_12164,N_13145);
and U14082 (N_14082,N_12790,N_12891);
nand U14083 (N_14083,N_12354,N_12636);
xor U14084 (N_14084,N_12944,N_12794);
xor U14085 (N_14085,N_12408,N_12839);
nor U14086 (N_14086,N_12323,N_12777);
nand U14087 (N_14087,N_12918,N_13096);
xnor U14088 (N_14088,N_12782,N_12270);
and U14089 (N_14089,N_12737,N_13348);
or U14090 (N_14090,N_12308,N_12210);
nand U14091 (N_14091,N_12823,N_12802);
and U14092 (N_14092,N_13149,N_12476);
nor U14093 (N_14093,N_13055,N_12808);
nand U14094 (N_14094,N_12601,N_13057);
xnor U14095 (N_14095,N_12778,N_13118);
and U14096 (N_14096,N_13345,N_12241);
and U14097 (N_14097,N_12166,N_12510);
or U14098 (N_14098,N_12637,N_12363);
nor U14099 (N_14099,N_12216,N_12251);
xnor U14100 (N_14100,N_12993,N_12699);
or U14101 (N_14101,N_12513,N_12213);
and U14102 (N_14102,N_12429,N_12958);
or U14103 (N_14103,N_12097,N_12329);
xor U14104 (N_14104,N_12502,N_12811);
or U14105 (N_14105,N_12252,N_12622);
nand U14106 (N_14106,N_12102,N_12557);
or U14107 (N_14107,N_13315,N_12532);
nor U14108 (N_14108,N_12258,N_12062);
and U14109 (N_14109,N_12304,N_12592);
nand U14110 (N_14110,N_12418,N_13004);
and U14111 (N_14111,N_12072,N_12669);
nor U14112 (N_14112,N_12212,N_12350);
and U14113 (N_14113,N_12752,N_12542);
or U14114 (N_14114,N_12541,N_13479);
nand U14115 (N_14115,N_13062,N_13210);
and U14116 (N_14116,N_12647,N_12809);
or U14117 (N_14117,N_12175,N_12160);
and U14118 (N_14118,N_12822,N_12814);
and U14119 (N_14119,N_12798,N_12835);
and U14120 (N_14120,N_12906,N_12868);
nor U14121 (N_14121,N_13085,N_12812);
nand U14122 (N_14122,N_13406,N_12438);
or U14123 (N_14123,N_13167,N_12413);
xor U14124 (N_14124,N_12006,N_13356);
or U14125 (N_14125,N_13204,N_12397);
nand U14126 (N_14126,N_12293,N_13256);
or U14127 (N_14127,N_12486,N_13009);
or U14128 (N_14128,N_12711,N_12420);
or U14129 (N_14129,N_12443,N_12465);
nor U14130 (N_14130,N_12202,N_13199);
nor U14131 (N_14131,N_12013,N_13354);
nand U14132 (N_14132,N_12645,N_13180);
or U14133 (N_14133,N_12314,N_12000);
or U14134 (N_14134,N_13421,N_12273);
or U14135 (N_14135,N_13229,N_13335);
xnor U14136 (N_14136,N_12660,N_12084);
nand U14137 (N_14137,N_12836,N_12992);
nor U14138 (N_14138,N_12088,N_12183);
nand U14139 (N_14139,N_12775,N_12426);
and U14140 (N_14140,N_12319,N_13220);
and U14141 (N_14141,N_12649,N_12058);
or U14142 (N_14142,N_12897,N_12278);
or U14143 (N_14143,N_13099,N_12686);
nor U14144 (N_14144,N_12456,N_12580);
nand U14145 (N_14145,N_12445,N_13150);
nor U14146 (N_14146,N_13030,N_12632);
or U14147 (N_14147,N_12528,N_12233);
and U14148 (N_14148,N_12127,N_12312);
nand U14149 (N_14149,N_12178,N_13001);
and U14150 (N_14150,N_12321,N_12274);
or U14151 (N_14151,N_13384,N_13177);
nand U14152 (N_14152,N_12478,N_12727);
and U14153 (N_14153,N_12229,N_12642);
and U14154 (N_14154,N_12655,N_12872);
and U14155 (N_14155,N_12746,N_13400);
nor U14156 (N_14156,N_12481,N_12569);
and U14157 (N_14157,N_12351,N_12530);
nand U14158 (N_14158,N_13143,N_13342);
nand U14159 (N_14159,N_13086,N_12903);
and U14160 (N_14160,N_12817,N_13190);
and U14161 (N_14161,N_12583,N_13316);
or U14162 (N_14162,N_12971,N_12120);
or U14163 (N_14163,N_12538,N_12844);
or U14164 (N_14164,N_12797,N_13028);
and U14165 (N_14165,N_12509,N_12197);
xnor U14166 (N_14166,N_12037,N_12198);
and U14167 (N_14167,N_13292,N_12975);
and U14168 (N_14168,N_13310,N_12124);
or U14169 (N_14169,N_12780,N_12765);
xnor U14170 (N_14170,N_12568,N_12879);
nor U14171 (N_14171,N_13311,N_13286);
or U14172 (N_14172,N_12880,N_12394);
or U14173 (N_14173,N_13130,N_12496);
xnor U14174 (N_14174,N_12862,N_12803);
nor U14175 (N_14175,N_12222,N_13215);
or U14176 (N_14176,N_12332,N_12544);
xor U14177 (N_14177,N_12349,N_13053);
nand U14178 (N_14178,N_12220,N_13179);
and U14179 (N_14179,N_12561,N_12247);
nor U14180 (N_14180,N_12152,N_12116);
and U14181 (N_14181,N_12825,N_13242);
or U14182 (N_14182,N_12810,N_12025);
nor U14183 (N_14183,N_12991,N_12208);
or U14184 (N_14184,N_12611,N_12105);
nor U14185 (N_14185,N_13058,N_13468);
nor U14186 (N_14186,N_13273,N_12717);
or U14187 (N_14187,N_13223,N_13090);
xor U14188 (N_14188,N_12695,N_12492);
and U14189 (N_14189,N_12979,N_12584);
nor U14190 (N_14190,N_12725,N_12156);
and U14191 (N_14191,N_12060,N_13274);
xor U14192 (N_14192,N_12942,N_12978);
and U14193 (N_14193,N_12913,N_12556);
nor U14194 (N_14194,N_12635,N_13424);
nand U14195 (N_14195,N_13027,N_12873);
nor U14196 (N_14196,N_12003,N_13378);
nand U14197 (N_14197,N_12694,N_12266);
nand U14198 (N_14198,N_12994,N_13443);
and U14199 (N_14199,N_12724,N_12843);
nor U14200 (N_14200,N_12049,N_13413);
and U14201 (N_14201,N_12577,N_12840);
xor U14202 (N_14202,N_12981,N_13003);
or U14203 (N_14203,N_13117,N_13365);
and U14204 (N_14204,N_13151,N_12316);
or U14205 (N_14205,N_12710,N_13066);
nand U14206 (N_14206,N_13399,N_12414);
and U14207 (N_14207,N_12117,N_13303);
or U14208 (N_14208,N_12909,N_13124);
nand U14209 (N_14209,N_12458,N_12337);
nor U14210 (N_14210,N_12518,N_13182);
nor U14211 (N_14211,N_12788,N_12614);
nand U14212 (N_14212,N_13440,N_12346);
and U14213 (N_14213,N_13078,N_13490);
nand U14214 (N_14214,N_13428,N_12996);
nand U14215 (N_14215,N_13125,N_13137);
or U14216 (N_14216,N_12625,N_12265);
nor U14217 (N_14217,N_12257,N_13277);
nand U14218 (N_14218,N_12800,N_12734);
nand U14219 (N_14219,N_12671,N_12453);
or U14220 (N_14220,N_13247,N_13461);
xnor U14221 (N_14221,N_13493,N_13012);
and U14222 (N_14222,N_12395,N_12679);
nor U14223 (N_14223,N_12057,N_12757);
and U14224 (N_14224,N_12858,N_13094);
xnor U14225 (N_14225,N_13482,N_13249);
xnor U14226 (N_14226,N_12255,N_12374);
nor U14227 (N_14227,N_12239,N_13077);
and U14228 (N_14228,N_12786,N_13355);
nor U14229 (N_14229,N_12631,N_13314);
xnor U14230 (N_14230,N_12761,N_13026);
nand U14231 (N_14231,N_13114,N_12585);
nor U14232 (N_14232,N_12444,N_13320);
or U14233 (N_14233,N_12499,N_13191);
nand U14234 (N_14234,N_12666,N_13006);
or U14235 (N_14235,N_12473,N_13203);
xor U14236 (N_14236,N_13049,N_12682);
or U14237 (N_14237,N_12384,N_12756);
or U14238 (N_14238,N_13289,N_12833);
nor U14239 (N_14239,N_12289,N_12471);
nand U14240 (N_14240,N_12537,N_12430);
or U14241 (N_14241,N_13121,N_12423);
xor U14242 (N_14242,N_12545,N_12619);
nor U14243 (N_14243,N_13227,N_13046);
and U14244 (N_14244,N_13069,N_12819);
nand U14245 (N_14245,N_13486,N_12990);
xnor U14246 (N_14246,N_12299,N_12617);
xnor U14247 (N_14247,N_12382,N_12747);
nor U14248 (N_14248,N_12249,N_13064);
and U14249 (N_14249,N_12527,N_12434);
or U14250 (N_14250,N_13192,N_13456);
nand U14251 (N_14251,N_12651,N_12205);
nor U14252 (N_14252,N_12677,N_12670);
nand U14253 (N_14253,N_12222,N_12379);
xor U14254 (N_14254,N_13003,N_12411);
and U14255 (N_14255,N_13381,N_13427);
or U14256 (N_14256,N_13486,N_12871);
or U14257 (N_14257,N_13402,N_13341);
nor U14258 (N_14258,N_13476,N_13475);
or U14259 (N_14259,N_13105,N_12951);
nand U14260 (N_14260,N_13398,N_12742);
or U14261 (N_14261,N_12877,N_12132);
nand U14262 (N_14262,N_13239,N_13392);
xnor U14263 (N_14263,N_13235,N_12976);
or U14264 (N_14264,N_12061,N_12650);
nand U14265 (N_14265,N_13483,N_12701);
xor U14266 (N_14266,N_12654,N_12813);
or U14267 (N_14267,N_12984,N_12947);
nand U14268 (N_14268,N_12603,N_13294);
xnor U14269 (N_14269,N_13375,N_12542);
and U14270 (N_14270,N_12284,N_13246);
xnor U14271 (N_14271,N_13070,N_13254);
and U14272 (N_14272,N_12404,N_13153);
or U14273 (N_14273,N_12959,N_12244);
nand U14274 (N_14274,N_12730,N_12397);
and U14275 (N_14275,N_12922,N_12809);
or U14276 (N_14276,N_13076,N_12059);
and U14277 (N_14277,N_13084,N_12747);
and U14278 (N_14278,N_12247,N_12921);
nand U14279 (N_14279,N_12114,N_13147);
or U14280 (N_14280,N_12917,N_12921);
nand U14281 (N_14281,N_12096,N_12637);
xnor U14282 (N_14282,N_12484,N_13205);
xnor U14283 (N_14283,N_13015,N_13068);
and U14284 (N_14284,N_12438,N_13234);
xor U14285 (N_14285,N_12816,N_12707);
or U14286 (N_14286,N_13232,N_12016);
or U14287 (N_14287,N_12466,N_12428);
or U14288 (N_14288,N_13353,N_13401);
or U14289 (N_14289,N_12305,N_12775);
nand U14290 (N_14290,N_12145,N_13239);
nand U14291 (N_14291,N_12881,N_12035);
nor U14292 (N_14292,N_12650,N_12097);
xnor U14293 (N_14293,N_12031,N_12199);
and U14294 (N_14294,N_12518,N_13083);
nor U14295 (N_14295,N_12272,N_13336);
or U14296 (N_14296,N_12593,N_13292);
xnor U14297 (N_14297,N_13135,N_13169);
and U14298 (N_14298,N_13420,N_12465);
nand U14299 (N_14299,N_13030,N_12690);
nand U14300 (N_14300,N_13383,N_12841);
or U14301 (N_14301,N_12257,N_12276);
xor U14302 (N_14302,N_13158,N_13163);
nor U14303 (N_14303,N_13057,N_12114);
and U14304 (N_14304,N_12248,N_13282);
xnor U14305 (N_14305,N_13338,N_13368);
and U14306 (N_14306,N_13007,N_13256);
xor U14307 (N_14307,N_12139,N_13375);
and U14308 (N_14308,N_13081,N_12355);
or U14309 (N_14309,N_12255,N_13386);
xor U14310 (N_14310,N_12298,N_12203);
and U14311 (N_14311,N_13192,N_12497);
xor U14312 (N_14312,N_12320,N_12889);
or U14313 (N_14313,N_12310,N_12707);
xor U14314 (N_14314,N_13213,N_12206);
xor U14315 (N_14315,N_12151,N_13462);
or U14316 (N_14316,N_13236,N_12109);
nand U14317 (N_14317,N_12295,N_13249);
nand U14318 (N_14318,N_12911,N_12550);
nor U14319 (N_14319,N_12058,N_12633);
nor U14320 (N_14320,N_12759,N_13135);
xor U14321 (N_14321,N_12406,N_12567);
and U14322 (N_14322,N_12896,N_13386);
or U14323 (N_14323,N_12921,N_12581);
and U14324 (N_14324,N_12052,N_13342);
nand U14325 (N_14325,N_13180,N_12787);
xnor U14326 (N_14326,N_13149,N_12367);
nand U14327 (N_14327,N_12423,N_12154);
nand U14328 (N_14328,N_12208,N_12921);
and U14329 (N_14329,N_12021,N_12389);
nor U14330 (N_14330,N_13069,N_12163);
and U14331 (N_14331,N_12704,N_13058);
or U14332 (N_14332,N_12041,N_12326);
xnor U14333 (N_14333,N_13065,N_12473);
nor U14334 (N_14334,N_12187,N_12202);
or U14335 (N_14335,N_13243,N_13255);
xnor U14336 (N_14336,N_13492,N_13028);
and U14337 (N_14337,N_13342,N_13252);
xnor U14338 (N_14338,N_12204,N_13408);
or U14339 (N_14339,N_13450,N_13373);
and U14340 (N_14340,N_13382,N_12007);
xor U14341 (N_14341,N_13064,N_12559);
and U14342 (N_14342,N_13055,N_12587);
xnor U14343 (N_14343,N_12402,N_13079);
and U14344 (N_14344,N_12920,N_13207);
xnor U14345 (N_14345,N_12504,N_13388);
xnor U14346 (N_14346,N_13302,N_13047);
or U14347 (N_14347,N_12541,N_12040);
nand U14348 (N_14348,N_12573,N_13475);
xor U14349 (N_14349,N_12834,N_12150);
or U14350 (N_14350,N_12145,N_13010);
nor U14351 (N_14351,N_12346,N_12988);
nor U14352 (N_14352,N_12956,N_13446);
and U14353 (N_14353,N_12319,N_12583);
xor U14354 (N_14354,N_12534,N_13372);
or U14355 (N_14355,N_12373,N_13101);
or U14356 (N_14356,N_13293,N_12668);
xnor U14357 (N_14357,N_13052,N_13110);
or U14358 (N_14358,N_13334,N_13224);
nand U14359 (N_14359,N_13197,N_12610);
xor U14360 (N_14360,N_13358,N_12960);
and U14361 (N_14361,N_12282,N_12482);
xnor U14362 (N_14362,N_12074,N_12306);
and U14363 (N_14363,N_13211,N_13364);
and U14364 (N_14364,N_12229,N_13257);
xor U14365 (N_14365,N_13462,N_13152);
xnor U14366 (N_14366,N_12871,N_12336);
or U14367 (N_14367,N_12740,N_13148);
xnor U14368 (N_14368,N_12103,N_12005);
and U14369 (N_14369,N_12084,N_12181);
and U14370 (N_14370,N_13067,N_12361);
xnor U14371 (N_14371,N_12197,N_13246);
xnor U14372 (N_14372,N_12699,N_12518);
or U14373 (N_14373,N_12461,N_12844);
xnor U14374 (N_14374,N_13360,N_12484);
and U14375 (N_14375,N_12772,N_13299);
nand U14376 (N_14376,N_12453,N_13118);
nand U14377 (N_14377,N_12433,N_12719);
or U14378 (N_14378,N_13498,N_12457);
nand U14379 (N_14379,N_12271,N_13442);
and U14380 (N_14380,N_12299,N_12494);
or U14381 (N_14381,N_12644,N_13146);
nand U14382 (N_14382,N_13055,N_13033);
xor U14383 (N_14383,N_13082,N_12379);
xor U14384 (N_14384,N_13174,N_12318);
nor U14385 (N_14385,N_13295,N_12029);
nor U14386 (N_14386,N_13464,N_13022);
nor U14387 (N_14387,N_13158,N_13443);
xnor U14388 (N_14388,N_12601,N_12142);
or U14389 (N_14389,N_12028,N_12020);
nand U14390 (N_14390,N_12593,N_12992);
and U14391 (N_14391,N_12872,N_13371);
and U14392 (N_14392,N_12838,N_13221);
nor U14393 (N_14393,N_12853,N_12173);
or U14394 (N_14394,N_13130,N_12278);
and U14395 (N_14395,N_12218,N_12476);
and U14396 (N_14396,N_13361,N_13441);
or U14397 (N_14397,N_12304,N_13097);
xnor U14398 (N_14398,N_12009,N_13255);
xor U14399 (N_14399,N_13477,N_12515);
nand U14400 (N_14400,N_12492,N_12667);
nand U14401 (N_14401,N_12945,N_12917);
nor U14402 (N_14402,N_12035,N_12400);
xor U14403 (N_14403,N_12756,N_12458);
nand U14404 (N_14404,N_12572,N_12753);
nor U14405 (N_14405,N_12575,N_12721);
and U14406 (N_14406,N_12888,N_12538);
nor U14407 (N_14407,N_12906,N_12008);
nand U14408 (N_14408,N_13168,N_12301);
nor U14409 (N_14409,N_12586,N_12993);
or U14410 (N_14410,N_12839,N_13057);
nand U14411 (N_14411,N_13121,N_13228);
nand U14412 (N_14412,N_13452,N_12492);
or U14413 (N_14413,N_12243,N_13309);
nand U14414 (N_14414,N_13021,N_12287);
xnor U14415 (N_14415,N_12583,N_12116);
and U14416 (N_14416,N_12340,N_12342);
xnor U14417 (N_14417,N_12981,N_12525);
or U14418 (N_14418,N_12507,N_13153);
xnor U14419 (N_14419,N_12298,N_12989);
nor U14420 (N_14420,N_13072,N_12425);
nor U14421 (N_14421,N_13005,N_13241);
or U14422 (N_14422,N_12772,N_13062);
nor U14423 (N_14423,N_12454,N_12431);
xnor U14424 (N_14424,N_13272,N_12119);
nor U14425 (N_14425,N_12374,N_12061);
xor U14426 (N_14426,N_13497,N_13233);
xor U14427 (N_14427,N_12710,N_13412);
or U14428 (N_14428,N_12802,N_12031);
xnor U14429 (N_14429,N_13407,N_12293);
and U14430 (N_14430,N_13453,N_13343);
xnor U14431 (N_14431,N_12102,N_12092);
xor U14432 (N_14432,N_13002,N_12095);
and U14433 (N_14433,N_13328,N_13387);
nor U14434 (N_14434,N_12958,N_12488);
nor U14435 (N_14435,N_13358,N_12435);
or U14436 (N_14436,N_13221,N_12936);
and U14437 (N_14437,N_12426,N_13123);
nand U14438 (N_14438,N_12724,N_13303);
nand U14439 (N_14439,N_13251,N_12851);
or U14440 (N_14440,N_12906,N_13139);
nor U14441 (N_14441,N_13205,N_12273);
or U14442 (N_14442,N_12037,N_12671);
or U14443 (N_14443,N_12624,N_12511);
nor U14444 (N_14444,N_13440,N_13030);
and U14445 (N_14445,N_12875,N_13392);
nor U14446 (N_14446,N_13153,N_12830);
and U14447 (N_14447,N_12565,N_12228);
nor U14448 (N_14448,N_12710,N_12161);
or U14449 (N_14449,N_12317,N_12990);
xnor U14450 (N_14450,N_12950,N_13257);
or U14451 (N_14451,N_12650,N_12330);
and U14452 (N_14452,N_13274,N_12763);
or U14453 (N_14453,N_13129,N_12098);
xor U14454 (N_14454,N_12726,N_12033);
nor U14455 (N_14455,N_13111,N_12960);
nand U14456 (N_14456,N_12477,N_12061);
xnor U14457 (N_14457,N_12165,N_12302);
nand U14458 (N_14458,N_12999,N_12234);
nor U14459 (N_14459,N_13283,N_13030);
nor U14460 (N_14460,N_12641,N_12374);
nand U14461 (N_14461,N_13234,N_12415);
nor U14462 (N_14462,N_12389,N_13424);
or U14463 (N_14463,N_12045,N_12554);
or U14464 (N_14464,N_12045,N_12578);
nor U14465 (N_14465,N_13447,N_12821);
or U14466 (N_14466,N_12032,N_13485);
xor U14467 (N_14467,N_12767,N_12763);
and U14468 (N_14468,N_12459,N_13211);
nor U14469 (N_14469,N_13187,N_12318);
nor U14470 (N_14470,N_12434,N_12814);
nor U14471 (N_14471,N_12874,N_12437);
nand U14472 (N_14472,N_12350,N_13489);
nor U14473 (N_14473,N_12935,N_13046);
nand U14474 (N_14474,N_12225,N_13339);
nand U14475 (N_14475,N_12793,N_12662);
and U14476 (N_14476,N_12489,N_12325);
and U14477 (N_14477,N_12277,N_13376);
xor U14478 (N_14478,N_13097,N_12007);
nand U14479 (N_14479,N_12434,N_12656);
nand U14480 (N_14480,N_12372,N_12221);
xnor U14481 (N_14481,N_12582,N_12170);
nor U14482 (N_14482,N_13363,N_12483);
and U14483 (N_14483,N_13216,N_12295);
nand U14484 (N_14484,N_12599,N_13319);
nand U14485 (N_14485,N_13346,N_12263);
nor U14486 (N_14486,N_13231,N_12650);
nor U14487 (N_14487,N_13365,N_13360);
xnor U14488 (N_14488,N_12843,N_13486);
xnor U14489 (N_14489,N_12021,N_12700);
xnor U14490 (N_14490,N_12318,N_12878);
nor U14491 (N_14491,N_12002,N_13436);
nor U14492 (N_14492,N_12573,N_12130);
nor U14493 (N_14493,N_12213,N_13402);
nor U14494 (N_14494,N_12568,N_12459);
and U14495 (N_14495,N_12268,N_12011);
or U14496 (N_14496,N_13254,N_12232);
nand U14497 (N_14497,N_12660,N_13263);
nor U14498 (N_14498,N_12959,N_12404);
and U14499 (N_14499,N_13463,N_12069);
nor U14500 (N_14500,N_12688,N_13079);
nor U14501 (N_14501,N_13161,N_12958);
and U14502 (N_14502,N_12612,N_13313);
and U14503 (N_14503,N_12017,N_12046);
or U14504 (N_14504,N_13004,N_12500);
nor U14505 (N_14505,N_12495,N_12117);
and U14506 (N_14506,N_12705,N_12163);
nor U14507 (N_14507,N_12435,N_13374);
xnor U14508 (N_14508,N_13339,N_12155);
nor U14509 (N_14509,N_13104,N_12441);
xnor U14510 (N_14510,N_12608,N_13071);
and U14511 (N_14511,N_12487,N_13160);
or U14512 (N_14512,N_13397,N_12045);
and U14513 (N_14513,N_13393,N_12927);
nor U14514 (N_14514,N_12949,N_12210);
or U14515 (N_14515,N_12482,N_12139);
nand U14516 (N_14516,N_12777,N_12404);
or U14517 (N_14517,N_12452,N_12360);
or U14518 (N_14518,N_12686,N_13395);
xor U14519 (N_14519,N_12011,N_13406);
or U14520 (N_14520,N_12475,N_13191);
nor U14521 (N_14521,N_12793,N_12082);
and U14522 (N_14522,N_12034,N_13367);
or U14523 (N_14523,N_12904,N_13386);
and U14524 (N_14524,N_12558,N_12283);
or U14525 (N_14525,N_12487,N_13390);
nor U14526 (N_14526,N_12731,N_12755);
nand U14527 (N_14527,N_12411,N_13109);
and U14528 (N_14528,N_12850,N_12244);
or U14529 (N_14529,N_12910,N_12203);
nand U14530 (N_14530,N_12261,N_12628);
nand U14531 (N_14531,N_12775,N_12063);
or U14532 (N_14532,N_12566,N_12162);
or U14533 (N_14533,N_13316,N_12981);
and U14534 (N_14534,N_12682,N_12949);
xnor U14535 (N_14535,N_13420,N_12233);
xnor U14536 (N_14536,N_12603,N_13410);
xor U14537 (N_14537,N_12208,N_13458);
nand U14538 (N_14538,N_13203,N_12026);
nor U14539 (N_14539,N_12444,N_12796);
nor U14540 (N_14540,N_13427,N_13447);
or U14541 (N_14541,N_12363,N_13408);
xor U14542 (N_14542,N_13305,N_13456);
nor U14543 (N_14543,N_13229,N_12848);
xor U14544 (N_14544,N_12456,N_12472);
and U14545 (N_14545,N_12390,N_12475);
xor U14546 (N_14546,N_13139,N_12242);
and U14547 (N_14547,N_12006,N_12852);
or U14548 (N_14548,N_12869,N_12097);
and U14549 (N_14549,N_12881,N_13494);
nand U14550 (N_14550,N_13018,N_12298);
xnor U14551 (N_14551,N_12756,N_13301);
nand U14552 (N_14552,N_13239,N_13157);
nor U14553 (N_14553,N_12316,N_13430);
or U14554 (N_14554,N_12196,N_13205);
nand U14555 (N_14555,N_13174,N_12791);
xor U14556 (N_14556,N_13306,N_12584);
nor U14557 (N_14557,N_12048,N_12224);
and U14558 (N_14558,N_12514,N_12508);
nor U14559 (N_14559,N_12044,N_12106);
nand U14560 (N_14560,N_13129,N_12448);
xor U14561 (N_14561,N_12555,N_13055);
and U14562 (N_14562,N_12930,N_12362);
nand U14563 (N_14563,N_13319,N_13255);
nand U14564 (N_14564,N_13044,N_12800);
or U14565 (N_14565,N_13011,N_13121);
xor U14566 (N_14566,N_13181,N_12821);
nand U14567 (N_14567,N_12530,N_13275);
xnor U14568 (N_14568,N_12888,N_12021);
or U14569 (N_14569,N_12482,N_12534);
nor U14570 (N_14570,N_13270,N_12414);
xor U14571 (N_14571,N_13225,N_12661);
xnor U14572 (N_14572,N_12993,N_13163);
xnor U14573 (N_14573,N_13285,N_12703);
nand U14574 (N_14574,N_12977,N_12996);
xnor U14575 (N_14575,N_13454,N_12623);
nor U14576 (N_14576,N_12765,N_12110);
and U14577 (N_14577,N_13065,N_12085);
and U14578 (N_14578,N_13377,N_13111);
or U14579 (N_14579,N_13390,N_12027);
nand U14580 (N_14580,N_12739,N_13129);
and U14581 (N_14581,N_12955,N_13327);
nor U14582 (N_14582,N_13106,N_13211);
nor U14583 (N_14583,N_12327,N_12089);
nand U14584 (N_14584,N_12832,N_13395);
and U14585 (N_14585,N_12845,N_12909);
xor U14586 (N_14586,N_13192,N_13232);
and U14587 (N_14587,N_12960,N_13146);
xnor U14588 (N_14588,N_12760,N_13113);
xnor U14589 (N_14589,N_12747,N_12341);
and U14590 (N_14590,N_12195,N_12171);
xor U14591 (N_14591,N_12168,N_12156);
xnor U14592 (N_14592,N_13367,N_13355);
or U14593 (N_14593,N_12424,N_12791);
xnor U14594 (N_14594,N_12192,N_13467);
or U14595 (N_14595,N_12843,N_13223);
or U14596 (N_14596,N_12432,N_12395);
nand U14597 (N_14597,N_12470,N_12015);
or U14598 (N_14598,N_13440,N_13424);
nor U14599 (N_14599,N_13488,N_12115);
and U14600 (N_14600,N_12467,N_13208);
and U14601 (N_14601,N_12636,N_12952);
nand U14602 (N_14602,N_12775,N_12409);
and U14603 (N_14603,N_12923,N_12941);
nor U14604 (N_14604,N_12569,N_13449);
or U14605 (N_14605,N_12362,N_12077);
and U14606 (N_14606,N_12781,N_12791);
nor U14607 (N_14607,N_12979,N_12680);
nand U14608 (N_14608,N_12055,N_12553);
and U14609 (N_14609,N_12053,N_12240);
nand U14610 (N_14610,N_13310,N_12104);
nand U14611 (N_14611,N_12879,N_12675);
nor U14612 (N_14612,N_12529,N_12842);
nand U14613 (N_14613,N_12588,N_12101);
xor U14614 (N_14614,N_12104,N_13287);
nor U14615 (N_14615,N_12624,N_12128);
nor U14616 (N_14616,N_13101,N_13018);
or U14617 (N_14617,N_12691,N_12781);
nor U14618 (N_14618,N_12753,N_13460);
nand U14619 (N_14619,N_13014,N_13096);
nand U14620 (N_14620,N_12090,N_13058);
or U14621 (N_14621,N_12323,N_12434);
or U14622 (N_14622,N_12558,N_12113);
nor U14623 (N_14623,N_13387,N_12483);
or U14624 (N_14624,N_12333,N_12021);
and U14625 (N_14625,N_12578,N_12863);
and U14626 (N_14626,N_12549,N_12380);
xor U14627 (N_14627,N_13195,N_12178);
nor U14628 (N_14628,N_12887,N_13357);
nand U14629 (N_14629,N_13439,N_12997);
xnor U14630 (N_14630,N_12285,N_13064);
nor U14631 (N_14631,N_13069,N_13065);
and U14632 (N_14632,N_13442,N_12757);
and U14633 (N_14633,N_13476,N_13179);
and U14634 (N_14634,N_12315,N_12328);
nand U14635 (N_14635,N_13141,N_12218);
or U14636 (N_14636,N_13121,N_13227);
nor U14637 (N_14637,N_12906,N_12901);
nand U14638 (N_14638,N_13247,N_13452);
nand U14639 (N_14639,N_12682,N_13413);
nand U14640 (N_14640,N_12619,N_12830);
and U14641 (N_14641,N_12731,N_12170);
nand U14642 (N_14642,N_12522,N_13319);
or U14643 (N_14643,N_12007,N_13322);
nand U14644 (N_14644,N_13329,N_12043);
nor U14645 (N_14645,N_12950,N_12311);
nand U14646 (N_14646,N_12979,N_13413);
nor U14647 (N_14647,N_13449,N_12882);
nand U14648 (N_14648,N_13194,N_13181);
or U14649 (N_14649,N_12916,N_13315);
nor U14650 (N_14650,N_12186,N_12325);
or U14651 (N_14651,N_12480,N_12371);
nor U14652 (N_14652,N_13117,N_13145);
nand U14653 (N_14653,N_12827,N_13175);
xnor U14654 (N_14654,N_12002,N_12363);
xnor U14655 (N_14655,N_12892,N_13315);
or U14656 (N_14656,N_13251,N_13086);
xor U14657 (N_14657,N_13196,N_12759);
nand U14658 (N_14658,N_12058,N_13473);
nor U14659 (N_14659,N_12880,N_12740);
nor U14660 (N_14660,N_12284,N_12424);
and U14661 (N_14661,N_13453,N_13430);
nor U14662 (N_14662,N_13367,N_12861);
xor U14663 (N_14663,N_12087,N_13335);
or U14664 (N_14664,N_12588,N_12914);
nand U14665 (N_14665,N_13152,N_13135);
xor U14666 (N_14666,N_12964,N_12140);
nor U14667 (N_14667,N_12019,N_12398);
xnor U14668 (N_14668,N_12498,N_12740);
xor U14669 (N_14669,N_13381,N_12769);
nand U14670 (N_14670,N_12951,N_12375);
nor U14671 (N_14671,N_13379,N_12350);
or U14672 (N_14672,N_12773,N_12277);
nor U14673 (N_14673,N_12856,N_12268);
nand U14674 (N_14674,N_12127,N_12527);
and U14675 (N_14675,N_13384,N_12876);
nand U14676 (N_14676,N_13391,N_12070);
or U14677 (N_14677,N_12649,N_12421);
xor U14678 (N_14678,N_12264,N_13476);
or U14679 (N_14679,N_12480,N_12059);
or U14680 (N_14680,N_12478,N_12816);
xnor U14681 (N_14681,N_13147,N_12421);
or U14682 (N_14682,N_12414,N_12008);
and U14683 (N_14683,N_12473,N_12357);
nor U14684 (N_14684,N_12301,N_12050);
xor U14685 (N_14685,N_12614,N_13017);
or U14686 (N_14686,N_12108,N_13392);
xor U14687 (N_14687,N_12752,N_12388);
or U14688 (N_14688,N_12238,N_12842);
and U14689 (N_14689,N_12209,N_12720);
xnor U14690 (N_14690,N_12146,N_12914);
and U14691 (N_14691,N_12453,N_12809);
and U14692 (N_14692,N_13126,N_13353);
nand U14693 (N_14693,N_12973,N_12969);
or U14694 (N_14694,N_12166,N_12230);
nand U14695 (N_14695,N_12670,N_12750);
nand U14696 (N_14696,N_12317,N_12739);
or U14697 (N_14697,N_13331,N_12860);
and U14698 (N_14698,N_13327,N_13187);
xor U14699 (N_14699,N_12567,N_12713);
nor U14700 (N_14700,N_13442,N_13196);
nor U14701 (N_14701,N_12645,N_12320);
nand U14702 (N_14702,N_12038,N_13270);
nor U14703 (N_14703,N_12421,N_12039);
or U14704 (N_14704,N_12728,N_12425);
or U14705 (N_14705,N_12181,N_12711);
and U14706 (N_14706,N_12282,N_12815);
nand U14707 (N_14707,N_13436,N_13489);
nor U14708 (N_14708,N_12238,N_12318);
or U14709 (N_14709,N_13150,N_12908);
nand U14710 (N_14710,N_13037,N_12649);
or U14711 (N_14711,N_12140,N_12499);
and U14712 (N_14712,N_12358,N_13293);
xor U14713 (N_14713,N_12468,N_12049);
nand U14714 (N_14714,N_12740,N_13196);
and U14715 (N_14715,N_12544,N_12491);
or U14716 (N_14716,N_12626,N_13198);
nand U14717 (N_14717,N_13478,N_12976);
nand U14718 (N_14718,N_12024,N_13439);
or U14719 (N_14719,N_12303,N_13125);
nand U14720 (N_14720,N_13468,N_12642);
and U14721 (N_14721,N_13407,N_13207);
nor U14722 (N_14722,N_13386,N_12380);
xor U14723 (N_14723,N_12658,N_13445);
or U14724 (N_14724,N_12444,N_13134);
or U14725 (N_14725,N_12741,N_12772);
xor U14726 (N_14726,N_12904,N_13116);
and U14727 (N_14727,N_12921,N_12071);
nand U14728 (N_14728,N_13461,N_12194);
xor U14729 (N_14729,N_12656,N_12760);
and U14730 (N_14730,N_12736,N_13391);
or U14731 (N_14731,N_12814,N_13270);
nand U14732 (N_14732,N_12975,N_12418);
xor U14733 (N_14733,N_12490,N_13141);
nor U14734 (N_14734,N_12917,N_12075);
and U14735 (N_14735,N_12451,N_12433);
and U14736 (N_14736,N_12273,N_12731);
nor U14737 (N_14737,N_12140,N_13203);
or U14738 (N_14738,N_13246,N_12363);
and U14739 (N_14739,N_13069,N_12813);
xnor U14740 (N_14740,N_12081,N_12180);
and U14741 (N_14741,N_13247,N_12152);
nand U14742 (N_14742,N_12670,N_13386);
nand U14743 (N_14743,N_12006,N_12649);
or U14744 (N_14744,N_13166,N_12802);
xor U14745 (N_14745,N_12214,N_13119);
nand U14746 (N_14746,N_12795,N_12574);
xor U14747 (N_14747,N_12227,N_12394);
or U14748 (N_14748,N_12807,N_12486);
and U14749 (N_14749,N_12763,N_12646);
xor U14750 (N_14750,N_13020,N_12347);
and U14751 (N_14751,N_12984,N_12453);
nand U14752 (N_14752,N_12647,N_12859);
or U14753 (N_14753,N_12611,N_12405);
nand U14754 (N_14754,N_12400,N_12738);
nand U14755 (N_14755,N_13431,N_12301);
nor U14756 (N_14756,N_12528,N_13221);
and U14757 (N_14757,N_12730,N_13406);
nor U14758 (N_14758,N_13090,N_12561);
xnor U14759 (N_14759,N_12400,N_12440);
or U14760 (N_14760,N_12359,N_13258);
xnor U14761 (N_14761,N_13353,N_13225);
xnor U14762 (N_14762,N_12626,N_13472);
nand U14763 (N_14763,N_12694,N_12788);
or U14764 (N_14764,N_13470,N_13086);
nand U14765 (N_14765,N_12492,N_13102);
nor U14766 (N_14766,N_12733,N_13113);
and U14767 (N_14767,N_13084,N_12011);
and U14768 (N_14768,N_12035,N_12766);
xnor U14769 (N_14769,N_13401,N_12400);
xor U14770 (N_14770,N_12238,N_13074);
or U14771 (N_14771,N_12158,N_12756);
or U14772 (N_14772,N_12655,N_13187);
or U14773 (N_14773,N_12267,N_13435);
or U14774 (N_14774,N_12146,N_12039);
nand U14775 (N_14775,N_12921,N_13293);
nand U14776 (N_14776,N_12803,N_12653);
nand U14777 (N_14777,N_13220,N_12104);
nor U14778 (N_14778,N_13196,N_12559);
or U14779 (N_14779,N_12230,N_13083);
or U14780 (N_14780,N_13186,N_12060);
and U14781 (N_14781,N_13053,N_13174);
nor U14782 (N_14782,N_12021,N_13295);
nor U14783 (N_14783,N_12345,N_12715);
and U14784 (N_14784,N_13466,N_12394);
and U14785 (N_14785,N_12734,N_12344);
nand U14786 (N_14786,N_12548,N_12500);
nand U14787 (N_14787,N_12716,N_12500);
xor U14788 (N_14788,N_13037,N_12856);
and U14789 (N_14789,N_12930,N_12635);
nand U14790 (N_14790,N_12626,N_12937);
and U14791 (N_14791,N_12468,N_12738);
or U14792 (N_14792,N_12231,N_12639);
or U14793 (N_14793,N_13298,N_12701);
xor U14794 (N_14794,N_12841,N_12211);
or U14795 (N_14795,N_12305,N_12545);
xnor U14796 (N_14796,N_12005,N_13298);
and U14797 (N_14797,N_12777,N_13358);
nand U14798 (N_14798,N_12044,N_12691);
and U14799 (N_14799,N_13241,N_13222);
and U14800 (N_14800,N_13406,N_12550);
nand U14801 (N_14801,N_12335,N_12007);
or U14802 (N_14802,N_12004,N_13401);
xor U14803 (N_14803,N_12029,N_13284);
nand U14804 (N_14804,N_12968,N_12494);
nand U14805 (N_14805,N_12611,N_13327);
and U14806 (N_14806,N_13378,N_12548);
or U14807 (N_14807,N_12386,N_12765);
or U14808 (N_14808,N_12288,N_12600);
xor U14809 (N_14809,N_12723,N_13188);
or U14810 (N_14810,N_12163,N_13029);
nor U14811 (N_14811,N_12330,N_12271);
nor U14812 (N_14812,N_13388,N_12005);
xnor U14813 (N_14813,N_13310,N_13475);
and U14814 (N_14814,N_12045,N_12970);
or U14815 (N_14815,N_12180,N_12657);
or U14816 (N_14816,N_13306,N_12280);
nand U14817 (N_14817,N_12417,N_12163);
nor U14818 (N_14818,N_12943,N_12292);
nand U14819 (N_14819,N_13443,N_13173);
nor U14820 (N_14820,N_12944,N_12616);
or U14821 (N_14821,N_13424,N_13446);
nor U14822 (N_14822,N_12167,N_13308);
and U14823 (N_14823,N_13142,N_12928);
or U14824 (N_14824,N_13055,N_12950);
xor U14825 (N_14825,N_12415,N_13049);
nor U14826 (N_14826,N_13099,N_12487);
nor U14827 (N_14827,N_13315,N_12893);
or U14828 (N_14828,N_12931,N_12523);
and U14829 (N_14829,N_12384,N_12998);
and U14830 (N_14830,N_12946,N_12304);
nor U14831 (N_14831,N_12605,N_12641);
xnor U14832 (N_14832,N_13091,N_12390);
nor U14833 (N_14833,N_12497,N_12667);
nand U14834 (N_14834,N_13411,N_13284);
nor U14835 (N_14835,N_12369,N_12239);
or U14836 (N_14836,N_12351,N_12937);
nand U14837 (N_14837,N_12756,N_13184);
or U14838 (N_14838,N_12220,N_12560);
nor U14839 (N_14839,N_12588,N_13251);
nor U14840 (N_14840,N_13481,N_13484);
and U14841 (N_14841,N_12165,N_13172);
nand U14842 (N_14842,N_12866,N_12191);
nor U14843 (N_14843,N_12191,N_13324);
or U14844 (N_14844,N_13006,N_13024);
and U14845 (N_14845,N_12326,N_12073);
nor U14846 (N_14846,N_12192,N_12762);
xnor U14847 (N_14847,N_13431,N_12742);
nand U14848 (N_14848,N_13297,N_13153);
nor U14849 (N_14849,N_13308,N_12195);
or U14850 (N_14850,N_13234,N_12329);
nand U14851 (N_14851,N_12236,N_12781);
and U14852 (N_14852,N_12973,N_12799);
nor U14853 (N_14853,N_13447,N_13391);
nand U14854 (N_14854,N_13331,N_13418);
nand U14855 (N_14855,N_12075,N_13102);
xnor U14856 (N_14856,N_12098,N_13101);
nand U14857 (N_14857,N_13105,N_13387);
xnor U14858 (N_14858,N_12366,N_12569);
and U14859 (N_14859,N_12310,N_13077);
and U14860 (N_14860,N_12560,N_13319);
and U14861 (N_14861,N_12204,N_13382);
nand U14862 (N_14862,N_12573,N_12937);
xor U14863 (N_14863,N_12660,N_13051);
and U14864 (N_14864,N_12002,N_12657);
nand U14865 (N_14865,N_12751,N_12395);
xnor U14866 (N_14866,N_12462,N_12403);
nor U14867 (N_14867,N_12578,N_12010);
nor U14868 (N_14868,N_13281,N_12552);
and U14869 (N_14869,N_12182,N_12762);
xor U14870 (N_14870,N_12221,N_12230);
and U14871 (N_14871,N_12998,N_12829);
and U14872 (N_14872,N_12661,N_12049);
and U14873 (N_14873,N_13319,N_13428);
nor U14874 (N_14874,N_13010,N_12367);
xnor U14875 (N_14875,N_13286,N_13041);
nand U14876 (N_14876,N_12559,N_12938);
xor U14877 (N_14877,N_12495,N_13177);
or U14878 (N_14878,N_13365,N_13489);
xor U14879 (N_14879,N_12409,N_12317);
nor U14880 (N_14880,N_12879,N_12730);
or U14881 (N_14881,N_12861,N_12654);
xnor U14882 (N_14882,N_12060,N_13027);
nor U14883 (N_14883,N_12694,N_12617);
or U14884 (N_14884,N_12307,N_13352);
nor U14885 (N_14885,N_13405,N_13298);
or U14886 (N_14886,N_13029,N_12907);
nor U14887 (N_14887,N_12867,N_13446);
nand U14888 (N_14888,N_12776,N_12745);
or U14889 (N_14889,N_13051,N_12688);
or U14890 (N_14890,N_13215,N_13422);
nand U14891 (N_14891,N_13099,N_13344);
and U14892 (N_14892,N_13042,N_12483);
and U14893 (N_14893,N_13203,N_12128);
nor U14894 (N_14894,N_12380,N_12139);
nand U14895 (N_14895,N_13418,N_12533);
or U14896 (N_14896,N_13368,N_12830);
nor U14897 (N_14897,N_12786,N_13433);
xnor U14898 (N_14898,N_12406,N_12586);
xnor U14899 (N_14899,N_12271,N_12505);
or U14900 (N_14900,N_13347,N_13331);
nor U14901 (N_14901,N_12768,N_12896);
xnor U14902 (N_14902,N_12043,N_12108);
xor U14903 (N_14903,N_12484,N_13199);
nor U14904 (N_14904,N_13230,N_13148);
or U14905 (N_14905,N_12877,N_12260);
xnor U14906 (N_14906,N_12214,N_12983);
and U14907 (N_14907,N_12891,N_12262);
and U14908 (N_14908,N_12588,N_12700);
nand U14909 (N_14909,N_13260,N_12474);
xor U14910 (N_14910,N_12128,N_12695);
nor U14911 (N_14911,N_13092,N_12577);
and U14912 (N_14912,N_12946,N_13245);
xor U14913 (N_14913,N_12073,N_12490);
xnor U14914 (N_14914,N_13131,N_13355);
nor U14915 (N_14915,N_12338,N_13473);
and U14916 (N_14916,N_12678,N_13104);
nand U14917 (N_14917,N_13315,N_12639);
and U14918 (N_14918,N_13362,N_12986);
xor U14919 (N_14919,N_12034,N_13287);
xnor U14920 (N_14920,N_13079,N_12374);
xor U14921 (N_14921,N_12361,N_12593);
or U14922 (N_14922,N_12432,N_12437);
nor U14923 (N_14923,N_12463,N_12623);
nor U14924 (N_14924,N_12047,N_12454);
nand U14925 (N_14925,N_13014,N_13350);
xnor U14926 (N_14926,N_13394,N_12005);
or U14927 (N_14927,N_13295,N_12518);
nor U14928 (N_14928,N_12771,N_12185);
nand U14929 (N_14929,N_13445,N_12495);
xor U14930 (N_14930,N_12627,N_12687);
nand U14931 (N_14931,N_12389,N_12853);
nand U14932 (N_14932,N_12319,N_12642);
nor U14933 (N_14933,N_12335,N_13262);
or U14934 (N_14934,N_12824,N_13017);
and U14935 (N_14935,N_12451,N_13161);
or U14936 (N_14936,N_12815,N_12533);
or U14937 (N_14937,N_12463,N_13027);
and U14938 (N_14938,N_13027,N_12768);
and U14939 (N_14939,N_12752,N_12139);
and U14940 (N_14940,N_12813,N_12717);
and U14941 (N_14941,N_13089,N_12346);
xor U14942 (N_14942,N_13439,N_12533);
nor U14943 (N_14943,N_12006,N_12247);
nand U14944 (N_14944,N_12043,N_12231);
and U14945 (N_14945,N_13120,N_12178);
nor U14946 (N_14946,N_13369,N_13364);
or U14947 (N_14947,N_13329,N_12213);
or U14948 (N_14948,N_13283,N_13209);
xnor U14949 (N_14949,N_12292,N_12845);
nand U14950 (N_14950,N_12611,N_13399);
and U14951 (N_14951,N_13019,N_13049);
and U14952 (N_14952,N_12859,N_12338);
and U14953 (N_14953,N_12813,N_13168);
nor U14954 (N_14954,N_12006,N_13298);
xnor U14955 (N_14955,N_12936,N_12192);
nand U14956 (N_14956,N_13142,N_13358);
or U14957 (N_14957,N_12598,N_13112);
and U14958 (N_14958,N_12204,N_12361);
or U14959 (N_14959,N_12400,N_13385);
nand U14960 (N_14960,N_12679,N_13494);
or U14961 (N_14961,N_13428,N_12687);
nand U14962 (N_14962,N_12405,N_12261);
xor U14963 (N_14963,N_12185,N_12205);
nor U14964 (N_14964,N_12221,N_12515);
nor U14965 (N_14965,N_13320,N_12459);
nor U14966 (N_14966,N_12940,N_13474);
or U14967 (N_14967,N_12841,N_12506);
or U14968 (N_14968,N_13086,N_12414);
nand U14969 (N_14969,N_13260,N_13240);
or U14970 (N_14970,N_12576,N_13116);
or U14971 (N_14971,N_12638,N_12441);
nand U14972 (N_14972,N_12646,N_12095);
and U14973 (N_14973,N_13228,N_12909);
and U14974 (N_14974,N_12776,N_13193);
nor U14975 (N_14975,N_12692,N_12306);
xor U14976 (N_14976,N_12389,N_12217);
nor U14977 (N_14977,N_12914,N_12222);
or U14978 (N_14978,N_12176,N_12079);
xor U14979 (N_14979,N_12696,N_13361);
xor U14980 (N_14980,N_13167,N_12689);
nand U14981 (N_14981,N_12387,N_12148);
or U14982 (N_14982,N_13293,N_13136);
or U14983 (N_14983,N_12332,N_12252);
nor U14984 (N_14984,N_13016,N_12516);
xor U14985 (N_14985,N_13159,N_13477);
or U14986 (N_14986,N_12124,N_13160);
and U14987 (N_14987,N_12801,N_12955);
xor U14988 (N_14988,N_12856,N_12091);
xnor U14989 (N_14989,N_12288,N_12413);
or U14990 (N_14990,N_12408,N_13433);
xor U14991 (N_14991,N_12037,N_13371);
xor U14992 (N_14992,N_13191,N_13449);
or U14993 (N_14993,N_12371,N_12030);
xor U14994 (N_14994,N_12474,N_12772);
nand U14995 (N_14995,N_13043,N_12817);
and U14996 (N_14996,N_13015,N_12279);
xor U14997 (N_14997,N_12804,N_13431);
and U14998 (N_14998,N_12756,N_12916);
nand U14999 (N_14999,N_13098,N_12711);
or UO_0 (O_0,N_14296,N_13618);
nor UO_1 (O_1,N_14096,N_14436);
xor UO_2 (O_2,N_13605,N_13651);
and UO_3 (O_3,N_14023,N_14622);
or UO_4 (O_4,N_14947,N_14599);
and UO_5 (O_5,N_13715,N_14458);
nor UO_6 (O_6,N_13761,N_14791);
nand UO_7 (O_7,N_13552,N_14564);
or UO_8 (O_8,N_14790,N_13892);
xor UO_9 (O_9,N_14219,N_14794);
or UO_10 (O_10,N_13989,N_14169);
or UO_11 (O_11,N_13908,N_14984);
nand UO_12 (O_12,N_14154,N_14756);
and UO_13 (O_13,N_14185,N_13671);
and UO_14 (O_14,N_13551,N_14806);
or UO_15 (O_15,N_14781,N_13673);
xnor UO_16 (O_16,N_14855,N_13562);
xnor UO_17 (O_17,N_14635,N_13950);
or UO_18 (O_18,N_14242,N_14792);
xor UO_19 (O_19,N_14659,N_13676);
nand UO_20 (O_20,N_13530,N_13579);
or UO_21 (O_21,N_13884,N_14042);
and UO_22 (O_22,N_14885,N_14537);
or UO_23 (O_23,N_13544,N_14893);
nor UO_24 (O_24,N_13799,N_14646);
xnor UO_25 (O_25,N_14064,N_14645);
nor UO_26 (O_26,N_14186,N_13636);
and UO_27 (O_27,N_13569,N_14323);
or UO_28 (O_28,N_14448,N_14009);
nor UO_29 (O_29,N_13638,N_13762);
and UO_30 (O_30,N_13999,N_13670);
nor UO_31 (O_31,N_13918,N_13801);
xor UO_32 (O_32,N_14500,N_14467);
nand UO_33 (O_33,N_14766,N_14069);
nor UO_34 (O_34,N_14521,N_14632);
xor UO_35 (O_35,N_13888,N_14229);
xnor UO_36 (O_36,N_14492,N_14471);
nor UO_37 (O_37,N_14502,N_14801);
or UO_38 (O_38,N_14285,N_14593);
and UO_39 (O_39,N_14282,N_13534);
or UO_40 (O_40,N_14385,N_13533);
xnor UO_41 (O_41,N_14916,N_14359);
xnor UO_42 (O_42,N_13719,N_13850);
xnor UO_43 (O_43,N_13927,N_14432);
or UO_44 (O_44,N_13868,N_14162);
xnor UO_45 (O_45,N_14172,N_14279);
or UO_46 (O_46,N_13933,N_14625);
nand UO_47 (O_47,N_14929,N_14444);
nor UO_48 (O_48,N_14982,N_14913);
nor UO_49 (O_49,N_14741,N_14680);
nand UO_50 (O_50,N_14433,N_14900);
nand UO_51 (O_51,N_14311,N_14674);
xor UO_52 (O_52,N_14539,N_14032);
or UO_53 (O_53,N_14991,N_14053);
and UO_54 (O_54,N_14063,N_14968);
xnor UO_55 (O_55,N_13856,N_13866);
nand UO_56 (O_56,N_14895,N_14113);
xnor UO_57 (O_57,N_14335,N_13796);
nand UO_58 (O_58,N_14347,N_14945);
and UO_59 (O_59,N_14591,N_14764);
nor UO_60 (O_60,N_14160,N_14253);
or UO_61 (O_61,N_14179,N_14938);
or UO_62 (O_62,N_13855,N_13596);
nand UO_63 (O_63,N_13541,N_14284);
nor UO_64 (O_64,N_14408,N_14830);
and UO_65 (O_65,N_13726,N_14532);
nand UO_66 (O_66,N_14905,N_14423);
nor UO_67 (O_67,N_14387,N_14760);
and UO_68 (O_68,N_14623,N_14611);
or UO_69 (O_69,N_14683,N_14030);
and UO_70 (O_70,N_14731,N_13641);
and UO_71 (O_71,N_13967,N_14758);
and UO_72 (O_72,N_14986,N_14034);
or UO_73 (O_73,N_14519,N_14059);
nor UO_74 (O_74,N_14515,N_13519);
or UO_75 (O_75,N_14943,N_14782);
xnor UO_76 (O_76,N_13807,N_14051);
or UO_77 (O_77,N_13996,N_14907);
nor UO_78 (O_78,N_14850,N_14803);
xnor UO_79 (O_79,N_14545,N_14001);
or UO_80 (O_80,N_14999,N_14283);
and UO_81 (O_81,N_13897,N_14522);
or UO_82 (O_82,N_14658,N_14816);
and UO_83 (O_83,N_13827,N_14906);
or UO_84 (O_84,N_14364,N_14925);
and UO_85 (O_85,N_13767,N_14894);
and UO_86 (O_86,N_14411,N_14404);
xnor UO_87 (O_87,N_13987,N_14429);
xor UO_88 (O_88,N_14763,N_14636);
or UO_89 (O_89,N_13830,N_14413);
or UO_90 (O_90,N_14221,N_13704);
nand UO_91 (O_91,N_14431,N_14144);
nand UO_92 (O_92,N_14380,N_14743);
nor UO_93 (O_93,N_14675,N_14990);
xor UO_94 (O_94,N_13648,N_14590);
or UO_95 (O_95,N_13935,N_14010);
nand UO_96 (O_96,N_14812,N_14531);
xnor UO_97 (O_97,N_14464,N_13786);
nand UO_98 (O_98,N_14274,N_14110);
xnor UO_99 (O_99,N_13802,N_14555);
nand UO_100 (O_100,N_14338,N_13581);
xor UO_101 (O_101,N_13733,N_14876);
nor UO_102 (O_102,N_13810,N_14739);
xor UO_103 (O_103,N_14316,N_13904);
xnor UO_104 (O_104,N_14556,N_13711);
xnor UO_105 (O_105,N_13663,N_14256);
nor UO_106 (O_106,N_13886,N_14665);
nor UO_107 (O_107,N_14588,N_14138);
xor UO_108 (O_108,N_14654,N_14871);
nand UO_109 (O_109,N_14414,N_13910);
or UO_110 (O_110,N_13893,N_13805);
nor UO_111 (O_111,N_13858,N_14882);
nand UO_112 (O_112,N_14437,N_14107);
nor UO_113 (O_113,N_13813,N_14570);
nor UO_114 (O_114,N_14852,N_14334);
nand UO_115 (O_115,N_14495,N_13609);
or UO_116 (O_116,N_14994,N_13571);
nand UO_117 (O_117,N_14506,N_14677);
or UO_118 (O_118,N_14525,N_13791);
or UO_119 (O_119,N_14161,N_14238);
nor UO_120 (O_120,N_14972,N_14040);
nand UO_121 (O_121,N_14870,N_14867);
nand UO_122 (O_122,N_14958,N_14027);
nand UO_123 (O_123,N_13578,N_14382);
nand UO_124 (O_124,N_14503,N_14696);
xnor UO_125 (O_125,N_14353,N_13896);
xor UO_126 (O_126,N_14980,N_13765);
and UO_127 (O_127,N_13758,N_14643);
nand UO_128 (O_128,N_13934,N_14148);
nand UO_129 (O_129,N_14018,N_14304);
xor UO_130 (O_130,N_13616,N_14526);
xor UO_131 (O_131,N_13575,N_14474);
and UO_132 (O_132,N_14576,N_14490);
or UO_133 (O_133,N_14839,N_13518);
nor UO_134 (O_134,N_14807,N_14046);
nand UO_135 (O_135,N_14045,N_14859);
nor UO_136 (O_136,N_14350,N_13646);
and UO_137 (O_137,N_14934,N_14657);
and UO_138 (O_138,N_13872,N_14552);
or UO_139 (O_139,N_14586,N_14793);
nand UO_140 (O_140,N_13943,N_14397);
or UO_141 (O_141,N_14286,N_13545);
xnor UO_142 (O_142,N_14134,N_13537);
and UO_143 (O_143,N_13859,N_14528);
or UO_144 (O_144,N_14076,N_14208);
xnor UO_145 (O_145,N_14785,N_14932);
and UO_146 (O_146,N_13845,N_13744);
nor UO_147 (O_147,N_14189,N_13693);
or UO_148 (O_148,N_14320,N_14226);
and UO_149 (O_149,N_14838,N_13559);
or UO_150 (O_150,N_13720,N_13783);
and UO_151 (O_151,N_14678,N_14339);
nor UO_152 (O_152,N_13828,N_14551);
nor UO_153 (O_153,N_14673,N_14033);
or UO_154 (O_154,N_14250,N_14390);
or UO_155 (O_155,N_14804,N_14846);
nand UO_156 (O_156,N_14459,N_14287);
xnor UO_157 (O_157,N_13548,N_14800);
and UO_158 (O_158,N_14100,N_14361);
xnor UO_159 (O_159,N_14773,N_13860);
xor UO_160 (O_160,N_14987,N_14384);
nand UO_161 (O_161,N_14888,N_13721);
or UO_162 (O_162,N_14853,N_13570);
nand UO_163 (O_163,N_14873,N_13808);
nand UO_164 (O_164,N_13949,N_13966);
or UO_165 (O_165,N_14641,N_14378);
and UO_166 (O_166,N_13956,N_14672);
xnor UO_167 (O_167,N_13546,N_13977);
or UO_168 (O_168,N_14857,N_13983);
xnor UO_169 (O_169,N_13524,N_13766);
nor UO_170 (O_170,N_13703,N_14554);
nand UO_171 (O_171,N_13611,N_14669);
nand UO_172 (O_172,N_14357,N_13675);
nor UO_173 (O_173,N_14629,N_14324);
or UO_174 (O_174,N_14689,N_13825);
and UO_175 (O_175,N_14610,N_14966);
nand UO_176 (O_176,N_13654,N_14465);
nor UO_177 (O_177,N_14967,N_13914);
nor UO_178 (O_178,N_14149,N_14187);
nand UO_179 (O_179,N_13574,N_14035);
nand UO_180 (O_180,N_14303,N_13599);
xor UO_181 (O_181,N_14094,N_13686);
nor UO_182 (O_182,N_13984,N_13925);
and UO_183 (O_183,N_14541,N_14604);
nand UO_184 (O_184,N_14057,N_14749);
nand UO_185 (O_185,N_14692,N_14892);
nor UO_186 (O_186,N_14542,N_13521);
or UO_187 (O_187,N_14970,N_14108);
xor UO_188 (O_188,N_13513,N_13839);
xnor UO_189 (O_189,N_13894,N_13591);
nor UO_190 (O_190,N_13577,N_14074);
or UO_191 (O_191,N_14575,N_14778);
or UO_192 (O_192,N_14720,N_13682);
or UO_193 (O_193,N_14137,N_14864);
or UO_194 (O_194,N_13895,N_14491);
or UO_195 (O_195,N_14068,N_14755);
xor UO_196 (O_196,N_14014,N_14174);
or UO_197 (O_197,N_14082,N_13504);
or UO_198 (O_198,N_13764,N_14159);
nand UO_199 (O_199,N_13771,N_14858);
nand UO_200 (O_200,N_13655,N_13653);
nor UO_201 (O_201,N_14922,N_13549);
xnor UO_202 (O_202,N_14469,N_14270);
nand UO_203 (O_203,N_13620,N_13916);
or UO_204 (O_204,N_14037,N_14571);
or UO_205 (O_205,N_14716,N_14964);
or UO_206 (O_206,N_13753,N_14275);
xor UO_207 (O_207,N_14292,N_13789);
nor UO_208 (O_208,N_13677,N_14322);
nor UO_209 (O_209,N_14662,N_14628);
nand UO_210 (O_210,N_14445,N_13710);
or UO_211 (O_211,N_13746,N_14737);
nand UO_212 (O_212,N_13992,N_14497);
xnor UO_213 (O_213,N_14881,N_14653);
xnor UO_214 (O_214,N_14862,N_14786);
nor UO_215 (O_215,N_14293,N_14637);
nand UO_216 (O_216,N_14239,N_14434);
xnor UO_217 (O_217,N_14209,N_14373);
and UO_218 (O_218,N_14681,N_13734);
xor UO_219 (O_219,N_14898,N_14548);
or UO_220 (O_220,N_14836,N_14199);
nand UO_221 (O_221,N_13612,N_13695);
or UO_222 (O_222,N_14252,N_14811);
and UO_223 (O_223,N_14146,N_14933);
and UO_224 (O_224,N_13728,N_13854);
xnor UO_225 (O_225,N_14241,N_13889);
or UO_226 (O_226,N_14188,N_13875);
and UO_227 (O_227,N_14823,N_14195);
xnor UO_228 (O_228,N_14860,N_14597);
nor UO_229 (O_229,N_14019,N_14487);
and UO_230 (O_230,N_14911,N_14071);
xnor UO_231 (O_231,N_14837,N_14721);
and UO_232 (O_232,N_13738,N_13660);
or UO_233 (O_233,N_14453,N_13946);
nand UO_234 (O_234,N_14524,N_14039);
xnor UO_235 (O_235,N_13566,N_14217);
or UO_236 (O_236,N_14544,N_13739);
nand UO_237 (O_237,N_13841,N_14054);
nor UO_238 (O_238,N_13532,N_14594);
nand UO_239 (O_239,N_13623,N_13523);
or UO_240 (O_240,N_14915,N_14992);
xnor UO_241 (O_241,N_14000,N_14928);
nand UO_242 (O_242,N_14299,N_14774);
nand UO_243 (O_243,N_13777,N_13852);
or UO_244 (O_244,N_14848,N_13742);
nand UO_245 (O_245,N_14639,N_14496);
and UO_246 (O_246,N_13773,N_14919);
or UO_247 (O_247,N_13668,N_14815);
or UO_248 (O_248,N_14167,N_13507);
or UO_249 (O_249,N_14602,N_13919);
xor UO_250 (O_250,N_14198,N_14482);
xor UO_251 (O_251,N_14826,N_14428);
xor UO_252 (O_252,N_14820,N_13775);
or UO_253 (O_253,N_13512,N_14003);
or UO_254 (O_254,N_14143,N_14573);
nand UO_255 (O_255,N_13818,N_14191);
or UO_256 (O_256,N_13874,N_14031);
nand UO_257 (O_257,N_13757,N_14557);
and UO_258 (O_258,N_13509,N_14917);
xnor UO_259 (O_259,N_14483,N_14395);
and UO_260 (O_260,N_14007,N_14751);
nor UO_261 (O_261,N_14321,N_13930);
or UO_262 (O_262,N_14374,N_14247);
nor UO_263 (O_263,N_14627,N_13716);
nand UO_264 (O_264,N_13691,N_14651);
xnor UO_265 (O_265,N_14608,N_14518);
and UO_266 (O_266,N_14394,N_13959);
nand UO_267 (O_267,N_14772,N_14485);
nand UO_268 (O_268,N_14438,N_14294);
or UO_269 (O_269,N_13941,N_13891);
and UO_270 (O_270,N_14723,N_14300);
xor UO_271 (O_271,N_13920,N_13661);
nor UO_272 (O_272,N_14310,N_14478);
and UO_273 (O_273,N_14440,N_13990);
nand UO_274 (O_274,N_14396,N_14668);
nor UO_275 (O_275,N_13698,N_13823);
or UO_276 (O_276,N_13560,N_14140);
nor UO_277 (O_277,N_13558,N_14372);
xor UO_278 (O_278,N_14523,N_13847);
nor UO_279 (O_279,N_14356,N_14463);
or UO_280 (O_280,N_14290,N_13610);
nor UO_281 (O_281,N_13740,N_13759);
nor UO_282 (O_282,N_13997,N_14684);
or UO_283 (O_283,N_14336,N_13981);
nor UO_284 (O_284,N_14200,N_14093);
or UO_285 (O_285,N_14297,N_14978);
xor UO_286 (O_286,N_13706,N_14998);
or UO_287 (O_287,N_14441,N_14719);
or UO_288 (O_288,N_14842,N_13760);
nor UO_289 (O_289,N_14333,N_14802);
or UO_290 (O_290,N_13628,N_14165);
xor UO_291 (O_291,N_14214,N_14784);
or UO_292 (O_292,N_14447,N_14343);
and UO_293 (O_293,N_14574,N_13602);
or UO_294 (O_294,N_13731,N_14952);
or UO_295 (O_295,N_14313,N_14914);
nand UO_296 (O_296,N_14201,N_13882);
nand UO_297 (O_297,N_14543,N_14017);
nand UO_298 (O_298,N_14462,N_14540);
nor UO_299 (O_299,N_14470,N_14312);
nand UO_300 (O_300,N_13754,N_14989);
and UO_301 (O_301,N_13785,N_13584);
nor UO_302 (O_302,N_14644,N_14798);
or UO_303 (O_303,N_14612,N_13717);
xnor UO_304 (O_304,N_14949,N_14702);
xnor UO_305 (O_305,N_13787,N_14975);
nand UO_306 (O_306,N_14566,N_13527);
and UO_307 (O_307,N_13643,N_14262);
xnor UO_308 (O_308,N_14583,N_14944);
nor UO_309 (O_309,N_14647,N_14666);
nand UO_310 (O_310,N_13926,N_14166);
or UO_311 (O_311,N_14358,N_14097);
or UO_312 (O_312,N_14732,N_13702);
or UO_313 (O_313,N_14747,N_14130);
or UO_314 (O_314,N_14155,N_13793);
and UO_315 (O_315,N_14289,N_14081);
and UO_316 (O_316,N_14302,N_13603);
xnor UO_317 (O_317,N_14461,N_14516);
and UO_318 (O_318,N_13582,N_14005);
xor UO_319 (O_319,N_13535,N_13763);
xnor UO_320 (O_320,N_14640,N_13741);
nand UO_321 (O_321,N_14595,N_13667);
and UO_322 (O_322,N_14379,N_14150);
or UO_323 (O_323,N_14101,N_14267);
nand UO_324 (O_324,N_13857,N_14585);
and UO_325 (O_325,N_14670,N_13873);
and UO_326 (O_326,N_13902,N_14430);
nand UO_327 (O_327,N_14769,N_13804);
or UO_328 (O_328,N_13712,N_14935);
nand UO_329 (O_329,N_14841,N_14912);
nand UO_330 (O_330,N_14349,N_13962);
and UO_331 (O_331,N_14550,N_13665);
or UO_332 (O_332,N_14115,N_14560);
nand UO_333 (O_333,N_14517,N_14207);
or UO_334 (O_334,N_14218,N_13672);
and UO_335 (O_335,N_13768,N_13851);
nor UO_336 (O_336,N_14193,N_14569);
or UO_337 (O_337,N_14762,N_14277);
nand UO_338 (O_338,N_14553,N_14809);
nand UO_339 (O_339,N_14733,N_14360);
xnor UO_340 (O_340,N_13540,N_13938);
or UO_341 (O_341,N_14204,N_14136);
nor UO_342 (O_342,N_14829,N_14479);
and UO_343 (O_343,N_13564,N_14828);
and UO_344 (O_344,N_13924,N_13606);
or UO_345 (O_345,N_13645,N_14326);
nand UO_346 (O_346,N_14163,N_14391);
xnor UO_347 (O_347,N_13639,N_14026);
xnor UO_348 (O_348,N_14142,N_13724);
xnor UO_349 (O_349,N_14488,N_14761);
nor UO_350 (O_350,N_14891,N_13678);
xnor UO_351 (O_351,N_14527,N_14260);
xor UO_352 (O_352,N_14703,N_14851);
nor UO_353 (O_353,N_13939,N_14685);
or UO_354 (O_354,N_13516,N_14183);
nand UO_355 (O_355,N_14559,N_14890);
and UO_356 (O_356,N_13862,N_14770);
or UO_357 (O_357,N_14997,N_14246);
xnor UO_358 (O_358,N_13652,N_14797);
xor UO_359 (O_359,N_14563,N_14718);
xor UO_360 (O_360,N_14887,N_13811);
and UO_361 (O_361,N_14472,N_14776);
xnor UO_362 (O_362,N_14810,N_13779);
and UO_363 (O_363,N_14814,N_14759);
or UO_364 (O_364,N_13713,N_14235);
or UO_365 (O_365,N_14607,N_14213);
nand UO_366 (O_366,N_14105,N_14319);
nor UO_367 (O_367,N_14969,N_14182);
or UO_368 (O_368,N_13978,N_14877);
nand UO_369 (O_369,N_14443,N_14314);
nor UO_370 (O_370,N_14415,N_14904);
nand UO_371 (O_371,N_14139,N_14258);
and UO_372 (O_372,N_14661,N_13844);
and UO_373 (O_373,N_14171,N_14631);
and UO_374 (O_374,N_13865,N_13501);
xnor UO_375 (O_375,N_14708,N_14796);
nand UO_376 (O_376,N_14771,N_14245);
or UO_377 (O_377,N_14352,N_14305);
or UO_378 (O_378,N_14288,N_14486);
xnor UO_379 (O_379,N_13631,N_13993);
xnor UO_380 (O_380,N_14399,N_14002);
or UO_381 (O_381,N_14538,N_13615);
and UO_382 (O_382,N_14176,N_14127);
and UO_383 (O_383,N_14125,N_14084);
and UO_384 (O_384,N_13506,N_13832);
nor UO_385 (O_385,N_14418,N_14618);
nand UO_386 (O_386,N_14642,N_13748);
nand UO_387 (O_387,N_14114,N_14029);
nand UO_388 (O_388,N_13630,N_14499);
xnor UO_389 (O_389,N_14577,N_14663);
nand UO_390 (O_390,N_13684,N_14974);
nand UO_391 (O_391,N_14164,N_14151);
nor UO_392 (O_392,N_14269,N_14401);
xnor UO_393 (O_393,N_13657,N_14092);
and UO_394 (O_394,N_14073,N_13913);
and UO_395 (O_395,N_13621,N_14098);
nor UO_396 (O_396,N_14249,N_13826);
and UO_397 (O_397,N_14298,N_13508);
or UO_398 (O_398,N_14170,N_14008);
nand UO_399 (O_399,N_13725,N_14050);
nand UO_400 (O_400,N_13593,N_14446);
xor UO_401 (O_401,N_13982,N_13705);
and UO_402 (O_402,N_14177,N_13557);
and UO_403 (O_403,N_14083,N_14753);
xor UO_404 (O_404,N_14493,N_14120);
xnor UO_405 (O_405,N_14942,N_13944);
nand UO_406 (O_406,N_14417,N_13975);
xor UO_407 (O_407,N_13869,N_13980);
or UO_408 (O_408,N_13538,N_14568);
or UO_409 (O_409,N_14504,N_14530);
and UO_410 (O_410,N_14318,N_14714);
xor UO_411 (O_411,N_13907,N_14927);
nor UO_412 (O_412,N_13502,N_14044);
xnor UO_413 (O_413,N_14567,N_13969);
or UO_414 (O_414,N_14308,N_14184);
nand UO_415 (O_415,N_14248,N_14449);
or UO_416 (O_416,N_14377,N_14808);
xor UO_417 (O_417,N_14365,N_14141);
and UO_418 (O_418,N_14874,N_14724);
and UO_419 (O_419,N_13567,N_13814);
and UO_420 (O_420,N_14070,N_13974);
or UO_421 (O_421,N_13688,N_14087);
and UO_422 (O_422,N_14909,N_14128);
nor UO_423 (O_423,N_14660,N_14799);
or UO_424 (O_424,N_14329,N_13842);
and UO_425 (O_425,N_14707,N_13968);
nor UO_426 (O_426,N_14734,N_14580);
nand UO_427 (O_427,N_13529,N_14147);
nand UO_428 (O_428,N_14687,N_14278);
nor UO_429 (O_429,N_14634,N_14727);
or UO_430 (O_430,N_14856,N_14402);
nand UO_431 (O_431,N_14960,N_14240);
or UO_432 (O_432,N_13780,N_14272);
nand UO_433 (O_433,N_14203,N_13572);
nor UO_434 (O_434,N_13942,N_13701);
or UO_435 (O_435,N_14866,N_14950);
nand UO_436 (O_436,N_13680,N_14896);
and UO_437 (O_437,N_14202,N_14648);
nor UO_438 (O_438,N_14697,N_14869);
and UO_439 (O_439,N_14362,N_13528);
xor UO_440 (O_440,N_13915,N_14015);
nand UO_441 (O_441,N_14959,N_13632);
xor UO_442 (O_442,N_13531,N_14745);
nand UO_443 (O_443,N_14620,N_13629);
and UO_444 (O_444,N_14133,N_13520);
and UO_445 (O_445,N_14789,N_13662);
or UO_446 (O_446,N_13622,N_13707);
nand UO_447 (O_447,N_14581,N_14509);
or UO_448 (O_448,N_13649,N_13554);
nand UO_449 (O_449,N_13752,N_13952);
and UO_450 (O_450,N_14152,N_14587);
or UO_451 (O_451,N_14765,N_14344);
and UO_452 (O_452,N_14536,N_14348);
nand UO_453 (O_453,N_14368,N_14407);
and UO_454 (O_454,N_14220,N_13835);
xnor UO_455 (O_455,N_14178,N_13817);
or UO_456 (O_456,N_14062,N_14060);
and UO_457 (O_457,N_14983,N_14937);
nor UO_458 (O_458,N_14398,N_14388);
or UO_459 (O_459,N_14600,N_14489);
or UO_460 (O_460,N_13563,N_14939);
nor UO_461 (O_461,N_14354,N_14480);
nor UO_462 (O_462,N_14834,N_13988);
or UO_463 (O_463,N_14041,N_14514);
nand UO_464 (O_464,N_13838,N_14117);
xnor UO_465 (O_465,N_13824,N_13834);
nand UO_466 (O_466,N_14234,N_14865);
or UO_467 (O_467,N_14617,N_14840);
nand UO_468 (O_468,N_14977,N_14157);
xor UO_469 (O_469,N_14251,N_13957);
nor UO_470 (O_470,N_14091,N_13899);
xnor UO_471 (O_471,N_14831,N_14730);
or UO_472 (O_472,N_14936,N_13539);
and UO_473 (O_473,N_14955,N_14746);
or UO_474 (O_474,N_14075,N_13870);
nor UO_475 (O_475,N_13666,N_13595);
and UO_476 (O_476,N_13737,N_13625);
xnor UO_477 (O_477,N_14729,N_14682);
or UO_478 (O_478,N_14351,N_13994);
and UO_479 (O_479,N_14210,N_13905);
xnor UO_480 (O_480,N_14706,N_13890);
or UO_481 (O_481,N_13751,N_14832);
or UO_482 (O_482,N_14833,N_14345);
nand UO_483 (O_483,N_14281,N_14847);
nand UO_484 (O_484,N_14513,N_14389);
nor UO_485 (O_485,N_14013,N_14589);
or UO_486 (O_486,N_13929,N_13976);
or UO_487 (O_487,N_13690,N_14923);
nor UO_488 (O_488,N_14456,N_14725);
or UO_489 (O_489,N_13644,N_14710);
nand UO_490 (O_490,N_14671,N_14036);
and UO_491 (O_491,N_13864,N_13792);
and UO_492 (O_492,N_13735,N_13515);
or UO_493 (O_493,N_13700,N_13960);
xnor UO_494 (O_494,N_13822,N_14422);
nor UO_495 (O_495,N_14156,N_14883);
nand UO_496 (O_496,N_14122,N_14346);
or UO_497 (O_497,N_14963,N_14940);
or UO_498 (O_498,N_14750,N_13536);
nand UO_499 (O_499,N_14233,N_14049);
and UO_500 (O_500,N_13576,N_14863);
and UO_501 (O_501,N_14630,N_14367);
and UO_502 (O_502,N_13776,N_14254);
nor UO_503 (O_503,N_13588,N_13945);
and UO_504 (O_504,N_14231,N_14973);
or UO_505 (O_505,N_14709,N_14505);
nor UO_506 (O_506,N_14613,N_14306);
xor UO_507 (O_507,N_13565,N_14340);
xnor UO_508 (O_508,N_13840,N_14616);
and UO_509 (O_509,N_14768,N_14592);
nor UO_510 (O_510,N_14902,N_14713);
xnor UO_511 (O_511,N_14255,N_14145);
and UO_512 (O_512,N_14403,N_13937);
nor UO_513 (O_513,N_14104,N_13782);
nand UO_514 (O_514,N_14918,N_14212);
nor UO_515 (O_515,N_14416,N_13517);
nor UO_516 (O_516,N_14868,N_13658);
nor UO_517 (O_517,N_13750,N_14331);
nand UO_518 (O_518,N_13723,N_13633);
nand UO_519 (O_519,N_14095,N_13881);
or UO_520 (O_520,N_14066,N_14609);
and UO_521 (O_521,N_13906,N_14072);
or UO_522 (O_522,N_13568,N_13747);
nor UO_523 (O_523,N_14123,N_13692);
and UO_524 (O_524,N_14897,N_14291);
or UO_525 (O_525,N_14244,N_14454);
nand UO_526 (O_526,N_14363,N_13542);
nor UO_527 (O_527,N_14501,N_13709);
nor UO_528 (O_528,N_14579,N_14024);
xnor UO_529 (O_529,N_14481,N_14926);
xnor UO_530 (O_530,N_14787,N_14817);
or UO_531 (O_531,N_14546,N_13998);
and UO_532 (O_532,N_14426,N_14822);
and UO_533 (O_533,N_13800,N_14711);
nor UO_534 (O_534,N_14225,N_13878);
xnor UO_535 (O_535,N_14473,N_13656);
nand UO_536 (O_536,N_14435,N_13697);
xnor UO_537 (O_537,N_14271,N_14827);
xnor UO_538 (O_538,N_13587,N_14206);
or UO_539 (O_539,N_14775,N_13848);
nor UO_540 (O_540,N_14656,N_14717);
and UO_541 (O_541,N_14295,N_13714);
or UO_542 (O_542,N_13635,N_14194);
nor UO_543 (O_543,N_14633,N_14930);
and UO_544 (O_544,N_14901,N_14924);
nor UO_545 (O_545,N_13965,N_14845);
and UO_546 (O_546,N_14954,N_14301);
xnor UO_547 (O_547,N_13556,N_13940);
nor UO_548 (O_548,N_14460,N_13580);
and UO_549 (O_549,N_13928,N_14124);
or UO_550 (O_550,N_13600,N_13583);
nand UO_551 (O_551,N_14406,N_13812);
or UO_552 (O_552,N_14061,N_13669);
nand UO_553 (O_553,N_14910,N_13745);
or UO_554 (O_554,N_14089,N_14819);
or UO_555 (O_555,N_13995,N_13932);
nand UO_556 (O_556,N_14004,N_14181);
xor UO_557 (O_557,N_14468,N_14257);
xor UO_558 (O_558,N_13585,N_13730);
xor UO_559 (O_559,N_14614,N_13592);
or UO_560 (O_560,N_13954,N_13708);
and UO_561 (O_561,N_13972,N_13729);
xnor UO_562 (O_562,N_13624,N_14861);
xor UO_563 (O_563,N_14705,N_13634);
and UO_564 (O_564,N_14126,N_14712);
or UO_565 (O_565,N_14701,N_14228);
nand UO_566 (O_566,N_13788,N_14695);
xnor UO_567 (O_567,N_14376,N_14263);
and UO_568 (O_568,N_14216,N_13831);
nand UO_569 (O_569,N_14921,N_14129);
nand UO_570 (O_570,N_14879,N_14561);
nand UO_571 (O_571,N_14369,N_14047);
nand UO_572 (O_572,N_13815,N_14016);
nand UO_573 (O_573,N_14196,N_13986);
and UO_574 (O_574,N_13696,N_14754);
nor UO_575 (O_575,N_14965,N_14596);
or UO_576 (O_576,N_13903,N_14520);
nand UO_577 (O_577,N_14985,N_14215);
xnor UO_578 (O_578,N_13505,N_14079);
nand UO_579 (O_579,N_14259,N_14276);
nor UO_580 (O_580,N_13749,N_14979);
xnor UO_581 (O_581,N_14562,N_13885);
nor UO_582 (O_582,N_14205,N_14386);
and UO_583 (O_583,N_13590,N_14941);
nand UO_584 (O_584,N_14450,N_13863);
and UO_585 (O_585,N_13991,N_13586);
or UO_586 (O_586,N_13522,N_14878);
nor UO_587 (O_587,N_13770,N_14715);
xnor UO_588 (O_588,N_14452,N_14268);
nor UO_589 (O_589,N_14605,N_14690);
and UO_590 (O_590,N_14058,N_13816);
xor UO_591 (O_591,N_14332,N_13970);
and UO_592 (O_592,N_14742,N_13642);
or UO_593 (O_593,N_14330,N_13550);
and UO_594 (O_594,N_14494,N_14844);
xnor UO_595 (O_595,N_14951,N_14190);
nor UO_596 (O_596,N_14821,N_13936);
or UO_597 (O_597,N_13922,N_14704);
and UO_598 (O_598,N_14649,N_14021);
and UO_599 (O_599,N_14650,N_14652);
or UO_600 (O_600,N_13901,N_13821);
nor UO_601 (O_601,N_13963,N_14976);
nand UO_602 (O_602,N_13503,N_14048);
and UO_603 (O_603,N_14236,N_14875);
nor UO_604 (O_604,N_14224,N_14598);
or UO_605 (O_605,N_13511,N_14006);
xnor UO_606 (O_606,N_13837,N_13853);
nor UO_607 (O_607,N_14679,N_14342);
and UO_608 (O_608,N_14371,N_14572);
and UO_609 (O_609,N_13561,N_13694);
xor UO_610 (O_610,N_14619,N_14783);
xnor UO_611 (O_611,N_13781,N_14835);
nor UO_612 (O_612,N_13769,N_14971);
and UO_613 (O_613,N_13961,N_14889);
or UO_614 (O_614,N_13846,N_14028);
or UO_615 (O_615,N_14090,N_14192);
nor UO_616 (O_616,N_13699,N_14366);
or UO_617 (O_617,N_14400,N_13555);
or UO_618 (O_618,N_13964,N_14813);
and UO_619 (O_619,N_13953,N_14410);
nor UO_620 (O_620,N_14956,N_14466);
nor UO_621 (O_621,N_13617,N_14584);
nand UO_622 (O_622,N_14843,N_14872);
nand UO_623 (O_623,N_14606,N_14056);
xnor UO_624 (O_624,N_14383,N_14788);
xor UO_625 (O_625,N_13778,N_14728);
or UO_626 (O_626,N_13951,N_13727);
and UO_627 (O_627,N_13722,N_14168);
xor UO_628 (O_628,N_14077,N_14777);
nor UO_629 (O_629,N_14582,N_14103);
nand UO_630 (O_630,N_13973,N_13795);
or UO_631 (O_631,N_14119,N_14099);
nor UO_632 (O_632,N_14993,N_14011);
or UO_633 (O_633,N_14370,N_14534);
nand UO_634 (O_634,N_13909,N_14694);
nand UO_635 (O_635,N_13500,N_14116);
nand UO_636 (O_636,N_14211,N_14655);
nor UO_637 (O_637,N_14779,N_13604);
xnor UO_638 (O_638,N_14419,N_13871);
nor UO_639 (O_639,N_13772,N_14337);
or UO_640 (O_640,N_14307,N_14222);
xor UO_641 (O_641,N_14726,N_13514);
and UO_642 (O_642,N_13843,N_14507);
nor UO_643 (O_643,N_14109,N_14825);
nor UO_644 (O_644,N_13627,N_14477);
or UO_645 (O_645,N_13647,N_13637);
nand UO_646 (O_646,N_13880,N_14529);
nand UO_647 (O_647,N_13685,N_14699);
nor UO_648 (O_648,N_14578,N_14425);
nand UO_649 (O_649,N_14736,N_14691);
xor UO_650 (O_650,N_14025,N_13689);
nand UO_651 (O_651,N_14676,N_14484);
and UO_652 (O_652,N_13601,N_14698);
and UO_653 (O_653,N_14439,N_14132);
and UO_654 (O_654,N_13598,N_14722);
or UO_655 (O_655,N_14744,N_14197);
xor UO_656 (O_656,N_14953,N_14638);
nand UO_657 (O_657,N_14512,N_14020);
nor UO_658 (O_658,N_14899,N_14884);
nand UO_659 (O_659,N_14854,N_14908);
nor UO_660 (O_660,N_13979,N_14442);
nor UO_661 (O_661,N_13833,N_14547);
and UO_662 (O_662,N_13755,N_14055);
nor UO_663 (O_663,N_14818,N_13797);
or UO_664 (O_664,N_13597,N_13674);
or UO_665 (O_665,N_14920,N_13829);
and UO_666 (O_666,N_14421,N_13947);
and UO_667 (O_667,N_14355,N_14412);
nand UO_668 (O_668,N_14393,N_14409);
and UO_669 (O_669,N_14981,N_14237);
nand UO_670 (O_670,N_14266,N_13867);
and UO_671 (O_671,N_13887,N_14931);
and UO_672 (O_672,N_13774,N_14535);
and UO_673 (O_673,N_14549,N_14309);
nand UO_674 (O_674,N_14392,N_13619);
and UO_675 (O_675,N_13664,N_14767);
nor UO_676 (O_676,N_14780,N_14153);
or UO_677 (O_677,N_14227,N_14424);
and UO_678 (O_678,N_14043,N_14085);
or UO_679 (O_679,N_13526,N_14230);
nor UO_680 (O_680,N_14420,N_13573);
nor UO_681 (O_681,N_13900,N_14664);
or UO_682 (O_682,N_14261,N_14086);
or UO_683 (O_683,N_14700,N_14065);
xnor UO_684 (O_684,N_13543,N_14824);
or UO_685 (O_685,N_13836,N_13819);
and UO_686 (O_686,N_14080,N_14022);
xnor UO_687 (O_687,N_13923,N_13732);
xnor UO_688 (O_688,N_14948,N_13784);
nand UO_689 (O_689,N_14405,N_14273);
or UO_690 (O_690,N_13883,N_14903);
nor UO_691 (O_691,N_14957,N_13948);
or UO_692 (O_692,N_13626,N_13820);
and UO_693 (O_693,N_13736,N_14455);
nor UO_694 (O_694,N_13798,N_14476);
or UO_695 (O_695,N_14688,N_14667);
xnor UO_696 (O_696,N_14078,N_13879);
and UO_697 (O_697,N_14315,N_14615);
xor UO_698 (O_698,N_13917,N_14849);
or UO_699 (O_699,N_14243,N_14131);
nor UO_700 (O_700,N_14102,N_13547);
nor UO_701 (O_701,N_13912,N_14988);
or UO_702 (O_702,N_13861,N_14748);
or UO_703 (O_703,N_14038,N_14475);
nand UO_704 (O_704,N_13659,N_14012);
or UO_705 (O_705,N_14735,N_14757);
xor UO_706 (O_706,N_13607,N_14601);
xnor UO_707 (O_707,N_13849,N_14052);
nand UO_708 (O_708,N_13594,N_13687);
nand UO_709 (O_709,N_14558,N_13681);
nand UO_710 (O_710,N_14280,N_14946);
and UO_711 (O_711,N_14375,N_14886);
nand UO_712 (O_712,N_13958,N_13679);
and UO_713 (O_713,N_13806,N_14327);
nor UO_714 (O_714,N_13683,N_14962);
and UO_715 (O_715,N_14328,N_14135);
nor UO_716 (O_716,N_13955,N_13898);
nand UO_717 (O_717,N_14457,N_14686);
nand UO_718 (O_718,N_14118,N_14880);
or UO_719 (O_719,N_13803,N_14175);
xor UO_720 (O_720,N_13985,N_14624);
nor UO_721 (O_721,N_13790,N_14533);
nand UO_722 (O_722,N_14173,N_13911);
nand UO_723 (O_723,N_14264,N_13640);
and UO_724 (O_724,N_14223,N_13877);
nor UO_725 (O_725,N_13589,N_14805);
or UO_726 (O_726,N_14995,N_14325);
or UO_727 (O_727,N_14067,N_13921);
nor UO_728 (O_728,N_13876,N_14381);
nor UO_729 (O_729,N_14621,N_14740);
nand UO_730 (O_730,N_14317,N_13971);
nand UO_731 (O_731,N_14121,N_14565);
and UO_732 (O_732,N_14451,N_13650);
and UO_733 (O_733,N_14795,N_14511);
xnor UO_734 (O_734,N_14510,N_14626);
or UO_735 (O_735,N_13743,N_13794);
and UO_736 (O_736,N_13510,N_14265);
nor UO_737 (O_737,N_14111,N_14427);
and UO_738 (O_738,N_14508,N_13613);
and UO_739 (O_739,N_13718,N_14180);
nand UO_740 (O_740,N_13931,N_14738);
and UO_741 (O_741,N_13614,N_13608);
nand UO_742 (O_742,N_14106,N_14112);
and UO_743 (O_743,N_14961,N_14603);
nand UO_744 (O_744,N_14996,N_13553);
or UO_745 (O_745,N_14232,N_14158);
nor UO_746 (O_746,N_13525,N_13756);
xnor UO_747 (O_747,N_13809,N_14341);
xor UO_748 (O_748,N_14752,N_14693);
nand UO_749 (O_749,N_14088,N_14498);
or UO_750 (O_750,N_14360,N_14306);
and UO_751 (O_751,N_14990,N_13834);
xnor UO_752 (O_752,N_14875,N_13969);
and UO_753 (O_753,N_14732,N_14460);
nor UO_754 (O_754,N_13691,N_14065);
and UO_755 (O_755,N_14492,N_13943);
xor UO_756 (O_756,N_13733,N_14608);
or UO_757 (O_757,N_14263,N_14374);
and UO_758 (O_758,N_14609,N_14606);
xor UO_759 (O_759,N_13731,N_13982);
and UO_760 (O_760,N_13826,N_14190);
nor UO_761 (O_761,N_14932,N_13503);
and UO_762 (O_762,N_14565,N_14205);
or UO_763 (O_763,N_13933,N_14471);
or UO_764 (O_764,N_14093,N_14629);
and UO_765 (O_765,N_14007,N_14699);
xor UO_766 (O_766,N_14517,N_14587);
nor UO_767 (O_767,N_14142,N_13895);
nor UO_768 (O_768,N_14027,N_14290);
and UO_769 (O_769,N_14088,N_14589);
or UO_770 (O_770,N_14251,N_14917);
xor UO_771 (O_771,N_14772,N_14406);
nor UO_772 (O_772,N_14184,N_13726);
nor UO_773 (O_773,N_13834,N_14921);
xor UO_774 (O_774,N_14880,N_14360);
nor UO_775 (O_775,N_13804,N_14399);
nand UO_776 (O_776,N_14312,N_14051);
or UO_777 (O_777,N_14789,N_14489);
nor UO_778 (O_778,N_13732,N_13984);
nor UO_779 (O_779,N_14052,N_14638);
nor UO_780 (O_780,N_13777,N_14362);
nor UO_781 (O_781,N_14783,N_13936);
or UO_782 (O_782,N_13865,N_14004);
or UO_783 (O_783,N_14402,N_14861);
and UO_784 (O_784,N_13921,N_13627);
xor UO_785 (O_785,N_13943,N_14165);
nor UO_786 (O_786,N_13821,N_13985);
and UO_787 (O_787,N_14341,N_14946);
nand UO_788 (O_788,N_13658,N_13660);
and UO_789 (O_789,N_14420,N_14324);
or UO_790 (O_790,N_14093,N_14141);
nand UO_791 (O_791,N_14443,N_14129);
and UO_792 (O_792,N_14704,N_14982);
nor UO_793 (O_793,N_14526,N_14549);
xor UO_794 (O_794,N_14966,N_14457);
nor UO_795 (O_795,N_14922,N_13761);
xor UO_796 (O_796,N_14202,N_14634);
and UO_797 (O_797,N_14525,N_13647);
and UO_798 (O_798,N_14991,N_13611);
xnor UO_799 (O_799,N_14076,N_13967);
nor UO_800 (O_800,N_14185,N_14580);
or UO_801 (O_801,N_14952,N_14583);
and UO_802 (O_802,N_13799,N_14728);
nand UO_803 (O_803,N_14670,N_13572);
or UO_804 (O_804,N_13812,N_13729);
nor UO_805 (O_805,N_14170,N_14057);
and UO_806 (O_806,N_14266,N_14872);
and UO_807 (O_807,N_13927,N_14696);
nor UO_808 (O_808,N_14935,N_14580);
xnor UO_809 (O_809,N_14400,N_13500);
and UO_810 (O_810,N_14515,N_14418);
nor UO_811 (O_811,N_14049,N_14737);
and UO_812 (O_812,N_14393,N_14069);
nor UO_813 (O_813,N_14854,N_13645);
nand UO_814 (O_814,N_14813,N_14640);
nand UO_815 (O_815,N_14921,N_14723);
nor UO_816 (O_816,N_13897,N_14851);
nor UO_817 (O_817,N_14182,N_13945);
nor UO_818 (O_818,N_14161,N_13654);
nand UO_819 (O_819,N_14569,N_14404);
nor UO_820 (O_820,N_14471,N_14486);
and UO_821 (O_821,N_13946,N_14838);
or UO_822 (O_822,N_14525,N_14683);
and UO_823 (O_823,N_14777,N_13725);
xor UO_824 (O_824,N_13645,N_14307);
nand UO_825 (O_825,N_14336,N_14355);
or UO_826 (O_826,N_14456,N_14838);
nand UO_827 (O_827,N_14731,N_13578);
nor UO_828 (O_828,N_14219,N_14811);
nand UO_829 (O_829,N_14754,N_14852);
xnor UO_830 (O_830,N_14552,N_13913);
or UO_831 (O_831,N_14555,N_14288);
nand UO_832 (O_832,N_14700,N_13532);
and UO_833 (O_833,N_14340,N_14678);
xnor UO_834 (O_834,N_14442,N_13830);
nor UO_835 (O_835,N_14038,N_14824);
and UO_836 (O_836,N_14693,N_13624);
nor UO_837 (O_837,N_14243,N_13755);
xnor UO_838 (O_838,N_13641,N_13726);
and UO_839 (O_839,N_14561,N_14478);
and UO_840 (O_840,N_14364,N_14798);
and UO_841 (O_841,N_14834,N_14197);
nor UO_842 (O_842,N_14180,N_14248);
nand UO_843 (O_843,N_13881,N_14882);
or UO_844 (O_844,N_14168,N_14104);
or UO_845 (O_845,N_14415,N_13919);
and UO_846 (O_846,N_14153,N_14609);
or UO_847 (O_847,N_13511,N_14842);
xor UO_848 (O_848,N_14041,N_13931);
xnor UO_849 (O_849,N_14253,N_14385);
nand UO_850 (O_850,N_14445,N_13708);
xor UO_851 (O_851,N_14062,N_14253);
nand UO_852 (O_852,N_14958,N_14485);
nand UO_853 (O_853,N_14011,N_14489);
and UO_854 (O_854,N_14902,N_14393);
nor UO_855 (O_855,N_13514,N_14297);
and UO_856 (O_856,N_14589,N_14889);
xor UO_857 (O_857,N_14495,N_13787);
xor UO_858 (O_858,N_14731,N_14189);
xor UO_859 (O_859,N_14823,N_13976);
nand UO_860 (O_860,N_13991,N_14938);
nand UO_861 (O_861,N_14928,N_14750);
nand UO_862 (O_862,N_14305,N_14898);
nand UO_863 (O_863,N_13568,N_14588);
and UO_864 (O_864,N_14508,N_14027);
and UO_865 (O_865,N_14296,N_14942);
nor UO_866 (O_866,N_13967,N_13534);
xnor UO_867 (O_867,N_14940,N_13511);
xnor UO_868 (O_868,N_14216,N_13679);
nor UO_869 (O_869,N_14404,N_14536);
or UO_870 (O_870,N_14570,N_13944);
nor UO_871 (O_871,N_14826,N_13796);
nand UO_872 (O_872,N_14690,N_14041);
xor UO_873 (O_873,N_13821,N_14770);
and UO_874 (O_874,N_13795,N_14411);
and UO_875 (O_875,N_14347,N_14126);
or UO_876 (O_876,N_14861,N_14108);
or UO_877 (O_877,N_14749,N_14445);
nand UO_878 (O_878,N_14452,N_14220);
xor UO_879 (O_879,N_14932,N_13883);
and UO_880 (O_880,N_14617,N_14349);
xor UO_881 (O_881,N_13741,N_14860);
nand UO_882 (O_882,N_14491,N_14765);
nor UO_883 (O_883,N_14201,N_14922);
nand UO_884 (O_884,N_14729,N_14044);
and UO_885 (O_885,N_14384,N_14260);
nand UO_886 (O_886,N_14842,N_13840);
nand UO_887 (O_887,N_14331,N_13653);
and UO_888 (O_888,N_14665,N_13888);
or UO_889 (O_889,N_14006,N_14090);
nand UO_890 (O_890,N_14277,N_13743);
or UO_891 (O_891,N_13636,N_14989);
xnor UO_892 (O_892,N_13610,N_13604);
and UO_893 (O_893,N_13815,N_13727);
xor UO_894 (O_894,N_14758,N_14966);
nand UO_895 (O_895,N_14515,N_14677);
or UO_896 (O_896,N_13853,N_14517);
nand UO_897 (O_897,N_13510,N_14515);
nand UO_898 (O_898,N_14219,N_14236);
xnor UO_899 (O_899,N_13899,N_14977);
or UO_900 (O_900,N_14043,N_14597);
and UO_901 (O_901,N_14523,N_14344);
nand UO_902 (O_902,N_14509,N_13708);
xnor UO_903 (O_903,N_14677,N_14089);
xnor UO_904 (O_904,N_14864,N_14075);
nor UO_905 (O_905,N_14694,N_13598);
nand UO_906 (O_906,N_13606,N_13857);
and UO_907 (O_907,N_14911,N_13809);
nand UO_908 (O_908,N_14030,N_14428);
or UO_909 (O_909,N_14521,N_14986);
nand UO_910 (O_910,N_14431,N_14467);
and UO_911 (O_911,N_14582,N_13504);
nor UO_912 (O_912,N_14438,N_13560);
or UO_913 (O_913,N_14897,N_14597);
xor UO_914 (O_914,N_13708,N_14249);
xnor UO_915 (O_915,N_14403,N_14117);
xnor UO_916 (O_916,N_14700,N_14448);
nor UO_917 (O_917,N_13577,N_13877);
nor UO_918 (O_918,N_14033,N_13549);
nor UO_919 (O_919,N_13543,N_14635);
xor UO_920 (O_920,N_13777,N_14497);
xnor UO_921 (O_921,N_14990,N_13786);
or UO_922 (O_922,N_14628,N_13941);
or UO_923 (O_923,N_13558,N_14063);
nor UO_924 (O_924,N_14887,N_14175);
nor UO_925 (O_925,N_13584,N_13963);
or UO_926 (O_926,N_14240,N_14440);
nor UO_927 (O_927,N_13936,N_14300);
nor UO_928 (O_928,N_14269,N_13675);
nand UO_929 (O_929,N_13566,N_14082);
and UO_930 (O_930,N_14630,N_14110);
nor UO_931 (O_931,N_13871,N_14193);
nor UO_932 (O_932,N_14609,N_14993);
nor UO_933 (O_933,N_14936,N_14527);
nor UO_934 (O_934,N_14881,N_13768);
xnor UO_935 (O_935,N_14353,N_14908);
or UO_936 (O_936,N_14312,N_14377);
or UO_937 (O_937,N_13760,N_14350);
nor UO_938 (O_938,N_13674,N_13917);
xor UO_939 (O_939,N_13591,N_13719);
nor UO_940 (O_940,N_14233,N_13797);
nand UO_941 (O_941,N_14483,N_13554);
nand UO_942 (O_942,N_13768,N_14792);
nor UO_943 (O_943,N_13728,N_13600);
and UO_944 (O_944,N_13894,N_14732);
xor UO_945 (O_945,N_14495,N_13747);
or UO_946 (O_946,N_14558,N_13735);
xnor UO_947 (O_947,N_13743,N_14351);
or UO_948 (O_948,N_14434,N_14412);
nor UO_949 (O_949,N_14068,N_14094);
nor UO_950 (O_950,N_14291,N_14642);
and UO_951 (O_951,N_14335,N_14834);
or UO_952 (O_952,N_14183,N_14420);
nand UO_953 (O_953,N_14142,N_14747);
or UO_954 (O_954,N_14836,N_14027);
nand UO_955 (O_955,N_14751,N_13955);
and UO_956 (O_956,N_13776,N_13594);
and UO_957 (O_957,N_13822,N_14508);
nor UO_958 (O_958,N_14421,N_13704);
nand UO_959 (O_959,N_13762,N_14923);
xnor UO_960 (O_960,N_13907,N_14520);
nor UO_961 (O_961,N_14266,N_13642);
and UO_962 (O_962,N_13735,N_14168);
or UO_963 (O_963,N_14853,N_13682);
or UO_964 (O_964,N_13549,N_14817);
nor UO_965 (O_965,N_13890,N_13605);
nor UO_966 (O_966,N_14032,N_14368);
nor UO_967 (O_967,N_13886,N_14787);
and UO_968 (O_968,N_14917,N_14684);
and UO_969 (O_969,N_14837,N_14312);
nand UO_970 (O_970,N_14236,N_13597);
nand UO_971 (O_971,N_13991,N_13647);
nand UO_972 (O_972,N_14411,N_14928);
nand UO_973 (O_973,N_14065,N_14303);
nand UO_974 (O_974,N_13954,N_14238);
nand UO_975 (O_975,N_14312,N_14677);
nor UO_976 (O_976,N_14272,N_14837);
or UO_977 (O_977,N_14707,N_14199);
and UO_978 (O_978,N_13553,N_14707);
and UO_979 (O_979,N_13599,N_14696);
or UO_980 (O_980,N_14334,N_14867);
and UO_981 (O_981,N_14258,N_13539);
xor UO_982 (O_982,N_14920,N_14558);
nor UO_983 (O_983,N_14827,N_14049);
xor UO_984 (O_984,N_14459,N_14618);
nand UO_985 (O_985,N_14682,N_14912);
and UO_986 (O_986,N_14033,N_13671);
nand UO_987 (O_987,N_14189,N_14031);
nor UO_988 (O_988,N_14398,N_13960);
and UO_989 (O_989,N_13981,N_14525);
xor UO_990 (O_990,N_13810,N_14239);
and UO_991 (O_991,N_14245,N_14902);
or UO_992 (O_992,N_13501,N_13751);
nor UO_993 (O_993,N_13945,N_14777);
or UO_994 (O_994,N_14356,N_14422);
nand UO_995 (O_995,N_14327,N_14822);
nand UO_996 (O_996,N_13647,N_13612);
and UO_997 (O_997,N_13987,N_13877);
nor UO_998 (O_998,N_13516,N_14695);
and UO_999 (O_999,N_14367,N_14961);
nor UO_1000 (O_1000,N_13698,N_14965);
xor UO_1001 (O_1001,N_13556,N_13723);
or UO_1002 (O_1002,N_13948,N_13631);
and UO_1003 (O_1003,N_14549,N_14773);
xnor UO_1004 (O_1004,N_14703,N_13724);
and UO_1005 (O_1005,N_13818,N_14936);
nor UO_1006 (O_1006,N_14130,N_14128);
or UO_1007 (O_1007,N_14042,N_14275);
xor UO_1008 (O_1008,N_14964,N_14027);
or UO_1009 (O_1009,N_14076,N_14732);
or UO_1010 (O_1010,N_14272,N_14579);
xor UO_1011 (O_1011,N_13978,N_14744);
nor UO_1012 (O_1012,N_14840,N_14344);
xor UO_1013 (O_1013,N_14245,N_14750);
nor UO_1014 (O_1014,N_13939,N_14190);
nor UO_1015 (O_1015,N_14796,N_13813);
and UO_1016 (O_1016,N_14205,N_14473);
xnor UO_1017 (O_1017,N_14955,N_14049);
nor UO_1018 (O_1018,N_13980,N_13724);
and UO_1019 (O_1019,N_13692,N_13506);
nand UO_1020 (O_1020,N_13667,N_14037);
and UO_1021 (O_1021,N_14965,N_14184);
or UO_1022 (O_1022,N_13666,N_14348);
or UO_1023 (O_1023,N_14563,N_14062);
nand UO_1024 (O_1024,N_13751,N_14275);
nand UO_1025 (O_1025,N_14658,N_14588);
or UO_1026 (O_1026,N_14088,N_14186);
and UO_1027 (O_1027,N_14022,N_14409);
nor UO_1028 (O_1028,N_14294,N_14443);
xor UO_1029 (O_1029,N_13589,N_14429);
and UO_1030 (O_1030,N_14565,N_14653);
xor UO_1031 (O_1031,N_13583,N_14632);
nand UO_1032 (O_1032,N_14330,N_14470);
nor UO_1033 (O_1033,N_14624,N_14039);
nor UO_1034 (O_1034,N_13906,N_14235);
xor UO_1035 (O_1035,N_13592,N_13878);
nand UO_1036 (O_1036,N_14930,N_14259);
and UO_1037 (O_1037,N_14413,N_14945);
xor UO_1038 (O_1038,N_14390,N_14826);
xnor UO_1039 (O_1039,N_14927,N_13731);
xnor UO_1040 (O_1040,N_14024,N_14938);
and UO_1041 (O_1041,N_14687,N_13858);
or UO_1042 (O_1042,N_14059,N_14751);
or UO_1043 (O_1043,N_14493,N_14294);
xor UO_1044 (O_1044,N_14660,N_14028);
xor UO_1045 (O_1045,N_14665,N_14766);
and UO_1046 (O_1046,N_13973,N_14348);
or UO_1047 (O_1047,N_14988,N_14072);
nand UO_1048 (O_1048,N_14361,N_13811);
nor UO_1049 (O_1049,N_14246,N_14423);
nor UO_1050 (O_1050,N_13535,N_14683);
nand UO_1051 (O_1051,N_13821,N_13595);
and UO_1052 (O_1052,N_13731,N_13768);
xnor UO_1053 (O_1053,N_14967,N_13682);
xnor UO_1054 (O_1054,N_14711,N_14921);
nor UO_1055 (O_1055,N_14742,N_14128);
nor UO_1056 (O_1056,N_14617,N_14715);
nor UO_1057 (O_1057,N_13519,N_13700);
xor UO_1058 (O_1058,N_14665,N_14615);
and UO_1059 (O_1059,N_13892,N_14892);
xor UO_1060 (O_1060,N_14795,N_13985);
nor UO_1061 (O_1061,N_13909,N_14491);
nor UO_1062 (O_1062,N_13664,N_14944);
and UO_1063 (O_1063,N_14548,N_14355);
xnor UO_1064 (O_1064,N_13501,N_13511);
nor UO_1065 (O_1065,N_13888,N_13823);
nor UO_1066 (O_1066,N_14073,N_13999);
xnor UO_1067 (O_1067,N_13810,N_14439);
or UO_1068 (O_1068,N_14650,N_14448);
nand UO_1069 (O_1069,N_14203,N_14745);
and UO_1070 (O_1070,N_13723,N_14496);
nand UO_1071 (O_1071,N_13973,N_13910);
nand UO_1072 (O_1072,N_14713,N_14132);
nand UO_1073 (O_1073,N_14931,N_14175);
and UO_1074 (O_1074,N_13648,N_14942);
nand UO_1075 (O_1075,N_13539,N_13550);
or UO_1076 (O_1076,N_14865,N_14852);
nor UO_1077 (O_1077,N_14962,N_13961);
xnor UO_1078 (O_1078,N_14391,N_14506);
nand UO_1079 (O_1079,N_14554,N_14091);
nand UO_1080 (O_1080,N_14866,N_13690);
nor UO_1081 (O_1081,N_14363,N_14165);
nand UO_1082 (O_1082,N_14088,N_13673);
or UO_1083 (O_1083,N_14690,N_13779);
or UO_1084 (O_1084,N_13699,N_14323);
nor UO_1085 (O_1085,N_14756,N_13702);
xor UO_1086 (O_1086,N_13896,N_14234);
or UO_1087 (O_1087,N_13948,N_14202);
nor UO_1088 (O_1088,N_13536,N_13988);
nor UO_1089 (O_1089,N_14964,N_13644);
or UO_1090 (O_1090,N_14873,N_14128);
xor UO_1091 (O_1091,N_14844,N_13980);
and UO_1092 (O_1092,N_14296,N_14640);
nand UO_1093 (O_1093,N_14301,N_14766);
xor UO_1094 (O_1094,N_13885,N_14960);
or UO_1095 (O_1095,N_13574,N_14115);
or UO_1096 (O_1096,N_14991,N_14726);
and UO_1097 (O_1097,N_14721,N_14259);
nand UO_1098 (O_1098,N_13819,N_13625);
or UO_1099 (O_1099,N_14792,N_13790);
or UO_1100 (O_1100,N_14527,N_13801);
and UO_1101 (O_1101,N_14703,N_14165);
xor UO_1102 (O_1102,N_14303,N_14559);
nand UO_1103 (O_1103,N_14725,N_14717);
nor UO_1104 (O_1104,N_13508,N_14680);
xnor UO_1105 (O_1105,N_13991,N_14808);
nor UO_1106 (O_1106,N_14469,N_13880);
or UO_1107 (O_1107,N_14156,N_13724);
nor UO_1108 (O_1108,N_14247,N_14218);
or UO_1109 (O_1109,N_14045,N_13956);
nor UO_1110 (O_1110,N_14653,N_14295);
nor UO_1111 (O_1111,N_14031,N_14290);
nand UO_1112 (O_1112,N_14927,N_13807);
xnor UO_1113 (O_1113,N_14570,N_14140);
and UO_1114 (O_1114,N_13819,N_13974);
xnor UO_1115 (O_1115,N_14935,N_14354);
nand UO_1116 (O_1116,N_13645,N_14327);
nand UO_1117 (O_1117,N_14699,N_14198);
nand UO_1118 (O_1118,N_14154,N_14713);
and UO_1119 (O_1119,N_13540,N_13900);
nor UO_1120 (O_1120,N_14135,N_14916);
nand UO_1121 (O_1121,N_13788,N_13534);
nor UO_1122 (O_1122,N_14655,N_13613);
nand UO_1123 (O_1123,N_14158,N_13854);
nand UO_1124 (O_1124,N_14610,N_14150);
nand UO_1125 (O_1125,N_13692,N_14246);
or UO_1126 (O_1126,N_14203,N_14051);
or UO_1127 (O_1127,N_14172,N_13867);
nor UO_1128 (O_1128,N_14331,N_14876);
or UO_1129 (O_1129,N_13699,N_14318);
nor UO_1130 (O_1130,N_14590,N_14117);
nor UO_1131 (O_1131,N_13870,N_13686);
nor UO_1132 (O_1132,N_14563,N_14933);
nand UO_1133 (O_1133,N_13816,N_14247);
nand UO_1134 (O_1134,N_14109,N_13716);
and UO_1135 (O_1135,N_14732,N_14955);
xor UO_1136 (O_1136,N_13908,N_14874);
and UO_1137 (O_1137,N_14724,N_14655);
nand UO_1138 (O_1138,N_13582,N_14133);
nor UO_1139 (O_1139,N_14605,N_14578);
and UO_1140 (O_1140,N_13933,N_13920);
nor UO_1141 (O_1141,N_14915,N_14808);
or UO_1142 (O_1142,N_14006,N_14369);
or UO_1143 (O_1143,N_13541,N_14383);
or UO_1144 (O_1144,N_13602,N_14275);
and UO_1145 (O_1145,N_13565,N_14608);
or UO_1146 (O_1146,N_14779,N_14850);
nor UO_1147 (O_1147,N_14231,N_13678);
and UO_1148 (O_1148,N_13833,N_14784);
and UO_1149 (O_1149,N_14480,N_14047);
nand UO_1150 (O_1150,N_13650,N_14140);
and UO_1151 (O_1151,N_14262,N_14584);
or UO_1152 (O_1152,N_13766,N_14612);
nor UO_1153 (O_1153,N_14043,N_13674);
xnor UO_1154 (O_1154,N_14608,N_13909);
nand UO_1155 (O_1155,N_13764,N_13657);
or UO_1156 (O_1156,N_14601,N_13760);
and UO_1157 (O_1157,N_13850,N_14691);
and UO_1158 (O_1158,N_13766,N_14837);
xnor UO_1159 (O_1159,N_13595,N_14505);
nand UO_1160 (O_1160,N_14308,N_14480);
nand UO_1161 (O_1161,N_14574,N_13587);
nor UO_1162 (O_1162,N_14509,N_14978);
and UO_1163 (O_1163,N_14323,N_13716);
xnor UO_1164 (O_1164,N_14339,N_14735);
and UO_1165 (O_1165,N_14473,N_14374);
xor UO_1166 (O_1166,N_14763,N_14114);
or UO_1167 (O_1167,N_14399,N_14094);
nand UO_1168 (O_1168,N_13621,N_14536);
nor UO_1169 (O_1169,N_14737,N_14756);
and UO_1170 (O_1170,N_14801,N_14633);
nand UO_1171 (O_1171,N_13584,N_14037);
and UO_1172 (O_1172,N_13757,N_14655);
or UO_1173 (O_1173,N_14825,N_13890);
nand UO_1174 (O_1174,N_14121,N_13752);
and UO_1175 (O_1175,N_13923,N_13974);
and UO_1176 (O_1176,N_14728,N_14808);
xnor UO_1177 (O_1177,N_14214,N_14180);
xnor UO_1178 (O_1178,N_14137,N_14468);
nand UO_1179 (O_1179,N_13837,N_14455);
and UO_1180 (O_1180,N_14553,N_14799);
and UO_1181 (O_1181,N_14456,N_14242);
nor UO_1182 (O_1182,N_14726,N_13754);
nor UO_1183 (O_1183,N_13693,N_14009);
xnor UO_1184 (O_1184,N_14918,N_14898);
nor UO_1185 (O_1185,N_14891,N_14500);
or UO_1186 (O_1186,N_13718,N_13690);
nand UO_1187 (O_1187,N_14202,N_14287);
nand UO_1188 (O_1188,N_14724,N_14562);
and UO_1189 (O_1189,N_13792,N_14238);
nand UO_1190 (O_1190,N_14324,N_14182);
and UO_1191 (O_1191,N_14933,N_14931);
nand UO_1192 (O_1192,N_13692,N_14238);
nand UO_1193 (O_1193,N_14171,N_14118);
nand UO_1194 (O_1194,N_14130,N_13547);
nor UO_1195 (O_1195,N_14532,N_14925);
nand UO_1196 (O_1196,N_14686,N_14521);
nor UO_1197 (O_1197,N_14203,N_13684);
xnor UO_1198 (O_1198,N_13732,N_14510);
xnor UO_1199 (O_1199,N_13521,N_14032);
and UO_1200 (O_1200,N_13926,N_14627);
nand UO_1201 (O_1201,N_14595,N_13860);
nor UO_1202 (O_1202,N_14659,N_14553);
nand UO_1203 (O_1203,N_13720,N_13832);
xor UO_1204 (O_1204,N_14621,N_14148);
nand UO_1205 (O_1205,N_14567,N_14987);
xor UO_1206 (O_1206,N_13936,N_13872);
nor UO_1207 (O_1207,N_14335,N_14313);
nand UO_1208 (O_1208,N_14054,N_14952);
nand UO_1209 (O_1209,N_13734,N_14071);
or UO_1210 (O_1210,N_14057,N_14199);
nand UO_1211 (O_1211,N_14373,N_14477);
nand UO_1212 (O_1212,N_14739,N_13903);
and UO_1213 (O_1213,N_14164,N_14536);
nand UO_1214 (O_1214,N_14216,N_14284);
nand UO_1215 (O_1215,N_14250,N_13521);
xor UO_1216 (O_1216,N_14476,N_14629);
and UO_1217 (O_1217,N_14201,N_13519);
and UO_1218 (O_1218,N_14295,N_13902);
xnor UO_1219 (O_1219,N_13679,N_13519);
nand UO_1220 (O_1220,N_14088,N_14923);
nand UO_1221 (O_1221,N_13912,N_13636);
or UO_1222 (O_1222,N_13739,N_13644);
nand UO_1223 (O_1223,N_14555,N_14850);
xor UO_1224 (O_1224,N_13830,N_14874);
or UO_1225 (O_1225,N_14441,N_14413);
nor UO_1226 (O_1226,N_14443,N_14223);
nor UO_1227 (O_1227,N_14642,N_13962);
nand UO_1228 (O_1228,N_14218,N_13586);
nor UO_1229 (O_1229,N_14042,N_13665);
and UO_1230 (O_1230,N_14999,N_14482);
and UO_1231 (O_1231,N_13687,N_13529);
or UO_1232 (O_1232,N_14992,N_13923);
nand UO_1233 (O_1233,N_14645,N_13950);
or UO_1234 (O_1234,N_14204,N_14590);
nand UO_1235 (O_1235,N_14193,N_13541);
xnor UO_1236 (O_1236,N_13643,N_14578);
xor UO_1237 (O_1237,N_14772,N_13792);
or UO_1238 (O_1238,N_14291,N_14997);
and UO_1239 (O_1239,N_13977,N_13720);
and UO_1240 (O_1240,N_13664,N_14989);
xnor UO_1241 (O_1241,N_14446,N_14469);
nand UO_1242 (O_1242,N_13950,N_13969);
xor UO_1243 (O_1243,N_14025,N_14729);
nand UO_1244 (O_1244,N_13845,N_14447);
nor UO_1245 (O_1245,N_13992,N_13586);
or UO_1246 (O_1246,N_14142,N_14924);
or UO_1247 (O_1247,N_14991,N_13687);
nor UO_1248 (O_1248,N_14169,N_14768);
nand UO_1249 (O_1249,N_14843,N_14521);
nor UO_1250 (O_1250,N_13973,N_13803);
or UO_1251 (O_1251,N_14729,N_14698);
or UO_1252 (O_1252,N_14457,N_13534);
or UO_1253 (O_1253,N_14577,N_14902);
and UO_1254 (O_1254,N_14042,N_13806);
or UO_1255 (O_1255,N_14965,N_13711);
and UO_1256 (O_1256,N_13855,N_13800);
xnor UO_1257 (O_1257,N_14885,N_14694);
xnor UO_1258 (O_1258,N_14495,N_13602);
or UO_1259 (O_1259,N_14600,N_13741);
or UO_1260 (O_1260,N_13633,N_14906);
xnor UO_1261 (O_1261,N_14535,N_13543);
xor UO_1262 (O_1262,N_14424,N_14544);
and UO_1263 (O_1263,N_14630,N_13968);
nor UO_1264 (O_1264,N_14130,N_13708);
or UO_1265 (O_1265,N_13822,N_14917);
nor UO_1266 (O_1266,N_13830,N_14474);
nor UO_1267 (O_1267,N_14854,N_13734);
nand UO_1268 (O_1268,N_13785,N_14972);
or UO_1269 (O_1269,N_14283,N_14713);
and UO_1270 (O_1270,N_14469,N_13523);
and UO_1271 (O_1271,N_13958,N_14584);
xor UO_1272 (O_1272,N_14957,N_13645);
nor UO_1273 (O_1273,N_14324,N_13755);
or UO_1274 (O_1274,N_13580,N_13814);
nor UO_1275 (O_1275,N_13778,N_13527);
xnor UO_1276 (O_1276,N_14558,N_13747);
nor UO_1277 (O_1277,N_14814,N_14739);
or UO_1278 (O_1278,N_14440,N_13850);
nand UO_1279 (O_1279,N_14488,N_13675);
nor UO_1280 (O_1280,N_14129,N_14793);
nand UO_1281 (O_1281,N_13524,N_14454);
nor UO_1282 (O_1282,N_13910,N_14123);
or UO_1283 (O_1283,N_14549,N_14222);
or UO_1284 (O_1284,N_14031,N_14651);
and UO_1285 (O_1285,N_14689,N_14440);
and UO_1286 (O_1286,N_14291,N_13908);
nand UO_1287 (O_1287,N_14589,N_14253);
nor UO_1288 (O_1288,N_14633,N_14804);
xor UO_1289 (O_1289,N_14982,N_13897);
xor UO_1290 (O_1290,N_14518,N_13537);
or UO_1291 (O_1291,N_13514,N_14190);
nor UO_1292 (O_1292,N_14292,N_14939);
nand UO_1293 (O_1293,N_14449,N_14416);
nand UO_1294 (O_1294,N_14287,N_14093);
xor UO_1295 (O_1295,N_14531,N_13690);
and UO_1296 (O_1296,N_13553,N_14131);
nor UO_1297 (O_1297,N_13646,N_14745);
nand UO_1298 (O_1298,N_13534,N_13934);
or UO_1299 (O_1299,N_13555,N_14825);
nand UO_1300 (O_1300,N_13654,N_14173);
xor UO_1301 (O_1301,N_14538,N_14303);
or UO_1302 (O_1302,N_13863,N_14229);
nand UO_1303 (O_1303,N_14754,N_14745);
xnor UO_1304 (O_1304,N_13829,N_14594);
xor UO_1305 (O_1305,N_14589,N_13598);
nor UO_1306 (O_1306,N_14100,N_14207);
nor UO_1307 (O_1307,N_14140,N_14063);
and UO_1308 (O_1308,N_14485,N_14923);
xor UO_1309 (O_1309,N_14306,N_14433);
xor UO_1310 (O_1310,N_14485,N_14576);
and UO_1311 (O_1311,N_14354,N_14137);
nor UO_1312 (O_1312,N_14771,N_14486);
nand UO_1313 (O_1313,N_14364,N_14458);
or UO_1314 (O_1314,N_14098,N_14888);
or UO_1315 (O_1315,N_14053,N_14596);
nand UO_1316 (O_1316,N_13537,N_14581);
nand UO_1317 (O_1317,N_14530,N_14422);
nand UO_1318 (O_1318,N_14250,N_14912);
xor UO_1319 (O_1319,N_13872,N_14095);
nor UO_1320 (O_1320,N_13756,N_13929);
xnor UO_1321 (O_1321,N_14447,N_14054);
nand UO_1322 (O_1322,N_14253,N_14243);
nor UO_1323 (O_1323,N_14229,N_13695);
xnor UO_1324 (O_1324,N_13797,N_14460);
or UO_1325 (O_1325,N_14147,N_14099);
nand UO_1326 (O_1326,N_14959,N_14162);
or UO_1327 (O_1327,N_14237,N_14261);
nand UO_1328 (O_1328,N_14438,N_13664);
nor UO_1329 (O_1329,N_14527,N_14268);
nor UO_1330 (O_1330,N_13706,N_13519);
nand UO_1331 (O_1331,N_13874,N_14417);
and UO_1332 (O_1332,N_14930,N_14552);
nand UO_1333 (O_1333,N_13955,N_14335);
or UO_1334 (O_1334,N_14767,N_13644);
nor UO_1335 (O_1335,N_13600,N_14869);
nand UO_1336 (O_1336,N_14762,N_14878);
nand UO_1337 (O_1337,N_13884,N_14212);
nand UO_1338 (O_1338,N_13874,N_14051);
nand UO_1339 (O_1339,N_14300,N_14612);
nand UO_1340 (O_1340,N_14352,N_14076);
and UO_1341 (O_1341,N_13980,N_14572);
nor UO_1342 (O_1342,N_13979,N_14853);
and UO_1343 (O_1343,N_13914,N_13721);
xor UO_1344 (O_1344,N_14845,N_14482);
xnor UO_1345 (O_1345,N_14851,N_14609);
nor UO_1346 (O_1346,N_14206,N_14495);
nand UO_1347 (O_1347,N_14205,N_14950);
and UO_1348 (O_1348,N_13814,N_14208);
nand UO_1349 (O_1349,N_14851,N_14172);
or UO_1350 (O_1350,N_14966,N_14917);
or UO_1351 (O_1351,N_14957,N_14209);
xnor UO_1352 (O_1352,N_14873,N_14078);
xnor UO_1353 (O_1353,N_13634,N_14503);
nor UO_1354 (O_1354,N_14246,N_13652);
nand UO_1355 (O_1355,N_14647,N_14374);
nand UO_1356 (O_1356,N_13529,N_14576);
and UO_1357 (O_1357,N_14953,N_14445);
nand UO_1358 (O_1358,N_14408,N_13603);
xnor UO_1359 (O_1359,N_13910,N_14004);
and UO_1360 (O_1360,N_13618,N_13549);
xor UO_1361 (O_1361,N_14515,N_14700);
nand UO_1362 (O_1362,N_14146,N_14648);
or UO_1363 (O_1363,N_14770,N_13688);
or UO_1364 (O_1364,N_13823,N_14550);
nor UO_1365 (O_1365,N_14218,N_13588);
nor UO_1366 (O_1366,N_14107,N_13845);
xor UO_1367 (O_1367,N_14148,N_14789);
nand UO_1368 (O_1368,N_13761,N_14021);
nand UO_1369 (O_1369,N_14370,N_14661);
nor UO_1370 (O_1370,N_13759,N_13717);
nor UO_1371 (O_1371,N_14705,N_14479);
and UO_1372 (O_1372,N_14821,N_14292);
xnor UO_1373 (O_1373,N_14340,N_13868);
xor UO_1374 (O_1374,N_14835,N_14877);
nand UO_1375 (O_1375,N_14132,N_13616);
and UO_1376 (O_1376,N_14490,N_13649);
and UO_1377 (O_1377,N_14816,N_14379);
and UO_1378 (O_1378,N_14271,N_14414);
xnor UO_1379 (O_1379,N_14385,N_14971);
nor UO_1380 (O_1380,N_13754,N_13860);
or UO_1381 (O_1381,N_14073,N_14764);
nand UO_1382 (O_1382,N_14464,N_14774);
nand UO_1383 (O_1383,N_13808,N_14453);
nor UO_1384 (O_1384,N_14858,N_14412);
and UO_1385 (O_1385,N_13870,N_13916);
or UO_1386 (O_1386,N_13617,N_13818);
nor UO_1387 (O_1387,N_13641,N_14314);
or UO_1388 (O_1388,N_14624,N_13964);
nor UO_1389 (O_1389,N_14862,N_14141);
nor UO_1390 (O_1390,N_14836,N_13608);
xnor UO_1391 (O_1391,N_14382,N_14605);
or UO_1392 (O_1392,N_14320,N_14544);
and UO_1393 (O_1393,N_14548,N_13786);
nor UO_1394 (O_1394,N_14648,N_14659);
or UO_1395 (O_1395,N_13961,N_14992);
or UO_1396 (O_1396,N_14566,N_13567);
nand UO_1397 (O_1397,N_14608,N_14535);
or UO_1398 (O_1398,N_13528,N_14318);
nor UO_1399 (O_1399,N_14014,N_14316);
or UO_1400 (O_1400,N_13918,N_13906);
xnor UO_1401 (O_1401,N_14527,N_13656);
or UO_1402 (O_1402,N_13969,N_14172);
or UO_1403 (O_1403,N_14046,N_14845);
xnor UO_1404 (O_1404,N_14886,N_13575);
nand UO_1405 (O_1405,N_14285,N_13560);
and UO_1406 (O_1406,N_14700,N_14245);
and UO_1407 (O_1407,N_14616,N_13711);
and UO_1408 (O_1408,N_14730,N_14654);
nor UO_1409 (O_1409,N_14973,N_13907);
and UO_1410 (O_1410,N_13730,N_14248);
nand UO_1411 (O_1411,N_13779,N_14494);
and UO_1412 (O_1412,N_14981,N_13591);
and UO_1413 (O_1413,N_14652,N_14877);
nor UO_1414 (O_1414,N_13815,N_14597);
or UO_1415 (O_1415,N_14395,N_14964);
and UO_1416 (O_1416,N_14785,N_14994);
nand UO_1417 (O_1417,N_14451,N_14515);
xor UO_1418 (O_1418,N_14094,N_14377);
nor UO_1419 (O_1419,N_13806,N_14471);
or UO_1420 (O_1420,N_13819,N_13710);
nand UO_1421 (O_1421,N_14026,N_13739);
and UO_1422 (O_1422,N_14512,N_14536);
or UO_1423 (O_1423,N_13699,N_14641);
and UO_1424 (O_1424,N_14206,N_13961);
xnor UO_1425 (O_1425,N_13916,N_13565);
and UO_1426 (O_1426,N_13777,N_14810);
nand UO_1427 (O_1427,N_14599,N_14163);
and UO_1428 (O_1428,N_13859,N_14199);
nand UO_1429 (O_1429,N_14145,N_14081);
xnor UO_1430 (O_1430,N_14437,N_13510);
xnor UO_1431 (O_1431,N_14304,N_14692);
nand UO_1432 (O_1432,N_14642,N_14278);
nor UO_1433 (O_1433,N_14877,N_13793);
nand UO_1434 (O_1434,N_14232,N_14027);
xor UO_1435 (O_1435,N_14510,N_13849);
and UO_1436 (O_1436,N_14581,N_14241);
nand UO_1437 (O_1437,N_14443,N_14832);
xor UO_1438 (O_1438,N_13504,N_14608);
xnor UO_1439 (O_1439,N_14807,N_13740);
or UO_1440 (O_1440,N_13519,N_14690);
and UO_1441 (O_1441,N_14241,N_14101);
nand UO_1442 (O_1442,N_13678,N_13732);
nor UO_1443 (O_1443,N_14616,N_13823);
and UO_1444 (O_1444,N_14666,N_14057);
xor UO_1445 (O_1445,N_14153,N_14229);
or UO_1446 (O_1446,N_13655,N_14731);
or UO_1447 (O_1447,N_14743,N_14751);
xor UO_1448 (O_1448,N_13880,N_13800);
and UO_1449 (O_1449,N_13619,N_14943);
or UO_1450 (O_1450,N_14364,N_14968);
nand UO_1451 (O_1451,N_14521,N_14613);
nor UO_1452 (O_1452,N_14018,N_13834);
nand UO_1453 (O_1453,N_14448,N_14818);
and UO_1454 (O_1454,N_14707,N_14368);
nor UO_1455 (O_1455,N_13705,N_13513);
nor UO_1456 (O_1456,N_14082,N_14159);
nor UO_1457 (O_1457,N_14437,N_14185);
and UO_1458 (O_1458,N_14758,N_13599);
nand UO_1459 (O_1459,N_14314,N_14810);
nand UO_1460 (O_1460,N_14439,N_14319);
nand UO_1461 (O_1461,N_13728,N_14424);
nand UO_1462 (O_1462,N_14495,N_14725);
xnor UO_1463 (O_1463,N_14181,N_13941);
and UO_1464 (O_1464,N_14087,N_13806);
nor UO_1465 (O_1465,N_14874,N_14212);
xor UO_1466 (O_1466,N_14205,N_14238);
nor UO_1467 (O_1467,N_14598,N_13735);
or UO_1468 (O_1468,N_14911,N_14124);
nor UO_1469 (O_1469,N_14521,N_14313);
or UO_1470 (O_1470,N_14578,N_14139);
nor UO_1471 (O_1471,N_13773,N_14385);
nand UO_1472 (O_1472,N_14259,N_14988);
nor UO_1473 (O_1473,N_13658,N_14225);
nor UO_1474 (O_1474,N_13912,N_13920);
nand UO_1475 (O_1475,N_14427,N_14733);
or UO_1476 (O_1476,N_14185,N_13894);
nor UO_1477 (O_1477,N_13553,N_14526);
xor UO_1478 (O_1478,N_13898,N_13535);
xor UO_1479 (O_1479,N_14303,N_14007);
nand UO_1480 (O_1480,N_14240,N_13586);
nand UO_1481 (O_1481,N_14757,N_13757);
and UO_1482 (O_1482,N_13752,N_14271);
nor UO_1483 (O_1483,N_13603,N_14493);
and UO_1484 (O_1484,N_13726,N_14752);
or UO_1485 (O_1485,N_14935,N_14873);
xnor UO_1486 (O_1486,N_13877,N_14644);
nand UO_1487 (O_1487,N_14888,N_14296);
xor UO_1488 (O_1488,N_14860,N_14859);
or UO_1489 (O_1489,N_14185,N_14575);
and UO_1490 (O_1490,N_14270,N_14457);
xor UO_1491 (O_1491,N_14158,N_14516);
and UO_1492 (O_1492,N_13759,N_14528);
or UO_1493 (O_1493,N_14075,N_14544);
and UO_1494 (O_1494,N_14620,N_14879);
or UO_1495 (O_1495,N_13862,N_13846);
nor UO_1496 (O_1496,N_13537,N_14871);
and UO_1497 (O_1497,N_14287,N_14241);
xor UO_1498 (O_1498,N_14502,N_14558);
nand UO_1499 (O_1499,N_14746,N_13810);
and UO_1500 (O_1500,N_14338,N_13580);
and UO_1501 (O_1501,N_14204,N_13685);
xor UO_1502 (O_1502,N_13667,N_14286);
xor UO_1503 (O_1503,N_14594,N_14060);
and UO_1504 (O_1504,N_14166,N_13972);
nand UO_1505 (O_1505,N_14417,N_14776);
nor UO_1506 (O_1506,N_13837,N_14584);
and UO_1507 (O_1507,N_13612,N_14599);
nand UO_1508 (O_1508,N_14862,N_13669);
nor UO_1509 (O_1509,N_13880,N_14819);
and UO_1510 (O_1510,N_14390,N_14477);
or UO_1511 (O_1511,N_13517,N_14453);
and UO_1512 (O_1512,N_14455,N_14155);
and UO_1513 (O_1513,N_14361,N_14035);
or UO_1514 (O_1514,N_13553,N_14833);
xor UO_1515 (O_1515,N_13633,N_14600);
nand UO_1516 (O_1516,N_14216,N_14569);
nor UO_1517 (O_1517,N_14175,N_14633);
and UO_1518 (O_1518,N_14613,N_14227);
nand UO_1519 (O_1519,N_13860,N_14051);
nor UO_1520 (O_1520,N_14758,N_14443);
and UO_1521 (O_1521,N_14704,N_14881);
nor UO_1522 (O_1522,N_14788,N_13740);
xnor UO_1523 (O_1523,N_13952,N_13641);
xor UO_1524 (O_1524,N_13682,N_13653);
nor UO_1525 (O_1525,N_14706,N_13705);
nand UO_1526 (O_1526,N_13856,N_14937);
and UO_1527 (O_1527,N_14279,N_14942);
and UO_1528 (O_1528,N_14226,N_14954);
nor UO_1529 (O_1529,N_13960,N_14966);
nor UO_1530 (O_1530,N_14200,N_13863);
and UO_1531 (O_1531,N_13749,N_13526);
xor UO_1532 (O_1532,N_14011,N_14708);
or UO_1533 (O_1533,N_13677,N_14460);
xor UO_1534 (O_1534,N_14959,N_13761);
and UO_1535 (O_1535,N_14213,N_14938);
or UO_1536 (O_1536,N_13719,N_13763);
or UO_1537 (O_1537,N_14067,N_14271);
and UO_1538 (O_1538,N_14347,N_14693);
xnor UO_1539 (O_1539,N_13867,N_13880);
xor UO_1540 (O_1540,N_14703,N_14793);
and UO_1541 (O_1541,N_14799,N_13572);
or UO_1542 (O_1542,N_13627,N_14902);
or UO_1543 (O_1543,N_14918,N_14538);
and UO_1544 (O_1544,N_13977,N_13582);
xor UO_1545 (O_1545,N_14435,N_13865);
xnor UO_1546 (O_1546,N_13771,N_14733);
nand UO_1547 (O_1547,N_14697,N_14059);
nor UO_1548 (O_1548,N_14416,N_13931);
and UO_1549 (O_1549,N_14674,N_14489);
and UO_1550 (O_1550,N_13843,N_13642);
and UO_1551 (O_1551,N_14961,N_13634);
or UO_1552 (O_1552,N_13571,N_13604);
nor UO_1553 (O_1553,N_14072,N_13981);
nand UO_1554 (O_1554,N_14316,N_13897);
nand UO_1555 (O_1555,N_14610,N_14958);
nand UO_1556 (O_1556,N_13976,N_14983);
nor UO_1557 (O_1557,N_13655,N_13557);
xor UO_1558 (O_1558,N_14375,N_13852);
and UO_1559 (O_1559,N_14722,N_13717);
or UO_1560 (O_1560,N_13890,N_14020);
and UO_1561 (O_1561,N_14649,N_13964);
nand UO_1562 (O_1562,N_14213,N_14695);
xnor UO_1563 (O_1563,N_14534,N_14502);
xnor UO_1564 (O_1564,N_14500,N_14299);
nand UO_1565 (O_1565,N_14100,N_14110);
or UO_1566 (O_1566,N_14183,N_14955);
or UO_1567 (O_1567,N_13703,N_13621);
nand UO_1568 (O_1568,N_14302,N_14111);
nand UO_1569 (O_1569,N_14456,N_13678);
or UO_1570 (O_1570,N_14147,N_14064);
nand UO_1571 (O_1571,N_14626,N_14456);
xnor UO_1572 (O_1572,N_14877,N_14378);
xor UO_1573 (O_1573,N_14636,N_13880);
or UO_1574 (O_1574,N_14641,N_14179);
xor UO_1575 (O_1575,N_14500,N_14641);
or UO_1576 (O_1576,N_14236,N_13723);
and UO_1577 (O_1577,N_14194,N_14057);
and UO_1578 (O_1578,N_13854,N_14892);
or UO_1579 (O_1579,N_14084,N_14757);
and UO_1580 (O_1580,N_13748,N_14407);
and UO_1581 (O_1581,N_13843,N_13815);
xnor UO_1582 (O_1582,N_14246,N_14625);
nor UO_1583 (O_1583,N_13992,N_13665);
or UO_1584 (O_1584,N_14005,N_14876);
xor UO_1585 (O_1585,N_14245,N_13816);
xnor UO_1586 (O_1586,N_13845,N_13580);
nand UO_1587 (O_1587,N_13703,N_14617);
nand UO_1588 (O_1588,N_13736,N_14698);
nor UO_1589 (O_1589,N_13994,N_14726);
or UO_1590 (O_1590,N_14932,N_14195);
and UO_1591 (O_1591,N_13615,N_13758);
xor UO_1592 (O_1592,N_14238,N_14159);
xor UO_1593 (O_1593,N_14012,N_14693);
and UO_1594 (O_1594,N_13965,N_13727);
or UO_1595 (O_1595,N_14457,N_14907);
and UO_1596 (O_1596,N_13582,N_13967);
xnor UO_1597 (O_1597,N_13617,N_14314);
nand UO_1598 (O_1598,N_14976,N_14685);
nand UO_1599 (O_1599,N_14075,N_13707);
nor UO_1600 (O_1600,N_14976,N_14893);
and UO_1601 (O_1601,N_13852,N_14359);
xor UO_1602 (O_1602,N_14410,N_14614);
nand UO_1603 (O_1603,N_14843,N_13848);
nor UO_1604 (O_1604,N_14223,N_14600);
nor UO_1605 (O_1605,N_13884,N_14831);
nor UO_1606 (O_1606,N_14099,N_13963);
xor UO_1607 (O_1607,N_14203,N_14681);
nand UO_1608 (O_1608,N_13888,N_14752);
or UO_1609 (O_1609,N_14398,N_13569);
xnor UO_1610 (O_1610,N_14600,N_14743);
nor UO_1611 (O_1611,N_13576,N_14457);
xnor UO_1612 (O_1612,N_14500,N_14960);
and UO_1613 (O_1613,N_14971,N_14779);
and UO_1614 (O_1614,N_14644,N_13616);
and UO_1615 (O_1615,N_14616,N_14953);
and UO_1616 (O_1616,N_13534,N_14672);
xor UO_1617 (O_1617,N_13745,N_14437);
xor UO_1618 (O_1618,N_13695,N_14371);
nor UO_1619 (O_1619,N_13732,N_14278);
nand UO_1620 (O_1620,N_13716,N_13848);
or UO_1621 (O_1621,N_14524,N_13766);
and UO_1622 (O_1622,N_14662,N_14961);
xor UO_1623 (O_1623,N_14981,N_13526);
or UO_1624 (O_1624,N_14670,N_14258);
xor UO_1625 (O_1625,N_14745,N_14216);
xnor UO_1626 (O_1626,N_13854,N_14065);
nor UO_1627 (O_1627,N_13616,N_14816);
or UO_1628 (O_1628,N_14076,N_14459);
xnor UO_1629 (O_1629,N_14469,N_14332);
nor UO_1630 (O_1630,N_14192,N_14067);
nand UO_1631 (O_1631,N_13998,N_13553);
nand UO_1632 (O_1632,N_14961,N_14738);
nand UO_1633 (O_1633,N_14806,N_13910);
xor UO_1634 (O_1634,N_13515,N_13549);
xor UO_1635 (O_1635,N_14105,N_14714);
xnor UO_1636 (O_1636,N_14690,N_13989);
and UO_1637 (O_1637,N_14502,N_13820);
nand UO_1638 (O_1638,N_13586,N_14406);
nand UO_1639 (O_1639,N_13699,N_14606);
nor UO_1640 (O_1640,N_14083,N_14178);
or UO_1641 (O_1641,N_13956,N_13616);
or UO_1642 (O_1642,N_14036,N_14324);
or UO_1643 (O_1643,N_14946,N_14943);
or UO_1644 (O_1644,N_14732,N_13967);
xor UO_1645 (O_1645,N_13598,N_14645);
and UO_1646 (O_1646,N_14043,N_13916);
nand UO_1647 (O_1647,N_13630,N_13919);
nand UO_1648 (O_1648,N_14898,N_14831);
nor UO_1649 (O_1649,N_14980,N_14186);
and UO_1650 (O_1650,N_14177,N_14817);
xor UO_1651 (O_1651,N_14529,N_13732);
nor UO_1652 (O_1652,N_14274,N_14587);
and UO_1653 (O_1653,N_13819,N_13658);
nor UO_1654 (O_1654,N_13950,N_14759);
xnor UO_1655 (O_1655,N_13828,N_14528);
nor UO_1656 (O_1656,N_13561,N_13839);
nand UO_1657 (O_1657,N_14070,N_14130);
nand UO_1658 (O_1658,N_14425,N_13864);
or UO_1659 (O_1659,N_13682,N_14784);
xor UO_1660 (O_1660,N_14060,N_14668);
or UO_1661 (O_1661,N_14903,N_14547);
nor UO_1662 (O_1662,N_14098,N_14833);
and UO_1663 (O_1663,N_13642,N_14574);
nor UO_1664 (O_1664,N_14798,N_14326);
and UO_1665 (O_1665,N_14413,N_13972);
nand UO_1666 (O_1666,N_14746,N_14187);
nand UO_1667 (O_1667,N_14282,N_14497);
xor UO_1668 (O_1668,N_13885,N_14953);
xnor UO_1669 (O_1669,N_14984,N_13924);
and UO_1670 (O_1670,N_14689,N_13844);
or UO_1671 (O_1671,N_14737,N_14793);
or UO_1672 (O_1672,N_14657,N_14385);
and UO_1673 (O_1673,N_14067,N_14879);
xnor UO_1674 (O_1674,N_13643,N_14306);
xor UO_1675 (O_1675,N_14592,N_13952);
or UO_1676 (O_1676,N_14341,N_13795);
nor UO_1677 (O_1677,N_14103,N_14686);
nor UO_1678 (O_1678,N_14023,N_14643);
and UO_1679 (O_1679,N_14071,N_14118);
nor UO_1680 (O_1680,N_13575,N_14186);
or UO_1681 (O_1681,N_14815,N_13558);
nor UO_1682 (O_1682,N_14320,N_14713);
nor UO_1683 (O_1683,N_14556,N_14736);
and UO_1684 (O_1684,N_14298,N_13601);
or UO_1685 (O_1685,N_14101,N_14076);
nand UO_1686 (O_1686,N_13772,N_13895);
nor UO_1687 (O_1687,N_14031,N_14759);
or UO_1688 (O_1688,N_14024,N_14662);
and UO_1689 (O_1689,N_14019,N_14845);
and UO_1690 (O_1690,N_14881,N_14993);
and UO_1691 (O_1691,N_14937,N_13637);
xnor UO_1692 (O_1692,N_14300,N_14418);
and UO_1693 (O_1693,N_13997,N_13947);
nand UO_1694 (O_1694,N_14807,N_14054);
xor UO_1695 (O_1695,N_14908,N_14050);
nor UO_1696 (O_1696,N_14325,N_13505);
or UO_1697 (O_1697,N_14169,N_14731);
xor UO_1698 (O_1698,N_14400,N_14982);
nor UO_1699 (O_1699,N_14438,N_13939);
nand UO_1700 (O_1700,N_13524,N_13786);
nand UO_1701 (O_1701,N_13597,N_14471);
nand UO_1702 (O_1702,N_14107,N_14557);
nand UO_1703 (O_1703,N_14503,N_14230);
nand UO_1704 (O_1704,N_13577,N_14857);
and UO_1705 (O_1705,N_13956,N_13815);
nand UO_1706 (O_1706,N_13957,N_14717);
nor UO_1707 (O_1707,N_14355,N_14892);
xnor UO_1708 (O_1708,N_14462,N_14155);
nand UO_1709 (O_1709,N_13800,N_14289);
nand UO_1710 (O_1710,N_14114,N_14159);
and UO_1711 (O_1711,N_14848,N_14221);
xnor UO_1712 (O_1712,N_13641,N_14806);
and UO_1713 (O_1713,N_14681,N_14487);
nor UO_1714 (O_1714,N_14648,N_14115);
nor UO_1715 (O_1715,N_14388,N_14847);
xor UO_1716 (O_1716,N_14143,N_14200);
xnor UO_1717 (O_1717,N_13520,N_13794);
nor UO_1718 (O_1718,N_13725,N_14969);
or UO_1719 (O_1719,N_13532,N_14111);
nor UO_1720 (O_1720,N_14297,N_14513);
xor UO_1721 (O_1721,N_14456,N_14672);
nor UO_1722 (O_1722,N_14358,N_14780);
nand UO_1723 (O_1723,N_14327,N_14422);
or UO_1724 (O_1724,N_14615,N_14225);
xor UO_1725 (O_1725,N_13938,N_14110);
and UO_1726 (O_1726,N_14582,N_14016);
xnor UO_1727 (O_1727,N_13556,N_13627);
xor UO_1728 (O_1728,N_14544,N_14981);
or UO_1729 (O_1729,N_14686,N_14216);
and UO_1730 (O_1730,N_13676,N_14567);
or UO_1731 (O_1731,N_13508,N_14629);
nand UO_1732 (O_1732,N_14833,N_14057);
xor UO_1733 (O_1733,N_14872,N_13519);
nand UO_1734 (O_1734,N_13737,N_13721);
nor UO_1735 (O_1735,N_14369,N_14872);
nor UO_1736 (O_1736,N_14699,N_13831);
and UO_1737 (O_1737,N_14004,N_14882);
or UO_1738 (O_1738,N_14239,N_13896);
nor UO_1739 (O_1739,N_14230,N_14464);
or UO_1740 (O_1740,N_14720,N_14607);
or UO_1741 (O_1741,N_13989,N_13751);
xnor UO_1742 (O_1742,N_14454,N_14385);
xnor UO_1743 (O_1743,N_13715,N_13705);
or UO_1744 (O_1744,N_14650,N_14306);
nor UO_1745 (O_1745,N_14875,N_13936);
xor UO_1746 (O_1746,N_14222,N_14955);
and UO_1747 (O_1747,N_14324,N_13614);
nor UO_1748 (O_1748,N_14243,N_13725);
or UO_1749 (O_1749,N_14000,N_13654);
nor UO_1750 (O_1750,N_14546,N_14070);
and UO_1751 (O_1751,N_14981,N_14595);
nand UO_1752 (O_1752,N_14095,N_13712);
nand UO_1753 (O_1753,N_13973,N_14656);
xnor UO_1754 (O_1754,N_14371,N_13801);
and UO_1755 (O_1755,N_13645,N_13980);
or UO_1756 (O_1756,N_14064,N_14848);
nand UO_1757 (O_1757,N_14156,N_14364);
nand UO_1758 (O_1758,N_14704,N_13960);
xnor UO_1759 (O_1759,N_13919,N_14978);
and UO_1760 (O_1760,N_13712,N_13745);
and UO_1761 (O_1761,N_14924,N_14388);
nand UO_1762 (O_1762,N_14263,N_14660);
and UO_1763 (O_1763,N_13616,N_13611);
nand UO_1764 (O_1764,N_14625,N_13660);
or UO_1765 (O_1765,N_13892,N_14611);
nor UO_1766 (O_1766,N_14059,N_14945);
nor UO_1767 (O_1767,N_14824,N_14452);
nand UO_1768 (O_1768,N_14907,N_14380);
nand UO_1769 (O_1769,N_14692,N_13771);
xnor UO_1770 (O_1770,N_14574,N_14038);
or UO_1771 (O_1771,N_13995,N_14118);
nand UO_1772 (O_1772,N_14589,N_13834);
xor UO_1773 (O_1773,N_14899,N_14893);
nand UO_1774 (O_1774,N_14871,N_14136);
or UO_1775 (O_1775,N_14578,N_13590);
and UO_1776 (O_1776,N_13552,N_14976);
and UO_1777 (O_1777,N_14656,N_13564);
xnor UO_1778 (O_1778,N_13946,N_14415);
and UO_1779 (O_1779,N_14535,N_14133);
xor UO_1780 (O_1780,N_13737,N_14774);
xor UO_1781 (O_1781,N_13683,N_14673);
and UO_1782 (O_1782,N_14566,N_13826);
nor UO_1783 (O_1783,N_13771,N_14826);
or UO_1784 (O_1784,N_14842,N_14884);
or UO_1785 (O_1785,N_14445,N_13588);
and UO_1786 (O_1786,N_14506,N_14496);
nor UO_1787 (O_1787,N_14354,N_14942);
or UO_1788 (O_1788,N_14922,N_13924);
or UO_1789 (O_1789,N_14656,N_14496);
nor UO_1790 (O_1790,N_14856,N_14729);
xnor UO_1791 (O_1791,N_14644,N_14711);
xnor UO_1792 (O_1792,N_13603,N_14131);
nand UO_1793 (O_1793,N_14307,N_13599);
xor UO_1794 (O_1794,N_13870,N_14216);
nand UO_1795 (O_1795,N_14165,N_14888);
or UO_1796 (O_1796,N_14275,N_14515);
xor UO_1797 (O_1797,N_14090,N_13793);
and UO_1798 (O_1798,N_13648,N_13595);
xnor UO_1799 (O_1799,N_14032,N_14154);
or UO_1800 (O_1800,N_13619,N_14060);
nor UO_1801 (O_1801,N_14218,N_14252);
and UO_1802 (O_1802,N_14757,N_14179);
xor UO_1803 (O_1803,N_13924,N_14081);
nor UO_1804 (O_1804,N_14574,N_14870);
xnor UO_1805 (O_1805,N_14243,N_14212);
and UO_1806 (O_1806,N_14007,N_13562);
and UO_1807 (O_1807,N_14820,N_14594);
or UO_1808 (O_1808,N_13817,N_13777);
nand UO_1809 (O_1809,N_13796,N_14775);
and UO_1810 (O_1810,N_13723,N_13590);
and UO_1811 (O_1811,N_14662,N_13645);
and UO_1812 (O_1812,N_14687,N_13981);
nor UO_1813 (O_1813,N_14465,N_13504);
and UO_1814 (O_1814,N_14172,N_14875);
nand UO_1815 (O_1815,N_14143,N_14667);
nor UO_1816 (O_1816,N_14634,N_14724);
and UO_1817 (O_1817,N_14215,N_14281);
or UO_1818 (O_1818,N_13846,N_13960);
xnor UO_1819 (O_1819,N_14558,N_14431);
nor UO_1820 (O_1820,N_14248,N_14356);
xor UO_1821 (O_1821,N_14360,N_14378);
or UO_1822 (O_1822,N_14811,N_14898);
nor UO_1823 (O_1823,N_13978,N_13837);
xnor UO_1824 (O_1824,N_14244,N_13889);
or UO_1825 (O_1825,N_14527,N_14791);
or UO_1826 (O_1826,N_13996,N_13842);
nand UO_1827 (O_1827,N_14627,N_13800);
nor UO_1828 (O_1828,N_14266,N_13966);
nand UO_1829 (O_1829,N_13505,N_14031);
or UO_1830 (O_1830,N_13782,N_14523);
nor UO_1831 (O_1831,N_14547,N_14659);
or UO_1832 (O_1832,N_14552,N_14895);
or UO_1833 (O_1833,N_13566,N_14150);
or UO_1834 (O_1834,N_14644,N_14627);
xor UO_1835 (O_1835,N_14471,N_13803);
xnor UO_1836 (O_1836,N_14262,N_13925);
nor UO_1837 (O_1837,N_14137,N_14558);
xnor UO_1838 (O_1838,N_14240,N_14417);
and UO_1839 (O_1839,N_14464,N_14252);
xnor UO_1840 (O_1840,N_14744,N_14245);
or UO_1841 (O_1841,N_14552,N_14880);
xnor UO_1842 (O_1842,N_13681,N_13936);
or UO_1843 (O_1843,N_14692,N_13743);
or UO_1844 (O_1844,N_14717,N_14564);
nand UO_1845 (O_1845,N_14538,N_13927);
and UO_1846 (O_1846,N_14072,N_14078);
nor UO_1847 (O_1847,N_14503,N_14201);
xnor UO_1848 (O_1848,N_13697,N_14484);
and UO_1849 (O_1849,N_14813,N_14379);
or UO_1850 (O_1850,N_13728,N_14020);
and UO_1851 (O_1851,N_14041,N_14358);
and UO_1852 (O_1852,N_14645,N_14516);
or UO_1853 (O_1853,N_14174,N_14769);
and UO_1854 (O_1854,N_14875,N_13671);
and UO_1855 (O_1855,N_14921,N_14197);
xnor UO_1856 (O_1856,N_13512,N_13645);
and UO_1857 (O_1857,N_14822,N_14848);
nor UO_1858 (O_1858,N_14757,N_13845);
and UO_1859 (O_1859,N_14711,N_13525);
nor UO_1860 (O_1860,N_14782,N_13850);
xnor UO_1861 (O_1861,N_14308,N_14045);
nand UO_1862 (O_1862,N_13745,N_14322);
nor UO_1863 (O_1863,N_14593,N_14930);
nor UO_1864 (O_1864,N_13805,N_13605);
or UO_1865 (O_1865,N_14486,N_13717);
nand UO_1866 (O_1866,N_13884,N_14944);
or UO_1867 (O_1867,N_14560,N_14628);
and UO_1868 (O_1868,N_14219,N_13504);
and UO_1869 (O_1869,N_14933,N_14799);
nand UO_1870 (O_1870,N_13645,N_14021);
xnor UO_1871 (O_1871,N_14118,N_14342);
nor UO_1872 (O_1872,N_14839,N_13918);
and UO_1873 (O_1873,N_13766,N_14638);
xnor UO_1874 (O_1874,N_14375,N_14285);
nand UO_1875 (O_1875,N_14498,N_13833);
xnor UO_1876 (O_1876,N_13506,N_14003);
xor UO_1877 (O_1877,N_14294,N_13656);
and UO_1878 (O_1878,N_14200,N_14862);
xor UO_1879 (O_1879,N_14170,N_14496);
and UO_1880 (O_1880,N_14263,N_14563);
nand UO_1881 (O_1881,N_14734,N_13675);
or UO_1882 (O_1882,N_13514,N_13848);
xnor UO_1883 (O_1883,N_14310,N_13567);
xnor UO_1884 (O_1884,N_14814,N_14779);
xnor UO_1885 (O_1885,N_14218,N_14890);
and UO_1886 (O_1886,N_13964,N_14229);
nand UO_1887 (O_1887,N_14159,N_14980);
and UO_1888 (O_1888,N_14603,N_13693);
nand UO_1889 (O_1889,N_14532,N_14684);
nand UO_1890 (O_1890,N_14928,N_14213);
or UO_1891 (O_1891,N_13561,N_14969);
or UO_1892 (O_1892,N_14590,N_14508);
or UO_1893 (O_1893,N_14160,N_14186);
xor UO_1894 (O_1894,N_14450,N_14644);
nand UO_1895 (O_1895,N_13602,N_14472);
and UO_1896 (O_1896,N_14342,N_14510);
or UO_1897 (O_1897,N_13695,N_14278);
nand UO_1898 (O_1898,N_13922,N_14526);
nor UO_1899 (O_1899,N_14175,N_14433);
and UO_1900 (O_1900,N_14860,N_13990);
and UO_1901 (O_1901,N_14839,N_14692);
nand UO_1902 (O_1902,N_13635,N_13926);
nor UO_1903 (O_1903,N_14836,N_14802);
xor UO_1904 (O_1904,N_13656,N_13985);
xnor UO_1905 (O_1905,N_14875,N_13581);
nor UO_1906 (O_1906,N_14093,N_13803);
or UO_1907 (O_1907,N_14953,N_13547);
nor UO_1908 (O_1908,N_13703,N_14523);
and UO_1909 (O_1909,N_14683,N_14573);
nor UO_1910 (O_1910,N_14434,N_13579);
nand UO_1911 (O_1911,N_13619,N_13814);
nand UO_1912 (O_1912,N_14028,N_13704);
xnor UO_1913 (O_1913,N_14024,N_14246);
or UO_1914 (O_1914,N_14785,N_14453);
nand UO_1915 (O_1915,N_14272,N_14362);
and UO_1916 (O_1916,N_13889,N_13581);
nor UO_1917 (O_1917,N_14619,N_14295);
nor UO_1918 (O_1918,N_14435,N_14746);
nor UO_1919 (O_1919,N_14945,N_14301);
and UO_1920 (O_1920,N_14168,N_14374);
xnor UO_1921 (O_1921,N_13728,N_14729);
nand UO_1922 (O_1922,N_13911,N_13874);
or UO_1923 (O_1923,N_13618,N_14839);
nor UO_1924 (O_1924,N_14012,N_14068);
or UO_1925 (O_1925,N_14864,N_14644);
nand UO_1926 (O_1926,N_14034,N_14557);
nand UO_1927 (O_1927,N_13993,N_14861);
nor UO_1928 (O_1928,N_14325,N_13717);
and UO_1929 (O_1929,N_14900,N_14497);
nor UO_1930 (O_1930,N_14205,N_14831);
nand UO_1931 (O_1931,N_14267,N_13847);
nor UO_1932 (O_1932,N_14097,N_13511);
nor UO_1933 (O_1933,N_14201,N_14498);
xor UO_1934 (O_1934,N_14691,N_14643);
xor UO_1935 (O_1935,N_14522,N_13863);
or UO_1936 (O_1936,N_14717,N_14318);
xor UO_1937 (O_1937,N_14748,N_13870);
or UO_1938 (O_1938,N_14142,N_14579);
and UO_1939 (O_1939,N_13697,N_14011);
nand UO_1940 (O_1940,N_14430,N_13893);
nand UO_1941 (O_1941,N_13580,N_13645);
xor UO_1942 (O_1942,N_14259,N_14149);
nand UO_1943 (O_1943,N_13523,N_14227);
nor UO_1944 (O_1944,N_14256,N_14189);
nand UO_1945 (O_1945,N_14583,N_14177);
xnor UO_1946 (O_1946,N_14609,N_13618);
nor UO_1947 (O_1947,N_14632,N_14166);
nand UO_1948 (O_1948,N_13631,N_14128);
nand UO_1949 (O_1949,N_14701,N_13567);
nand UO_1950 (O_1950,N_14398,N_14630);
nand UO_1951 (O_1951,N_14639,N_14019);
nand UO_1952 (O_1952,N_14820,N_14318);
nand UO_1953 (O_1953,N_13660,N_14917);
or UO_1954 (O_1954,N_13975,N_13591);
nand UO_1955 (O_1955,N_14594,N_14189);
xnor UO_1956 (O_1956,N_14647,N_13946);
nand UO_1957 (O_1957,N_13884,N_14862);
xnor UO_1958 (O_1958,N_14754,N_13786);
nand UO_1959 (O_1959,N_14038,N_13519);
xnor UO_1960 (O_1960,N_14604,N_14368);
nand UO_1961 (O_1961,N_14286,N_13752);
and UO_1962 (O_1962,N_13793,N_13960);
nor UO_1963 (O_1963,N_14015,N_13682);
or UO_1964 (O_1964,N_14347,N_14003);
xnor UO_1965 (O_1965,N_13783,N_14134);
or UO_1966 (O_1966,N_14926,N_13856);
xnor UO_1967 (O_1967,N_14947,N_14001);
or UO_1968 (O_1968,N_14820,N_13981);
nand UO_1969 (O_1969,N_14325,N_14094);
nor UO_1970 (O_1970,N_13561,N_13803);
nor UO_1971 (O_1971,N_14235,N_14408);
or UO_1972 (O_1972,N_13573,N_13896);
nand UO_1973 (O_1973,N_14450,N_14342);
and UO_1974 (O_1974,N_14847,N_14546);
and UO_1975 (O_1975,N_14441,N_14941);
nor UO_1976 (O_1976,N_13703,N_14255);
or UO_1977 (O_1977,N_14419,N_14594);
nand UO_1978 (O_1978,N_13680,N_13702);
and UO_1979 (O_1979,N_14354,N_14745);
nor UO_1980 (O_1980,N_13569,N_14947);
or UO_1981 (O_1981,N_14947,N_14882);
and UO_1982 (O_1982,N_13900,N_13666);
nor UO_1983 (O_1983,N_14634,N_14807);
or UO_1984 (O_1984,N_14951,N_14927);
and UO_1985 (O_1985,N_14540,N_13958);
nor UO_1986 (O_1986,N_14536,N_14870);
nor UO_1987 (O_1987,N_14112,N_14649);
xnor UO_1988 (O_1988,N_14212,N_14946);
nand UO_1989 (O_1989,N_13740,N_14708);
or UO_1990 (O_1990,N_13894,N_14552);
nand UO_1991 (O_1991,N_14928,N_13725);
or UO_1992 (O_1992,N_14174,N_14789);
or UO_1993 (O_1993,N_14780,N_13556);
nand UO_1994 (O_1994,N_14437,N_14416);
nor UO_1995 (O_1995,N_13716,N_14879);
nand UO_1996 (O_1996,N_14157,N_14522);
nand UO_1997 (O_1997,N_14331,N_14230);
and UO_1998 (O_1998,N_13581,N_13786);
and UO_1999 (O_1999,N_14640,N_14262);
endmodule