module basic_750_5000_1000_25_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
xnor U0 (N_0,In_210,In_336);
or U1 (N_1,In_537,In_280);
nand U2 (N_2,In_675,In_161);
nand U3 (N_3,In_410,In_163);
or U4 (N_4,In_439,In_729);
xor U5 (N_5,In_368,In_631);
xnor U6 (N_6,In_86,In_718);
nand U7 (N_7,In_618,In_355);
nor U8 (N_8,In_571,In_424);
nor U9 (N_9,In_349,In_674);
or U10 (N_10,In_38,In_331);
or U11 (N_11,In_185,In_353);
xnor U12 (N_12,In_712,In_141);
xor U13 (N_13,In_722,In_427);
xor U14 (N_14,In_447,In_272);
nand U15 (N_15,In_79,In_364);
and U16 (N_16,In_232,In_545);
or U17 (N_17,In_189,In_226);
or U18 (N_18,In_714,In_154);
xnor U19 (N_19,In_463,In_68);
nand U20 (N_20,In_651,In_291);
nand U21 (N_21,In_170,In_602);
nand U22 (N_22,In_159,In_107);
nor U23 (N_23,In_670,In_337);
xor U24 (N_24,In_378,In_274);
xnor U25 (N_25,In_564,In_322);
xnor U26 (N_26,In_743,In_438);
nand U27 (N_27,In_307,In_190);
nor U28 (N_28,In_739,In_487);
or U29 (N_29,In_339,In_301);
or U30 (N_30,In_153,In_299);
nand U31 (N_31,In_333,In_471);
nor U32 (N_32,In_453,In_483);
xor U33 (N_33,In_741,In_746);
and U34 (N_34,In_318,In_546);
nand U35 (N_35,In_166,In_91);
or U36 (N_36,In_199,In_476);
and U37 (N_37,In_366,In_112);
xnor U38 (N_38,In_541,In_628);
nand U39 (N_39,In_17,In_623);
nor U40 (N_40,In_691,In_576);
nand U41 (N_41,In_127,In_627);
xor U42 (N_42,In_397,In_48);
xor U43 (N_43,In_491,In_32);
nand U44 (N_44,In_694,In_417);
and U45 (N_45,In_432,In_281);
and U46 (N_46,In_401,In_367);
and U47 (N_47,In_237,In_229);
and U48 (N_48,In_109,In_589);
nand U49 (N_49,In_196,In_707);
xnor U50 (N_50,In_300,In_225);
nand U51 (N_51,In_309,In_180);
nor U52 (N_52,In_239,In_358);
nor U53 (N_53,In_70,In_55);
xnor U54 (N_54,In_634,In_136);
or U55 (N_55,In_332,In_202);
or U56 (N_56,In_535,In_678);
or U57 (N_57,In_516,In_24);
or U58 (N_58,In_175,In_108);
nand U59 (N_59,In_494,In_5);
xnor U60 (N_60,In_591,In_615);
xor U61 (N_61,In_636,In_482);
nand U62 (N_62,In_104,In_523);
or U63 (N_63,In_560,In_134);
xor U64 (N_64,In_744,In_46);
nor U65 (N_65,In_182,In_611);
and U66 (N_66,In_408,In_446);
and U67 (N_67,In_128,In_29);
or U68 (N_68,In_305,In_548);
xor U69 (N_69,In_0,In_215);
or U70 (N_70,In_462,In_216);
nand U71 (N_71,In_220,In_735);
or U72 (N_72,In_486,In_533);
nor U73 (N_73,In_177,In_413);
nor U74 (N_74,In_686,In_534);
nor U75 (N_75,In_635,In_688);
and U76 (N_76,In_121,In_713);
or U77 (N_77,In_525,In_458);
xor U78 (N_78,In_49,In_478);
and U79 (N_79,In_261,In_338);
nand U80 (N_80,In_664,In_363);
nor U81 (N_81,In_372,In_450);
xnor U82 (N_82,In_371,In_573);
or U83 (N_83,In_479,In_47);
xor U84 (N_84,In_286,In_71);
nor U85 (N_85,In_633,In_143);
or U86 (N_86,In_257,In_164);
nand U87 (N_87,In_357,In_96);
nand U88 (N_88,In_666,In_474);
nand U89 (N_89,In_467,In_724);
and U90 (N_90,In_391,In_85);
or U91 (N_91,In_477,In_461);
and U92 (N_92,In_704,In_61);
nor U93 (N_93,In_640,In_661);
nor U94 (N_94,In_81,In_431);
nand U95 (N_95,In_264,In_122);
and U96 (N_96,In_552,In_579);
xor U97 (N_97,In_437,In_749);
and U98 (N_98,In_76,In_659);
or U99 (N_99,In_470,In_64);
nor U100 (N_100,In_39,In_6);
nand U101 (N_101,In_245,In_53);
nand U102 (N_102,In_99,In_456);
and U103 (N_103,In_669,In_130);
or U104 (N_104,In_473,In_97);
nand U105 (N_105,In_673,In_587);
xnor U106 (N_106,In_619,In_303);
xnor U107 (N_107,In_208,In_649);
and U108 (N_108,In_599,In_582);
nor U109 (N_109,In_510,In_517);
nor U110 (N_110,In_379,In_279);
nand U111 (N_111,In_147,In_736);
xor U112 (N_112,In_296,In_551);
xnor U113 (N_113,In_526,In_335);
xor U114 (N_114,In_621,In_711);
nor U115 (N_115,In_205,In_341);
nor U116 (N_116,In_359,In_35);
xnor U117 (N_117,In_186,In_455);
nand U118 (N_118,In_65,In_62);
and U119 (N_119,In_69,In_183);
nand U120 (N_120,In_209,In_464);
nand U121 (N_121,In_43,In_689);
nand U122 (N_122,In_740,In_402);
nor U123 (N_123,In_100,In_265);
xnor U124 (N_124,In_643,In_558);
nor U125 (N_125,In_601,In_441);
or U126 (N_126,In_387,In_681);
nor U127 (N_127,In_512,In_313);
nor U128 (N_128,In_256,In_652);
or U129 (N_129,In_481,In_683);
xnor U130 (N_130,In_241,In_613);
and U131 (N_131,In_319,In_422);
nand U132 (N_132,In_668,In_416);
nand U133 (N_133,In_728,In_234);
xor U134 (N_134,In_275,In_298);
xor U135 (N_135,In_50,In_259);
nand U136 (N_136,In_734,In_562);
or U137 (N_137,In_197,In_568);
nor U138 (N_138,In_88,In_213);
or U139 (N_139,In_733,In_547);
and U140 (N_140,In_556,In_608);
nor U141 (N_141,In_224,In_513);
nand U142 (N_142,In_521,In_263);
nand U143 (N_143,In_382,In_30);
xnor U144 (N_144,In_529,In_14);
or U145 (N_145,In_472,In_444);
xnor U146 (N_146,In_16,In_460);
nand U147 (N_147,In_351,In_609);
and U148 (N_148,In_87,In_114);
nand U149 (N_149,In_41,In_110);
nor U150 (N_150,In_191,In_699);
nor U151 (N_151,In_373,In_346);
nor U152 (N_152,In_392,In_612);
or U153 (N_153,In_594,In_252);
nand U154 (N_154,In_705,In_129);
nor U155 (N_155,In_721,In_505);
xor U156 (N_156,In_747,In_95);
and U157 (N_157,In_409,In_327);
nand U158 (N_158,In_414,In_13);
or U159 (N_159,In_730,In_420);
nand U160 (N_160,In_187,In_273);
nor U161 (N_161,In_266,In_44);
xnor U162 (N_162,In_403,In_555);
nand U163 (N_163,In_42,In_503);
or U164 (N_164,In_680,In_51);
or U165 (N_165,In_698,In_146);
or U166 (N_166,In_126,In_550);
nand U167 (N_167,In_287,In_421);
and U168 (N_168,In_459,In_231);
xnor U169 (N_169,In_246,In_727);
nor U170 (N_170,In_433,In_198);
nand U171 (N_171,In_221,In_277);
or U172 (N_172,In_26,In_235);
xnor U173 (N_173,In_7,In_243);
nor U174 (N_174,In_250,In_696);
nand U175 (N_175,In_192,In_34);
and U176 (N_176,In_278,In_148);
or U177 (N_177,In_646,In_748);
nand U178 (N_178,In_394,In_11);
xor U179 (N_179,In_247,In_524);
xnor U180 (N_180,In_742,In_536);
nand U181 (N_181,In_329,In_701);
xnor U182 (N_182,In_285,In_518);
and U183 (N_183,In_574,In_12);
and U184 (N_184,In_625,In_629);
or U185 (N_185,In_267,In_253);
or U186 (N_186,In_15,In_345);
nand U187 (N_187,In_78,In_726);
and U188 (N_188,In_632,In_554);
and U189 (N_189,In_489,In_667);
xor U190 (N_190,In_36,In_106);
and U191 (N_191,In_706,In_124);
nor U192 (N_192,In_268,In_18);
and U193 (N_193,In_238,In_665);
nand U194 (N_194,In_288,In_223);
and U195 (N_195,In_290,In_607);
and U196 (N_196,In_151,In_425);
nor U197 (N_197,In_93,In_142);
and U198 (N_198,In_448,In_436);
or U199 (N_199,In_644,In_2);
nand U200 (N_200,N_74,In_375);
xor U201 (N_201,In_328,N_69);
nand U202 (N_202,In_119,In_655);
xor U203 (N_203,In_527,In_181);
nand U204 (N_204,In_600,N_53);
and U205 (N_205,N_190,In_731);
nand U206 (N_206,N_156,N_64);
xor U207 (N_207,N_130,N_5);
nor U208 (N_208,In_501,N_114);
nand U209 (N_209,In_693,N_164);
or U210 (N_210,In_67,In_228);
nor U211 (N_211,N_175,In_138);
xor U212 (N_212,In_217,N_50);
nor U213 (N_213,In_588,N_16);
xnor U214 (N_214,In_384,In_271);
xnor U215 (N_215,In_380,N_124);
or U216 (N_216,N_36,N_117);
nand U217 (N_217,In_679,In_73);
nor U218 (N_218,N_63,In_630);
nor U219 (N_219,In_567,In_9);
xnor U220 (N_220,In_398,In_738);
or U221 (N_221,N_67,In_155);
and U222 (N_222,N_60,N_177);
xor U223 (N_223,In_492,In_74);
or U224 (N_224,N_176,In_411);
nor U225 (N_225,In_145,In_393);
and U226 (N_226,N_111,In_212);
nor U227 (N_227,In_395,N_86);
nor U228 (N_228,In_654,N_187);
and U229 (N_229,N_195,N_140);
nand U230 (N_230,In_101,In_519);
and U231 (N_231,In_412,N_71);
or U232 (N_232,N_101,N_192);
nor U233 (N_233,In_449,In_314);
and U234 (N_234,In_248,In_317);
nand U235 (N_235,In_311,In_330);
xor U236 (N_236,In_572,N_57);
nand U237 (N_237,In_348,In_687);
nor U238 (N_238,In_703,In_528);
or U239 (N_239,In_222,In_484);
and U240 (N_240,In_639,In_28);
nor U241 (N_241,N_49,In_137);
xor U242 (N_242,N_30,In_566);
and U243 (N_243,In_430,N_72);
nand U244 (N_244,N_158,In_658);
and U245 (N_245,In_542,N_70);
xor U246 (N_246,N_39,In_140);
nor U247 (N_247,In_139,In_720);
nand U248 (N_248,In_475,N_55);
xor U249 (N_249,N_99,N_149);
or U250 (N_250,N_38,In_451);
or U251 (N_251,In_496,N_35);
or U252 (N_252,In_3,In_544);
xnor U253 (N_253,In_52,In_227);
xor U254 (N_254,N_107,In_376);
or U255 (N_255,In_258,N_17);
nand U256 (N_256,N_155,In_648);
xnor U257 (N_257,In_169,In_206);
or U258 (N_258,N_106,In_115);
nor U259 (N_259,In_662,In_125);
nand U260 (N_260,N_85,N_79);
nor U261 (N_261,In_719,N_29);
xnor U262 (N_262,In_581,In_63);
nor U263 (N_263,In_506,In_56);
xnor U264 (N_264,N_137,N_24);
nand U265 (N_265,In_251,In_435);
nand U266 (N_266,In_157,N_198);
nor U267 (N_267,In_321,In_428);
xor U268 (N_268,N_51,In_236);
nand U269 (N_269,N_47,In_709);
xor U270 (N_270,In_171,N_4);
nand U271 (N_271,In_660,In_406);
xnor U272 (N_272,N_142,In_624);
or U273 (N_273,N_73,In_653);
nor U274 (N_274,In_304,In_493);
and U275 (N_275,N_95,In_334);
or U276 (N_276,In_80,N_109);
nor U277 (N_277,N_185,In_57);
or U278 (N_278,N_128,In_324);
and U279 (N_279,N_143,In_443);
nor U280 (N_280,In_66,N_19);
nor U281 (N_281,In_116,In_715);
nand U282 (N_282,N_15,In_559);
or U283 (N_283,In_295,In_203);
nor U284 (N_284,In_539,In_89);
xor U285 (N_285,N_62,In_174);
xor U286 (N_286,In_495,In_214);
and U287 (N_287,In_504,In_72);
and U288 (N_288,In_45,In_585);
nand U289 (N_289,N_126,In_452);
xnor U290 (N_290,N_112,In_19);
nor U291 (N_291,In_242,N_148);
nor U292 (N_292,N_160,In_350);
or U293 (N_293,In_656,In_400);
nor U294 (N_294,In_75,In_604);
nor U295 (N_295,In_593,N_1);
nand U296 (N_296,N_196,In_194);
nor U297 (N_297,In_343,N_171);
nor U298 (N_298,In_440,N_27);
nand U299 (N_299,In_407,N_75);
and U300 (N_300,N_8,N_90);
nor U301 (N_301,In_383,In_162);
and U302 (N_302,In_284,N_32);
nand U303 (N_303,In_270,In_1);
or U304 (N_304,In_514,In_21);
or U305 (N_305,N_59,N_102);
xnor U306 (N_306,In_173,N_173);
or U307 (N_307,In_282,In_293);
nand U308 (N_308,In_60,In_603);
xnor U309 (N_309,N_129,In_294);
and U310 (N_310,N_34,In_429);
nor U311 (N_311,In_418,In_94);
and U312 (N_312,In_240,In_82);
or U313 (N_313,In_365,In_188);
and U314 (N_314,In_302,In_732);
and U315 (N_315,In_480,In_549);
xor U316 (N_316,N_123,In_283);
or U317 (N_317,N_121,In_445);
nor U318 (N_318,In_207,In_710);
and U319 (N_319,In_316,In_133);
and U320 (N_320,In_276,N_12);
and U321 (N_321,In_386,In_507);
xnor U322 (N_322,N_76,N_81);
or U323 (N_323,N_84,In_320);
xor U324 (N_324,In_465,In_176);
and U325 (N_325,N_197,In_59);
or U326 (N_326,In_325,N_108);
xnor U327 (N_327,In_637,In_399);
nand U328 (N_328,In_531,In_626);
nor U329 (N_329,N_98,N_23);
xnor U330 (N_330,In_538,N_163);
or U331 (N_331,In_158,In_614);
or U332 (N_332,In_672,In_310);
xnor U333 (N_333,In_415,N_25);
xor U334 (N_334,In_340,In_219);
xor U335 (N_335,N_159,N_166);
or U336 (N_336,N_181,In_168);
or U337 (N_337,In_111,In_356);
nand U338 (N_338,In_23,N_152);
xor U339 (N_339,In_388,In_377);
nand U340 (N_340,In_716,N_44);
nor U341 (N_341,N_116,In_565);
xnor U342 (N_342,In_700,In_717);
nand U343 (N_343,In_113,In_499);
nand U344 (N_344,In_262,In_702);
and U345 (N_345,In_605,In_255);
nand U346 (N_346,In_434,N_87);
and U347 (N_347,In_369,In_269);
and U348 (N_348,N_7,In_543);
and U349 (N_349,N_33,In_58);
and U350 (N_350,In_557,In_598);
or U351 (N_351,In_360,In_583);
or U352 (N_352,In_532,In_561);
nand U353 (N_353,N_122,In_150);
xnor U354 (N_354,N_151,In_200);
and U355 (N_355,In_354,In_502);
and U356 (N_356,In_254,N_172);
nand U357 (N_357,N_184,In_22);
xnor U358 (N_358,In_663,N_9);
nor U359 (N_359,In_165,N_189);
xnor U360 (N_360,In_500,In_485);
and U361 (N_361,N_144,In_160);
xnor U362 (N_362,In_201,In_468);
nor U363 (N_363,N_131,In_563);
or U364 (N_364,In_211,In_570);
nand U365 (N_365,In_676,In_260);
nand U366 (N_366,In_520,In_620);
nand U367 (N_367,In_490,N_120);
xor U368 (N_368,In_144,N_3);
nand U369 (N_369,In_4,In_244);
or U370 (N_370,In_396,N_165);
xnor U371 (N_371,N_21,In_578);
or U372 (N_372,N_88,In_606);
nor U373 (N_373,In_149,N_147);
nand U374 (N_374,In_497,In_361);
nor U375 (N_375,In_645,N_119);
nand U376 (N_376,In_515,In_385);
or U377 (N_377,In_117,In_671);
nor U378 (N_378,In_616,In_657);
or U379 (N_379,In_592,In_131);
nand U380 (N_380,N_45,N_2);
or U381 (N_381,In_33,In_84);
nor U382 (N_382,In_347,In_423);
and U383 (N_383,N_54,N_167);
nand U384 (N_384,In_25,In_374);
or U385 (N_385,In_610,In_83);
and U386 (N_386,N_48,In_426);
and U387 (N_387,N_103,In_381);
and U388 (N_388,In_530,In_178);
nand U389 (N_389,In_580,N_191);
nand U390 (N_390,In_156,N_26);
and U391 (N_391,N_93,N_125);
nor U392 (N_392,In_90,In_723);
and U393 (N_393,N_65,In_195);
or U394 (N_394,In_697,In_184);
or U395 (N_395,N_133,In_362);
nor U396 (N_396,In_289,N_153);
nand U397 (N_397,In_204,N_96);
and U398 (N_398,N_83,N_10);
nor U399 (N_399,N_115,N_14);
or U400 (N_400,In_575,N_356);
or U401 (N_401,In_682,In_10);
or U402 (N_402,In_193,In_540);
xnor U403 (N_403,In_622,In_509);
nor U404 (N_404,N_350,N_274);
and U405 (N_405,In_553,N_247);
nor U406 (N_406,N_337,In_326);
nand U407 (N_407,N_391,N_234);
or U408 (N_408,N_135,N_328);
nand U409 (N_409,N_299,N_304);
nor U410 (N_410,N_20,N_218);
xor U411 (N_411,N_235,N_6);
nor U412 (N_412,N_310,N_217);
and U413 (N_413,N_221,N_344);
nand U414 (N_414,In_233,N_208);
nand U415 (N_415,N_272,In_249);
and U416 (N_416,N_56,N_361);
nor U417 (N_417,N_238,N_316);
or U418 (N_418,N_150,In_695);
xnor U419 (N_419,N_105,N_355);
nor U420 (N_420,N_216,N_389);
or U421 (N_421,N_286,N_209);
or U422 (N_422,In_27,In_469);
or U423 (N_423,N_275,N_385);
nand U424 (N_424,N_306,N_338);
or U425 (N_425,N_94,N_319);
xnor U426 (N_426,N_359,N_395);
and U427 (N_427,In_737,N_118);
or U428 (N_428,N_349,N_314);
or U429 (N_429,N_254,N_97);
or U430 (N_430,N_297,N_229);
or U431 (N_431,N_265,N_82);
xnor U432 (N_432,N_301,N_264);
nor U433 (N_433,N_322,In_442);
nor U434 (N_434,N_291,N_320);
xnor U435 (N_435,N_179,N_292);
or U436 (N_436,In_650,In_323);
nor U437 (N_437,N_362,N_373);
xnor U438 (N_438,N_382,N_226);
xor U439 (N_439,N_113,N_266);
xnor U440 (N_440,N_242,In_312);
and U441 (N_441,N_186,In_522);
nor U442 (N_442,In_586,In_152);
xnor U443 (N_443,N_332,N_146);
and U444 (N_444,In_8,N_245);
or U445 (N_445,In_488,In_306);
nand U446 (N_446,N_341,N_222);
xor U447 (N_447,N_379,N_110);
and U448 (N_448,N_330,N_295);
or U449 (N_449,N_255,N_296);
or U450 (N_450,In_120,N_225);
nor U451 (N_451,N_298,N_41);
or U452 (N_452,N_280,N_288);
xnor U453 (N_453,N_326,In_577);
nor U454 (N_454,In_105,N_240);
or U455 (N_455,N_154,N_368);
and U456 (N_456,N_244,N_258);
xor U457 (N_457,N_270,N_346);
and U458 (N_458,In_617,In_31);
nand U459 (N_459,N_46,N_308);
nand U460 (N_460,N_227,N_228);
and U461 (N_461,N_357,N_251);
and U462 (N_462,N_232,N_215);
nor U463 (N_463,N_268,N_61);
xor U464 (N_464,N_243,In_40);
or U465 (N_465,N_327,N_100);
or U466 (N_466,N_397,In_596);
nor U467 (N_467,N_263,N_277);
and U468 (N_468,N_206,N_211);
nor U469 (N_469,N_31,N_18);
nand U470 (N_470,N_388,In_230);
or U471 (N_471,N_241,N_269);
nor U472 (N_472,N_139,N_366);
or U473 (N_473,N_205,N_220);
and U474 (N_474,N_77,N_313);
and U475 (N_475,N_348,N_178);
and U476 (N_476,N_22,N_210);
or U477 (N_477,N_374,N_334);
nor U478 (N_478,N_300,N_194);
or U479 (N_479,In_390,N_257);
or U480 (N_480,N_305,N_261);
xor U481 (N_481,In_37,N_207);
and U482 (N_482,In_167,N_260);
nor U483 (N_483,N_342,N_352);
and U484 (N_484,In_135,N_294);
nand U485 (N_485,N_145,In_419);
or U486 (N_486,N_287,N_360);
xor U487 (N_487,N_293,N_170);
nand U488 (N_488,In_677,N_239);
and U489 (N_489,N_284,N_302);
nor U490 (N_490,N_384,N_283);
nand U491 (N_491,N_315,N_399);
nand U492 (N_492,In_389,In_685);
xor U493 (N_493,In_692,N_246);
or U494 (N_494,N_335,N_138);
or U495 (N_495,N_347,N_252);
xor U496 (N_496,N_324,N_136);
nor U497 (N_497,N_230,N_289);
nand U498 (N_498,N_168,N_13);
nor U499 (N_499,N_202,N_68);
nand U500 (N_500,In_584,N_392);
or U501 (N_501,N_312,N_345);
nand U502 (N_502,N_219,N_303);
or U503 (N_503,In_595,In_54);
or U504 (N_504,N_58,N_253);
xor U505 (N_505,N_398,N_193);
and U506 (N_506,In_344,N_372);
nand U507 (N_507,N_231,N_89);
and U508 (N_508,In_132,In_745);
or U509 (N_509,In_218,N_378);
nor U510 (N_510,N_351,In_297);
nor U511 (N_511,N_354,In_641);
nor U512 (N_512,N_11,N_162);
and U513 (N_513,N_267,In_102);
nand U514 (N_514,In_308,N_281);
nor U515 (N_515,N_317,N_157);
xnor U516 (N_516,N_141,N_381);
or U517 (N_517,In_708,N_376);
xnor U518 (N_518,In_457,N_183);
and U519 (N_519,N_199,N_329);
and U520 (N_520,N_212,In_352);
and U521 (N_521,N_307,N_200);
or U522 (N_522,N_278,N_224);
nor U523 (N_523,In_690,N_237);
and U524 (N_524,In_511,N_375);
nand U525 (N_525,N_396,N_182);
or U526 (N_526,N_37,N_259);
nand U527 (N_527,In_684,N_276);
and U528 (N_528,N_311,N_369);
nor U529 (N_529,In_370,N_250);
nor U530 (N_530,N_365,In_342);
and U531 (N_531,In_638,N_333);
nor U532 (N_532,N_380,N_248);
nor U533 (N_533,N_367,N_256);
or U534 (N_534,N_390,N_386);
nand U535 (N_535,N_358,In_123);
or U536 (N_536,N_309,N_370);
nand U537 (N_537,N_214,N_364);
nor U538 (N_538,N_127,In_569);
and U539 (N_539,N_174,N_28);
and U540 (N_540,In_597,N_132);
xnor U541 (N_541,N_290,N_262);
xor U542 (N_542,N_161,In_172);
and U543 (N_543,N_387,N_91);
and U544 (N_544,N_340,In_498);
xor U545 (N_545,In_642,N_134);
nor U546 (N_546,In_647,N_282);
xnor U547 (N_547,N_223,N_279);
nor U548 (N_548,N_249,In_98);
nand U549 (N_549,N_0,In_404);
nand U550 (N_550,N_180,N_393);
nor U551 (N_551,In_179,N_394);
xnor U552 (N_552,N_339,N_188);
nor U553 (N_553,N_201,N_92);
xor U554 (N_554,N_66,In_20);
or U555 (N_555,In_315,N_323);
and U556 (N_556,In_292,N_377);
xor U557 (N_557,N_321,In_454);
xnor U558 (N_558,N_371,N_169);
xor U559 (N_559,N_236,N_353);
nand U560 (N_560,N_43,In_92);
or U561 (N_561,N_203,N_363);
or U562 (N_562,N_78,N_42);
nor U563 (N_563,N_285,In_77);
and U564 (N_564,In_466,N_40);
or U565 (N_565,N_383,In_103);
and U566 (N_566,N_213,N_104);
nand U567 (N_567,N_336,N_80);
nand U568 (N_568,N_331,N_52);
nand U569 (N_569,N_325,In_590);
nand U570 (N_570,N_233,In_405);
xnor U571 (N_571,In_118,N_204);
xnor U572 (N_572,N_318,N_343);
and U573 (N_573,N_273,In_508);
nor U574 (N_574,N_271,In_725);
nand U575 (N_575,N_182,In_695);
xor U576 (N_576,In_584,In_641);
or U577 (N_577,N_325,In_466);
or U578 (N_578,N_300,N_249);
nor U579 (N_579,In_172,N_346);
or U580 (N_580,N_345,In_27);
or U581 (N_581,N_280,N_203);
nor U582 (N_582,N_241,N_261);
nand U583 (N_583,N_388,N_300);
nor U584 (N_584,N_372,N_246);
or U585 (N_585,N_344,N_292);
nand U586 (N_586,N_313,N_235);
or U587 (N_587,N_330,N_46);
nor U588 (N_588,N_334,N_221);
and U589 (N_589,N_292,N_240);
or U590 (N_590,N_110,N_295);
or U591 (N_591,N_323,N_309);
and U592 (N_592,N_343,In_522);
nand U593 (N_593,N_276,N_332);
nor U594 (N_594,In_390,N_274);
xnor U595 (N_595,N_246,N_284);
and U596 (N_596,N_346,In_708);
nor U597 (N_597,In_454,N_317);
and U598 (N_598,In_692,N_347);
xor U599 (N_599,N_399,N_288);
or U600 (N_600,N_466,N_538);
nand U601 (N_601,N_486,N_498);
and U602 (N_602,N_435,N_437);
nor U603 (N_603,N_467,N_500);
xor U604 (N_604,N_406,N_463);
nor U605 (N_605,N_457,N_413);
or U606 (N_606,N_442,N_520);
nand U607 (N_607,N_459,N_598);
nor U608 (N_608,N_562,N_454);
xnor U609 (N_609,N_560,N_495);
nor U610 (N_610,N_576,N_582);
or U611 (N_611,N_402,N_419);
xnor U612 (N_612,N_439,N_533);
xor U613 (N_613,N_557,N_556);
xor U614 (N_614,N_455,N_438);
xnor U615 (N_615,N_541,N_404);
nand U616 (N_616,N_528,N_501);
or U617 (N_617,N_480,N_471);
nand U618 (N_618,N_496,N_552);
nand U619 (N_619,N_436,N_405);
or U620 (N_620,N_555,N_563);
and U621 (N_621,N_474,N_523);
and U622 (N_622,N_542,N_526);
and U623 (N_623,N_477,N_579);
and U624 (N_624,N_570,N_519);
xnor U625 (N_625,N_478,N_452);
nand U626 (N_626,N_529,N_517);
or U627 (N_627,N_456,N_532);
nor U628 (N_628,N_583,N_574);
nor U629 (N_629,N_535,N_482);
or U630 (N_630,N_411,N_472);
xnor U631 (N_631,N_580,N_485);
xor U632 (N_632,N_548,N_539);
or U633 (N_633,N_503,N_515);
nand U634 (N_634,N_420,N_481);
nor U635 (N_635,N_527,N_588);
xor U636 (N_636,N_427,N_475);
or U637 (N_637,N_429,N_468);
xnor U638 (N_638,N_561,N_508);
or U639 (N_639,N_446,N_421);
xnor U640 (N_640,N_423,N_566);
xnor U641 (N_641,N_531,N_403);
or U642 (N_642,N_537,N_569);
xnor U643 (N_643,N_502,N_441);
or U644 (N_644,N_511,N_567);
xnor U645 (N_645,N_543,N_564);
nand U646 (N_646,N_587,N_476);
and U647 (N_647,N_451,N_453);
xor U648 (N_648,N_469,N_492);
nand U649 (N_649,N_493,N_479);
xor U650 (N_650,N_445,N_595);
nor U651 (N_651,N_408,N_489);
or U652 (N_652,N_586,N_443);
nand U653 (N_653,N_449,N_521);
nor U654 (N_654,N_545,N_572);
nor U655 (N_655,N_447,N_464);
or U656 (N_656,N_575,N_462);
xor U657 (N_657,N_505,N_581);
or U658 (N_658,N_589,N_473);
xor U659 (N_659,N_510,N_596);
xor U660 (N_660,N_428,N_409);
xor U661 (N_661,N_460,N_544);
nand U662 (N_662,N_509,N_584);
xnor U663 (N_663,N_513,N_424);
or U664 (N_664,N_571,N_430);
and U665 (N_665,N_578,N_434);
xnor U666 (N_666,N_487,N_410);
or U667 (N_667,N_516,N_522);
and U668 (N_668,N_426,N_512);
nor U669 (N_669,N_534,N_416);
and U670 (N_670,N_490,N_553);
and U671 (N_671,N_431,N_558);
nor U672 (N_672,N_432,N_549);
nor U673 (N_673,N_577,N_497);
xor U674 (N_674,N_414,N_546);
xnor U675 (N_675,N_594,N_450);
nand U676 (N_676,N_568,N_524);
nor U677 (N_677,N_507,N_551);
and U678 (N_678,N_585,N_590);
nand U679 (N_679,N_565,N_483);
nor U680 (N_680,N_491,N_440);
xnor U681 (N_681,N_591,N_525);
nand U682 (N_682,N_412,N_407);
or U683 (N_683,N_592,N_550);
and U684 (N_684,N_506,N_499);
and U685 (N_685,N_461,N_417);
nand U686 (N_686,N_444,N_593);
nor U687 (N_687,N_488,N_418);
nand U688 (N_688,N_425,N_554);
nand U689 (N_689,N_433,N_401);
nand U690 (N_690,N_514,N_458);
nor U691 (N_691,N_400,N_530);
and U692 (N_692,N_484,N_599);
xnor U693 (N_693,N_597,N_448);
nor U694 (N_694,N_573,N_540);
or U695 (N_695,N_536,N_518);
nand U696 (N_696,N_422,N_415);
xnor U697 (N_697,N_470,N_547);
xnor U698 (N_698,N_504,N_494);
xor U699 (N_699,N_559,N_465);
or U700 (N_700,N_525,N_555);
xor U701 (N_701,N_409,N_572);
xor U702 (N_702,N_571,N_483);
nor U703 (N_703,N_529,N_549);
and U704 (N_704,N_493,N_554);
or U705 (N_705,N_593,N_538);
xor U706 (N_706,N_541,N_530);
xnor U707 (N_707,N_480,N_567);
and U708 (N_708,N_520,N_496);
and U709 (N_709,N_580,N_542);
nor U710 (N_710,N_441,N_541);
nand U711 (N_711,N_534,N_517);
xor U712 (N_712,N_584,N_425);
or U713 (N_713,N_561,N_569);
or U714 (N_714,N_511,N_441);
or U715 (N_715,N_599,N_481);
nor U716 (N_716,N_490,N_528);
xnor U717 (N_717,N_514,N_419);
nand U718 (N_718,N_537,N_567);
nand U719 (N_719,N_598,N_479);
and U720 (N_720,N_585,N_546);
nor U721 (N_721,N_539,N_467);
or U722 (N_722,N_413,N_515);
and U723 (N_723,N_537,N_452);
nor U724 (N_724,N_566,N_534);
nand U725 (N_725,N_485,N_475);
nor U726 (N_726,N_595,N_436);
or U727 (N_727,N_436,N_500);
nand U728 (N_728,N_414,N_563);
xnor U729 (N_729,N_522,N_541);
nand U730 (N_730,N_458,N_526);
or U731 (N_731,N_570,N_478);
nor U732 (N_732,N_569,N_442);
xnor U733 (N_733,N_514,N_598);
xor U734 (N_734,N_456,N_493);
and U735 (N_735,N_552,N_532);
nand U736 (N_736,N_558,N_546);
nand U737 (N_737,N_556,N_535);
and U738 (N_738,N_528,N_503);
or U739 (N_739,N_488,N_507);
nor U740 (N_740,N_434,N_449);
nor U741 (N_741,N_577,N_538);
nor U742 (N_742,N_428,N_578);
or U743 (N_743,N_437,N_595);
nand U744 (N_744,N_470,N_558);
or U745 (N_745,N_404,N_563);
nand U746 (N_746,N_527,N_530);
xor U747 (N_747,N_467,N_515);
nor U748 (N_748,N_485,N_527);
xor U749 (N_749,N_574,N_576);
or U750 (N_750,N_541,N_598);
xor U751 (N_751,N_572,N_460);
xor U752 (N_752,N_487,N_497);
xnor U753 (N_753,N_467,N_589);
or U754 (N_754,N_530,N_497);
nand U755 (N_755,N_407,N_548);
xnor U756 (N_756,N_423,N_561);
and U757 (N_757,N_584,N_547);
xnor U758 (N_758,N_401,N_597);
nor U759 (N_759,N_513,N_431);
or U760 (N_760,N_431,N_459);
nor U761 (N_761,N_564,N_597);
nor U762 (N_762,N_503,N_500);
nor U763 (N_763,N_553,N_518);
or U764 (N_764,N_559,N_534);
nand U765 (N_765,N_525,N_576);
or U766 (N_766,N_580,N_486);
xor U767 (N_767,N_443,N_524);
xor U768 (N_768,N_582,N_579);
xnor U769 (N_769,N_515,N_593);
or U770 (N_770,N_467,N_559);
nand U771 (N_771,N_444,N_408);
or U772 (N_772,N_455,N_544);
and U773 (N_773,N_457,N_422);
nor U774 (N_774,N_475,N_416);
xnor U775 (N_775,N_520,N_516);
nand U776 (N_776,N_400,N_536);
xor U777 (N_777,N_491,N_597);
nor U778 (N_778,N_526,N_468);
and U779 (N_779,N_417,N_595);
and U780 (N_780,N_509,N_548);
or U781 (N_781,N_418,N_433);
xnor U782 (N_782,N_463,N_500);
xor U783 (N_783,N_469,N_545);
and U784 (N_784,N_525,N_506);
nand U785 (N_785,N_540,N_428);
and U786 (N_786,N_455,N_543);
nor U787 (N_787,N_412,N_506);
xnor U788 (N_788,N_591,N_559);
nand U789 (N_789,N_416,N_564);
xor U790 (N_790,N_441,N_478);
nor U791 (N_791,N_427,N_516);
nor U792 (N_792,N_483,N_566);
or U793 (N_793,N_410,N_467);
nor U794 (N_794,N_446,N_567);
and U795 (N_795,N_499,N_463);
and U796 (N_796,N_556,N_596);
and U797 (N_797,N_513,N_467);
nor U798 (N_798,N_473,N_455);
nand U799 (N_799,N_522,N_457);
xnor U800 (N_800,N_721,N_671);
or U801 (N_801,N_623,N_787);
nand U802 (N_802,N_762,N_793);
nor U803 (N_803,N_622,N_741);
or U804 (N_804,N_690,N_694);
or U805 (N_805,N_669,N_699);
and U806 (N_806,N_778,N_604);
xnor U807 (N_807,N_666,N_737);
and U808 (N_808,N_620,N_766);
xor U809 (N_809,N_618,N_645);
xnor U810 (N_810,N_715,N_697);
and U811 (N_811,N_726,N_719);
nand U812 (N_812,N_689,N_722);
and U813 (N_813,N_747,N_750);
nand U814 (N_814,N_706,N_608);
and U815 (N_815,N_765,N_771);
xor U816 (N_816,N_630,N_643);
nand U817 (N_817,N_667,N_716);
xor U818 (N_818,N_711,N_703);
xor U819 (N_819,N_639,N_744);
nor U820 (N_820,N_635,N_627);
nand U821 (N_821,N_743,N_610);
xor U822 (N_822,N_712,N_634);
xnor U823 (N_823,N_674,N_767);
nand U824 (N_824,N_795,N_688);
and U825 (N_825,N_708,N_638);
and U826 (N_826,N_756,N_751);
or U827 (N_827,N_692,N_729);
and U828 (N_828,N_700,N_788);
and U829 (N_829,N_631,N_609);
and U830 (N_830,N_796,N_685);
and U831 (N_831,N_745,N_702);
or U832 (N_832,N_647,N_763);
and U833 (N_833,N_710,N_779);
and U834 (N_834,N_782,N_777);
nand U835 (N_835,N_728,N_730);
xor U836 (N_836,N_611,N_769);
xor U837 (N_837,N_676,N_601);
xor U838 (N_838,N_640,N_772);
and U839 (N_839,N_695,N_600);
xnor U840 (N_840,N_753,N_705);
and U841 (N_841,N_736,N_658);
and U842 (N_842,N_755,N_681);
and U843 (N_843,N_783,N_790);
nor U844 (N_844,N_785,N_748);
and U845 (N_845,N_642,N_625);
xor U846 (N_846,N_749,N_792);
xnor U847 (N_847,N_646,N_682);
nand U848 (N_848,N_607,N_636);
nand U849 (N_849,N_653,N_773);
xor U850 (N_850,N_686,N_780);
nor U851 (N_851,N_701,N_731);
xnor U852 (N_852,N_621,N_663);
nor U853 (N_853,N_675,N_746);
nand U854 (N_854,N_616,N_770);
or U855 (N_855,N_670,N_673);
xnor U856 (N_856,N_648,N_661);
nor U857 (N_857,N_678,N_735);
or U858 (N_858,N_624,N_633);
or U859 (N_859,N_628,N_776);
xor U860 (N_860,N_704,N_775);
or U861 (N_861,N_680,N_734);
and U862 (N_862,N_629,N_687);
or U863 (N_863,N_696,N_764);
nor U864 (N_864,N_717,N_672);
nand U865 (N_865,N_768,N_797);
and U866 (N_866,N_698,N_742);
nand U867 (N_867,N_794,N_709);
xor U868 (N_868,N_789,N_739);
nand U869 (N_869,N_752,N_761);
nand U870 (N_870,N_656,N_637);
xnor U871 (N_871,N_651,N_684);
nor U872 (N_872,N_665,N_727);
or U873 (N_873,N_732,N_664);
and U874 (N_874,N_791,N_798);
xnor U875 (N_875,N_723,N_774);
and U876 (N_876,N_724,N_654);
nor U877 (N_877,N_612,N_652);
nor U878 (N_878,N_693,N_668);
xnor U879 (N_879,N_786,N_660);
nand U880 (N_880,N_649,N_626);
or U881 (N_881,N_707,N_759);
and U882 (N_882,N_655,N_613);
nand U883 (N_883,N_781,N_677);
nand U884 (N_884,N_718,N_641);
and U885 (N_885,N_720,N_657);
or U886 (N_886,N_760,N_659);
nor U887 (N_887,N_679,N_757);
and U888 (N_888,N_606,N_615);
nand U889 (N_889,N_738,N_754);
nand U890 (N_890,N_714,N_683);
or U891 (N_891,N_784,N_619);
nand U892 (N_892,N_644,N_602);
and U893 (N_893,N_799,N_650);
xnor U894 (N_894,N_603,N_614);
or U895 (N_895,N_632,N_758);
xnor U896 (N_896,N_605,N_662);
or U897 (N_897,N_713,N_725);
and U898 (N_898,N_691,N_733);
or U899 (N_899,N_617,N_740);
and U900 (N_900,N_788,N_601);
nand U901 (N_901,N_708,N_667);
nor U902 (N_902,N_790,N_768);
and U903 (N_903,N_745,N_738);
xnor U904 (N_904,N_775,N_630);
nand U905 (N_905,N_754,N_714);
nand U906 (N_906,N_797,N_673);
or U907 (N_907,N_742,N_615);
and U908 (N_908,N_684,N_654);
nor U909 (N_909,N_689,N_762);
or U910 (N_910,N_657,N_755);
and U911 (N_911,N_783,N_782);
xor U912 (N_912,N_736,N_642);
or U913 (N_913,N_660,N_792);
xor U914 (N_914,N_658,N_621);
nor U915 (N_915,N_739,N_649);
nor U916 (N_916,N_618,N_783);
or U917 (N_917,N_634,N_720);
nor U918 (N_918,N_797,N_693);
xnor U919 (N_919,N_765,N_603);
and U920 (N_920,N_784,N_722);
nor U921 (N_921,N_676,N_635);
nor U922 (N_922,N_759,N_624);
nand U923 (N_923,N_629,N_659);
nor U924 (N_924,N_714,N_758);
or U925 (N_925,N_645,N_765);
nand U926 (N_926,N_756,N_613);
xnor U927 (N_927,N_632,N_673);
nand U928 (N_928,N_744,N_717);
or U929 (N_929,N_726,N_785);
or U930 (N_930,N_714,N_682);
and U931 (N_931,N_702,N_693);
and U932 (N_932,N_781,N_687);
nor U933 (N_933,N_765,N_732);
nand U934 (N_934,N_673,N_683);
and U935 (N_935,N_752,N_747);
nand U936 (N_936,N_635,N_678);
or U937 (N_937,N_694,N_711);
nand U938 (N_938,N_763,N_725);
nor U939 (N_939,N_787,N_708);
or U940 (N_940,N_793,N_765);
nand U941 (N_941,N_631,N_746);
nor U942 (N_942,N_741,N_787);
nor U943 (N_943,N_750,N_791);
xor U944 (N_944,N_692,N_695);
and U945 (N_945,N_758,N_797);
or U946 (N_946,N_677,N_672);
nor U947 (N_947,N_708,N_681);
xor U948 (N_948,N_762,N_773);
or U949 (N_949,N_722,N_668);
or U950 (N_950,N_767,N_775);
or U951 (N_951,N_741,N_792);
nand U952 (N_952,N_777,N_746);
nor U953 (N_953,N_659,N_702);
xor U954 (N_954,N_667,N_741);
xnor U955 (N_955,N_701,N_748);
nand U956 (N_956,N_732,N_747);
nor U957 (N_957,N_602,N_696);
nor U958 (N_958,N_730,N_623);
or U959 (N_959,N_666,N_796);
or U960 (N_960,N_715,N_764);
nor U961 (N_961,N_659,N_651);
or U962 (N_962,N_625,N_746);
and U963 (N_963,N_663,N_604);
xnor U964 (N_964,N_675,N_684);
xor U965 (N_965,N_703,N_675);
and U966 (N_966,N_613,N_740);
xnor U967 (N_967,N_605,N_732);
and U968 (N_968,N_710,N_652);
nand U969 (N_969,N_796,N_724);
and U970 (N_970,N_731,N_638);
nand U971 (N_971,N_691,N_739);
or U972 (N_972,N_660,N_670);
nand U973 (N_973,N_752,N_697);
nand U974 (N_974,N_702,N_610);
nand U975 (N_975,N_771,N_657);
nor U976 (N_976,N_750,N_660);
nor U977 (N_977,N_661,N_631);
nand U978 (N_978,N_692,N_632);
nand U979 (N_979,N_783,N_754);
or U980 (N_980,N_683,N_766);
nand U981 (N_981,N_607,N_673);
nand U982 (N_982,N_666,N_792);
or U983 (N_983,N_787,N_711);
and U984 (N_984,N_777,N_713);
nand U985 (N_985,N_671,N_621);
xor U986 (N_986,N_744,N_663);
and U987 (N_987,N_619,N_749);
or U988 (N_988,N_700,N_628);
nand U989 (N_989,N_612,N_604);
xnor U990 (N_990,N_662,N_754);
or U991 (N_991,N_762,N_710);
nand U992 (N_992,N_690,N_692);
and U993 (N_993,N_603,N_791);
nand U994 (N_994,N_767,N_600);
xor U995 (N_995,N_756,N_674);
or U996 (N_996,N_660,N_731);
nand U997 (N_997,N_766,N_758);
nand U998 (N_998,N_722,N_672);
nand U999 (N_999,N_714,N_681);
nand U1000 (N_1000,N_892,N_855);
nand U1001 (N_1001,N_831,N_947);
or U1002 (N_1002,N_896,N_980);
xnor U1003 (N_1003,N_827,N_894);
and U1004 (N_1004,N_978,N_888);
nand U1005 (N_1005,N_904,N_950);
xnor U1006 (N_1006,N_987,N_852);
xor U1007 (N_1007,N_971,N_990);
and U1008 (N_1008,N_865,N_966);
or U1009 (N_1009,N_840,N_999);
xnor U1010 (N_1010,N_908,N_948);
and U1011 (N_1011,N_870,N_905);
and U1012 (N_1012,N_997,N_820);
xor U1013 (N_1013,N_801,N_841);
and U1014 (N_1014,N_805,N_928);
xor U1015 (N_1015,N_880,N_961);
or U1016 (N_1016,N_810,N_906);
and U1017 (N_1017,N_926,N_834);
xor U1018 (N_1018,N_984,N_854);
and U1019 (N_1019,N_969,N_844);
xor U1020 (N_1020,N_821,N_995);
xor U1021 (N_1021,N_932,N_991);
xnor U1022 (N_1022,N_845,N_937);
nand U1023 (N_1023,N_815,N_863);
and U1024 (N_1024,N_998,N_806);
nor U1025 (N_1025,N_960,N_949);
xnor U1026 (N_1026,N_972,N_889);
and U1027 (N_1027,N_804,N_954);
xnor U1028 (N_1028,N_917,N_858);
and U1029 (N_1029,N_857,N_900);
and U1030 (N_1030,N_847,N_924);
and U1031 (N_1031,N_837,N_938);
xnor U1032 (N_1032,N_862,N_976);
nor U1033 (N_1033,N_802,N_989);
xnor U1034 (N_1034,N_903,N_835);
or U1035 (N_1035,N_881,N_945);
or U1036 (N_1036,N_901,N_920);
xor U1037 (N_1037,N_970,N_927);
or U1038 (N_1038,N_982,N_955);
and U1039 (N_1039,N_890,N_816);
or U1040 (N_1040,N_877,N_872);
nand U1041 (N_1041,N_957,N_964);
xnor U1042 (N_1042,N_823,N_981);
xor U1043 (N_1043,N_873,N_853);
xor U1044 (N_1044,N_883,N_811);
xnor U1045 (N_1045,N_848,N_897);
xor U1046 (N_1046,N_974,N_914);
xnor U1047 (N_1047,N_952,N_992);
xor U1048 (N_1048,N_922,N_887);
or U1049 (N_1049,N_986,N_979);
nand U1050 (N_1050,N_959,N_958);
or U1051 (N_1051,N_882,N_833);
nor U1052 (N_1052,N_910,N_830);
nor U1053 (N_1053,N_934,N_996);
nor U1054 (N_1054,N_867,N_921);
xnor U1055 (N_1055,N_838,N_916);
xor U1056 (N_1056,N_951,N_879);
nand U1057 (N_1057,N_943,N_925);
xor U1058 (N_1058,N_850,N_931);
xnor U1059 (N_1059,N_915,N_918);
or U1060 (N_1060,N_864,N_826);
xnor U1061 (N_1061,N_967,N_941);
nand U1062 (N_1062,N_907,N_983);
nand U1063 (N_1063,N_859,N_843);
xnor U1064 (N_1064,N_956,N_817);
xnor U1065 (N_1065,N_912,N_953);
nand U1066 (N_1066,N_885,N_860);
xnor U1067 (N_1067,N_936,N_836);
and U1068 (N_1068,N_993,N_869);
xnor U1069 (N_1069,N_876,N_994);
or U1070 (N_1070,N_962,N_985);
xor U1071 (N_1071,N_808,N_946);
nor U1072 (N_1072,N_988,N_828);
xor U1073 (N_1073,N_871,N_933);
nand U1074 (N_1074,N_824,N_891);
or U1075 (N_1075,N_803,N_944);
xnor U1076 (N_1076,N_913,N_800);
or U1077 (N_1077,N_814,N_919);
nor U1078 (N_1078,N_886,N_861);
nor U1079 (N_1079,N_930,N_973);
or U1080 (N_1080,N_893,N_968);
xor U1081 (N_1081,N_874,N_822);
and U1082 (N_1082,N_878,N_963);
nor U1083 (N_1083,N_832,N_809);
nand U1084 (N_1084,N_807,N_849);
nand U1085 (N_1085,N_813,N_899);
and U1086 (N_1086,N_965,N_929);
and U1087 (N_1087,N_942,N_923);
nor U1088 (N_1088,N_939,N_975);
or U1089 (N_1089,N_898,N_902);
or U1090 (N_1090,N_842,N_818);
and U1091 (N_1091,N_911,N_846);
and U1092 (N_1092,N_819,N_829);
nand U1093 (N_1093,N_977,N_851);
nor U1094 (N_1094,N_884,N_868);
nor U1095 (N_1095,N_825,N_856);
nor U1096 (N_1096,N_895,N_935);
xnor U1097 (N_1097,N_940,N_812);
or U1098 (N_1098,N_839,N_909);
or U1099 (N_1099,N_875,N_866);
and U1100 (N_1100,N_815,N_893);
and U1101 (N_1101,N_903,N_940);
nand U1102 (N_1102,N_898,N_928);
or U1103 (N_1103,N_934,N_819);
nor U1104 (N_1104,N_897,N_870);
nand U1105 (N_1105,N_939,N_868);
xor U1106 (N_1106,N_975,N_922);
or U1107 (N_1107,N_912,N_992);
or U1108 (N_1108,N_812,N_873);
nand U1109 (N_1109,N_851,N_815);
and U1110 (N_1110,N_902,N_801);
or U1111 (N_1111,N_865,N_846);
or U1112 (N_1112,N_869,N_962);
and U1113 (N_1113,N_808,N_952);
and U1114 (N_1114,N_933,N_829);
nor U1115 (N_1115,N_883,N_928);
nor U1116 (N_1116,N_803,N_812);
nor U1117 (N_1117,N_849,N_947);
or U1118 (N_1118,N_827,N_847);
nand U1119 (N_1119,N_946,N_851);
or U1120 (N_1120,N_853,N_924);
xor U1121 (N_1121,N_881,N_912);
or U1122 (N_1122,N_986,N_843);
nand U1123 (N_1123,N_992,N_977);
or U1124 (N_1124,N_829,N_967);
or U1125 (N_1125,N_839,N_871);
xor U1126 (N_1126,N_902,N_823);
and U1127 (N_1127,N_818,N_912);
nor U1128 (N_1128,N_968,N_857);
and U1129 (N_1129,N_803,N_874);
xnor U1130 (N_1130,N_896,N_804);
xor U1131 (N_1131,N_834,N_898);
xor U1132 (N_1132,N_957,N_976);
nand U1133 (N_1133,N_893,N_944);
nor U1134 (N_1134,N_949,N_993);
nand U1135 (N_1135,N_800,N_817);
and U1136 (N_1136,N_899,N_939);
nor U1137 (N_1137,N_895,N_810);
nand U1138 (N_1138,N_832,N_964);
xor U1139 (N_1139,N_850,N_814);
xor U1140 (N_1140,N_818,N_896);
or U1141 (N_1141,N_832,N_991);
xnor U1142 (N_1142,N_877,N_840);
or U1143 (N_1143,N_981,N_880);
or U1144 (N_1144,N_819,N_895);
nand U1145 (N_1145,N_814,N_959);
xnor U1146 (N_1146,N_978,N_937);
nor U1147 (N_1147,N_896,N_978);
or U1148 (N_1148,N_808,N_948);
nor U1149 (N_1149,N_967,N_955);
or U1150 (N_1150,N_819,N_970);
nand U1151 (N_1151,N_814,N_907);
and U1152 (N_1152,N_939,N_827);
nand U1153 (N_1153,N_899,N_866);
or U1154 (N_1154,N_929,N_874);
nor U1155 (N_1155,N_880,N_924);
xnor U1156 (N_1156,N_928,N_810);
xor U1157 (N_1157,N_902,N_907);
xnor U1158 (N_1158,N_839,N_948);
and U1159 (N_1159,N_909,N_942);
nand U1160 (N_1160,N_856,N_969);
nor U1161 (N_1161,N_939,N_937);
xnor U1162 (N_1162,N_857,N_850);
nand U1163 (N_1163,N_880,N_949);
nor U1164 (N_1164,N_926,N_939);
nor U1165 (N_1165,N_945,N_880);
nor U1166 (N_1166,N_941,N_901);
nor U1167 (N_1167,N_883,N_866);
nand U1168 (N_1168,N_856,N_895);
xnor U1169 (N_1169,N_967,N_943);
xor U1170 (N_1170,N_849,N_926);
and U1171 (N_1171,N_995,N_973);
and U1172 (N_1172,N_913,N_911);
nor U1173 (N_1173,N_821,N_892);
or U1174 (N_1174,N_904,N_892);
nand U1175 (N_1175,N_928,N_972);
nand U1176 (N_1176,N_897,N_948);
and U1177 (N_1177,N_875,N_948);
nand U1178 (N_1178,N_988,N_990);
nor U1179 (N_1179,N_968,N_838);
or U1180 (N_1180,N_877,N_957);
nor U1181 (N_1181,N_898,N_931);
xnor U1182 (N_1182,N_914,N_940);
nand U1183 (N_1183,N_826,N_861);
or U1184 (N_1184,N_955,N_947);
and U1185 (N_1185,N_972,N_893);
xor U1186 (N_1186,N_932,N_956);
xnor U1187 (N_1187,N_829,N_916);
and U1188 (N_1188,N_945,N_927);
nand U1189 (N_1189,N_847,N_810);
or U1190 (N_1190,N_961,N_970);
or U1191 (N_1191,N_833,N_915);
and U1192 (N_1192,N_801,N_812);
nor U1193 (N_1193,N_932,N_877);
nand U1194 (N_1194,N_846,N_993);
and U1195 (N_1195,N_841,N_945);
nand U1196 (N_1196,N_831,N_819);
nor U1197 (N_1197,N_854,N_906);
or U1198 (N_1198,N_949,N_953);
nor U1199 (N_1199,N_878,N_875);
xnor U1200 (N_1200,N_1171,N_1160);
nor U1201 (N_1201,N_1162,N_1099);
xor U1202 (N_1202,N_1066,N_1035);
xnor U1203 (N_1203,N_1033,N_1012);
nand U1204 (N_1204,N_1187,N_1190);
or U1205 (N_1205,N_1068,N_1036);
nand U1206 (N_1206,N_1023,N_1146);
and U1207 (N_1207,N_1089,N_1108);
xor U1208 (N_1208,N_1007,N_1060);
nand U1209 (N_1209,N_1085,N_1049);
nand U1210 (N_1210,N_1105,N_1013);
nand U1211 (N_1211,N_1073,N_1010);
nand U1212 (N_1212,N_1058,N_1167);
or U1213 (N_1213,N_1134,N_1186);
xnor U1214 (N_1214,N_1124,N_1079);
or U1215 (N_1215,N_1143,N_1014);
or U1216 (N_1216,N_1070,N_1178);
xor U1217 (N_1217,N_1080,N_1118);
nand U1218 (N_1218,N_1093,N_1074);
and U1219 (N_1219,N_1081,N_1110);
nand U1220 (N_1220,N_1192,N_1156);
nand U1221 (N_1221,N_1075,N_1133);
and U1222 (N_1222,N_1042,N_1140);
xnor U1223 (N_1223,N_1179,N_1153);
and U1224 (N_1224,N_1001,N_1083);
and U1225 (N_1225,N_1173,N_1164);
nand U1226 (N_1226,N_1127,N_1009);
or U1227 (N_1227,N_1177,N_1185);
and U1228 (N_1228,N_1102,N_1027);
nor U1229 (N_1229,N_1120,N_1022);
and U1230 (N_1230,N_1157,N_1098);
nand U1231 (N_1231,N_1182,N_1091);
xnor U1232 (N_1232,N_1053,N_1090);
xnor U1233 (N_1233,N_1125,N_1176);
nand U1234 (N_1234,N_1055,N_1024);
nand U1235 (N_1235,N_1130,N_1094);
and U1236 (N_1236,N_1155,N_1002);
xor U1237 (N_1237,N_1030,N_1109);
xnor U1238 (N_1238,N_1117,N_1154);
or U1239 (N_1239,N_1015,N_1142);
xor U1240 (N_1240,N_1062,N_1019);
nand U1241 (N_1241,N_1151,N_1034);
nand U1242 (N_1242,N_1113,N_1052);
and U1243 (N_1243,N_1038,N_1039);
nor U1244 (N_1244,N_1149,N_1065);
nor U1245 (N_1245,N_1037,N_1054);
nand U1246 (N_1246,N_1000,N_1112);
and U1247 (N_1247,N_1092,N_1017);
nand U1248 (N_1248,N_1181,N_1020);
nand U1249 (N_1249,N_1121,N_1132);
or U1250 (N_1250,N_1107,N_1197);
or U1251 (N_1251,N_1137,N_1006);
xor U1252 (N_1252,N_1072,N_1048);
xor U1253 (N_1253,N_1040,N_1064);
and U1254 (N_1254,N_1199,N_1077);
and U1255 (N_1255,N_1194,N_1170);
nor U1256 (N_1256,N_1016,N_1114);
and U1257 (N_1257,N_1100,N_1135);
or U1258 (N_1258,N_1097,N_1139);
nor U1259 (N_1259,N_1059,N_1032);
and U1260 (N_1260,N_1138,N_1163);
and U1261 (N_1261,N_1101,N_1018);
or U1262 (N_1262,N_1082,N_1061);
xor U1263 (N_1263,N_1086,N_1180);
nor U1264 (N_1264,N_1123,N_1115);
nand U1265 (N_1265,N_1184,N_1046);
nand U1266 (N_1266,N_1152,N_1095);
nor U1267 (N_1267,N_1172,N_1195);
and U1268 (N_1268,N_1158,N_1128);
and U1269 (N_1269,N_1169,N_1147);
nand U1270 (N_1270,N_1026,N_1193);
xnor U1271 (N_1271,N_1057,N_1111);
or U1272 (N_1272,N_1045,N_1165);
nand U1273 (N_1273,N_1198,N_1069);
nand U1274 (N_1274,N_1087,N_1196);
xnor U1275 (N_1275,N_1136,N_1078);
or U1276 (N_1276,N_1126,N_1076);
or U1277 (N_1277,N_1106,N_1104);
and U1278 (N_1278,N_1144,N_1029);
and U1279 (N_1279,N_1071,N_1047);
xnor U1280 (N_1280,N_1044,N_1063);
and U1281 (N_1281,N_1129,N_1084);
and U1282 (N_1282,N_1189,N_1008);
or U1283 (N_1283,N_1056,N_1159);
or U1284 (N_1284,N_1041,N_1148);
or U1285 (N_1285,N_1028,N_1168);
xor U1286 (N_1286,N_1005,N_1051);
and U1287 (N_1287,N_1067,N_1004);
nand U1288 (N_1288,N_1161,N_1050);
nor U1289 (N_1289,N_1088,N_1166);
nand U1290 (N_1290,N_1043,N_1141);
or U1291 (N_1291,N_1183,N_1096);
nand U1292 (N_1292,N_1021,N_1031);
or U1293 (N_1293,N_1188,N_1131);
nor U1294 (N_1294,N_1025,N_1145);
xnor U1295 (N_1295,N_1003,N_1119);
or U1296 (N_1296,N_1103,N_1150);
or U1297 (N_1297,N_1175,N_1122);
nand U1298 (N_1298,N_1011,N_1116);
nand U1299 (N_1299,N_1191,N_1174);
or U1300 (N_1300,N_1051,N_1172);
nand U1301 (N_1301,N_1060,N_1070);
or U1302 (N_1302,N_1062,N_1076);
or U1303 (N_1303,N_1053,N_1167);
nand U1304 (N_1304,N_1186,N_1167);
xnor U1305 (N_1305,N_1067,N_1015);
nor U1306 (N_1306,N_1062,N_1058);
and U1307 (N_1307,N_1047,N_1178);
xnor U1308 (N_1308,N_1191,N_1002);
or U1309 (N_1309,N_1012,N_1115);
or U1310 (N_1310,N_1065,N_1098);
nor U1311 (N_1311,N_1062,N_1038);
and U1312 (N_1312,N_1178,N_1129);
nor U1313 (N_1313,N_1030,N_1191);
or U1314 (N_1314,N_1064,N_1123);
nand U1315 (N_1315,N_1066,N_1018);
nor U1316 (N_1316,N_1054,N_1077);
nand U1317 (N_1317,N_1135,N_1080);
nor U1318 (N_1318,N_1098,N_1061);
nor U1319 (N_1319,N_1086,N_1155);
xnor U1320 (N_1320,N_1180,N_1112);
xor U1321 (N_1321,N_1054,N_1047);
nor U1322 (N_1322,N_1036,N_1007);
nand U1323 (N_1323,N_1002,N_1121);
xor U1324 (N_1324,N_1113,N_1070);
nor U1325 (N_1325,N_1089,N_1055);
nand U1326 (N_1326,N_1070,N_1076);
nand U1327 (N_1327,N_1040,N_1156);
or U1328 (N_1328,N_1025,N_1166);
nand U1329 (N_1329,N_1059,N_1124);
and U1330 (N_1330,N_1081,N_1099);
nand U1331 (N_1331,N_1046,N_1130);
or U1332 (N_1332,N_1170,N_1027);
nor U1333 (N_1333,N_1028,N_1139);
nand U1334 (N_1334,N_1168,N_1063);
nor U1335 (N_1335,N_1128,N_1166);
nand U1336 (N_1336,N_1012,N_1069);
or U1337 (N_1337,N_1013,N_1003);
and U1338 (N_1338,N_1070,N_1119);
and U1339 (N_1339,N_1004,N_1044);
nand U1340 (N_1340,N_1124,N_1137);
nand U1341 (N_1341,N_1007,N_1090);
and U1342 (N_1342,N_1099,N_1111);
xor U1343 (N_1343,N_1122,N_1144);
xor U1344 (N_1344,N_1136,N_1108);
nor U1345 (N_1345,N_1155,N_1000);
xor U1346 (N_1346,N_1110,N_1050);
or U1347 (N_1347,N_1066,N_1140);
nand U1348 (N_1348,N_1175,N_1133);
or U1349 (N_1349,N_1090,N_1129);
or U1350 (N_1350,N_1120,N_1168);
nor U1351 (N_1351,N_1019,N_1113);
nor U1352 (N_1352,N_1093,N_1071);
nor U1353 (N_1353,N_1142,N_1086);
xor U1354 (N_1354,N_1083,N_1039);
nand U1355 (N_1355,N_1127,N_1077);
nand U1356 (N_1356,N_1190,N_1122);
nand U1357 (N_1357,N_1175,N_1072);
and U1358 (N_1358,N_1073,N_1174);
nor U1359 (N_1359,N_1151,N_1007);
and U1360 (N_1360,N_1022,N_1145);
nand U1361 (N_1361,N_1026,N_1179);
or U1362 (N_1362,N_1122,N_1096);
and U1363 (N_1363,N_1182,N_1044);
nand U1364 (N_1364,N_1129,N_1108);
xor U1365 (N_1365,N_1001,N_1077);
and U1366 (N_1366,N_1104,N_1164);
xnor U1367 (N_1367,N_1183,N_1027);
nor U1368 (N_1368,N_1082,N_1189);
nand U1369 (N_1369,N_1090,N_1118);
and U1370 (N_1370,N_1038,N_1150);
nor U1371 (N_1371,N_1165,N_1070);
nand U1372 (N_1372,N_1127,N_1070);
xnor U1373 (N_1373,N_1072,N_1013);
nor U1374 (N_1374,N_1102,N_1056);
nor U1375 (N_1375,N_1154,N_1162);
and U1376 (N_1376,N_1003,N_1075);
nand U1377 (N_1377,N_1066,N_1138);
nand U1378 (N_1378,N_1043,N_1155);
nand U1379 (N_1379,N_1147,N_1040);
or U1380 (N_1380,N_1100,N_1050);
or U1381 (N_1381,N_1105,N_1164);
nand U1382 (N_1382,N_1091,N_1002);
and U1383 (N_1383,N_1022,N_1109);
or U1384 (N_1384,N_1025,N_1198);
or U1385 (N_1385,N_1046,N_1054);
and U1386 (N_1386,N_1113,N_1152);
xor U1387 (N_1387,N_1194,N_1049);
xor U1388 (N_1388,N_1140,N_1151);
nand U1389 (N_1389,N_1052,N_1098);
nor U1390 (N_1390,N_1131,N_1055);
nand U1391 (N_1391,N_1194,N_1089);
xor U1392 (N_1392,N_1120,N_1078);
and U1393 (N_1393,N_1009,N_1177);
nand U1394 (N_1394,N_1069,N_1160);
nand U1395 (N_1395,N_1186,N_1073);
or U1396 (N_1396,N_1047,N_1044);
and U1397 (N_1397,N_1183,N_1131);
xnor U1398 (N_1398,N_1101,N_1147);
or U1399 (N_1399,N_1051,N_1095);
nor U1400 (N_1400,N_1320,N_1325);
nand U1401 (N_1401,N_1226,N_1259);
nand U1402 (N_1402,N_1204,N_1352);
and U1403 (N_1403,N_1236,N_1215);
xnor U1404 (N_1404,N_1266,N_1237);
nand U1405 (N_1405,N_1323,N_1265);
nand U1406 (N_1406,N_1216,N_1290);
nand U1407 (N_1407,N_1356,N_1208);
nor U1408 (N_1408,N_1328,N_1337);
nand U1409 (N_1409,N_1366,N_1277);
xnor U1410 (N_1410,N_1217,N_1304);
xnor U1411 (N_1411,N_1264,N_1317);
nand U1412 (N_1412,N_1293,N_1294);
nand U1413 (N_1413,N_1345,N_1244);
or U1414 (N_1414,N_1256,N_1297);
and U1415 (N_1415,N_1349,N_1371);
nor U1416 (N_1416,N_1348,N_1380);
xor U1417 (N_1417,N_1276,N_1260);
xnor U1418 (N_1418,N_1246,N_1372);
and U1419 (N_1419,N_1258,N_1285);
nor U1420 (N_1420,N_1339,N_1335);
xnor U1421 (N_1421,N_1239,N_1238);
nor U1422 (N_1422,N_1281,N_1207);
and U1423 (N_1423,N_1212,N_1309);
nor U1424 (N_1424,N_1318,N_1291);
and U1425 (N_1425,N_1223,N_1347);
or U1426 (N_1426,N_1200,N_1338);
nor U1427 (N_1427,N_1311,N_1295);
and U1428 (N_1428,N_1301,N_1334);
nor U1429 (N_1429,N_1283,N_1298);
nand U1430 (N_1430,N_1343,N_1365);
nor U1431 (N_1431,N_1396,N_1395);
xnor U1432 (N_1432,N_1274,N_1279);
xnor U1433 (N_1433,N_1242,N_1201);
xnor U1434 (N_1434,N_1303,N_1327);
nor U1435 (N_1435,N_1230,N_1233);
nor U1436 (N_1436,N_1261,N_1252);
or U1437 (N_1437,N_1210,N_1333);
or U1438 (N_1438,N_1227,N_1245);
nand U1439 (N_1439,N_1219,N_1286);
and U1440 (N_1440,N_1341,N_1322);
or U1441 (N_1441,N_1267,N_1386);
or U1442 (N_1442,N_1313,N_1379);
nor U1443 (N_1443,N_1344,N_1271);
or U1444 (N_1444,N_1273,N_1397);
and U1445 (N_1445,N_1319,N_1247);
and U1446 (N_1446,N_1361,N_1257);
nor U1447 (N_1447,N_1287,N_1292);
or U1448 (N_1448,N_1213,N_1316);
and U1449 (N_1449,N_1367,N_1332);
nand U1450 (N_1450,N_1382,N_1384);
nor U1451 (N_1451,N_1373,N_1222);
nor U1452 (N_1452,N_1314,N_1221);
nand U1453 (N_1453,N_1374,N_1275);
and U1454 (N_1454,N_1306,N_1398);
xnor U1455 (N_1455,N_1268,N_1358);
nor U1456 (N_1456,N_1302,N_1235);
nand U1457 (N_1457,N_1305,N_1224);
and U1458 (N_1458,N_1342,N_1378);
nor U1459 (N_1459,N_1326,N_1255);
nand U1460 (N_1460,N_1299,N_1350);
xnor U1461 (N_1461,N_1262,N_1312);
nor U1462 (N_1462,N_1394,N_1288);
nand U1463 (N_1463,N_1228,N_1354);
nor U1464 (N_1464,N_1392,N_1389);
xor U1465 (N_1465,N_1240,N_1351);
nor U1466 (N_1466,N_1383,N_1203);
nand U1467 (N_1467,N_1241,N_1270);
xnor U1468 (N_1468,N_1315,N_1360);
xor U1469 (N_1469,N_1346,N_1330);
xnor U1470 (N_1470,N_1218,N_1214);
or U1471 (N_1471,N_1385,N_1355);
or U1472 (N_1472,N_1376,N_1307);
or U1473 (N_1473,N_1243,N_1272);
or U1474 (N_1474,N_1377,N_1282);
xor U1475 (N_1475,N_1364,N_1399);
or U1476 (N_1476,N_1284,N_1369);
and U1477 (N_1477,N_1253,N_1340);
xor U1478 (N_1478,N_1251,N_1363);
nor U1479 (N_1479,N_1388,N_1232);
or U1480 (N_1480,N_1336,N_1205);
xor U1481 (N_1481,N_1300,N_1368);
and U1482 (N_1482,N_1324,N_1250);
nor U1483 (N_1483,N_1202,N_1278);
xnor U1484 (N_1484,N_1225,N_1362);
nor U1485 (N_1485,N_1375,N_1248);
nand U1486 (N_1486,N_1211,N_1370);
nand U1487 (N_1487,N_1359,N_1331);
nor U1488 (N_1488,N_1289,N_1254);
or U1489 (N_1489,N_1209,N_1329);
xnor U1490 (N_1490,N_1220,N_1381);
xnor U1491 (N_1491,N_1357,N_1231);
or U1492 (N_1492,N_1310,N_1391);
or U1493 (N_1493,N_1387,N_1308);
or U1494 (N_1494,N_1280,N_1321);
nand U1495 (N_1495,N_1353,N_1263);
or U1496 (N_1496,N_1229,N_1269);
xnor U1497 (N_1497,N_1249,N_1234);
nor U1498 (N_1498,N_1393,N_1390);
nor U1499 (N_1499,N_1296,N_1206);
nor U1500 (N_1500,N_1207,N_1309);
xor U1501 (N_1501,N_1216,N_1331);
nor U1502 (N_1502,N_1304,N_1358);
or U1503 (N_1503,N_1344,N_1233);
nand U1504 (N_1504,N_1207,N_1223);
nor U1505 (N_1505,N_1337,N_1286);
or U1506 (N_1506,N_1212,N_1342);
nand U1507 (N_1507,N_1396,N_1211);
or U1508 (N_1508,N_1341,N_1308);
and U1509 (N_1509,N_1288,N_1319);
and U1510 (N_1510,N_1270,N_1398);
nor U1511 (N_1511,N_1312,N_1353);
and U1512 (N_1512,N_1399,N_1307);
or U1513 (N_1513,N_1361,N_1210);
and U1514 (N_1514,N_1225,N_1353);
nor U1515 (N_1515,N_1355,N_1254);
nor U1516 (N_1516,N_1243,N_1205);
and U1517 (N_1517,N_1226,N_1367);
and U1518 (N_1518,N_1359,N_1368);
xnor U1519 (N_1519,N_1246,N_1310);
nor U1520 (N_1520,N_1350,N_1336);
nor U1521 (N_1521,N_1235,N_1237);
or U1522 (N_1522,N_1359,N_1272);
nor U1523 (N_1523,N_1342,N_1332);
nand U1524 (N_1524,N_1385,N_1263);
and U1525 (N_1525,N_1321,N_1356);
and U1526 (N_1526,N_1282,N_1314);
nand U1527 (N_1527,N_1291,N_1362);
nor U1528 (N_1528,N_1284,N_1233);
nor U1529 (N_1529,N_1246,N_1315);
nand U1530 (N_1530,N_1255,N_1329);
nor U1531 (N_1531,N_1336,N_1297);
xor U1532 (N_1532,N_1351,N_1395);
xnor U1533 (N_1533,N_1293,N_1356);
and U1534 (N_1534,N_1368,N_1229);
or U1535 (N_1535,N_1303,N_1246);
or U1536 (N_1536,N_1288,N_1275);
xnor U1537 (N_1537,N_1370,N_1364);
or U1538 (N_1538,N_1369,N_1252);
or U1539 (N_1539,N_1356,N_1310);
and U1540 (N_1540,N_1366,N_1356);
nand U1541 (N_1541,N_1225,N_1219);
nor U1542 (N_1542,N_1267,N_1224);
and U1543 (N_1543,N_1327,N_1343);
and U1544 (N_1544,N_1229,N_1304);
nand U1545 (N_1545,N_1319,N_1223);
or U1546 (N_1546,N_1243,N_1297);
or U1547 (N_1547,N_1346,N_1389);
nor U1548 (N_1548,N_1236,N_1279);
nand U1549 (N_1549,N_1309,N_1238);
xnor U1550 (N_1550,N_1387,N_1212);
and U1551 (N_1551,N_1352,N_1260);
and U1552 (N_1552,N_1217,N_1278);
xnor U1553 (N_1553,N_1395,N_1347);
or U1554 (N_1554,N_1296,N_1240);
nand U1555 (N_1555,N_1372,N_1350);
nor U1556 (N_1556,N_1310,N_1215);
nor U1557 (N_1557,N_1391,N_1337);
and U1558 (N_1558,N_1344,N_1238);
and U1559 (N_1559,N_1392,N_1371);
and U1560 (N_1560,N_1339,N_1246);
or U1561 (N_1561,N_1240,N_1389);
nand U1562 (N_1562,N_1352,N_1289);
or U1563 (N_1563,N_1238,N_1207);
nand U1564 (N_1564,N_1219,N_1252);
nand U1565 (N_1565,N_1233,N_1220);
xnor U1566 (N_1566,N_1298,N_1252);
xnor U1567 (N_1567,N_1212,N_1294);
or U1568 (N_1568,N_1383,N_1238);
nand U1569 (N_1569,N_1234,N_1237);
and U1570 (N_1570,N_1372,N_1308);
nor U1571 (N_1571,N_1389,N_1306);
or U1572 (N_1572,N_1324,N_1302);
and U1573 (N_1573,N_1381,N_1378);
nor U1574 (N_1574,N_1380,N_1345);
or U1575 (N_1575,N_1394,N_1267);
nand U1576 (N_1576,N_1343,N_1295);
or U1577 (N_1577,N_1216,N_1345);
xor U1578 (N_1578,N_1310,N_1295);
or U1579 (N_1579,N_1209,N_1255);
and U1580 (N_1580,N_1316,N_1308);
xnor U1581 (N_1581,N_1304,N_1227);
nand U1582 (N_1582,N_1259,N_1212);
nor U1583 (N_1583,N_1332,N_1226);
and U1584 (N_1584,N_1279,N_1235);
or U1585 (N_1585,N_1365,N_1288);
nand U1586 (N_1586,N_1250,N_1330);
or U1587 (N_1587,N_1348,N_1212);
or U1588 (N_1588,N_1242,N_1321);
and U1589 (N_1589,N_1297,N_1264);
and U1590 (N_1590,N_1341,N_1216);
and U1591 (N_1591,N_1227,N_1320);
xnor U1592 (N_1592,N_1234,N_1340);
or U1593 (N_1593,N_1250,N_1288);
or U1594 (N_1594,N_1319,N_1364);
xor U1595 (N_1595,N_1232,N_1377);
or U1596 (N_1596,N_1298,N_1216);
nand U1597 (N_1597,N_1325,N_1308);
xnor U1598 (N_1598,N_1204,N_1319);
or U1599 (N_1599,N_1224,N_1315);
and U1600 (N_1600,N_1524,N_1508);
nor U1601 (N_1601,N_1589,N_1463);
nor U1602 (N_1602,N_1569,N_1473);
nor U1603 (N_1603,N_1467,N_1594);
nand U1604 (N_1604,N_1492,N_1411);
or U1605 (N_1605,N_1424,N_1442);
and U1606 (N_1606,N_1468,N_1481);
and U1607 (N_1607,N_1507,N_1578);
nor U1608 (N_1608,N_1584,N_1572);
and U1609 (N_1609,N_1576,N_1443);
nand U1610 (N_1610,N_1489,N_1546);
xnor U1611 (N_1611,N_1414,N_1509);
xor U1612 (N_1612,N_1462,N_1552);
xor U1613 (N_1613,N_1593,N_1420);
xor U1614 (N_1614,N_1458,N_1567);
or U1615 (N_1615,N_1441,N_1598);
or U1616 (N_1616,N_1418,N_1556);
nor U1617 (N_1617,N_1547,N_1581);
xor U1618 (N_1618,N_1499,N_1599);
nand U1619 (N_1619,N_1422,N_1521);
and U1620 (N_1620,N_1526,N_1446);
nor U1621 (N_1621,N_1416,N_1579);
nand U1622 (N_1622,N_1533,N_1440);
or U1623 (N_1623,N_1563,N_1503);
or U1624 (N_1624,N_1565,N_1511);
and U1625 (N_1625,N_1548,N_1537);
or U1626 (N_1626,N_1403,N_1482);
or U1627 (N_1627,N_1591,N_1469);
or U1628 (N_1628,N_1493,N_1496);
and U1629 (N_1629,N_1459,N_1423);
and U1630 (N_1630,N_1497,N_1592);
nor U1631 (N_1631,N_1501,N_1505);
nor U1632 (N_1632,N_1412,N_1532);
xnor U1633 (N_1633,N_1425,N_1417);
nand U1634 (N_1634,N_1530,N_1439);
xor U1635 (N_1635,N_1456,N_1510);
and U1636 (N_1636,N_1564,N_1574);
nor U1637 (N_1637,N_1434,N_1485);
xnor U1638 (N_1638,N_1553,N_1504);
or U1639 (N_1639,N_1568,N_1519);
and U1640 (N_1640,N_1419,N_1520);
and U1641 (N_1641,N_1555,N_1477);
xor U1642 (N_1642,N_1597,N_1494);
xnor U1643 (N_1643,N_1402,N_1538);
and U1644 (N_1644,N_1498,N_1429);
xnor U1645 (N_1645,N_1539,N_1449);
nor U1646 (N_1646,N_1483,N_1409);
and U1647 (N_1647,N_1536,N_1476);
nor U1648 (N_1648,N_1438,N_1466);
nand U1649 (N_1649,N_1545,N_1580);
nor U1650 (N_1650,N_1444,N_1406);
and U1651 (N_1651,N_1488,N_1528);
xnor U1652 (N_1652,N_1535,N_1415);
nor U1653 (N_1653,N_1437,N_1518);
xor U1654 (N_1654,N_1551,N_1454);
or U1655 (N_1655,N_1460,N_1490);
nor U1656 (N_1656,N_1514,N_1487);
or U1657 (N_1657,N_1575,N_1453);
or U1658 (N_1658,N_1582,N_1465);
and U1659 (N_1659,N_1527,N_1522);
nor U1660 (N_1660,N_1502,N_1404);
or U1661 (N_1661,N_1495,N_1472);
xor U1662 (N_1662,N_1554,N_1405);
and U1663 (N_1663,N_1428,N_1450);
nand U1664 (N_1664,N_1525,N_1471);
nand U1665 (N_1665,N_1596,N_1408);
nand U1666 (N_1666,N_1474,N_1431);
nand U1667 (N_1667,N_1541,N_1515);
xor U1668 (N_1668,N_1531,N_1430);
nand U1669 (N_1669,N_1475,N_1513);
and U1670 (N_1670,N_1585,N_1523);
nor U1671 (N_1671,N_1590,N_1587);
nand U1672 (N_1672,N_1583,N_1562);
or U1673 (N_1673,N_1421,N_1506);
and U1674 (N_1674,N_1480,N_1451);
or U1675 (N_1675,N_1571,N_1543);
and U1676 (N_1676,N_1512,N_1550);
nor U1677 (N_1677,N_1500,N_1577);
and U1678 (N_1678,N_1557,N_1560);
nor U1679 (N_1679,N_1549,N_1479);
nand U1680 (N_1680,N_1401,N_1413);
nor U1681 (N_1681,N_1595,N_1461);
or U1682 (N_1682,N_1486,N_1432);
xor U1683 (N_1683,N_1534,N_1457);
or U1684 (N_1684,N_1407,N_1447);
or U1685 (N_1685,N_1464,N_1570);
xor U1686 (N_1686,N_1445,N_1561);
nand U1687 (N_1687,N_1478,N_1540);
and U1688 (N_1688,N_1544,N_1573);
and U1689 (N_1689,N_1470,N_1433);
nand U1690 (N_1690,N_1517,N_1588);
nor U1691 (N_1691,N_1566,N_1435);
xor U1692 (N_1692,N_1529,N_1426);
or U1693 (N_1693,N_1448,N_1452);
and U1694 (N_1694,N_1400,N_1558);
nor U1695 (N_1695,N_1410,N_1586);
xor U1696 (N_1696,N_1491,N_1542);
xnor U1697 (N_1697,N_1455,N_1559);
or U1698 (N_1698,N_1427,N_1516);
nand U1699 (N_1699,N_1484,N_1436);
nor U1700 (N_1700,N_1426,N_1486);
and U1701 (N_1701,N_1583,N_1528);
nor U1702 (N_1702,N_1530,N_1575);
and U1703 (N_1703,N_1515,N_1466);
nand U1704 (N_1704,N_1572,N_1437);
nand U1705 (N_1705,N_1461,N_1418);
and U1706 (N_1706,N_1421,N_1569);
or U1707 (N_1707,N_1575,N_1515);
nand U1708 (N_1708,N_1480,N_1413);
xnor U1709 (N_1709,N_1472,N_1449);
nand U1710 (N_1710,N_1421,N_1505);
xor U1711 (N_1711,N_1511,N_1448);
nand U1712 (N_1712,N_1575,N_1525);
nand U1713 (N_1713,N_1590,N_1435);
xnor U1714 (N_1714,N_1539,N_1427);
xor U1715 (N_1715,N_1539,N_1473);
or U1716 (N_1716,N_1562,N_1496);
nand U1717 (N_1717,N_1516,N_1557);
nor U1718 (N_1718,N_1409,N_1494);
xor U1719 (N_1719,N_1414,N_1468);
nand U1720 (N_1720,N_1505,N_1529);
xnor U1721 (N_1721,N_1460,N_1402);
and U1722 (N_1722,N_1455,N_1454);
nand U1723 (N_1723,N_1410,N_1411);
or U1724 (N_1724,N_1537,N_1415);
nand U1725 (N_1725,N_1503,N_1406);
xnor U1726 (N_1726,N_1437,N_1423);
xor U1727 (N_1727,N_1431,N_1453);
nand U1728 (N_1728,N_1594,N_1562);
and U1729 (N_1729,N_1439,N_1440);
nand U1730 (N_1730,N_1542,N_1583);
nor U1731 (N_1731,N_1569,N_1568);
and U1732 (N_1732,N_1497,N_1577);
xnor U1733 (N_1733,N_1572,N_1593);
or U1734 (N_1734,N_1530,N_1533);
nand U1735 (N_1735,N_1558,N_1522);
xnor U1736 (N_1736,N_1545,N_1412);
nor U1737 (N_1737,N_1556,N_1516);
and U1738 (N_1738,N_1561,N_1529);
nand U1739 (N_1739,N_1437,N_1461);
or U1740 (N_1740,N_1584,N_1445);
nand U1741 (N_1741,N_1447,N_1455);
nand U1742 (N_1742,N_1494,N_1467);
and U1743 (N_1743,N_1415,N_1409);
xor U1744 (N_1744,N_1403,N_1427);
nand U1745 (N_1745,N_1455,N_1593);
nand U1746 (N_1746,N_1415,N_1479);
nor U1747 (N_1747,N_1533,N_1596);
nand U1748 (N_1748,N_1498,N_1575);
nand U1749 (N_1749,N_1522,N_1447);
nand U1750 (N_1750,N_1593,N_1556);
nand U1751 (N_1751,N_1580,N_1583);
xnor U1752 (N_1752,N_1569,N_1482);
and U1753 (N_1753,N_1564,N_1515);
nand U1754 (N_1754,N_1593,N_1445);
nor U1755 (N_1755,N_1524,N_1463);
nor U1756 (N_1756,N_1466,N_1480);
nor U1757 (N_1757,N_1590,N_1499);
nor U1758 (N_1758,N_1409,N_1580);
nor U1759 (N_1759,N_1509,N_1592);
xnor U1760 (N_1760,N_1502,N_1535);
nor U1761 (N_1761,N_1541,N_1522);
and U1762 (N_1762,N_1463,N_1585);
and U1763 (N_1763,N_1507,N_1493);
xor U1764 (N_1764,N_1453,N_1580);
or U1765 (N_1765,N_1519,N_1587);
nor U1766 (N_1766,N_1484,N_1587);
and U1767 (N_1767,N_1533,N_1416);
nor U1768 (N_1768,N_1426,N_1571);
xor U1769 (N_1769,N_1547,N_1421);
nand U1770 (N_1770,N_1506,N_1554);
and U1771 (N_1771,N_1433,N_1429);
or U1772 (N_1772,N_1470,N_1444);
or U1773 (N_1773,N_1419,N_1513);
and U1774 (N_1774,N_1424,N_1501);
or U1775 (N_1775,N_1469,N_1545);
nand U1776 (N_1776,N_1568,N_1586);
xor U1777 (N_1777,N_1444,N_1590);
and U1778 (N_1778,N_1473,N_1545);
and U1779 (N_1779,N_1520,N_1568);
nor U1780 (N_1780,N_1578,N_1430);
and U1781 (N_1781,N_1465,N_1541);
nor U1782 (N_1782,N_1568,N_1532);
nor U1783 (N_1783,N_1566,N_1551);
nand U1784 (N_1784,N_1519,N_1494);
or U1785 (N_1785,N_1449,N_1550);
nand U1786 (N_1786,N_1491,N_1595);
nor U1787 (N_1787,N_1495,N_1505);
xnor U1788 (N_1788,N_1515,N_1441);
or U1789 (N_1789,N_1402,N_1544);
xnor U1790 (N_1790,N_1400,N_1478);
nor U1791 (N_1791,N_1592,N_1559);
nand U1792 (N_1792,N_1460,N_1583);
or U1793 (N_1793,N_1400,N_1406);
nand U1794 (N_1794,N_1553,N_1593);
nor U1795 (N_1795,N_1489,N_1575);
or U1796 (N_1796,N_1543,N_1482);
and U1797 (N_1797,N_1540,N_1564);
nor U1798 (N_1798,N_1405,N_1546);
or U1799 (N_1799,N_1525,N_1445);
nand U1800 (N_1800,N_1669,N_1733);
or U1801 (N_1801,N_1694,N_1725);
nand U1802 (N_1802,N_1646,N_1663);
and U1803 (N_1803,N_1657,N_1609);
xor U1804 (N_1804,N_1616,N_1712);
or U1805 (N_1805,N_1651,N_1781);
nand U1806 (N_1806,N_1772,N_1673);
and U1807 (N_1807,N_1726,N_1763);
nor U1808 (N_1808,N_1792,N_1610);
nor U1809 (N_1809,N_1723,N_1751);
nor U1810 (N_1810,N_1688,N_1630);
and U1811 (N_1811,N_1777,N_1639);
and U1812 (N_1812,N_1691,N_1615);
nand U1813 (N_1813,N_1698,N_1714);
or U1814 (N_1814,N_1721,N_1677);
nor U1815 (N_1815,N_1658,N_1749);
or U1816 (N_1816,N_1748,N_1703);
nor U1817 (N_1817,N_1685,N_1624);
xor U1818 (N_1818,N_1793,N_1641);
or U1819 (N_1819,N_1640,N_1617);
or U1820 (N_1820,N_1774,N_1668);
xnor U1821 (N_1821,N_1730,N_1759);
and U1822 (N_1822,N_1627,N_1728);
and U1823 (N_1823,N_1702,N_1742);
and U1824 (N_1824,N_1700,N_1783);
nand U1825 (N_1825,N_1608,N_1690);
xor U1826 (N_1826,N_1791,N_1765);
and U1827 (N_1827,N_1718,N_1746);
or U1828 (N_1828,N_1629,N_1631);
nor U1829 (N_1829,N_1788,N_1604);
nor U1830 (N_1830,N_1671,N_1734);
xnor U1831 (N_1831,N_1649,N_1655);
or U1832 (N_1832,N_1750,N_1789);
and U1833 (N_1833,N_1761,N_1705);
xor U1834 (N_1834,N_1612,N_1686);
and U1835 (N_1835,N_1695,N_1745);
or U1836 (N_1836,N_1707,N_1650);
nor U1837 (N_1837,N_1626,N_1618);
or U1838 (N_1838,N_1779,N_1764);
and U1839 (N_1839,N_1758,N_1635);
or U1840 (N_1840,N_1778,N_1744);
and U1841 (N_1841,N_1797,N_1656);
and U1842 (N_1842,N_1760,N_1741);
xor U1843 (N_1843,N_1672,N_1636);
xnor U1844 (N_1844,N_1770,N_1667);
xor U1845 (N_1845,N_1664,N_1790);
nor U1846 (N_1846,N_1699,N_1637);
nand U1847 (N_1847,N_1753,N_1676);
nor U1848 (N_1848,N_1755,N_1687);
xor U1849 (N_1849,N_1785,N_1743);
and U1850 (N_1850,N_1738,N_1642);
and U1851 (N_1851,N_1711,N_1796);
nor U1852 (N_1852,N_1740,N_1737);
nor U1853 (N_1853,N_1645,N_1697);
nand U1854 (N_1854,N_1621,N_1784);
and U1855 (N_1855,N_1766,N_1706);
nand U1856 (N_1856,N_1782,N_1692);
nor U1857 (N_1857,N_1653,N_1652);
nand U1858 (N_1858,N_1601,N_1681);
nor U1859 (N_1859,N_1775,N_1622);
nand U1860 (N_1860,N_1701,N_1732);
or U1861 (N_1861,N_1666,N_1607);
nor U1862 (N_1862,N_1623,N_1715);
or U1863 (N_1863,N_1661,N_1717);
or U1864 (N_1864,N_1754,N_1654);
and U1865 (N_1865,N_1606,N_1680);
and U1866 (N_1866,N_1768,N_1620);
nand U1867 (N_1867,N_1710,N_1719);
or U1868 (N_1868,N_1716,N_1739);
and U1869 (N_1869,N_1795,N_1709);
or U1870 (N_1870,N_1780,N_1633);
and U1871 (N_1871,N_1648,N_1794);
xor U1872 (N_1872,N_1665,N_1693);
nor U1873 (N_1873,N_1659,N_1638);
and U1874 (N_1874,N_1647,N_1786);
or U1875 (N_1875,N_1600,N_1762);
and U1876 (N_1876,N_1660,N_1683);
nand U1877 (N_1877,N_1776,N_1720);
xnor U1878 (N_1878,N_1613,N_1603);
or U1879 (N_1879,N_1625,N_1736);
nor U1880 (N_1880,N_1769,N_1787);
nor U1881 (N_1881,N_1704,N_1674);
and U1882 (N_1882,N_1735,N_1628);
or U1883 (N_1883,N_1708,N_1722);
xor U1884 (N_1884,N_1643,N_1713);
xnor U1885 (N_1885,N_1682,N_1644);
xnor U1886 (N_1886,N_1670,N_1619);
xnor U1887 (N_1887,N_1724,N_1731);
nand U1888 (N_1888,N_1747,N_1773);
and U1889 (N_1889,N_1602,N_1771);
xnor U1890 (N_1890,N_1675,N_1679);
nand U1891 (N_1891,N_1799,N_1696);
nor U1892 (N_1892,N_1757,N_1611);
nor U1893 (N_1893,N_1767,N_1689);
or U1894 (N_1894,N_1798,N_1678);
and U1895 (N_1895,N_1729,N_1605);
nor U1896 (N_1896,N_1634,N_1727);
nor U1897 (N_1897,N_1662,N_1614);
or U1898 (N_1898,N_1752,N_1632);
and U1899 (N_1899,N_1756,N_1684);
or U1900 (N_1900,N_1781,N_1687);
and U1901 (N_1901,N_1772,N_1779);
or U1902 (N_1902,N_1796,N_1788);
or U1903 (N_1903,N_1692,N_1718);
nand U1904 (N_1904,N_1723,N_1757);
nor U1905 (N_1905,N_1703,N_1650);
nand U1906 (N_1906,N_1684,N_1691);
xnor U1907 (N_1907,N_1658,N_1676);
and U1908 (N_1908,N_1621,N_1795);
nand U1909 (N_1909,N_1694,N_1615);
nand U1910 (N_1910,N_1620,N_1660);
nor U1911 (N_1911,N_1672,N_1611);
nand U1912 (N_1912,N_1683,N_1709);
or U1913 (N_1913,N_1792,N_1661);
nor U1914 (N_1914,N_1729,N_1745);
nand U1915 (N_1915,N_1764,N_1667);
or U1916 (N_1916,N_1694,N_1733);
xnor U1917 (N_1917,N_1783,N_1735);
and U1918 (N_1918,N_1783,N_1776);
nand U1919 (N_1919,N_1657,N_1762);
xor U1920 (N_1920,N_1744,N_1693);
xnor U1921 (N_1921,N_1762,N_1658);
and U1922 (N_1922,N_1701,N_1697);
and U1923 (N_1923,N_1658,N_1779);
nand U1924 (N_1924,N_1714,N_1777);
or U1925 (N_1925,N_1779,N_1744);
nand U1926 (N_1926,N_1790,N_1778);
or U1927 (N_1927,N_1785,N_1637);
xor U1928 (N_1928,N_1732,N_1753);
and U1929 (N_1929,N_1728,N_1600);
nand U1930 (N_1930,N_1778,N_1751);
and U1931 (N_1931,N_1702,N_1737);
xnor U1932 (N_1932,N_1647,N_1672);
or U1933 (N_1933,N_1731,N_1652);
and U1934 (N_1934,N_1673,N_1675);
xor U1935 (N_1935,N_1756,N_1717);
or U1936 (N_1936,N_1726,N_1790);
and U1937 (N_1937,N_1791,N_1714);
nor U1938 (N_1938,N_1659,N_1713);
xnor U1939 (N_1939,N_1644,N_1730);
nand U1940 (N_1940,N_1622,N_1617);
or U1941 (N_1941,N_1677,N_1764);
xnor U1942 (N_1942,N_1631,N_1647);
nor U1943 (N_1943,N_1671,N_1670);
xor U1944 (N_1944,N_1713,N_1702);
xnor U1945 (N_1945,N_1792,N_1603);
xor U1946 (N_1946,N_1612,N_1712);
nand U1947 (N_1947,N_1739,N_1656);
nand U1948 (N_1948,N_1740,N_1608);
nor U1949 (N_1949,N_1615,N_1637);
and U1950 (N_1950,N_1675,N_1665);
and U1951 (N_1951,N_1656,N_1669);
xnor U1952 (N_1952,N_1779,N_1706);
nand U1953 (N_1953,N_1774,N_1747);
or U1954 (N_1954,N_1711,N_1764);
and U1955 (N_1955,N_1664,N_1782);
xnor U1956 (N_1956,N_1626,N_1658);
xor U1957 (N_1957,N_1675,N_1775);
nor U1958 (N_1958,N_1794,N_1663);
or U1959 (N_1959,N_1618,N_1686);
or U1960 (N_1960,N_1708,N_1768);
nor U1961 (N_1961,N_1613,N_1690);
or U1962 (N_1962,N_1621,N_1625);
or U1963 (N_1963,N_1793,N_1687);
or U1964 (N_1964,N_1627,N_1776);
xnor U1965 (N_1965,N_1786,N_1666);
nor U1966 (N_1966,N_1771,N_1706);
xnor U1967 (N_1967,N_1741,N_1644);
xnor U1968 (N_1968,N_1768,N_1653);
nand U1969 (N_1969,N_1727,N_1601);
nor U1970 (N_1970,N_1725,N_1635);
and U1971 (N_1971,N_1619,N_1798);
nand U1972 (N_1972,N_1614,N_1772);
nor U1973 (N_1973,N_1728,N_1658);
and U1974 (N_1974,N_1651,N_1744);
xor U1975 (N_1975,N_1609,N_1709);
and U1976 (N_1976,N_1769,N_1611);
or U1977 (N_1977,N_1719,N_1677);
nor U1978 (N_1978,N_1637,N_1697);
nand U1979 (N_1979,N_1670,N_1722);
or U1980 (N_1980,N_1643,N_1665);
nand U1981 (N_1981,N_1769,N_1731);
and U1982 (N_1982,N_1602,N_1704);
or U1983 (N_1983,N_1607,N_1679);
nor U1984 (N_1984,N_1628,N_1699);
or U1985 (N_1985,N_1734,N_1668);
xor U1986 (N_1986,N_1718,N_1638);
xnor U1987 (N_1987,N_1722,N_1620);
xnor U1988 (N_1988,N_1760,N_1613);
xnor U1989 (N_1989,N_1721,N_1609);
xor U1990 (N_1990,N_1733,N_1716);
or U1991 (N_1991,N_1651,N_1791);
or U1992 (N_1992,N_1690,N_1705);
xor U1993 (N_1993,N_1633,N_1785);
nor U1994 (N_1994,N_1771,N_1786);
nand U1995 (N_1995,N_1719,N_1727);
xnor U1996 (N_1996,N_1734,N_1771);
xor U1997 (N_1997,N_1617,N_1758);
xnor U1998 (N_1998,N_1790,N_1639);
and U1999 (N_1999,N_1731,N_1743);
or U2000 (N_2000,N_1996,N_1891);
xor U2001 (N_2001,N_1813,N_1976);
or U2002 (N_2002,N_1984,N_1854);
and U2003 (N_2003,N_1929,N_1972);
nand U2004 (N_2004,N_1889,N_1806);
and U2005 (N_2005,N_1946,N_1981);
nor U2006 (N_2006,N_1948,N_1954);
nand U2007 (N_2007,N_1884,N_1825);
or U2008 (N_2008,N_1843,N_1800);
and U2009 (N_2009,N_1844,N_1905);
or U2010 (N_2010,N_1966,N_1974);
or U2011 (N_2011,N_1969,N_1838);
nand U2012 (N_2012,N_1895,N_1842);
or U2013 (N_2013,N_1949,N_1918);
or U2014 (N_2014,N_1814,N_1898);
xor U2015 (N_2015,N_1935,N_1923);
xor U2016 (N_2016,N_1956,N_1882);
and U2017 (N_2017,N_1989,N_1963);
xor U2018 (N_2018,N_1967,N_1965);
nor U2019 (N_2019,N_1836,N_1916);
nor U2020 (N_2020,N_1851,N_1933);
or U2021 (N_2021,N_1901,N_1823);
xor U2022 (N_2022,N_1805,N_1925);
nand U2023 (N_2023,N_1924,N_1870);
xnor U2024 (N_2024,N_1865,N_1970);
nand U2025 (N_2025,N_1907,N_1863);
nand U2026 (N_2026,N_1821,N_1826);
and U2027 (N_2027,N_1926,N_1928);
nor U2028 (N_2028,N_1808,N_1847);
nand U2029 (N_2029,N_1837,N_1910);
nand U2030 (N_2030,N_1846,N_1961);
and U2031 (N_2031,N_1906,N_1861);
xnor U2032 (N_2032,N_1862,N_1912);
nand U2033 (N_2033,N_1818,N_1899);
or U2034 (N_2034,N_1968,N_1932);
nand U2035 (N_2035,N_1943,N_1885);
nor U2036 (N_2036,N_1975,N_1950);
nand U2037 (N_2037,N_1883,N_1804);
nand U2038 (N_2038,N_1921,N_1915);
and U2039 (N_2039,N_1940,N_1858);
nand U2040 (N_2040,N_1845,N_1902);
nand U2041 (N_2041,N_1992,N_1913);
nor U2042 (N_2042,N_1829,N_1831);
nand U2043 (N_2043,N_1815,N_1816);
and U2044 (N_2044,N_1993,N_1822);
nand U2045 (N_2045,N_1802,N_1834);
or U2046 (N_2046,N_1876,N_1897);
nor U2047 (N_2047,N_1850,N_1985);
nand U2048 (N_2048,N_1994,N_1980);
or U2049 (N_2049,N_1840,N_1962);
and U2050 (N_2050,N_1922,N_1807);
or U2051 (N_2051,N_1881,N_1927);
and U2052 (N_2052,N_1958,N_1971);
and U2053 (N_2053,N_1860,N_1887);
xor U2054 (N_2054,N_1812,N_1857);
xor U2055 (N_2055,N_1973,N_1855);
and U2056 (N_2056,N_1896,N_1991);
nor U2057 (N_2057,N_1978,N_1936);
nor U2058 (N_2058,N_1864,N_1903);
nand U2059 (N_2059,N_1911,N_1839);
nand U2060 (N_2060,N_1904,N_1877);
and U2061 (N_2061,N_1833,N_1977);
or U2062 (N_2062,N_1830,N_1873);
nand U2063 (N_2063,N_1939,N_1890);
or U2064 (N_2064,N_1809,N_1811);
nor U2065 (N_2065,N_1869,N_1953);
xor U2066 (N_2066,N_1859,N_1832);
xor U2067 (N_2067,N_1892,N_1900);
nand U2068 (N_2068,N_1908,N_1879);
nor U2069 (N_2069,N_1995,N_1872);
xnor U2070 (N_2070,N_1874,N_1867);
xor U2071 (N_2071,N_1982,N_1820);
xnor U2072 (N_2072,N_1917,N_1817);
nand U2073 (N_2073,N_1937,N_1852);
nor U2074 (N_2074,N_1947,N_1959);
nor U2075 (N_2075,N_1841,N_1848);
and U2076 (N_2076,N_1803,N_1952);
nand U2077 (N_2077,N_1824,N_1951);
xnor U2078 (N_2078,N_1888,N_1827);
nand U2079 (N_2079,N_1944,N_1931);
nor U2080 (N_2080,N_1990,N_1979);
xnor U2081 (N_2081,N_1886,N_1810);
nor U2082 (N_2082,N_1878,N_1871);
or U2083 (N_2083,N_1964,N_1998);
nor U2084 (N_2084,N_1868,N_1942);
nor U2085 (N_2085,N_1801,N_1875);
and U2086 (N_2086,N_1988,N_1930);
and U2087 (N_2087,N_1893,N_1880);
xor U2088 (N_2088,N_1934,N_1941);
xnor U2089 (N_2089,N_1914,N_1849);
nand U2090 (N_2090,N_1957,N_1955);
and U2091 (N_2091,N_1945,N_1920);
nand U2092 (N_2092,N_1828,N_1866);
and U2093 (N_2093,N_1835,N_1986);
or U2094 (N_2094,N_1919,N_1909);
nand U2095 (N_2095,N_1894,N_1960);
and U2096 (N_2096,N_1997,N_1856);
and U2097 (N_2097,N_1853,N_1983);
nand U2098 (N_2098,N_1819,N_1938);
nand U2099 (N_2099,N_1999,N_1987);
nor U2100 (N_2100,N_1992,N_1831);
nand U2101 (N_2101,N_1821,N_1869);
xor U2102 (N_2102,N_1931,N_1975);
nand U2103 (N_2103,N_1845,N_1994);
nor U2104 (N_2104,N_1949,N_1879);
nor U2105 (N_2105,N_1900,N_1936);
nor U2106 (N_2106,N_1939,N_1863);
nand U2107 (N_2107,N_1884,N_1857);
xor U2108 (N_2108,N_1879,N_1800);
nand U2109 (N_2109,N_1824,N_1998);
nand U2110 (N_2110,N_1871,N_1918);
and U2111 (N_2111,N_1992,N_1802);
xor U2112 (N_2112,N_1945,N_1864);
xnor U2113 (N_2113,N_1907,N_1967);
nor U2114 (N_2114,N_1830,N_1919);
nor U2115 (N_2115,N_1941,N_1981);
xor U2116 (N_2116,N_1893,N_1967);
nor U2117 (N_2117,N_1962,N_1941);
or U2118 (N_2118,N_1928,N_1800);
xor U2119 (N_2119,N_1868,N_1858);
and U2120 (N_2120,N_1842,N_1901);
or U2121 (N_2121,N_1900,N_1977);
and U2122 (N_2122,N_1854,N_1844);
xnor U2123 (N_2123,N_1894,N_1979);
or U2124 (N_2124,N_1928,N_1839);
xor U2125 (N_2125,N_1852,N_1881);
and U2126 (N_2126,N_1849,N_1888);
nand U2127 (N_2127,N_1856,N_1940);
xor U2128 (N_2128,N_1941,N_1894);
xnor U2129 (N_2129,N_1838,N_1870);
nand U2130 (N_2130,N_1888,N_1945);
xnor U2131 (N_2131,N_1817,N_1920);
xor U2132 (N_2132,N_1970,N_1984);
xnor U2133 (N_2133,N_1875,N_1865);
and U2134 (N_2134,N_1878,N_1994);
nand U2135 (N_2135,N_1874,N_1908);
nor U2136 (N_2136,N_1895,N_1976);
or U2137 (N_2137,N_1890,N_1987);
nand U2138 (N_2138,N_1891,N_1868);
and U2139 (N_2139,N_1995,N_1821);
and U2140 (N_2140,N_1990,N_1966);
nand U2141 (N_2141,N_1961,N_1836);
and U2142 (N_2142,N_1811,N_1907);
nor U2143 (N_2143,N_1933,N_1801);
or U2144 (N_2144,N_1939,N_1826);
and U2145 (N_2145,N_1897,N_1982);
nand U2146 (N_2146,N_1896,N_1890);
and U2147 (N_2147,N_1878,N_1954);
nand U2148 (N_2148,N_1893,N_1819);
nand U2149 (N_2149,N_1911,N_1982);
nor U2150 (N_2150,N_1878,N_1969);
nand U2151 (N_2151,N_1807,N_1972);
and U2152 (N_2152,N_1910,N_1847);
and U2153 (N_2153,N_1808,N_1809);
or U2154 (N_2154,N_1923,N_1833);
nand U2155 (N_2155,N_1903,N_1917);
or U2156 (N_2156,N_1917,N_1923);
or U2157 (N_2157,N_1980,N_1804);
xnor U2158 (N_2158,N_1806,N_1926);
or U2159 (N_2159,N_1953,N_1842);
nand U2160 (N_2160,N_1991,N_1901);
and U2161 (N_2161,N_1847,N_1881);
or U2162 (N_2162,N_1829,N_1998);
and U2163 (N_2163,N_1845,N_1972);
and U2164 (N_2164,N_1838,N_1957);
xor U2165 (N_2165,N_1958,N_1932);
and U2166 (N_2166,N_1830,N_1983);
or U2167 (N_2167,N_1960,N_1885);
or U2168 (N_2168,N_1902,N_1892);
nand U2169 (N_2169,N_1894,N_1909);
nor U2170 (N_2170,N_1845,N_1895);
or U2171 (N_2171,N_1866,N_1814);
xor U2172 (N_2172,N_1817,N_1996);
and U2173 (N_2173,N_1963,N_1843);
or U2174 (N_2174,N_1911,N_1812);
xnor U2175 (N_2175,N_1868,N_1898);
xor U2176 (N_2176,N_1984,N_1955);
or U2177 (N_2177,N_1986,N_1806);
xor U2178 (N_2178,N_1906,N_1853);
xnor U2179 (N_2179,N_1933,N_1929);
xor U2180 (N_2180,N_1835,N_1902);
nand U2181 (N_2181,N_1807,N_1895);
xnor U2182 (N_2182,N_1807,N_1878);
or U2183 (N_2183,N_1907,N_1815);
or U2184 (N_2184,N_1810,N_1892);
nand U2185 (N_2185,N_1887,N_1986);
xnor U2186 (N_2186,N_1898,N_1833);
or U2187 (N_2187,N_1860,N_1841);
nand U2188 (N_2188,N_1924,N_1946);
nand U2189 (N_2189,N_1965,N_1825);
and U2190 (N_2190,N_1830,N_1964);
and U2191 (N_2191,N_1818,N_1902);
nand U2192 (N_2192,N_1988,N_1894);
or U2193 (N_2193,N_1802,N_1847);
or U2194 (N_2194,N_1802,N_1879);
or U2195 (N_2195,N_1893,N_1956);
nand U2196 (N_2196,N_1947,N_1970);
xnor U2197 (N_2197,N_1988,N_1929);
nand U2198 (N_2198,N_1938,N_1862);
and U2199 (N_2199,N_1898,N_1947);
nor U2200 (N_2200,N_2025,N_2106);
nand U2201 (N_2201,N_2154,N_2089);
xnor U2202 (N_2202,N_2000,N_2037);
xnor U2203 (N_2203,N_2052,N_2074);
nor U2204 (N_2204,N_2149,N_2158);
or U2205 (N_2205,N_2161,N_2076);
and U2206 (N_2206,N_2028,N_2031);
or U2207 (N_2207,N_2040,N_2193);
xor U2208 (N_2208,N_2088,N_2012);
xor U2209 (N_2209,N_2116,N_2094);
nand U2210 (N_2210,N_2046,N_2062);
xor U2211 (N_2211,N_2050,N_2068);
and U2212 (N_2212,N_2199,N_2023);
and U2213 (N_2213,N_2035,N_2159);
or U2214 (N_2214,N_2093,N_2067);
or U2215 (N_2215,N_2188,N_2143);
and U2216 (N_2216,N_2181,N_2121);
xnor U2217 (N_2217,N_2174,N_2078);
nand U2218 (N_2218,N_2118,N_2080);
xnor U2219 (N_2219,N_2160,N_2058);
or U2220 (N_2220,N_2103,N_2087);
and U2221 (N_2221,N_2086,N_2126);
nand U2222 (N_2222,N_2108,N_2085);
or U2223 (N_2223,N_2195,N_2018);
xnor U2224 (N_2224,N_2186,N_2022);
xor U2225 (N_2225,N_2044,N_2135);
xor U2226 (N_2226,N_2138,N_2079);
nand U2227 (N_2227,N_2100,N_2069);
xnor U2228 (N_2228,N_2101,N_2075);
nand U2229 (N_2229,N_2110,N_2197);
xnor U2230 (N_2230,N_2027,N_2082);
nor U2231 (N_2231,N_2130,N_2041);
nand U2232 (N_2232,N_2125,N_2163);
xor U2233 (N_2233,N_2141,N_2051);
or U2234 (N_2234,N_2152,N_2166);
xor U2235 (N_2235,N_2001,N_2104);
and U2236 (N_2236,N_2169,N_2172);
nor U2237 (N_2237,N_2131,N_2147);
nand U2238 (N_2238,N_2115,N_2060);
and U2239 (N_2239,N_2179,N_2029);
and U2240 (N_2240,N_2055,N_2008);
nor U2241 (N_2241,N_2064,N_2002);
or U2242 (N_2242,N_2117,N_2170);
or U2243 (N_2243,N_2184,N_2081);
or U2244 (N_2244,N_2146,N_2043);
and U2245 (N_2245,N_2003,N_2155);
or U2246 (N_2246,N_2190,N_2173);
and U2247 (N_2247,N_2175,N_2164);
xnor U2248 (N_2248,N_2016,N_2083);
or U2249 (N_2249,N_2059,N_2033);
nand U2250 (N_2250,N_2127,N_2053);
xor U2251 (N_2251,N_2057,N_2180);
nand U2252 (N_2252,N_2054,N_2198);
nand U2253 (N_2253,N_2134,N_2151);
or U2254 (N_2254,N_2133,N_2178);
nand U2255 (N_2255,N_2061,N_2038);
nor U2256 (N_2256,N_2098,N_2020);
nor U2257 (N_2257,N_2030,N_2063);
nand U2258 (N_2258,N_2036,N_2049);
and U2259 (N_2259,N_2096,N_2091);
xnor U2260 (N_2260,N_2010,N_2182);
nand U2261 (N_2261,N_2191,N_2119);
nor U2262 (N_2262,N_2015,N_2132);
xnor U2263 (N_2263,N_2153,N_2092);
and U2264 (N_2264,N_2021,N_2072);
nand U2265 (N_2265,N_2007,N_2129);
or U2266 (N_2266,N_2148,N_2113);
xor U2267 (N_2267,N_2009,N_2168);
xor U2268 (N_2268,N_2066,N_2124);
or U2269 (N_2269,N_2090,N_2165);
nor U2270 (N_2270,N_2144,N_2019);
nor U2271 (N_2271,N_2192,N_2128);
xor U2272 (N_2272,N_2048,N_2039);
nand U2273 (N_2273,N_2006,N_2084);
and U2274 (N_2274,N_2196,N_2157);
nor U2275 (N_2275,N_2187,N_2167);
or U2276 (N_2276,N_2099,N_2139);
nand U2277 (N_2277,N_2026,N_2034);
nor U2278 (N_2278,N_2013,N_2183);
and U2279 (N_2279,N_2189,N_2095);
nor U2280 (N_2280,N_2077,N_2145);
or U2281 (N_2281,N_2045,N_2004);
and U2282 (N_2282,N_2065,N_2011);
xnor U2283 (N_2283,N_2194,N_2014);
xnor U2284 (N_2284,N_2056,N_2122);
xor U2285 (N_2285,N_2112,N_2123);
or U2286 (N_2286,N_2073,N_2114);
xnor U2287 (N_2287,N_2005,N_2032);
nor U2288 (N_2288,N_2042,N_2017);
and U2289 (N_2289,N_2102,N_2185);
xnor U2290 (N_2290,N_2176,N_2024);
nand U2291 (N_2291,N_2120,N_2105);
and U2292 (N_2292,N_2140,N_2070);
nor U2293 (N_2293,N_2156,N_2177);
and U2294 (N_2294,N_2137,N_2150);
xnor U2295 (N_2295,N_2162,N_2142);
nand U2296 (N_2296,N_2071,N_2111);
nand U2297 (N_2297,N_2047,N_2171);
nand U2298 (N_2298,N_2109,N_2097);
nand U2299 (N_2299,N_2136,N_2107);
xor U2300 (N_2300,N_2056,N_2002);
xnor U2301 (N_2301,N_2138,N_2175);
xnor U2302 (N_2302,N_2046,N_2174);
and U2303 (N_2303,N_2182,N_2004);
nor U2304 (N_2304,N_2049,N_2098);
nand U2305 (N_2305,N_2034,N_2007);
xnor U2306 (N_2306,N_2038,N_2107);
nand U2307 (N_2307,N_2083,N_2065);
or U2308 (N_2308,N_2060,N_2053);
and U2309 (N_2309,N_2188,N_2109);
or U2310 (N_2310,N_2194,N_2106);
or U2311 (N_2311,N_2093,N_2121);
nor U2312 (N_2312,N_2065,N_2097);
xnor U2313 (N_2313,N_2147,N_2137);
nand U2314 (N_2314,N_2125,N_2044);
xnor U2315 (N_2315,N_2033,N_2183);
and U2316 (N_2316,N_2073,N_2142);
or U2317 (N_2317,N_2146,N_2139);
nor U2318 (N_2318,N_2072,N_2160);
or U2319 (N_2319,N_2162,N_2143);
nand U2320 (N_2320,N_2172,N_2188);
nor U2321 (N_2321,N_2041,N_2009);
and U2322 (N_2322,N_2127,N_2132);
nand U2323 (N_2323,N_2140,N_2105);
or U2324 (N_2324,N_2007,N_2122);
xnor U2325 (N_2325,N_2075,N_2085);
or U2326 (N_2326,N_2181,N_2020);
nand U2327 (N_2327,N_2047,N_2155);
or U2328 (N_2328,N_2069,N_2006);
or U2329 (N_2329,N_2116,N_2093);
nand U2330 (N_2330,N_2166,N_2180);
xor U2331 (N_2331,N_2051,N_2135);
nor U2332 (N_2332,N_2122,N_2009);
and U2333 (N_2333,N_2022,N_2196);
nand U2334 (N_2334,N_2135,N_2084);
xnor U2335 (N_2335,N_2088,N_2170);
or U2336 (N_2336,N_2156,N_2179);
or U2337 (N_2337,N_2092,N_2113);
and U2338 (N_2338,N_2190,N_2148);
nand U2339 (N_2339,N_2048,N_2052);
and U2340 (N_2340,N_2197,N_2180);
and U2341 (N_2341,N_2030,N_2107);
xor U2342 (N_2342,N_2184,N_2148);
or U2343 (N_2343,N_2116,N_2179);
nor U2344 (N_2344,N_2125,N_2094);
and U2345 (N_2345,N_2189,N_2192);
nor U2346 (N_2346,N_2024,N_2142);
nand U2347 (N_2347,N_2182,N_2145);
and U2348 (N_2348,N_2173,N_2130);
and U2349 (N_2349,N_2123,N_2021);
or U2350 (N_2350,N_2135,N_2086);
xor U2351 (N_2351,N_2176,N_2061);
nand U2352 (N_2352,N_2176,N_2183);
xor U2353 (N_2353,N_2193,N_2166);
nor U2354 (N_2354,N_2100,N_2186);
nand U2355 (N_2355,N_2022,N_2073);
and U2356 (N_2356,N_2028,N_2132);
nand U2357 (N_2357,N_2037,N_2067);
nand U2358 (N_2358,N_2161,N_2030);
nor U2359 (N_2359,N_2006,N_2031);
xnor U2360 (N_2360,N_2026,N_2116);
nand U2361 (N_2361,N_2000,N_2062);
and U2362 (N_2362,N_2111,N_2197);
nor U2363 (N_2363,N_2067,N_2170);
or U2364 (N_2364,N_2158,N_2132);
or U2365 (N_2365,N_2157,N_2122);
nor U2366 (N_2366,N_2190,N_2139);
or U2367 (N_2367,N_2054,N_2190);
nand U2368 (N_2368,N_2066,N_2163);
xor U2369 (N_2369,N_2026,N_2085);
nor U2370 (N_2370,N_2059,N_2046);
nand U2371 (N_2371,N_2082,N_2180);
xnor U2372 (N_2372,N_2194,N_2048);
nand U2373 (N_2373,N_2003,N_2172);
nand U2374 (N_2374,N_2022,N_2177);
nand U2375 (N_2375,N_2171,N_2122);
and U2376 (N_2376,N_2194,N_2193);
or U2377 (N_2377,N_2122,N_2046);
nor U2378 (N_2378,N_2137,N_2084);
nand U2379 (N_2379,N_2176,N_2078);
xnor U2380 (N_2380,N_2094,N_2089);
nand U2381 (N_2381,N_2132,N_2114);
nor U2382 (N_2382,N_2095,N_2019);
xor U2383 (N_2383,N_2131,N_2169);
and U2384 (N_2384,N_2106,N_2116);
or U2385 (N_2385,N_2115,N_2113);
and U2386 (N_2386,N_2081,N_2115);
and U2387 (N_2387,N_2051,N_2064);
xnor U2388 (N_2388,N_2108,N_2011);
xnor U2389 (N_2389,N_2152,N_2074);
and U2390 (N_2390,N_2015,N_2083);
and U2391 (N_2391,N_2180,N_2059);
and U2392 (N_2392,N_2124,N_2126);
nor U2393 (N_2393,N_2158,N_2017);
and U2394 (N_2394,N_2179,N_2110);
nor U2395 (N_2395,N_2164,N_2159);
and U2396 (N_2396,N_2142,N_2082);
or U2397 (N_2397,N_2068,N_2117);
nand U2398 (N_2398,N_2148,N_2059);
nor U2399 (N_2399,N_2059,N_2000);
nor U2400 (N_2400,N_2343,N_2386);
nor U2401 (N_2401,N_2375,N_2301);
or U2402 (N_2402,N_2272,N_2310);
or U2403 (N_2403,N_2232,N_2329);
nand U2404 (N_2404,N_2210,N_2393);
xor U2405 (N_2405,N_2308,N_2366);
and U2406 (N_2406,N_2291,N_2239);
nand U2407 (N_2407,N_2280,N_2256);
nand U2408 (N_2408,N_2251,N_2389);
nor U2409 (N_2409,N_2219,N_2303);
or U2410 (N_2410,N_2316,N_2344);
nand U2411 (N_2411,N_2306,N_2346);
and U2412 (N_2412,N_2276,N_2286);
nand U2413 (N_2413,N_2244,N_2296);
or U2414 (N_2414,N_2294,N_2322);
nor U2415 (N_2415,N_2222,N_2265);
and U2416 (N_2416,N_2289,N_2277);
nor U2417 (N_2417,N_2388,N_2279);
nand U2418 (N_2418,N_2230,N_2227);
and U2419 (N_2419,N_2284,N_2309);
nor U2420 (N_2420,N_2337,N_2361);
or U2421 (N_2421,N_2332,N_2338);
nor U2422 (N_2422,N_2311,N_2245);
nand U2423 (N_2423,N_2398,N_2274);
nor U2424 (N_2424,N_2395,N_2328);
xor U2425 (N_2425,N_2313,N_2266);
and U2426 (N_2426,N_2243,N_2257);
nand U2427 (N_2427,N_2317,N_2369);
xnor U2428 (N_2428,N_2209,N_2318);
nor U2429 (N_2429,N_2267,N_2224);
nand U2430 (N_2430,N_2249,N_2264);
xor U2431 (N_2431,N_2233,N_2390);
xnor U2432 (N_2432,N_2370,N_2312);
or U2433 (N_2433,N_2285,N_2391);
or U2434 (N_2434,N_2207,N_2215);
and U2435 (N_2435,N_2324,N_2283);
or U2436 (N_2436,N_2359,N_2340);
and U2437 (N_2437,N_2315,N_2213);
and U2438 (N_2438,N_2342,N_2260);
nor U2439 (N_2439,N_2208,N_2278);
nand U2440 (N_2440,N_2360,N_2218);
and U2441 (N_2441,N_2392,N_2238);
nor U2442 (N_2442,N_2206,N_2374);
nand U2443 (N_2443,N_2226,N_2211);
nor U2444 (N_2444,N_2259,N_2216);
xnor U2445 (N_2445,N_2353,N_2368);
and U2446 (N_2446,N_2247,N_2348);
nand U2447 (N_2447,N_2268,N_2304);
nand U2448 (N_2448,N_2205,N_2383);
or U2449 (N_2449,N_2203,N_2378);
xnor U2450 (N_2450,N_2221,N_2293);
xnor U2451 (N_2451,N_2214,N_2335);
nand U2452 (N_2452,N_2326,N_2349);
or U2453 (N_2453,N_2352,N_2292);
nor U2454 (N_2454,N_2365,N_2380);
or U2455 (N_2455,N_2347,N_2307);
nand U2456 (N_2456,N_2220,N_2282);
nand U2457 (N_2457,N_2382,N_2297);
or U2458 (N_2458,N_2248,N_2364);
nand U2459 (N_2459,N_2362,N_2331);
xor U2460 (N_2460,N_2202,N_2397);
or U2461 (N_2461,N_2235,N_2254);
nor U2462 (N_2462,N_2258,N_2363);
and U2463 (N_2463,N_2354,N_2288);
nor U2464 (N_2464,N_2201,N_2261);
xnor U2465 (N_2465,N_2334,N_2229);
nor U2466 (N_2466,N_2379,N_2394);
nor U2467 (N_2467,N_2355,N_2305);
nor U2468 (N_2468,N_2381,N_2270);
or U2469 (N_2469,N_2336,N_2341);
and U2470 (N_2470,N_2200,N_2314);
nor U2471 (N_2471,N_2384,N_2236);
xnor U2472 (N_2472,N_2217,N_2387);
or U2473 (N_2473,N_2357,N_2295);
nand U2474 (N_2474,N_2319,N_2320);
xnor U2475 (N_2475,N_2358,N_2399);
nor U2476 (N_2476,N_2298,N_2263);
xor U2477 (N_2477,N_2376,N_2253);
and U2478 (N_2478,N_2275,N_2255);
nor U2479 (N_2479,N_2273,N_2350);
nand U2480 (N_2480,N_2250,N_2237);
nand U2481 (N_2481,N_2351,N_2302);
nand U2482 (N_2482,N_2373,N_2262);
nand U2483 (N_2483,N_2204,N_2345);
and U2484 (N_2484,N_2300,N_2234);
and U2485 (N_2485,N_2228,N_2299);
and U2486 (N_2486,N_2356,N_2367);
or U2487 (N_2487,N_2281,N_2325);
and U2488 (N_2488,N_2231,N_2269);
nor U2489 (N_2489,N_2271,N_2371);
and U2490 (N_2490,N_2323,N_2223);
nand U2491 (N_2491,N_2290,N_2212);
xor U2492 (N_2492,N_2385,N_2287);
xnor U2493 (N_2493,N_2225,N_2241);
and U2494 (N_2494,N_2246,N_2339);
xnor U2495 (N_2495,N_2242,N_2327);
nand U2496 (N_2496,N_2240,N_2321);
nor U2497 (N_2497,N_2252,N_2396);
and U2498 (N_2498,N_2377,N_2330);
nor U2499 (N_2499,N_2333,N_2372);
nand U2500 (N_2500,N_2386,N_2364);
nor U2501 (N_2501,N_2308,N_2290);
nand U2502 (N_2502,N_2369,N_2288);
and U2503 (N_2503,N_2390,N_2241);
nor U2504 (N_2504,N_2362,N_2261);
nand U2505 (N_2505,N_2226,N_2384);
xnor U2506 (N_2506,N_2252,N_2389);
nand U2507 (N_2507,N_2322,N_2323);
and U2508 (N_2508,N_2386,N_2244);
nor U2509 (N_2509,N_2276,N_2320);
and U2510 (N_2510,N_2202,N_2362);
nor U2511 (N_2511,N_2336,N_2316);
nor U2512 (N_2512,N_2288,N_2278);
or U2513 (N_2513,N_2318,N_2293);
or U2514 (N_2514,N_2261,N_2390);
nor U2515 (N_2515,N_2239,N_2235);
xnor U2516 (N_2516,N_2273,N_2345);
xnor U2517 (N_2517,N_2277,N_2276);
xnor U2518 (N_2518,N_2395,N_2211);
nor U2519 (N_2519,N_2283,N_2318);
and U2520 (N_2520,N_2315,N_2310);
or U2521 (N_2521,N_2237,N_2388);
or U2522 (N_2522,N_2237,N_2357);
and U2523 (N_2523,N_2300,N_2243);
nor U2524 (N_2524,N_2367,N_2274);
nor U2525 (N_2525,N_2304,N_2271);
or U2526 (N_2526,N_2347,N_2260);
nor U2527 (N_2527,N_2392,N_2334);
xor U2528 (N_2528,N_2397,N_2341);
nor U2529 (N_2529,N_2306,N_2207);
or U2530 (N_2530,N_2285,N_2222);
xor U2531 (N_2531,N_2347,N_2257);
or U2532 (N_2532,N_2231,N_2393);
nand U2533 (N_2533,N_2294,N_2245);
nor U2534 (N_2534,N_2264,N_2301);
xor U2535 (N_2535,N_2266,N_2336);
xnor U2536 (N_2536,N_2221,N_2204);
and U2537 (N_2537,N_2216,N_2388);
and U2538 (N_2538,N_2257,N_2239);
nand U2539 (N_2539,N_2322,N_2209);
or U2540 (N_2540,N_2243,N_2348);
nand U2541 (N_2541,N_2337,N_2247);
and U2542 (N_2542,N_2320,N_2261);
and U2543 (N_2543,N_2264,N_2266);
nor U2544 (N_2544,N_2213,N_2265);
nor U2545 (N_2545,N_2313,N_2328);
xnor U2546 (N_2546,N_2218,N_2294);
nand U2547 (N_2547,N_2229,N_2294);
nand U2548 (N_2548,N_2255,N_2220);
xor U2549 (N_2549,N_2214,N_2299);
and U2550 (N_2550,N_2204,N_2229);
nand U2551 (N_2551,N_2280,N_2364);
xor U2552 (N_2552,N_2352,N_2382);
xor U2553 (N_2553,N_2361,N_2232);
and U2554 (N_2554,N_2237,N_2229);
nand U2555 (N_2555,N_2374,N_2283);
xor U2556 (N_2556,N_2321,N_2290);
nand U2557 (N_2557,N_2367,N_2331);
and U2558 (N_2558,N_2317,N_2347);
and U2559 (N_2559,N_2389,N_2373);
nand U2560 (N_2560,N_2233,N_2222);
and U2561 (N_2561,N_2369,N_2290);
nand U2562 (N_2562,N_2374,N_2295);
xor U2563 (N_2563,N_2273,N_2223);
nand U2564 (N_2564,N_2201,N_2288);
and U2565 (N_2565,N_2250,N_2262);
xnor U2566 (N_2566,N_2376,N_2336);
and U2567 (N_2567,N_2350,N_2342);
nand U2568 (N_2568,N_2328,N_2239);
and U2569 (N_2569,N_2310,N_2279);
nor U2570 (N_2570,N_2247,N_2396);
nor U2571 (N_2571,N_2362,N_2249);
nand U2572 (N_2572,N_2387,N_2393);
or U2573 (N_2573,N_2236,N_2284);
xnor U2574 (N_2574,N_2352,N_2221);
nand U2575 (N_2575,N_2230,N_2205);
and U2576 (N_2576,N_2300,N_2301);
nor U2577 (N_2577,N_2324,N_2352);
and U2578 (N_2578,N_2216,N_2234);
and U2579 (N_2579,N_2391,N_2281);
xnor U2580 (N_2580,N_2250,N_2390);
nand U2581 (N_2581,N_2336,N_2390);
nor U2582 (N_2582,N_2308,N_2352);
nand U2583 (N_2583,N_2366,N_2352);
and U2584 (N_2584,N_2261,N_2258);
or U2585 (N_2585,N_2391,N_2219);
and U2586 (N_2586,N_2231,N_2252);
xnor U2587 (N_2587,N_2355,N_2251);
nor U2588 (N_2588,N_2301,N_2340);
xnor U2589 (N_2589,N_2291,N_2206);
and U2590 (N_2590,N_2399,N_2309);
xor U2591 (N_2591,N_2267,N_2323);
nor U2592 (N_2592,N_2338,N_2378);
or U2593 (N_2593,N_2340,N_2289);
xor U2594 (N_2594,N_2375,N_2320);
xor U2595 (N_2595,N_2242,N_2316);
and U2596 (N_2596,N_2313,N_2212);
and U2597 (N_2597,N_2206,N_2336);
xor U2598 (N_2598,N_2293,N_2309);
or U2599 (N_2599,N_2267,N_2309);
and U2600 (N_2600,N_2504,N_2475);
xnor U2601 (N_2601,N_2592,N_2441);
nand U2602 (N_2602,N_2521,N_2543);
xor U2603 (N_2603,N_2505,N_2477);
and U2604 (N_2604,N_2414,N_2501);
xnor U2605 (N_2605,N_2489,N_2553);
or U2606 (N_2606,N_2582,N_2541);
xnor U2607 (N_2607,N_2495,N_2406);
and U2608 (N_2608,N_2470,N_2481);
and U2609 (N_2609,N_2528,N_2454);
xnor U2610 (N_2610,N_2448,N_2415);
xor U2611 (N_2611,N_2591,N_2588);
and U2612 (N_2612,N_2514,N_2532);
or U2613 (N_2613,N_2416,N_2427);
or U2614 (N_2614,N_2485,N_2438);
and U2615 (N_2615,N_2584,N_2422);
nand U2616 (N_2616,N_2431,N_2516);
nand U2617 (N_2617,N_2542,N_2443);
and U2618 (N_2618,N_2401,N_2418);
nand U2619 (N_2619,N_2417,N_2439);
or U2620 (N_2620,N_2435,N_2434);
nand U2621 (N_2621,N_2508,N_2529);
xor U2622 (N_2622,N_2594,N_2590);
nand U2623 (N_2623,N_2445,N_2507);
and U2624 (N_2624,N_2420,N_2493);
nor U2625 (N_2625,N_2460,N_2536);
or U2626 (N_2626,N_2500,N_2570);
xnor U2627 (N_2627,N_2535,N_2565);
and U2628 (N_2628,N_2465,N_2599);
xnor U2629 (N_2629,N_2469,N_2474);
and U2630 (N_2630,N_2423,N_2523);
and U2631 (N_2631,N_2513,N_2517);
nor U2632 (N_2632,N_2561,N_2597);
nor U2633 (N_2633,N_2581,N_2412);
xnor U2634 (N_2634,N_2544,N_2425);
xor U2635 (N_2635,N_2539,N_2571);
or U2636 (N_2636,N_2569,N_2440);
and U2637 (N_2637,N_2442,N_2555);
or U2638 (N_2638,N_2506,N_2446);
and U2639 (N_2639,N_2540,N_2518);
nand U2640 (N_2640,N_2486,N_2547);
nor U2641 (N_2641,N_2464,N_2545);
or U2642 (N_2642,N_2436,N_2566);
or U2643 (N_2643,N_2548,N_2429);
nand U2644 (N_2644,N_2538,N_2476);
xor U2645 (N_2645,N_2478,N_2527);
or U2646 (N_2646,N_2549,N_2575);
xor U2647 (N_2647,N_2578,N_2428);
nor U2648 (N_2648,N_2473,N_2519);
nor U2649 (N_2649,N_2410,N_2558);
nand U2650 (N_2650,N_2403,N_2444);
or U2651 (N_2651,N_2499,N_2580);
nor U2652 (N_2652,N_2522,N_2596);
and U2653 (N_2653,N_2573,N_2509);
or U2654 (N_2654,N_2466,N_2472);
or U2655 (N_2655,N_2494,N_2408);
or U2656 (N_2656,N_2576,N_2463);
nor U2657 (N_2657,N_2451,N_2430);
and U2658 (N_2658,N_2490,N_2562);
nor U2659 (N_2659,N_2526,N_2595);
or U2660 (N_2660,N_2559,N_2450);
and U2661 (N_2661,N_2447,N_2471);
xnor U2662 (N_2662,N_2492,N_2552);
and U2663 (N_2663,N_2409,N_2402);
xor U2664 (N_2664,N_2583,N_2534);
xnor U2665 (N_2665,N_2498,N_2564);
nand U2666 (N_2666,N_2491,N_2511);
and U2667 (N_2667,N_2587,N_2468);
xnor U2668 (N_2668,N_2457,N_2512);
nor U2669 (N_2669,N_2586,N_2598);
or U2670 (N_2670,N_2574,N_2531);
xnor U2671 (N_2671,N_2426,N_2515);
xor U2672 (N_2672,N_2589,N_2482);
xor U2673 (N_2673,N_2537,N_2449);
or U2674 (N_2674,N_2567,N_2497);
nor U2675 (N_2675,N_2487,N_2405);
xnor U2676 (N_2676,N_2568,N_2467);
and U2677 (N_2677,N_2550,N_2433);
or U2678 (N_2678,N_2437,N_2453);
or U2679 (N_2679,N_2452,N_2413);
or U2680 (N_2680,N_2502,N_2458);
nor U2681 (N_2681,N_2419,N_2563);
xor U2682 (N_2682,N_2560,N_2455);
or U2683 (N_2683,N_2459,N_2483);
xor U2684 (N_2684,N_2551,N_2456);
nand U2685 (N_2685,N_2432,N_2546);
or U2686 (N_2686,N_2407,N_2488);
or U2687 (N_2687,N_2533,N_2593);
or U2688 (N_2688,N_2525,N_2530);
xnor U2689 (N_2689,N_2400,N_2510);
nand U2690 (N_2690,N_2585,N_2461);
xor U2691 (N_2691,N_2484,N_2554);
nand U2692 (N_2692,N_2462,N_2520);
nor U2693 (N_2693,N_2524,N_2421);
xnor U2694 (N_2694,N_2572,N_2424);
and U2695 (N_2695,N_2577,N_2556);
nor U2696 (N_2696,N_2557,N_2496);
or U2697 (N_2697,N_2579,N_2404);
nand U2698 (N_2698,N_2479,N_2480);
and U2699 (N_2699,N_2411,N_2503);
nor U2700 (N_2700,N_2422,N_2416);
nor U2701 (N_2701,N_2486,N_2527);
xor U2702 (N_2702,N_2506,N_2513);
nor U2703 (N_2703,N_2563,N_2593);
xor U2704 (N_2704,N_2459,N_2511);
nand U2705 (N_2705,N_2440,N_2465);
nand U2706 (N_2706,N_2448,N_2523);
nand U2707 (N_2707,N_2468,N_2452);
or U2708 (N_2708,N_2447,N_2552);
or U2709 (N_2709,N_2478,N_2549);
nor U2710 (N_2710,N_2550,N_2513);
and U2711 (N_2711,N_2452,N_2547);
or U2712 (N_2712,N_2559,N_2542);
nor U2713 (N_2713,N_2423,N_2506);
nor U2714 (N_2714,N_2429,N_2422);
or U2715 (N_2715,N_2591,N_2460);
nor U2716 (N_2716,N_2558,N_2582);
nor U2717 (N_2717,N_2438,N_2592);
nor U2718 (N_2718,N_2540,N_2570);
or U2719 (N_2719,N_2542,N_2581);
nor U2720 (N_2720,N_2500,N_2582);
or U2721 (N_2721,N_2404,N_2411);
nand U2722 (N_2722,N_2406,N_2550);
nor U2723 (N_2723,N_2474,N_2501);
nand U2724 (N_2724,N_2491,N_2418);
nand U2725 (N_2725,N_2536,N_2564);
xnor U2726 (N_2726,N_2457,N_2539);
xnor U2727 (N_2727,N_2410,N_2514);
xor U2728 (N_2728,N_2485,N_2596);
nand U2729 (N_2729,N_2537,N_2591);
nor U2730 (N_2730,N_2438,N_2498);
and U2731 (N_2731,N_2427,N_2403);
and U2732 (N_2732,N_2573,N_2564);
nand U2733 (N_2733,N_2579,N_2567);
or U2734 (N_2734,N_2539,N_2495);
and U2735 (N_2735,N_2430,N_2521);
or U2736 (N_2736,N_2463,N_2400);
xor U2737 (N_2737,N_2504,N_2448);
xor U2738 (N_2738,N_2572,N_2512);
nor U2739 (N_2739,N_2549,N_2435);
xor U2740 (N_2740,N_2510,N_2414);
or U2741 (N_2741,N_2406,N_2405);
nand U2742 (N_2742,N_2410,N_2598);
xor U2743 (N_2743,N_2502,N_2545);
nand U2744 (N_2744,N_2459,N_2463);
nand U2745 (N_2745,N_2487,N_2479);
nor U2746 (N_2746,N_2517,N_2441);
and U2747 (N_2747,N_2519,N_2565);
and U2748 (N_2748,N_2593,N_2425);
or U2749 (N_2749,N_2423,N_2528);
and U2750 (N_2750,N_2442,N_2469);
xnor U2751 (N_2751,N_2442,N_2467);
nand U2752 (N_2752,N_2495,N_2522);
xor U2753 (N_2753,N_2453,N_2599);
and U2754 (N_2754,N_2562,N_2523);
and U2755 (N_2755,N_2475,N_2506);
xnor U2756 (N_2756,N_2566,N_2591);
nor U2757 (N_2757,N_2508,N_2593);
xnor U2758 (N_2758,N_2497,N_2518);
nor U2759 (N_2759,N_2451,N_2482);
or U2760 (N_2760,N_2403,N_2564);
and U2761 (N_2761,N_2452,N_2462);
nand U2762 (N_2762,N_2461,N_2565);
nor U2763 (N_2763,N_2419,N_2555);
nor U2764 (N_2764,N_2441,N_2466);
nand U2765 (N_2765,N_2477,N_2537);
or U2766 (N_2766,N_2401,N_2476);
or U2767 (N_2767,N_2530,N_2597);
or U2768 (N_2768,N_2460,N_2522);
nand U2769 (N_2769,N_2543,N_2472);
nand U2770 (N_2770,N_2472,N_2563);
nor U2771 (N_2771,N_2520,N_2478);
nor U2772 (N_2772,N_2469,N_2523);
nor U2773 (N_2773,N_2509,N_2413);
or U2774 (N_2774,N_2434,N_2568);
or U2775 (N_2775,N_2575,N_2433);
and U2776 (N_2776,N_2508,N_2518);
or U2777 (N_2777,N_2563,N_2549);
nor U2778 (N_2778,N_2534,N_2586);
xnor U2779 (N_2779,N_2473,N_2449);
nor U2780 (N_2780,N_2432,N_2553);
nor U2781 (N_2781,N_2561,N_2430);
xnor U2782 (N_2782,N_2585,N_2503);
nand U2783 (N_2783,N_2453,N_2455);
xnor U2784 (N_2784,N_2491,N_2563);
nand U2785 (N_2785,N_2571,N_2453);
xnor U2786 (N_2786,N_2523,N_2532);
nand U2787 (N_2787,N_2499,N_2433);
and U2788 (N_2788,N_2440,N_2558);
nand U2789 (N_2789,N_2445,N_2433);
nor U2790 (N_2790,N_2541,N_2556);
xnor U2791 (N_2791,N_2536,N_2594);
nand U2792 (N_2792,N_2410,N_2486);
xnor U2793 (N_2793,N_2449,N_2542);
nor U2794 (N_2794,N_2519,N_2413);
nor U2795 (N_2795,N_2473,N_2563);
and U2796 (N_2796,N_2503,N_2547);
and U2797 (N_2797,N_2595,N_2459);
nor U2798 (N_2798,N_2564,N_2426);
nand U2799 (N_2799,N_2440,N_2437);
nand U2800 (N_2800,N_2624,N_2629);
and U2801 (N_2801,N_2715,N_2781);
xor U2802 (N_2802,N_2708,N_2759);
xnor U2803 (N_2803,N_2681,N_2679);
nand U2804 (N_2804,N_2793,N_2655);
and U2805 (N_2805,N_2642,N_2769);
xnor U2806 (N_2806,N_2664,N_2635);
and U2807 (N_2807,N_2660,N_2620);
xor U2808 (N_2808,N_2745,N_2724);
or U2809 (N_2809,N_2764,N_2782);
nor U2810 (N_2810,N_2658,N_2728);
or U2811 (N_2811,N_2773,N_2630);
or U2812 (N_2812,N_2619,N_2799);
and U2813 (N_2813,N_2657,N_2792);
nor U2814 (N_2814,N_2699,N_2718);
nand U2815 (N_2815,N_2682,N_2632);
and U2816 (N_2816,N_2663,N_2779);
xor U2817 (N_2817,N_2787,N_2711);
and U2818 (N_2818,N_2771,N_2768);
or U2819 (N_2819,N_2694,N_2780);
nor U2820 (N_2820,N_2791,N_2696);
or U2821 (N_2821,N_2680,N_2614);
xnor U2822 (N_2822,N_2601,N_2735);
xor U2823 (N_2823,N_2672,N_2778);
and U2824 (N_2824,N_2637,N_2688);
nor U2825 (N_2825,N_2723,N_2640);
nand U2826 (N_2826,N_2703,N_2650);
nor U2827 (N_2827,N_2713,N_2656);
nor U2828 (N_2828,N_2740,N_2761);
nand U2829 (N_2829,N_2602,N_2751);
xor U2830 (N_2830,N_2727,N_2686);
xor U2831 (N_2831,N_2706,N_2653);
and U2832 (N_2832,N_2754,N_2702);
and U2833 (N_2833,N_2608,N_2704);
and U2834 (N_2834,N_2646,N_2733);
xor U2835 (N_2835,N_2644,N_2670);
nand U2836 (N_2836,N_2692,N_2665);
nand U2837 (N_2837,N_2677,N_2603);
and U2838 (N_2838,N_2638,N_2683);
and U2839 (N_2839,N_2750,N_2641);
nand U2840 (N_2840,N_2742,N_2714);
nor U2841 (N_2841,N_2690,N_2610);
or U2842 (N_2842,N_2676,N_2798);
or U2843 (N_2843,N_2671,N_2693);
nor U2844 (N_2844,N_2760,N_2662);
nor U2845 (N_2845,N_2748,N_2765);
nand U2846 (N_2846,N_2795,N_2772);
nand U2847 (N_2847,N_2776,N_2625);
nor U2848 (N_2848,N_2648,N_2757);
xnor U2849 (N_2849,N_2651,N_2775);
nand U2850 (N_2850,N_2636,N_2721);
nand U2851 (N_2851,N_2719,N_2684);
xor U2852 (N_2852,N_2730,N_2674);
and U2853 (N_2853,N_2732,N_2604);
nand U2854 (N_2854,N_2743,N_2675);
and U2855 (N_2855,N_2678,N_2720);
nor U2856 (N_2856,N_2689,N_2628);
nand U2857 (N_2857,N_2758,N_2726);
nor U2858 (N_2858,N_2729,N_2673);
and U2859 (N_2859,N_2770,N_2607);
or U2860 (N_2860,N_2634,N_2627);
nand U2861 (N_2861,N_2717,N_2788);
xor U2862 (N_2862,N_2701,N_2783);
nand U2863 (N_2863,N_2667,N_2649);
nor U2864 (N_2864,N_2797,N_2777);
nor U2865 (N_2865,N_2767,N_2645);
and U2866 (N_2866,N_2666,N_2616);
or U2867 (N_2867,N_2609,N_2697);
nand U2868 (N_2868,N_2691,N_2774);
nand U2869 (N_2869,N_2739,N_2685);
nor U2870 (N_2870,N_2741,N_2600);
xor U2871 (N_2871,N_2710,N_2606);
nand U2872 (N_2872,N_2762,N_2661);
or U2873 (N_2873,N_2756,N_2639);
xnor U2874 (N_2874,N_2631,N_2613);
nand U2875 (N_2875,N_2709,N_2790);
nand U2876 (N_2876,N_2698,N_2763);
or U2877 (N_2877,N_2789,N_2796);
or U2878 (N_2878,N_2659,N_2695);
xnor U2879 (N_2879,N_2785,N_2734);
and U2880 (N_2880,N_2784,N_2736);
nand U2881 (N_2881,N_2700,N_2652);
nand U2882 (N_2882,N_2617,N_2746);
xnor U2883 (N_2883,N_2786,N_2605);
nand U2884 (N_2884,N_2707,N_2766);
nor U2885 (N_2885,N_2612,N_2731);
nor U2886 (N_2886,N_2626,N_2633);
nor U2887 (N_2887,N_2669,N_2615);
nand U2888 (N_2888,N_2753,N_2712);
nor U2889 (N_2889,N_2737,N_2654);
nand U2890 (N_2890,N_2749,N_2725);
nor U2891 (N_2891,N_2687,N_2647);
xor U2892 (N_2892,N_2618,N_2611);
nor U2893 (N_2893,N_2668,N_2755);
xnor U2894 (N_2894,N_2752,N_2747);
and U2895 (N_2895,N_2716,N_2705);
xor U2896 (N_2896,N_2794,N_2622);
and U2897 (N_2897,N_2722,N_2738);
and U2898 (N_2898,N_2744,N_2623);
and U2899 (N_2899,N_2643,N_2621);
nor U2900 (N_2900,N_2717,N_2720);
or U2901 (N_2901,N_2739,N_2723);
nand U2902 (N_2902,N_2636,N_2701);
and U2903 (N_2903,N_2660,N_2773);
xnor U2904 (N_2904,N_2745,N_2600);
nand U2905 (N_2905,N_2748,N_2674);
xor U2906 (N_2906,N_2621,N_2684);
nor U2907 (N_2907,N_2766,N_2614);
xor U2908 (N_2908,N_2739,N_2766);
and U2909 (N_2909,N_2696,N_2705);
or U2910 (N_2910,N_2612,N_2649);
nand U2911 (N_2911,N_2657,N_2696);
xor U2912 (N_2912,N_2651,N_2690);
or U2913 (N_2913,N_2737,N_2682);
and U2914 (N_2914,N_2631,N_2694);
xor U2915 (N_2915,N_2637,N_2728);
and U2916 (N_2916,N_2758,N_2696);
nand U2917 (N_2917,N_2721,N_2629);
and U2918 (N_2918,N_2772,N_2610);
and U2919 (N_2919,N_2758,N_2740);
xor U2920 (N_2920,N_2717,N_2766);
nor U2921 (N_2921,N_2656,N_2720);
or U2922 (N_2922,N_2777,N_2725);
and U2923 (N_2923,N_2621,N_2733);
and U2924 (N_2924,N_2645,N_2741);
nand U2925 (N_2925,N_2624,N_2744);
and U2926 (N_2926,N_2707,N_2751);
nor U2927 (N_2927,N_2758,N_2755);
and U2928 (N_2928,N_2750,N_2716);
xnor U2929 (N_2929,N_2716,N_2621);
xnor U2930 (N_2930,N_2649,N_2647);
xor U2931 (N_2931,N_2664,N_2652);
nand U2932 (N_2932,N_2668,N_2748);
nand U2933 (N_2933,N_2753,N_2760);
nor U2934 (N_2934,N_2726,N_2606);
nand U2935 (N_2935,N_2648,N_2742);
xnor U2936 (N_2936,N_2613,N_2748);
nor U2937 (N_2937,N_2766,N_2632);
xor U2938 (N_2938,N_2709,N_2637);
nor U2939 (N_2939,N_2614,N_2687);
xor U2940 (N_2940,N_2672,N_2683);
or U2941 (N_2941,N_2739,N_2640);
or U2942 (N_2942,N_2785,N_2771);
xor U2943 (N_2943,N_2779,N_2772);
and U2944 (N_2944,N_2715,N_2729);
and U2945 (N_2945,N_2606,N_2612);
or U2946 (N_2946,N_2684,N_2643);
xnor U2947 (N_2947,N_2793,N_2736);
nand U2948 (N_2948,N_2611,N_2733);
or U2949 (N_2949,N_2726,N_2689);
and U2950 (N_2950,N_2765,N_2726);
nor U2951 (N_2951,N_2741,N_2729);
and U2952 (N_2952,N_2754,N_2651);
xor U2953 (N_2953,N_2757,N_2784);
nor U2954 (N_2954,N_2738,N_2712);
nand U2955 (N_2955,N_2795,N_2784);
nor U2956 (N_2956,N_2608,N_2617);
nor U2957 (N_2957,N_2626,N_2781);
or U2958 (N_2958,N_2626,N_2638);
and U2959 (N_2959,N_2610,N_2640);
and U2960 (N_2960,N_2674,N_2773);
nor U2961 (N_2961,N_2637,N_2773);
nand U2962 (N_2962,N_2720,N_2602);
nor U2963 (N_2963,N_2693,N_2710);
nor U2964 (N_2964,N_2703,N_2614);
nand U2965 (N_2965,N_2637,N_2699);
and U2966 (N_2966,N_2625,N_2760);
or U2967 (N_2967,N_2698,N_2685);
nor U2968 (N_2968,N_2750,N_2721);
xnor U2969 (N_2969,N_2702,N_2751);
nand U2970 (N_2970,N_2729,N_2762);
and U2971 (N_2971,N_2607,N_2602);
nor U2972 (N_2972,N_2795,N_2641);
nor U2973 (N_2973,N_2679,N_2643);
xor U2974 (N_2974,N_2764,N_2699);
and U2975 (N_2975,N_2688,N_2671);
and U2976 (N_2976,N_2759,N_2715);
or U2977 (N_2977,N_2729,N_2681);
xnor U2978 (N_2978,N_2764,N_2703);
and U2979 (N_2979,N_2694,N_2719);
nand U2980 (N_2980,N_2621,N_2607);
nand U2981 (N_2981,N_2798,N_2651);
nor U2982 (N_2982,N_2601,N_2665);
or U2983 (N_2983,N_2773,N_2638);
xnor U2984 (N_2984,N_2697,N_2781);
and U2985 (N_2985,N_2710,N_2748);
and U2986 (N_2986,N_2798,N_2613);
xor U2987 (N_2987,N_2785,N_2671);
xnor U2988 (N_2988,N_2695,N_2665);
xor U2989 (N_2989,N_2708,N_2628);
nand U2990 (N_2990,N_2779,N_2661);
and U2991 (N_2991,N_2744,N_2751);
or U2992 (N_2992,N_2611,N_2660);
xnor U2993 (N_2993,N_2613,N_2780);
xor U2994 (N_2994,N_2781,N_2640);
xor U2995 (N_2995,N_2773,N_2677);
xor U2996 (N_2996,N_2623,N_2705);
xor U2997 (N_2997,N_2676,N_2682);
nand U2998 (N_2998,N_2713,N_2658);
xor U2999 (N_2999,N_2677,N_2606);
or U3000 (N_3000,N_2846,N_2919);
nand U3001 (N_3001,N_2820,N_2824);
and U3002 (N_3002,N_2883,N_2922);
or U3003 (N_3003,N_2897,N_2810);
and U3004 (N_3004,N_2925,N_2985);
or U3005 (N_3005,N_2839,N_2943);
nand U3006 (N_3006,N_2944,N_2869);
nor U3007 (N_3007,N_2804,N_2859);
xnor U3008 (N_3008,N_2989,N_2923);
and U3009 (N_3009,N_2902,N_2888);
and U3010 (N_3010,N_2990,N_2834);
or U3011 (N_3011,N_2930,N_2849);
nand U3012 (N_3012,N_2837,N_2952);
nand U3013 (N_3013,N_2965,N_2968);
nor U3014 (N_3014,N_2874,N_2958);
nand U3015 (N_3015,N_2953,N_2949);
or U3016 (N_3016,N_2871,N_2962);
nand U3017 (N_3017,N_2969,N_2867);
nand U3018 (N_3018,N_2893,N_2833);
xnor U3019 (N_3019,N_2911,N_2811);
and U3020 (N_3020,N_2948,N_2827);
and U3021 (N_3021,N_2979,N_2817);
nand U3022 (N_3022,N_2964,N_2939);
or U3023 (N_3023,N_2987,N_2975);
xor U3024 (N_3024,N_2894,N_2860);
xor U3025 (N_3025,N_2994,N_2908);
or U3026 (N_3026,N_2829,N_2855);
xnor U3027 (N_3027,N_2899,N_2864);
nor U3028 (N_3028,N_2933,N_2854);
and U3029 (N_3029,N_2870,N_2805);
and U3030 (N_3030,N_2848,N_2938);
nor U3031 (N_3031,N_2887,N_2844);
or U3032 (N_3032,N_2845,N_2928);
nor U3033 (N_3033,N_2977,N_2889);
nand U3034 (N_3034,N_2957,N_2835);
nor U3035 (N_3035,N_2880,N_2921);
and U3036 (N_3036,N_2997,N_2822);
and U3037 (N_3037,N_2896,N_2825);
nand U3038 (N_3038,N_2882,N_2950);
xor U3039 (N_3039,N_2927,N_2981);
or U3040 (N_3040,N_2912,N_2879);
nor U3041 (N_3041,N_2826,N_2856);
and U3042 (N_3042,N_2838,N_2935);
or U3043 (N_3043,N_2976,N_2967);
or U3044 (N_3044,N_2842,N_2830);
or U3045 (N_3045,N_2906,N_2926);
or U3046 (N_3046,N_2904,N_2821);
xnor U3047 (N_3047,N_2861,N_2993);
nand U3048 (N_3048,N_2914,N_2918);
or U3049 (N_3049,N_2900,N_2818);
or U3050 (N_3050,N_2801,N_2951);
nor U3051 (N_3051,N_2960,N_2988);
nand U3052 (N_3052,N_2823,N_2892);
or U3053 (N_3053,N_2812,N_2998);
xnor U3054 (N_3054,N_2966,N_2866);
nor U3055 (N_3055,N_2913,N_2907);
xnor U3056 (N_3056,N_2999,N_2898);
or U3057 (N_3057,N_2932,N_2991);
and U3058 (N_3058,N_2862,N_2831);
and U3059 (N_3059,N_2802,N_2857);
or U3060 (N_3060,N_2982,N_2929);
or U3061 (N_3061,N_2901,N_2800);
nor U3062 (N_3062,N_2876,N_2995);
or U3063 (N_3063,N_2885,N_2836);
xnor U3064 (N_3064,N_2905,N_2963);
nand U3065 (N_3065,N_2891,N_2881);
nor U3066 (N_3066,N_2910,N_2946);
or U3067 (N_3067,N_2947,N_2890);
xor U3068 (N_3068,N_2852,N_2983);
and U3069 (N_3069,N_2940,N_2974);
nor U3070 (N_3070,N_2814,N_2850);
and U3071 (N_3071,N_2813,N_2984);
or U3072 (N_3072,N_2954,N_2956);
nor U3073 (N_3073,N_2819,N_2808);
xnor U3074 (N_3074,N_2816,N_2865);
nand U3075 (N_3075,N_2916,N_2955);
and U3076 (N_3076,N_2959,N_2941);
xor U3077 (N_3077,N_2872,N_2992);
nand U3078 (N_3078,N_2843,N_2895);
nand U3079 (N_3079,N_2873,N_2971);
nand U3080 (N_3080,N_2936,N_2858);
nor U3081 (N_3081,N_2934,N_2840);
nor U3082 (N_3082,N_2945,N_2973);
or U3083 (N_3083,N_2903,N_2875);
nand U3084 (N_3084,N_2970,N_2868);
or U3085 (N_3085,N_2917,N_2807);
nand U3086 (N_3086,N_2972,N_2986);
or U3087 (N_3087,N_2851,N_2884);
xor U3088 (N_3088,N_2806,N_2847);
nand U3089 (N_3089,N_2915,N_2853);
xor U3090 (N_3090,N_2877,N_2996);
nor U3091 (N_3091,N_2931,N_2920);
or U3092 (N_3092,N_2909,N_2832);
nor U3093 (N_3093,N_2828,N_2815);
nand U3094 (N_3094,N_2961,N_2978);
xnor U3095 (N_3095,N_2924,N_2878);
nor U3096 (N_3096,N_2980,N_2886);
and U3097 (N_3097,N_2841,N_2809);
nand U3098 (N_3098,N_2942,N_2937);
or U3099 (N_3099,N_2863,N_2803);
xor U3100 (N_3100,N_2844,N_2948);
and U3101 (N_3101,N_2966,N_2939);
xnor U3102 (N_3102,N_2843,N_2897);
or U3103 (N_3103,N_2866,N_2876);
or U3104 (N_3104,N_2937,N_2871);
xor U3105 (N_3105,N_2914,N_2944);
or U3106 (N_3106,N_2961,N_2959);
and U3107 (N_3107,N_2996,N_2830);
or U3108 (N_3108,N_2997,N_2858);
or U3109 (N_3109,N_2976,N_2996);
nand U3110 (N_3110,N_2945,N_2960);
and U3111 (N_3111,N_2932,N_2948);
nor U3112 (N_3112,N_2953,N_2979);
xnor U3113 (N_3113,N_2943,N_2949);
or U3114 (N_3114,N_2883,N_2942);
nand U3115 (N_3115,N_2879,N_2963);
or U3116 (N_3116,N_2915,N_2926);
and U3117 (N_3117,N_2802,N_2804);
or U3118 (N_3118,N_2997,N_2893);
and U3119 (N_3119,N_2811,N_2827);
xnor U3120 (N_3120,N_2907,N_2908);
nor U3121 (N_3121,N_2864,N_2942);
or U3122 (N_3122,N_2817,N_2997);
xnor U3123 (N_3123,N_2996,N_2890);
xor U3124 (N_3124,N_2840,N_2857);
nor U3125 (N_3125,N_2892,N_2927);
and U3126 (N_3126,N_2830,N_2875);
nand U3127 (N_3127,N_2810,N_2961);
and U3128 (N_3128,N_2811,N_2898);
nor U3129 (N_3129,N_2946,N_2862);
nand U3130 (N_3130,N_2882,N_2801);
nand U3131 (N_3131,N_2861,N_2838);
nand U3132 (N_3132,N_2996,N_2949);
nand U3133 (N_3133,N_2957,N_2926);
and U3134 (N_3134,N_2923,N_2983);
and U3135 (N_3135,N_2895,N_2917);
and U3136 (N_3136,N_2859,N_2985);
nor U3137 (N_3137,N_2964,N_2973);
or U3138 (N_3138,N_2940,N_2945);
nand U3139 (N_3139,N_2917,N_2956);
and U3140 (N_3140,N_2834,N_2876);
and U3141 (N_3141,N_2926,N_2986);
nor U3142 (N_3142,N_2942,N_2826);
xnor U3143 (N_3143,N_2881,N_2824);
nand U3144 (N_3144,N_2914,N_2814);
xor U3145 (N_3145,N_2804,N_2902);
nand U3146 (N_3146,N_2954,N_2951);
and U3147 (N_3147,N_2937,N_2997);
and U3148 (N_3148,N_2931,N_2826);
nand U3149 (N_3149,N_2881,N_2849);
xnor U3150 (N_3150,N_2842,N_2862);
or U3151 (N_3151,N_2847,N_2989);
xnor U3152 (N_3152,N_2956,N_2873);
and U3153 (N_3153,N_2912,N_2869);
nor U3154 (N_3154,N_2933,N_2831);
or U3155 (N_3155,N_2852,N_2892);
or U3156 (N_3156,N_2858,N_2911);
nand U3157 (N_3157,N_2950,N_2896);
xnor U3158 (N_3158,N_2990,N_2882);
and U3159 (N_3159,N_2899,N_2971);
or U3160 (N_3160,N_2903,N_2814);
or U3161 (N_3161,N_2960,N_2981);
xnor U3162 (N_3162,N_2805,N_2887);
or U3163 (N_3163,N_2904,N_2910);
and U3164 (N_3164,N_2856,N_2832);
nand U3165 (N_3165,N_2801,N_2865);
or U3166 (N_3166,N_2840,N_2973);
xor U3167 (N_3167,N_2922,N_2995);
nand U3168 (N_3168,N_2933,N_2945);
nand U3169 (N_3169,N_2969,N_2854);
and U3170 (N_3170,N_2932,N_2997);
nand U3171 (N_3171,N_2933,N_2825);
xor U3172 (N_3172,N_2923,N_2934);
or U3173 (N_3173,N_2804,N_2831);
and U3174 (N_3174,N_2915,N_2955);
or U3175 (N_3175,N_2859,N_2838);
nor U3176 (N_3176,N_2944,N_2950);
nand U3177 (N_3177,N_2976,N_2964);
and U3178 (N_3178,N_2955,N_2919);
nand U3179 (N_3179,N_2965,N_2842);
or U3180 (N_3180,N_2927,N_2953);
xor U3181 (N_3181,N_2926,N_2817);
nand U3182 (N_3182,N_2854,N_2849);
nor U3183 (N_3183,N_2832,N_2838);
and U3184 (N_3184,N_2957,N_2853);
and U3185 (N_3185,N_2988,N_2951);
xor U3186 (N_3186,N_2853,N_2916);
nor U3187 (N_3187,N_2979,N_2970);
xnor U3188 (N_3188,N_2951,N_2879);
nor U3189 (N_3189,N_2855,N_2948);
nand U3190 (N_3190,N_2891,N_2906);
or U3191 (N_3191,N_2812,N_2906);
nor U3192 (N_3192,N_2858,N_2806);
or U3193 (N_3193,N_2911,N_2898);
nand U3194 (N_3194,N_2883,N_2839);
and U3195 (N_3195,N_2822,N_2887);
or U3196 (N_3196,N_2871,N_2939);
nor U3197 (N_3197,N_2803,N_2853);
nor U3198 (N_3198,N_2927,N_2950);
or U3199 (N_3199,N_2976,N_2956);
nor U3200 (N_3200,N_3160,N_3082);
and U3201 (N_3201,N_3198,N_3013);
nor U3202 (N_3202,N_3076,N_3021);
or U3203 (N_3203,N_3107,N_3025);
nor U3204 (N_3204,N_3079,N_3156);
and U3205 (N_3205,N_3129,N_3031);
nor U3206 (N_3206,N_3086,N_3091);
or U3207 (N_3207,N_3078,N_3012);
and U3208 (N_3208,N_3149,N_3102);
nor U3209 (N_3209,N_3023,N_3015);
and U3210 (N_3210,N_3118,N_3033);
xor U3211 (N_3211,N_3074,N_3037);
and U3212 (N_3212,N_3081,N_3043);
nor U3213 (N_3213,N_3073,N_3057);
nand U3214 (N_3214,N_3194,N_3159);
and U3215 (N_3215,N_3008,N_3070);
nor U3216 (N_3216,N_3146,N_3111);
xnor U3217 (N_3217,N_3117,N_3121);
xnor U3218 (N_3218,N_3109,N_3032);
xnor U3219 (N_3219,N_3143,N_3084);
xor U3220 (N_3220,N_3014,N_3132);
and U3221 (N_3221,N_3191,N_3182);
xnor U3222 (N_3222,N_3113,N_3016);
or U3223 (N_3223,N_3150,N_3062);
nand U3224 (N_3224,N_3034,N_3048);
nor U3225 (N_3225,N_3166,N_3155);
nor U3226 (N_3226,N_3036,N_3180);
nor U3227 (N_3227,N_3099,N_3060);
or U3228 (N_3228,N_3069,N_3197);
xnor U3229 (N_3229,N_3001,N_3046);
or U3230 (N_3230,N_3105,N_3085);
nand U3231 (N_3231,N_3067,N_3050);
nand U3232 (N_3232,N_3126,N_3135);
xor U3233 (N_3233,N_3110,N_3130);
nand U3234 (N_3234,N_3190,N_3028);
and U3235 (N_3235,N_3186,N_3038);
nor U3236 (N_3236,N_3176,N_3195);
xnor U3237 (N_3237,N_3145,N_3140);
nor U3238 (N_3238,N_3196,N_3175);
nand U3239 (N_3239,N_3122,N_3125);
nor U3240 (N_3240,N_3047,N_3088);
nand U3241 (N_3241,N_3040,N_3051);
nand U3242 (N_3242,N_3128,N_3171);
and U3243 (N_3243,N_3096,N_3167);
or U3244 (N_3244,N_3127,N_3178);
and U3245 (N_3245,N_3007,N_3018);
nand U3246 (N_3246,N_3049,N_3000);
and U3247 (N_3247,N_3041,N_3030);
nor U3248 (N_3248,N_3147,N_3170);
and U3249 (N_3249,N_3002,N_3089);
nand U3250 (N_3250,N_3029,N_3172);
xor U3251 (N_3251,N_3095,N_3045);
nor U3252 (N_3252,N_3063,N_3154);
and U3253 (N_3253,N_3164,N_3024);
nor U3254 (N_3254,N_3192,N_3093);
or U3255 (N_3255,N_3183,N_3003);
nor U3256 (N_3256,N_3071,N_3022);
and U3257 (N_3257,N_3061,N_3065);
nand U3258 (N_3258,N_3165,N_3112);
nor U3259 (N_3259,N_3177,N_3056);
nor U3260 (N_3260,N_3148,N_3052);
or U3261 (N_3261,N_3035,N_3068);
and U3262 (N_3262,N_3199,N_3158);
or U3263 (N_3263,N_3054,N_3027);
and U3264 (N_3264,N_3185,N_3142);
nor U3265 (N_3265,N_3004,N_3098);
nor U3266 (N_3266,N_3162,N_3020);
nor U3267 (N_3267,N_3169,N_3100);
nand U3268 (N_3268,N_3077,N_3136);
nand U3269 (N_3269,N_3153,N_3131);
and U3270 (N_3270,N_3101,N_3174);
xnor U3271 (N_3271,N_3179,N_3087);
and U3272 (N_3272,N_3075,N_3124);
or U3273 (N_3273,N_3173,N_3053);
nand U3274 (N_3274,N_3161,N_3103);
nor U3275 (N_3275,N_3092,N_3116);
xnor U3276 (N_3276,N_3066,N_3184);
or U3277 (N_3277,N_3083,N_3157);
nand U3278 (N_3278,N_3044,N_3163);
and U3279 (N_3279,N_3139,N_3017);
and U3280 (N_3280,N_3151,N_3090);
xnor U3281 (N_3281,N_3108,N_3039);
xnor U3282 (N_3282,N_3042,N_3106);
nor U3283 (N_3283,N_3123,N_3152);
nor U3284 (N_3284,N_3104,N_3188);
and U3285 (N_3285,N_3114,N_3138);
and U3286 (N_3286,N_3137,N_3094);
or U3287 (N_3287,N_3010,N_3187);
and U3288 (N_3288,N_3120,N_3141);
xnor U3289 (N_3289,N_3009,N_3181);
nor U3290 (N_3290,N_3005,N_3058);
nand U3291 (N_3291,N_3133,N_3072);
or U3292 (N_3292,N_3119,N_3097);
nor U3293 (N_3293,N_3080,N_3011);
xnor U3294 (N_3294,N_3019,N_3193);
xnor U3295 (N_3295,N_3115,N_3144);
or U3296 (N_3296,N_3006,N_3189);
nor U3297 (N_3297,N_3134,N_3064);
and U3298 (N_3298,N_3168,N_3059);
nand U3299 (N_3299,N_3055,N_3026);
nand U3300 (N_3300,N_3085,N_3192);
or U3301 (N_3301,N_3194,N_3037);
or U3302 (N_3302,N_3114,N_3097);
nor U3303 (N_3303,N_3193,N_3014);
xnor U3304 (N_3304,N_3115,N_3160);
or U3305 (N_3305,N_3048,N_3191);
nand U3306 (N_3306,N_3145,N_3060);
xnor U3307 (N_3307,N_3010,N_3018);
and U3308 (N_3308,N_3134,N_3001);
xor U3309 (N_3309,N_3170,N_3023);
nand U3310 (N_3310,N_3129,N_3051);
or U3311 (N_3311,N_3185,N_3113);
and U3312 (N_3312,N_3044,N_3115);
nor U3313 (N_3313,N_3150,N_3191);
or U3314 (N_3314,N_3166,N_3161);
nor U3315 (N_3315,N_3013,N_3099);
xnor U3316 (N_3316,N_3135,N_3032);
nand U3317 (N_3317,N_3115,N_3159);
xnor U3318 (N_3318,N_3009,N_3169);
nor U3319 (N_3319,N_3084,N_3112);
nand U3320 (N_3320,N_3101,N_3016);
or U3321 (N_3321,N_3167,N_3038);
nor U3322 (N_3322,N_3050,N_3008);
or U3323 (N_3323,N_3038,N_3126);
nand U3324 (N_3324,N_3083,N_3190);
or U3325 (N_3325,N_3094,N_3065);
xnor U3326 (N_3326,N_3098,N_3144);
xor U3327 (N_3327,N_3081,N_3029);
nand U3328 (N_3328,N_3137,N_3013);
nand U3329 (N_3329,N_3187,N_3122);
nor U3330 (N_3330,N_3023,N_3064);
xnor U3331 (N_3331,N_3089,N_3147);
or U3332 (N_3332,N_3098,N_3052);
nor U3333 (N_3333,N_3152,N_3156);
xor U3334 (N_3334,N_3195,N_3001);
and U3335 (N_3335,N_3140,N_3046);
nor U3336 (N_3336,N_3171,N_3129);
and U3337 (N_3337,N_3101,N_3031);
or U3338 (N_3338,N_3179,N_3190);
nor U3339 (N_3339,N_3180,N_3178);
or U3340 (N_3340,N_3057,N_3053);
nor U3341 (N_3341,N_3098,N_3110);
nor U3342 (N_3342,N_3046,N_3048);
and U3343 (N_3343,N_3182,N_3099);
and U3344 (N_3344,N_3139,N_3141);
and U3345 (N_3345,N_3005,N_3075);
nor U3346 (N_3346,N_3170,N_3117);
or U3347 (N_3347,N_3094,N_3124);
nor U3348 (N_3348,N_3155,N_3078);
nand U3349 (N_3349,N_3089,N_3111);
nor U3350 (N_3350,N_3005,N_3140);
xor U3351 (N_3351,N_3044,N_3095);
nor U3352 (N_3352,N_3029,N_3025);
nand U3353 (N_3353,N_3100,N_3178);
nand U3354 (N_3354,N_3060,N_3022);
xnor U3355 (N_3355,N_3105,N_3106);
and U3356 (N_3356,N_3046,N_3114);
nor U3357 (N_3357,N_3008,N_3098);
xor U3358 (N_3358,N_3110,N_3129);
and U3359 (N_3359,N_3003,N_3069);
nor U3360 (N_3360,N_3164,N_3048);
nor U3361 (N_3361,N_3169,N_3061);
nor U3362 (N_3362,N_3059,N_3056);
nor U3363 (N_3363,N_3006,N_3101);
xor U3364 (N_3364,N_3039,N_3170);
xor U3365 (N_3365,N_3001,N_3038);
nand U3366 (N_3366,N_3035,N_3055);
or U3367 (N_3367,N_3002,N_3111);
nand U3368 (N_3368,N_3130,N_3196);
and U3369 (N_3369,N_3142,N_3051);
and U3370 (N_3370,N_3099,N_3118);
and U3371 (N_3371,N_3147,N_3112);
xor U3372 (N_3372,N_3086,N_3126);
or U3373 (N_3373,N_3034,N_3073);
or U3374 (N_3374,N_3133,N_3046);
and U3375 (N_3375,N_3051,N_3089);
xor U3376 (N_3376,N_3147,N_3067);
and U3377 (N_3377,N_3117,N_3089);
xor U3378 (N_3378,N_3175,N_3168);
xor U3379 (N_3379,N_3137,N_3177);
xnor U3380 (N_3380,N_3100,N_3180);
nand U3381 (N_3381,N_3096,N_3023);
or U3382 (N_3382,N_3194,N_3056);
and U3383 (N_3383,N_3128,N_3077);
and U3384 (N_3384,N_3010,N_3046);
nor U3385 (N_3385,N_3182,N_3183);
or U3386 (N_3386,N_3076,N_3036);
nor U3387 (N_3387,N_3009,N_3013);
xor U3388 (N_3388,N_3196,N_3042);
or U3389 (N_3389,N_3057,N_3090);
xor U3390 (N_3390,N_3029,N_3032);
nor U3391 (N_3391,N_3079,N_3171);
and U3392 (N_3392,N_3018,N_3016);
xnor U3393 (N_3393,N_3098,N_3122);
nor U3394 (N_3394,N_3089,N_3049);
xnor U3395 (N_3395,N_3047,N_3074);
and U3396 (N_3396,N_3005,N_3116);
and U3397 (N_3397,N_3100,N_3145);
and U3398 (N_3398,N_3143,N_3024);
nand U3399 (N_3399,N_3096,N_3194);
nand U3400 (N_3400,N_3313,N_3326);
or U3401 (N_3401,N_3301,N_3303);
nor U3402 (N_3402,N_3357,N_3248);
nor U3403 (N_3403,N_3293,N_3335);
or U3404 (N_3404,N_3224,N_3352);
xor U3405 (N_3405,N_3306,N_3383);
xnor U3406 (N_3406,N_3289,N_3251);
xor U3407 (N_3407,N_3279,N_3286);
or U3408 (N_3408,N_3377,N_3360);
nor U3409 (N_3409,N_3356,N_3227);
or U3410 (N_3410,N_3317,N_3380);
xor U3411 (N_3411,N_3259,N_3372);
or U3412 (N_3412,N_3222,N_3237);
xor U3413 (N_3413,N_3294,N_3217);
nand U3414 (N_3414,N_3260,N_3391);
and U3415 (N_3415,N_3275,N_3327);
nand U3416 (N_3416,N_3291,N_3340);
or U3417 (N_3417,N_3263,N_3284);
nor U3418 (N_3418,N_3334,N_3280);
or U3419 (N_3419,N_3220,N_3239);
and U3420 (N_3420,N_3201,N_3389);
or U3421 (N_3421,N_3381,N_3349);
or U3422 (N_3422,N_3249,N_3320);
and U3423 (N_3423,N_3242,N_3244);
nand U3424 (N_3424,N_3221,N_3304);
and U3425 (N_3425,N_3385,N_3392);
nor U3426 (N_3426,N_3281,N_3209);
nor U3427 (N_3427,N_3319,N_3394);
and U3428 (N_3428,N_3228,N_3374);
nand U3429 (N_3429,N_3210,N_3332);
xnor U3430 (N_3430,N_3364,N_3252);
xor U3431 (N_3431,N_3225,N_3328);
and U3432 (N_3432,N_3215,N_3343);
nand U3433 (N_3433,N_3367,N_3316);
nand U3434 (N_3434,N_3308,N_3370);
nand U3435 (N_3435,N_3287,N_3321);
nand U3436 (N_3436,N_3322,N_3393);
or U3437 (N_3437,N_3229,N_3363);
nand U3438 (N_3438,N_3331,N_3231);
nor U3439 (N_3439,N_3246,N_3254);
and U3440 (N_3440,N_3345,N_3366);
nand U3441 (N_3441,N_3307,N_3212);
nand U3442 (N_3442,N_3230,N_3346);
and U3443 (N_3443,N_3213,N_3205);
nor U3444 (N_3444,N_3208,N_3368);
nor U3445 (N_3445,N_3271,N_3395);
and U3446 (N_3446,N_3333,N_3302);
and U3447 (N_3447,N_3298,N_3398);
nor U3448 (N_3448,N_3247,N_3348);
and U3449 (N_3449,N_3369,N_3314);
or U3450 (N_3450,N_3270,N_3351);
nor U3451 (N_3451,N_3382,N_3347);
xor U3452 (N_3452,N_3329,N_3255);
nor U3453 (N_3453,N_3354,N_3310);
xor U3454 (N_3454,N_3226,N_3300);
nand U3455 (N_3455,N_3365,N_3267);
xor U3456 (N_3456,N_3214,N_3223);
nor U3457 (N_3457,N_3337,N_3324);
nand U3458 (N_3458,N_3203,N_3243);
nor U3459 (N_3459,N_3297,N_3236);
nand U3460 (N_3460,N_3384,N_3305);
nand U3461 (N_3461,N_3344,N_3283);
xnor U3462 (N_3462,N_3218,N_3268);
and U3463 (N_3463,N_3387,N_3375);
nor U3464 (N_3464,N_3350,N_3202);
xnor U3465 (N_3465,N_3261,N_3257);
xor U3466 (N_3466,N_3362,N_3399);
and U3467 (N_3467,N_3342,N_3318);
and U3468 (N_3468,N_3200,N_3378);
xnor U3469 (N_3469,N_3341,N_3386);
nand U3470 (N_3470,N_3336,N_3204);
xnor U3471 (N_3471,N_3250,N_3296);
or U3472 (N_3472,N_3312,N_3376);
nand U3473 (N_3473,N_3330,N_3258);
and U3474 (N_3474,N_3273,N_3265);
nand U3475 (N_3475,N_3299,N_3233);
and U3476 (N_3476,N_3234,N_3216);
nor U3477 (N_3477,N_3276,N_3256);
or U3478 (N_3478,N_3272,N_3355);
xnor U3479 (N_3479,N_3361,N_3338);
nand U3480 (N_3480,N_3253,N_3245);
xor U3481 (N_3481,N_3207,N_3397);
or U3482 (N_3482,N_3371,N_3323);
xnor U3483 (N_3483,N_3325,N_3358);
xor U3484 (N_3484,N_3288,N_3262);
xnor U3485 (N_3485,N_3388,N_3359);
and U3486 (N_3486,N_3390,N_3278);
or U3487 (N_3487,N_3396,N_3295);
or U3488 (N_3488,N_3311,N_3315);
nor U3489 (N_3489,N_3373,N_3269);
xor U3490 (N_3490,N_3339,N_3292);
xor U3491 (N_3491,N_3232,N_3274);
and U3492 (N_3492,N_3238,N_3379);
nand U3493 (N_3493,N_3309,N_3235);
nor U3494 (N_3494,N_3211,N_3219);
nor U3495 (N_3495,N_3277,N_3353);
and U3496 (N_3496,N_3264,N_3240);
or U3497 (N_3497,N_3290,N_3241);
and U3498 (N_3498,N_3282,N_3266);
nor U3499 (N_3499,N_3285,N_3206);
nor U3500 (N_3500,N_3224,N_3338);
or U3501 (N_3501,N_3338,N_3295);
or U3502 (N_3502,N_3250,N_3266);
and U3503 (N_3503,N_3315,N_3345);
nor U3504 (N_3504,N_3229,N_3384);
nor U3505 (N_3505,N_3397,N_3370);
or U3506 (N_3506,N_3327,N_3361);
nand U3507 (N_3507,N_3362,N_3227);
nor U3508 (N_3508,N_3249,N_3391);
xor U3509 (N_3509,N_3315,N_3385);
or U3510 (N_3510,N_3278,N_3221);
nor U3511 (N_3511,N_3354,N_3381);
and U3512 (N_3512,N_3372,N_3269);
and U3513 (N_3513,N_3317,N_3345);
xor U3514 (N_3514,N_3304,N_3389);
xor U3515 (N_3515,N_3263,N_3314);
xor U3516 (N_3516,N_3218,N_3228);
nand U3517 (N_3517,N_3282,N_3364);
xor U3518 (N_3518,N_3278,N_3276);
nor U3519 (N_3519,N_3283,N_3374);
xnor U3520 (N_3520,N_3361,N_3270);
nor U3521 (N_3521,N_3234,N_3398);
nor U3522 (N_3522,N_3298,N_3218);
xnor U3523 (N_3523,N_3217,N_3214);
nand U3524 (N_3524,N_3374,N_3244);
nor U3525 (N_3525,N_3201,N_3214);
nand U3526 (N_3526,N_3386,N_3259);
nor U3527 (N_3527,N_3314,N_3242);
and U3528 (N_3528,N_3383,N_3235);
and U3529 (N_3529,N_3324,N_3359);
xor U3530 (N_3530,N_3206,N_3332);
nor U3531 (N_3531,N_3264,N_3389);
and U3532 (N_3532,N_3356,N_3214);
xnor U3533 (N_3533,N_3334,N_3270);
xnor U3534 (N_3534,N_3317,N_3202);
nor U3535 (N_3535,N_3380,N_3308);
xor U3536 (N_3536,N_3242,N_3325);
and U3537 (N_3537,N_3282,N_3269);
nand U3538 (N_3538,N_3285,N_3304);
and U3539 (N_3539,N_3209,N_3254);
nand U3540 (N_3540,N_3333,N_3326);
nand U3541 (N_3541,N_3363,N_3399);
nor U3542 (N_3542,N_3241,N_3272);
and U3543 (N_3543,N_3278,N_3333);
nand U3544 (N_3544,N_3298,N_3365);
nand U3545 (N_3545,N_3360,N_3286);
nor U3546 (N_3546,N_3229,N_3365);
nand U3547 (N_3547,N_3214,N_3312);
xnor U3548 (N_3548,N_3386,N_3330);
and U3549 (N_3549,N_3227,N_3256);
or U3550 (N_3550,N_3386,N_3318);
xor U3551 (N_3551,N_3266,N_3374);
nand U3552 (N_3552,N_3238,N_3322);
and U3553 (N_3553,N_3288,N_3351);
nand U3554 (N_3554,N_3324,N_3301);
or U3555 (N_3555,N_3372,N_3309);
and U3556 (N_3556,N_3375,N_3216);
and U3557 (N_3557,N_3311,N_3346);
nor U3558 (N_3558,N_3347,N_3264);
nand U3559 (N_3559,N_3385,N_3396);
xnor U3560 (N_3560,N_3228,N_3369);
and U3561 (N_3561,N_3335,N_3392);
nor U3562 (N_3562,N_3328,N_3352);
or U3563 (N_3563,N_3347,N_3359);
xnor U3564 (N_3564,N_3235,N_3343);
and U3565 (N_3565,N_3258,N_3277);
or U3566 (N_3566,N_3281,N_3261);
and U3567 (N_3567,N_3224,N_3205);
nor U3568 (N_3568,N_3283,N_3288);
and U3569 (N_3569,N_3203,N_3328);
xor U3570 (N_3570,N_3308,N_3353);
xor U3571 (N_3571,N_3225,N_3394);
nor U3572 (N_3572,N_3340,N_3279);
nor U3573 (N_3573,N_3323,N_3200);
nor U3574 (N_3574,N_3399,N_3381);
or U3575 (N_3575,N_3279,N_3216);
or U3576 (N_3576,N_3279,N_3382);
xnor U3577 (N_3577,N_3274,N_3253);
or U3578 (N_3578,N_3348,N_3340);
or U3579 (N_3579,N_3288,N_3325);
and U3580 (N_3580,N_3392,N_3345);
or U3581 (N_3581,N_3251,N_3327);
and U3582 (N_3582,N_3315,N_3317);
xnor U3583 (N_3583,N_3362,N_3285);
nor U3584 (N_3584,N_3348,N_3305);
nand U3585 (N_3585,N_3352,N_3272);
and U3586 (N_3586,N_3368,N_3335);
or U3587 (N_3587,N_3273,N_3282);
and U3588 (N_3588,N_3288,N_3238);
nand U3589 (N_3589,N_3317,N_3265);
nor U3590 (N_3590,N_3262,N_3372);
and U3591 (N_3591,N_3395,N_3205);
nor U3592 (N_3592,N_3325,N_3359);
and U3593 (N_3593,N_3254,N_3284);
nor U3594 (N_3594,N_3275,N_3288);
nand U3595 (N_3595,N_3311,N_3340);
or U3596 (N_3596,N_3289,N_3260);
nand U3597 (N_3597,N_3348,N_3311);
or U3598 (N_3598,N_3340,N_3346);
or U3599 (N_3599,N_3388,N_3308);
or U3600 (N_3600,N_3503,N_3587);
and U3601 (N_3601,N_3426,N_3460);
nor U3602 (N_3602,N_3518,N_3496);
nand U3603 (N_3603,N_3586,N_3441);
xor U3604 (N_3604,N_3444,N_3439);
or U3605 (N_3605,N_3412,N_3470);
nor U3606 (N_3606,N_3514,N_3565);
and U3607 (N_3607,N_3471,N_3490);
and U3608 (N_3608,N_3599,N_3474);
and U3609 (N_3609,N_3433,N_3593);
and U3610 (N_3610,N_3403,N_3532);
nor U3611 (N_3611,N_3447,N_3458);
xor U3612 (N_3612,N_3548,N_3469);
nand U3613 (N_3613,N_3453,N_3451);
or U3614 (N_3614,N_3547,N_3544);
xor U3615 (N_3615,N_3494,N_3425);
xor U3616 (N_3616,N_3522,N_3524);
nand U3617 (N_3617,N_3450,N_3545);
nor U3618 (N_3618,N_3546,N_3584);
nand U3619 (N_3619,N_3574,N_3459);
or U3620 (N_3620,N_3594,N_3568);
xor U3621 (N_3621,N_3417,N_3517);
and U3622 (N_3622,N_3486,N_3509);
nor U3623 (N_3623,N_3499,N_3432);
nand U3624 (N_3624,N_3498,N_3483);
and U3625 (N_3625,N_3402,N_3549);
nor U3626 (N_3626,N_3598,N_3415);
and U3627 (N_3627,N_3575,N_3409);
or U3628 (N_3628,N_3579,N_3562);
nand U3629 (N_3629,N_3516,N_3523);
nor U3630 (N_3630,N_3407,N_3559);
xnor U3631 (N_3631,N_3489,N_3467);
nor U3632 (N_3632,N_3481,N_3478);
or U3633 (N_3633,N_3406,N_3477);
nand U3634 (N_3634,N_3421,N_3405);
xnor U3635 (N_3635,N_3527,N_3495);
nor U3636 (N_3636,N_3414,N_3502);
nor U3637 (N_3637,N_3475,N_3510);
xor U3638 (N_3638,N_3573,N_3479);
and U3639 (N_3639,N_3535,N_3526);
nand U3640 (N_3640,N_3497,N_3513);
xnor U3641 (N_3641,N_3591,N_3442);
nand U3642 (N_3642,N_3555,N_3468);
xnor U3643 (N_3643,N_3446,N_3539);
and U3644 (N_3644,N_3588,N_3519);
or U3645 (N_3645,N_3551,N_3578);
and U3646 (N_3646,N_3529,N_3572);
or U3647 (N_3647,N_3457,N_3520);
xnor U3648 (N_3648,N_3418,N_3500);
or U3649 (N_3649,N_3400,N_3465);
or U3650 (N_3650,N_3476,N_3567);
nand U3651 (N_3651,N_3589,N_3564);
nor U3652 (N_3652,N_3485,N_3511);
nor U3653 (N_3653,N_3556,N_3454);
xor U3654 (N_3654,N_3515,N_3512);
or U3655 (N_3655,N_3435,N_3416);
nand U3656 (N_3656,N_3576,N_3437);
or U3657 (N_3657,N_3569,N_3595);
and U3658 (N_3658,N_3530,N_3423);
nor U3659 (N_3659,N_3506,N_3445);
nor U3660 (N_3660,N_3427,N_3521);
or U3661 (N_3661,N_3420,N_3508);
nand U3662 (N_3662,N_3443,N_3566);
or U3663 (N_3663,N_3438,N_3550);
nand U3664 (N_3664,N_3596,N_3431);
nand U3665 (N_3665,N_3585,N_3401);
nor U3666 (N_3666,N_3552,N_3558);
xor U3667 (N_3667,N_3580,N_3505);
and U3668 (N_3668,N_3541,N_3424);
or U3669 (N_3669,N_3404,N_3429);
xor U3670 (N_3670,N_3484,N_3504);
or U3671 (N_3671,N_3462,N_3577);
nor U3672 (N_3672,N_3473,N_3472);
or U3673 (N_3673,N_3507,N_3456);
nand U3674 (N_3674,N_3597,N_3482);
xor U3675 (N_3675,N_3413,N_3449);
or U3676 (N_3676,N_3411,N_3428);
xnor U3677 (N_3677,N_3592,N_3410);
nor U3678 (N_3678,N_3533,N_3525);
or U3679 (N_3679,N_3583,N_3536);
nor U3680 (N_3680,N_3492,N_3488);
and U3681 (N_3681,N_3464,N_3538);
nor U3682 (N_3682,N_3582,N_3434);
xor U3683 (N_3683,N_3466,N_3590);
or U3684 (N_3684,N_3480,N_3561);
nor U3685 (N_3685,N_3531,N_3542);
xor U3686 (N_3686,N_3543,N_3422);
nand U3687 (N_3687,N_3408,N_3528);
nor U3688 (N_3688,N_3419,N_3448);
and U3689 (N_3689,N_3440,N_3571);
or U3690 (N_3690,N_3557,N_3570);
nor U3691 (N_3691,N_3581,N_3452);
nor U3692 (N_3692,N_3540,N_3501);
or U3693 (N_3693,N_3463,N_3461);
nor U3694 (N_3694,N_3554,N_3493);
nand U3695 (N_3695,N_3491,N_3436);
and U3696 (N_3696,N_3455,N_3534);
xnor U3697 (N_3697,N_3487,N_3560);
nand U3698 (N_3698,N_3553,N_3563);
xor U3699 (N_3699,N_3537,N_3430);
nand U3700 (N_3700,N_3560,N_3530);
xnor U3701 (N_3701,N_3479,N_3533);
nand U3702 (N_3702,N_3494,N_3432);
or U3703 (N_3703,N_3495,N_3437);
or U3704 (N_3704,N_3458,N_3497);
and U3705 (N_3705,N_3463,N_3465);
nand U3706 (N_3706,N_3462,N_3572);
xnor U3707 (N_3707,N_3498,N_3430);
nand U3708 (N_3708,N_3505,N_3453);
and U3709 (N_3709,N_3554,N_3483);
nor U3710 (N_3710,N_3434,N_3567);
nand U3711 (N_3711,N_3421,N_3563);
or U3712 (N_3712,N_3546,N_3449);
xnor U3713 (N_3713,N_3496,N_3492);
or U3714 (N_3714,N_3538,N_3590);
nor U3715 (N_3715,N_3562,N_3549);
and U3716 (N_3716,N_3577,N_3536);
or U3717 (N_3717,N_3558,N_3461);
xnor U3718 (N_3718,N_3437,N_3453);
xnor U3719 (N_3719,N_3441,N_3453);
nand U3720 (N_3720,N_3586,N_3512);
nor U3721 (N_3721,N_3455,N_3475);
xnor U3722 (N_3722,N_3420,N_3503);
xor U3723 (N_3723,N_3463,N_3538);
and U3724 (N_3724,N_3444,N_3483);
nor U3725 (N_3725,N_3422,N_3554);
and U3726 (N_3726,N_3446,N_3524);
nand U3727 (N_3727,N_3504,N_3404);
or U3728 (N_3728,N_3546,N_3510);
or U3729 (N_3729,N_3550,N_3458);
or U3730 (N_3730,N_3581,N_3556);
nor U3731 (N_3731,N_3466,N_3588);
nor U3732 (N_3732,N_3407,N_3547);
nand U3733 (N_3733,N_3464,N_3423);
nor U3734 (N_3734,N_3495,N_3558);
nand U3735 (N_3735,N_3500,N_3530);
and U3736 (N_3736,N_3544,N_3499);
and U3737 (N_3737,N_3536,N_3504);
xor U3738 (N_3738,N_3506,N_3566);
and U3739 (N_3739,N_3403,N_3461);
nor U3740 (N_3740,N_3502,N_3419);
and U3741 (N_3741,N_3561,N_3416);
nand U3742 (N_3742,N_3561,N_3511);
or U3743 (N_3743,N_3536,N_3469);
and U3744 (N_3744,N_3523,N_3529);
nor U3745 (N_3745,N_3400,N_3598);
and U3746 (N_3746,N_3465,N_3557);
xnor U3747 (N_3747,N_3543,N_3563);
xnor U3748 (N_3748,N_3488,N_3584);
or U3749 (N_3749,N_3428,N_3474);
and U3750 (N_3750,N_3469,N_3487);
and U3751 (N_3751,N_3505,N_3491);
and U3752 (N_3752,N_3448,N_3427);
and U3753 (N_3753,N_3518,N_3406);
nor U3754 (N_3754,N_3587,N_3481);
xnor U3755 (N_3755,N_3540,N_3595);
nor U3756 (N_3756,N_3545,N_3452);
xor U3757 (N_3757,N_3405,N_3443);
nor U3758 (N_3758,N_3430,N_3415);
xnor U3759 (N_3759,N_3475,N_3548);
nor U3760 (N_3760,N_3550,N_3432);
nand U3761 (N_3761,N_3566,N_3500);
nand U3762 (N_3762,N_3490,N_3460);
and U3763 (N_3763,N_3468,N_3500);
or U3764 (N_3764,N_3483,N_3411);
and U3765 (N_3765,N_3593,N_3422);
nor U3766 (N_3766,N_3407,N_3556);
nor U3767 (N_3767,N_3477,N_3469);
or U3768 (N_3768,N_3428,N_3483);
or U3769 (N_3769,N_3540,N_3539);
xor U3770 (N_3770,N_3576,N_3518);
xnor U3771 (N_3771,N_3532,N_3497);
xor U3772 (N_3772,N_3435,N_3509);
xor U3773 (N_3773,N_3442,N_3541);
nor U3774 (N_3774,N_3516,N_3502);
or U3775 (N_3775,N_3449,N_3462);
and U3776 (N_3776,N_3506,N_3516);
nand U3777 (N_3777,N_3591,N_3437);
xor U3778 (N_3778,N_3596,N_3433);
or U3779 (N_3779,N_3561,N_3457);
nor U3780 (N_3780,N_3569,N_3434);
and U3781 (N_3781,N_3552,N_3463);
nand U3782 (N_3782,N_3470,N_3402);
or U3783 (N_3783,N_3557,N_3533);
and U3784 (N_3784,N_3531,N_3592);
and U3785 (N_3785,N_3489,N_3544);
or U3786 (N_3786,N_3503,N_3431);
nor U3787 (N_3787,N_3467,N_3466);
or U3788 (N_3788,N_3437,N_3463);
or U3789 (N_3789,N_3481,N_3597);
nand U3790 (N_3790,N_3434,N_3435);
or U3791 (N_3791,N_3529,N_3404);
nor U3792 (N_3792,N_3431,N_3553);
or U3793 (N_3793,N_3538,N_3532);
or U3794 (N_3794,N_3537,N_3483);
or U3795 (N_3795,N_3545,N_3459);
nor U3796 (N_3796,N_3581,N_3591);
nor U3797 (N_3797,N_3595,N_3433);
and U3798 (N_3798,N_3415,N_3481);
xnor U3799 (N_3799,N_3412,N_3507);
xnor U3800 (N_3800,N_3602,N_3792);
nand U3801 (N_3801,N_3766,N_3759);
xor U3802 (N_3802,N_3798,N_3769);
and U3803 (N_3803,N_3658,N_3690);
nand U3804 (N_3804,N_3712,N_3780);
nand U3805 (N_3805,N_3771,N_3773);
nand U3806 (N_3806,N_3654,N_3737);
and U3807 (N_3807,N_3621,N_3666);
or U3808 (N_3808,N_3692,N_3776);
or U3809 (N_3809,N_3628,N_3642);
nand U3810 (N_3810,N_3603,N_3696);
nor U3811 (N_3811,N_3615,N_3634);
and U3812 (N_3812,N_3717,N_3695);
nor U3813 (N_3813,N_3707,N_3700);
and U3814 (N_3814,N_3752,N_3736);
and U3815 (N_3815,N_3777,N_3799);
xnor U3816 (N_3816,N_3793,N_3622);
nand U3817 (N_3817,N_3650,N_3703);
and U3818 (N_3818,N_3686,N_3785);
and U3819 (N_3819,N_3627,N_3768);
or U3820 (N_3820,N_3649,N_3770);
nor U3821 (N_3821,N_3775,N_3623);
xnor U3822 (N_3822,N_3683,N_3699);
and U3823 (N_3823,N_3612,N_3675);
nor U3824 (N_3824,N_3709,N_3697);
or U3825 (N_3825,N_3786,N_3757);
and U3826 (N_3826,N_3730,N_3632);
nand U3827 (N_3827,N_3754,N_3681);
xor U3828 (N_3828,N_3747,N_3617);
xor U3829 (N_3829,N_3610,N_3755);
xor U3830 (N_3830,N_3667,N_3758);
nor U3831 (N_3831,N_3735,N_3680);
and U3832 (N_3832,N_3608,N_3641);
xnor U3833 (N_3833,N_3783,N_3745);
or U3834 (N_3834,N_3796,N_3740);
xnor U3835 (N_3835,N_3601,N_3657);
xor U3836 (N_3836,N_3646,N_3716);
xnor U3837 (N_3837,N_3763,N_3721);
nand U3838 (N_3838,N_3715,N_3613);
nor U3839 (N_3839,N_3787,N_3772);
nand U3840 (N_3840,N_3710,N_3668);
nand U3841 (N_3841,N_3674,N_3633);
xor U3842 (N_3842,N_3784,N_3767);
or U3843 (N_3843,N_3714,N_3669);
and U3844 (N_3844,N_3645,N_3708);
xor U3845 (N_3845,N_3724,N_3729);
xor U3846 (N_3846,N_3694,N_3778);
nand U3847 (N_3847,N_3713,N_3739);
or U3848 (N_3848,N_3660,N_3620);
nand U3849 (N_3849,N_3614,N_3698);
xnor U3850 (N_3850,N_3679,N_3746);
or U3851 (N_3851,N_3779,N_3644);
or U3852 (N_3852,N_3677,N_3676);
and U3853 (N_3853,N_3616,N_3704);
nor U3854 (N_3854,N_3691,N_3722);
xor U3855 (N_3855,N_3790,N_3689);
and U3856 (N_3856,N_3693,N_3652);
or U3857 (N_3857,N_3753,N_3727);
xnor U3858 (N_3858,N_3618,N_3673);
xor U3859 (N_3859,N_3607,N_3636);
nand U3860 (N_3860,N_3665,N_3635);
and U3861 (N_3861,N_3605,N_3797);
xnor U3862 (N_3862,N_3600,N_3670);
and U3863 (N_3863,N_3606,N_3664);
and U3864 (N_3864,N_3738,N_3626);
or U3865 (N_3865,N_3688,N_3725);
nor U3866 (N_3866,N_3647,N_3630);
xor U3867 (N_3867,N_3731,N_3656);
and U3868 (N_3868,N_3748,N_3631);
nor U3869 (N_3869,N_3719,N_3732);
xnor U3870 (N_3870,N_3662,N_3604);
nand U3871 (N_3871,N_3765,N_3705);
nor U3872 (N_3872,N_3625,N_3685);
and U3873 (N_3873,N_3720,N_3743);
and U3874 (N_3874,N_3611,N_3624);
nor U3875 (N_3875,N_3781,N_3671);
nor U3876 (N_3876,N_3640,N_3762);
and U3877 (N_3877,N_3651,N_3655);
or U3878 (N_3878,N_3749,N_3760);
nand U3879 (N_3879,N_3751,N_3782);
and U3880 (N_3880,N_3609,N_3756);
nor U3881 (N_3881,N_3661,N_3711);
or U3882 (N_3882,N_3726,N_3682);
or U3883 (N_3883,N_3678,N_3687);
or U3884 (N_3884,N_3702,N_3734);
xor U3885 (N_3885,N_3774,N_3663);
nor U3886 (N_3886,N_3742,N_3744);
and U3887 (N_3887,N_3648,N_3706);
xnor U3888 (N_3888,N_3637,N_3653);
xor U3889 (N_3889,N_3761,N_3728);
or U3890 (N_3890,N_3643,N_3795);
nand U3891 (N_3891,N_3794,N_3723);
xor U3892 (N_3892,N_3718,N_3791);
and U3893 (N_3893,N_3789,N_3701);
xnor U3894 (N_3894,N_3638,N_3788);
xnor U3895 (N_3895,N_3733,N_3741);
nor U3896 (N_3896,N_3639,N_3659);
or U3897 (N_3897,N_3684,N_3750);
xnor U3898 (N_3898,N_3672,N_3764);
or U3899 (N_3899,N_3619,N_3629);
nand U3900 (N_3900,N_3714,N_3725);
or U3901 (N_3901,N_3743,N_3737);
and U3902 (N_3902,N_3718,N_3722);
nand U3903 (N_3903,N_3795,N_3747);
or U3904 (N_3904,N_3693,N_3607);
xor U3905 (N_3905,N_3689,N_3662);
nor U3906 (N_3906,N_3709,N_3675);
nand U3907 (N_3907,N_3622,N_3643);
xnor U3908 (N_3908,N_3714,N_3623);
and U3909 (N_3909,N_3613,N_3760);
or U3910 (N_3910,N_3626,N_3631);
nand U3911 (N_3911,N_3746,N_3773);
and U3912 (N_3912,N_3729,N_3657);
and U3913 (N_3913,N_3775,N_3687);
and U3914 (N_3914,N_3750,N_3672);
nand U3915 (N_3915,N_3795,N_3783);
or U3916 (N_3916,N_3783,N_3721);
or U3917 (N_3917,N_3766,N_3630);
nand U3918 (N_3918,N_3615,N_3782);
xnor U3919 (N_3919,N_3726,N_3773);
and U3920 (N_3920,N_3774,N_3621);
and U3921 (N_3921,N_3695,N_3778);
or U3922 (N_3922,N_3701,N_3638);
nand U3923 (N_3923,N_3663,N_3773);
nand U3924 (N_3924,N_3789,N_3782);
or U3925 (N_3925,N_3634,N_3793);
or U3926 (N_3926,N_3748,N_3797);
nand U3927 (N_3927,N_3656,N_3787);
nor U3928 (N_3928,N_3776,N_3798);
and U3929 (N_3929,N_3687,N_3648);
and U3930 (N_3930,N_3793,N_3688);
nand U3931 (N_3931,N_3662,N_3783);
and U3932 (N_3932,N_3754,N_3759);
nand U3933 (N_3933,N_3771,N_3620);
xor U3934 (N_3934,N_3799,N_3688);
nand U3935 (N_3935,N_3799,N_3759);
xor U3936 (N_3936,N_3712,N_3683);
nor U3937 (N_3937,N_3751,N_3786);
nor U3938 (N_3938,N_3740,N_3741);
xnor U3939 (N_3939,N_3680,N_3711);
or U3940 (N_3940,N_3658,N_3604);
or U3941 (N_3941,N_3769,N_3704);
nor U3942 (N_3942,N_3650,N_3662);
and U3943 (N_3943,N_3732,N_3606);
and U3944 (N_3944,N_3667,N_3753);
and U3945 (N_3945,N_3741,N_3652);
and U3946 (N_3946,N_3675,N_3766);
and U3947 (N_3947,N_3763,N_3701);
or U3948 (N_3948,N_3616,N_3740);
and U3949 (N_3949,N_3628,N_3784);
nand U3950 (N_3950,N_3646,N_3677);
nor U3951 (N_3951,N_3793,N_3618);
or U3952 (N_3952,N_3778,N_3655);
and U3953 (N_3953,N_3625,N_3628);
xnor U3954 (N_3954,N_3670,N_3636);
or U3955 (N_3955,N_3751,N_3686);
or U3956 (N_3956,N_3716,N_3724);
and U3957 (N_3957,N_3604,N_3624);
xnor U3958 (N_3958,N_3723,N_3783);
and U3959 (N_3959,N_3701,N_3629);
and U3960 (N_3960,N_3711,N_3781);
or U3961 (N_3961,N_3663,N_3656);
nand U3962 (N_3962,N_3635,N_3612);
xor U3963 (N_3963,N_3773,N_3697);
nor U3964 (N_3964,N_3782,N_3793);
or U3965 (N_3965,N_3730,N_3696);
nor U3966 (N_3966,N_3686,N_3723);
xor U3967 (N_3967,N_3601,N_3652);
or U3968 (N_3968,N_3781,N_3771);
or U3969 (N_3969,N_3648,N_3767);
or U3970 (N_3970,N_3775,N_3795);
or U3971 (N_3971,N_3660,N_3609);
xor U3972 (N_3972,N_3690,N_3720);
and U3973 (N_3973,N_3747,N_3647);
nand U3974 (N_3974,N_3624,N_3662);
xnor U3975 (N_3975,N_3746,N_3628);
nor U3976 (N_3976,N_3632,N_3636);
and U3977 (N_3977,N_3634,N_3770);
nand U3978 (N_3978,N_3705,N_3615);
nand U3979 (N_3979,N_3737,N_3767);
and U3980 (N_3980,N_3770,N_3793);
xnor U3981 (N_3981,N_3723,N_3617);
or U3982 (N_3982,N_3772,N_3705);
or U3983 (N_3983,N_3749,N_3628);
xor U3984 (N_3984,N_3716,N_3661);
and U3985 (N_3985,N_3715,N_3625);
or U3986 (N_3986,N_3643,N_3607);
xor U3987 (N_3987,N_3696,N_3609);
and U3988 (N_3988,N_3722,N_3795);
nor U3989 (N_3989,N_3797,N_3721);
xor U3990 (N_3990,N_3648,N_3779);
nor U3991 (N_3991,N_3756,N_3710);
or U3992 (N_3992,N_3637,N_3672);
nor U3993 (N_3993,N_3645,N_3692);
and U3994 (N_3994,N_3673,N_3645);
nor U3995 (N_3995,N_3710,N_3789);
xor U3996 (N_3996,N_3615,N_3687);
nor U3997 (N_3997,N_3682,N_3733);
or U3998 (N_3998,N_3617,N_3798);
nand U3999 (N_3999,N_3688,N_3700);
xnor U4000 (N_4000,N_3888,N_3989);
and U4001 (N_4001,N_3903,N_3800);
nor U4002 (N_4002,N_3890,N_3933);
or U4003 (N_4003,N_3885,N_3832);
or U4004 (N_4004,N_3994,N_3869);
nor U4005 (N_4005,N_3921,N_3884);
or U4006 (N_4006,N_3872,N_3844);
and U4007 (N_4007,N_3806,N_3906);
and U4008 (N_4008,N_3986,N_3914);
and U4009 (N_4009,N_3980,N_3870);
and U4010 (N_4010,N_3947,N_3949);
nor U4011 (N_4011,N_3871,N_3831);
nand U4012 (N_4012,N_3856,N_3905);
and U4013 (N_4013,N_3957,N_3984);
and U4014 (N_4014,N_3912,N_3883);
xor U4015 (N_4015,N_3891,N_3878);
and U4016 (N_4016,N_3995,N_3930);
nand U4017 (N_4017,N_3932,N_3810);
or U4018 (N_4018,N_3849,N_3899);
or U4019 (N_4019,N_3911,N_3961);
nor U4020 (N_4020,N_3898,N_3972);
nor U4021 (N_4021,N_3838,N_3946);
and U4022 (N_4022,N_3965,N_3877);
and U4023 (N_4023,N_3900,N_3979);
xor U4024 (N_4024,N_3804,N_3845);
or U4025 (N_4025,N_3978,N_3808);
nand U4026 (N_4026,N_3850,N_3915);
or U4027 (N_4027,N_3812,N_3881);
xnor U4028 (N_4028,N_3920,N_3853);
nor U4029 (N_4029,N_3822,N_3807);
and U4030 (N_4030,N_3834,N_3981);
nor U4031 (N_4031,N_3862,N_3817);
and U4032 (N_4032,N_3931,N_3910);
or U4033 (N_4033,N_3815,N_3969);
nand U4034 (N_4034,N_3923,N_3959);
nor U4035 (N_4035,N_3860,N_3828);
and U4036 (N_4036,N_3892,N_3889);
nor U4037 (N_4037,N_3814,N_3945);
and U4038 (N_4038,N_3970,N_3854);
xnor U4039 (N_4039,N_3934,N_3897);
nand U4040 (N_4040,N_3967,N_3985);
or U4041 (N_4041,N_3936,N_3955);
xnor U4042 (N_4042,N_3996,N_3880);
and U4043 (N_4043,N_3827,N_3913);
nand U4044 (N_4044,N_3937,N_3848);
nand U4045 (N_4045,N_3858,N_3960);
or U4046 (N_4046,N_3837,N_3924);
xor U4047 (N_4047,N_3802,N_3823);
or U4048 (N_4048,N_3864,N_3939);
or U4049 (N_4049,N_3847,N_3865);
and U4050 (N_4050,N_3968,N_3958);
or U4051 (N_4051,N_3895,N_3942);
nand U4052 (N_4052,N_3974,N_3971);
and U4053 (N_4053,N_3840,N_3855);
or U4054 (N_4054,N_3927,N_3940);
nor U4055 (N_4055,N_3821,N_3917);
nor U4056 (N_4056,N_3824,N_3833);
nand U4057 (N_4057,N_3830,N_3902);
nor U4058 (N_4058,N_3825,N_3963);
or U4059 (N_4059,N_3992,N_3803);
nand U4060 (N_4060,N_3819,N_3962);
and U4061 (N_4061,N_3809,N_3861);
xnor U4062 (N_4062,N_3964,N_3852);
and U4063 (N_4063,N_3846,N_3901);
nand U4064 (N_4064,N_3938,N_3820);
xor U4065 (N_4065,N_3935,N_3987);
or U4066 (N_4066,N_3925,N_3999);
xnor U4067 (N_4067,N_3868,N_3907);
nand U4068 (N_4068,N_3966,N_3863);
xor U4069 (N_4069,N_3977,N_3908);
xnor U4070 (N_4070,N_3926,N_3918);
nor U4071 (N_4071,N_3909,N_3950);
or U4072 (N_4072,N_3952,N_3813);
nor U4073 (N_4073,N_3983,N_3842);
nor U4074 (N_4074,N_3988,N_3886);
or U4075 (N_4075,N_3816,N_3973);
nand U4076 (N_4076,N_3867,N_3976);
nand U4077 (N_4077,N_3982,N_3818);
nor U4078 (N_4078,N_3873,N_3836);
and U4079 (N_4079,N_3929,N_3882);
xnor U4080 (N_4080,N_3916,N_3887);
xnor U4081 (N_4081,N_3839,N_3997);
and U4082 (N_4082,N_3801,N_3875);
xnor U4083 (N_4083,N_3829,N_3990);
or U4084 (N_4084,N_3904,N_3851);
nand U4085 (N_4085,N_3879,N_3928);
nor U4086 (N_4086,N_3975,N_3859);
or U4087 (N_4087,N_3874,N_3805);
or U4088 (N_4088,N_3998,N_3894);
xnor U4089 (N_4089,N_3954,N_3944);
and U4090 (N_4090,N_3893,N_3876);
xnor U4091 (N_4091,N_3993,N_3943);
nor U4092 (N_4092,N_3956,N_3991);
or U4093 (N_4093,N_3953,N_3948);
nor U4094 (N_4094,N_3919,N_3896);
xor U4095 (N_4095,N_3843,N_3941);
xor U4096 (N_4096,N_3835,N_3826);
nor U4097 (N_4097,N_3811,N_3841);
or U4098 (N_4098,N_3922,N_3857);
or U4099 (N_4099,N_3951,N_3866);
or U4100 (N_4100,N_3843,N_3980);
nor U4101 (N_4101,N_3858,N_3840);
nand U4102 (N_4102,N_3950,N_3835);
xor U4103 (N_4103,N_3930,N_3948);
nor U4104 (N_4104,N_3857,N_3808);
nand U4105 (N_4105,N_3954,N_3808);
xor U4106 (N_4106,N_3831,N_3994);
nor U4107 (N_4107,N_3832,N_3923);
xor U4108 (N_4108,N_3918,N_3899);
nand U4109 (N_4109,N_3983,N_3847);
or U4110 (N_4110,N_3891,N_3852);
or U4111 (N_4111,N_3813,N_3988);
or U4112 (N_4112,N_3841,N_3971);
or U4113 (N_4113,N_3808,N_3820);
xnor U4114 (N_4114,N_3923,N_3883);
and U4115 (N_4115,N_3892,N_3974);
nand U4116 (N_4116,N_3902,N_3929);
or U4117 (N_4117,N_3993,N_3813);
nand U4118 (N_4118,N_3978,N_3964);
or U4119 (N_4119,N_3939,N_3995);
or U4120 (N_4120,N_3899,N_3871);
or U4121 (N_4121,N_3945,N_3845);
nor U4122 (N_4122,N_3894,N_3845);
nand U4123 (N_4123,N_3832,N_3819);
or U4124 (N_4124,N_3997,N_3924);
nor U4125 (N_4125,N_3907,N_3901);
nand U4126 (N_4126,N_3921,N_3847);
nor U4127 (N_4127,N_3875,N_3951);
nand U4128 (N_4128,N_3970,N_3918);
nor U4129 (N_4129,N_3877,N_3848);
xor U4130 (N_4130,N_3887,N_3949);
nand U4131 (N_4131,N_3835,N_3948);
xnor U4132 (N_4132,N_3825,N_3930);
nand U4133 (N_4133,N_3954,N_3853);
and U4134 (N_4134,N_3879,N_3906);
or U4135 (N_4135,N_3919,N_3898);
or U4136 (N_4136,N_3985,N_3982);
or U4137 (N_4137,N_3944,N_3860);
nand U4138 (N_4138,N_3882,N_3932);
xnor U4139 (N_4139,N_3834,N_3866);
nand U4140 (N_4140,N_3857,N_3975);
or U4141 (N_4141,N_3888,N_3950);
nor U4142 (N_4142,N_3803,N_3856);
and U4143 (N_4143,N_3825,N_3817);
nor U4144 (N_4144,N_3978,N_3972);
nor U4145 (N_4145,N_3842,N_3812);
nand U4146 (N_4146,N_3890,N_3884);
or U4147 (N_4147,N_3911,N_3924);
or U4148 (N_4148,N_3835,N_3968);
xor U4149 (N_4149,N_3841,N_3962);
xnor U4150 (N_4150,N_3853,N_3898);
xnor U4151 (N_4151,N_3834,N_3921);
nand U4152 (N_4152,N_3823,N_3887);
and U4153 (N_4153,N_3822,N_3867);
nand U4154 (N_4154,N_3883,N_3827);
xnor U4155 (N_4155,N_3936,N_3845);
nor U4156 (N_4156,N_3857,N_3960);
nor U4157 (N_4157,N_3820,N_3866);
and U4158 (N_4158,N_3883,N_3930);
xor U4159 (N_4159,N_3959,N_3810);
nand U4160 (N_4160,N_3825,N_3866);
xnor U4161 (N_4161,N_3880,N_3956);
or U4162 (N_4162,N_3907,N_3997);
xor U4163 (N_4163,N_3958,N_3881);
nand U4164 (N_4164,N_3960,N_3992);
and U4165 (N_4165,N_3801,N_3904);
xor U4166 (N_4166,N_3830,N_3999);
xnor U4167 (N_4167,N_3901,N_3997);
nand U4168 (N_4168,N_3804,N_3814);
nor U4169 (N_4169,N_3928,N_3823);
nand U4170 (N_4170,N_3962,N_3918);
or U4171 (N_4171,N_3968,N_3931);
nor U4172 (N_4172,N_3989,N_3886);
or U4173 (N_4173,N_3817,N_3849);
xnor U4174 (N_4174,N_3824,N_3937);
and U4175 (N_4175,N_3961,N_3865);
nor U4176 (N_4176,N_3883,N_3971);
or U4177 (N_4177,N_3953,N_3804);
and U4178 (N_4178,N_3849,N_3843);
nand U4179 (N_4179,N_3917,N_3942);
and U4180 (N_4180,N_3834,N_3963);
nand U4181 (N_4181,N_3904,N_3963);
nand U4182 (N_4182,N_3867,N_3985);
and U4183 (N_4183,N_3880,N_3947);
xor U4184 (N_4184,N_3992,N_3809);
and U4185 (N_4185,N_3941,N_3824);
nor U4186 (N_4186,N_3967,N_3810);
and U4187 (N_4187,N_3986,N_3916);
nand U4188 (N_4188,N_3842,N_3908);
nand U4189 (N_4189,N_3852,N_3914);
or U4190 (N_4190,N_3996,N_3986);
and U4191 (N_4191,N_3831,N_3878);
nand U4192 (N_4192,N_3902,N_3842);
xor U4193 (N_4193,N_3916,N_3962);
xor U4194 (N_4194,N_3880,N_3836);
nand U4195 (N_4195,N_3938,N_3844);
and U4196 (N_4196,N_3862,N_3812);
nand U4197 (N_4197,N_3834,N_3858);
or U4198 (N_4198,N_3805,N_3883);
nand U4199 (N_4199,N_3802,N_3816);
and U4200 (N_4200,N_4193,N_4063);
and U4201 (N_4201,N_4106,N_4069);
nand U4202 (N_4202,N_4189,N_4140);
nor U4203 (N_4203,N_4139,N_4013);
and U4204 (N_4204,N_4177,N_4035);
or U4205 (N_4205,N_4095,N_4173);
xnor U4206 (N_4206,N_4159,N_4129);
or U4207 (N_4207,N_4084,N_4008);
nor U4208 (N_4208,N_4163,N_4015);
or U4209 (N_4209,N_4056,N_4142);
or U4210 (N_4210,N_4104,N_4179);
nand U4211 (N_4211,N_4157,N_4103);
or U4212 (N_4212,N_4018,N_4098);
xnor U4213 (N_4213,N_4100,N_4114);
and U4214 (N_4214,N_4057,N_4121);
xnor U4215 (N_4215,N_4158,N_4178);
nand U4216 (N_4216,N_4006,N_4077);
and U4217 (N_4217,N_4074,N_4164);
nand U4218 (N_4218,N_4079,N_4170);
or U4219 (N_4219,N_4032,N_4083);
xnor U4220 (N_4220,N_4148,N_4071);
nor U4221 (N_4221,N_4132,N_4045);
xnor U4222 (N_4222,N_4089,N_4105);
nor U4223 (N_4223,N_4010,N_4182);
or U4224 (N_4224,N_4168,N_4138);
xnor U4225 (N_4225,N_4065,N_4119);
nand U4226 (N_4226,N_4186,N_4017);
nand U4227 (N_4227,N_4194,N_4060);
nor U4228 (N_4228,N_4149,N_4120);
or U4229 (N_4229,N_4090,N_4183);
nor U4230 (N_4230,N_4144,N_4123);
and U4231 (N_4231,N_4038,N_4094);
xnor U4232 (N_4232,N_4175,N_4027);
or U4233 (N_4233,N_4117,N_4002);
nor U4234 (N_4234,N_4001,N_4188);
xor U4235 (N_4235,N_4147,N_4047);
and U4236 (N_4236,N_4191,N_4185);
or U4237 (N_4237,N_4033,N_4097);
xor U4238 (N_4238,N_4118,N_4022);
nand U4239 (N_4239,N_4176,N_4125);
xor U4240 (N_4240,N_4196,N_4034);
and U4241 (N_4241,N_4126,N_4054);
nand U4242 (N_4242,N_4052,N_4135);
and U4243 (N_4243,N_4145,N_4153);
or U4244 (N_4244,N_4025,N_4092);
nand U4245 (N_4245,N_4101,N_4146);
and U4246 (N_4246,N_4143,N_4066);
xor U4247 (N_4247,N_4174,N_4005);
nand U4248 (N_4248,N_4059,N_4091);
or U4249 (N_4249,N_4102,N_4112);
and U4250 (N_4250,N_4046,N_4042);
nor U4251 (N_4251,N_4070,N_4136);
or U4252 (N_4252,N_4156,N_4093);
or U4253 (N_4253,N_4151,N_4037);
or U4254 (N_4254,N_4080,N_4050);
and U4255 (N_4255,N_4044,N_4048);
xor U4256 (N_4256,N_4150,N_4058);
nor U4257 (N_4257,N_4012,N_4049);
or U4258 (N_4258,N_4130,N_4064);
or U4259 (N_4259,N_4021,N_4085);
nand U4260 (N_4260,N_4075,N_4113);
or U4261 (N_4261,N_4082,N_4029);
or U4262 (N_4262,N_4108,N_4127);
xor U4263 (N_4263,N_4004,N_4116);
or U4264 (N_4264,N_4169,N_4026);
or U4265 (N_4265,N_4086,N_4133);
xor U4266 (N_4266,N_4198,N_4111);
or U4267 (N_4267,N_4115,N_4078);
xnor U4268 (N_4268,N_4141,N_4199);
and U4269 (N_4269,N_4014,N_4166);
xor U4270 (N_4270,N_4197,N_4195);
and U4271 (N_4271,N_4162,N_4154);
xor U4272 (N_4272,N_4020,N_4011);
xor U4273 (N_4273,N_4072,N_4000);
and U4274 (N_4274,N_4187,N_4088);
and U4275 (N_4275,N_4131,N_4067);
or U4276 (N_4276,N_4181,N_4028);
nand U4277 (N_4277,N_4081,N_4184);
or U4278 (N_4278,N_4062,N_4055);
nor U4279 (N_4279,N_4161,N_4030);
and U4280 (N_4280,N_4053,N_4172);
nor U4281 (N_4281,N_4031,N_4190);
xnor U4282 (N_4282,N_4043,N_4076);
or U4283 (N_4283,N_4024,N_4099);
or U4284 (N_4284,N_4124,N_4128);
nor U4285 (N_4285,N_4107,N_4040);
xnor U4286 (N_4286,N_4087,N_4036);
xor U4287 (N_4287,N_4171,N_4003);
or U4288 (N_4288,N_4019,N_4051);
xor U4289 (N_4289,N_4096,N_4152);
nor U4290 (N_4290,N_4041,N_4007);
nand U4291 (N_4291,N_4068,N_4167);
nand U4292 (N_4292,N_4192,N_4180);
or U4293 (N_4293,N_4137,N_4039);
nor U4294 (N_4294,N_4160,N_4155);
and U4295 (N_4295,N_4009,N_4061);
nand U4296 (N_4296,N_4016,N_4023);
or U4297 (N_4297,N_4110,N_4165);
nand U4298 (N_4298,N_4134,N_4073);
nand U4299 (N_4299,N_4122,N_4109);
nand U4300 (N_4300,N_4138,N_4151);
xor U4301 (N_4301,N_4041,N_4094);
and U4302 (N_4302,N_4197,N_4122);
or U4303 (N_4303,N_4022,N_4192);
nor U4304 (N_4304,N_4162,N_4049);
or U4305 (N_4305,N_4044,N_4023);
or U4306 (N_4306,N_4161,N_4014);
nor U4307 (N_4307,N_4186,N_4073);
xnor U4308 (N_4308,N_4101,N_4111);
nor U4309 (N_4309,N_4018,N_4055);
or U4310 (N_4310,N_4061,N_4103);
nor U4311 (N_4311,N_4082,N_4138);
or U4312 (N_4312,N_4125,N_4111);
nor U4313 (N_4313,N_4005,N_4187);
and U4314 (N_4314,N_4097,N_4013);
nand U4315 (N_4315,N_4121,N_4078);
or U4316 (N_4316,N_4091,N_4165);
nand U4317 (N_4317,N_4044,N_4189);
and U4318 (N_4318,N_4165,N_4118);
nand U4319 (N_4319,N_4028,N_4039);
xor U4320 (N_4320,N_4190,N_4147);
nor U4321 (N_4321,N_4140,N_4118);
and U4322 (N_4322,N_4077,N_4047);
and U4323 (N_4323,N_4045,N_4142);
and U4324 (N_4324,N_4070,N_4150);
nand U4325 (N_4325,N_4143,N_4120);
nand U4326 (N_4326,N_4068,N_4000);
and U4327 (N_4327,N_4144,N_4192);
and U4328 (N_4328,N_4165,N_4037);
nor U4329 (N_4329,N_4195,N_4145);
or U4330 (N_4330,N_4091,N_4124);
or U4331 (N_4331,N_4182,N_4101);
or U4332 (N_4332,N_4158,N_4193);
or U4333 (N_4333,N_4004,N_4049);
nand U4334 (N_4334,N_4154,N_4059);
and U4335 (N_4335,N_4078,N_4052);
or U4336 (N_4336,N_4146,N_4035);
and U4337 (N_4337,N_4159,N_4047);
and U4338 (N_4338,N_4087,N_4164);
nand U4339 (N_4339,N_4076,N_4161);
nor U4340 (N_4340,N_4011,N_4142);
and U4341 (N_4341,N_4058,N_4021);
and U4342 (N_4342,N_4157,N_4092);
nand U4343 (N_4343,N_4146,N_4044);
or U4344 (N_4344,N_4123,N_4193);
nor U4345 (N_4345,N_4133,N_4106);
and U4346 (N_4346,N_4048,N_4110);
or U4347 (N_4347,N_4106,N_4048);
or U4348 (N_4348,N_4168,N_4157);
nand U4349 (N_4349,N_4139,N_4060);
nand U4350 (N_4350,N_4018,N_4101);
nand U4351 (N_4351,N_4013,N_4050);
or U4352 (N_4352,N_4056,N_4107);
xnor U4353 (N_4353,N_4002,N_4031);
or U4354 (N_4354,N_4012,N_4001);
and U4355 (N_4355,N_4104,N_4110);
and U4356 (N_4356,N_4144,N_4109);
nor U4357 (N_4357,N_4078,N_4028);
or U4358 (N_4358,N_4119,N_4132);
nor U4359 (N_4359,N_4161,N_4016);
or U4360 (N_4360,N_4170,N_4123);
nand U4361 (N_4361,N_4089,N_4043);
nor U4362 (N_4362,N_4032,N_4145);
or U4363 (N_4363,N_4144,N_4150);
or U4364 (N_4364,N_4074,N_4193);
or U4365 (N_4365,N_4008,N_4009);
nand U4366 (N_4366,N_4148,N_4041);
nor U4367 (N_4367,N_4117,N_4017);
nand U4368 (N_4368,N_4057,N_4032);
and U4369 (N_4369,N_4199,N_4091);
nand U4370 (N_4370,N_4035,N_4101);
nor U4371 (N_4371,N_4069,N_4146);
xnor U4372 (N_4372,N_4024,N_4104);
or U4373 (N_4373,N_4127,N_4166);
nand U4374 (N_4374,N_4031,N_4019);
or U4375 (N_4375,N_4032,N_4097);
or U4376 (N_4376,N_4125,N_4142);
nor U4377 (N_4377,N_4133,N_4052);
or U4378 (N_4378,N_4070,N_4021);
nand U4379 (N_4379,N_4188,N_4089);
nand U4380 (N_4380,N_4132,N_4199);
and U4381 (N_4381,N_4100,N_4155);
or U4382 (N_4382,N_4169,N_4147);
nand U4383 (N_4383,N_4046,N_4072);
nand U4384 (N_4384,N_4058,N_4105);
nor U4385 (N_4385,N_4132,N_4130);
or U4386 (N_4386,N_4132,N_4072);
xor U4387 (N_4387,N_4120,N_4075);
and U4388 (N_4388,N_4082,N_4053);
nand U4389 (N_4389,N_4178,N_4010);
and U4390 (N_4390,N_4078,N_4015);
and U4391 (N_4391,N_4096,N_4125);
and U4392 (N_4392,N_4005,N_4110);
or U4393 (N_4393,N_4160,N_4078);
or U4394 (N_4394,N_4154,N_4043);
nor U4395 (N_4395,N_4049,N_4181);
nand U4396 (N_4396,N_4032,N_4189);
or U4397 (N_4397,N_4144,N_4079);
xnor U4398 (N_4398,N_4139,N_4177);
xnor U4399 (N_4399,N_4007,N_4065);
and U4400 (N_4400,N_4307,N_4315);
nand U4401 (N_4401,N_4215,N_4338);
nor U4402 (N_4402,N_4369,N_4263);
xor U4403 (N_4403,N_4225,N_4312);
nor U4404 (N_4404,N_4216,N_4289);
nor U4405 (N_4405,N_4398,N_4249);
xnor U4406 (N_4406,N_4282,N_4300);
nor U4407 (N_4407,N_4275,N_4294);
nand U4408 (N_4408,N_4280,N_4299);
nand U4409 (N_4409,N_4291,N_4269);
xnor U4410 (N_4410,N_4359,N_4351);
xnor U4411 (N_4411,N_4335,N_4332);
and U4412 (N_4412,N_4247,N_4256);
or U4413 (N_4413,N_4266,N_4203);
nand U4414 (N_4414,N_4232,N_4229);
or U4415 (N_4415,N_4322,N_4234);
or U4416 (N_4416,N_4394,N_4213);
xor U4417 (N_4417,N_4255,N_4377);
or U4418 (N_4418,N_4257,N_4328);
xor U4419 (N_4419,N_4314,N_4251);
and U4420 (N_4420,N_4325,N_4310);
nor U4421 (N_4421,N_4302,N_4278);
xnor U4422 (N_4422,N_4270,N_4358);
nor U4423 (N_4423,N_4217,N_4205);
and U4424 (N_4424,N_4250,N_4318);
and U4425 (N_4425,N_4349,N_4274);
xnor U4426 (N_4426,N_4371,N_4220);
and U4427 (N_4427,N_4341,N_4397);
and U4428 (N_4428,N_4352,N_4285);
or U4429 (N_4429,N_4372,N_4242);
and U4430 (N_4430,N_4378,N_4379);
and U4431 (N_4431,N_4283,N_4383);
and U4432 (N_4432,N_4262,N_4260);
or U4433 (N_4433,N_4284,N_4287);
nor U4434 (N_4434,N_4393,N_4355);
nand U4435 (N_4435,N_4243,N_4237);
and U4436 (N_4436,N_4373,N_4226);
xor U4437 (N_4437,N_4384,N_4389);
and U4438 (N_4438,N_4221,N_4375);
and U4439 (N_4439,N_4253,N_4347);
or U4440 (N_4440,N_4345,N_4340);
nor U4441 (N_4441,N_4254,N_4392);
nand U4442 (N_4442,N_4381,N_4252);
nand U4443 (N_4443,N_4235,N_4222);
nor U4444 (N_4444,N_4301,N_4200);
nor U4445 (N_4445,N_4277,N_4321);
xnor U4446 (N_4446,N_4391,N_4380);
xnor U4447 (N_4447,N_4201,N_4334);
nor U4448 (N_4448,N_4376,N_4390);
xnor U4449 (N_4449,N_4268,N_4236);
nand U4450 (N_4450,N_4308,N_4303);
and U4451 (N_4451,N_4218,N_4223);
xor U4452 (N_4452,N_4292,N_4239);
nand U4453 (N_4453,N_4210,N_4360);
nand U4454 (N_4454,N_4357,N_4233);
nand U4455 (N_4455,N_4382,N_4343);
nand U4456 (N_4456,N_4202,N_4336);
nor U4457 (N_4457,N_4259,N_4388);
or U4458 (N_4458,N_4261,N_4309);
xor U4459 (N_4459,N_4241,N_4330);
or U4460 (N_4460,N_4272,N_4333);
nor U4461 (N_4461,N_4374,N_4396);
or U4462 (N_4462,N_4317,N_4366);
or U4463 (N_4463,N_4208,N_4385);
nand U4464 (N_4464,N_4219,N_4342);
xor U4465 (N_4465,N_4363,N_4207);
nor U4466 (N_4466,N_4264,N_4395);
nand U4467 (N_4467,N_4231,N_4387);
xor U4468 (N_4468,N_4246,N_4295);
nor U4469 (N_4469,N_4290,N_4311);
nand U4470 (N_4470,N_4364,N_4297);
nand U4471 (N_4471,N_4368,N_4286);
nor U4472 (N_4472,N_4327,N_4367);
nor U4473 (N_4473,N_4209,N_4313);
and U4474 (N_4474,N_4204,N_4271);
nand U4475 (N_4475,N_4354,N_4362);
nand U4476 (N_4476,N_4306,N_4326);
nand U4477 (N_4477,N_4296,N_4288);
nor U4478 (N_4478,N_4324,N_4248);
nand U4479 (N_4479,N_4344,N_4323);
and U4480 (N_4480,N_4365,N_4206);
nand U4481 (N_4481,N_4212,N_4265);
nand U4482 (N_4482,N_4245,N_4230);
nor U4483 (N_4483,N_4273,N_4227);
and U4484 (N_4484,N_4281,N_4320);
nor U4485 (N_4485,N_4346,N_4353);
nor U4486 (N_4486,N_4276,N_4331);
xnor U4487 (N_4487,N_4240,N_4350);
nor U4488 (N_4488,N_4337,N_4267);
xor U4489 (N_4489,N_4370,N_4228);
nor U4490 (N_4490,N_4386,N_4339);
xor U4491 (N_4491,N_4258,N_4329);
or U4492 (N_4492,N_4319,N_4304);
nand U4493 (N_4493,N_4361,N_4298);
xnor U4494 (N_4494,N_4211,N_4279);
nor U4495 (N_4495,N_4214,N_4348);
xor U4496 (N_4496,N_4293,N_4305);
or U4497 (N_4497,N_4316,N_4244);
and U4498 (N_4498,N_4224,N_4399);
nand U4499 (N_4499,N_4356,N_4238);
nor U4500 (N_4500,N_4293,N_4322);
xor U4501 (N_4501,N_4372,N_4290);
or U4502 (N_4502,N_4363,N_4270);
nor U4503 (N_4503,N_4221,N_4374);
xnor U4504 (N_4504,N_4376,N_4287);
or U4505 (N_4505,N_4339,N_4354);
xnor U4506 (N_4506,N_4303,N_4338);
and U4507 (N_4507,N_4200,N_4317);
or U4508 (N_4508,N_4370,N_4358);
nor U4509 (N_4509,N_4331,N_4234);
nand U4510 (N_4510,N_4212,N_4357);
xnor U4511 (N_4511,N_4371,N_4361);
nand U4512 (N_4512,N_4264,N_4269);
nor U4513 (N_4513,N_4306,N_4375);
and U4514 (N_4514,N_4245,N_4263);
nor U4515 (N_4515,N_4279,N_4308);
and U4516 (N_4516,N_4279,N_4248);
nor U4517 (N_4517,N_4383,N_4324);
or U4518 (N_4518,N_4249,N_4223);
nor U4519 (N_4519,N_4258,N_4344);
and U4520 (N_4520,N_4386,N_4266);
or U4521 (N_4521,N_4292,N_4367);
nand U4522 (N_4522,N_4351,N_4205);
nor U4523 (N_4523,N_4228,N_4221);
nand U4524 (N_4524,N_4211,N_4287);
nand U4525 (N_4525,N_4273,N_4389);
nor U4526 (N_4526,N_4377,N_4256);
and U4527 (N_4527,N_4262,N_4322);
or U4528 (N_4528,N_4311,N_4225);
xnor U4529 (N_4529,N_4208,N_4262);
nand U4530 (N_4530,N_4271,N_4299);
and U4531 (N_4531,N_4297,N_4230);
xnor U4532 (N_4532,N_4341,N_4371);
xor U4533 (N_4533,N_4271,N_4392);
nor U4534 (N_4534,N_4202,N_4363);
nor U4535 (N_4535,N_4399,N_4238);
and U4536 (N_4536,N_4261,N_4222);
or U4537 (N_4537,N_4301,N_4234);
or U4538 (N_4538,N_4383,N_4396);
or U4539 (N_4539,N_4249,N_4359);
nor U4540 (N_4540,N_4240,N_4288);
nor U4541 (N_4541,N_4291,N_4203);
or U4542 (N_4542,N_4346,N_4314);
and U4543 (N_4543,N_4276,N_4235);
and U4544 (N_4544,N_4393,N_4296);
nor U4545 (N_4545,N_4221,N_4203);
nor U4546 (N_4546,N_4277,N_4236);
and U4547 (N_4547,N_4363,N_4377);
or U4548 (N_4548,N_4305,N_4233);
nor U4549 (N_4549,N_4276,N_4382);
nand U4550 (N_4550,N_4270,N_4303);
xor U4551 (N_4551,N_4225,N_4231);
nor U4552 (N_4552,N_4266,N_4355);
nand U4553 (N_4553,N_4243,N_4287);
nand U4554 (N_4554,N_4306,N_4399);
nor U4555 (N_4555,N_4208,N_4310);
xnor U4556 (N_4556,N_4352,N_4377);
nor U4557 (N_4557,N_4290,N_4320);
or U4558 (N_4558,N_4271,N_4290);
and U4559 (N_4559,N_4295,N_4396);
xor U4560 (N_4560,N_4281,N_4317);
xor U4561 (N_4561,N_4232,N_4384);
and U4562 (N_4562,N_4372,N_4322);
nand U4563 (N_4563,N_4274,N_4363);
or U4564 (N_4564,N_4208,N_4281);
xor U4565 (N_4565,N_4319,N_4336);
nand U4566 (N_4566,N_4327,N_4232);
and U4567 (N_4567,N_4248,N_4235);
and U4568 (N_4568,N_4378,N_4258);
nand U4569 (N_4569,N_4399,N_4239);
and U4570 (N_4570,N_4246,N_4249);
xnor U4571 (N_4571,N_4305,N_4220);
xnor U4572 (N_4572,N_4236,N_4316);
nor U4573 (N_4573,N_4378,N_4271);
nor U4574 (N_4574,N_4381,N_4225);
or U4575 (N_4575,N_4214,N_4218);
xnor U4576 (N_4576,N_4241,N_4292);
xor U4577 (N_4577,N_4338,N_4234);
or U4578 (N_4578,N_4236,N_4319);
and U4579 (N_4579,N_4207,N_4257);
nand U4580 (N_4580,N_4314,N_4352);
and U4581 (N_4581,N_4319,N_4310);
xnor U4582 (N_4582,N_4239,N_4393);
nand U4583 (N_4583,N_4252,N_4317);
nor U4584 (N_4584,N_4373,N_4347);
xnor U4585 (N_4585,N_4296,N_4339);
and U4586 (N_4586,N_4301,N_4208);
or U4587 (N_4587,N_4334,N_4343);
xor U4588 (N_4588,N_4340,N_4297);
and U4589 (N_4589,N_4289,N_4266);
nand U4590 (N_4590,N_4355,N_4327);
or U4591 (N_4591,N_4274,N_4353);
and U4592 (N_4592,N_4300,N_4307);
nand U4593 (N_4593,N_4282,N_4218);
or U4594 (N_4594,N_4371,N_4358);
or U4595 (N_4595,N_4302,N_4298);
nand U4596 (N_4596,N_4350,N_4223);
xnor U4597 (N_4597,N_4385,N_4397);
and U4598 (N_4598,N_4222,N_4382);
xnor U4599 (N_4599,N_4353,N_4326);
nand U4600 (N_4600,N_4582,N_4543);
nor U4601 (N_4601,N_4480,N_4545);
xnor U4602 (N_4602,N_4525,N_4571);
xnor U4603 (N_4603,N_4404,N_4414);
xnor U4604 (N_4604,N_4458,N_4454);
nand U4605 (N_4605,N_4503,N_4415);
and U4606 (N_4606,N_4511,N_4565);
nor U4607 (N_4607,N_4470,N_4475);
xnor U4608 (N_4608,N_4455,N_4595);
nand U4609 (N_4609,N_4485,N_4497);
xnor U4610 (N_4610,N_4590,N_4574);
nor U4611 (N_4611,N_4563,N_4459);
and U4612 (N_4612,N_4561,N_4416);
nor U4613 (N_4613,N_4438,N_4538);
and U4614 (N_4614,N_4473,N_4424);
and U4615 (N_4615,N_4558,N_4486);
and U4616 (N_4616,N_4578,N_4434);
and U4617 (N_4617,N_4507,N_4586);
nand U4618 (N_4618,N_4527,N_4544);
xnor U4619 (N_4619,N_4477,N_4429);
xnor U4620 (N_4620,N_4488,N_4401);
nor U4621 (N_4621,N_4426,N_4554);
nand U4622 (N_4622,N_4496,N_4583);
and U4623 (N_4623,N_4425,N_4483);
nor U4624 (N_4624,N_4594,N_4461);
nand U4625 (N_4625,N_4508,N_4474);
nand U4626 (N_4626,N_4411,N_4552);
xnor U4627 (N_4627,N_4541,N_4575);
and U4628 (N_4628,N_4421,N_4437);
nand U4629 (N_4629,N_4514,N_4494);
and U4630 (N_4630,N_4419,N_4519);
nor U4631 (N_4631,N_4417,N_4481);
or U4632 (N_4632,N_4442,N_4448);
and U4633 (N_4633,N_4431,N_4418);
xnor U4634 (N_4634,N_4524,N_4515);
or U4635 (N_4635,N_4478,N_4462);
nor U4636 (N_4636,N_4509,N_4567);
nand U4637 (N_4637,N_4439,N_4484);
or U4638 (N_4638,N_4526,N_4435);
nand U4639 (N_4639,N_4569,N_4550);
or U4640 (N_4640,N_4498,N_4579);
nand U4641 (N_4641,N_4451,N_4531);
nand U4642 (N_4642,N_4467,N_4585);
nand U4643 (N_4643,N_4542,N_4557);
nand U4644 (N_4644,N_4482,N_4407);
xnor U4645 (N_4645,N_4433,N_4555);
nor U4646 (N_4646,N_4537,N_4492);
and U4647 (N_4647,N_4469,N_4553);
or U4648 (N_4648,N_4589,N_4540);
and U4649 (N_4649,N_4568,N_4529);
or U4650 (N_4650,N_4562,N_4500);
and U4651 (N_4651,N_4539,N_4428);
nand U4652 (N_4652,N_4546,N_4587);
or U4653 (N_4653,N_4573,N_4533);
xnor U4654 (N_4654,N_4560,N_4491);
nand U4655 (N_4655,N_4593,N_4460);
or U4656 (N_4656,N_4599,N_4532);
nor U4657 (N_4657,N_4523,N_4577);
xnor U4658 (N_4658,N_4452,N_4410);
nor U4659 (N_4659,N_4406,N_4534);
and U4660 (N_4660,N_4464,N_4598);
or U4661 (N_4661,N_4430,N_4597);
nand U4662 (N_4662,N_4408,N_4495);
and U4663 (N_4663,N_4450,N_4463);
nand U4664 (N_4664,N_4427,N_4570);
xnor U4665 (N_4665,N_4521,N_4591);
or U4666 (N_4666,N_4512,N_4466);
or U4667 (N_4667,N_4528,N_4412);
and U4668 (N_4668,N_4449,N_4489);
or U4669 (N_4669,N_4517,N_4465);
or U4670 (N_4670,N_4581,N_4580);
or U4671 (N_4671,N_4518,N_4501);
or U4672 (N_4672,N_4468,N_4403);
nand U4673 (N_4673,N_4444,N_4409);
nand U4674 (N_4674,N_4490,N_4592);
and U4675 (N_4675,N_4446,N_4476);
and U4676 (N_4676,N_4441,N_4516);
and U4677 (N_4677,N_4457,N_4566);
nand U4678 (N_4678,N_4572,N_4453);
and U4679 (N_4679,N_4502,N_4400);
xor U4680 (N_4680,N_4402,N_4436);
and U4681 (N_4681,N_4440,N_4535);
nor U4682 (N_4682,N_4413,N_4422);
nor U4683 (N_4683,N_4445,N_4505);
xnor U4684 (N_4684,N_4443,N_4522);
nor U4685 (N_4685,N_4506,N_4530);
xor U4686 (N_4686,N_4548,N_4423);
nand U4687 (N_4687,N_4471,N_4576);
nand U4688 (N_4688,N_4556,N_4479);
nand U4689 (N_4689,N_4504,N_4559);
and U4690 (N_4690,N_4549,N_4513);
nor U4691 (N_4691,N_4547,N_4432);
xor U4692 (N_4692,N_4405,N_4520);
and U4693 (N_4693,N_4456,N_4472);
nand U4694 (N_4694,N_4493,N_4596);
and U4695 (N_4695,N_4564,N_4510);
nand U4696 (N_4696,N_4584,N_4487);
and U4697 (N_4697,N_4447,N_4420);
or U4698 (N_4698,N_4499,N_4551);
or U4699 (N_4699,N_4588,N_4536);
nand U4700 (N_4700,N_4580,N_4427);
and U4701 (N_4701,N_4432,N_4550);
or U4702 (N_4702,N_4486,N_4460);
xor U4703 (N_4703,N_4590,N_4501);
and U4704 (N_4704,N_4430,N_4576);
nor U4705 (N_4705,N_4467,N_4524);
nor U4706 (N_4706,N_4406,N_4548);
or U4707 (N_4707,N_4486,N_4532);
or U4708 (N_4708,N_4539,N_4412);
nand U4709 (N_4709,N_4406,N_4588);
nor U4710 (N_4710,N_4506,N_4572);
nand U4711 (N_4711,N_4596,N_4403);
xor U4712 (N_4712,N_4594,N_4560);
and U4713 (N_4713,N_4428,N_4479);
nand U4714 (N_4714,N_4411,N_4444);
nor U4715 (N_4715,N_4427,N_4452);
and U4716 (N_4716,N_4500,N_4595);
nor U4717 (N_4717,N_4476,N_4513);
xor U4718 (N_4718,N_4402,N_4458);
nor U4719 (N_4719,N_4488,N_4446);
and U4720 (N_4720,N_4520,N_4485);
nor U4721 (N_4721,N_4498,N_4486);
nand U4722 (N_4722,N_4474,N_4500);
and U4723 (N_4723,N_4533,N_4568);
and U4724 (N_4724,N_4534,N_4459);
nand U4725 (N_4725,N_4535,N_4455);
nand U4726 (N_4726,N_4545,N_4414);
xnor U4727 (N_4727,N_4439,N_4573);
nand U4728 (N_4728,N_4551,N_4466);
and U4729 (N_4729,N_4595,N_4593);
nand U4730 (N_4730,N_4566,N_4417);
nand U4731 (N_4731,N_4514,N_4581);
or U4732 (N_4732,N_4563,N_4407);
or U4733 (N_4733,N_4440,N_4403);
and U4734 (N_4734,N_4461,N_4522);
xor U4735 (N_4735,N_4416,N_4598);
xor U4736 (N_4736,N_4523,N_4426);
and U4737 (N_4737,N_4497,N_4524);
nand U4738 (N_4738,N_4557,N_4590);
nand U4739 (N_4739,N_4408,N_4508);
nor U4740 (N_4740,N_4462,N_4526);
and U4741 (N_4741,N_4439,N_4429);
and U4742 (N_4742,N_4526,N_4459);
nand U4743 (N_4743,N_4596,N_4513);
nand U4744 (N_4744,N_4414,N_4514);
xnor U4745 (N_4745,N_4589,N_4528);
nand U4746 (N_4746,N_4598,N_4576);
xor U4747 (N_4747,N_4410,N_4404);
xnor U4748 (N_4748,N_4493,N_4585);
or U4749 (N_4749,N_4473,N_4564);
nor U4750 (N_4750,N_4424,N_4534);
nor U4751 (N_4751,N_4480,N_4521);
nor U4752 (N_4752,N_4549,N_4402);
nand U4753 (N_4753,N_4537,N_4514);
xnor U4754 (N_4754,N_4430,N_4571);
and U4755 (N_4755,N_4453,N_4499);
or U4756 (N_4756,N_4541,N_4474);
and U4757 (N_4757,N_4454,N_4567);
or U4758 (N_4758,N_4538,N_4423);
or U4759 (N_4759,N_4459,N_4583);
or U4760 (N_4760,N_4472,N_4410);
or U4761 (N_4761,N_4455,N_4559);
or U4762 (N_4762,N_4571,N_4599);
nand U4763 (N_4763,N_4519,N_4434);
nor U4764 (N_4764,N_4492,N_4432);
nor U4765 (N_4765,N_4556,N_4406);
nand U4766 (N_4766,N_4503,N_4472);
nor U4767 (N_4767,N_4415,N_4486);
and U4768 (N_4768,N_4460,N_4492);
xnor U4769 (N_4769,N_4487,N_4592);
nand U4770 (N_4770,N_4587,N_4561);
or U4771 (N_4771,N_4567,N_4520);
nor U4772 (N_4772,N_4496,N_4441);
xor U4773 (N_4773,N_4477,N_4596);
or U4774 (N_4774,N_4508,N_4527);
nand U4775 (N_4775,N_4543,N_4406);
nor U4776 (N_4776,N_4511,N_4536);
and U4777 (N_4777,N_4408,N_4558);
nand U4778 (N_4778,N_4443,N_4563);
nand U4779 (N_4779,N_4491,N_4540);
and U4780 (N_4780,N_4471,N_4414);
nand U4781 (N_4781,N_4555,N_4488);
nor U4782 (N_4782,N_4411,N_4537);
and U4783 (N_4783,N_4500,N_4567);
xnor U4784 (N_4784,N_4470,N_4538);
and U4785 (N_4785,N_4502,N_4462);
xnor U4786 (N_4786,N_4442,N_4464);
and U4787 (N_4787,N_4459,N_4404);
and U4788 (N_4788,N_4561,N_4466);
xnor U4789 (N_4789,N_4562,N_4597);
nor U4790 (N_4790,N_4453,N_4546);
and U4791 (N_4791,N_4454,N_4588);
nand U4792 (N_4792,N_4469,N_4588);
xor U4793 (N_4793,N_4514,N_4589);
and U4794 (N_4794,N_4531,N_4460);
nor U4795 (N_4795,N_4408,N_4434);
or U4796 (N_4796,N_4570,N_4551);
xnor U4797 (N_4797,N_4583,N_4434);
and U4798 (N_4798,N_4407,N_4595);
and U4799 (N_4799,N_4453,N_4589);
nor U4800 (N_4800,N_4702,N_4782);
nor U4801 (N_4801,N_4681,N_4713);
or U4802 (N_4802,N_4679,N_4611);
and U4803 (N_4803,N_4755,N_4762);
or U4804 (N_4804,N_4682,N_4663);
and U4805 (N_4805,N_4699,N_4780);
xnor U4806 (N_4806,N_4658,N_4622);
or U4807 (N_4807,N_4676,N_4778);
xor U4808 (N_4808,N_4765,N_4756);
nand U4809 (N_4809,N_4701,N_4612);
or U4810 (N_4810,N_4752,N_4725);
or U4811 (N_4811,N_4609,N_4601);
or U4812 (N_4812,N_4630,N_4645);
and U4813 (N_4813,N_4749,N_4721);
and U4814 (N_4814,N_4792,N_4600);
nor U4815 (N_4815,N_4641,N_4714);
nand U4816 (N_4816,N_4656,N_4728);
nor U4817 (N_4817,N_4718,N_4649);
or U4818 (N_4818,N_4716,N_4690);
and U4819 (N_4819,N_4693,N_4621);
or U4820 (N_4820,N_4674,N_4614);
or U4821 (N_4821,N_4795,N_4738);
nor U4822 (N_4822,N_4736,N_4624);
and U4823 (N_4823,N_4683,N_4769);
nor U4824 (N_4824,N_4720,N_4618);
or U4825 (N_4825,N_4710,N_4760);
nor U4826 (N_4826,N_4629,N_4766);
and U4827 (N_4827,N_4711,N_4633);
and U4828 (N_4828,N_4632,N_4745);
xnor U4829 (N_4829,N_4647,N_4610);
nand U4830 (N_4830,N_4793,N_4734);
xnor U4831 (N_4831,N_4664,N_4653);
nand U4832 (N_4832,N_4626,N_4746);
nor U4833 (N_4833,N_4668,N_4726);
or U4834 (N_4834,N_4787,N_4636);
xor U4835 (N_4835,N_4731,N_4770);
or U4836 (N_4836,N_4730,N_4703);
or U4837 (N_4837,N_4779,N_4771);
and U4838 (N_4838,N_4659,N_4747);
or U4839 (N_4839,N_4741,N_4735);
nand U4840 (N_4840,N_4724,N_4648);
and U4841 (N_4841,N_4605,N_4774);
nor U4842 (N_4842,N_4739,N_4619);
nand U4843 (N_4843,N_4796,N_4744);
nand U4844 (N_4844,N_4603,N_4661);
nand U4845 (N_4845,N_4785,N_4788);
and U4846 (N_4846,N_4727,N_4764);
xnor U4847 (N_4847,N_4650,N_4617);
or U4848 (N_4848,N_4705,N_4722);
nor U4849 (N_4849,N_4662,N_4783);
nand U4850 (N_4850,N_4737,N_4775);
nand U4851 (N_4851,N_4784,N_4761);
xnor U4852 (N_4852,N_4640,N_4798);
or U4853 (N_4853,N_4794,N_4673);
xor U4854 (N_4854,N_4763,N_4773);
and U4855 (N_4855,N_4672,N_4628);
nor U4856 (N_4856,N_4695,N_4768);
and U4857 (N_4857,N_4712,N_4602);
and U4858 (N_4858,N_4657,N_4689);
nor U4859 (N_4859,N_4753,N_4651);
and U4860 (N_4860,N_4772,N_4607);
nor U4861 (N_4861,N_4743,N_4789);
and U4862 (N_4862,N_4758,N_4709);
and U4863 (N_4863,N_4750,N_4667);
or U4864 (N_4864,N_4706,N_4684);
nand U4865 (N_4865,N_4687,N_4697);
xor U4866 (N_4866,N_4688,N_4615);
and U4867 (N_4867,N_4694,N_4678);
or U4868 (N_4868,N_4767,N_4644);
and U4869 (N_4869,N_4665,N_4719);
nand U4870 (N_4870,N_4627,N_4740);
xnor U4871 (N_4871,N_4691,N_4613);
nand U4872 (N_4872,N_4637,N_4616);
nor U4873 (N_4873,N_4666,N_4733);
xnor U4874 (N_4874,N_4634,N_4692);
or U4875 (N_4875,N_4604,N_4655);
or U4876 (N_4876,N_4620,N_4677);
and U4877 (N_4877,N_4707,N_4700);
nor U4878 (N_4878,N_4638,N_4786);
xor U4879 (N_4879,N_4751,N_4723);
nand U4880 (N_4880,N_4708,N_4623);
nor U4881 (N_4881,N_4654,N_4606);
nor U4882 (N_4882,N_4631,N_4670);
xnor U4883 (N_4883,N_4642,N_4639);
and U4884 (N_4884,N_4732,N_4686);
or U4885 (N_4885,N_4680,N_4669);
and U4886 (N_4886,N_4790,N_4675);
nor U4887 (N_4887,N_4759,N_4643);
and U4888 (N_4888,N_4625,N_4777);
nand U4889 (N_4889,N_4742,N_4696);
xor U4890 (N_4890,N_4704,N_4791);
or U4891 (N_4891,N_4748,N_4646);
xor U4892 (N_4892,N_4608,N_4729);
and U4893 (N_4893,N_4797,N_4671);
and U4894 (N_4894,N_4660,N_4685);
and U4895 (N_4895,N_4754,N_4635);
and U4896 (N_4896,N_4781,N_4757);
xor U4897 (N_4897,N_4776,N_4715);
and U4898 (N_4898,N_4799,N_4698);
nor U4899 (N_4899,N_4717,N_4652);
nand U4900 (N_4900,N_4794,N_4677);
and U4901 (N_4901,N_4719,N_4603);
and U4902 (N_4902,N_4791,N_4672);
or U4903 (N_4903,N_4796,N_4699);
nor U4904 (N_4904,N_4720,N_4668);
nor U4905 (N_4905,N_4648,N_4686);
nand U4906 (N_4906,N_4780,N_4799);
and U4907 (N_4907,N_4737,N_4699);
nand U4908 (N_4908,N_4786,N_4685);
xnor U4909 (N_4909,N_4760,N_4713);
nor U4910 (N_4910,N_4652,N_4734);
and U4911 (N_4911,N_4694,N_4748);
nand U4912 (N_4912,N_4797,N_4663);
nand U4913 (N_4913,N_4733,N_4704);
nand U4914 (N_4914,N_4704,N_4660);
xor U4915 (N_4915,N_4683,N_4665);
nand U4916 (N_4916,N_4665,N_4716);
nand U4917 (N_4917,N_4657,N_4730);
nand U4918 (N_4918,N_4774,N_4729);
nor U4919 (N_4919,N_4787,N_4649);
nor U4920 (N_4920,N_4797,N_4677);
and U4921 (N_4921,N_4666,N_4773);
nand U4922 (N_4922,N_4608,N_4752);
xnor U4923 (N_4923,N_4703,N_4603);
and U4924 (N_4924,N_4762,N_4723);
nor U4925 (N_4925,N_4783,N_4715);
nor U4926 (N_4926,N_4674,N_4629);
nor U4927 (N_4927,N_4620,N_4660);
nand U4928 (N_4928,N_4701,N_4710);
nor U4929 (N_4929,N_4738,N_4630);
nand U4930 (N_4930,N_4657,N_4604);
nand U4931 (N_4931,N_4794,N_4636);
nor U4932 (N_4932,N_4713,N_4791);
nor U4933 (N_4933,N_4790,N_4691);
nor U4934 (N_4934,N_4605,N_4653);
nand U4935 (N_4935,N_4694,N_4615);
or U4936 (N_4936,N_4796,N_4727);
xnor U4937 (N_4937,N_4790,N_4638);
nand U4938 (N_4938,N_4727,N_4671);
nand U4939 (N_4939,N_4609,N_4627);
or U4940 (N_4940,N_4625,N_4629);
and U4941 (N_4941,N_4755,N_4676);
and U4942 (N_4942,N_4623,N_4713);
nor U4943 (N_4943,N_4631,N_4780);
nor U4944 (N_4944,N_4679,N_4781);
nand U4945 (N_4945,N_4788,N_4721);
nand U4946 (N_4946,N_4709,N_4779);
nor U4947 (N_4947,N_4764,N_4769);
nor U4948 (N_4948,N_4631,N_4714);
nor U4949 (N_4949,N_4656,N_4729);
nand U4950 (N_4950,N_4762,N_4630);
or U4951 (N_4951,N_4759,N_4765);
or U4952 (N_4952,N_4731,N_4703);
nor U4953 (N_4953,N_4752,N_4706);
nor U4954 (N_4954,N_4671,N_4755);
or U4955 (N_4955,N_4634,N_4633);
nor U4956 (N_4956,N_4750,N_4748);
or U4957 (N_4957,N_4612,N_4640);
xnor U4958 (N_4958,N_4664,N_4651);
nor U4959 (N_4959,N_4670,N_4764);
and U4960 (N_4960,N_4690,N_4661);
nor U4961 (N_4961,N_4756,N_4727);
nand U4962 (N_4962,N_4686,N_4751);
or U4963 (N_4963,N_4638,N_4754);
nand U4964 (N_4964,N_4754,N_4748);
nand U4965 (N_4965,N_4671,N_4621);
nand U4966 (N_4966,N_4669,N_4799);
xor U4967 (N_4967,N_4682,N_4680);
nor U4968 (N_4968,N_4720,N_4691);
nor U4969 (N_4969,N_4614,N_4766);
and U4970 (N_4970,N_4793,N_4744);
nor U4971 (N_4971,N_4790,N_4795);
xnor U4972 (N_4972,N_4618,N_4604);
nand U4973 (N_4973,N_4707,N_4667);
and U4974 (N_4974,N_4653,N_4686);
and U4975 (N_4975,N_4667,N_4702);
and U4976 (N_4976,N_4696,N_4665);
nor U4977 (N_4977,N_4742,N_4730);
nand U4978 (N_4978,N_4766,N_4723);
xor U4979 (N_4979,N_4725,N_4628);
and U4980 (N_4980,N_4672,N_4600);
or U4981 (N_4981,N_4659,N_4685);
and U4982 (N_4982,N_4743,N_4703);
nand U4983 (N_4983,N_4794,N_4792);
and U4984 (N_4984,N_4711,N_4706);
and U4985 (N_4985,N_4746,N_4643);
or U4986 (N_4986,N_4795,N_4707);
xnor U4987 (N_4987,N_4647,N_4602);
nor U4988 (N_4988,N_4669,N_4653);
nor U4989 (N_4989,N_4647,N_4768);
or U4990 (N_4990,N_4674,N_4736);
nor U4991 (N_4991,N_4707,N_4617);
xnor U4992 (N_4992,N_4755,N_4642);
nand U4993 (N_4993,N_4618,N_4747);
nand U4994 (N_4994,N_4789,N_4783);
nor U4995 (N_4995,N_4639,N_4733);
and U4996 (N_4996,N_4755,N_4626);
and U4997 (N_4997,N_4685,N_4652);
or U4998 (N_4998,N_4760,N_4700);
nand U4999 (N_4999,N_4632,N_4778);
or UO_0 (O_0,N_4868,N_4929);
nand UO_1 (O_1,N_4841,N_4931);
nor UO_2 (O_2,N_4821,N_4921);
nor UO_3 (O_3,N_4934,N_4919);
or UO_4 (O_4,N_4851,N_4988);
nor UO_5 (O_5,N_4888,N_4806);
or UO_6 (O_6,N_4886,N_4999);
xor UO_7 (O_7,N_4915,N_4913);
nand UO_8 (O_8,N_4838,N_4980);
xor UO_9 (O_9,N_4803,N_4866);
xor UO_10 (O_10,N_4958,N_4849);
nand UO_11 (O_11,N_4860,N_4940);
and UO_12 (O_12,N_4847,N_4876);
nand UO_13 (O_13,N_4908,N_4971);
and UO_14 (O_14,N_4943,N_4948);
nor UO_15 (O_15,N_4974,N_4998);
or UO_16 (O_16,N_4989,N_4852);
and UO_17 (O_17,N_4961,N_4896);
xnor UO_18 (O_18,N_4832,N_4899);
nand UO_19 (O_19,N_4882,N_4986);
nor UO_20 (O_20,N_4842,N_4939);
xor UO_21 (O_21,N_4885,N_4926);
nand UO_22 (O_22,N_4981,N_4825);
or UO_23 (O_23,N_4970,N_4815);
nor UO_24 (O_24,N_4905,N_4972);
nand UO_25 (O_25,N_4897,N_4912);
nor UO_26 (O_26,N_4904,N_4973);
nor UO_27 (O_27,N_4992,N_4833);
nand UO_28 (O_28,N_4870,N_4834);
and UO_29 (O_29,N_4889,N_4829);
xor UO_30 (O_30,N_4867,N_4903);
xor UO_31 (O_31,N_4839,N_4865);
nor UO_32 (O_32,N_4922,N_4819);
and UO_33 (O_33,N_4898,N_4848);
or UO_34 (O_34,N_4923,N_4810);
nor UO_35 (O_35,N_4987,N_4859);
and UO_36 (O_36,N_4930,N_4954);
nor UO_37 (O_37,N_4862,N_4996);
or UO_38 (O_38,N_4968,N_4850);
and UO_39 (O_39,N_4846,N_4877);
or UO_40 (O_40,N_4966,N_4937);
or UO_41 (O_41,N_4950,N_4944);
xnor UO_42 (O_42,N_4936,N_4924);
nor UO_43 (O_43,N_4873,N_4802);
xor UO_44 (O_44,N_4854,N_4959);
xor UO_45 (O_45,N_4977,N_4836);
nand UO_46 (O_46,N_4979,N_4828);
nor UO_47 (O_47,N_4875,N_4813);
nor UO_48 (O_48,N_4946,N_4843);
xnor UO_49 (O_49,N_4880,N_4890);
nand UO_50 (O_50,N_4969,N_4891);
and UO_51 (O_51,N_4960,N_4932);
nor UO_52 (O_52,N_4938,N_4894);
and UO_53 (O_53,N_4893,N_4857);
and UO_54 (O_54,N_4800,N_4823);
xor UO_55 (O_55,N_4827,N_4984);
nand UO_56 (O_56,N_4812,N_4928);
xor UO_57 (O_57,N_4941,N_4820);
xor UO_58 (O_58,N_4900,N_4807);
or UO_59 (O_59,N_4945,N_4962);
nor UO_60 (O_60,N_4978,N_4955);
or UO_61 (O_61,N_4990,N_4952);
nand UO_62 (O_62,N_4814,N_4925);
xnor UO_63 (O_63,N_4895,N_4911);
xnor UO_64 (O_64,N_4957,N_4918);
and UO_65 (O_65,N_4864,N_4951);
nand UO_66 (O_66,N_4887,N_4909);
nand UO_67 (O_67,N_4965,N_4976);
nand UO_68 (O_68,N_4914,N_4995);
or UO_69 (O_69,N_4872,N_4845);
nor UO_70 (O_70,N_4910,N_4871);
and UO_71 (O_71,N_4964,N_4855);
or UO_72 (O_72,N_4826,N_4963);
nand UO_73 (O_73,N_4982,N_4874);
nor UO_74 (O_74,N_4835,N_4861);
or UO_75 (O_75,N_4869,N_4837);
and UO_76 (O_76,N_4902,N_4975);
and UO_77 (O_77,N_4991,N_4892);
nand UO_78 (O_78,N_4906,N_4994);
nor UO_79 (O_79,N_4808,N_4879);
or UO_80 (O_80,N_4884,N_4844);
or UO_81 (O_81,N_4901,N_4818);
nor UO_82 (O_82,N_4878,N_4927);
xor UO_83 (O_83,N_4947,N_4997);
and UO_84 (O_84,N_4863,N_4858);
or UO_85 (O_85,N_4916,N_4953);
xnor UO_86 (O_86,N_4831,N_4816);
and UO_87 (O_87,N_4993,N_4809);
and UO_88 (O_88,N_4805,N_4804);
xnor UO_89 (O_89,N_4853,N_4933);
and UO_90 (O_90,N_4856,N_4983);
nor UO_91 (O_91,N_4920,N_4907);
nor UO_92 (O_92,N_4840,N_4949);
xor UO_93 (O_93,N_4942,N_4881);
xnor UO_94 (O_94,N_4917,N_4935);
or UO_95 (O_95,N_4817,N_4822);
or UO_96 (O_96,N_4830,N_4801);
or UO_97 (O_97,N_4985,N_4883);
or UO_98 (O_98,N_4824,N_4811);
nor UO_99 (O_99,N_4956,N_4967);
nor UO_100 (O_100,N_4811,N_4951);
and UO_101 (O_101,N_4837,N_4890);
or UO_102 (O_102,N_4834,N_4802);
nor UO_103 (O_103,N_4941,N_4922);
or UO_104 (O_104,N_4984,N_4978);
xnor UO_105 (O_105,N_4992,N_4812);
nor UO_106 (O_106,N_4876,N_4849);
nand UO_107 (O_107,N_4997,N_4852);
or UO_108 (O_108,N_4840,N_4894);
xor UO_109 (O_109,N_4995,N_4990);
nor UO_110 (O_110,N_4920,N_4913);
nand UO_111 (O_111,N_4809,N_4930);
xor UO_112 (O_112,N_4907,N_4860);
nand UO_113 (O_113,N_4859,N_4963);
and UO_114 (O_114,N_4878,N_4946);
and UO_115 (O_115,N_4819,N_4951);
and UO_116 (O_116,N_4899,N_4834);
and UO_117 (O_117,N_4897,N_4948);
or UO_118 (O_118,N_4964,N_4956);
or UO_119 (O_119,N_4876,N_4963);
or UO_120 (O_120,N_4888,N_4900);
or UO_121 (O_121,N_4935,N_4948);
nor UO_122 (O_122,N_4849,N_4866);
xor UO_123 (O_123,N_4934,N_4950);
nor UO_124 (O_124,N_4839,N_4912);
nand UO_125 (O_125,N_4921,N_4977);
or UO_126 (O_126,N_4825,N_4827);
nor UO_127 (O_127,N_4834,N_4903);
nor UO_128 (O_128,N_4857,N_4974);
nor UO_129 (O_129,N_4873,N_4819);
nand UO_130 (O_130,N_4834,N_4893);
or UO_131 (O_131,N_4887,N_4971);
and UO_132 (O_132,N_4842,N_4897);
or UO_133 (O_133,N_4983,N_4861);
nor UO_134 (O_134,N_4857,N_4988);
nand UO_135 (O_135,N_4837,N_4860);
and UO_136 (O_136,N_4817,N_4870);
nand UO_137 (O_137,N_4885,N_4934);
nor UO_138 (O_138,N_4915,N_4922);
xnor UO_139 (O_139,N_4891,N_4992);
or UO_140 (O_140,N_4921,N_4919);
nor UO_141 (O_141,N_4971,N_4842);
nor UO_142 (O_142,N_4821,N_4816);
xnor UO_143 (O_143,N_4925,N_4831);
nor UO_144 (O_144,N_4957,N_4962);
xor UO_145 (O_145,N_4908,N_4919);
nor UO_146 (O_146,N_4917,N_4959);
nand UO_147 (O_147,N_4959,N_4826);
xor UO_148 (O_148,N_4851,N_4999);
nor UO_149 (O_149,N_4974,N_4964);
or UO_150 (O_150,N_4948,N_4870);
nand UO_151 (O_151,N_4882,N_4951);
or UO_152 (O_152,N_4852,N_4958);
xnor UO_153 (O_153,N_4966,N_4969);
and UO_154 (O_154,N_4801,N_4951);
and UO_155 (O_155,N_4903,N_4950);
nand UO_156 (O_156,N_4989,N_4863);
or UO_157 (O_157,N_4901,N_4983);
or UO_158 (O_158,N_4852,N_4977);
and UO_159 (O_159,N_4858,N_4902);
nor UO_160 (O_160,N_4953,N_4826);
or UO_161 (O_161,N_4862,N_4829);
or UO_162 (O_162,N_4870,N_4859);
and UO_163 (O_163,N_4998,N_4916);
nor UO_164 (O_164,N_4945,N_4851);
and UO_165 (O_165,N_4840,N_4878);
and UO_166 (O_166,N_4925,N_4930);
and UO_167 (O_167,N_4921,N_4972);
xnor UO_168 (O_168,N_4916,N_4928);
or UO_169 (O_169,N_4977,N_4989);
or UO_170 (O_170,N_4981,N_4845);
and UO_171 (O_171,N_4903,N_4947);
nor UO_172 (O_172,N_4901,N_4841);
nor UO_173 (O_173,N_4811,N_4948);
and UO_174 (O_174,N_4812,N_4976);
nor UO_175 (O_175,N_4896,N_4930);
xor UO_176 (O_176,N_4855,N_4983);
xor UO_177 (O_177,N_4961,N_4898);
nor UO_178 (O_178,N_4942,N_4841);
or UO_179 (O_179,N_4878,N_4819);
xnor UO_180 (O_180,N_4912,N_4883);
xnor UO_181 (O_181,N_4982,N_4856);
or UO_182 (O_182,N_4902,N_4929);
xnor UO_183 (O_183,N_4923,N_4880);
xnor UO_184 (O_184,N_4957,N_4960);
nand UO_185 (O_185,N_4986,N_4969);
and UO_186 (O_186,N_4821,N_4867);
nor UO_187 (O_187,N_4986,N_4955);
nand UO_188 (O_188,N_4850,N_4893);
nor UO_189 (O_189,N_4934,N_4958);
xnor UO_190 (O_190,N_4942,N_4983);
nand UO_191 (O_191,N_4821,N_4917);
nor UO_192 (O_192,N_4861,N_4955);
nor UO_193 (O_193,N_4859,N_4877);
or UO_194 (O_194,N_4951,N_4820);
and UO_195 (O_195,N_4947,N_4940);
and UO_196 (O_196,N_4938,N_4923);
or UO_197 (O_197,N_4957,N_4971);
xnor UO_198 (O_198,N_4808,N_4981);
and UO_199 (O_199,N_4813,N_4961);
xor UO_200 (O_200,N_4950,N_4925);
xor UO_201 (O_201,N_4927,N_4954);
nand UO_202 (O_202,N_4868,N_4967);
or UO_203 (O_203,N_4993,N_4905);
nand UO_204 (O_204,N_4839,N_4881);
xnor UO_205 (O_205,N_4936,N_4888);
xor UO_206 (O_206,N_4969,N_4932);
nor UO_207 (O_207,N_4860,N_4878);
and UO_208 (O_208,N_4879,N_4904);
or UO_209 (O_209,N_4873,N_4864);
or UO_210 (O_210,N_4985,N_4850);
nor UO_211 (O_211,N_4840,N_4870);
nor UO_212 (O_212,N_4933,N_4875);
and UO_213 (O_213,N_4905,N_4987);
nand UO_214 (O_214,N_4924,N_4928);
or UO_215 (O_215,N_4929,N_4811);
nor UO_216 (O_216,N_4935,N_4980);
xor UO_217 (O_217,N_4851,N_4869);
xor UO_218 (O_218,N_4979,N_4827);
or UO_219 (O_219,N_4931,N_4969);
nor UO_220 (O_220,N_4996,N_4871);
xnor UO_221 (O_221,N_4825,N_4978);
nor UO_222 (O_222,N_4817,N_4994);
nand UO_223 (O_223,N_4987,N_4895);
xor UO_224 (O_224,N_4855,N_4912);
and UO_225 (O_225,N_4922,N_4901);
xnor UO_226 (O_226,N_4947,N_4877);
xor UO_227 (O_227,N_4812,N_4866);
or UO_228 (O_228,N_4844,N_4865);
nand UO_229 (O_229,N_4902,N_4953);
nor UO_230 (O_230,N_4950,N_4835);
nand UO_231 (O_231,N_4807,N_4991);
nand UO_232 (O_232,N_4884,N_4974);
nand UO_233 (O_233,N_4905,N_4876);
or UO_234 (O_234,N_4822,N_4876);
nand UO_235 (O_235,N_4804,N_4875);
nor UO_236 (O_236,N_4877,N_4882);
xor UO_237 (O_237,N_4978,N_4973);
nand UO_238 (O_238,N_4999,N_4823);
or UO_239 (O_239,N_4838,N_4985);
and UO_240 (O_240,N_4948,N_4838);
xor UO_241 (O_241,N_4973,N_4923);
xor UO_242 (O_242,N_4867,N_4854);
nand UO_243 (O_243,N_4911,N_4883);
nand UO_244 (O_244,N_4983,N_4833);
nor UO_245 (O_245,N_4927,N_4888);
xnor UO_246 (O_246,N_4961,N_4911);
and UO_247 (O_247,N_4985,N_4901);
and UO_248 (O_248,N_4975,N_4887);
or UO_249 (O_249,N_4884,N_4865);
xor UO_250 (O_250,N_4950,N_4997);
nand UO_251 (O_251,N_4919,N_4914);
nor UO_252 (O_252,N_4894,N_4846);
nand UO_253 (O_253,N_4931,N_4983);
nand UO_254 (O_254,N_4876,N_4820);
xnor UO_255 (O_255,N_4921,N_4956);
and UO_256 (O_256,N_4830,N_4992);
xnor UO_257 (O_257,N_4926,N_4942);
xor UO_258 (O_258,N_4975,N_4906);
and UO_259 (O_259,N_4834,N_4808);
and UO_260 (O_260,N_4850,N_4904);
or UO_261 (O_261,N_4844,N_4820);
nand UO_262 (O_262,N_4822,N_4980);
and UO_263 (O_263,N_4925,N_4901);
nor UO_264 (O_264,N_4873,N_4910);
nor UO_265 (O_265,N_4845,N_4906);
nor UO_266 (O_266,N_4931,N_4835);
nor UO_267 (O_267,N_4971,N_4841);
or UO_268 (O_268,N_4818,N_4871);
nor UO_269 (O_269,N_4893,N_4931);
xor UO_270 (O_270,N_4950,N_4824);
or UO_271 (O_271,N_4804,N_4891);
and UO_272 (O_272,N_4854,N_4887);
and UO_273 (O_273,N_4812,N_4966);
and UO_274 (O_274,N_4999,N_4970);
nand UO_275 (O_275,N_4912,N_4852);
xnor UO_276 (O_276,N_4999,N_4930);
or UO_277 (O_277,N_4805,N_4832);
nand UO_278 (O_278,N_4933,N_4869);
and UO_279 (O_279,N_4812,N_4872);
and UO_280 (O_280,N_4845,N_4822);
and UO_281 (O_281,N_4905,N_4844);
xor UO_282 (O_282,N_4909,N_4852);
or UO_283 (O_283,N_4920,N_4835);
and UO_284 (O_284,N_4978,N_4931);
or UO_285 (O_285,N_4921,N_4922);
or UO_286 (O_286,N_4945,N_4866);
and UO_287 (O_287,N_4996,N_4958);
or UO_288 (O_288,N_4818,N_4949);
xnor UO_289 (O_289,N_4968,N_4808);
xnor UO_290 (O_290,N_4991,N_4917);
xnor UO_291 (O_291,N_4958,N_4951);
xor UO_292 (O_292,N_4963,N_4824);
and UO_293 (O_293,N_4822,N_4804);
and UO_294 (O_294,N_4884,N_4979);
xor UO_295 (O_295,N_4853,N_4929);
xor UO_296 (O_296,N_4928,N_4811);
xor UO_297 (O_297,N_4858,N_4929);
nand UO_298 (O_298,N_4858,N_4889);
nand UO_299 (O_299,N_4916,N_4942);
nand UO_300 (O_300,N_4974,N_4802);
xor UO_301 (O_301,N_4871,N_4906);
nand UO_302 (O_302,N_4821,N_4965);
nand UO_303 (O_303,N_4980,N_4862);
or UO_304 (O_304,N_4969,N_4892);
nand UO_305 (O_305,N_4954,N_4952);
nor UO_306 (O_306,N_4985,N_4886);
or UO_307 (O_307,N_4880,N_4968);
nor UO_308 (O_308,N_4804,N_4874);
and UO_309 (O_309,N_4915,N_4808);
nand UO_310 (O_310,N_4874,N_4999);
nor UO_311 (O_311,N_4823,N_4835);
xor UO_312 (O_312,N_4827,N_4843);
and UO_313 (O_313,N_4945,N_4838);
xnor UO_314 (O_314,N_4914,N_4825);
and UO_315 (O_315,N_4973,N_4994);
and UO_316 (O_316,N_4971,N_4922);
or UO_317 (O_317,N_4849,N_4957);
nand UO_318 (O_318,N_4804,N_4867);
nand UO_319 (O_319,N_4880,N_4892);
or UO_320 (O_320,N_4882,N_4866);
or UO_321 (O_321,N_4959,N_4820);
xnor UO_322 (O_322,N_4993,N_4983);
nand UO_323 (O_323,N_4928,N_4974);
nand UO_324 (O_324,N_4904,N_4830);
and UO_325 (O_325,N_4861,N_4840);
or UO_326 (O_326,N_4815,N_4802);
nor UO_327 (O_327,N_4806,N_4862);
and UO_328 (O_328,N_4942,N_4993);
xor UO_329 (O_329,N_4922,N_4838);
xnor UO_330 (O_330,N_4878,N_4991);
xnor UO_331 (O_331,N_4951,N_4912);
and UO_332 (O_332,N_4833,N_4896);
nor UO_333 (O_333,N_4946,N_4976);
xnor UO_334 (O_334,N_4824,N_4880);
nand UO_335 (O_335,N_4891,N_4815);
xnor UO_336 (O_336,N_4848,N_4869);
xor UO_337 (O_337,N_4941,N_4845);
nor UO_338 (O_338,N_4933,N_4847);
xor UO_339 (O_339,N_4956,N_4962);
and UO_340 (O_340,N_4939,N_4809);
nand UO_341 (O_341,N_4984,N_4912);
xor UO_342 (O_342,N_4950,N_4899);
nand UO_343 (O_343,N_4902,N_4994);
nor UO_344 (O_344,N_4882,N_4980);
and UO_345 (O_345,N_4806,N_4936);
nor UO_346 (O_346,N_4917,N_4983);
xnor UO_347 (O_347,N_4903,N_4803);
and UO_348 (O_348,N_4946,N_4982);
and UO_349 (O_349,N_4823,N_4951);
or UO_350 (O_350,N_4848,N_4978);
or UO_351 (O_351,N_4974,N_4953);
or UO_352 (O_352,N_4923,N_4999);
and UO_353 (O_353,N_4819,N_4856);
nor UO_354 (O_354,N_4854,N_4875);
nor UO_355 (O_355,N_4825,N_4904);
nor UO_356 (O_356,N_4936,N_4825);
or UO_357 (O_357,N_4816,N_4818);
xor UO_358 (O_358,N_4957,N_4825);
xnor UO_359 (O_359,N_4909,N_4874);
nor UO_360 (O_360,N_4993,N_4839);
or UO_361 (O_361,N_4968,N_4829);
xor UO_362 (O_362,N_4974,N_4950);
or UO_363 (O_363,N_4828,N_4862);
xor UO_364 (O_364,N_4866,N_4838);
or UO_365 (O_365,N_4958,N_4944);
xnor UO_366 (O_366,N_4911,N_4807);
nor UO_367 (O_367,N_4990,N_4807);
nor UO_368 (O_368,N_4820,N_4990);
or UO_369 (O_369,N_4934,N_4916);
nor UO_370 (O_370,N_4805,N_4853);
or UO_371 (O_371,N_4924,N_4818);
nor UO_372 (O_372,N_4851,N_4977);
nor UO_373 (O_373,N_4848,N_4934);
and UO_374 (O_374,N_4821,N_4958);
nor UO_375 (O_375,N_4830,N_4964);
nor UO_376 (O_376,N_4953,N_4910);
or UO_377 (O_377,N_4964,N_4809);
nor UO_378 (O_378,N_4974,N_4989);
or UO_379 (O_379,N_4840,N_4924);
and UO_380 (O_380,N_4885,N_4804);
and UO_381 (O_381,N_4910,N_4900);
nand UO_382 (O_382,N_4808,N_4844);
xor UO_383 (O_383,N_4994,N_4835);
or UO_384 (O_384,N_4939,N_4847);
and UO_385 (O_385,N_4987,N_4921);
and UO_386 (O_386,N_4954,N_4856);
and UO_387 (O_387,N_4991,N_4986);
nand UO_388 (O_388,N_4885,N_4826);
and UO_389 (O_389,N_4804,N_4936);
nand UO_390 (O_390,N_4930,N_4980);
nand UO_391 (O_391,N_4929,N_4842);
nor UO_392 (O_392,N_4840,N_4810);
nor UO_393 (O_393,N_4832,N_4948);
xnor UO_394 (O_394,N_4859,N_4898);
nor UO_395 (O_395,N_4904,N_4878);
xor UO_396 (O_396,N_4986,N_4900);
nor UO_397 (O_397,N_4917,N_4825);
or UO_398 (O_398,N_4959,N_4962);
nand UO_399 (O_399,N_4819,N_4832);
nor UO_400 (O_400,N_4983,N_4905);
xor UO_401 (O_401,N_4807,N_4836);
and UO_402 (O_402,N_4850,N_4832);
xor UO_403 (O_403,N_4950,N_4937);
or UO_404 (O_404,N_4949,N_4908);
nand UO_405 (O_405,N_4889,N_4929);
or UO_406 (O_406,N_4841,N_4824);
nand UO_407 (O_407,N_4926,N_4869);
or UO_408 (O_408,N_4855,N_4925);
and UO_409 (O_409,N_4934,N_4807);
xnor UO_410 (O_410,N_4872,N_4871);
nand UO_411 (O_411,N_4982,N_4978);
nor UO_412 (O_412,N_4805,N_4848);
and UO_413 (O_413,N_4819,N_4881);
nor UO_414 (O_414,N_4877,N_4968);
xor UO_415 (O_415,N_4875,N_4900);
or UO_416 (O_416,N_4923,N_4910);
nand UO_417 (O_417,N_4904,N_4815);
nand UO_418 (O_418,N_4973,N_4872);
nor UO_419 (O_419,N_4844,N_4917);
and UO_420 (O_420,N_4803,N_4840);
and UO_421 (O_421,N_4956,N_4880);
nor UO_422 (O_422,N_4976,N_4986);
nor UO_423 (O_423,N_4900,N_4865);
or UO_424 (O_424,N_4809,N_4824);
nor UO_425 (O_425,N_4935,N_4854);
nand UO_426 (O_426,N_4818,N_4902);
nor UO_427 (O_427,N_4985,N_4820);
and UO_428 (O_428,N_4973,N_4835);
nand UO_429 (O_429,N_4881,N_4897);
nand UO_430 (O_430,N_4850,N_4880);
nand UO_431 (O_431,N_4894,N_4924);
nand UO_432 (O_432,N_4856,N_4934);
or UO_433 (O_433,N_4886,N_4820);
nor UO_434 (O_434,N_4834,N_4920);
and UO_435 (O_435,N_4861,N_4932);
nor UO_436 (O_436,N_4913,N_4840);
xnor UO_437 (O_437,N_4912,N_4825);
nand UO_438 (O_438,N_4951,N_4910);
nand UO_439 (O_439,N_4917,N_4961);
nor UO_440 (O_440,N_4857,N_4892);
nor UO_441 (O_441,N_4950,N_4989);
nor UO_442 (O_442,N_4808,N_4806);
nand UO_443 (O_443,N_4950,N_4820);
and UO_444 (O_444,N_4956,N_4871);
or UO_445 (O_445,N_4990,N_4827);
nor UO_446 (O_446,N_4895,N_4909);
or UO_447 (O_447,N_4944,N_4980);
or UO_448 (O_448,N_4989,N_4850);
or UO_449 (O_449,N_4923,N_4886);
nand UO_450 (O_450,N_4806,N_4954);
nand UO_451 (O_451,N_4928,N_4827);
nand UO_452 (O_452,N_4914,N_4927);
and UO_453 (O_453,N_4864,N_4949);
nor UO_454 (O_454,N_4870,N_4976);
nor UO_455 (O_455,N_4967,N_4908);
and UO_456 (O_456,N_4983,N_4928);
nand UO_457 (O_457,N_4940,N_4991);
and UO_458 (O_458,N_4825,N_4855);
nor UO_459 (O_459,N_4832,N_4919);
nor UO_460 (O_460,N_4946,N_4988);
and UO_461 (O_461,N_4837,N_4931);
or UO_462 (O_462,N_4933,N_4924);
and UO_463 (O_463,N_4849,N_4865);
nor UO_464 (O_464,N_4860,N_4921);
and UO_465 (O_465,N_4932,N_4887);
nor UO_466 (O_466,N_4885,N_4842);
xnor UO_467 (O_467,N_4876,N_4805);
or UO_468 (O_468,N_4916,N_4886);
and UO_469 (O_469,N_4967,N_4820);
or UO_470 (O_470,N_4855,N_4881);
xnor UO_471 (O_471,N_4845,N_4821);
or UO_472 (O_472,N_4850,N_4983);
or UO_473 (O_473,N_4962,N_4986);
and UO_474 (O_474,N_4893,N_4993);
and UO_475 (O_475,N_4985,N_4910);
and UO_476 (O_476,N_4811,N_4974);
or UO_477 (O_477,N_4820,N_4978);
or UO_478 (O_478,N_4888,N_4929);
or UO_479 (O_479,N_4842,N_4872);
and UO_480 (O_480,N_4919,N_4955);
nand UO_481 (O_481,N_4988,N_4969);
xnor UO_482 (O_482,N_4919,N_4822);
and UO_483 (O_483,N_4817,N_4876);
nand UO_484 (O_484,N_4986,N_4815);
nand UO_485 (O_485,N_4826,N_4857);
nand UO_486 (O_486,N_4869,N_4989);
nor UO_487 (O_487,N_4855,N_4973);
nand UO_488 (O_488,N_4945,N_4994);
and UO_489 (O_489,N_4937,N_4981);
or UO_490 (O_490,N_4980,N_4858);
and UO_491 (O_491,N_4886,N_4892);
or UO_492 (O_492,N_4802,N_4922);
and UO_493 (O_493,N_4835,N_4934);
or UO_494 (O_494,N_4921,N_4938);
xor UO_495 (O_495,N_4977,N_4831);
and UO_496 (O_496,N_4814,N_4976);
or UO_497 (O_497,N_4937,N_4847);
xnor UO_498 (O_498,N_4987,N_4996);
nor UO_499 (O_499,N_4963,N_4955);
and UO_500 (O_500,N_4841,N_4843);
nand UO_501 (O_501,N_4962,N_4874);
xnor UO_502 (O_502,N_4937,N_4831);
nor UO_503 (O_503,N_4938,N_4808);
and UO_504 (O_504,N_4987,N_4874);
or UO_505 (O_505,N_4959,N_4864);
nor UO_506 (O_506,N_4943,N_4934);
or UO_507 (O_507,N_4805,N_4887);
nand UO_508 (O_508,N_4972,N_4854);
nand UO_509 (O_509,N_4932,N_4970);
nand UO_510 (O_510,N_4915,N_4926);
and UO_511 (O_511,N_4988,N_4913);
xor UO_512 (O_512,N_4995,N_4814);
and UO_513 (O_513,N_4959,N_4830);
or UO_514 (O_514,N_4961,N_4849);
or UO_515 (O_515,N_4869,N_4971);
xnor UO_516 (O_516,N_4828,N_4962);
nor UO_517 (O_517,N_4998,N_4995);
xnor UO_518 (O_518,N_4879,N_4919);
nand UO_519 (O_519,N_4891,N_4800);
xnor UO_520 (O_520,N_4893,N_4943);
xnor UO_521 (O_521,N_4871,N_4882);
and UO_522 (O_522,N_4812,N_4886);
nand UO_523 (O_523,N_4996,N_4927);
xor UO_524 (O_524,N_4920,N_4846);
and UO_525 (O_525,N_4852,N_4875);
and UO_526 (O_526,N_4853,N_4813);
and UO_527 (O_527,N_4898,N_4943);
xnor UO_528 (O_528,N_4897,N_4978);
or UO_529 (O_529,N_4913,N_4967);
and UO_530 (O_530,N_4808,N_4858);
or UO_531 (O_531,N_4901,N_4889);
nand UO_532 (O_532,N_4969,N_4930);
xor UO_533 (O_533,N_4899,N_4901);
or UO_534 (O_534,N_4956,N_4920);
and UO_535 (O_535,N_4850,N_4915);
nor UO_536 (O_536,N_4805,N_4899);
xor UO_537 (O_537,N_4855,N_4888);
nand UO_538 (O_538,N_4808,N_4856);
nor UO_539 (O_539,N_4907,N_4802);
or UO_540 (O_540,N_4926,N_4920);
and UO_541 (O_541,N_4813,N_4974);
nand UO_542 (O_542,N_4917,N_4951);
and UO_543 (O_543,N_4810,N_4876);
and UO_544 (O_544,N_4944,N_4993);
nand UO_545 (O_545,N_4915,N_4963);
and UO_546 (O_546,N_4921,N_4960);
or UO_547 (O_547,N_4824,N_4842);
nor UO_548 (O_548,N_4883,N_4907);
nor UO_549 (O_549,N_4824,N_4866);
nor UO_550 (O_550,N_4879,N_4851);
nand UO_551 (O_551,N_4894,N_4880);
xor UO_552 (O_552,N_4887,N_4811);
nand UO_553 (O_553,N_4939,N_4811);
and UO_554 (O_554,N_4878,N_4919);
nor UO_555 (O_555,N_4976,N_4934);
nor UO_556 (O_556,N_4865,N_4984);
nand UO_557 (O_557,N_4945,N_4906);
nand UO_558 (O_558,N_4911,N_4842);
nand UO_559 (O_559,N_4879,N_4974);
and UO_560 (O_560,N_4995,N_4838);
nand UO_561 (O_561,N_4924,N_4874);
or UO_562 (O_562,N_4936,N_4929);
nor UO_563 (O_563,N_4814,N_4895);
nor UO_564 (O_564,N_4954,N_4912);
nand UO_565 (O_565,N_4944,N_4934);
or UO_566 (O_566,N_4808,N_4947);
nor UO_567 (O_567,N_4928,N_4884);
nor UO_568 (O_568,N_4843,N_4910);
nor UO_569 (O_569,N_4887,N_4878);
nor UO_570 (O_570,N_4995,N_4932);
or UO_571 (O_571,N_4876,N_4836);
nand UO_572 (O_572,N_4922,N_4809);
or UO_573 (O_573,N_4806,N_4907);
nor UO_574 (O_574,N_4916,N_4903);
or UO_575 (O_575,N_4923,N_4818);
and UO_576 (O_576,N_4810,N_4903);
or UO_577 (O_577,N_4941,N_4895);
nor UO_578 (O_578,N_4862,N_4976);
nor UO_579 (O_579,N_4808,N_4878);
xnor UO_580 (O_580,N_4953,N_4980);
or UO_581 (O_581,N_4956,N_4909);
xnor UO_582 (O_582,N_4993,N_4913);
and UO_583 (O_583,N_4832,N_4985);
nand UO_584 (O_584,N_4827,N_4858);
nand UO_585 (O_585,N_4824,N_4839);
xnor UO_586 (O_586,N_4813,N_4978);
nand UO_587 (O_587,N_4917,N_4956);
nand UO_588 (O_588,N_4841,N_4975);
xor UO_589 (O_589,N_4864,N_4903);
and UO_590 (O_590,N_4964,N_4932);
nor UO_591 (O_591,N_4987,N_4947);
nor UO_592 (O_592,N_4804,N_4807);
and UO_593 (O_593,N_4985,N_4924);
nand UO_594 (O_594,N_4935,N_4837);
xor UO_595 (O_595,N_4889,N_4807);
and UO_596 (O_596,N_4867,N_4801);
nand UO_597 (O_597,N_4950,N_4853);
and UO_598 (O_598,N_4836,N_4816);
xnor UO_599 (O_599,N_4984,N_4826);
or UO_600 (O_600,N_4920,N_4864);
or UO_601 (O_601,N_4885,N_4946);
and UO_602 (O_602,N_4999,N_4933);
or UO_603 (O_603,N_4905,N_4999);
and UO_604 (O_604,N_4861,N_4908);
and UO_605 (O_605,N_4821,N_4814);
or UO_606 (O_606,N_4962,N_4844);
nor UO_607 (O_607,N_4809,N_4841);
xnor UO_608 (O_608,N_4977,N_4902);
xnor UO_609 (O_609,N_4919,N_4985);
xnor UO_610 (O_610,N_4984,N_4942);
xor UO_611 (O_611,N_4893,N_4887);
xnor UO_612 (O_612,N_4832,N_4933);
nor UO_613 (O_613,N_4951,N_4841);
or UO_614 (O_614,N_4875,N_4817);
xnor UO_615 (O_615,N_4804,N_4815);
and UO_616 (O_616,N_4839,N_4990);
nor UO_617 (O_617,N_4890,N_4986);
nor UO_618 (O_618,N_4901,N_4897);
nand UO_619 (O_619,N_4833,N_4960);
nor UO_620 (O_620,N_4840,N_4821);
nor UO_621 (O_621,N_4926,N_4887);
and UO_622 (O_622,N_4979,N_4965);
nand UO_623 (O_623,N_4878,N_4854);
or UO_624 (O_624,N_4821,N_4879);
and UO_625 (O_625,N_4887,N_4939);
and UO_626 (O_626,N_4820,N_4875);
and UO_627 (O_627,N_4901,N_4932);
nor UO_628 (O_628,N_4815,N_4958);
xor UO_629 (O_629,N_4866,N_4881);
nor UO_630 (O_630,N_4981,N_4855);
and UO_631 (O_631,N_4852,N_4800);
xnor UO_632 (O_632,N_4879,N_4859);
xor UO_633 (O_633,N_4881,N_4851);
nand UO_634 (O_634,N_4903,N_4937);
xnor UO_635 (O_635,N_4942,N_4915);
nor UO_636 (O_636,N_4896,N_4922);
and UO_637 (O_637,N_4842,N_4959);
xnor UO_638 (O_638,N_4938,N_4840);
nand UO_639 (O_639,N_4841,N_4941);
nor UO_640 (O_640,N_4816,N_4891);
nand UO_641 (O_641,N_4880,N_4821);
and UO_642 (O_642,N_4935,N_4825);
and UO_643 (O_643,N_4849,N_4901);
nor UO_644 (O_644,N_4961,N_4812);
nor UO_645 (O_645,N_4816,N_4955);
nor UO_646 (O_646,N_4884,N_4836);
nand UO_647 (O_647,N_4993,N_4996);
nand UO_648 (O_648,N_4800,N_4838);
or UO_649 (O_649,N_4977,N_4992);
nand UO_650 (O_650,N_4856,N_4866);
and UO_651 (O_651,N_4869,N_4844);
nand UO_652 (O_652,N_4889,N_4824);
nand UO_653 (O_653,N_4802,N_4865);
xnor UO_654 (O_654,N_4880,N_4938);
xor UO_655 (O_655,N_4944,N_4854);
xor UO_656 (O_656,N_4911,N_4946);
or UO_657 (O_657,N_4853,N_4839);
or UO_658 (O_658,N_4961,N_4943);
xnor UO_659 (O_659,N_4820,N_4917);
nand UO_660 (O_660,N_4828,N_4815);
or UO_661 (O_661,N_4942,N_4939);
and UO_662 (O_662,N_4911,N_4897);
or UO_663 (O_663,N_4959,N_4900);
xnor UO_664 (O_664,N_4965,N_4811);
nand UO_665 (O_665,N_4812,N_4939);
nor UO_666 (O_666,N_4978,N_4950);
xor UO_667 (O_667,N_4813,N_4999);
nor UO_668 (O_668,N_4975,N_4916);
nand UO_669 (O_669,N_4876,N_4902);
nor UO_670 (O_670,N_4992,N_4845);
xnor UO_671 (O_671,N_4973,N_4965);
nor UO_672 (O_672,N_4996,N_4925);
and UO_673 (O_673,N_4818,N_4995);
xnor UO_674 (O_674,N_4861,N_4852);
and UO_675 (O_675,N_4878,N_4833);
and UO_676 (O_676,N_4939,N_4912);
or UO_677 (O_677,N_4826,N_4994);
and UO_678 (O_678,N_4826,N_4917);
and UO_679 (O_679,N_4830,N_4911);
xor UO_680 (O_680,N_4843,N_4963);
or UO_681 (O_681,N_4989,N_4924);
and UO_682 (O_682,N_4808,N_4907);
nand UO_683 (O_683,N_4865,N_4887);
and UO_684 (O_684,N_4960,N_4998);
xor UO_685 (O_685,N_4905,N_4871);
xor UO_686 (O_686,N_4860,N_4856);
and UO_687 (O_687,N_4932,N_4915);
or UO_688 (O_688,N_4811,N_4912);
nor UO_689 (O_689,N_4997,N_4888);
nand UO_690 (O_690,N_4852,N_4833);
nor UO_691 (O_691,N_4987,N_4870);
xnor UO_692 (O_692,N_4854,N_4846);
nor UO_693 (O_693,N_4858,N_4825);
nor UO_694 (O_694,N_4960,N_4867);
or UO_695 (O_695,N_4813,N_4971);
and UO_696 (O_696,N_4869,N_4923);
nor UO_697 (O_697,N_4988,N_4846);
or UO_698 (O_698,N_4999,N_4902);
or UO_699 (O_699,N_4940,N_4959);
xor UO_700 (O_700,N_4843,N_4995);
nor UO_701 (O_701,N_4951,N_4849);
or UO_702 (O_702,N_4840,N_4857);
nand UO_703 (O_703,N_4807,N_4971);
or UO_704 (O_704,N_4950,N_4851);
or UO_705 (O_705,N_4959,N_4812);
or UO_706 (O_706,N_4862,N_4971);
and UO_707 (O_707,N_4837,N_4891);
xor UO_708 (O_708,N_4881,N_4858);
xor UO_709 (O_709,N_4860,N_4869);
nor UO_710 (O_710,N_4859,N_4944);
and UO_711 (O_711,N_4911,N_4894);
nand UO_712 (O_712,N_4922,N_4912);
nor UO_713 (O_713,N_4830,N_4802);
or UO_714 (O_714,N_4811,N_4930);
or UO_715 (O_715,N_4987,N_4936);
nand UO_716 (O_716,N_4978,N_4993);
and UO_717 (O_717,N_4916,N_4855);
nand UO_718 (O_718,N_4910,N_4901);
nand UO_719 (O_719,N_4900,N_4961);
xor UO_720 (O_720,N_4818,N_4936);
nor UO_721 (O_721,N_4993,N_4952);
and UO_722 (O_722,N_4930,N_4859);
nor UO_723 (O_723,N_4973,N_4886);
xor UO_724 (O_724,N_4853,N_4966);
xor UO_725 (O_725,N_4894,N_4833);
and UO_726 (O_726,N_4917,N_4993);
xor UO_727 (O_727,N_4962,N_4890);
nor UO_728 (O_728,N_4957,N_4864);
xor UO_729 (O_729,N_4886,N_4860);
and UO_730 (O_730,N_4896,N_4981);
xor UO_731 (O_731,N_4826,N_4996);
nand UO_732 (O_732,N_4960,N_4827);
xor UO_733 (O_733,N_4950,N_4909);
nor UO_734 (O_734,N_4956,N_4994);
or UO_735 (O_735,N_4952,N_4995);
or UO_736 (O_736,N_4897,N_4955);
nand UO_737 (O_737,N_4919,N_4965);
xor UO_738 (O_738,N_4940,N_4877);
nand UO_739 (O_739,N_4945,N_4844);
nor UO_740 (O_740,N_4985,N_4898);
nand UO_741 (O_741,N_4857,N_4847);
and UO_742 (O_742,N_4881,N_4862);
or UO_743 (O_743,N_4800,N_4874);
nand UO_744 (O_744,N_4933,N_4804);
and UO_745 (O_745,N_4865,N_4853);
xnor UO_746 (O_746,N_4966,N_4940);
and UO_747 (O_747,N_4941,N_4929);
nor UO_748 (O_748,N_4945,N_4855);
nor UO_749 (O_749,N_4856,N_4922);
nand UO_750 (O_750,N_4978,N_4842);
and UO_751 (O_751,N_4837,N_4919);
nor UO_752 (O_752,N_4814,N_4954);
nand UO_753 (O_753,N_4984,N_4948);
or UO_754 (O_754,N_4939,N_4890);
nor UO_755 (O_755,N_4878,N_4814);
or UO_756 (O_756,N_4842,N_4889);
nand UO_757 (O_757,N_4925,N_4907);
and UO_758 (O_758,N_4810,N_4979);
and UO_759 (O_759,N_4831,N_4975);
or UO_760 (O_760,N_4896,N_4931);
nand UO_761 (O_761,N_4943,N_4834);
and UO_762 (O_762,N_4853,N_4993);
nand UO_763 (O_763,N_4882,N_4800);
or UO_764 (O_764,N_4848,N_4837);
xor UO_765 (O_765,N_4877,N_4890);
or UO_766 (O_766,N_4948,N_4880);
or UO_767 (O_767,N_4854,N_4917);
nor UO_768 (O_768,N_4951,N_4925);
or UO_769 (O_769,N_4950,N_4860);
nor UO_770 (O_770,N_4876,N_4894);
nor UO_771 (O_771,N_4801,N_4805);
nand UO_772 (O_772,N_4906,N_4816);
nand UO_773 (O_773,N_4917,N_4851);
nand UO_774 (O_774,N_4968,N_4862);
nor UO_775 (O_775,N_4963,N_4817);
nor UO_776 (O_776,N_4959,N_4868);
xor UO_777 (O_777,N_4933,N_4926);
nand UO_778 (O_778,N_4960,N_4877);
or UO_779 (O_779,N_4971,N_4925);
or UO_780 (O_780,N_4834,N_4845);
and UO_781 (O_781,N_4925,N_4862);
and UO_782 (O_782,N_4919,N_4854);
and UO_783 (O_783,N_4839,N_4891);
nand UO_784 (O_784,N_4921,N_4997);
nor UO_785 (O_785,N_4904,N_4874);
xor UO_786 (O_786,N_4964,N_4825);
nor UO_787 (O_787,N_4896,N_4821);
and UO_788 (O_788,N_4810,N_4975);
xor UO_789 (O_789,N_4871,N_4937);
nor UO_790 (O_790,N_4931,N_4981);
and UO_791 (O_791,N_4818,N_4845);
nand UO_792 (O_792,N_4919,N_4893);
nor UO_793 (O_793,N_4976,N_4919);
and UO_794 (O_794,N_4900,N_4804);
or UO_795 (O_795,N_4933,N_4971);
nor UO_796 (O_796,N_4851,N_4922);
and UO_797 (O_797,N_4832,N_4940);
xor UO_798 (O_798,N_4988,N_4982);
or UO_799 (O_799,N_4953,N_4820);
xor UO_800 (O_800,N_4994,N_4880);
xnor UO_801 (O_801,N_4899,N_4853);
and UO_802 (O_802,N_4953,N_4844);
nor UO_803 (O_803,N_4907,N_4908);
nor UO_804 (O_804,N_4821,N_4844);
nor UO_805 (O_805,N_4982,N_4800);
xor UO_806 (O_806,N_4974,N_4882);
nor UO_807 (O_807,N_4858,N_4843);
nor UO_808 (O_808,N_4969,N_4901);
nand UO_809 (O_809,N_4925,N_4827);
nand UO_810 (O_810,N_4954,N_4823);
and UO_811 (O_811,N_4870,N_4833);
xnor UO_812 (O_812,N_4972,N_4994);
or UO_813 (O_813,N_4808,N_4813);
nor UO_814 (O_814,N_4858,N_4840);
xnor UO_815 (O_815,N_4981,N_4946);
or UO_816 (O_816,N_4828,N_4855);
nand UO_817 (O_817,N_4961,N_4840);
nor UO_818 (O_818,N_4920,N_4900);
nor UO_819 (O_819,N_4951,N_4856);
xnor UO_820 (O_820,N_4967,N_4819);
xor UO_821 (O_821,N_4885,N_4819);
nand UO_822 (O_822,N_4835,N_4895);
xnor UO_823 (O_823,N_4910,N_4800);
and UO_824 (O_824,N_4869,N_4911);
and UO_825 (O_825,N_4889,N_4936);
or UO_826 (O_826,N_4807,N_4843);
and UO_827 (O_827,N_4800,N_4900);
nor UO_828 (O_828,N_4983,N_4838);
or UO_829 (O_829,N_4852,N_4840);
or UO_830 (O_830,N_4938,N_4847);
nor UO_831 (O_831,N_4862,N_4901);
and UO_832 (O_832,N_4859,N_4803);
nor UO_833 (O_833,N_4838,N_4992);
nor UO_834 (O_834,N_4886,N_4993);
xnor UO_835 (O_835,N_4977,N_4871);
nor UO_836 (O_836,N_4835,N_4919);
nor UO_837 (O_837,N_4977,N_4853);
and UO_838 (O_838,N_4943,N_4880);
xor UO_839 (O_839,N_4966,N_4912);
and UO_840 (O_840,N_4835,N_4921);
and UO_841 (O_841,N_4895,N_4810);
and UO_842 (O_842,N_4850,N_4963);
nor UO_843 (O_843,N_4804,N_4881);
nand UO_844 (O_844,N_4986,N_4998);
nand UO_845 (O_845,N_4983,N_4873);
xnor UO_846 (O_846,N_4943,N_4849);
or UO_847 (O_847,N_4885,N_4852);
or UO_848 (O_848,N_4949,N_4873);
nor UO_849 (O_849,N_4921,N_4999);
xnor UO_850 (O_850,N_4883,N_4940);
nand UO_851 (O_851,N_4871,N_4870);
nor UO_852 (O_852,N_4959,N_4980);
and UO_853 (O_853,N_4902,N_4932);
and UO_854 (O_854,N_4978,N_4866);
and UO_855 (O_855,N_4848,N_4836);
and UO_856 (O_856,N_4815,N_4988);
or UO_857 (O_857,N_4895,N_4886);
and UO_858 (O_858,N_4883,N_4869);
nand UO_859 (O_859,N_4818,N_4898);
nor UO_860 (O_860,N_4939,N_4808);
xor UO_861 (O_861,N_4802,N_4862);
nor UO_862 (O_862,N_4901,N_4870);
nand UO_863 (O_863,N_4970,N_4867);
nand UO_864 (O_864,N_4914,N_4969);
and UO_865 (O_865,N_4937,N_4842);
and UO_866 (O_866,N_4962,N_4976);
nor UO_867 (O_867,N_4849,N_4906);
or UO_868 (O_868,N_4923,N_4962);
or UO_869 (O_869,N_4989,N_4855);
and UO_870 (O_870,N_4993,N_4918);
or UO_871 (O_871,N_4987,N_4823);
xnor UO_872 (O_872,N_4827,N_4876);
xnor UO_873 (O_873,N_4857,N_4973);
and UO_874 (O_874,N_4878,N_4976);
nand UO_875 (O_875,N_4836,N_4911);
and UO_876 (O_876,N_4840,N_4847);
and UO_877 (O_877,N_4805,N_4817);
or UO_878 (O_878,N_4882,N_4907);
nor UO_879 (O_879,N_4825,N_4954);
xor UO_880 (O_880,N_4831,N_4830);
xor UO_881 (O_881,N_4814,N_4904);
xor UO_882 (O_882,N_4955,N_4825);
nor UO_883 (O_883,N_4859,N_4916);
xor UO_884 (O_884,N_4964,N_4811);
or UO_885 (O_885,N_4875,N_4948);
nor UO_886 (O_886,N_4907,N_4971);
and UO_887 (O_887,N_4911,N_4866);
nor UO_888 (O_888,N_4958,N_4928);
and UO_889 (O_889,N_4967,N_4917);
nand UO_890 (O_890,N_4819,N_4872);
and UO_891 (O_891,N_4877,N_4905);
or UO_892 (O_892,N_4968,N_4990);
nor UO_893 (O_893,N_4984,N_4864);
nand UO_894 (O_894,N_4942,N_4876);
nor UO_895 (O_895,N_4886,N_4868);
and UO_896 (O_896,N_4960,N_4819);
xor UO_897 (O_897,N_4837,N_4976);
xnor UO_898 (O_898,N_4857,N_4863);
nand UO_899 (O_899,N_4807,N_4841);
xnor UO_900 (O_900,N_4889,N_4981);
xor UO_901 (O_901,N_4950,N_4831);
xor UO_902 (O_902,N_4916,N_4960);
or UO_903 (O_903,N_4896,N_4880);
nand UO_904 (O_904,N_4863,N_4940);
nand UO_905 (O_905,N_4841,N_4818);
or UO_906 (O_906,N_4823,N_4819);
xnor UO_907 (O_907,N_4845,N_4900);
or UO_908 (O_908,N_4982,N_4880);
nand UO_909 (O_909,N_4845,N_4961);
or UO_910 (O_910,N_4806,N_4855);
nor UO_911 (O_911,N_4946,N_4820);
xor UO_912 (O_912,N_4885,N_4907);
and UO_913 (O_913,N_4815,N_4948);
xnor UO_914 (O_914,N_4961,N_4802);
or UO_915 (O_915,N_4877,N_4986);
xor UO_916 (O_916,N_4803,N_4969);
and UO_917 (O_917,N_4859,N_4970);
nand UO_918 (O_918,N_4937,N_4841);
and UO_919 (O_919,N_4807,N_4868);
or UO_920 (O_920,N_4805,N_4972);
nor UO_921 (O_921,N_4997,N_4996);
and UO_922 (O_922,N_4952,N_4809);
nor UO_923 (O_923,N_4809,N_4997);
or UO_924 (O_924,N_4884,N_4830);
and UO_925 (O_925,N_4885,N_4881);
and UO_926 (O_926,N_4944,N_4826);
xor UO_927 (O_927,N_4808,N_4934);
or UO_928 (O_928,N_4848,N_4880);
or UO_929 (O_929,N_4867,N_4897);
or UO_930 (O_930,N_4953,N_4927);
nor UO_931 (O_931,N_4836,N_4843);
nor UO_932 (O_932,N_4803,N_4825);
nor UO_933 (O_933,N_4963,N_4970);
or UO_934 (O_934,N_4950,N_4983);
or UO_935 (O_935,N_4808,N_4841);
or UO_936 (O_936,N_4840,N_4856);
or UO_937 (O_937,N_4914,N_4810);
nand UO_938 (O_938,N_4944,N_4820);
or UO_939 (O_939,N_4915,N_4805);
and UO_940 (O_940,N_4809,N_4878);
or UO_941 (O_941,N_4892,N_4938);
nor UO_942 (O_942,N_4882,N_4950);
nand UO_943 (O_943,N_4877,N_4848);
xnor UO_944 (O_944,N_4961,N_4819);
nor UO_945 (O_945,N_4998,N_4859);
or UO_946 (O_946,N_4971,N_4837);
or UO_947 (O_947,N_4809,N_4954);
xor UO_948 (O_948,N_4819,N_4896);
xor UO_949 (O_949,N_4969,N_4960);
xor UO_950 (O_950,N_4870,N_4949);
xnor UO_951 (O_951,N_4836,N_4874);
nand UO_952 (O_952,N_4870,N_4962);
xnor UO_953 (O_953,N_4935,N_4882);
nor UO_954 (O_954,N_4858,N_4850);
nor UO_955 (O_955,N_4878,N_4877);
nor UO_956 (O_956,N_4872,N_4817);
xnor UO_957 (O_957,N_4933,N_4803);
nor UO_958 (O_958,N_4922,N_4928);
nand UO_959 (O_959,N_4949,N_4930);
and UO_960 (O_960,N_4812,N_4894);
and UO_961 (O_961,N_4929,N_4908);
xnor UO_962 (O_962,N_4959,N_4957);
nor UO_963 (O_963,N_4939,N_4990);
or UO_964 (O_964,N_4873,N_4967);
nor UO_965 (O_965,N_4977,N_4804);
xor UO_966 (O_966,N_4976,N_4802);
or UO_967 (O_967,N_4959,N_4865);
nand UO_968 (O_968,N_4863,N_4903);
nor UO_969 (O_969,N_4927,N_4979);
or UO_970 (O_970,N_4863,N_4854);
or UO_971 (O_971,N_4993,N_4851);
xnor UO_972 (O_972,N_4820,N_4814);
nand UO_973 (O_973,N_4921,N_4955);
xnor UO_974 (O_974,N_4811,N_4845);
nand UO_975 (O_975,N_4871,N_4911);
or UO_976 (O_976,N_4908,N_4807);
xnor UO_977 (O_977,N_4954,N_4998);
xnor UO_978 (O_978,N_4896,N_4820);
and UO_979 (O_979,N_4977,N_4812);
xor UO_980 (O_980,N_4981,N_4909);
and UO_981 (O_981,N_4989,N_4904);
or UO_982 (O_982,N_4966,N_4880);
nor UO_983 (O_983,N_4826,N_4863);
xnor UO_984 (O_984,N_4858,N_4909);
or UO_985 (O_985,N_4914,N_4836);
or UO_986 (O_986,N_4994,N_4841);
nor UO_987 (O_987,N_4867,N_4832);
nand UO_988 (O_988,N_4825,N_4961);
xor UO_989 (O_989,N_4895,N_4853);
nand UO_990 (O_990,N_4832,N_4887);
or UO_991 (O_991,N_4845,N_4838);
nor UO_992 (O_992,N_4873,N_4932);
nor UO_993 (O_993,N_4855,N_4846);
nand UO_994 (O_994,N_4891,N_4805);
xnor UO_995 (O_995,N_4921,N_4981);
nor UO_996 (O_996,N_4866,N_4840);
xor UO_997 (O_997,N_4937,N_4826);
xor UO_998 (O_998,N_4856,N_4913);
and UO_999 (O_999,N_4848,N_4865);
endmodule